module basic_750_5000_1000_10_levels_5xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
and U0 (N_0,In_536,In_431);
nor U1 (N_1,In_231,In_144);
nand U2 (N_2,In_639,In_171);
or U3 (N_3,In_617,In_381);
and U4 (N_4,In_553,In_629);
and U5 (N_5,In_335,In_628);
xor U6 (N_6,In_296,In_519);
and U7 (N_7,In_138,In_408);
or U8 (N_8,In_413,In_581);
or U9 (N_9,In_475,In_569);
or U10 (N_10,In_0,In_507);
or U11 (N_11,In_266,In_331);
nor U12 (N_12,In_115,In_270);
and U13 (N_13,In_533,In_33);
and U14 (N_14,In_557,In_438);
nand U15 (N_15,In_31,In_717);
nand U16 (N_16,In_517,In_538);
nand U17 (N_17,In_703,In_540);
and U18 (N_18,In_73,In_55);
nand U19 (N_19,In_549,In_460);
or U20 (N_20,In_715,In_94);
nor U21 (N_21,In_72,In_30);
or U22 (N_22,In_319,In_136);
nor U23 (N_23,In_156,In_19);
and U24 (N_24,In_347,In_669);
or U25 (N_25,In_133,In_297);
nor U26 (N_26,In_423,In_178);
or U27 (N_27,In_678,In_742);
nand U28 (N_28,In_2,In_532);
xnor U29 (N_29,In_106,In_101);
nor U30 (N_30,In_340,In_98);
xnor U31 (N_31,In_672,In_359);
nor U32 (N_32,In_68,In_479);
and U33 (N_33,In_422,In_470);
nand U34 (N_34,In_50,In_258);
nor U35 (N_35,In_725,In_530);
nor U36 (N_36,In_34,In_449);
or U37 (N_37,In_706,In_738);
nand U38 (N_38,In_459,In_370);
nor U39 (N_39,In_587,In_46);
xor U40 (N_40,In_315,In_642);
xor U41 (N_41,In_485,In_405);
xor U42 (N_42,In_62,In_656);
and U43 (N_43,In_209,In_32);
and U44 (N_44,In_379,In_372);
nand U45 (N_45,In_303,In_747);
and U46 (N_46,In_337,In_245);
nand U47 (N_47,In_329,In_127);
or U48 (N_48,In_518,In_516);
xnor U49 (N_49,In_609,In_406);
nand U50 (N_50,In_43,In_74);
and U51 (N_51,In_263,In_239);
or U52 (N_52,In_570,In_24);
nor U53 (N_53,In_154,In_304);
nand U54 (N_54,In_17,In_183);
nand U55 (N_55,In_621,In_66);
nor U56 (N_56,In_634,In_698);
or U57 (N_57,In_710,In_99);
nor U58 (N_58,In_116,In_524);
and U59 (N_59,In_456,In_436);
nand U60 (N_60,In_293,In_463);
nor U61 (N_61,In_177,In_11);
nor U62 (N_62,In_421,In_282);
and U63 (N_63,In_583,In_616);
xnor U64 (N_64,In_54,In_22);
or U65 (N_65,In_588,In_633);
or U66 (N_66,In_102,In_313);
nor U67 (N_67,In_264,In_442);
and U68 (N_68,In_220,In_743);
nor U69 (N_69,In_145,In_185);
nand U70 (N_70,In_192,In_573);
and U71 (N_71,In_501,In_534);
or U72 (N_72,In_396,In_499);
nand U73 (N_73,In_654,In_724);
and U74 (N_74,In_733,In_146);
xor U75 (N_75,In_322,In_57);
xnor U76 (N_76,In_486,In_595);
or U77 (N_77,In_615,In_555);
xnor U78 (N_78,In_464,In_23);
nand U79 (N_79,In_492,In_650);
and U80 (N_80,In_212,In_551);
and U81 (N_81,In_346,In_348);
or U82 (N_82,In_197,In_166);
xnor U83 (N_83,In_637,In_179);
nor U84 (N_84,In_167,In_605);
nand U85 (N_85,In_56,In_748);
and U86 (N_86,In_675,In_607);
xnor U87 (N_87,In_497,In_417);
nor U88 (N_88,In_202,In_207);
nor U89 (N_89,In_150,In_172);
and U90 (N_90,In_623,In_376);
nor U91 (N_91,In_276,In_249);
or U92 (N_92,In_28,In_673);
nand U93 (N_93,In_309,In_671);
nand U94 (N_94,In_435,In_502);
or U95 (N_95,In_451,In_478);
xnor U96 (N_96,In_389,In_18);
and U97 (N_97,In_283,In_565);
or U98 (N_98,In_424,In_8);
nand U99 (N_99,In_728,In_250);
nand U100 (N_100,In_221,In_467);
nor U101 (N_101,In_9,In_606);
nand U102 (N_102,In_471,In_638);
and U103 (N_103,In_281,In_520);
nor U104 (N_104,In_692,In_614);
nand U105 (N_105,In_584,In_388);
and U106 (N_106,In_195,In_139);
nor U107 (N_107,In_320,In_203);
nand U108 (N_108,In_600,In_739);
nor U109 (N_109,In_407,In_448);
and U110 (N_110,In_361,In_187);
nor U111 (N_111,In_67,In_380);
or U112 (N_112,In_416,In_147);
nand U113 (N_113,In_493,In_613);
and U114 (N_114,In_240,In_465);
and U115 (N_115,In_174,In_664);
nor U116 (N_116,In_472,In_445);
nor U117 (N_117,In_545,In_686);
nor U118 (N_118,In_82,In_469);
or U119 (N_119,In_740,In_151);
nand U120 (N_120,In_323,In_399);
or U121 (N_121,In_10,In_114);
and U122 (N_122,In_326,In_306);
nand U123 (N_123,In_180,In_229);
nor U124 (N_124,In_257,In_602);
nor U125 (N_125,In_41,In_420);
and U126 (N_126,In_230,In_119);
and U127 (N_127,In_487,In_414);
and U128 (N_128,In_412,In_109);
and U129 (N_129,In_676,In_120);
nand U130 (N_130,In_333,In_59);
nand U131 (N_131,In_241,In_375);
nor U132 (N_132,In_318,In_419);
nand U133 (N_133,In_367,In_87);
or U134 (N_134,In_437,In_394);
and U135 (N_135,In_208,In_103);
xnor U136 (N_136,In_400,In_97);
or U137 (N_137,In_344,In_38);
and U138 (N_138,In_29,In_425);
xor U139 (N_139,In_188,In_374);
nand U140 (N_140,In_369,In_679);
xor U141 (N_141,In_117,In_196);
xor U142 (N_142,In_100,In_705);
nor U143 (N_143,In_35,In_491);
nor U144 (N_144,In_129,In_392);
or U145 (N_145,In_622,In_163);
nor U146 (N_146,In_560,In_291);
nor U147 (N_147,In_691,In_135);
or U148 (N_148,In_288,In_746);
or U149 (N_149,In_578,In_426);
nand U150 (N_150,In_75,In_182);
nor U151 (N_151,In_681,In_336);
xnor U152 (N_152,In_591,In_40);
and U153 (N_153,In_730,In_526);
and U154 (N_154,In_744,In_726);
or U155 (N_155,In_184,In_648);
or U156 (N_156,In_153,In_697);
or U157 (N_157,In_558,In_722);
or U158 (N_158,In_51,In_342);
nand U159 (N_159,In_734,In_317);
and U160 (N_160,In_49,In_599);
and U161 (N_161,In_44,In_47);
nand U162 (N_162,In_299,In_711);
nand U163 (N_163,In_217,In_636);
nand U164 (N_164,In_732,In_531);
or U165 (N_165,In_140,In_358);
or U166 (N_166,In_363,In_130);
or U167 (N_167,In_53,In_60);
or U168 (N_168,In_658,In_537);
nor U169 (N_169,In_301,In_6);
nand U170 (N_170,In_528,In_494);
or U171 (N_171,In_554,In_237);
and U172 (N_172,In_290,In_640);
or U173 (N_173,In_198,In_77);
nor U174 (N_174,In_660,In_398);
and U175 (N_175,In_37,In_111);
or U176 (N_176,In_736,In_611);
and U177 (N_177,In_521,In_158);
nor U178 (N_178,In_618,In_58);
or U179 (N_179,In_328,In_162);
and U180 (N_180,In_657,In_210);
nor U181 (N_181,In_384,In_619);
or U182 (N_182,In_149,In_527);
nor U183 (N_183,In_125,In_434);
nor U184 (N_184,In_123,In_383);
or U185 (N_185,In_401,In_556);
nand U186 (N_186,In_121,In_727);
and U187 (N_187,In_509,In_688);
or U188 (N_188,In_542,In_741);
or U189 (N_189,In_351,In_265);
nor U190 (N_190,In_289,In_176);
nor U191 (N_191,In_324,In_513);
nand U192 (N_192,In_696,In_577);
and U193 (N_193,In_511,In_409);
nor U194 (N_194,In_690,In_218);
and U195 (N_195,In_215,In_362);
or U196 (N_196,In_548,In_484);
and U197 (N_197,In_593,In_368);
or U198 (N_198,In_685,In_134);
or U199 (N_199,In_277,In_477);
nor U200 (N_200,In_271,In_723);
nor U201 (N_201,In_88,In_65);
nor U202 (N_202,In_439,In_311);
or U203 (N_203,In_397,In_25);
and U204 (N_204,In_48,In_693);
nand U205 (N_205,In_563,In_709);
nor U206 (N_206,In_76,In_226);
and U207 (N_207,In_256,In_700);
nand U208 (N_208,In_204,In_223);
nand U209 (N_209,In_16,In_122);
and U210 (N_210,In_143,In_356);
or U211 (N_211,In_107,In_255);
and U212 (N_212,In_663,In_3);
and U213 (N_213,In_371,In_70);
and U214 (N_214,In_300,In_745);
xnor U215 (N_215,In_458,In_128);
nand U216 (N_216,In_701,In_390);
nand U217 (N_217,In_393,In_680);
or U218 (N_218,In_253,In_428);
or U219 (N_219,In_168,In_720);
nand U220 (N_220,In_468,In_339);
and U221 (N_221,In_476,In_539);
and U222 (N_222,In_211,In_395);
and U223 (N_223,In_5,In_170);
xnor U224 (N_224,In_261,In_645);
and U225 (N_225,In_7,In_199);
nor U226 (N_226,In_544,In_225);
or U227 (N_227,In_391,In_444);
xor U228 (N_228,In_505,In_666);
nand U229 (N_229,In_1,In_525);
nand U230 (N_230,In_205,In_78);
or U231 (N_231,In_452,In_63);
or U232 (N_232,In_718,In_446);
nand U233 (N_233,In_643,In_330);
and U234 (N_234,In_546,In_161);
nor U235 (N_235,In_535,In_164);
nor U236 (N_236,In_552,In_729);
xor U237 (N_237,In_473,In_36);
nand U238 (N_238,In_308,In_699);
nor U239 (N_239,In_108,In_731);
or U240 (N_240,In_357,In_214);
nor U241 (N_241,In_21,In_332);
and U242 (N_242,In_110,In_105);
xor U243 (N_243,In_343,In_286);
and U244 (N_244,In_278,In_81);
nor U245 (N_245,In_547,In_626);
nor U246 (N_246,In_126,In_719);
or U247 (N_247,In_382,In_677);
or U248 (N_248,In_181,In_267);
nand U249 (N_249,In_651,In_42);
nor U250 (N_250,In_496,In_284);
nor U251 (N_251,In_550,In_659);
or U252 (N_252,In_440,In_137);
nand U253 (N_253,In_118,In_576);
xor U254 (N_254,In_191,In_232);
xor U255 (N_255,In_222,In_104);
and U256 (N_256,In_378,In_612);
nand U257 (N_257,In_441,In_352);
nand U258 (N_258,In_490,In_314);
nor U259 (N_259,In_589,In_26);
nor U260 (N_260,In_349,In_355);
and U261 (N_261,In_603,In_620);
nor U262 (N_262,In_341,In_579);
and U263 (N_263,In_189,In_334);
nand U264 (N_264,In_242,In_429);
nor U265 (N_265,In_175,In_236);
xor U266 (N_266,In_345,In_641);
nand U267 (N_267,In_604,In_280);
and U268 (N_268,In_387,In_321);
xor U269 (N_269,In_160,In_541);
or U270 (N_270,In_273,In_80);
nor U271 (N_271,In_410,In_694);
and U272 (N_272,In_272,In_235);
xnor U273 (N_273,In_206,In_704);
nor U274 (N_274,In_353,In_27);
xnor U275 (N_275,In_489,In_173);
xnor U276 (N_276,In_512,In_737);
nor U277 (N_277,In_402,In_403);
or U278 (N_278,In_590,In_586);
xnor U279 (N_279,In_86,In_132);
nor U280 (N_280,In_508,In_260);
xor U281 (N_281,In_562,In_702);
nand U282 (N_282,In_707,In_113);
and U283 (N_283,In_522,In_92);
nand U284 (N_284,In_186,In_597);
nor U285 (N_285,In_95,In_682);
or U286 (N_286,In_238,In_12);
xor U287 (N_287,In_275,In_495);
nand U288 (N_288,In_354,In_433);
nor U289 (N_289,In_287,In_712);
and U290 (N_290,In_4,In_52);
xor U291 (N_291,In_112,In_200);
nand U292 (N_292,In_649,In_244);
nand U293 (N_293,In_695,In_85);
nand U294 (N_294,In_247,In_432);
xor U295 (N_295,In_466,In_503);
or U296 (N_296,In_453,In_385);
or U297 (N_297,In_141,In_601);
xnor U298 (N_298,In_455,In_124);
or U299 (N_299,In_274,In_305);
nand U300 (N_300,In_500,In_561);
or U301 (N_301,In_592,In_668);
nand U302 (N_302,In_159,In_152);
nand U303 (N_303,In_450,In_504);
nor U304 (N_304,In_373,In_262);
xor U305 (N_305,In_316,In_716);
or U306 (N_306,In_683,In_646);
nand U307 (N_307,In_83,In_566);
or U308 (N_308,In_148,In_365);
nor U309 (N_309,In_430,In_662);
and U310 (N_310,In_93,In_14);
nand U311 (N_311,In_404,In_514);
xnor U312 (N_312,In_213,In_447);
nor U313 (N_313,In_631,In_157);
and U314 (N_314,In_571,In_131);
nand U315 (N_315,In_635,In_598);
xor U316 (N_316,In_625,In_251);
xnor U317 (N_317,In_481,In_285);
or U318 (N_318,In_510,In_39);
nand U319 (N_319,In_366,In_377);
nor U320 (N_320,In_294,In_415);
or U321 (N_321,In_193,In_575);
nor U322 (N_322,In_674,In_292);
or U323 (N_323,In_325,In_653);
nor U324 (N_324,In_310,In_687);
and U325 (N_325,In_543,In_248);
nor U326 (N_326,In_96,In_610);
or U327 (N_327,In_652,In_254);
nor U328 (N_328,In_714,In_228);
xor U329 (N_329,In_190,In_84);
nor U330 (N_330,In_482,In_227);
and U331 (N_331,In_219,In_708);
nand U332 (N_332,In_252,In_411);
nor U333 (N_333,In_364,In_523);
nand U334 (N_334,In_559,In_462);
nor U335 (N_335,In_749,In_268);
nor U336 (N_336,In_574,In_582);
and U337 (N_337,In_529,In_644);
or U338 (N_338,In_624,In_64);
or U339 (N_339,In_307,In_350);
nand U340 (N_340,In_302,In_568);
nand U341 (N_341,In_91,In_90);
and U342 (N_342,In_647,In_20);
nand U343 (N_343,In_713,In_89);
and U344 (N_344,In_259,In_224);
and U345 (N_345,In_564,In_443);
and U346 (N_346,In_661,In_461);
nand U347 (N_347,In_312,In_295);
nand U348 (N_348,In_735,In_608);
or U349 (N_349,In_418,In_45);
nand U350 (N_350,In_246,In_216);
or U351 (N_351,In_165,In_585);
or U352 (N_352,In_457,In_627);
nand U353 (N_353,In_670,In_721);
or U354 (N_354,In_684,In_498);
nor U355 (N_355,In_201,In_632);
xor U356 (N_356,In_233,In_665);
or U357 (N_357,In_515,In_234);
nor U358 (N_358,In_194,In_79);
nand U359 (N_359,In_71,In_630);
or U360 (N_360,In_454,In_142);
nand U361 (N_361,In_15,In_655);
nor U362 (N_362,In_483,In_386);
nor U363 (N_363,In_338,In_580);
nand U364 (N_364,In_427,In_474);
or U365 (N_365,In_61,In_298);
nor U366 (N_366,In_279,In_360);
nand U367 (N_367,In_155,In_667);
nor U368 (N_368,In_488,In_269);
nor U369 (N_369,In_594,In_567);
nand U370 (N_370,In_13,In_596);
or U371 (N_371,In_689,In_69);
nor U372 (N_372,In_327,In_480);
nor U373 (N_373,In_506,In_169);
nor U374 (N_374,In_572,In_243);
or U375 (N_375,In_176,In_485);
and U376 (N_376,In_684,In_540);
xnor U377 (N_377,In_604,In_367);
xor U378 (N_378,In_230,In_156);
nand U379 (N_379,In_57,In_218);
nor U380 (N_380,In_614,In_473);
or U381 (N_381,In_42,In_241);
nor U382 (N_382,In_516,In_196);
and U383 (N_383,In_4,In_74);
and U384 (N_384,In_222,In_725);
or U385 (N_385,In_102,In_308);
xnor U386 (N_386,In_388,In_99);
or U387 (N_387,In_135,In_79);
xnor U388 (N_388,In_675,In_730);
nand U389 (N_389,In_62,In_246);
nand U390 (N_390,In_260,In_373);
and U391 (N_391,In_517,In_490);
and U392 (N_392,In_458,In_75);
or U393 (N_393,In_452,In_276);
or U394 (N_394,In_464,In_81);
or U395 (N_395,In_136,In_188);
and U396 (N_396,In_668,In_607);
or U397 (N_397,In_580,In_514);
xnor U398 (N_398,In_384,In_317);
and U399 (N_399,In_219,In_681);
or U400 (N_400,In_240,In_609);
nor U401 (N_401,In_219,In_593);
nor U402 (N_402,In_580,In_158);
nor U403 (N_403,In_178,In_367);
or U404 (N_404,In_569,In_29);
nand U405 (N_405,In_422,In_731);
or U406 (N_406,In_226,In_26);
nor U407 (N_407,In_244,In_655);
nor U408 (N_408,In_682,In_167);
nor U409 (N_409,In_180,In_481);
nor U410 (N_410,In_295,In_606);
nor U411 (N_411,In_245,In_703);
and U412 (N_412,In_353,In_436);
nand U413 (N_413,In_350,In_670);
xor U414 (N_414,In_715,In_392);
nand U415 (N_415,In_632,In_131);
or U416 (N_416,In_701,In_131);
nand U417 (N_417,In_221,In_60);
nand U418 (N_418,In_521,In_458);
or U419 (N_419,In_563,In_444);
nand U420 (N_420,In_521,In_421);
nor U421 (N_421,In_400,In_366);
or U422 (N_422,In_352,In_157);
nand U423 (N_423,In_506,In_554);
or U424 (N_424,In_522,In_524);
or U425 (N_425,In_209,In_239);
xnor U426 (N_426,In_189,In_545);
nor U427 (N_427,In_26,In_131);
and U428 (N_428,In_158,In_244);
nand U429 (N_429,In_115,In_481);
and U430 (N_430,In_384,In_394);
and U431 (N_431,In_181,In_695);
nor U432 (N_432,In_182,In_250);
nand U433 (N_433,In_489,In_178);
and U434 (N_434,In_496,In_304);
xor U435 (N_435,In_286,In_190);
and U436 (N_436,In_714,In_398);
nand U437 (N_437,In_604,In_644);
and U438 (N_438,In_493,In_130);
or U439 (N_439,In_444,In_637);
and U440 (N_440,In_492,In_288);
nor U441 (N_441,In_621,In_23);
nor U442 (N_442,In_146,In_475);
and U443 (N_443,In_738,In_268);
or U444 (N_444,In_574,In_9);
nand U445 (N_445,In_246,In_75);
or U446 (N_446,In_383,In_277);
and U447 (N_447,In_682,In_89);
xnor U448 (N_448,In_458,In_665);
or U449 (N_449,In_624,In_548);
nand U450 (N_450,In_524,In_737);
nor U451 (N_451,In_385,In_216);
nand U452 (N_452,In_219,In_423);
xor U453 (N_453,In_555,In_549);
or U454 (N_454,In_108,In_187);
and U455 (N_455,In_462,In_489);
xor U456 (N_456,In_229,In_90);
nand U457 (N_457,In_344,In_472);
and U458 (N_458,In_312,In_703);
and U459 (N_459,In_22,In_595);
xnor U460 (N_460,In_603,In_78);
xor U461 (N_461,In_238,In_640);
and U462 (N_462,In_738,In_330);
xnor U463 (N_463,In_518,In_586);
nor U464 (N_464,In_195,In_680);
or U465 (N_465,In_454,In_320);
and U466 (N_466,In_215,In_94);
and U467 (N_467,In_553,In_546);
or U468 (N_468,In_19,In_259);
nor U469 (N_469,In_651,In_83);
nand U470 (N_470,In_693,In_145);
and U471 (N_471,In_149,In_268);
nor U472 (N_472,In_351,In_219);
and U473 (N_473,In_253,In_627);
nor U474 (N_474,In_691,In_736);
nand U475 (N_475,In_101,In_463);
or U476 (N_476,In_160,In_529);
or U477 (N_477,In_108,In_679);
and U478 (N_478,In_680,In_404);
and U479 (N_479,In_519,In_716);
nand U480 (N_480,In_340,In_345);
nor U481 (N_481,In_203,In_83);
and U482 (N_482,In_385,In_460);
and U483 (N_483,In_205,In_190);
or U484 (N_484,In_380,In_505);
nor U485 (N_485,In_229,In_588);
and U486 (N_486,In_697,In_672);
nand U487 (N_487,In_381,In_461);
and U488 (N_488,In_29,In_483);
xor U489 (N_489,In_493,In_480);
nand U490 (N_490,In_360,In_402);
nand U491 (N_491,In_242,In_53);
or U492 (N_492,In_391,In_385);
and U493 (N_493,In_16,In_209);
nand U494 (N_494,In_172,In_397);
and U495 (N_495,In_151,In_252);
nor U496 (N_496,In_200,In_287);
and U497 (N_497,In_252,In_544);
and U498 (N_498,In_464,In_553);
and U499 (N_499,In_582,In_339);
nor U500 (N_500,N_232,N_268);
and U501 (N_501,N_477,N_83);
and U502 (N_502,N_68,N_470);
nor U503 (N_503,N_362,N_177);
and U504 (N_504,N_246,N_230);
nor U505 (N_505,N_270,N_72);
and U506 (N_506,N_158,N_264);
nor U507 (N_507,N_408,N_236);
and U508 (N_508,N_152,N_441);
nor U509 (N_509,N_340,N_314);
xnor U510 (N_510,N_492,N_315);
nand U511 (N_511,N_222,N_198);
nor U512 (N_512,N_214,N_52);
and U513 (N_513,N_128,N_143);
xor U514 (N_514,N_61,N_175);
nor U515 (N_515,N_107,N_226);
nand U516 (N_516,N_131,N_469);
and U517 (N_517,N_355,N_280);
nor U518 (N_518,N_167,N_378);
nor U519 (N_519,N_407,N_133);
nand U520 (N_520,N_365,N_259);
nand U521 (N_521,N_425,N_93);
nor U522 (N_522,N_377,N_217);
nor U523 (N_523,N_460,N_58);
xnor U524 (N_524,N_276,N_458);
nand U525 (N_525,N_38,N_242);
nor U526 (N_526,N_307,N_115);
xor U527 (N_527,N_162,N_266);
nand U528 (N_528,N_433,N_326);
and U529 (N_529,N_216,N_211);
and U530 (N_530,N_130,N_79);
and U531 (N_531,N_453,N_112);
xnor U532 (N_532,N_185,N_209);
or U533 (N_533,N_244,N_106);
and U534 (N_534,N_406,N_389);
nand U535 (N_535,N_105,N_339);
nand U536 (N_536,N_27,N_431);
or U537 (N_537,N_60,N_289);
nor U538 (N_538,N_284,N_486);
nand U539 (N_539,N_301,N_239);
xor U540 (N_540,N_159,N_456);
and U541 (N_541,N_450,N_403);
nor U542 (N_542,N_138,N_50);
nor U543 (N_543,N_415,N_135);
xor U544 (N_544,N_480,N_76);
xnor U545 (N_545,N_99,N_25);
nand U546 (N_546,N_464,N_325);
and U547 (N_547,N_430,N_300);
or U548 (N_548,N_41,N_288);
and U549 (N_549,N_191,N_54);
nor U550 (N_550,N_95,N_488);
nor U551 (N_551,N_279,N_0);
or U552 (N_552,N_74,N_468);
nand U553 (N_553,N_420,N_240);
or U554 (N_554,N_479,N_33);
nor U555 (N_555,N_418,N_461);
and U556 (N_556,N_328,N_364);
nor U557 (N_557,N_146,N_102);
and U558 (N_558,N_67,N_118);
nor U559 (N_559,N_385,N_11);
xor U560 (N_560,N_207,N_64);
xnor U561 (N_561,N_134,N_168);
nand U562 (N_562,N_21,N_332);
nor U563 (N_563,N_234,N_275);
and U564 (N_564,N_44,N_14);
and U565 (N_565,N_117,N_59);
and U566 (N_566,N_353,N_17);
and U567 (N_567,N_104,N_84);
or U568 (N_568,N_229,N_97);
and U569 (N_569,N_394,N_87);
nand U570 (N_570,N_195,N_210);
or U571 (N_571,N_132,N_243);
xor U572 (N_572,N_161,N_205);
or U573 (N_573,N_449,N_475);
nand U574 (N_574,N_111,N_125);
and U575 (N_575,N_145,N_483);
nor U576 (N_576,N_457,N_184);
nand U577 (N_577,N_178,N_150);
nand U578 (N_578,N_272,N_291);
and U579 (N_579,N_327,N_192);
nand U580 (N_580,N_422,N_330);
or U581 (N_581,N_429,N_71);
or U582 (N_582,N_305,N_2);
nand U583 (N_583,N_361,N_452);
nor U584 (N_584,N_320,N_400);
nor U585 (N_585,N_271,N_421);
nor U586 (N_586,N_379,N_487);
nor U587 (N_587,N_194,N_7);
and U588 (N_588,N_108,N_174);
xnor U589 (N_589,N_251,N_18);
nor U590 (N_590,N_81,N_447);
nand U591 (N_591,N_472,N_366);
nor U592 (N_592,N_42,N_395);
nor U593 (N_593,N_160,N_293);
and U594 (N_594,N_173,N_169);
xor U595 (N_595,N_485,N_48);
nand U596 (N_596,N_181,N_70);
nor U597 (N_597,N_380,N_298);
and U598 (N_598,N_345,N_16);
nor U599 (N_599,N_490,N_215);
nor U600 (N_600,N_374,N_85);
and U601 (N_601,N_120,N_176);
or U602 (N_602,N_22,N_318);
and U603 (N_603,N_75,N_333);
xnor U604 (N_604,N_156,N_122);
nor U605 (N_605,N_261,N_297);
or U606 (N_606,N_423,N_113);
and U607 (N_607,N_121,N_166);
nor U608 (N_608,N_204,N_454);
or U609 (N_609,N_98,N_155);
nor U610 (N_610,N_89,N_390);
nor U611 (N_611,N_193,N_393);
nand U612 (N_612,N_123,N_474);
nand U613 (N_613,N_416,N_5);
and U614 (N_614,N_187,N_428);
or U615 (N_615,N_283,N_331);
nor U616 (N_616,N_248,N_13);
nor U617 (N_617,N_46,N_322);
nand U618 (N_618,N_323,N_182);
or U619 (N_619,N_317,N_308);
and U620 (N_620,N_252,N_43);
nor U621 (N_621,N_90,N_281);
and U622 (N_622,N_496,N_45);
and U623 (N_623,N_412,N_459);
or U624 (N_624,N_258,N_218);
and U625 (N_625,N_201,N_373);
and U626 (N_626,N_199,N_171);
xnor U627 (N_627,N_249,N_88);
or U628 (N_628,N_338,N_260);
and U629 (N_629,N_354,N_294);
nor U630 (N_630,N_419,N_212);
and U631 (N_631,N_286,N_147);
nor U632 (N_632,N_381,N_263);
or U633 (N_633,N_219,N_6);
and U634 (N_634,N_274,N_140);
xnor U635 (N_635,N_144,N_91);
nand U636 (N_636,N_269,N_278);
and U637 (N_637,N_141,N_186);
nand U638 (N_638,N_273,N_387);
and U639 (N_639,N_376,N_228);
nor U640 (N_640,N_304,N_164);
xnor U641 (N_641,N_179,N_348);
nand U642 (N_642,N_28,N_329);
nor U643 (N_643,N_129,N_398);
nor U644 (N_644,N_321,N_440);
and U645 (N_645,N_473,N_324);
xor U646 (N_646,N_335,N_336);
nand U647 (N_647,N_342,N_445);
nor U648 (N_648,N_465,N_96);
nor U649 (N_649,N_388,N_78);
or U650 (N_650,N_489,N_55);
nand U651 (N_651,N_165,N_9);
nor U652 (N_652,N_221,N_39);
or U653 (N_653,N_53,N_495);
or U654 (N_654,N_316,N_358);
or U655 (N_655,N_312,N_63);
or U656 (N_656,N_344,N_357);
or U657 (N_657,N_392,N_383);
nor U658 (N_658,N_56,N_200);
xnor U659 (N_659,N_265,N_127);
or U660 (N_660,N_206,N_92);
nand U661 (N_661,N_466,N_65);
or U662 (N_662,N_346,N_148);
and U663 (N_663,N_334,N_116);
nor U664 (N_664,N_73,N_413);
and U665 (N_665,N_153,N_227);
nand U666 (N_666,N_247,N_8);
and U667 (N_667,N_391,N_47);
nand U668 (N_668,N_23,N_220);
nor U669 (N_669,N_292,N_31);
or U670 (N_670,N_463,N_1);
xor U671 (N_671,N_94,N_402);
nand U672 (N_672,N_223,N_208);
nor U673 (N_673,N_36,N_302);
or U674 (N_674,N_444,N_497);
nand U675 (N_675,N_313,N_409);
nor U676 (N_676,N_319,N_238);
nor U677 (N_677,N_352,N_434);
nand U678 (N_678,N_3,N_436);
nor U679 (N_679,N_375,N_396);
or U680 (N_680,N_494,N_349);
or U681 (N_681,N_371,N_277);
and U682 (N_682,N_382,N_233);
xor U683 (N_683,N_424,N_399);
nor U684 (N_684,N_401,N_157);
xor U685 (N_685,N_196,N_267);
and U686 (N_686,N_19,N_109);
xnor U687 (N_687,N_149,N_435);
or U688 (N_688,N_411,N_467);
or U689 (N_689,N_310,N_341);
and U690 (N_690,N_484,N_438);
nor U691 (N_691,N_427,N_356);
or U692 (N_692,N_237,N_69);
and U693 (N_693,N_190,N_367);
nor U694 (N_694,N_347,N_476);
nor U695 (N_695,N_363,N_482);
or U696 (N_696,N_369,N_197);
nand U697 (N_697,N_82,N_303);
xnor U698 (N_698,N_410,N_180);
or U699 (N_699,N_245,N_493);
nand U700 (N_700,N_372,N_241);
nand U701 (N_701,N_255,N_110);
nand U702 (N_702,N_163,N_126);
xnor U703 (N_703,N_405,N_359);
nand U704 (N_704,N_124,N_350);
and U705 (N_705,N_462,N_451);
nor U706 (N_706,N_231,N_80);
nor U707 (N_707,N_290,N_235);
and U708 (N_708,N_437,N_360);
and U709 (N_709,N_417,N_491);
nand U710 (N_710,N_32,N_103);
or U711 (N_711,N_285,N_287);
nand U712 (N_712,N_426,N_225);
and U713 (N_713,N_202,N_35);
nor U714 (N_714,N_498,N_296);
nor U715 (N_715,N_370,N_256);
nor U716 (N_716,N_337,N_343);
or U717 (N_717,N_101,N_309);
nor U718 (N_718,N_282,N_142);
nand U719 (N_719,N_448,N_170);
nand U720 (N_720,N_10,N_114);
and U721 (N_721,N_100,N_29);
or U722 (N_722,N_30,N_137);
or U723 (N_723,N_203,N_49);
nand U724 (N_724,N_34,N_24);
nor U725 (N_725,N_254,N_20);
xor U726 (N_726,N_183,N_213);
nor U727 (N_727,N_119,N_15);
or U728 (N_728,N_188,N_12);
and U729 (N_729,N_40,N_62);
or U730 (N_730,N_37,N_478);
nor U731 (N_731,N_139,N_439);
nand U732 (N_732,N_224,N_136);
and U733 (N_733,N_295,N_57);
nand U734 (N_734,N_250,N_257);
nor U735 (N_735,N_154,N_262);
xnor U736 (N_736,N_443,N_432);
nand U737 (N_737,N_26,N_306);
or U738 (N_738,N_66,N_414);
nand U739 (N_739,N_384,N_172);
or U740 (N_740,N_151,N_442);
nor U741 (N_741,N_189,N_455);
xor U742 (N_742,N_397,N_446);
nor U743 (N_743,N_253,N_299);
xnor U744 (N_744,N_86,N_481);
nor U745 (N_745,N_368,N_351);
nand U746 (N_746,N_499,N_404);
or U747 (N_747,N_77,N_471);
and U748 (N_748,N_4,N_311);
and U749 (N_749,N_386,N_51);
nand U750 (N_750,N_473,N_79);
nand U751 (N_751,N_143,N_6);
nand U752 (N_752,N_139,N_160);
or U753 (N_753,N_226,N_163);
nand U754 (N_754,N_131,N_278);
and U755 (N_755,N_379,N_472);
or U756 (N_756,N_23,N_466);
and U757 (N_757,N_481,N_299);
or U758 (N_758,N_415,N_169);
nand U759 (N_759,N_257,N_339);
or U760 (N_760,N_177,N_74);
and U761 (N_761,N_42,N_352);
and U762 (N_762,N_127,N_302);
and U763 (N_763,N_269,N_124);
and U764 (N_764,N_287,N_166);
xnor U765 (N_765,N_322,N_168);
or U766 (N_766,N_217,N_371);
nor U767 (N_767,N_52,N_365);
nand U768 (N_768,N_341,N_5);
or U769 (N_769,N_292,N_309);
nor U770 (N_770,N_484,N_379);
or U771 (N_771,N_285,N_463);
nand U772 (N_772,N_340,N_382);
or U773 (N_773,N_70,N_194);
and U774 (N_774,N_331,N_358);
nor U775 (N_775,N_173,N_60);
and U776 (N_776,N_434,N_261);
nand U777 (N_777,N_437,N_409);
nor U778 (N_778,N_67,N_231);
xor U779 (N_779,N_208,N_410);
nor U780 (N_780,N_334,N_117);
nor U781 (N_781,N_438,N_203);
or U782 (N_782,N_9,N_17);
nor U783 (N_783,N_309,N_303);
nor U784 (N_784,N_91,N_408);
nand U785 (N_785,N_350,N_102);
nand U786 (N_786,N_317,N_280);
nor U787 (N_787,N_436,N_222);
or U788 (N_788,N_101,N_282);
nand U789 (N_789,N_84,N_316);
and U790 (N_790,N_498,N_494);
nor U791 (N_791,N_200,N_431);
or U792 (N_792,N_389,N_152);
nor U793 (N_793,N_288,N_302);
nor U794 (N_794,N_483,N_496);
nor U795 (N_795,N_164,N_69);
nand U796 (N_796,N_238,N_147);
nand U797 (N_797,N_332,N_293);
nor U798 (N_798,N_222,N_248);
and U799 (N_799,N_285,N_457);
and U800 (N_800,N_237,N_122);
nand U801 (N_801,N_494,N_209);
nand U802 (N_802,N_96,N_241);
xnor U803 (N_803,N_409,N_101);
nor U804 (N_804,N_422,N_433);
nor U805 (N_805,N_414,N_469);
nor U806 (N_806,N_392,N_467);
nand U807 (N_807,N_37,N_303);
and U808 (N_808,N_332,N_91);
or U809 (N_809,N_439,N_387);
nand U810 (N_810,N_51,N_214);
or U811 (N_811,N_145,N_409);
xor U812 (N_812,N_23,N_162);
nor U813 (N_813,N_290,N_461);
nand U814 (N_814,N_360,N_296);
and U815 (N_815,N_328,N_210);
nor U816 (N_816,N_8,N_483);
nor U817 (N_817,N_267,N_450);
and U818 (N_818,N_78,N_99);
nand U819 (N_819,N_211,N_198);
nor U820 (N_820,N_40,N_59);
and U821 (N_821,N_494,N_361);
and U822 (N_822,N_242,N_63);
nand U823 (N_823,N_487,N_33);
nor U824 (N_824,N_19,N_107);
nand U825 (N_825,N_268,N_78);
xor U826 (N_826,N_132,N_316);
or U827 (N_827,N_381,N_247);
or U828 (N_828,N_496,N_404);
nand U829 (N_829,N_462,N_465);
xor U830 (N_830,N_243,N_402);
and U831 (N_831,N_389,N_379);
and U832 (N_832,N_283,N_475);
or U833 (N_833,N_83,N_396);
nor U834 (N_834,N_183,N_342);
nand U835 (N_835,N_51,N_275);
and U836 (N_836,N_135,N_449);
or U837 (N_837,N_328,N_142);
xor U838 (N_838,N_242,N_444);
or U839 (N_839,N_403,N_436);
nand U840 (N_840,N_77,N_342);
nor U841 (N_841,N_22,N_496);
nor U842 (N_842,N_280,N_327);
and U843 (N_843,N_355,N_84);
xnor U844 (N_844,N_170,N_56);
nand U845 (N_845,N_62,N_319);
nand U846 (N_846,N_7,N_159);
and U847 (N_847,N_88,N_196);
or U848 (N_848,N_9,N_195);
and U849 (N_849,N_42,N_434);
nand U850 (N_850,N_151,N_303);
nor U851 (N_851,N_468,N_243);
or U852 (N_852,N_327,N_244);
and U853 (N_853,N_491,N_269);
and U854 (N_854,N_5,N_411);
xor U855 (N_855,N_366,N_491);
or U856 (N_856,N_69,N_298);
nor U857 (N_857,N_432,N_232);
and U858 (N_858,N_145,N_155);
xor U859 (N_859,N_246,N_446);
and U860 (N_860,N_294,N_283);
nor U861 (N_861,N_61,N_401);
and U862 (N_862,N_374,N_255);
nor U863 (N_863,N_465,N_40);
nor U864 (N_864,N_104,N_483);
nand U865 (N_865,N_336,N_141);
nor U866 (N_866,N_40,N_331);
xor U867 (N_867,N_483,N_369);
or U868 (N_868,N_472,N_9);
nor U869 (N_869,N_41,N_384);
nor U870 (N_870,N_9,N_201);
or U871 (N_871,N_263,N_134);
or U872 (N_872,N_186,N_71);
xor U873 (N_873,N_443,N_72);
or U874 (N_874,N_416,N_485);
xor U875 (N_875,N_433,N_475);
nand U876 (N_876,N_241,N_305);
nand U877 (N_877,N_91,N_131);
and U878 (N_878,N_474,N_194);
xnor U879 (N_879,N_97,N_39);
and U880 (N_880,N_394,N_140);
and U881 (N_881,N_293,N_482);
and U882 (N_882,N_360,N_429);
and U883 (N_883,N_195,N_248);
or U884 (N_884,N_57,N_267);
nand U885 (N_885,N_86,N_220);
and U886 (N_886,N_111,N_424);
or U887 (N_887,N_148,N_166);
and U888 (N_888,N_13,N_156);
and U889 (N_889,N_280,N_173);
and U890 (N_890,N_475,N_439);
or U891 (N_891,N_203,N_221);
xnor U892 (N_892,N_293,N_155);
xnor U893 (N_893,N_280,N_193);
or U894 (N_894,N_431,N_355);
and U895 (N_895,N_342,N_352);
and U896 (N_896,N_59,N_494);
and U897 (N_897,N_176,N_490);
nand U898 (N_898,N_451,N_5);
nand U899 (N_899,N_340,N_85);
and U900 (N_900,N_72,N_448);
nor U901 (N_901,N_130,N_9);
nand U902 (N_902,N_43,N_221);
nor U903 (N_903,N_53,N_463);
xnor U904 (N_904,N_458,N_483);
and U905 (N_905,N_243,N_147);
and U906 (N_906,N_490,N_486);
nor U907 (N_907,N_436,N_341);
nand U908 (N_908,N_381,N_380);
nand U909 (N_909,N_336,N_329);
or U910 (N_910,N_217,N_350);
nor U911 (N_911,N_307,N_108);
and U912 (N_912,N_463,N_374);
and U913 (N_913,N_365,N_153);
xnor U914 (N_914,N_112,N_196);
nand U915 (N_915,N_92,N_72);
and U916 (N_916,N_263,N_453);
or U917 (N_917,N_219,N_497);
or U918 (N_918,N_187,N_345);
or U919 (N_919,N_386,N_241);
nand U920 (N_920,N_273,N_399);
nand U921 (N_921,N_462,N_343);
nor U922 (N_922,N_112,N_444);
xor U923 (N_923,N_170,N_487);
nand U924 (N_924,N_162,N_240);
nand U925 (N_925,N_106,N_47);
nor U926 (N_926,N_112,N_96);
nand U927 (N_927,N_4,N_27);
xor U928 (N_928,N_429,N_46);
or U929 (N_929,N_441,N_317);
nor U930 (N_930,N_449,N_105);
nand U931 (N_931,N_349,N_372);
nor U932 (N_932,N_18,N_158);
nand U933 (N_933,N_279,N_158);
xor U934 (N_934,N_154,N_490);
nor U935 (N_935,N_393,N_373);
nor U936 (N_936,N_79,N_380);
and U937 (N_937,N_425,N_167);
nor U938 (N_938,N_183,N_4);
and U939 (N_939,N_308,N_368);
xnor U940 (N_940,N_465,N_216);
or U941 (N_941,N_52,N_289);
nor U942 (N_942,N_145,N_397);
nand U943 (N_943,N_299,N_257);
nor U944 (N_944,N_43,N_345);
and U945 (N_945,N_76,N_119);
xnor U946 (N_946,N_298,N_251);
nor U947 (N_947,N_389,N_225);
xor U948 (N_948,N_387,N_154);
nand U949 (N_949,N_331,N_13);
and U950 (N_950,N_208,N_363);
nor U951 (N_951,N_243,N_199);
nand U952 (N_952,N_74,N_490);
nor U953 (N_953,N_185,N_419);
or U954 (N_954,N_312,N_310);
nand U955 (N_955,N_387,N_12);
nand U956 (N_956,N_184,N_130);
or U957 (N_957,N_198,N_429);
nand U958 (N_958,N_3,N_52);
or U959 (N_959,N_461,N_120);
nor U960 (N_960,N_205,N_399);
and U961 (N_961,N_11,N_265);
nand U962 (N_962,N_360,N_225);
and U963 (N_963,N_79,N_52);
nor U964 (N_964,N_4,N_148);
nor U965 (N_965,N_220,N_247);
and U966 (N_966,N_86,N_123);
or U967 (N_967,N_107,N_84);
or U968 (N_968,N_283,N_244);
nand U969 (N_969,N_84,N_285);
xnor U970 (N_970,N_419,N_21);
nand U971 (N_971,N_36,N_334);
nand U972 (N_972,N_285,N_115);
nand U973 (N_973,N_59,N_318);
nor U974 (N_974,N_411,N_457);
nand U975 (N_975,N_381,N_249);
or U976 (N_976,N_375,N_458);
nand U977 (N_977,N_451,N_326);
nor U978 (N_978,N_89,N_458);
nor U979 (N_979,N_213,N_53);
nor U980 (N_980,N_100,N_13);
nand U981 (N_981,N_485,N_245);
or U982 (N_982,N_352,N_296);
nor U983 (N_983,N_106,N_12);
nand U984 (N_984,N_340,N_112);
or U985 (N_985,N_303,N_498);
nor U986 (N_986,N_462,N_337);
or U987 (N_987,N_387,N_151);
and U988 (N_988,N_223,N_37);
and U989 (N_989,N_227,N_456);
nand U990 (N_990,N_294,N_290);
nand U991 (N_991,N_497,N_140);
or U992 (N_992,N_341,N_490);
and U993 (N_993,N_483,N_49);
and U994 (N_994,N_457,N_346);
or U995 (N_995,N_367,N_384);
or U996 (N_996,N_278,N_95);
or U997 (N_997,N_453,N_121);
and U998 (N_998,N_367,N_448);
and U999 (N_999,N_302,N_435);
nor U1000 (N_1000,N_736,N_632);
nor U1001 (N_1001,N_567,N_819);
and U1002 (N_1002,N_816,N_780);
nand U1003 (N_1003,N_617,N_501);
nand U1004 (N_1004,N_626,N_708);
nand U1005 (N_1005,N_600,N_956);
or U1006 (N_1006,N_767,N_504);
nor U1007 (N_1007,N_815,N_875);
xnor U1008 (N_1008,N_846,N_987);
nand U1009 (N_1009,N_863,N_661);
nand U1010 (N_1010,N_986,N_768);
nand U1011 (N_1011,N_784,N_518);
or U1012 (N_1012,N_836,N_868);
nand U1013 (N_1013,N_637,N_893);
and U1014 (N_1014,N_603,N_786);
nor U1015 (N_1015,N_817,N_998);
and U1016 (N_1016,N_562,N_579);
and U1017 (N_1017,N_520,N_808);
nand U1018 (N_1018,N_720,N_828);
xor U1019 (N_1019,N_545,N_939);
and U1020 (N_1020,N_787,N_920);
or U1021 (N_1021,N_781,N_599);
and U1022 (N_1022,N_728,N_739);
and U1023 (N_1023,N_552,N_914);
and U1024 (N_1024,N_902,N_872);
nand U1025 (N_1025,N_740,N_764);
or U1026 (N_1026,N_591,N_992);
and U1027 (N_1027,N_905,N_649);
and U1028 (N_1028,N_578,N_548);
nand U1029 (N_1029,N_732,N_832);
and U1030 (N_1030,N_703,N_702);
or U1031 (N_1031,N_970,N_514);
xnor U1032 (N_1032,N_722,N_916);
nor U1033 (N_1033,N_978,N_789);
nand U1034 (N_1034,N_745,N_964);
nand U1035 (N_1035,N_766,N_934);
nor U1036 (N_1036,N_800,N_926);
or U1037 (N_1037,N_509,N_754);
nor U1038 (N_1038,N_560,N_952);
or U1039 (N_1039,N_891,N_746);
nor U1040 (N_1040,N_625,N_663);
nand U1041 (N_1041,N_593,N_719);
and U1042 (N_1042,N_762,N_575);
or U1043 (N_1043,N_553,N_790);
and U1044 (N_1044,N_627,N_761);
xor U1045 (N_1045,N_750,N_997);
or U1046 (N_1046,N_515,N_707);
nor U1047 (N_1047,N_500,N_915);
nor U1048 (N_1048,N_644,N_782);
or U1049 (N_1049,N_733,N_948);
nand U1050 (N_1050,N_711,N_531);
and U1051 (N_1051,N_512,N_674);
and U1052 (N_1052,N_540,N_859);
nor U1053 (N_1053,N_508,N_933);
nand U1054 (N_1054,N_931,N_641);
nor U1055 (N_1055,N_801,N_831);
or U1056 (N_1056,N_601,N_555);
nand U1057 (N_1057,N_568,N_797);
nand U1058 (N_1058,N_855,N_994);
and U1059 (N_1059,N_587,N_658);
or U1060 (N_1060,N_772,N_670);
and U1061 (N_1061,N_922,N_731);
xor U1062 (N_1062,N_536,N_791);
or U1063 (N_1063,N_660,N_543);
nor U1064 (N_1064,N_506,N_995);
and U1065 (N_1065,N_608,N_984);
nand U1066 (N_1066,N_615,N_597);
nor U1067 (N_1067,N_752,N_982);
nand U1068 (N_1068,N_770,N_849);
nand U1069 (N_1069,N_737,N_643);
nand U1070 (N_1070,N_699,N_877);
nor U1071 (N_1071,N_897,N_847);
nand U1072 (N_1072,N_908,N_581);
and U1073 (N_1073,N_704,N_673);
or U1074 (N_1074,N_503,N_941);
xor U1075 (N_1075,N_590,N_651);
and U1076 (N_1076,N_687,N_843);
nand U1077 (N_1077,N_694,N_585);
or U1078 (N_1078,N_979,N_974);
xor U1079 (N_1079,N_813,N_633);
and U1080 (N_1080,N_814,N_901);
and U1081 (N_1081,N_717,N_577);
or U1082 (N_1082,N_713,N_550);
or U1083 (N_1083,N_676,N_785);
or U1084 (N_1084,N_534,N_944);
nor U1085 (N_1085,N_796,N_692);
or U1086 (N_1086,N_923,N_885);
and U1087 (N_1087,N_878,N_793);
or U1088 (N_1088,N_876,N_613);
nand U1089 (N_1089,N_924,N_822);
nand U1090 (N_1090,N_749,N_530);
and U1091 (N_1091,N_844,N_748);
nor U1092 (N_1092,N_610,N_758);
and U1093 (N_1093,N_773,N_630);
and U1094 (N_1094,N_912,N_738);
or U1095 (N_1095,N_946,N_654);
and U1096 (N_1096,N_678,N_918);
nand U1097 (N_1097,N_873,N_525);
and U1098 (N_1098,N_857,N_693);
nor U1099 (N_1099,N_958,N_624);
and U1100 (N_1100,N_806,N_892);
and U1101 (N_1101,N_835,N_842);
or U1102 (N_1102,N_913,N_642);
and U1103 (N_1103,N_963,N_726);
nor U1104 (N_1104,N_535,N_932);
nand U1105 (N_1105,N_852,N_742);
nor U1106 (N_1106,N_664,N_689);
or U1107 (N_1107,N_950,N_966);
nor U1108 (N_1108,N_517,N_904);
nand U1109 (N_1109,N_606,N_975);
or U1110 (N_1110,N_554,N_820);
and U1111 (N_1111,N_823,N_710);
xor U1112 (N_1112,N_690,N_821);
or U1113 (N_1113,N_803,N_866);
xor U1114 (N_1114,N_727,N_840);
nor U1115 (N_1115,N_779,N_989);
nand U1116 (N_1116,N_516,N_935);
and U1117 (N_1117,N_705,N_735);
nor U1118 (N_1118,N_700,N_594);
nor U1119 (N_1119,N_596,N_869);
xnor U1120 (N_1120,N_839,N_672);
nand U1121 (N_1121,N_561,N_804);
nor U1122 (N_1122,N_684,N_522);
and U1123 (N_1123,N_653,N_943);
nand U1124 (N_1124,N_580,N_629);
nor U1125 (N_1125,N_883,N_871);
or U1126 (N_1126,N_854,N_675);
nor U1127 (N_1127,N_917,N_861);
xor U1128 (N_1128,N_583,N_775);
nor U1129 (N_1129,N_524,N_756);
nand U1130 (N_1130,N_698,N_906);
xnor U1131 (N_1131,N_755,N_774);
nand U1132 (N_1132,N_695,N_896);
and U1133 (N_1133,N_955,N_993);
or U1134 (N_1134,N_810,N_930);
and U1135 (N_1135,N_688,N_841);
nor U1136 (N_1136,N_715,N_763);
or U1137 (N_1137,N_682,N_851);
and U1138 (N_1138,N_716,N_751);
or U1139 (N_1139,N_765,N_856);
nor U1140 (N_1140,N_592,N_928);
nand U1141 (N_1141,N_874,N_771);
and U1142 (N_1142,N_622,N_798);
nand U1143 (N_1143,N_718,N_894);
or U1144 (N_1144,N_881,N_650);
and U1145 (N_1145,N_598,N_620);
and U1146 (N_1146,N_954,N_638);
nor U1147 (N_1147,N_879,N_827);
xor U1148 (N_1148,N_667,N_563);
and U1149 (N_1149,N_967,N_890);
and U1150 (N_1150,N_947,N_811);
and U1151 (N_1151,N_976,N_584);
nand U1152 (N_1152,N_539,N_988);
nor U1153 (N_1153,N_953,N_971);
and U1154 (N_1154,N_942,N_741);
and U1155 (N_1155,N_968,N_645);
and U1156 (N_1156,N_623,N_502);
nor U1157 (N_1157,N_677,N_805);
nand U1158 (N_1158,N_867,N_895);
nand U1159 (N_1159,N_569,N_903);
nand U1160 (N_1160,N_604,N_659);
and U1161 (N_1161,N_576,N_729);
and U1162 (N_1162,N_521,N_628);
xnor U1163 (N_1163,N_513,N_656);
nand U1164 (N_1164,N_616,N_712);
or U1165 (N_1165,N_671,N_753);
nand U1166 (N_1166,N_607,N_959);
nor U1167 (N_1167,N_961,N_636);
nand U1168 (N_1168,N_884,N_864);
nor U1169 (N_1169,N_595,N_794);
nand U1170 (N_1170,N_635,N_734);
nor U1171 (N_1171,N_949,N_777);
and U1172 (N_1172,N_542,N_611);
xnor U1173 (N_1173,N_723,N_640);
or U1174 (N_1174,N_657,N_602);
or U1175 (N_1175,N_647,N_911);
and U1176 (N_1176,N_662,N_899);
or U1177 (N_1177,N_582,N_991);
nor U1178 (N_1178,N_614,N_646);
nor U1179 (N_1179,N_759,N_747);
and U1180 (N_1180,N_527,N_544);
nor U1181 (N_1181,N_829,N_529);
and U1182 (N_1182,N_696,N_837);
nor U1183 (N_1183,N_900,N_706);
and U1184 (N_1184,N_783,N_679);
or U1185 (N_1185,N_634,N_532);
nand U1186 (N_1186,N_860,N_691);
and U1187 (N_1187,N_927,N_519);
and U1188 (N_1188,N_809,N_566);
nor U1189 (N_1189,N_969,N_744);
nand U1190 (N_1190,N_802,N_639);
or U1191 (N_1191,N_730,N_724);
or U1192 (N_1192,N_697,N_951);
nand U1193 (N_1193,N_919,N_619);
xnor U1194 (N_1194,N_666,N_850);
xnor U1195 (N_1195,N_760,N_605);
nor U1196 (N_1196,N_848,N_865);
nor U1197 (N_1197,N_686,N_962);
xnor U1198 (N_1198,N_778,N_996);
nand U1199 (N_1199,N_556,N_570);
nand U1200 (N_1200,N_609,N_826);
nand U1201 (N_1201,N_631,N_757);
nor U1202 (N_1202,N_558,N_547);
nor U1203 (N_1203,N_977,N_907);
nor U1204 (N_1204,N_612,N_565);
and U1205 (N_1205,N_557,N_888);
and U1206 (N_1206,N_936,N_870);
and U1207 (N_1207,N_511,N_889);
nand U1208 (N_1208,N_769,N_960);
or U1209 (N_1209,N_652,N_799);
xor U1210 (N_1210,N_795,N_571);
nand U1211 (N_1211,N_648,N_546);
and U1212 (N_1212,N_818,N_586);
or U1213 (N_1213,N_510,N_589);
nor U1214 (N_1214,N_981,N_945);
or U1215 (N_1215,N_938,N_588);
nand U1216 (N_1216,N_834,N_807);
and U1217 (N_1217,N_882,N_973);
and U1218 (N_1218,N_909,N_725);
and U1219 (N_1219,N_523,N_858);
nor U1220 (N_1220,N_999,N_526);
nor U1221 (N_1221,N_507,N_833);
or U1222 (N_1222,N_721,N_655);
or U1223 (N_1223,N_538,N_618);
or U1224 (N_1224,N_573,N_668);
nand U1225 (N_1225,N_709,N_965);
nand U1226 (N_1226,N_680,N_551);
and U1227 (N_1227,N_559,N_990);
nor U1228 (N_1228,N_825,N_886);
nand U1229 (N_1229,N_862,N_665);
and U1230 (N_1230,N_898,N_549);
or U1231 (N_1231,N_669,N_937);
xnor U1232 (N_1232,N_830,N_788);
nor U1233 (N_1233,N_845,N_985);
and U1234 (N_1234,N_792,N_533);
xor U1235 (N_1235,N_743,N_528);
nand U1236 (N_1236,N_505,N_812);
xor U1237 (N_1237,N_683,N_537);
and U1238 (N_1238,N_621,N_681);
nand U1239 (N_1239,N_925,N_957);
nor U1240 (N_1240,N_685,N_701);
nor U1241 (N_1241,N_921,N_880);
or U1242 (N_1242,N_824,N_929);
and U1243 (N_1243,N_541,N_887);
or U1244 (N_1244,N_574,N_940);
and U1245 (N_1245,N_776,N_572);
or U1246 (N_1246,N_972,N_983);
or U1247 (N_1247,N_980,N_564);
nand U1248 (N_1248,N_714,N_910);
nor U1249 (N_1249,N_853,N_838);
nand U1250 (N_1250,N_955,N_585);
nor U1251 (N_1251,N_776,N_781);
nor U1252 (N_1252,N_967,N_704);
xnor U1253 (N_1253,N_814,N_835);
nand U1254 (N_1254,N_853,N_612);
nand U1255 (N_1255,N_990,N_594);
or U1256 (N_1256,N_881,N_730);
nand U1257 (N_1257,N_809,N_642);
nand U1258 (N_1258,N_533,N_821);
or U1259 (N_1259,N_763,N_516);
nand U1260 (N_1260,N_569,N_616);
or U1261 (N_1261,N_783,N_616);
and U1262 (N_1262,N_762,N_645);
and U1263 (N_1263,N_992,N_682);
nor U1264 (N_1264,N_711,N_616);
nand U1265 (N_1265,N_558,N_660);
nand U1266 (N_1266,N_895,N_646);
or U1267 (N_1267,N_706,N_898);
nand U1268 (N_1268,N_871,N_770);
nor U1269 (N_1269,N_568,N_528);
and U1270 (N_1270,N_769,N_940);
nand U1271 (N_1271,N_749,N_796);
xnor U1272 (N_1272,N_635,N_744);
nor U1273 (N_1273,N_679,N_535);
nand U1274 (N_1274,N_869,N_899);
nor U1275 (N_1275,N_707,N_972);
nand U1276 (N_1276,N_708,N_898);
or U1277 (N_1277,N_643,N_500);
and U1278 (N_1278,N_517,N_988);
nand U1279 (N_1279,N_524,N_552);
or U1280 (N_1280,N_882,N_946);
and U1281 (N_1281,N_794,N_834);
and U1282 (N_1282,N_968,N_818);
or U1283 (N_1283,N_946,N_727);
and U1284 (N_1284,N_691,N_734);
or U1285 (N_1285,N_697,N_963);
nor U1286 (N_1286,N_619,N_887);
and U1287 (N_1287,N_822,N_543);
nor U1288 (N_1288,N_935,N_693);
nand U1289 (N_1289,N_854,N_692);
nand U1290 (N_1290,N_968,N_889);
or U1291 (N_1291,N_909,N_867);
nand U1292 (N_1292,N_712,N_536);
and U1293 (N_1293,N_560,N_786);
nand U1294 (N_1294,N_588,N_942);
and U1295 (N_1295,N_998,N_659);
xnor U1296 (N_1296,N_993,N_623);
or U1297 (N_1297,N_975,N_762);
and U1298 (N_1298,N_769,N_677);
xnor U1299 (N_1299,N_571,N_945);
nor U1300 (N_1300,N_693,N_704);
nand U1301 (N_1301,N_569,N_868);
xor U1302 (N_1302,N_859,N_906);
nand U1303 (N_1303,N_599,N_671);
and U1304 (N_1304,N_537,N_952);
or U1305 (N_1305,N_665,N_913);
nand U1306 (N_1306,N_916,N_967);
nor U1307 (N_1307,N_604,N_713);
nor U1308 (N_1308,N_613,N_636);
or U1309 (N_1309,N_623,N_873);
nand U1310 (N_1310,N_670,N_634);
nand U1311 (N_1311,N_580,N_614);
or U1312 (N_1312,N_843,N_699);
nand U1313 (N_1313,N_986,N_960);
nor U1314 (N_1314,N_781,N_543);
and U1315 (N_1315,N_845,N_679);
nand U1316 (N_1316,N_970,N_748);
or U1317 (N_1317,N_548,N_897);
or U1318 (N_1318,N_678,N_568);
nor U1319 (N_1319,N_543,N_679);
nand U1320 (N_1320,N_950,N_562);
nor U1321 (N_1321,N_503,N_639);
or U1322 (N_1322,N_983,N_916);
and U1323 (N_1323,N_679,N_741);
xnor U1324 (N_1324,N_994,N_577);
and U1325 (N_1325,N_921,N_840);
nand U1326 (N_1326,N_588,N_829);
or U1327 (N_1327,N_757,N_984);
xor U1328 (N_1328,N_810,N_864);
nand U1329 (N_1329,N_855,N_716);
nor U1330 (N_1330,N_762,N_763);
or U1331 (N_1331,N_847,N_600);
and U1332 (N_1332,N_592,N_528);
nand U1333 (N_1333,N_884,N_535);
or U1334 (N_1334,N_985,N_983);
nand U1335 (N_1335,N_959,N_874);
xnor U1336 (N_1336,N_530,N_671);
nor U1337 (N_1337,N_642,N_910);
xnor U1338 (N_1338,N_684,N_992);
and U1339 (N_1339,N_950,N_801);
and U1340 (N_1340,N_906,N_712);
nor U1341 (N_1341,N_682,N_650);
nand U1342 (N_1342,N_681,N_528);
nor U1343 (N_1343,N_819,N_806);
nor U1344 (N_1344,N_955,N_758);
nor U1345 (N_1345,N_527,N_805);
nor U1346 (N_1346,N_760,N_878);
and U1347 (N_1347,N_638,N_634);
nor U1348 (N_1348,N_653,N_867);
nor U1349 (N_1349,N_894,N_856);
nand U1350 (N_1350,N_874,N_581);
nand U1351 (N_1351,N_829,N_676);
or U1352 (N_1352,N_905,N_935);
or U1353 (N_1353,N_504,N_587);
and U1354 (N_1354,N_828,N_590);
or U1355 (N_1355,N_633,N_609);
and U1356 (N_1356,N_935,N_511);
nand U1357 (N_1357,N_815,N_554);
xnor U1358 (N_1358,N_978,N_601);
nand U1359 (N_1359,N_982,N_569);
nand U1360 (N_1360,N_641,N_504);
xnor U1361 (N_1361,N_504,N_878);
or U1362 (N_1362,N_518,N_563);
or U1363 (N_1363,N_909,N_745);
nand U1364 (N_1364,N_898,N_751);
or U1365 (N_1365,N_983,N_890);
and U1366 (N_1366,N_616,N_571);
and U1367 (N_1367,N_735,N_765);
nor U1368 (N_1368,N_739,N_543);
nand U1369 (N_1369,N_687,N_640);
nor U1370 (N_1370,N_856,N_846);
or U1371 (N_1371,N_731,N_837);
nor U1372 (N_1372,N_722,N_776);
nand U1373 (N_1373,N_748,N_782);
or U1374 (N_1374,N_681,N_976);
xnor U1375 (N_1375,N_924,N_876);
nand U1376 (N_1376,N_546,N_525);
nand U1377 (N_1377,N_994,N_688);
nand U1378 (N_1378,N_533,N_801);
nor U1379 (N_1379,N_520,N_833);
nor U1380 (N_1380,N_595,N_911);
xor U1381 (N_1381,N_809,N_652);
nand U1382 (N_1382,N_957,N_941);
nand U1383 (N_1383,N_833,N_676);
xnor U1384 (N_1384,N_553,N_907);
and U1385 (N_1385,N_611,N_595);
and U1386 (N_1386,N_940,N_507);
or U1387 (N_1387,N_899,N_586);
nor U1388 (N_1388,N_737,N_625);
and U1389 (N_1389,N_738,N_769);
and U1390 (N_1390,N_870,N_745);
nand U1391 (N_1391,N_577,N_829);
nand U1392 (N_1392,N_755,N_734);
xor U1393 (N_1393,N_603,N_802);
nand U1394 (N_1394,N_547,N_500);
nand U1395 (N_1395,N_697,N_977);
nor U1396 (N_1396,N_748,N_729);
nand U1397 (N_1397,N_552,N_843);
or U1398 (N_1398,N_627,N_675);
nand U1399 (N_1399,N_508,N_924);
nor U1400 (N_1400,N_604,N_594);
nor U1401 (N_1401,N_907,N_847);
or U1402 (N_1402,N_559,N_966);
or U1403 (N_1403,N_620,N_903);
nor U1404 (N_1404,N_556,N_916);
nor U1405 (N_1405,N_786,N_605);
nand U1406 (N_1406,N_634,N_749);
nor U1407 (N_1407,N_537,N_539);
or U1408 (N_1408,N_966,N_629);
nand U1409 (N_1409,N_897,N_531);
nor U1410 (N_1410,N_586,N_677);
or U1411 (N_1411,N_797,N_689);
nor U1412 (N_1412,N_659,N_826);
or U1413 (N_1413,N_535,N_709);
nor U1414 (N_1414,N_935,N_770);
or U1415 (N_1415,N_795,N_836);
nor U1416 (N_1416,N_709,N_773);
nand U1417 (N_1417,N_866,N_864);
and U1418 (N_1418,N_777,N_711);
and U1419 (N_1419,N_689,N_747);
nand U1420 (N_1420,N_771,N_553);
or U1421 (N_1421,N_988,N_601);
nand U1422 (N_1422,N_638,N_997);
and U1423 (N_1423,N_885,N_882);
xor U1424 (N_1424,N_910,N_997);
nor U1425 (N_1425,N_884,N_613);
nand U1426 (N_1426,N_525,N_702);
nand U1427 (N_1427,N_855,N_691);
or U1428 (N_1428,N_522,N_600);
or U1429 (N_1429,N_557,N_794);
or U1430 (N_1430,N_729,N_608);
xor U1431 (N_1431,N_705,N_631);
nor U1432 (N_1432,N_693,N_595);
nor U1433 (N_1433,N_606,N_684);
and U1434 (N_1434,N_900,N_855);
nand U1435 (N_1435,N_712,N_716);
nor U1436 (N_1436,N_551,N_719);
and U1437 (N_1437,N_759,N_731);
nand U1438 (N_1438,N_797,N_770);
nand U1439 (N_1439,N_948,N_629);
nor U1440 (N_1440,N_613,N_937);
nand U1441 (N_1441,N_952,N_788);
nor U1442 (N_1442,N_724,N_673);
nand U1443 (N_1443,N_818,N_977);
nand U1444 (N_1444,N_775,N_645);
or U1445 (N_1445,N_698,N_674);
nor U1446 (N_1446,N_812,N_704);
nor U1447 (N_1447,N_998,N_865);
xnor U1448 (N_1448,N_666,N_852);
nor U1449 (N_1449,N_792,N_503);
or U1450 (N_1450,N_936,N_938);
nor U1451 (N_1451,N_853,N_947);
and U1452 (N_1452,N_972,N_684);
and U1453 (N_1453,N_998,N_534);
nand U1454 (N_1454,N_696,N_717);
or U1455 (N_1455,N_637,N_981);
nor U1456 (N_1456,N_775,N_647);
and U1457 (N_1457,N_507,N_597);
nor U1458 (N_1458,N_932,N_884);
nor U1459 (N_1459,N_919,N_587);
or U1460 (N_1460,N_853,N_801);
nor U1461 (N_1461,N_990,N_945);
xor U1462 (N_1462,N_533,N_532);
nand U1463 (N_1463,N_830,N_701);
or U1464 (N_1464,N_982,N_685);
nand U1465 (N_1465,N_749,N_651);
nand U1466 (N_1466,N_732,N_722);
nand U1467 (N_1467,N_828,N_786);
and U1468 (N_1468,N_746,N_931);
and U1469 (N_1469,N_670,N_659);
and U1470 (N_1470,N_509,N_965);
and U1471 (N_1471,N_931,N_536);
or U1472 (N_1472,N_978,N_906);
and U1473 (N_1473,N_675,N_552);
or U1474 (N_1474,N_779,N_644);
or U1475 (N_1475,N_763,N_594);
and U1476 (N_1476,N_530,N_808);
and U1477 (N_1477,N_749,N_550);
or U1478 (N_1478,N_926,N_952);
xnor U1479 (N_1479,N_862,N_777);
nand U1480 (N_1480,N_725,N_815);
or U1481 (N_1481,N_908,N_612);
and U1482 (N_1482,N_924,N_826);
and U1483 (N_1483,N_884,N_963);
and U1484 (N_1484,N_905,N_964);
nand U1485 (N_1485,N_547,N_518);
or U1486 (N_1486,N_958,N_799);
nand U1487 (N_1487,N_500,N_679);
or U1488 (N_1488,N_661,N_573);
nor U1489 (N_1489,N_757,N_855);
and U1490 (N_1490,N_821,N_608);
and U1491 (N_1491,N_783,N_994);
or U1492 (N_1492,N_536,N_685);
xnor U1493 (N_1493,N_761,N_856);
and U1494 (N_1494,N_822,N_729);
or U1495 (N_1495,N_954,N_788);
nor U1496 (N_1496,N_829,N_718);
and U1497 (N_1497,N_712,N_731);
nand U1498 (N_1498,N_990,N_644);
or U1499 (N_1499,N_908,N_995);
and U1500 (N_1500,N_1330,N_1309);
or U1501 (N_1501,N_1324,N_1406);
nor U1502 (N_1502,N_1062,N_1233);
or U1503 (N_1503,N_1241,N_1442);
nand U1504 (N_1504,N_1074,N_1011);
and U1505 (N_1505,N_1432,N_1239);
or U1506 (N_1506,N_1351,N_1075);
nor U1507 (N_1507,N_1322,N_1262);
nor U1508 (N_1508,N_1169,N_1146);
or U1509 (N_1509,N_1257,N_1336);
or U1510 (N_1510,N_1467,N_1054);
xor U1511 (N_1511,N_1398,N_1460);
xnor U1512 (N_1512,N_1323,N_1431);
or U1513 (N_1513,N_1109,N_1219);
xor U1514 (N_1514,N_1349,N_1188);
and U1515 (N_1515,N_1053,N_1279);
nor U1516 (N_1516,N_1457,N_1270);
and U1517 (N_1517,N_1275,N_1373);
nand U1518 (N_1518,N_1212,N_1413);
nand U1519 (N_1519,N_1091,N_1113);
nor U1520 (N_1520,N_1181,N_1415);
or U1521 (N_1521,N_1229,N_1046);
nor U1522 (N_1522,N_1186,N_1447);
or U1523 (N_1523,N_1087,N_1428);
nand U1524 (N_1524,N_1244,N_1020);
or U1525 (N_1525,N_1476,N_1164);
or U1526 (N_1526,N_1409,N_1190);
nand U1527 (N_1527,N_1217,N_1385);
or U1528 (N_1528,N_1490,N_1359);
nor U1529 (N_1529,N_1363,N_1289);
and U1530 (N_1530,N_1080,N_1214);
and U1531 (N_1531,N_1378,N_1434);
nor U1532 (N_1532,N_1086,N_1176);
and U1533 (N_1533,N_1374,N_1215);
and U1534 (N_1534,N_1421,N_1228);
nand U1535 (N_1535,N_1450,N_1313);
nor U1536 (N_1536,N_1052,N_1369);
nor U1537 (N_1537,N_1366,N_1499);
nand U1538 (N_1538,N_1397,N_1250);
nor U1539 (N_1539,N_1041,N_1165);
or U1540 (N_1540,N_1106,N_1225);
or U1541 (N_1541,N_1193,N_1491);
nand U1542 (N_1542,N_1222,N_1364);
and U1543 (N_1543,N_1158,N_1178);
or U1544 (N_1544,N_1472,N_1372);
nor U1545 (N_1545,N_1043,N_1051);
and U1546 (N_1546,N_1458,N_1353);
or U1547 (N_1547,N_1312,N_1333);
nand U1548 (N_1548,N_1145,N_1267);
nand U1549 (N_1549,N_1402,N_1037);
nor U1550 (N_1550,N_1433,N_1104);
or U1551 (N_1551,N_1057,N_1039);
or U1552 (N_1552,N_1329,N_1185);
or U1553 (N_1553,N_1357,N_1276);
and U1554 (N_1554,N_1069,N_1101);
and U1555 (N_1555,N_1471,N_1187);
or U1556 (N_1556,N_1288,N_1355);
and U1557 (N_1557,N_1044,N_1105);
or U1558 (N_1558,N_1390,N_1002);
nand U1559 (N_1559,N_1059,N_1419);
nand U1560 (N_1560,N_1412,N_1466);
nand U1561 (N_1561,N_1138,N_1142);
nor U1562 (N_1562,N_1468,N_1456);
nor U1563 (N_1563,N_1108,N_1480);
nand U1564 (N_1564,N_1337,N_1157);
nand U1565 (N_1565,N_1098,N_1026);
and U1566 (N_1566,N_1110,N_1301);
nor U1567 (N_1567,N_1266,N_1114);
and U1568 (N_1568,N_1271,N_1141);
and U1569 (N_1569,N_1498,N_1201);
nor U1570 (N_1570,N_1200,N_1341);
and U1571 (N_1571,N_1277,N_1462);
nor U1572 (N_1572,N_1208,N_1064);
or U1573 (N_1573,N_1345,N_1029);
and U1574 (N_1574,N_1487,N_1430);
nor U1575 (N_1575,N_1386,N_1420);
nor U1576 (N_1576,N_1206,N_1147);
and U1577 (N_1577,N_1417,N_1172);
nor U1578 (N_1578,N_1038,N_1151);
nor U1579 (N_1579,N_1122,N_1081);
nand U1580 (N_1580,N_1300,N_1477);
or U1581 (N_1581,N_1066,N_1166);
nor U1582 (N_1582,N_1231,N_1482);
or U1583 (N_1583,N_1036,N_1112);
nand U1584 (N_1584,N_1048,N_1015);
or U1585 (N_1585,N_1174,N_1342);
nor U1586 (N_1586,N_1168,N_1137);
xnor U1587 (N_1587,N_1092,N_1023);
nand U1588 (N_1588,N_1278,N_1116);
nand U1589 (N_1589,N_1311,N_1260);
or U1590 (N_1590,N_1042,N_1383);
xor U1591 (N_1591,N_1132,N_1263);
and U1592 (N_1592,N_1177,N_1014);
nand U1593 (N_1593,N_1354,N_1134);
nor U1594 (N_1594,N_1230,N_1405);
nand U1595 (N_1595,N_1247,N_1461);
nand U1596 (N_1596,N_1148,N_1088);
or U1597 (N_1597,N_1005,N_1096);
nor U1598 (N_1598,N_1484,N_1140);
nor U1599 (N_1599,N_1454,N_1416);
nand U1600 (N_1600,N_1310,N_1259);
nor U1601 (N_1601,N_1258,N_1335);
or U1602 (N_1602,N_1334,N_1326);
nor U1603 (N_1603,N_1221,N_1189);
and U1604 (N_1604,N_1006,N_1443);
nand U1605 (N_1605,N_1360,N_1197);
or U1606 (N_1606,N_1426,N_1017);
nor U1607 (N_1607,N_1389,N_1379);
xnor U1608 (N_1608,N_1317,N_1045);
nor U1609 (N_1609,N_1242,N_1209);
or U1610 (N_1610,N_1124,N_1024);
or U1611 (N_1611,N_1403,N_1144);
nand U1612 (N_1612,N_1294,N_1459);
xnor U1613 (N_1613,N_1479,N_1131);
or U1614 (N_1614,N_1129,N_1035);
or U1615 (N_1615,N_1286,N_1224);
nand U1616 (N_1616,N_1365,N_1440);
and U1617 (N_1617,N_1202,N_1232);
and U1618 (N_1618,N_1380,N_1469);
and U1619 (N_1619,N_1033,N_1155);
xor U1620 (N_1620,N_1444,N_1115);
nand U1621 (N_1621,N_1400,N_1465);
xnor U1622 (N_1622,N_1156,N_1285);
nand U1623 (N_1623,N_1424,N_1305);
and U1624 (N_1624,N_1414,N_1304);
nor U1625 (N_1625,N_1295,N_1254);
nor U1626 (N_1626,N_1475,N_1198);
nand U1627 (N_1627,N_1255,N_1003);
or U1628 (N_1628,N_1143,N_1159);
or U1629 (N_1629,N_1411,N_1248);
nand U1630 (N_1630,N_1325,N_1287);
or U1631 (N_1631,N_1094,N_1371);
or U1632 (N_1632,N_1281,N_1030);
or U1633 (N_1633,N_1246,N_1418);
xnor U1634 (N_1634,N_1284,N_1034);
and U1635 (N_1635,N_1216,N_1280);
nor U1636 (N_1636,N_1089,N_1394);
xnor U1637 (N_1637,N_1265,N_1408);
nor U1638 (N_1638,N_1382,N_1436);
or U1639 (N_1639,N_1210,N_1404);
nor U1640 (N_1640,N_1302,N_1211);
or U1641 (N_1641,N_1347,N_1226);
nand U1642 (N_1642,N_1021,N_1455);
or U1643 (N_1643,N_1422,N_1274);
nor U1644 (N_1644,N_1388,N_1474);
nand U1645 (N_1645,N_1207,N_1316);
or U1646 (N_1646,N_1032,N_1031);
nand U1647 (N_1647,N_1249,N_1154);
nand U1648 (N_1648,N_1387,N_1435);
nand U1649 (N_1649,N_1119,N_1152);
nand U1650 (N_1650,N_1162,N_1047);
nor U1651 (N_1651,N_1494,N_1150);
and U1652 (N_1652,N_1204,N_1290);
xor U1653 (N_1653,N_1127,N_1315);
and U1654 (N_1654,N_1196,N_1478);
nand U1655 (N_1655,N_1410,N_1481);
xnor U1656 (N_1656,N_1076,N_1245);
nor U1657 (N_1657,N_1027,N_1083);
and U1658 (N_1658,N_1299,N_1049);
nand U1659 (N_1659,N_1437,N_1375);
nor U1660 (N_1660,N_1077,N_1446);
nand U1661 (N_1661,N_1384,N_1213);
nand U1662 (N_1662,N_1283,N_1269);
nand U1663 (N_1663,N_1488,N_1019);
nor U1664 (N_1664,N_1327,N_1451);
and U1665 (N_1665,N_1438,N_1293);
nand U1666 (N_1666,N_1332,N_1040);
nor U1667 (N_1667,N_1381,N_1028);
and U1668 (N_1668,N_1370,N_1180);
nor U1669 (N_1669,N_1120,N_1439);
nand U1670 (N_1670,N_1307,N_1130);
nor U1671 (N_1671,N_1022,N_1393);
or U1672 (N_1672,N_1448,N_1073);
or U1673 (N_1673,N_1067,N_1427);
or U1674 (N_1674,N_1182,N_1055);
nand U1675 (N_1675,N_1203,N_1356);
nand U1676 (N_1676,N_1399,N_1496);
xnor U1677 (N_1677,N_1012,N_1179);
and U1678 (N_1678,N_1167,N_1252);
nand U1679 (N_1679,N_1194,N_1061);
nand U1680 (N_1680,N_1236,N_1346);
or U1681 (N_1681,N_1331,N_1063);
xor U1682 (N_1682,N_1396,N_1340);
or U1683 (N_1683,N_1493,N_1100);
or U1684 (N_1684,N_1362,N_1093);
and U1685 (N_1685,N_1199,N_1161);
and U1686 (N_1686,N_1306,N_1321);
and U1687 (N_1687,N_1358,N_1483);
and U1688 (N_1688,N_1445,N_1060);
xor U1689 (N_1689,N_1495,N_1025);
nor U1690 (N_1690,N_1205,N_1253);
and U1691 (N_1691,N_1234,N_1352);
nor U1692 (N_1692,N_1084,N_1183);
and U1693 (N_1693,N_1010,N_1001);
or U1694 (N_1694,N_1135,N_1298);
and U1695 (N_1695,N_1308,N_1125);
nor U1696 (N_1696,N_1121,N_1065);
and U1697 (N_1697,N_1184,N_1441);
nor U1698 (N_1698,N_1009,N_1268);
xnor U1699 (N_1699,N_1272,N_1401);
nor U1700 (N_1700,N_1079,N_1473);
nor U1701 (N_1701,N_1292,N_1078);
nor U1702 (N_1702,N_1082,N_1103);
nand U1703 (N_1703,N_1395,N_1238);
or U1704 (N_1704,N_1470,N_1016);
and U1705 (N_1705,N_1220,N_1175);
or U1706 (N_1706,N_1218,N_1282);
nand U1707 (N_1707,N_1452,N_1492);
nand U1708 (N_1708,N_1343,N_1068);
or U1709 (N_1709,N_1377,N_1264);
or U1710 (N_1710,N_1489,N_1391);
or U1711 (N_1711,N_1139,N_1171);
and U1712 (N_1712,N_1071,N_1425);
nand U1713 (N_1713,N_1173,N_1107);
or U1714 (N_1714,N_1338,N_1118);
nand U1715 (N_1715,N_1235,N_1133);
nand U1716 (N_1716,N_1018,N_1123);
nand U1717 (N_1717,N_1339,N_1243);
or U1718 (N_1718,N_1297,N_1007);
or U1719 (N_1719,N_1485,N_1237);
and U1720 (N_1720,N_1256,N_1102);
and U1721 (N_1721,N_1170,N_1111);
nand U1722 (N_1722,N_1128,N_1085);
or U1723 (N_1723,N_1350,N_1097);
xor U1724 (N_1724,N_1008,N_1273);
nor U1725 (N_1725,N_1251,N_1429);
or U1726 (N_1726,N_1303,N_1195);
and U1727 (N_1727,N_1497,N_1126);
or U1728 (N_1728,N_1348,N_1328);
or U1729 (N_1729,N_1240,N_1227);
nand U1730 (N_1730,N_1000,N_1072);
or U1731 (N_1731,N_1058,N_1191);
or U1732 (N_1732,N_1149,N_1319);
nor U1733 (N_1733,N_1423,N_1013);
or U1734 (N_1734,N_1392,N_1070);
and U1735 (N_1735,N_1095,N_1160);
and U1736 (N_1736,N_1361,N_1368);
or U1737 (N_1737,N_1136,N_1463);
nand U1738 (N_1738,N_1344,N_1314);
or U1739 (N_1739,N_1153,N_1192);
and U1740 (N_1740,N_1376,N_1291);
nand U1741 (N_1741,N_1223,N_1453);
xor U1742 (N_1742,N_1486,N_1099);
nand U1743 (N_1743,N_1464,N_1449);
or U1744 (N_1744,N_1261,N_1056);
and U1745 (N_1745,N_1090,N_1050);
nand U1746 (N_1746,N_1004,N_1296);
nand U1747 (N_1747,N_1117,N_1320);
or U1748 (N_1748,N_1163,N_1407);
and U1749 (N_1749,N_1318,N_1367);
or U1750 (N_1750,N_1111,N_1301);
nand U1751 (N_1751,N_1426,N_1305);
nor U1752 (N_1752,N_1041,N_1287);
nor U1753 (N_1753,N_1186,N_1400);
nor U1754 (N_1754,N_1167,N_1336);
nor U1755 (N_1755,N_1127,N_1354);
nor U1756 (N_1756,N_1344,N_1255);
and U1757 (N_1757,N_1336,N_1243);
xor U1758 (N_1758,N_1037,N_1436);
nand U1759 (N_1759,N_1435,N_1197);
nand U1760 (N_1760,N_1242,N_1189);
and U1761 (N_1761,N_1384,N_1175);
nand U1762 (N_1762,N_1495,N_1464);
and U1763 (N_1763,N_1199,N_1377);
nor U1764 (N_1764,N_1451,N_1361);
and U1765 (N_1765,N_1427,N_1264);
or U1766 (N_1766,N_1301,N_1083);
xnor U1767 (N_1767,N_1494,N_1002);
nor U1768 (N_1768,N_1220,N_1181);
nand U1769 (N_1769,N_1196,N_1203);
or U1770 (N_1770,N_1114,N_1039);
and U1771 (N_1771,N_1318,N_1335);
nor U1772 (N_1772,N_1243,N_1315);
or U1773 (N_1773,N_1360,N_1276);
and U1774 (N_1774,N_1151,N_1220);
nand U1775 (N_1775,N_1231,N_1131);
and U1776 (N_1776,N_1074,N_1114);
nor U1777 (N_1777,N_1306,N_1341);
and U1778 (N_1778,N_1468,N_1060);
nor U1779 (N_1779,N_1280,N_1462);
and U1780 (N_1780,N_1075,N_1190);
nor U1781 (N_1781,N_1263,N_1186);
xnor U1782 (N_1782,N_1253,N_1140);
or U1783 (N_1783,N_1160,N_1234);
and U1784 (N_1784,N_1313,N_1136);
and U1785 (N_1785,N_1113,N_1107);
or U1786 (N_1786,N_1202,N_1298);
nand U1787 (N_1787,N_1139,N_1311);
and U1788 (N_1788,N_1191,N_1407);
or U1789 (N_1789,N_1041,N_1079);
and U1790 (N_1790,N_1226,N_1296);
and U1791 (N_1791,N_1188,N_1252);
or U1792 (N_1792,N_1352,N_1235);
nor U1793 (N_1793,N_1433,N_1150);
nor U1794 (N_1794,N_1324,N_1158);
and U1795 (N_1795,N_1392,N_1065);
or U1796 (N_1796,N_1169,N_1379);
and U1797 (N_1797,N_1136,N_1380);
nor U1798 (N_1798,N_1355,N_1163);
nor U1799 (N_1799,N_1451,N_1085);
or U1800 (N_1800,N_1282,N_1255);
nand U1801 (N_1801,N_1007,N_1455);
or U1802 (N_1802,N_1471,N_1220);
nand U1803 (N_1803,N_1436,N_1367);
nor U1804 (N_1804,N_1029,N_1330);
or U1805 (N_1805,N_1174,N_1268);
nand U1806 (N_1806,N_1387,N_1088);
or U1807 (N_1807,N_1176,N_1268);
and U1808 (N_1808,N_1295,N_1284);
nor U1809 (N_1809,N_1074,N_1323);
xnor U1810 (N_1810,N_1002,N_1490);
nor U1811 (N_1811,N_1312,N_1396);
nand U1812 (N_1812,N_1075,N_1172);
and U1813 (N_1813,N_1335,N_1344);
or U1814 (N_1814,N_1228,N_1067);
nor U1815 (N_1815,N_1400,N_1298);
and U1816 (N_1816,N_1001,N_1147);
or U1817 (N_1817,N_1009,N_1168);
and U1818 (N_1818,N_1202,N_1337);
and U1819 (N_1819,N_1294,N_1131);
and U1820 (N_1820,N_1232,N_1471);
nand U1821 (N_1821,N_1466,N_1408);
nor U1822 (N_1822,N_1326,N_1073);
xnor U1823 (N_1823,N_1429,N_1323);
nand U1824 (N_1824,N_1318,N_1279);
xnor U1825 (N_1825,N_1299,N_1398);
or U1826 (N_1826,N_1108,N_1120);
nor U1827 (N_1827,N_1414,N_1229);
nand U1828 (N_1828,N_1311,N_1449);
nor U1829 (N_1829,N_1215,N_1105);
and U1830 (N_1830,N_1488,N_1482);
and U1831 (N_1831,N_1398,N_1441);
or U1832 (N_1832,N_1081,N_1340);
nor U1833 (N_1833,N_1425,N_1222);
nor U1834 (N_1834,N_1441,N_1193);
nand U1835 (N_1835,N_1330,N_1328);
nor U1836 (N_1836,N_1145,N_1363);
and U1837 (N_1837,N_1288,N_1364);
and U1838 (N_1838,N_1396,N_1175);
xnor U1839 (N_1839,N_1299,N_1287);
nand U1840 (N_1840,N_1384,N_1046);
or U1841 (N_1841,N_1489,N_1479);
nor U1842 (N_1842,N_1236,N_1294);
nor U1843 (N_1843,N_1033,N_1355);
nand U1844 (N_1844,N_1132,N_1400);
and U1845 (N_1845,N_1074,N_1280);
and U1846 (N_1846,N_1008,N_1490);
nor U1847 (N_1847,N_1016,N_1386);
nand U1848 (N_1848,N_1436,N_1300);
nand U1849 (N_1849,N_1409,N_1132);
nor U1850 (N_1850,N_1208,N_1187);
nor U1851 (N_1851,N_1464,N_1036);
and U1852 (N_1852,N_1090,N_1048);
nor U1853 (N_1853,N_1220,N_1184);
or U1854 (N_1854,N_1006,N_1286);
and U1855 (N_1855,N_1067,N_1153);
nor U1856 (N_1856,N_1030,N_1200);
xor U1857 (N_1857,N_1289,N_1031);
and U1858 (N_1858,N_1087,N_1134);
or U1859 (N_1859,N_1348,N_1139);
and U1860 (N_1860,N_1336,N_1376);
nand U1861 (N_1861,N_1102,N_1056);
or U1862 (N_1862,N_1297,N_1092);
or U1863 (N_1863,N_1316,N_1457);
xnor U1864 (N_1864,N_1120,N_1139);
nor U1865 (N_1865,N_1214,N_1319);
or U1866 (N_1866,N_1491,N_1234);
xor U1867 (N_1867,N_1041,N_1167);
and U1868 (N_1868,N_1245,N_1465);
or U1869 (N_1869,N_1365,N_1463);
or U1870 (N_1870,N_1043,N_1120);
and U1871 (N_1871,N_1201,N_1407);
nor U1872 (N_1872,N_1333,N_1462);
and U1873 (N_1873,N_1319,N_1318);
and U1874 (N_1874,N_1117,N_1423);
or U1875 (N_1875,N_1270,N_1427);
and U1876 (N_1876,N_1452,N_1221);
or U1877 (N_1877,N_1271,N_1390);
nand U1878 (N_1878,N_1095,N_1303);
nand U1879 (N_1879,N_1390,N_1208);
and U1880 (N_1880,N_1290,N_1086);
nor U1881 (N_1881,N_1150,N_1070);
and U1882 (N_1882,N_1484,N_1317);
nor U1883 (N_1883,N_1313,N_1093);
nor U1884 (N_1884,N_1453,N_1427);
nor U1885 (N_1885,N_1390,N_1138);
or U1886 (N_1886,N_1298,N_1146);
nand U1887 (N_1887,N_1369,N_1260);
xnor U1888 (N_1888,N_1150,N_1075);
nand U1889 (N_1889,N_1483,N_1169);
nand U1890 (N_1890,N_1492,N_1101);
nor U1891 (N_1891,N_1259,N_1066);
nor U1892 (N_1892,N_1220,N_1268);
xnor U1893 (N_1893,N_1189,N_1178);
nand U1894 (N_1894,N_1479,N_1449);
nor U1895 (N_1895,N_1268,N_1413);
nor U1896 (N_1896,N_1186,N_1260);
or U1897 (N_1897,N_1265,N_1404);
nor U1898 (N_1898,N_1076,N_1122);
or U1899 (N_1899,N_1225,N_1284);
and U1900 (N_1900,N_1230,N_1038);
and U1901 (N_1901,N_1093,N_1111);
and U1902 (N_1902,N_1098,N_1278);
nand U1903 (N_1903,N_1366,N_1158);
or U1904 (N_1904,N_1421,N_1063);
nor U1905 (N_1905,N_1389,N_1457);
nand U1906 (N_1906,N_1459,N_1284);
and U1907 (N_1907,N_1134,N_1404);
nand U1908 (N_1908,N_1229,N_1061);
nand U1909 (N_1909,N_1239,N_1317);
and U1910 (N_1910,N_1053,N_1473);
nor U1911 (N_1911,N_1277,N_1324);
nor U1912 (N_1912,N_1491,N_1023);
or U1913 (N_1913,N_1410,N_1094);
nand U1914 (N_1914,N_1016,N_1104);
and U1915 (N_1915,N_1135,N_1193);
and U1916 (N_1916,N_1391,N_1418);
and U1917 (N_1917,N_1250,N_1174);
nor U1918 (N_1918,N_1481,N_1208);
nand U1919 (N_1919,N_1095,N_1127);
xnor U1920 (N_1920,N_1206,N_1043);
and U1921 (N_1921,N_1066,N_1162);
and U1922 (N_1922,N_1072,N_1140);
and U1923 (N_1923,N_1033,N_1249);
xor U1924 (N_1924,N_1265,N_1120);
nor U1925 (N_1925,N_1346,N_1355);
and U1926 (N_1926,N_1167,N_1389);
xor U1927 (N_1927,N_1022,N_1469);
nand U1928 (N_1928,N_1044,N_1476);
and U1929 (N_1929,N_1432,N_1027);
nor U1930 (N_1930,N_1320,N_1285);
and U1931 (N_1931,N_1092,N_1159);
xnor U1932 (N_1932,N_1263,N_1007);
nor U1933 (N_1933,N_1321,N_1032);
and U1934 (N_1934,N_1211,N_1405);
or U1935 (N_1935,N_1190,N_1338);
or U1936 (N_1936,N_1246,N_1072);
or U1937 (N_1937,N_1436,N_1133);
and U1938 (N_1938,N_1105,N_1128);
or U1939 (N_1939,N_1335,N_1233);
nor U1940 (N_1940,N_1098,N_1047);
nand U1941 (N_1941,N_1175,N_1158);
xor U1942 (N_1942,N_1248,N_1323);
and U1943 (N_1943,N_1168,N_1240);
or U1944 (N_1944,N_1309,N_1153);
nor U1945 (N_1945,N_1154,N_1058);
nand U1946 (N_1946,N_1430,N_1136);
or U1947 (N_1947,N_1451,N_1059);
nand U1948 (N_1948,N_1015,N_1074);
and U1949 (N_1949,N_1409,N_1241);
and U1950 (N_1950,N_1485,N_1228);
or U1951 (N_1951,N_1156,N_1002);
and U1952 (N_1952,N_1016,N_1485);
or U1953 (N_1953,N_1050,N_1382);
and U1954 (N_1954,N_1264,N_1195);
nor U1955 (N_1955,N_1238,N_1390);
nor U1956 (N_1956,N_1262,N_1330);
and U1957 (N_1957,N_1172,N_1118);
nand U1958 (N_1958,N_1311,N_1397);
or U1959 (N_1959,N_1116,N_1313);
nand U1960 (N_1960,N_1079,N_1424);
nor U1961 (N_1961,N_1454,N_1089);
and U1962 (N_1962,N_1158,N_1425);
nand U1963 (N_1963,N_1003,N_1230);
or U1964 (N_1964,N_1143,N_1343);
nor U1965 (N_1965,N_1445,N_1188);
nand U1966 (N_1966,N_1301,N_1258);
or U1967 (N_1967,N_1430,N_1384);
and U1968 (N_1968,N_1240,N_1175);
or U1969 (N_1969,N_1288,N_1403);
and U1970 (N_1970,N_1385,N_1234);
nor U1971 (N_1971,N_1074,N_1109);
or U1972 (N_1972,N_1253,N_1098);
or U1973 (N_1973,N_1330,N_1260);
and U1974 (N_1974,N_1487,N_1093);
nand U1975 (N_1975,N_1064,N_1030);
or U1976 (N_1976,N_1485,N_1208);
and U1977 (N_1977,N_1016,N_1260);
nor U1978 (N_1978,N_1028,N_1177);
or U1979 (N_1979,N_1030,N_1469);
or U1980 (N_1980,N_1311,N_1467);
and U1981 (N_1981,N_1343,N_1318);
and U1982 (N_1982,N_1140,N_1483);
nand U1983 (N_1983,N_1235,N_1413);
nand U1984 (N_1984,N_1348,N_1469);
nand U1985 (N_1985,N_1133,N_1222);
or U1986 (N_1986,N_1493,N_1175);
nand U1987 (N_1987,N_1183,N_1004);
nand U1988 (N_1988,N_1376,N_1279);
nor U1989 (N_1989,N_1037,N_1492);
or U1990 (N_1990,N_1076,N_1261);
xor U1991 (N_1991,N_1410,N_1110);
xor U1992 (N_1992,N_1171,N_1096);
and U1993 (N_1993,N_1309,N_1366);
nor U1994 (N_1994,N_1324,N_1190);
or U1995 (N_1995,N_1117,N_1104);
nor U1996 (N_1996,N_1217,N_1243);
nand U1997 (N_1997,N_1321,N_1385);
nor U1998 (N_1998,N_1146,N_1149);
and U1999 (N_1999,N_1467,N_1412);
nand U2000 (N_2000,N_1660,N_1996);
or U2001 (N_2001,N_1775,N_1909);
xor U2002 (N_2002,N_1718,N_1702);
nor U2003 (N_2003,N_1872,N_1721);
nand U2004 (N_2004,N_1841,N_1740);
or U2005 (N_2005,N_1683,N_1539);
nand U2006 (N_2006,N_1679,N_1670);
and U2007 (N_2007,N_1845,N_1929);
or U2008 (N_2008,N_1981,N_1587);
nor U2009 (N_2009,N_1635,N_1533);
and U2010 (N_2010,N_1859,N_1680);
or U2011 (N_2011,N_1638,N_1887);
or U2012 (N_2012,N_1623,N_1770);
or U2013 (N_2013,N_1944,N_1863);
nor U2014 (N_2014,N_1585,N_1963);
and U2015 (N_2015,N_1643,N_1554);
or U2016 (N_2016,N_1945,N_1608);
nor U2017 (N_2017,N_1516,N_1550);
or U2018 (N_2018,N_1584,N_1960);
or U2019 (N_2019,N_1649,N_1890);
nor U2020 (N_2020,N_1631,N_1777);
or U2021 (N_2021,N_1742,N_1618);
or U2022 (N_2022,N_1738,N_1757);
or U2023 (N_2023,N_1878,N_1778);
and U2024 (N_2024,N_1789,N_1595);
or U2025 (N_2025,N_1568,N_1682);
nand U2026 (N_2026,N_1946,N_1606);
nand U2027 (N_2027,N_1813,N_1604);
and U2028 (N_2028,N_1528,N_1575);
or U2029 (N_2029,N_1684,N_1801);
nor U2030 (N_2030,N_1629,N_1959);
or U2031 (N_2031,N_1936,N_1990);
nor U2032 (N_2032,N_1931,N_1833);
xnor U2033 (N_2033,N_1821,N_1949);
or U2034 (N_2034,N_1676,N_1545);
and U2035 (N_2035,N_1612,N_1995);
or U2036 (N_2036,N_1647,N_1527);
nand U2037 (N_2037,N_1637,N_1529);
nor U2038 (N_2038,N_1885,N_1988);
or U2039 (N_2039,N_1715,N_1985);
or U2040 (N_2040,N_1734,N_1835);
nor U2041 (N_2041,N_1817,N_1669);
nand U2042 (N_2042,N_1819,N_1883);
nor U2043 (N_2043,N_1849,N_1611);
or U2044 (N_2044,N_1766,N_1888);
xnor U2045 (N_2045,N_1706,N_1621);
or U2046 (N_2046,N_1544,N_1593);
xnor U2047 (N_2047,N_1799,N_1722);
and U2048 (N_2048,N_1865,N_1563);
and U2049 (N_2049,N_1502,N_1724);
or U2050 (N_2050,N_1923,N_1930);
nor U2051 (N_2051,N_1681,N_1615);
xor U2052 (N_2052,N_1814,N_1573);
nand U2053 (N_2053,N_1927,N_1614);
or U2054 (N_2054,N_1654,N_1696);
nand U2055 (N_2055,N_1852,N_1751);
nand U2056 (N_2056,N_1505,N_1795);
nand U2057 (N_2057,N_1965,N_1639);
nand U2058 (N_2058,N_1521,N_1752);
nand U2059 (N_2059,N_1762,N_1882);
nor U2060 (N_2060,N_1871,N_1656);
and U2061 (N_2061,N_1727,N_1735);
nand U2062 (N_2062,N_1524,N_1553);
or U2063 (N_2063,N_1761,N_1576);
nand U2064 (N_2064,N_1806,N_1747);
nand U2065 (N_2065,N_1954,N_1517);
xor U2066 (N_2066,N_1627,N_1520);
and U2067 (N_2067,N_1601,N_1840);
or U2068 (N_2068,N_1815,N_1624);
and U2069 (N_2069,N_1699,N_1860);
xnor U2070 (N_2070,N_1707,N_1847);
xnor U2071 (N_2071,N_1597,N_1805);
nor U2072 (N_2072,N_1774,N_1879);
nand U2073 (N_2073,N_1744,N_1515);
nor U2074 (N_2074,N_1736,N_1519);
nand U2075 (N_2075,N_1672,N_1894);
nand U2076 (N_2076,N_1993,N_1832);
xor U2077 (N_2077,N_1809,N_1725);
nor U2078 (N_2078,N_1901,N_1561);
and U2079 (N_2079,N_1678,N_1934);
xnor U2080 (N_2080,N_1782,N_1763);
nand U2081 (N_2081,N_1663,N_1535);
and U2082 (N_2082,N_1961,N_1975);
or U2083 (N_2083,N_1896,N_1969);
nor U2084 (N_2084,N_1746,N_1594);
xor U2085 (N_2085,N_1552,N_1537);
nand U2086 (N_2086,N_1987,N_1820);
or U2087 (N_2087,N_1636,N_1500);
nor U2088 (N_2088,N_1864,N_1912);
nand U2089 (N_2089,N_1977,N_1773);
or U2090 (N_2090,N_1844,N_1791);
nand U2091 (N_2091,N_1753,N_1562);
nor U2092 (N_2092,N_1645,N_1915);
or U2093 (N_2093,N_1939,N_1571);
nand U2094 (N_2094,N_1677,N_1810);
nand U2095 (N_2095,N_1632,N_1857);
and U2096 (N_2096,N_1754,N_1708);
or U2097 (N_2097,N_1967,N_1530);
or U2098 (N_2098,N_1962,N_1523);
nor U2099 (N_2099,N_1951,N_1673);
nand U2100 (N_2100,N_1880,N_1551);
nand U2101 (N_2101,N_1732,N_1602);
and U2102 (N_2102,N_1626,N_1916);
nand U2103 (N_2103,N_1855,N_1698);
nor U2104 (N_2104,N_1633,N_1514);
nand U2105 (N_2105,N_1572,N_1589);
or U2106 (N_2106,N_1566,N_1688);
or U2107 (N_2107,N_1997,N_1943);
and U2108 (N_2108,N_1513,N_1846);
and U2109 (N_2109,N_1803,N_1641);
and U2110 (N_2110,N_1532,N_1812);
or U2111 (N_2111,N_1522,N_1827);
nand U2112 (N_2112,N_1902,N_1919);
nand U2113 (N_2113,N_1876,N_1854);
nor U2114 (N_2114,N_1994,N_1991);
and U2115 (N_2115,N_1549,N_1829);
or U2116 (N_2116,N_1978,N_1652);
or U2117 (N_2117,N_1657,N_1512);
and U2118 (N_2118,N_1560,N_1570);
or U2119 (N_2119,N_1913,N_1893);
nand U2120 (N_2120,N_1583,N_1619);
or U2121 (N_2121,N_1664,N_1726);
nor U2122 (N_2122,N_1870,N_1907);
nor U2123 (N_2123,N_1613,N_1824);
or U2124 (N_2124,N_1924,N_1947);
and U2125 (N_2125,N_1784,N_1596);
or U2126 (N_2126,N_1701,N_1556);
nor U2127 (N_2127,N_1668,N_1733);
xor U2128 (N_2128,N_1675,N_1980);
or U2129 (N_2129,N_1651,N_1536);
nor U2130 (N_2130,N_1794,N_1942);
nor U2131 (N_2131,N_1869,N_1765);
and U2132 (N_2132,N_1759,N_1546);
nand U2133 (N_2133,N_1692,N_1578);
and U2134 (N_2134,N_1848,N_1653);
nand U2135 (N_2135,N_1973,N_1889);
nor U2136 (N_2136,N_1822,N_1843);
and U2137 (N_2137,N_1581,N_1525);
nor U2138 (N_2138,N_1720,N_1866);
and U2139 (N_2139,N_1900,N_1650);
and U2140 (N_2140,N_1694,N_1592);
or U2141 (N_2141,N_1755,N_1504);
nor U2142 (N_2142,N_1966,N_1695);
or U2143 (N_2143,N_1640,N_1825);
nor U2144 (N_2144,N_1507,N_1783);
xor U2145 (N_2145,N_1714,N_1712);
and U2146 (N_2146,N_1964,N_1999);
or U2147 (N_2147,N_1796,N_1998);
or U2148 (N_2148,N_1767,N_1772);
or U2149 (N_2149,N_1590,N_1538);
xor U2150 (N_2150,N_1986,N_1582);
or U2151 (N_2151,N_1926,N_1737);
nand U2152 (N_2152,N_1970,N_1972);
and U2153 (N_2153,N_1713,N_1548);
and U2154 (N_2154,N_1598,N_1605);
nor U2155 (N_2155,N_1823,N_1620);
nor U2156 (N_2156,N_1937,N_1600);
nor U2157 (N_2157,N_1790,N_1910);
nor U2158 (N_2158,N_1874,N_1933);
and U2159 (N_2159,N_1719,N_1567);
or U2160 (N_2160,N_1957,N_1758);
and U2161 (N_2161,N_1983,N_1904);
nand U2162 (N_2162,N_1802,N_1591);
nand U2163 (N_2163,N_1974,N_1704);
or U2164 (N_2164,N_1674,N_1666);
nand U2165 (N_2165,N_1661,N_1716);
or U2166 (N_2166,N_1940,N_1897);
and U2167 (N_2167,N_1749,N_1886);
nor U2168 (N_2168,N_1800,N_1580);
nand U2169 (N_2169,N_1569,N_1792);
or U2170 (N_2170,N_1780,N_1984);
or U2171 (N_2171,N_1830,N_1793);
nor U2172 (N_2172,N_1510,N_1728);
or U2173 (N_2173,N_1911,N_1764);
nor U2174 (N_2174,N_1992,N_1642);
nor U2175 (N_2175,N_1828,N_1917);
or U2176 (N_2176,N_1577,N_1950);
or U2177 (N_2177,N_1531,N_1771);
or U2178 (N_2178,N_1982,N_1839);
nor U2179 (N_2179,N_1630,N_1616);
and U2180 (N_2180,N_1856,N_1555);
xor U2181 (N_2181,N_1729,N_1644);
nor U2182 (N_2182,N_1685,N_1873);
xor U2183 (N_2183,N_1776,N_1625);
nor U2184 (N_2184,N_1971,N_1700);
nor U2185 (N_2185,N_1646,N_1804);
and U2186 (N_2186,N_1586,N_1807);
xnor U2187 (N_2187,N_1834,N_1686);
nand U2188 (N_2188,N_1503,N_1785);
and U2189 (N_2189,N_1671,N_1895);
xor U2190 (N_2190,N_1941,N_1739);
nor U2191 (N_2191,N_1884,N_1508);
or U2192 (N_2192,N_1850,N_1842);
nand U2193 (N_2193,N_1607,N_1687);
xnor U2194 (N_2194,N_1748,N_1952);
nor U2195 (N_2195,N_1659,N_1797);
nor U2196 (N_2196,N_1922,N_1603);
or U2197 (N_2197,N_1976,N_1689);
or U2198 (N_2198,N_1918,N_1559);
nand U2199 (N_2199,N_1588,N_1609);
xnor U2200 (N_2200,N_1914,N_1534);
nand U2201 (N_2201,N_1731,N_1690);
nor U2202 (N_2202,N_1541,N_1634);
xor U2203 (N_2203,N_1557,N_1948);
or U2204 (N_2204,N_1705,N_1665);
nor U2205 (N_2205,N_1768,N_1798);
and U2206 (N_2206,N_1877,N_1921);
nand U2207 (N_2207,N_1655,N_1506);
nand U2208 (N_2208,N_1906,N_1542);
or U2209 (N_2209,N_1853,N_1979);
or U2210 (N_2210,N_1565,N_1938);
or U2211 (N_2211,N_1622,N_1861);
and U2212 (N_2212,N_1892,N_1697);
or U2213 (N_2213,N_1925,N_1501);
nand U2214 (N_2214,N_1811,N_1509);
and U2215 (N_2215,N_1838,N_1920);
nand U2216 (N_2216,N_1658,N_1511);
or U2217 (N_2217,N_1891,N_1543);
and U2218 (N_2218,N_1932,N_1745);
or U2219 (N_2219,N_1610,N_1908);
or U2220 (N_2220,N_1781,N_1717);
xnor U2221 (N_2221,N_1667,N_1691);
or U2222 (N_2222,N_1711,N_1905);
nor U2223 (N_2223,N_1760,N_1858);
nor U2224 (N_2224,N_1709,N_1928);
or U2225 (N_2225,N_1518,N_1837);
and U2226 (N_2226,N_1628,N_1741);
and U2227 (N_2227,N_1662,N_1836);
nor U2228 (N_2228,N_1955,N_1703);
nand U2229 (N_2229,N_1851,N_1898);
and U2230 (N_2230,N_1903,N_1935);
nand U2231 (N_2231,N_1743,N_1730);
and U2232 (N_2232,N_1750,N_1574);
nor U2233 (N_2233,N_1816,N_1558);
and U2234 (N_2234,N_1723,N_1958);
and U2235 (N_2235,N_1526,N_1710);
or U2236 (N_2236,N_1540,N_1953);
and U2237 (N_2237,N_1564,N_1867);
or U2238 (N_2238,N_1779,N_1881);
and U2239 (N_2239,N_1956,N_1808);
and U2240 (N_2240,N_1831,N_1599);
or U2241 (N_2241,N_1875,N_1769);
and U2242 (N_2242,N_1579,N_1989);
and U2243 (N_2243,N_1968,N_1788);
nand U2244 (N_2244,N_1648,N_1547);
nor U2245 (N_2245,N_1826,N_1868);
nor U2246 (N_2246,N_1818,N_1756);
and U2247 (N_2247,N_1899,N_1693);
xnor U2248 (N_2248,N_1862,N_1786);
nor U2249 (N_2249,N_1617,N_1787);
nand U2250 (N_2250,N_1901,N_1855);
nor U2251 (N_2251,N_1931,N_1939);
or U2252 (N_2252,N_1623,N_1941);
nor U2253 (N_2253,N_1731,N_1584);
nand U2254 (N_2254,N_1965,N_1885);
nand U2255 (N_2255,N_1981,N_1858);
xor U2256 (N_2256,N_1788,N_1564);
nand U2257 (N_2257,N_1644,N_1537);
and U2258 (N_2258,N_1734,N_1733);
or U2259 (N_2259,N_1907,N_1528);
and U2260 (N_2260,N_1686,N_1696);
and U2261 (N_2261,N_1687,N_1615);
and U2262 (N_2262,N_1530,N_1560);
or U2263 (N_2263,N_1939,N_1786);
nor U2264 (N_2264,N_1784,N_1698);
nor U2265 (N_2265,N_1923,N_1835);
and U2266 (N_2266,N_1957,N_1782);
xnor U2267 (N_2267,N_1943,N_1971);
nor U2268 (N_2268,N_1997,N_1635);
and U2269 (N_2269,N_1580,N_1635);
nor U2270 (N_2270,N_1861,N_1540);
and U2271 (N_2271,N_1697,N_1765);
and U2272 (N_2272,N_1615,N_1931);
and U2273 (N_2273,N_1775,N_1963);
nor U2274 (N_2274,N_1964,N_1913);
and U2275 (N_2275,N_1934,N_1946);
and U2276 (N_2276,N_1842,N_1858);
nor U2277 (N_2277,N_1745,N_1568);
or U2278 (N_2278,N_1993,N_1901);
nand U2279 (N_2279,N_1905,N_1640);
nand U2280 (N_2280,N_1611,N_1713);
xor U2281 (N_2281,N_1783,N_1768);
nand U2282 (N_2282,N_1506,N_1919);
nor U2283 (N_2283,N_1676,N_1839);
nor U2284 (N_2284,N_1558,N_1523);
xor U2285 (N_2285,N_1842,N_1753);
nand U2286 (N_2286,N_1510,N_1688);
nand U2287 (N_2287,N_1813,N_1985);
xor U2288 (N_2288,N_1807,N_1821);
nor U2289 (N_2289,N_1891,N_1792);
xnor U2290 (N_2290,N_1544,N_1877);
and U2291 (N_2291,N_1710,N_1662);
and U2292 (N_2292,N_1957,N_1872);
and U2293 (N_2293,N_1784,N_1766);
or U2294 (N_2294,N_1979,N_1859);
nor U2295 (N_2295,N_1528,N_1884);
and U2296 (N_2296,N_1579,N_1991);
and U2297 (N_2297,N_1755,N_1940);
nor U2298 (N_2298,N_1620,N_1655);
nand U2299 (N_2299,N_1848,N_1892);
and U2300 (N_2300,N_1770,N_1580);
nand U2301 (N_2301,N_1747,N_1945);
nor U2302 (N_2302,N_1743,N_1772);
nand U2303 (N_2303,N_1993,N_1610);
and U2304 (N_2304,N_1880,N_1706);
or U2305 (N_2305,N_1675,N_1590);
and U2306 (N_2306,N_1882,N_1509);
nand U2307 (N_2307,N_1823,N_1807);
nor U2308 (N_2308,N_1752,N_1986);
or U2309 (N_2309,N_1597,N_1601);
nand U2310 (N_2310,N_1733,N_1583);
and U2311 (N_2311,N_1632,N_1825);
xor U2312 (N_2312,N_1572,N_1788);
or U2313 (N_2313,N_1500,N_1705);
nor U2314 (N_2314,N_1753,N_1657);
nand U2315 (N_2315,N_1989,N_1688);
nand U2316 (N_2316,N_1934,N_1906);
and U2317 (N_2317,N_1901,N_1958);
and U2318 (N_2318,N_1775,N_1876);
nand U2319 (N_2319,N_1567,N_1547);
nor U2320 (N_2320,N_1795,N_1927);
and U2321 (N_2321,N_1911,N_1591);
nor U2322 (N_2322,N_1692,N_1876);
and U2323 (N_2323,N_1948,N_1660);
or U2324 (N_2324,N_1501,N_1560);
xnor U2325 (N_2325,N_1703,N_1901);
nor U2326 (N_2326,N_1942,N_1980);
and U2327 (N_2327,N_1757,N_1692);
and U2328 (N_2328,N_1907,N_1578);
and U2329 (N_2329,N_1577,N_1968);
xnor U2330 (N_2330,N_1826,N_1656);
nor U2331 (N_2331,N_1914,N_1756);
or U2332 (N_2332,N_1808,N_1796);
nand U2333 (N_2333,N_1604,N_1964);
or U2334 (N_2334,N_1829,N_1580);
nor U2335 (N_2335,N_1696,N_1729);
nor U2336 (N_2336,N_1581,N_1882);
and U2337 (N_2337,N_1916,N_1790);
nor U2338 (N_2338,N_1844,N_1821);
or U2339 (N_2339,N_1705,N_1990);
or U2340 (N_2340,N_1512,N_1931);
nor U2341 (N_2341,N_1766,N_1728);
nand U2342 (N_2342,N_1815,N_1504);
nor U2343 (N_2343,N_1723,N_1959);
nor U2344 (N_2344,N_1585,N_1517);
and U2345 (N_2345,N_1568,N_1948);
nand U2346 (N_2346,N_1962,N_1820);
and U2347 (N_2347,N_1717,N_1673);
and U2348 (N_2348,N_1822,N_1851);
xor U2349 (N_2349,N_1692,N_1514);
nand U2350 (N_2350,N_1529,N_1537);
nor U2351 (N_2351,N_1548,N_1941);
nand U2352 (N_2352,N_1842,N_1794);
or U2353 (N_2353,N_1846,N_1993);
nor U2354 (N_2354,N_1791,N_1663);
and U2355 (N_2355,N_1962,N_1884);
xnor U2356 (N_2356,N_1811,N_1902);
or U2357 (N_2357,N_1647,N_1701);
xor U2358 (N_2358,N_1765,N_1684);
nor U2359 (N_2359,N_1571,N_1963);
nand U2360 (N_2360,N_1796,N_1644);
nand U2361 (N_2361,N_1571,N_1705);
xnor U2362 (N_2362,N_1763,N_1636);
and U2363 (N_2363,N_1580,N_1771);
or U2364 (N_2364,N_1897,N_1943);
nand U2365 (N_2365,N_1887,N_1649);
nor U2366 (N_2366,N_1726,N_1914);
nand U2367 (N_2367,N_1987,N_1676);
nor U2368 (N_2368,N_1900,N_1857);
nand U2369 (N_2369,N_1533,N_1841);
nor U2370 (N_2370,N_1905,N_1729);
and U2371 (N_2371,N_1619,N_1645);
xnor U2372 (N_2372,N_1972,N_1926);
and U2373 (N_2373,N_1633,N_1811);
nand U2374 (N_2374,N_1586,N_1768);
nor U2375 (N_2375,N_1678,N_1980);
nand U2376 (N_2376,N_1585,N_1769);
xor U2377 (N_2377,N_1780,N_1832);
nor U2378 (N_2378,N_1582,N_1560);
and U2379 (N_2379,N_1580,N_1563);
nand U2380 (N_2380,N_1544,N_1951);
nor U2381 (N_2381,N_1630,N_1557);
nor U2382 (N_2382,N_1910,N_1832);
nand U2383 (N_2383,N_1852,N_1899);
xnor U2384 (N_2384,N_1543,N_1720);
or U2385 (N_2385,N_1990,N_1589);
and U2386 (N_2386,N_1502,N_1973);
or U2387 (N_2387,N_1518,N_1791);
and U2388 (N_2388,N_1500,N_1987);
and U2389 (N_2389,N_1901,N_1728);
nand U2390 (N_2390,N_1625,N_1879);
or U2391 (N_2391,N_1645,N_1901);
or U2392 (N_2392,N_1647,N_1551);
nor U2393 (N_2393,N_1934,N_1623);
nand U2394 (N_2394,N_1518,N_1808);
or U2395 (N_2395,N_1710,N_1726);
and U2396 (N_2396,N_1582,N_1662);
or U2397 (N_2397,N_1519,N_1856);
nor U2398 (N_2398,N_1653,N_1872);
or U2399 (N_2399,N_1948,N_1874);
nand U2400 (N_2400,N_1659,N_1533);
or U2401 (N_2401,N_1675,N_1990);
or U2402 (N_2402,N_1525,N_1803);
xnor U2403 (N_2403,N_1969,N_1794);
or U2404 (N_2404,N_1674,N_1988);
nand U2405 (N_2405,N_1913,N_1864);
nand U2406 (N_2406,N_1703,N_1554);
nor U2407 (N_2407,N_1704,N_1714);
nor U2408 (N_2408,N_1906,N_1791);
and U2409 (N_2409,N_1577,N_1619);
nand U2410 (N_2410,N_1521,N_1881);
nand U2411 (N_2411,N_1912,N_1804);
or U2412 (N_2412,N_1555,N_1997);
nor U2413 (N_2413,N_1905,N_1947);
and U2414 (N_2414,N_1835,N_1919);
nand U2415 (N_2415,N_1872,N_1963);
nor U2416 (N_2416,N_1582,N_1503);
nor U2417 (N_2417,N_1962,N_1763);
nand U2418 (N_2418,N_1763,N_1684);
or U2419 (N_2419,N_1805,N_1804);
nand U2420 (N_2420,N_1886,N_1812);
and U2421 (N_2421,N_1777,N_1739);
nor U2422 (N_2422,N_1840,N_1814);
or U2423 (N_2423,N_1553,N_1988);
or U2424 (N_2424,N_1660,N_1708);
nor U2425 (N_2425,N_1987,N_1611);
xor U2426 (N_2426,N_1655,N_1878);
or U2427 (N_2427,N_1868,N_1904);
nand U2428 (N_2428,N_1636,N_1842);
nor U2429 (N_2429,N_1771,N_1821);
and U2430 (N_2430,N_1782,N_1680);
xnor U2431 (N_2431,N_1701,N_1552);
nor U2432 (N_2432,N_1779,N_1687);
nor U2433 (N_2433,N_1737,N_1902);
nor U2434 (N_2434,N_1642,N_1951);
nor U2435 (N_2435,N_1866,N_1943);
nor U2436 (N_2436,N_1839,N_1606);
xor U2437 (N_2437,N_1561,N_1828);
nand U2438 (N_2438,N_1741,N_1508);
nand U2439 (N_2439,N_1536,N_1692);
nor U2440 (N_2440,N_1731,N_1679);
or U2441 (N_2441,N_1650,N_1914);
nor U2442 (N_2442,N_1674,N_1813);
and U2443 (N_2443,N_1588,N_1883);
nor U2444 (N_2444,N_1941,N_1764);
nor U2445 (N_2445,N_1514,N_1705);
nor U2446 (N_2446,N_1742,N_1709);
nand U2447 (N_2447,N_1902,N_1762);
and U2448 (N_2448,N_1589,N_1660);
nand U2449 (N_2449,N_1872,N_1596);
or U2450 (N_2450,N_1756,N_1960);
or U2451 (N_2451,N_1923,N_1733);
nor U2452 (N_2452,N_1617,N_1518);
nand U2453 (N_2453,N_1795,N_1554);
nand U2454 (N_2454,N_1725,N_1797);
and U2455 (N_2455,N_1597,N_1899);
or U2456 (N_2456,N_1657,N_1785);
and U2457 (N_2457,N_1902,N_1780);
or U2458 (N_2458,N_1774,N_1793);
or U2459 (N_2459,N_1567,N_1634);
nor U2460 (N_2460,N_1941,N_1874);
nand U2461 (N_2461,N_1664,N_1865);
nor U2462 (N_2462,N_1699,N_1656);
xor U2463 (N_2463,N_1503,N_1772);
nor U2464 (N_2464,N_1922,N_1812);
nand U2465 (N_2465,N_1663,N_1576);
nand U2466 (N_2466,N_1870,N_1929);
nand U2467 (N_2467,N_1546,N_1508);
and U2468 (N_2468,N_1985,N_1645);
and U2469 (N_2469,N_1914,N_1665);
and U2470 (N_2470,N_1825,N_1822);
nand U2471 (N_2471,N_1784,N_1545);
xor U2472 (N_2472,N_1914,N_1520);
nor U2473 (N_2473,N_1917,N_1748);
or U2474 (N_2474,N_1799,N_1528);
and U2475 (N_2475,N_1822,N_1688);
xor U2476 (N_2476,N_1865,N_1652);
or U2477 (N_2477,N_1869,N_1615);
nor U2478 (N_2478,N_1670,N_1849);
nor U2479 (N_2479,N_1633,N_1595);
or U2480 (N_2480,N_1602,N_1505);
or U2481 (N_2481,N_1804,N_1503);
nand U2482 (N_2482,N_1974,N_1644);
nor U2483 (N_2483,N_1882,N_1655);
nor U2484 (N_2484,N_1585,N_1908);
nor U2485 (N_2485,N_1812,N_1821);
and U2486 (N_2486,N_1910,N_1808);
and U2487 (N_2487,N_1985,N_1839);
or U2488 (N_2488,N_1780,N_1724);
nor U2489 (N_2489,N_1823,N_1619);
nand U2490 (N_2490,N_1631,N_1563);
nand U2491 (N_2491,N_1906,N_1531);
and U2492 (N_2492,N_1927,N_1883);
and U2493 (N_2493,N_1792,N_1578);
and U2494 (N_2494,N_1509,N_1649);
and U2495 (N_2495,N_1605,N_1826);
or U2496 (N_2496,N_1632,N_1642);
or U2497 (N_2497,N_1676,N_1695);
nand U2498 (N_2498,N_1797,N_1812);
or U2499 (N_2499,N_1639,N_1605);
nor U2500 (N_2500,N_2049,N_2097);
nor U2501 (N_2501,N_2161,N_2480);
or U2502 (N_2502,N_2260,N_2268);
nand U2503 (N_2503,N_2026,N_2245);
nand U2504 (N_2504,N_2218,N_2335);
and U2505 (N_2505,N_2415,N_2076);
and U2506 (N_2506,N_2212,N_2347);
nand U2507 (N_2507,N_2020,N_2429);
and U2508 (N_2508,N_2146,N_2185);
or U2509 (N_2509,N_2267,N_2265);
and U2510 (N_2510,N_2457,N_2287);
nor U2511 (N_2511,N_2277,N_2246);
or U2512 (N_2512,N_2010,N_2223);
and U2513 (N_2513,N_2148,N_2001);
nor U2514 (N_2514,N_2015,N_2176);
nor U2515 (N_2515,N_2012,N_2380);
nand U2516 (N_2516,N_2052,N_2111);
or U2517 (N_2517,N_2116,N_2203);
or U2518 (N_2518,N_2235,N_2110);
nand U2519 (N_2519,N_2201,N_2058);
or U2520 (N_2520,N_2389,N_2056);
and U2521 (N_2521,N_2135,N_2204);
and U2522 (N_2522,N_2120,N_2248);
nor U2523 (N_2523,N_2200,N_2048);
nor U2524 (N_2524,N_2392,N_2397);
or U2525 (N_2525,N_2388,N_2441);
xor U2526 (N_2526,N_2222,N_2450);
and U2527 (N_2527,N_2198,N_2408);
nor U2528 (N_2528,N_2409,N_2172);
nor U2529 (N_2529,N_2124,N_2394);
nor U2530 (N_2530,N_2381,N_2371);
nand U2531 (N_2531,N_2065,N_2121);
or U2532 (N_2532,N_2239,N_2206);
and U2533 (N_2533,N_2227,N_2313);
nor U2534 (N_2534,N_2241,N_2259);
and U2535 (N_2535,N_2150,N_2028);
or U2536 (N_2536,N_2363,N_2437);
or U2537 (N_2537,N_2168,N_2063);
nor U2538 (N_2538,N_2112,N_2413);
nor U2539 (N_2539,N_2411,N_2035);
nand U2540 (N_2540,N_2162,N_2432);
nand U2541 (N_2541,N_2333,N_2468);
nor U2542 (N_2542,N_2396,N_2405);
nand U2543 (N_2543,N_2329,N_2027);
and U2544 (N_2544,N_2194,N_2034);
nand U2545 (N_2545,N_2467,N_2122);
nand U2546 (N_2546,N_2127,N_2359);
nor U2547 (N_2547,N_2322,N_2266);
nor U2548 (N_2548,N_2365,N_2079);
nand U2549 (N_2549,N_2482,N_2354);
and U2550 (N_2550,N_2387,N_2478);
nand U2551 (N_2551,N_2103,N_2017);
nor U2552 (N_2552,N_2244,N_2033);
xnor U2553 (N_2553,N_2059,N_2226);
nor U2554 (N_2554,N_2327,N_2296);
and U2555 (N_2555,N_2062,N_2158);
nor U2556 (N_2556,N_2102,N_2153);
and U2557 (N_2557,N_2473,N_2350);
and U2558 (N_2558,N_2231,N_2283);
nor U2559 (N_2559,N_2126,N_2487);
nor U2560 (N_2560,N_2300,N_2298);
nand U2561 (N_2561,N_2323,N_2434);
or U2562 (N_2562,N_2175,N_2188);
or U2563 (N_2563,N_2317,N_2439);
or U2564 (N_2564,N_2495,N_2321);
nor U2565 (N_2565,N_2195,N_2237);
and U2566 (N_2566,N_2293,N_2332);
or U2567 (N_2567,N_2316,N_2009);
nand U2568 (N_2568,N_2319,N_2104);
and U2569 (N_2569,N_2479,N_2067);
nor U2570 (N_2570,N_2025,N_2073);
nor U2571 (N_2571,N_2207,N_2367);
nor U2572 (N_2572,N_2082,N_2159);
nor U2573 (N_2573,N_2419,N_2310);
nand U2574 (N_2574,N_2324,N_2081);
nor U2575 (N_2575,N_2431,N_2352);
nor U2576 (N_2576,N_2485,N_2414);
xor U2577 (N_2577,N_2088,N_2136);
and U2578 (N_2578,N_2286,N_2374);
nor U2579 (N_2579,N_2236,N_2118);
nand U2580 (N_2580,N_2433,N_2357);
nand U2581 (N_2581,N_2156,N_2232);
and U2582 (N_2582,N_2358,N_2233);
xor U2583 (N_2583,N_2336,N_2132);
and U2584 (N_2584,N_2092,N_2289);
or U2585 (N_2585,N_2100,N_2416);
nor U2586 (N_2586,N_2379,N_2094);
nand U2587 (N_2587,N_2217,N_2364);
nand U2588 (N_2588,N_2045,N_2421);
xor U2589 (N_2589,N_2472,N_2040);
xor U2590 (N_2590,N_2253,N_2403);
or U2591 (N_2591,N_2117,N_2187);
or U2592 (N_2592,N_2166,N_2279);
xnor U2593 (N_2593,N_2464,N_2004);
nand U2594 (N_2594,N_2474,N_2284);
or U2595 (N_2595,N_2054,N_2318);
and U2596 (N_2596,N_2440,N_2167);
nor U2597 (N_2597,N_2261,N_2142);
or U2598 (N_2598,N_2098,N_2143);
xor U2599 (N_2599,N_2077,N_2060);
nor U2600 (N_2600,N_2275,N_2171);
xnor U2601 (N_2601,N_2247,N_2447);
nand U2602 (N_2602,N_2230,N_2448);
xor U2603 (N_2603,N_2134,N_2210);
and U2604 (N_2604,N_2280,N_2084);
and U2605 (N_2605,N_2486,N_2193);
and U2606 (N_2606,N_2404,N_2443);
nor U2607 (N_2607,N_2196,N_2091);
nor U2608 (N_2608,N_2254,N_2177);
nor U2609 (N_2609,N_2471,N_2070);
or U2610 (N_2610,N_2240,N_2263);
and U2611 (N_2611,N_2356,N_2046);
nor U2612 (N_2612,N_2139,N_2490);
nand U2613 (N_2613,N_2024,N_2303);
nand U2614 (N_2614,N_2488,N_2055);
xnor U2615 (N_2615,N_2219,N_2007);
nand U2616 (N_2616,N_2368,N_2325);
and U2617 (N_2617,N_2191,N_2406);
nand U2618 (N_2618,N_2288,N_2256);
and U2619 (N_2619,N_2360,N_2087);
nor U2620 (N_2620,N_2013,N_2257);
nor U2621 (N_2621,N_2243,N_2407);
or U2622 (N_2622,N_2211,N_2197);
nor U2623 (N_2623,N_2453,N_2083);
nand U2624 (N_2624,N_2494,N_2221);
or U2625 (N_2625,N_2086,N_2469);
nor U2626 (N_2626,N_2216,N_2057);
nand U2627 (N_2627,N_2101,N_2115);
nor U2628 (N_2628,N_2229,N_2271);
nor U2629 (N_2629,N_2458,N_2163);
nand U2630 (N_2630,N_2242,N_2498);
and U2631 (N_2631,N_2308,N_2465);
nand U2632 (N_2632,N_2497,N_2064);
nor U2633 (N_2633,N_2138,N_2238);
nor U2634 (N_2634,N_2032,N_2080);
and U2635 (N_2635,N_2209,N_2170);
or U2636 (N_2636,N_2165,N_2186);
nor U2637 (N_2637,N_2422,N_2023);
nand U2638 (N_2638,N_2290,N_2192);
nand U2639 (N_2639,N_2330,N_2320);
nor U2640 (N_2640,N_2306,N_2011);
nor U2641 (N_2641,N_2400,N_2131);
or U2642 (N_2642,N_2003,N_2160);
nand U2643 (N_2643,N_2130,N_2305);
nor U2644 (N_2644,N_2022,N_2438);
or U2645 (N_2645,N_2152,N_2355);
xor U2646 (N_2646,N_2331,N_2029);
and U2647 (N_2647,N_2157,N_2382);
and U2648 (N_2648,N_2208,N_2466);
nand U2649 (N_2649,N_2493,N_2147);
xnor U2650 (N_2650,N_2425,N_2449);
xnor U2651 (N_2651,N_2018,N_2372);
and U2652 (N_2652,N_2395,N_2270);
xor U2653 (N_2653,N_2484,N_2169);
nor U2654 (N_2654,N_2285,N_2294);
and U2655 (N_2655,N_2462,N_2264);
xor U2656 (N_2656,N_2144,N_2050);
or U2657 (N_2657,N_2089,N_2299);
nor U2658 (N_2658,N_2417,N_2315);
or U2659 (N_2659,N_2068,N_2251);
or U2660 (N_2660,N_2002,N_2334);
and U2661 (N_2661,N_2053,N_2295);
and U2662 (N_2662,N_2398,N_2383);
and U2663 (N_2663,N_2436,N_2499);
nor U2664 (N_2664,N_2214,N_2399);
and U2665 (N_2665,N_2426,N_2173);
and U2666 (N_2666,N_2014,N_2456);
xnor U2667 (N_2667,N_2442,N_2039);
or U2668 (N_2668,N_2341,N_2427);
and U2669 (N_2669,N_2297,N_2113);
nor U2670 (N_2670,N_2307,N_2178);
nor U2671 (N_2671,N_2129,N_2326);
xor U2672 (N_2672,N_2038,N_2078);
nand U2673 (N_2673,N_2312,N_2224);
nor U2674 (N_2674,N_2149,N_2281);
nor U2675 (N_2675,N_2346,N_2071);
nor U2676 (N_2676,N_2107,N_2489);
and U2677 (N_2677,N_2154,N_2114);
nand U2678 (N_2678,N_2047,N_2314);
nor U2679 (N_2679,N_2301,N_2491);
nor U2680 (N_2680,N_2074,N_2483);
xnor U2681 (N_2681,N_2075,N_2199);
and U2682 (N_2682,N_2095,N_2037);
or U2683 (N_2683,N_2043,N_2444);
or U2684 (N_2684,N_2339,N_2430);
or U2685 (N_2685,N_2373,N_2292);
xnor U2686 (N_2686,N_2151,N_2402);
nand U2687 (N_2687,N_2386,N_2362);
or U2688 (N_2688,N_2338,N_2460);
xnor U2689 (N_2689,N_2435,N_2291);
nor U2690 (N_2690,N_2361,N_2492);
or U2691 (N_2691,N_2202,N_2390);
nor U2692 (N_2692,N_2328,N_2349);
xor U2693 (N_2693,N_2481,N_2424);
and U2694 (N_2694,N_2269,N_2133);
xnor U2695 (N_2695,N_2030,N_2476);
xnor U2696 (N_2696,N_2213,N_2125);
and U2697 (N_2697,N_2477,N_2446);
or U2698 (N_2698,N_2451,N_2377);
nand U2699 (N_2699,N_2343,N_2423);
and U2700 (N_2700,N_2181,N_2273);
xor U2701 (N_2701,N_2258,N_2096);
nor U2702 (N_2702,N_2378,N_2475);
nor U2703 (N_2703,N_2182,N_2385);
or U2704 (N_2704,N_2109,N_2412);
nand U2705 (N_2705,N_2042,N_2340);
nor U2706 (N_2706,N_2145,N_2179);
or U2707 (N_2707,N_2000,N_2418);
xor U2708 (N_2708,N_2044,N_2282);
or U2709 (N_2709,N_2189,N_2249);
xnor U2710 (N_2710,N_2375,N_2366);
nor U2711 (N_2711,N_2190,N_2250);
nand U2712 (N_2712,N_2345,N_2225);
or U2713 (N_2713,N_2351,N_2090);
and U2714 (N_2714,N_2452,N_2410);
nor U2715 (N_2715,N_2384,N_2106);
nor U2716 (N_2716,N_2344,N_2041);
nand U2717 (N_2717,N_2105,N_2278);
or U2718 (N_2718,N_2069,N_2093);
and U2719 (N_2719,N_2184,N_2348);
nor U2720 (N_2720,N_2459,N_2234);
nor U2721 (N_2721,N_2302,N_2141);
xnor U2722 (N_2722,N_2274,N_2183);
and U2723 (N_2723,N_2123,N_2016);
and U2724 (N_2724,N_2006,N_2463);
or U2725 (N_2725,N_2470,N_2137);
nor U2726 (N_2726,N_2304,N_2376);
or U2727 (N_2727,N_2337,N_2128);
and U2728 (N_2728,N_2461,N_2085);
and U2729 (N_2729,N_2496,N_2072);
or U2730 (N_2730,N_2255,N_2005);
nand U2731 (N_2731,N_2445,N_2262);
and U2732 (N_2732,N_2369,N_2220);
nand U2733 (N_2733,N_2099,N_2205);
nand U2734 (N_2734,N_2276,N_2008);
xor U2735 (N_2735,N_2140,N_2066);
or U2736 (N_2736,N_2342,N_2108);
or U2737 (N_2737,N_2180,N_2119);
and U2738 (N_2738,N_2021,N_2019);
and U2739 (N_2739,N_2174,N_2391);
xnor U2740 (N_2740,N_2353,N_2454);
nand U2741 (N_2741,N_2311,N_2309);
xor U2742 (N_2742,N_2164,N_2252);
xnor U2743 (N_2743,N_2215,N_2051);
or U2744 (N_2744,N_2031,N_2061);
nor U2745 (N_2745,N_2228,N_2455);
or U2746 (N_2746,N_2370,N_2272);
xnor U2747 (N_2747,N_2036,N_2420);
and U2748 (N_2748,N_2393,N_2401);
nor U2749 (N_2749,N_2155,N_2428);
or U2750 (N_2750,N_2435,N_2237);
nor U2751 (N_2751,N_2029,N_2236);
or U2752 (N_2752,N_2430,N_2004);
nor U2753 (N_2753,N_2190,N_2216);
and U2754 (N_2754,N_2455,N_2049);
or U2755 (N_2755,N_2004,N_2015);
nand U2756 (N_2756,N_2230,N_2485);
xnor U2757 (N_2757,N_2072,N_2123);
nand U2758 (N_2758,N_2225,N_2309);
nor U2759 (N_2759,N_2092,N_2367);
xnor U2760 (N_2760,N_2294,N_2128);
nor U2761 (N_2761,N_2204,N_2029);
nor U2762 (N_2762,N_2499,N_2111);
and U2763 (N_2763,N_2024,N_2119);
nor U2764 (N_2764,N_2453,N_2305);
nand U2765 (N_2765,N_2265,N_2200);
nor U2766 (N_2766,N_2069,N_2123);
and U2767 (N_2767,N_2424,N_2165);
xnor U2768 (N_2768,N_2323,N_2431);
or U2769 (N_2769,N_2401,N_2451);
or U2770 (N_2770,N_2464,N_2309);
nand U2771 (N_2771,N_2097,N_2191);
and U2772 (N_2772,N_2087,N_2090);
xor U2773 (N_2773,N_2272,N_2337);
nor U2774 (N_2774,N_2252,N_2340);
and U2775 (N_2775,N_2075,N_2437);
nor U2776 (N_2776,N_2336,N_2244);
or U2777 (N_2777,N_2247,N_2118);
and U2778 (N_2778,N_2021,N_2368);
xor U2779 (N_2779,N_2495,N_2194);
nor U2780 (N_2780,N_2416,N_2231);
nand U2781 (N_2781,N_2364,N_2381);
nand U2782 (N_2782,N_2151,N_2428);
or U2783 (N_2783,N_2328,N_2300);
or U2784 (N_2784,N_2255,N_2365);
nor U2785 (N_2785,N_2420,N_2278);
nand U2786 (N_2786,N_2419,N_2262);
and U2787 (N_2787,N_2345,N_2060);
and U2788 (N_2788,N_2250,N_2387);
nand U2789 (N_2789,N_2033,N_2141);
or U2790 (N_2790,N_2025,N_2004);
nand U2791 (N_2791,N_2112,N_2251);
nor U2792 (N_2792,N_2325,N_2263);
and U2793 (N_2793,N_2388,N_2111);
and U2794 (N_2794,N_2181,N_2281);
nand U2795 (N_2795,N_2152,N_2264);
nand U2796 (N_2796,N_2056,N_2209);
nand U2797 (N_2797,N_2131,N_2339);
nor U2798 (N_2798,N_2063,N_2099);
or U2799 (N_2799,N_2350,N_2465);
and U2800 (N_2800,N_2325,N_2436);
or U2801 (N_2801,N_2088,N_2121);
nor U2802 (N_2802,N_2074,N_2283);
nand U2803 (N_2803,N_2016,N_2159);
and U2804 (N_2804,N_2167,N_2230);
nor U2805 (N_2805,N_2479,N_2415);
nor U2806 (N_2806,N_2326,N_2316);
and U2807 (N_2807,N_2344,N_2257);
or U2808 (N_2808,N_2120,N_2018);
nand U2809 (N_2809,N_2363,N_2378);
or U2810 (N_2810,N_2473,N_2278);
and U2811 (N_2811,N_2089,N_2324);
nor U2812 (N_2812,N_2484,N_2303);
nor U2813 (N_2813,N_2490,N_2063);
nor U2814 (N_2814,N_2152,N_2301);
nand U2815 (N_2815,N_2014,N_2239);
nand U2816 (N_2816,N_2028,N_2105);
or U2817 (N_2817,N_2006,N_2146);
and U2818 (N_2818,N_2345,N_2003);
nand U2819 (N_2819,N_2086,N_2139);
or U2820 (N_2820,N_2286,N_2236);
nand U2821 (N_2821,N_2381,N_2471);
nand U2822 (N_2822,N_2435,N_2337);
and U2823 (N_2823,N_2444,N_2290);
nor U2824 (N_2824,N_2427,N_2183);
or U2825 (N_2825,N_2145,N_2131);
xnor U2826 (N_2826,N_2340,N_2458);
and U2827 (N_2827,N_2452,N_2082);
nand U2828 (N_2828,N_2356,N_2017);
and U2829 (N_2829,N_2040,N_2378);
nor U2830 (N_2830,N_2390,N_2103);
nor U2831 (N_2831,N_2381,N_2133);
nor U2832 (N_2832,N_2066,N_2106);
and U2833 (N_2833,N_2355,N_2421);
or U2834 (N_2834,N_2189,N_2277);
and U2835 (N_2835,N_2275,N_2073);
nor U2836 (N_2836,N_2106,N_2348);
nand U2837 (N_2837,N_2301,N_2458);
nor U2838 (N_2838,N_2100,N_2437);
nand U2839 (N_2839,N_2496,N_2056);
and U2840 (N_2840,N_2026,N_2203);
nand U2841 (N_2841,N_2098,N_2364);
and U2842 (N_2842,N_2442,N_2393);
nor U2843 (N_2843,N_2019,N_2168);
and U2844 (N_2844,N_2280,N_2424);
nor U2845 (N_2845,N_2221,N_2087);
and U2846 (N_2846,N_2262,N_2455);
xnor U2847 (N_2847,N_2032,N_2053);
or U2848 (N_2848,N_2218,N_2125);
nor U2849 (N_2849,N_2357,N_2180);
xor U2850 (N_2850,N_2418,N_2372);
and U2851 (N_2851,N_2117,N_2047);
nor U2852 (N_2852,N_2153,N_2416);
nand U2853 (N_2853,N_2234,N_2274);
and U2854 (N_2854,N_2063,N_2339);
xor U2855 (N_2855,N_2255,N_2208);
or U2856 (N_2856,N_2194,N_2479);
nor U2857 (N_2857,N_2256,N_2078);
nor U2858 (N_2858,N_2115,N_2460);
nand U2859 (N_2859,N_2229,N_2103);
nor U2860 (N_2860,N_2477,N_2245);
xor U2861 (N_2861,N_2168,N_2485);
nand U2862 (N_2862,N_2130,N_2495);
or U2863 (N_2863,N_2334,N_2090);
and U2864 (N_2864,N_2267,N_2354);
xnor U2865 (N_2865,N_2209,N_2231);
or U2866 (N_2866,N_2181,N_2147);
or U2867 (N_2867,N_2040,N_2157);
xnor U2868 (N_2868,N_2482,N_2016);
nor U2869 (N_2869,N_2059,N_2330);
nor U2870 (N_2870,N_2187,N_2093);
or U2871 (N_2871,N_2338,N_2328);
or U2872 (N_2872,N_2190,N_2385);
or U2873 (N_2873,N_2053,N_2382);
or U2874 (N_2874,N_2128,N_2490);
or U2875 (N_2875,N_2268,N_2157);
or U2876 (N_2876,N_2486,N_2007);
nor U2877 (N_2877,N_2283,N_2430);
nor U2878 (N_2878,N_2252,N_2432);
and U2879 (N_2879,N_2021,N_2154);
nand U2880 (N_2880,N_2038,N_2226);
and U2881 (N_2881,N_2220,N_2165);
xor U2882 (N_2882,N_2481,N_2016);
or U2883 (N_2883,N_2005,N_2026);
nand U2884 (N_2884,N_2073,N_2432);
nand U2885 (N_2885,N_2353,N_2008);
nor U2886 (N_2886,N_2376,N_2065);
or U2887 (N_2887,N_2211,N_2390);
nand U2888 (N_2888,N_2454,N_2277);
xor U2889 (N_2889,N_2431,N_2415);
and U2890 (N_2890,N_2245,N_2436);
nand U2891 (N_2891,N_2152,N_2456);
or U2892 (N_2892,N_2120,N_2250);
nand U2893 (N_2893,N_2325,N_2014);
xor U2894 (N_2894,N_2041,N_2439);
or U2895 (N_2895,N_2236,N_2034);
nand U2896 (N_2896,N_2401,N_2486);
or U2897 (N_2897,N_2441,N_2242);
or U2898 (N_2898,N_2193,N_2466);
and U2899 (N_2899,N_2091,N_2345);
and U2900 (N_2900,N_2177,N_2145);
and U2901 (N_2901,N_2342,N_2083);
nor U2902 (N_2902,N_2229,N_2043);
or U2903 (N_2903,N_2004,N_2165);
or U2904 (N_2904,N_2017,N_2142);
nand U2905 (N_2905,N_2176,N_2113);
and U2906 (N_2906,N_2050,N_2279);
nand U2907 (N_2907,N_2458,N_2298);
nor U2908 (N_2908,N_2451,N_2095);
and U2909 (N_2909,N_2142,N_2426);
or U2910 (N_2910,N_2309,N_2028);
nor U2911 (N_2911,N_2041,N_2117);
or U2912 (N_2912,N_2171,N_2305);
or U2913 (N_2913,N_2488,N_2415);
and U2914 (N_2914,N_2210,N_2398);
and U2915 (N_2915,N_2148,N_2285);
and U2916 (N_2916,N_2274,N_2158);
or U2917 (N_2917,N_2334,N_2073);
and U2918 (N_2918,N_2137,N_2152);
nor U2919 (N_2919,N_2237,N_2203);
nor U2920 (N_2920,N_2193,N_2075);
or U2921 (N_2921,N_2083,N_2355);
nor U2922 (N_2922,N_2292,N_2283);
and U2923 (N_2923,N_2403,N_2483);
xor U2924 (N_2924,N_2078,N_2277);
nand U2925 (N_2925,N_2234,N_2179);
or U2926 (N_2926,N_2370,N_2201);
nand U2927 (N_2927,N_2097,N_2098);
nor U2928 (N_2928,N_2443,N_2328);
and U2929 (N_2929,N_2442,N_2394);
xnor U2930 (N_2930,N_2308,N_2399);
or U2931 (N_2931,N_2458,N_2030);
nor U2932 (N_2932,N_2294,N_2174);
xnor U2933 (N_2933,N_2339,N_2247);
nor U2934 (N_2934,N_2262,N_2054);
nand U2935 (N_2935,N_2037,N_2438);
nor U2936 (N_2936,N_2080,N_2394);
nor U2937 (N_2937,N_2048,N_2439);
or U2938 (N_2938,N_2112,N_2435);
xnor U2939 (N_2939,N_2258,N_2436);
nor U2940 (N_2940,N_2341,N_2005);
or U2941 (N_2941,N_2470,N_2189);
or U2942 (N_2942,N_2318,N_2341);
and U2943 (N_2943,N_2443,N_2419);
nand U2944 (N_2944,N_2234,N_2214);
or U2945 (N_2945,N_2372,N_2312);
and U2946 (N_2946,N_2477,N_2189);
nand U2947 (N_2947,N_2007,N_2199);
nand U2948 (N_2948,N_2397,N_2093);
nand U2949 (N_2949,N_2202,N_2349);
or U2950 (N_2950,N_2399,N_2133);
or U2951 (N_2951,N_2368,N_2278);
or U2952 (N_2952,N_2238,N_2197);
or U2953 (N_2953,N_2135,N_2385);
xnor U2954 (N_2954,N_2191,N_2232);
nand U2955 (N_2955,N_2365,N_2279);
and U2956 (N_2956,N_2219,N_2145);
or U2957 (N_2957,N_2378,N_2025);
nand U2958 (N_2958,N_2286,N_2301);
nand U2959 (N_2959,N_2353,N_2135);
nor U2960 (N_2960,N_2130,N_2203);
nand U2961 (N_2961,N_2484,N_2441);
nor U2962 (N_2962,N_2261,N_2141);
nand U2963 (N_2963,N_2069,N_2089);
or U2964 (N_2964,N_2298,N_2473);
nor U2965 (N_2965,N_2167,N_2275);
xor U2966 (N_2966,N_2108,N_2290);
or U2967 (N_2967,N_2175,N_2484);
xnor U2968 (N_2968,N_2038,N_2404);
or U2969 (N_2969,N_2381,N_2027);
nand U2970 (N_2970,N_2286,N_2335);
nor U2971 (N_2971,N_2351,N_2367);
nor U2972 (N_2972,N_2238,N_2097);
or U2973 (N_2973,N_2068,N_2062);
and U2974 (N_2974,N_2396,N_2134);
nand U2975 (N_2975,N_2302,N_2373);
or U2976 (N_2976,N_2017,N_2481);
and U2977 (N_2977,N_2393,N_2297);
or U2978 (N_2978,N_2424,N_2498);
and U2979 (N_2979,N_2435,N_2441);
nand U2980 (N_2980,N_2275,N_2358);
and U2981 (N_2981,N_2252,N_2457);
nand U2982 (N_2982,N_2265,N_2037);
xnor U2983 (N_2983,N_2047,N_2459);
nor U2984 (N_2984,N_2151,N_2000);
xor U2985 (N_2985,N_2031,N_2434);
nor U2986 (N_2986,N_2255,N_2242);
nand U2987 (N_2987,N_2191,N_2342);
or U2988 (N_2988,N_2407,N_2106);
nand U2989 (N_2989,N_2063,N_2297);
or U2990 (N_2990,N_2432,N_2462);
and U2991 (N_2991,N_2217,N_2035);
xnor U2992 (N_2992,N_2273,N_2347);
nor U2993 (N_2993,N_2267,N_2311);
nand U2994 (N_2994,N_2087,N_2017);
and U2995 (N_2995,N_2215,N_2328);
or U2996 (N_2996,N_2057,N_2294);
or U2997 (N_2997,N_2332,N_2071);
or U2998 (N_2998,N_2360,N_2002);
and U2999 (N_2999,N_2183,N_2472);
nor U3000 (N_3000,N_2924,N_2631);
nor U3001 (N_3001,N_2986,N_2560);
nor U3002 (N_3002,N_2863,N_2927);
nor U3003 (N_3003,N_2868,N_2992);
and U3004 (N_3004,N_2996,N_2871);
and U3005 (N_3005,N_2659,N_2858);
nor U3006 (N_3006,N_2831,N_2643);
nand U3007 (N_3007,N_2591,N_2714);
or U3008 (N_3008,N_2964,N_2800);
nor U3009 (N_3009,N_2755,N_2592);
and U3010 (N_3010,N_2567,N_2564);
nor U3011 (N_3011,N_2570,N_2849);
xnor U3012 (N_3012,N_2799,N_2937);
or U3013 (N_3013,N_2874,N_2953);
or U3014 (N_3014,N_2517,N_2847);
or U3015 (N_3015,N_2782,N_2982);
nand U3016 (N_3016,N_2722,N_2754);
or U3017 (N_3017,N_2861,N_2683);
and U3018 (N_3018,N_2784,N_2597);
xor U3019 (N_3019,N_2575,N_2817);
nand U3020 (N_3020,N_2940,N_2795);
nand U3021 (N_3021,N_2700,N_2828);
nor U3022 (N_3022,N_2882,N_2619);
nor U3023 (N_3023,N_2712,N_2845);
nor U3024 (N_3024,N_2599,N_2840);
nand U3025 (N_3025,N_2688,N_2635);
or U3026 (N_3026,N_2743,N_2623);
nor U3027 (N_3027,N_2834,N_2933);
nor U3028 (N_3028,N_2629,N_2837);
or U3029 (N_3029,N_2565,N_2549);
nand U3030 (N_3030,N_2644,N_2864);
xnor U3031 (N_3031,N_2734,N_2855);
nor U3032 (N_3032,N_2595,N_2798);
xor U3033 (N_3033,N_2520,N_2785);
nor U3034 (N_3034,N_2757,N_2732);
xor U3035 (N_3035,N_2775,N_2507);
xnor U3036 (N_3036,N_2691,N_2690);
or U3037 (N_3037,N_2725,N_2534);
and U3038 (N_3038,N_2990,N_2848);
nor U3039 (N_3039,N_2749,N_2913);
nor U3040 (N_3040,N_2969,N_2918);
nor U3041 (N_3041,N_2931,N_2669);
or U3042 (N_3042,N_2970,N_2747);
nand U3043 (N_3043,N_2791,N_2949);
or U3044 (N_3044,N_2998,N_2668);
nor U3045 (N_3045,N_2952,N_2707);
or U3046 (N_3046,N_2822,N_2892);
xor U3047 (N_3047,N_2981,N_2706);
or U3048 (N_3048,N_2765,N_2737);
nor U3049 (N_3049,N_2720,N_2829);
nor U3050 (N_3050,N_2899,N_2955);
and U3051 (N_3051,N_2950,N_2508);
nand U3052 (N_3052,N_2699,N_2993);
nor U3053 (N_3053,N_2762,N_2652);
and U3054 (N_3054,N_2751,N_2917);
xnor U3055 (N_3055,N_2852,N_2671);
nor U3056 (N_3056,N_2793,N_2675);
or U3057 (N_3057,N_2532,N_2593);
or U3058 (N_3058,N_2803,N_2711);
and U3059 (N_3059,N_2729,N_2813);
nor U3060 (N_3060,N_2571,N_2826);
and U3061 (N_3061,N_2881,N_2735);
nand U3062 (N_3062,N_2963,N_2548);
nor U3063 (N_3063,N_2617,N_2736);
or U3064 (N_3064,N_2836,N_2985);
xor U3065 (N_3065,N_2502,N_2738);
or U3066 (N_3066,N_2854,N_2649);
or U3067 (N_3067,N_2514,N_2640);
xor U3068 (N_3068,N_2694,N_2503);
and U3069 (N_3069,N_2621,N_2606);
nand U3070 (N_3070,N_2862,N_2541);
and U3071 (N_3071,N_2760,N_2756);
and U3072 (N_3072,N_2883,N_2584);
nor U3073 (N_3073,N_2806,N_2512);
or U3074 (N_3074,N_2914,N_2995);
nor U3075 (N_3075,N_2824,N_2594);
nand U3076 (N_3076,N_2865,N_2632);
nor U3077 (N_3077,N_2947,N_2956);
and U3078 (N_3078,N_2523,N_2815);
nor U3079 (N_3079,N_2904,N_2888);
and U3080 (N_3080,N_2513,N_2609);
nand U3081 (N_3081,N_2544,N_2999);
and U3082 (N_3082,N_2919,N_2814);
nor U3083 (N_3083,N_2946,N_2976);
nor U3084 (N_3084,N_2681,N_2766);
nand U3085 (N_3085,N_2807,N_2586);
and U3086 (N_3086,N_2610,N_2596);
nor U3087 (N_3087,N_2884,N_2797);
and U3088 (N_3088,N_2979,N_2971);
xor U3089 (N_3089,N_2835,N_2604);
or U3090 (N_3090,N_2866,N_2587);
and U3091 (N_3091,N_2536,N_2524);
or U3092 (N_3092,N_2941,N_2618);
and U3093 (N_3093,N_2843,N_2769);
nand U3094 (N_3094,N_2670,N_2639);
nand U3095 (N_3095,N_2516,N_2857);
or U3096 (N_3096,N_2509,N_2601);
or U3097 (N_3097,N_2590,N_2771);
nand U3098 (N_3098,N_2958,N_2713);
xnor U3099 (N_3099,N_2891,N_2853);
or U3100 (N_3100,N_2501,N_2566);
xnor U3101 (N_3101,N_2821,N_2576);
and U3102 (N_3102,N_2518,N_2526);
xor U3103 (N_3103,N_2636,N_2702);
or U3104 (N_3104,N_2577,N_2960);
nand U3105 (N_3105,N_2530,N_2646);
and U3106 (N_3106,N_2569,N_2539);
nor U3107 (N_3107,N_2902,N_2653);
and U3108 (N_3108,N_2588,N_2948);
nor U3109 (N_3109,N_2647,N_2521);
xor U3110 (N_3110,N_2870,N_2889);
nand U3111 (N_3111,N_2708,N_2838);
and U3112 (N_3112,N_2574,N_2934);
nor U3113 (N_3113,N_2938,N_2731);
nor U3114 (N_3114,N_2908,N_2578);
nor U3115 (N_3115,N_2607,N_2562);
and U3116 (N_3116,N_2790,N_2974);
or U3117 (N_3117,N_2816,N_2906);
nor U3118 (N_3118,N_2978,N_2930);
nand U3119 (N_3119,N_2951,N_2867);
xnor U3120 (N_3120,N_2750,N_2580);
and U3121 (N_3121,N_2844,N_2638);
nor U3122 (N_3122,N_2959,N_2920);
nand U3123 (N_3123,N_2878,N_2825);
xnor U3124 (N_3124,N_2615,N_2774);
and U3125 (N_3125,N_2641,N_2833);
or U3126 (N_3126,N_2894,N_2678);
and U3127 (N_3127,N_2819,N_2674);
or U3128 (N_3128,N_2943,N_2905);
nand U3129 (N_3129,N_2783,N_2695);
or U3130 (N_3130,N_2812,N_2598);
and U3131 (N_3131,N_2616,N_2546);
nor U3132 (N_3132,N_2611,N_2925);
nor U3133 (N_3133,N_2528,N_2811);
and U3134 (N_3134,N_2525,N_2645);
nand U3135 (N_3135,N_2954,N_2667);
or U3136 (N_3136,N_2942,N_2733);
or U3137 (N_3137,N_2746,N_2657);
nor U3138 (N_3138,N_2748,N_2991);
nand U3139 (N_3139,N_2911,N_2701);
nand U3140 (N_3140,N_2781,N_2557);
nor U3141 (N_3141,N_2563,N_2697);
and U3142 (N_3142,N_2936,N_2910);
and U3143 (N_3143,N_2945,N_2801);
nand U3144 (N_3144,N_2551,N_2926);
and U3145 (N_3145,N_2921,N_2531);
or U3146 (N_3146,N_2778,N_2656);
or U3147 (N_3147,N_2552,N_2901);
and U3148 (N_3148,N_2535,N_2922);
and U3149 (N_3149,N_2624,N_2692);
nand U3150 (N_3150,N_2585,N_2608);
nor U3151 (N_3151,N_2772,N_2665);
nor U3152 (N_3152,N_2794,N_2686);
or U3153 (N_3153,N_2787,N_2500);
and U3154 (N_3154,N_2770,N_2676);
or U3155 (N_3155,N_2637,N_2543);
xor U3156 (N_3156,N_2988,N_2704);
and U3157 (N_3157,N_2573,N_2932);
xor U3158 (N_3158,N_2776,N_2510);
and U3159 (N_3159,N_2915,N_2581);
and U3160 (N_3160,N_2511,N_2547);
or U3161 (N_3161,N_2709,N_2809);
and U3162 (N_3162,N_2873,N_2506);
or U3163 (N_3163,N_2839,N_2630);
nand U3164 (N_3164,N_2987,N_2550);
nor U3165 (N_3165,N_2758,N_2684);
nand U3166 (N_3166,N_2880,N_2879);
nor U3167 (N_3167,N_2877,N_2529);
nor U3168 (N_3168,N_2582,N_2627);
or U3169 (N_3169,N_2851,N_2568);
xor U3170 (N_3170,N_2540,N_2850);
xor U3171 (N_3171,N_2710,N_2846);
nand U3172 (N_3172,N_2673,N_2788);
nand U3173 (N_3173,N_2648,N_2742);
or U3174 (N_3174,N_2808,N_2832);
xnor U3175 (N_3175,N_2962,N_2980);
or U3176 (N_3176,N_2537,N_2689);
and U3177 (N_3177,N_2898,N_2728);
and U3178 (N_3178,N_2759,N_2792);
xnor U3179 (N_3179,N_2763,N_2997);
or U3180 (N_3180,N_2715,N_2723);
or U3181 (N_3181,N_2764,N_2504);
or U3182 (N_3182,N_2698,N_2538);
and U3183 (N_3183,N_2869,N_2786);
or U3184 (N_3184,N_2890,N_2994);
and U3185 (N_3185,N_2796,N_2605);
nor U3186 (N_3186,N_2967,N_2827);
xor U3187 (N_3187,N_2730,N_2555);
and U3188 (N_3188,N_2944,N_2741);
or U3189 (N_3189,N_2693,N_2628);
nor U3190 (N_3190,N_2612,N_2753);
nor U3191 (N_3191,N_2841,N_2687);
xor U3192 (N_3192,N_2556,N_2777);
and U3193 (N_3193,N_2727,N_2533);
or U3194 (N_3194,N_2522,N_2802);
nand U3195 (N_3195,N_2716,N_2744);
nor U3196 (N_3196,N_2972,N_2527);
or U3197 (N_3197,N_2554,N_2872);
or U3198 (N_3198,N_2779,N_2705);
or U3199 (N_3199,N_2572,N_2859);
and U3200 (N_3200,N_2626,N_2957);
nor U3201 (N_3201,N_2696,N_2660);
nand U3202 (N_3202,N_2515,N_2614);
nor U3203 (N_3203,N_2966,N_2887);
nand U3204 (N_3204,N_2860,N_2625);
nand U3205 (N_3205,N_2789,N_2968);
or U3206 (N_3206,N_2897,N_2875);
nor U3207 (N_3207,N_2703,N_2558);
nand U3208 (N_3208,N_2654,N_2842);
nor U3209 (N_3209,N_2651,N_2885);
nor U3210 (N_3210,N_2896,N_2780);
or U3211 (N_3211,N_2583,N_2685);
nand U3212 (N_3212,N_2804,N_2900);
xnor U3213 (N_3213,N_2767,N_2909);
nor U3214 (N_3214,N_2893,N_2745);
or U3215 (N_3215,N_2672,N_2600);
nand U3216 (N_3216,N_2740,N_2907);
nand U3217 (N_3217,N_2724,N_2719);
xor U3218 (N_3218,N_2983,N_2561);
and U3219 (N_3219,N_2726,N_2886);
and U3220 (N_3220,N_2939,N_2622);
xor U3221 (N_3221,N_2805,N_2856);
nand U3222 (N_3222,N_2661,N_2663);
nor U3223 (N_3223,N_2929,N_2613);
nor U3224 (N_3224,N_2935,N_2545);
and U3225 (N_3225,N_2620,N_2677);
nand U3226 (N_3226,N_2752,N_2634);
and U3227 (N_3227,N_2721,N_2823);
nor U3228 (N_3228,N_2895,N_2989);
or U3229 (N_3229,N_2559,N_2923);
and U3230 (N_3230,N_2820,N_2658);
nand U3231 (N_3231,N_2680,N_2984);
and U3232 (N_3232,N_2662,N_2768);
or U3233 (N_3233,N_2977,N_2542);
or U3234 (N_3234,N_2718,N_2519);
xor U3235 (N_3235,N_2761,N_2912);
nor U3236 (N_3236,N_2633,N_2664);
nand U3237 (N_3237,N_2603,N_2975);
and U3238 (N_3238,N_2679,N_2965);
and U3239 (N_3239,N_2655,N_2666);
xor U3240 (N_3240,N_2773,N_2602);
nor U3241 (N_3241,N_2876,N_2650);
nand U3242 (N_3242,N_2682,N_2642);
or U3243 (N_3243,N_2830,N_2553);
nand U3244 (N_3244,N_2589,N_2505);
and U3245 (N_3245,N_2579,N_2961);
or U3246 (N_3246,N_2903,N_2717);
nor U3247 (N_3247,N_2973,N_2916);
and U3248 (N_3248,N_2739,N_2818);
or U3249 (N_3249,N_2928,N_2810);
and U3250 (N_3250,N_2684,N_2805);
or U3251 (N_3251,N_2625,N_2988);
nor U3252 (N_3252,N_2556,N_2692);
nor U3253 (N_3253,N_2759,N_2890);
and U3254 (N_3254,N_2976,N_2660);
nand U3255 (N_3255,N_2781,N_2823);
and U3256 (N_3256,N_2564,N_2720);
or U3257 (N_3257,N_2645,N_2619);
nand U3258 (N_3258,N_2885,N_2501);
or U3259 (N_3259,N_2766,N_2938);
nor U3260 (N_3260,N_2929,N_2673);
or U3261 (N_3261,N_2890,N_2696);
xor U3262 (N_3262,N_2517,N_2562);
or U3263 (N_3263,N_2985,N_2695);
and U3264 (N_3264,N_2896,N_2961);
nand U3265 (N_3265,N_2963,N_2986);
or U3266 (N_3266,N_2918,N_2585);
nor U3267 (N_3267,N_2976,N_2556);
nor U3268 (N_3268,N_2634,N_2985);
or U3269 (N_3269,N_2677,N_2700);
nand U3270 (N_3270,N_2546,N_2720);
nand U3271 (N_3271,N_2799,N_2845);
or U3272 (N_3272,N_2642,N_2885);
and U3273 (N_3273,N_2974,N_2708);
and U3274 (N_3274,N_2825,N_2642);
or U3275 (N_3275,N_2978,N_2965);
nor U3276 (N_3276,N_2911,N_2674);
and U3277 (N_3277,N_2817,N_2522);
and U3278 (N_3278,N_2759,N_2633);
and U3279 (N_3279,N_2905,N_2984);
and U3280 (N_3280,N_2827,N_2583);
and U3281 (N_3281,N_2981,N_2678);
or U3282 (N_3282,N_2525,N_2855);
nor U3283 (N_3283,N_2875,N_2843);
nand U3284 (N_3284,N_2728,N_2963);
xnor U3285 (N_3285,N_2549,N_2614);
and U3286 (N_3286,N_2935,N_2916);
and U3287 (N_3287,N_2901,N_2542);
nand U3288 (N_3288,N_2850,N_2861);
nor U3289 (N_3289,N_2631,N_2775);
and U3290 (N_3290,N_2987,N_2714);
nor U3291 (N_3291,N_2889,N_2926);
nor U3292 (N_3292,N_2523,N_2579);
nand U3293 (N_3293,N_2665,N_2783);
nor U3294 (N_3294,N_2933,N_2533);
or U3295 (N_3295,N_2561,N_2544);
xnor U3296 (N_3296,N_2789,N_2965);
and U3297 (N_3297,N_2567,N_2948);
nand U3298 (N_3298,N_2870,N_2752);
xnor U3299 (N_3299,N_2531,N_2883);
or U3300 (N_3300,N_2924,N_2659);
and U3301 (N_3301,N_2921,N_2740);
xnor U3302 (N_3302,N_2993,N_2882);
and U3303 (N_3303,N_2671,N_2550);
nand U3304 (N_3304,N_2872,N_2926);
and U3305 (N_3305,N_2727,N_2887);
nor U3306 (N_3306,N_2804,N_2922);
nor U3307 (N_3307,N_2925,N_2929);
nand U3308 (N_3308,N_2835,N_2564);
nor U3309 (N_3309,N_2982,N_2594);
and U3310 (N_3310,N_2938,N_2550);
and U3311 (N_3311,N_2862,N_2537);
nor U3312 (N_3312,N_2936,N_2725);
nand U3313 (N_3313,N_2709,N_2685);
nand U3314 (N_3314,N_2632,N_2501);
or U3315 (N_3315,N_2665,N_2626);
nand U3316 (N_3316,N_2890,N_2865);
and U3317 (N_3317,N_2972,N_2561);
or U3318 (N_3318,N_2911,N_2537);
nand U3319 (N_3319,N_2992,N_2921);
nor U3320 (N_3320,N_2769,N_2973);
and U3321 (N_3321,N_2808,N_2630);
or U3322 (N_3322,N_2706,N_2700);
nand U3323 (N_3323,N_2791,N_2596);
nand U3324 (N_3324,N_2906,N_2558);
and U3325 (N_3325,N_2608,N_2501);
xnor U3326 (N_3326,N_2710,N_2832);
or U3327 (N_3327,N_2936,N_2524);
and U3328 (N_3328,N_2865,N_2554);
or U3329 (N_3329,N_2798,N_2530);
nor U3330 (N_3330,N_2858,N_2785);
and U3331 (N_3331,N_2537,N_2515);
or U3332 (N_3332,N_2789,N_2978);
nand U3333 (N_3333,N_2640,N_2879);
xor U3334 (N_3334,N_2991,N_2727);
nor U3335 (N_3335,N_2880,N_2504);
nor U3336 (N_3336,N_2684,N_2827);
or U3337 (N_3337,N_2962,N_2522);
xnor U3338 (N_3338,N_2567,N_2599);
nand U3339 (N_3339,N_2685,N_2599);
or U3340 (N_3340,N_2858,N_2733);
nand U3341 (N_3341,N_2750,N_2759);
nand U3342 (N_3342,N_2863,N_2643);
nand U3343 (N_3343,N_2739,N_2654);
nand U3344 (N_3344,N_2614,N_2870);
nand U3345 (N_3345,N_2797,N_2905);
nand U3346 (N_3346,N_2633,N_2978);
nand U3347 (N_3347,N_2679,N_2842);
or U3348 (N_3348,N_2964,N_2806);
or U3349 (N_3349,N_2806,N_2864);
and U3350 (N_3350,N_2795,N_2979);
and U3351 (N_3351,N_2981,N_2684);
and U3352 (N_3352,N_2827,N_2615);
or U3353 (N_3353,N_2872,N_2691);
and U3354 (N_3354,N_2547,N_2891);
or U3355 (N_3355,N_2583,N_2844);
nand U3356 (N_3356,N_2568,N_2698);
xnor U3357 (N_3357,N_2971,N_2564);
xor U3358 (N_3358,N_2884,N_2760);
or U3359 (N_3359,N_2806,N_2611);
or U3360 (N_3360,N_2903,N_2841);
and U3361 (N_3361,N_2906,N_2808);
nand U3362 (N_3362,N_2737,N_2628);
nand U3363 (N_3363,N_2958,N_2595);
or U3364 (N_3364,N_2887,N_2866);
or U3365 (N_3365,N_2804,N_2535);
nor U3366 (N_3366,N_2769,N_2939);
or U3367 (N_3367,N_2890,N_2574);
nand U3368 (N_3368,N_2781,N_2980);
nand U3369 (N_3369,N_2707,N_2564);
nor U3370 (N_3370,N_2989,N_2909);
nand U3371 (N_3371,N_2905,N_2786);
and U3372 (N_3372,N_2639,N_2745);
and U3373 (N_3373,N_2852,N_2865);
or U3374 (N_3374,N_2678,N_2758);
xor U3375 (N_3375,N_2826,N_2851);
and U3376 (N_3376,N_2962,N_2975);
nand U3377 (N_3377,N_2610,N_2674);
or U3378 (N_3378,N_2502,N_2943);
nor U3379 (N_3379,N_2947,N_2619);
or U3380 (N_3380,N_2576,N_2765);
and U3381 (N_3381,N_2679,N_2777);
nor U3382 (N_3382,N_2551,N_2740);
and U3383 (N_3383,N_2677,N_2509);
xnor U3384 (N_3384,N_2872,N_2737);
and U3385 (N_3385,N_2869,N_2659);
xor U3386 (N_3386,N_2738,N_2890);
and U3387 (N_3387,N_2873,N_2881);
nand U3388 (N_3388,N_2894,N_2995);
and U3389 (N_3389,N_2807,N_2759);
and U3390 (N_3390,N_2544,N_2939);
nand U3391 (N_3391,N_2507,N_2948);
nor U3392 (N_3392,N_2825,N_2509);
nand U3393 (N_3393,N_2551,N_2540);
and U3394 (N_3394,N_2615,N_2826);
nand U3395 (N_3395,N_2817,N_2753);
or U3396 (N_3396,N_2688,N_2928);
or U3397 (N_3397,N_2758,N_2754);
nor U3398 (N_3398,N_2946,N_2649);
xor U3399 (N_3399,N_2826,N_2724);
or U3400 (N_3400,N_2830,N_2930);
nor U3401 (N_3401,N_2981,N_2665);
nand U3402 (N_3402,N_2824,N_2703);
or U3403 (N_3403,N_2769,N_2906);
nand U3404 (N_3404,N_2831,N_2506);
and U3405 (N_3405,N_2769,N_2852);
or U3406 (N_3406,N_2965,N_2623);
or U3407 (N_3407,N_2680,N_2864);
xnor U3408 (N_3408,N_2720,N_2623);
nor U3409 (N_3409,N_2555,N_2675);
nor U3410 (N_3410,N_2764,N_2918);
and U3411 (N_3411,N_2981,N_2809);
nor U3412 (N_3412,N_2585,N_2582);
xnor U3413 (N_3413,N_2625,N_2685);
and U3414 (N_3414,N_2986,N_2960);
nor U3415 (N_3415,N_2656,N_2826);
nand U3416 (N_3416,N_2547,N_2756);
and U3417 (N_3417,N_2566,N_2710);
nor U3418 (N_3418,N_2958,N_2842);
and U3419 (N_3419,N_2841,N_2923);
and U3420 (N_3420,N_2602,N_2786);
nor U3421 (N_3421,N_2783,N_2645);
or U3422 (N_3422,N_2756,N_2717);
or U3423 (N_3423,N_2917,N_2950);
and U3424 (N_3424,N_2685,N_2843);
xor U3425 (N_3425,N_2798,N_2503);
nand U3426 (N_3426,N_2723,N_2535);
or U3427 (N_3427,N_2884,N_2945);
or U3428 (N_3428,N_2743,N_2828);
nand U3429 (N_3429,N_2882,N_2527);
nand U3430 (N_3430,N_2595,N_2688);
nor U3431 (N_3431,N_2777,N_2552);
nand U3432 (N_3432,N_2526,N_2701);
nor U3433 (N_3433,N_2726,N_2927);
nand U3434 (N_3434,N_2694,N_2838);
or U3435 (N_3435,N_2800,N_2799);
nor U3436 (N_3436,N_2968,N_2788);
nand U3437 (N_3437,N_2895,N_2534);
nand U3438 (N_3438,N_2901,N_2926);
nand U3439 (N_3439,N_2831,N_2952);
nand U3440 (N_3440,N_2627,N_2639);
nand U3441 (N_3441,N_2736,N_2752);
or U3442 (N_3442,N_2570,N_2607);
xnor U3443 (N_3443,N_2696,N_2558);
and U3444 (N_3444,N_2878,N_2889);
nand U3445 (N_3445,N_2626,N_2602);
nand U3446 (N_3446,N_2982,N_2990);
and U3447 (N_3447,N_2938,N_2553);
xor U3448 (N_3448,N_2921,N_2807);
and U3449 (N_3449,N_2516,N_2518);
and U3450 (N_3450,N_2562,N_2915);
nand U3451 (N_3451,N_2792,N_2621);
nor U3452 (N_3452,N_2927,N_2743);
nand U3453 (N_3453,N_2995,N_2904);
nand U3454 (N_3454,N_2873,N_2818);
xor U3455 (N_3455,N_2883,N_2782);
nand U3456 (N_3456,N_2779,N_2928);
and U3457 (N_3457,N_2546,N_2935);
nor U3458 (N_3458,N_2663,N_2630);
and U3459 (N_3459,N_2741,N_2742);
and U3460 (N_3460,N_2705,N_2877);
nand U3461 (N_3461,N_2889,N_2991);
or U3462 (N_3462,N_2984,N_2799);
and U3463 (N_3463,N_2883,N_2724);
and U3464 (N_3464,N_2636,N_2645);
and U3465 (N_3465,N_2798,N_2836);
and U3466 (N_3466,N_2996,N_2954);
or U3467 (N_3467,N_2985,N_2666);
and U3468 (N_3468,N_2952,N_2930);
and U3469 (N_3469,N_2931,N_2649);
nand U3470 (N_3470,N_2986,N_2590);
and U3471 (N_3471,N_2977,N_2720);
nor U3472 (N_3472,N_2596,N_2834);
nor U3473 (N_3473,N_2819,N_2614);
nor U3474 (N_3474,N_2768,N_2635);
nor U3475 (N_3475,N_2910,N_2643);
or U3476 (N_3476,N_2909,N_2596);
and U3477 (N_3477,N_2822,N_2772);
and U3478 (N_3478,N_2510,N_2819);
nor U3479 (N_3479,N_2569,N_2659);
or U3480 (N_3480,N_2671,N_2891);
nand U3481 (N_3481,N_2732,N_2832);
and U3482 (N_3482,N_2698,N_2861);
or U3483 (N_3483,N_2785,N_2868);
and U3484 (N_3484,N_2712,N_2903);
nand U3485 (N_3485,N_2697,N_2789);
nor U3486 (N_3486,N_2991,N_2804);
xnor U3487 (N_3487,N_2696,N_2742);
nand U3488 (N_3488,N_2945,N_2755);
nor U3489 (N_3489,N_2764,N_2631);
nor U3490 (N_3490,N_2723,N_2714);
xnor U3491 (N_3491,N_2758,N_2834);
nand U3492 (N_3492,N_2559,N_2994);
nand U3493 (N_3493,N_2977,N_2622);
nor U3494 (N_3494,N_2716,N_2821);
nand U3495 (N_3495,N_2558,N_2974);
and U3496 (N_3496,N_2538,N_2869);
and U3497 (N_3497,N_2691,N_2682);
nor U3498 (N_3498,N_2712,N_2774);
and U3499 (N_3499,N_2717,N_2844);
nand U3500 (N_3500,N_3126,N_3273);
or U3501 (N_3501,N_3478,N_3060);
nor U3502 (N_3502,N_3074,N_3247);
nand U3503 (N_3503,N_3193,N_3169);
nor U3504 (N_3504,N_3113,N_3076);
or U3505 (N_3505,N_3174,N_3218);
and U3506 (N_3506,N_3456,N_3410);
nor U3507 (N_3507,N_3110,N_3133);
nand U3508 (N_3508,N_3122,N_3042);
nor U3509 (N_3509,N_3233,N_3062);
xnor U3510 (N_3510,N_3470,N_3085);
and U3511 (N_3511,N_3008,N_3214);
nor U3512 (N_3512,N_3031,N_3321);
xor U3513 (N_3513,N_3150,N_3418);
or U3514 (N_3514,N_3316,N_3070);
nor U3515 (N_3515,N_3088,N_3323);
nor U3516 (N_3516,N_3364,N_3403);
xnor U3517 (N_3517,N_3494,N_3077);
and U3518 (N_3518,N_3231,N_3275);
or U3519 (N_3519,N_3068,N_3017);
and U3520 (N_3520,N_3467,N_3400);
or U3521 (N_3521,N_3069,N_3151);
or U3522 (N_3522,N_3407,N_3288);
nor U3523 (N_3523,N_3251,N_3455);
or U3524 (N_3524,N_3472,N_3199);
xnor U3525 (N_3525,N_3004,N_3480);
xnor U3526 (N_3526,N_3277,N_3311);
or U3527 (N_3527,N_3454,N_3206);
nand U3528 (N_3528,N_3477,N_3191);
nand U3529 (N_3529,N_3237,N_3284);
nand U3530 (N_3530,N_3458,N_3269);
and U3531 (N_3531,N_3462,N_3268);
nor U3532 (N_3532,N_3302,N_3476);
or U3533 (N_3533,N_3198,N_3419);
and U3534 (N_3534,N_3356,N_3106);
or U3535 (N_3535,N_3125,N_3361);
or U3536 (N_3536,N_3224,N_3390);
nand U3537 (N_3537,N_3005,N_3227);
nand U3538 (N_3538,N_3093,N_3280);
xnor U3539 (N_3539,N_3200,N_3286);
nor U3540 (N_3540,N_3424,N_3406);
nor U3541 (N_3541,N_3378,N_3210);
nor U3542 (N_3542,N_3143,N_3234);
and U3543 (N_3543,N_3100,N_3355);
or U3544 (N_3544,N_3483,N_3160);
nand U3545 (N_3545,N_3437,N_3397);
xor U3546 (N_3546,N_3291,N_3059);
nor U3547 (N_3547,N_3440,N_3439);
or U3548 (N_3548,N_3033,N_3243);
nand U3549 (N_3549,N_3246,N_3282);
and U3550 (N_3550,N_3228,N_3072);
nand U3551 (N_3551,N_3138,N_3236);
nor U3552 (N_3552,N_3463,N_3026);
xor U3553 (N_3553,N_3117,N_3381);
nand U3554 (N_3554,N_3194,N_3444);
nand U3555 (N_3555,N_3149,N_3022);
nor U3556 (N_3556,N_3248,N_3445);
and U3557 (N_3557,N_3441,N_3057);
nor U3558 (N_3558,N_3166,N_3132);
or U3559 (N_3559,N_3036,N_3298);
nand U3560 (N_3560,N_3428,N_3091);
nand U3561 (N_3561,N_3384,N_3181);
nand U3562 (N_3562,N_3431,N_3482);
nor U3563 (N_3563,N_3207,N_3119);
nor U3564 (N_3564,N_3252,N_3346);
or U3565 (N_3565,N_3278,N_3197);
xnor U3566 (N_3566,N_3216,N_3367);
xnor U3567 (N_3567,N_3202,N_3374);
and U3568 (N_3568,N_3262,N_3087);
nand U3569 (N_3569,N_3489,N_3348);
nand U3570 (N_3570,N_3089,N_3493);
nor U3571 (N_3571,N_3308,N_3343);
or U3572 (N_3572,N_3305,N_3399);
xor U3573 (N_3573,N_3357,N_3156);
nor U3574 (N_3574,N_3449,N_3046);
xnor U3575 (N_3575,N_3289,N_3183);
xor U3576 (N_3576,N_3129,N_3433);
or U3577 (N_3577,N_3095,N_3195);
nor U3578 (N_3578,N_3386,N_3436);
nand U3579 (N_3579,N_3238,N_3351);
nand U3580 (N_3580,N_3371,N_3179);
nor U3581 (N_3581,N_3474,N_3242);
nor U3582 (N_3582,N_3137,N_3067);
or U3583 (N_3583,N_3063,N_3209);
and U3584 (N_3584,N_3263,N_3304);
or U3585 (N_3585,N_3294,N_3053);
and U3586 (N_3586,N_3312,N_3287);
or U3587 (N_3587,N_3297,N_3498);
or U3588 (N_3588,N_3421,N_3171);
nand U3589 (N_3589,N_3336,N_3239);
or U3590 (N_3590,N_3415,N_3338);
nor U3591 (N_3591,N_3468,N_3016);
and U3592 (N_3592,N_3081,N_3058);
nand U3593 (N_3593,N_3352,N_3230);
and U3594 (N_3594,N_3244,N_3101);
nand U3595 (N_3595,N_3054,N_3044);
nand U3596 (N_3596,N_3362,N_3011);
and U3597 (N_3597,N_3334,N_3222);
nor U3598 (N_3598,N_3028,N_3250);
nand U3599 (N_3599,N_3486,N_3414);
nand U3600 (N_3600,N_3385,N_3299);
or U3601 (N_3601,N_3102,N_3446);
or U3602 (N_3602,N_3354,N_3184);
nor U3603 (N_3603,N_3413,N_3182);
and U3604 (N_3604,N_3041,N_3189);
nor U3605 (N_3605,N_3145,N_3108);
or U3606 (N_3606,N_3372,N_3148);
and U3607 (N_3607,N_3034,N_3188);
nand U3608 (N_3608,N_3285,N_3073);
and U3609 (N_3609,N_3349,N_3377);
nand U3610 (N_3610,N_3303,N_3065);
and U3611 (N_3611,N_3394,N_3328);
xor U3612 (N_3612,N_3092,N_3121);
nand U3613 (N_3613,N_3382,N_3075);
nor U3614 (N_3614,N_3159,N_3154);
nand U3615 (N_3615,N_3043,N_3098);
and U3616 (N_3616,N_3429,N_3452);
and U3617 (N_3617,N_3442,N_3203);
and U3618 (N_3618,N_3499,N_3339);
nand U3619 (N_3619,N_3090,N_3315);
nor U3620 (N_3620,N_3164,N_3208);
and U3621 (N_3621,N_3422,N_3116);
and U3622 (N_3622,N_3003,N_3453);
and U3623 (N_3623,N_3322,N_3114);
and U3624 (N_3624,N_3411,N_3080);
or U3625 (N_3625,N_3402,N_3219);
nand U3626 (N_3626,N_3274,N_3459);
nand U3627 (N_3627,N_3387,N_3232);
nand U3628 (N_3628,N_3363,N_3438);
xor U3629 (N_3629,N_3401,N_3379);
and U3630 (N_3630,N_3450,N_3301);
xor U3631 (N_3631,N_3443,N_3490);
and U3632 (N_3632,N_3001,N_3404);
and U3633 (N_3633,N_3391,N_3084);
nor U3634 (N_3634,N_3358,N_3192);
xor U3635 (N_3635,N_3380,N_3327);
or U3636 (N_3636,N_3215,N_3395);
nand U3637 (N_3637,N_3266,N_3186);
and U3638 (N_3638,N_3447,N_3255);
xnor U3639 (N_3639,N_3405,N_3196);
or U3640 (N_3640,N_3479,N_3000);
and U3641 (N_3641,N_3465,N_3225);
nand U3642 (N_3642,N_3448,N_3120);
nor U3643 (N_3643,N_3333,N_3161);
and U3644 (N_3644,N_3375,N_3204);
and U3645 (N_3645,N_3165,N_3457);
nor U3646 (N_3646,N_3048,N_3146);
nor U3647 (N_3647,N_3078,N_3071);
xnor U3648 (N_3648,N_3006,N_3344);
and U3649 (N_3649,N_3290,N_3226);
xnor U3650 (N_3650,N_3221,N_3259);
or U3651 (N_3651,N_3013,N_3141);
nand U3652 (N_3652,N_3130,N_3432);
nor U3653 (N_3653,N_3331,N_3267);
nor U3654 (N_3654,N_3347,N_3396);
and U3655 (N_3655,N_3272,N_3389);
and U3656 (N_3656,N_3373,N_3383);
and U3657 (N_3657,N_3324,N_3134);
xor U3658 (N_3658,N_3366,N_3365);
or U3659 (N_3659,N_3061,N_3417);
nor U3660 (N_3660,N_3370,N_3025);
or U3661 (N_3661,N_3427,N_3020);
nor U3662 (N_3662,N_3103,N_3021);
and U3663 (N_3663,N_3083,N_3487);
or U3664 (N_3664,N_3435,N_3099);
and U3665 (N_3665,N_3050,N_3279);
nor U3666 (N_3666,N_3313,N_3350);
nor U3667 (N_3667,N_3292,N_3056);
xor U3668 (N_3668,N_3425,N_3131);
or U3669 (N_3669,N_3066,N_3475);
and U3670 (N_3670,N_3035,N_3241);
or U3671 (N_3671,N_3111,N_3270);
nand U3672 (N_3672,N_3388,N_3485);
nor U3673 (N_3673,N_3256,N_3167);
and U3674 (N_3674,N_3423,N_3326);
and U3675 (N_3675,N_3306,N_3109);
and U3676 (N_3676,N_3158,N_3329);
nor U3677 (N_3677,N_3140,N_3157);
xnor U3678 (N_3678,N_3086,N_3127);
nand U3679 (N_3679,N_3162,N_3155);
and U3680 (N_3680,N_3019,N_3332);
and U3681 (N_3681,N_3105,N_3420);
nand U3682 (N_3682,N_3045,N_3029);
nor U3683 (N_3683,N_3112,N_3293);
and U3684 (N_3684,N_3201,N_3211);
nor U3685 (N_3685,N_3369,N_3359);
and U3686 (N_3686,N_3296,N_3094);
and U3687 (N_3687,N_3104,N_3205);
nor U3688 (N_3688,N_3257,N_3253);
nor U3689 (N_3689,N_3314,N_3051);
nor U3690 (N_3690,N_3492,N_3317);
nand U3691 (N_3691,N_3055,N_3318);
and U3692 (N_3692,N_3039,N_3064);
or U3693 (N_3693,N_3220,N_3409);
nand U3694 (N_3694,N_3172,N_3037);
or U3695 (N_3695,N_3097,N_3027);
or U3696 (N_3696,N_3229,N_3049);
nor U3697 (N_3697,N_3281,N_3330);
or U3698 (N_3698,N_3002,N_3147);
or U3699 (N_3699,N_3177,N_3176);
nor U3700 (N_3700,N_3320,N_3124);
and U3701 (N_3701,N_3018,N_3142);
or U3702 (N_3702,N_3135,N_3310);
nand U3703 (N_3703,N_3325,N_3340);
xnor U3704 (N_3704,N_3096,N_3376);
and U3705 (N_3705,N_3024,N_3217);
nor U3706 (N_3706,N_3335,N_3212);
or U3707 (N_3707,N_3471,N_3190);
and U3708 (N_3708,N_3249,N_3283);
and U3709 (N_3709,N_3300,N_3258);
or U3710 (N_3710,N_3170,N_3223);
and U3711 (N_3711,N_3213,N_3144);
nor U3712 (N_3712,N_3342,N_3264);
nor U3713 (N_3713,N_3271,N_3240);
nand U3714 (N_3714,N_3168,N_3416);
xnor U3715 (N_3715,N_3015,N_3052);
nand U3716 (N_3716,N_3488,N_3497);
and U3717 (N_3717,N_3023,N_3464);
and U3718 (N_3718,N_3412,N_3175);
nand U3719 (N_3719,N_3163,N_3481);
nor U3720 (N_3720,N_3007,N_3484);
xor U3721 (N_3721,N_3152,N_3040);
xor U3722 (N_3722,N_3235,N_3260);
nand U3723 (N_3723,N_3451,N_3368);
or U3724 (N_3724,N_3265,N_3254);
or U3725 (N_3725,N_3360,N_3461);
nor U3726 (N_3726,N_3153,N_3139);
nand U3727 (N_3727,N_3012,N_3010);
and U3728 (N_3728,N_3460,N_3473);
xor U3729 (N_3729,N_3178,N_3187);
nor U3730 (N_3730,N_3495,N_3185);
nand U3731 (N_3731,N_3469,N_3115);
or U3732 (N_3732,N_3082,N_3295);
nand U3733 (N_3733,N_3276,N_3496);
and U3734 (N_3734,N_3107,N_3123);
or U3735 (N_3735,N_3309,N_3079);
or U3736 (N_3736,N_3408,N_3128);
nor U3737 (N_3737,N_3430,N_3319);
and U3738 (N_3738,N_3392,N_3491);
nor U3739 (N_3739,N_3261,N_3136);
and U3740 (N_3740,N_3180,N_3118);
nor U3741 (N_3741,N_3426,N_3434);
nand U3742 (N_3742,N_3398,N_3032);
xnor U3743 (N_3743,N_3014,N_3341);
and U3744 (N_3744,N_3337,N_3466);
and U3745 (N_3745,N_3353,N_3345);
xor U3746 (N_3746,N_3173,N_3030);
xor U3747 (N_3747,N_3047,N_3009);
nor U3748 (N_3748,N_3307,N_3393);
nor U3749 (N_3749,N_3245,N_3038);
nand U3750 (N_3750,N_3173,N_3411);
or U3751 (N_3751,N_3272,N_3059);
nor U3752 (N_3752,N_3283,N_3487);
and U3753 (N_3753,N_3403,N_3197);
nand U3754 (N_3754,N_3396,N_3202);
xnor U3755 (N_3755,N_3305,N_3307);
xor U3756 (N_3756,N_3387,N_3484);
and U3757 (N_3757,N_3351,N_3384);
or U3758 (N_3758,N_3294,N_3341);
and U3759 (N_3759,N_3152,N_3089);
nor U3760 (N_3760,N_3044,N_3055);
or U3761 (N_3761,N_3474,N_3362);
xnor U3762 (N_3762,N_3059,N_3070);
nor U3763 (N_3763,N_3339,N_3363);
nor U3764 (N_3764,N_3362,N_3275);
nor U3765 (N_3765,N_3290,N_3153);
nand U3766 (N_3766,N_3382,N_3082);
or U3767 (N_3767,N_3296,N_3203);
or U3768 (N_3768,N_3031,N_3134);
xor U3769 (N_3769,N_3197,N_3453);
and U3770 (N_3770,N_3082,N_3008);
xnor U3771 (N_3771,N_3419,N_3183);
nand U3772 (N_3772,N_3099,N_3315);
nor U3773 (N_3773,N_3380,N_3289);
nand U3774 (N_3774,N_3122,N_3175);
and U3775 (N_3775,N_3121,N_3298);
nor U3776 (N_3776,N_3198,N_3487);
and U3777 (N_3777,N_3239,N_3303);
nand U3778 (N_3778,N_3315,N_3043);
nor U3779 (N_3779,N_3130,N_3400);
and U3780 (N_3780,N_3095,N_3015);
xnor U3781 (N_3781,N_3211,N_3406);
nor U3782 (N_3782,N_3316,N_3320);
nand U3783 (N_3783,N_3165,N_3300);
nand U3784 (N_3784,N_3258,N_3339);
nor U3785 (N_3785,N_3184,N_3198);
and U3786 (N_3786,N_3248,N_3165);
or U3787 (N_3787,N_3465,N_3170);
nand U3788 (N_3788,N_3203,N_3421);
xor U3789 (N_3789,N_3408,N_3135);
nor U3790 (N_3790,N_3488,N_3120);
or U3791 (N_3791,N_3391,N_3186);
nor U3792 (N_3792,N_3027,N_3452);
nand U3793 (N_3793,N_3278,N_3057);
nand U3794 (N_3794,N_3355,N_3071);
or U3795 (N_3795,N_3269,N_3080);
nor U3796 (N_3796,N_3260,N_3283);
xor U3797 (N_3797,N_3041,N_3057);
nor U3798 (N_3798,N_3059,N_3370);
or U3799 (N_3799,N_3471,N_3128);
nand U3800 (N_3800,N_3263,N_3258);
or U3801 (N_3801,N_3152,N_3488);
nor U3802 (N_3802,N_3167,N_3243);
or U3803 (N_3803,N_3261,N_3108);
nand U3804 (N_3804,N_3495,N_3186);
or U3805 (N_3805,N_3221,N_3212);
nand U3806 (N_3806,N_3247,N_3251);
or U3807 (N_3807,N_3425,N_3038);
nand U3808 (N_3808,N_3257,N_3368);
xor U3809 (N_3809,N_3119,N_3302);
nand U3810 (N_3810,N_3145,N_3339);
nand U3811 (N_3811,N_3293,N_3358);
nor U3812 (N_3812,N_3393,N_3183);
or U3813 (N_3813,N_3256,N_3329);
nor U3814 (N_3814,N_3314,N_3313);
and U3815 (N_3815,N_3282,N_3168);
nor U3816 (N_3816,N_3244,N_3152);
nand U3817 (N_3817,N_3088,N_3171);
or U3818 (N_3818,N_3180,N_3318);
xnor U3819 (N_3819,N_3344,N_3300);
or U3820 (N_3820,N_3018,N_3099);
or U3821 (N_3821,N_3357,N_3210);
nor U3822 (N_3822,N_3245,N_3098);
nor U3823 (N_3823,N_3172,N_3428);
or U3824 (N_3824,N_3080,N_3002);
and U3825 (N_3825,N_3354,N_3000);
and U3826 (N_3826,N_3001,N_3483);
nor U3827 (N_3827,N_3015,N_3049);
or U3828 (N_3828,N_3318,N_3128);
xnor U3829 (N_3829,N_3140,N_3435);
or U3830 (N_3830,N_3219,N_3008);
xnor U3831 (N_3831,N_3419,N_3308);
nor U3832 (N_3832,N_3262,N_3025);
or U3833 (N_3833,N_3445,N_3104);
nand U3834 (N_3834,N_3015,N_3230);
and U3835 (N_3835,N_3369,N_3158);
nor U3836 (N_3836,N_3261,N_3467);
nand U3837 (N_3837,N_3220,N_3018);
and U3838 (N_3838,N_3377,N_3433);
and U3839 (N_3839,N_3015,N_3268);
or U3840 (N_3840,N_3023,N_3201);
nand U3841 (N_3841,N_3365,N_3049);
nand U3842 (N_3842,N_3184,N_3154);
and U3843 (N_3843,N_3064,N_3167);
or U3844 (N_3844,N_3031,N_3027);
xor U3845 (N_3845,N_3451,N_3142);
nor U3846 (N_3846,N_3300,N_3332);
and U3847 (N_3847,N_3219,N_3133);
or U3848 (N_3848,N_3367,N_3229);
or U3849 (N_3849,N_3170,N_3257);
nand U3850 (N_3850,N_3493,N_3421);
or U3851 (N_3851,N_3319,N_3093);
nand U3852 (N_3852,N_3073,N_3344);
and U3853 (N_3853,N_3050,N_3094);
or U3854 (N_3854,N_3212,N_3387);
nand U3855 (N_3855,N_3391,N_3287);
nand U3856 (N_3856,N_3134,N_3188);
nand U3857 (N_3857,N_3165,N_3211);
and U3858 (N_3858,N_3129,N_3301);
or U3859 (N_3859,N_3471,N_3423);
nor U3860 (N_3860,N_3113,N_3069);
or U3861 (N_3861,N_3029,N_3247);
nand U3862 (N_3862,N_3324,N_3275);
and U3863 (N_3863,N_3253,N_3074);
nand U3864 (N_3864,N_3105,N_3200);
nor U3865 (N_3865,N_3322,N_3423);
and U3866 (N_3866,N_3016,N_3327);
or U3867 (N_3867,N_3209,N_3343);
and U3868 (N_3868,N_3468,N_3099);
nand U3869 (N_3869,N_3223,N_3320);
nand U3870 (N_3870,N_3218,N_3496);
or U3871 (N_3871,N_3180,N_3179);
nor U3872 (N_3872,N_3295,N_3193);
or U3873 (N_3873,N_3429,N_3309);
and U3874 (N_3874,N_3037,N_3109);
nand U3875 (N_3875,N_3366,N_3445);
xor U3876 (N_3876,N_3197,N_3206);
and U3877 (N_3877,N_3085,N_3453);
or U3878 (N_3878,N_3463,N_3102);
xnor U3879 (N_3879,N_3152,N_3202);
nor U3880 (N_3880,N_3450,N_3361);
or U3881 (N_3881,N_3217,N_3498);
nor U3882 (N_3882,N_3250,N_3123);
xor U3883 (N_3883,N_3058,N_3387);
or U3884 (N_3884,N_3020,N_3496);
nor U3885 (N_3885,N_3387,N_3228);
and U3886 (N_3886,N_3035,N_3068);
nand U3887 (N_3887,N_3285,N_3474);
or U3888 (N_3888,N_3177,N_3194);
or U3889 (N_3889,N_3260,N_3132);
and U3890 (N_3890,N_3473,N_3026);
xnor U3891 (N_3891,N_3468,N_3226);
nor U3892 (N_3892,N_3399,N_3019);
xnor U3893 (N_3893,N_3095,N_3484);
and U3894 (N_3894,N_3287,N_3434);
and U3895 (N_3895,N_3360,N_3265);
or U3896 (N_3896,N_3224,N_3059);
or U3897 (N_3897,N_3093,N_3155);
or U3898 (N_3898,N_3299,N_3113);
nand U3899 (N_3899,N_3004,N_3139);
nor U3900 (N_3900,N_3183,N_3318);
nor U3901 (N_3901,N_3306,N_3072);
xor U3902 (N_3902,N_3482,N_3043);
or U3903 (N_3903,N_3329,N_3262);
and U3904 (N_3904,N_3205,N_3256);
nand U3905 (N_3905,N_3436,N_3301);
or U3906 (N_3906,N_3400,N_3426);
or U3907 (N_3907,N_3349,N_3452);
or U3908 (N_3908,N_3329,N_3270);
and U3909 (N_3909,N_3026,N_3317);
and U3910 (N_3910,N_3152,N_3228);
and U3911 (N_3911,N_3429,N_3005);
or U3912 (N_3912,N_3291,N_3372);
nand U3913 (N_3913,N_3309,N_3021);
and U3914 (N_3914,N_3336,N_3135);
xnor U3915 (N_3915,N_3333,N_3406);
or U3916 (N_3916,N_3120,N_3357);
nand U3917 (N_3917,N_3239,N_3217);
xor U3918 (N_3918,N_3127,N_3082);
and U3919 (N_3919,N_3009,N_3182);
and U3920 (N_3920,N_3266,N_3393);
or U3921 (N_3921,N_3248,N_3346);
nand U3922 (N_3922,N_3290,N_3340);
nor U3923 (N_3923,N_3213,N_3418);
nor U3924 (N_3924,N_3403,N_3200);
nor U3925 (N_3925,N_3353,N_3107);
nand U3926 (N_3926,N_3479,N_3292);
or U3927 (N_3927,N_3113,N_3302);
nand U3928 (N_3928,N_3201,N_3392);
nor U3929 (N_3929,N_3175,N_3100);
and U3930 (N_3930,N_3241,N_3112);
nor U3931 (N_3931,N_3013,N_3237);
or U3932 (N_3932,N_3497,N_3395);
nor U3933 (N_3933,N_3407,N_3099);
nor U3934 (N_3934,N_3416,N_3102);
or U3935 (N_3935,N_3458,N_3307);
and U3936 (N_3936,N_3402,N_3253);
nand U3937 (N_3937,N_3300,N_3130);
nand U3938 (N_3938,N_3369,N_3473);
xnor U3939 (N_3939,N_3462,N_3348);
or U3940 (N_3940,N_3129,N_3288);
nor U3941 (N_3941,N_3401,N_3150);
nand U3942 (N_3942,N_3013,N_3008);
nor U3943 (N_3943,N_3493,N_3015);
nand U3944 (N_3944,N_3314,N_3383);
nor U3945 (N_3945,N_3313,N_3375);
nand U3946 (N_3946,N_3261,N_3139);
and U3947 (N_3947,N_3112,N_3376);
or U3948 (N_3948,N_3010,N_3350);
and U3949 (N_3949,N_3297,N_3306);
nand U3950 (N_3950,N_3484,N_3200);
nor U3951 (N_3951,N_3375,N_3259);
nand U3952 (N_3952,N_3296,N_3353);
or U3953 (N_3953,N_3062,N_3060);
and U3954 (N_3954,N_3487,N_3484);
nor U3955 (N_3955,N_3413,N_3269);
nor U3956 (N_3956,N_3302,N_3330);
or U3957 (N_3957,N_3326,N_3447);
nand U3958 (N_3958,N_3256,N_3274);
nor U3959 (N_3959,N_3412,N_3320);
or U3960 (N_3960,N_3338,N_3293);
and U3961 (N_3961,N_3296,N_3455);
nor U3962 (N_3962,N_3447,N_3118);
and U3963 (N_3963,N_3118,N_3377);
and U3964 (N_3964,N_3362,N_3071);
nand U3965 (N_3965,N_3174,N_3394);
or U3966 (N_3966,N_3370,N_3450);
nor U3967 (N_3967,N_3046,N_3169);
or U3968 (N_3968,N_3430,N_3333);
and U3969 (N_3969,N_3086,N_3324);
nand U3970 (N_3970,N_3029,N_3020);
and U3971 (N_3971,N_3130,N_3284);
xor U3972 (N_3972,N_3051,N_3384);
xor U3973 (N_3973,N_3038,N_3341);
and U3974 (N_3974,N_3129,N_3304);
and U3975 (N_3975,N_3096,N_3337);
nand U3976 (N_3976,N_3407,N_3429);
or U3977 (N_3977,N_3466,N_3105);
xor U3978 (N_3978,N_3082,N_3344);
or U3979 (N_3979,N_3320,N_3108);
nand U3980 (N_3980,N_3403,N_3464);
nor U3981 (N_3981,N_3411,N_3278);
nor U3982 (N_3982,N_3298,N_3261);
nand U3983 (N_3983,N_3460,N_3213);
and U3984 (N_3984,N_3103,N_3176);
xnor U3985 (N_3985,N_3277,N_3034);
and U3986 (N_3986,N_3216,N_3376);
or U3987 (N_3987,N_3256,N_3330);
or U3988 (N_3988,N_3311,N_3086);
nor U3989 (N_3989,N_3417,N_3120);
or U3990 (N_3990,N_3185,N_3042);
and U3991 (N_3991,N_3340,N_3017);
nor U3992 (N_3992,N_3364,N_3354);
or U3993 (N_3993,N_3019,N_3016);
nor U3994 (N_3994,N_3337,N_3042);
or U3995 (N_3995,N_3285,N_3245);
and U3996 (N_3996,N_3089,N_3415);
and U3997 (N_3997,N_3215,N_3225);
and U3998 (N_3998,N_3492,N_3025);
and U3999 (N_3999,N_3132,N_3334);
nor U4000 (N_4000,N_3605,N_3819);
and U4001 (N_4001,N_3574,N_3554);
and U4002 (N_4002,N_3657,N_3851);
nor U4003 (N_4003,N_3993,N_3744);
xnor U4004 (N_4004,N_3955,N_3615);
or U4005 (N_4005,N_3603,N_3628);
and U4006 (N_4006,N_3613,N_3806);
xor U4007 (N_4007,N_3917,N_3811);
nand U4008 (N_4008,N_3751,N_3903);
nor U4009 (N_4009,N_3589,N_3681);
nor U4010 (N_4010,N_3975,N_3698);
nor U4011 (N_4011,N_3757,N_3976);
nand U4012 (N_4012,N_3969,N_3720);
or U4013 (N_4013,N_3511,N_3943);
or U4014 (N_4014,N_3640,N_3668);
xnor U4015 (N_4015,N_3826,N_3904);
and U4016 (N_4016,N_3716,N_3769);
and U4017 (N_4017,N_3669,N_3807);
nand U4018 (N_4018,N_3924,N_3521);
nor U4019 (N_4019,N_3643,N_3518);
and U4020 (N_4020,N_3753,N_3779);
nor U4021 (N_4021,N_3813,N_3771);
or U4022 (N_4022,N_3638,N_3763);
or U4023 (N_4023,N_3952,N_3877);
xnor U4024 (N_4024,N_3514,N_3503);
and U4025 (N_4025,N_3703,N_3506);
xor U4026 (N_4026,N_3876,N_3990);
and U4027 (N_4027,N_3540,N_3662);
nand U4028 (N_4028,N_3982,N_3983);
nor U4029 (N_4029,N_3792,N_3937);
and U4030 (N_4030,N_3594,N_3883);
and U4031 (N_4031,N_3998,N_3617);
or U4032 (N_4032,N_3833,N_3900);
xnor U4033 (N_4033,N_3596,N_3897);
nor U4034 (N_4034,N_3823,N_3762);
and U4035 (N_4035,N_3938,N_3765);
nor U4036 (N_4036,N_3967,N_3507);
and U4037 (N_4037,N_3670,N_3735);
or U4038 (N_4038,N_3542,N_3558);
or U4039 (N_4039,N_3634,N_3761);
nor U4040 (N_4040,N_3557,N_3799);
nor U4041 (N_4041,N_3738,N_3693);
xor U4042 (N_4042,N_3646,N_3855);
nand U4043 (N_4043,N_3785,N_3631);
nor U4044 (N_4044,N_3567,N_3838);
nand U4045 (N_4045,N_3986,N_3997);
xor U4046 (N_4046,N_3817,N_3915);
and U4047 (N_4047,N_3679,N_3930);
and U4048 (N_4048,N_3582,N_3641);
nand U4049 (N_4049,N_3798,N_3944);
nor U4050 (N_4050,N_3568,N_3630);
and U4051 (N_4051,N_3537,N_3885);
or U4052 (N_4052,N_3707,N_3754);
or U4053 (N_4053,N_3774,N_3687);
nand U4054 (N_4054,N_3690,N_3795);
and U4055 (N_4055,N_3783,N_3869);
nand U4056 (N_4056,N_3673,N_3614);
or U4057 (N_4057,N_3834,N_3674);
xor U4058 (N_4058,N_3538,N_3936);
or U4059 (N_4059,N_3736,N_3505);
nand U4060 (N_4060,N_3931,N_3878);
xor U4061 (N_4061,N_3595,N_3652);
xnor U4062 (N_4062,N_3750,N_3721);
xor U4063 (N_4063,N_3742,N_3991);
and U4064 (N_4064,N_3797,N_3841);
or U4065 (N_4065,N_3886,N_3760);
xnor U4066 (N_4066,N_3665,N_3803);
nand U4067 (N_4067,N_3780,N_3921);
nor U4068 (N_4068,N_3913,N_3724);
or U4069 (N_4069,N_3644,N_3545);
and U4070 (N_4070,N_3701,N_3859);
nor U4071 (N_4071,N_3896,N_3602);
nand U4072 (N_4072,N_3768,N_3905);
xnor U4073 (N_4073,N_3525,N_3844);
or U4074 (N_4074,N_3666,N_3529);
nand U4075 (N_4075,N_3516,N_3572);
and U4076 (N_4076,N_3714,N_3965);
xnor U4077 (N_4077,N_3879,N_3848);
nor U4078 (N_4078,N_3894,N_3898);
xor U4079 (N_4079,N_3950,N_3627);
xor U4080 (N_4080,N_3852,N_3973);
or U4081 (N_4081,N_3988,N_3947);
nor U4082 (N_4082,N_3692,N_3995);
or U4083 (N_4083,N_3712,N_3732);
nand U4084 (N_4084,N_3580,N_3565);
and U4085 (N_4085,N_3677,N_3637);
and U4086 (N_4086,N_3932,N_3512);
and U4087 (N_4087,N_3777,N_3658);
nor U4088 (N_4088,N_3981,N_3923);
and U4089 (N_4089,N_3942,N_3685);
nor U4090 (N_4090,N_3561,N_3906);
and U4091 (N_4091,N_3645,N_3513);
and U4092 (N_4092,N_3633,N_3578);
nand U4093 (N_4093,N_3840,N_3862);
and U4094 (N_4094,N_3680,N_3810);
nor U4095 (N_4095,N_3928,N_3961);
nor U4096 (N_4096,N_3532,N_3541);
nand U4097 (N_4097,N_3660,N_3620);
nor U4098 (N_4098,N_3782,N_3586);
nor U4099 (N_4099,N_3600,N_3935);
nor U4100 (N_4100,N_3530,N_3908);
nor U4101 (N_4101,N_3970,N_3555);
nor U4102 (N_4102,N_3764,N_3825);
and U4103 (N_4103,N_3684,N_3508);
and U4104 (N_4104,N_3718,N_3544);
nand U4105 (N_4105,N_3836,N_3543);
and U4106 (N_4106,N_3676,N_3749);
or U4107 (N_4107,N_3739,N_3767);
or U4108 (N_4108,N_3536,N_3748);
and U4109 (N_4109,N_3966,N_3925);
and U4110 (N_4110,N_3816,N_3667);
and U4111 (N_4111,N_3994,N_3746);
and U4112 (N_4112,N_3912,N_3711);
nor U4113 (N_4113,N_3927,N_3974);
xor U4114 (N_4114,N_3837,N_3728);
nand U4115 (N_4115,N_3881,N_3654);
xnor U4116 (N_4116,N_3522,N_3773);
or U4117 (N_4117,N_3534,N_3726);
and U4118 (N_4118,N_3733,N_3548);
nor U4119 (N_4119,N_3968,N_3978);
and U4120 (N_4120,N_3550,N_3664);
and U4121 (N_4121,N_3625,N_3672);
xor U4122 (N_4122,N_3571,N_3829);
xnor U4123 (N_4123,N_3846,N_3624);
nor U4124 (N_4124,N_3590,N_3651);
or U4125 (N_4125,N_3868,N_3926);
or U4126 (N_4126,N_3717,N_3700);
nand U4127 (N_4127,N_3989,N_3863);
or U4128 (N_4128,N_3688,N_3980);
nor U4129 (N_4129,N_3790,N_3719);
or U4130 (N_4130,N_3704,N_3585);
or U4131 (N_4131,N_3650,N_3891);
or U4132 (N_4132,N_3918,N_3832);
nor U4133 (N_4133,N_3963,N_3691);
nand U4134 (N_4134,N_3709,N_3830);
or U4135 (N_4135,N_3815,N_3710);
or U4136 (N_4136,N_3867,N_3575);
and U4137 (N_4137,N_3682,N_3941);
and U4138 (N_4138,N_3895,N_3737);
or U4139 (N_4139,N_3787,N_3962);
nand U4140 (N_4140,N_3598,N_3839);
and U4141 (N_4141,N_3500,N_3706);
and U4142 (N_4142,N_3591,N_3889);
xor U4143 (N_4143,N_3907,N_3547);
and U4144 (N_4144,N_3527,N_3656);
nor U4145 (N_4145,N_3653,N_3812);
xnor U4146 (N_4146,N_3636,N_3888);
nand U4147 (N_4147,N_3985,N_3861);
nand U4148 (N_4148,N_3729,N_3875);
and U4149 (N_4149,N_3880,N_3804);
or U4150 (N_4150,N_3610,N_3946);
nor U4151 (N_4151,N_3914,N_3805);
nand U4152 (N_4152,N_3933,N_3910);
nand U4153 (N_4153,N_3694,N_3501);
and U4154 (N_4154,N_3697,N_3874);
or U4155 (N_4155,N_3515,N_3526);
nor U4156 (N_4156,N_3911,N_3954);
or U4157 (N_4157,N_3919,N_3902);
or U4158 (N_4158,N_3597,N_3621);
xor U4159 (N_4159,N_3577,N_3854);
and U4160 (N_4160,N_3663,N_3971);
and U4161 (N_4161,N_3999,N_3964);
nor U4162 (N_4162,N_3678,N_3916);
nor U4163 (N_4163,N_3563,N_3722);
or U4164 (N_4164,N_3675,N_3642);
or U4165 (N_4165,N_3609,N_3996);
or U4166 (N_4166,N_3865,N_3979);
nand U4167 (N_4167,N_3551,N_3871);
or U4168 (N_4168,N_3699,N_3901);
and U4169 (N_4169,N_3593,N_3956);
nor U4170 (N_4170,N_3929,N_3899);
or U4171 (N_4171,N_3622,N_3570);
nand U4172 (N_4172,N_3922,N_3528);
xor U4173 (N_4173,N_3655,N_3647);
nand U4174 (N_4174,N_3853,N_3531);
and U4175 (N_4175,N_3629,N_3611);
or U4176 (N_4176,N_3781,N_3553);
nand U4177 (N_4177,N_3759,N_3820);
xnor U4178 (N_4178,N_3958,N_3581);
or U4179 (N_4179,N_3870,N_3766);
xor U4180 (N_4180,N_3835,N_3616);
nor U4181 (N_4181,N_3856,N_3794);
and U4182 (N_4182,N_3713,N_3770);
nand U4183 (N_4183,N_3793,N_3520);
or U4184 (N_4184,N_3909,N_3705);
nor U4185 (N_4185,N_3802,N_3573);
nand U4186 (N_4186,N_3623,N_3951);
and U4187 (N_4187,N_3731,N_3509);
xnor U4188 (N_4188,N_3519,N_3892);
nor U4189 (N_4189,N_3984,N_3758);
nor U4190 (N_4190,N_3887,N_3523);
nand U4191 (N_4191,N_3756,N_3510);
xnor U4192 (N_4192,N_3725,N_3784);
and U4193 (N_4193,N_3884,N_3619);
nor U4194 (N_4194,N_3775,N_3648);
nor U4195 (N_4195,N_3827,N_3727);
nor U4196 (N_4196,N_3639,N_3800);
or U4197 (N_4197,N_3940,N_3517);
and U4198 (N_4198,N_3945,N_3612);
and U4199 (N_4199,N_3893,N_3960);
nand U4200 (N_4200,N_3873,N_3576);
nand U4201 (N_4201,N_3850,N_3743);
nor U4202 (N_4202,N_3702,N_3659);
or U4203 (N_4203,N_3649,N_3708);
nand U4204 (N_4204,N_3755,N_3776);
nor U4205 (N_4205,N_3814,N_3745);
or U4206 (N_4206,N_3723,N_3824);
nor U4207 (N_4207,N_3552,N_3864);
and U4208 (N_4208,N_3959,N_3579);
nand U4209 (N_4209,N_3972,N_3987);
and U4210 (N_4210,N_3564,N_3524);
or U4211 (N_4211,N_3788,N_3546);
xnor U4212 (N_4212,N_3872,N_3858);
nand U4213 (N_4213,N_3796,N_3566);
and U4214 (N_4214,N_3671,N_3977);
and U4215 (N_4215,N_3696,N_3601);
nand U4216 (N_4216,N_3502,N_3556);
nor U4217 (N_4217,N_3730,N_3953);
and U4218 (N_4218,N_3604,N_3828);
and U4219 (N_4219,N_3618,N_3778);
nand U4220 (N_4220,N_3635,N_3822);
nand U4221 (N_4221,N_3842,N_3808);
nand U4222 (N_4222,N_3632,N_3801);
nand U4223 (N_4223,N_3584,N_3741);
nand U4224 (N_4224,N_3686,N_3847);
nand U4225 (N_4225,N_3569,N_3821);
nand U4226 (N_4226,N_3583,N_3866);
or U4227 (N_4227,N_3626,N_3890);
or U4228 (N_4228,N_3606,N_3809);
nand U4229 (N_4229,N_3789,N_3939);
or U4230 (N_4230,N_3740,N_3957);
and U4231 (N_4231,N_3549,N_3772);
and U4232 (N_4232,N_3831,N_3845);
nor U4233 (N_4233,N_3592,N_3535);
or U4234 (N_4234,N_3949,N_3948);
nor U4235 (N_4235,N_3695,N_3588);
nor U4236 (N_4236,N_3533,N_3608);
nand U4237 (N_4237,N_3934,N_3607);
or U4238 (N_4238,N_3661,N_3752);
nand U4239 (N_4239,N_3857,N_3504);
and U4240 (N_4240,N_3599,N_3791);
or U4241 (N_4241,N_3882,N_3920);
nand U4242 (N_4242,N_3734,N_3715);
and U4243 (N_4243,N_3689,N_3849);
nand U4244 (N_4244,N_3587,N_3747);
nand U4245 (N_4245,N_3683,N_3860);
or U4246 (N_4246,N_3786,N_3818);
and U4247 (N_4247,N_3559,N_3843);
xor U4248 (N_4248,N_3992,N_3539);
and U4249 (N_4249,N_3562,N_3560);
nand U4250 (N_4250,N_3621,N_3799);
or U4251 (N_4251,N_3709,N_3726);
nor U4252 (N_4252,N_3954,N_3979);
nand U4253 (N_4253,N_3693,N_3575);
and U4254 (N_4254,N_3904,N_3856);
or U4255 (N_4255,N_3833,N_3774);
or U4256 (N_4256,N_3989,N_3630);
and U4257 (N_4257,N_3760,N_3820);
and U4258 (N_4258,N_3532,N_3638);
xor U4259 (N_4259,N_3884,N_3953);
and U4260 (N_4260,N_3875,N_3690);
nand U4261 (N_4261,N_3590,N_3664);
or U4262 (N_4262,N_3667,N_3910);
or U4263 (N_4263,N_3732,N_3682);
nor U4264 (N_4264,N_3601,N_3967);
or U4265 (N_4265,N_3695,N_3587);
or U4266 (N_4266,N_3973,N_3551);
or U4267 (N_4267,N_3653,N_3904);
nor U4268 (N_4268,N_3603,N_3945);
and U4269 (N_4269,N_3886,N_3516);
nor U4270 (N_4270,N_3500,N_3937);
nand U4271 (N_4271,N_3710,N_3894);
or U4272 (N_4272,N_3847,N_3749);
nand U4273 (N_4273,N_3940,N_3841);
and U4274 (N_4274,N_3780,N_3905);
and U4275 (N_4275,N_3852,N_3788);
or U4276 (N_4276,N_3847,N_3858);
nand U4277 (N_4277,N_3608,N_3817);
and U4278 (N_4278,N_3676,N_3549);
or U4279 (N_4279,N_3755,N_3688);
and U4280 (N_4280,N_3641,N_3851);
or U4281 (N_4281,N_3719,N_3632);
nor U4282 (N_4282,N_3778,N_3748);
nor U4283 (N_4283,N_3918,N_3649);
and U4284 (N_4284,N_3618,N_3842);
or U4285 (N_4285,N_3937,N_3896);
xnor U4286 (N_4286,N_3537,N_3792);
nor U4287 (N_4287,N_3701,N_3887);
or U4288 (N_4288,N_3680,N_3649);
nor U4289 (N_4289,N_3560,N_3809);
and U4290 (N_4290,N_3514,N_3637);
nor U4291 (N_4291,N_3812,N_3793);
or U4292 (N_4292,N_3639,N_3811);
nor U4293 (N_4293,N_3964,N_3735);
and U4294 (N_4294,N_3508,N_3570);
nor U4295 (N_4295,N_3730,N_3676);
and U4296 (N_4296,N_3931,N_3990);
nand U4297 (N_4297,N_3872,N_3697);
nand U4298 (N_4298,N_3749,N_3833);
nand U4299 (N_4299,N_3948,N_3524);
and U4300 (N_4300,N_3520,N_3897);
and U4301 (N_4301,N_3503,N_3682);
or U4302 (N_4302,N_3529,N_3537);
nor U4303 (N_4303,N_3890,N_3539);
xor U4304 (N_4304,N_3769,N_3880);
xnor U4305 (N_4305,N_3683,N_3760);
nor U4306 (N_4306,N_3899,N_3900);
or U4307 (N_4307,N_3989,N_3865);
and U4308 (N_4308,N_3996,N_3541);
or U4309 (N_4309,N_3503,N_3670);
and U4310 (N_4310,N_3744,N_3873);
or U4311 (N_4311,N_3681,N_3783);
nor U4312 (N_4312,N_3888,N_3987);
or U4313 (N_4313,N_3694,N_3610);
nand U4314 (N_4314,N_3805,N_3727);
and U4315 (N_4315,N_3710,N_3911);
and U4316 (N_4316,N_3507,N_3965);
xnor U4317 (N_4317,N_3590,N_3673);
or U4318 (N_4318,N_3791,N_3601);
nand U4319 (N_4319,N_3744,N_3601);
nor U4320 (N_4320,N_3997,N_3644);
nand U4321 (N_4321,N_3723,N_3942);
nor U4322 (N_4322,N_3792,N_3827);
xor U4323 (N_4323,N_3775,N_3855);
nor U4324 (N_4324,N_3874,N_3794);
and U4325 (N_4325,N_3811,N_3633);
xnor U4326 (N_4326,N_3904,N_3764);
or U4327 (N_4327,N_3508,N_3587);
nand U4328 (N_4328,N_3853,N_3727);
xor U4329 (N_4329,N_3522,N_3524);
and U4330 (N_4330,N_3917,N_3745);
and U4331 (N_4331,N_3814,N_3828);
or U4332 (N_4332,N_3520,N_3922);
nor U4333 (N_4333,N_3614,N_3516);
or U4334 (N_4334,N_3681,N_3525);
nand U4335 (N_4335,N_3692,N_3697);
nand U4336 (N_4336,N_3858,N_3808);
and U4337 (N_4337,N_3837,N_3527);
or U4338 (N_4338,N_3837,N_3982);
and U4339 (N_4339,N_3573,N_3851);
nand U4340 (N_4340,N_3837,N_3509);
nor U4341 (N_4341,N_3937,N_3599);
or U4342 (N_4342,N_3753,N_3867);
or U4343 (N_4343,N_3950,N_3624);
nand U4344 (N_4344,N_3650,N_3593);
and U4345 (N_4345,N_3938,N_3912);
or U4346 (N_4346,N_3677,N_3630);
and U4347 (N_4347,N_3689,N_3698);
nand U4348 (N_4348,N_3533,N_3841);
and U4349 (N_4349,N_3796,N_3679);
xnor U4350 (N_4350,N_3938,N_3852);
nor U4351 (N_4351,N_3618,N_3579);
and U4352 (N_4352,N_3719,N_3950);
nand U4353 (N_4353,N_3621,N_3508);
nor U4354 (N_4354,N_3547,N_3694);
nand U4355 (N_4355,N_3546,N_3946);
nand U4356 (N_4356,N_3848,N_3888);
and U4357 (N_4357,N_3817,N_3772);
or U4358 (N_4358,N_3811,N_3964);
nor U4359 (N_4359,N_3998,N_3542);
or U4360 (N_4360,N_3748,N_3519);
nand U4361 (N_4361,N_3608,N_3753);
nor U4362 (N_4362,N_3917,N_3987);
and U4363 (N_4363,N_3908,N_3697);
xnor U4364 (N_4364,N_3897,N_3667);
and U4365 (N_4365,N_3833,N_3796);
and U4366 (N_4366,N_3903,N_3784);
or U4367 (N_4367,N_3771,N_3777);
or U4368 (N_4368,N_3721,N_3984);
nand U4369 (N_4369,N_3785,N_3889);
nor U4370 (N_4370,N_3600,N_3664);
xor U4371 (N_4371,N_3574,N_3851);
xnor U4372 (N_4372,N_3590,N_3611);
nor U4373 (N_4373,N_3858,N_3771);
nand U4374 (N_4374,N_3977,N_3731);
nand U4375 (N_4375,N_3624,N_3520);
xor U4376 (N_4376,N_3567,N_3734);
nor U4377 (N_4377,N_3738,N_3524);
and U4378 (N_4378,N_3796,N_3509);
or U4379 (N_4379,N_3804,N_3931);
or U4380 (N_4380,N_3936,N_3851);
or U4381 (N_4381,N_3822,N_3517);
or U4382 (N_4382,N_3853,N_3932);
nand U4383 (N_4383,N_3890,N_3849);
nor U4384 (N_4384,N_3676,N_3637);
nand U4385 (N_4385,N_3582,N_3894);
or U4386 (N_4386,N_3835,N_3549);
nand U4387 (N_4387,N_3631,N_3667);
xor U4388 (N_4388,N_3739,N_3556);
and U4389 (N_4389,N_3865,N_3747);
nand U4390 (N_4390,N_3669,N_3923);
or U4391 (N_4391,N_3967,N_3646);
and U4392 (N_4392,N_3506,N_3835);
xnor U4393 (N_4393,N_3884,N_3580);
or U4394 (N_4394,N_3571,N_3649);
nand U4395 (N_4395,N_3994,N_3505);
and U4396 (N_4396,N_3791,N_3507);
nor U4397 (N_4397,N_3806,N_3686);
and U4398 (N_4398,N_3659,N_3563);
nand U4399 (N_4399,N_3597,N_3803);
nand U4400 (N_4400,N_3508,N_3606);
or U4401 (N_4401,N_3762,N_3890);
nor U4402 (N_4402,N_3757,N_3656);
xor U4403 (N_4403,N_3641,N_3643);
or U4404 (N_4404,N_3642,N_3596);
or U4405 (N_4405,N_3910,N_3510);
nand U4406 (N_4406,N_3704,N_3831);
nand U4407 (N_4407,N_3757,N_3950);
or U4408 (N_4408,N_3767,N_3990);
and U4409 (N_4409,N_3735,N_3922);
and U4410 (N_4410,N_3841,N_3920);
or U4411 (N_4411,N_3692,N_3767);
nor U4412 (N_4412,N_3946,N_3951);
or U4413 (N_4413,N_3690,N_3810);
nor U4414 (N_4414,N_3887,N_3512);
nor U4415 (N_4415,N_3546,N_3623);
xor U4416 (N_4416,N_3954,N_3800);
and U4417 (N_4417,N_3699,N_3858);
and U4418 (N_4418,N_3830,N_3615);
or U4419 (N_4419,N_3877,N_3948);
and U4420 (N_4420,N_3702,N_3848);
nor U4421 (N_4421,N_3993,N_3593);
nor U4422 (N_4422,N_3524,N_3554);
nand U4423 (N_4423,N_3846,N_3611);
nor U4424 (N_4424,N_3818,N_3921);
nand U4425 (N_4425,N_3613,N_3860);
and U4426 (N_4426,N_3696,N_3544);
or U4427 (N_4427,N_3943,N_3576);
and U4428 (N_4428,N_3553,N_3531);
nor U4429 (N_4429,N_3875,N_3820);
nand U4430 (N_4430,N_3580,N_3809);
and U4431 (N_4431,N_3868,N_3602);
nor U4432 (N_4432,N_3522,N_3765);
and U4433 (N_4433,N_3733,N_3799);
or U4434 (N_4434,N_3668,N_3675);
and U4435 (N_4435,N_3596,N_3810);
nor U4436 (N_4436,N_3823,N_3691);
and U4437 (N_4437,N_3951,N_3910);
nand U4438 (N_4438,N_3967,N_3522);
xnor U4439 (N_4439,N_3921,N_3618);
or U4440 (N_4440,N_3833,N_3921);
nor U4441 (N_4441,N_3607,N_3544);
xnor U4442 (N_4442,N_3527,N_3661);
nand U4443 (N_4443,N_3986,N_3613);
and U4444 (N_4444,N_3987,N_3675);
nor U4445 (N_4445,N_3557,N_3730);
nand U4446 (N_4446,N_3889,N_3637);
or U4447 (N_4447,N_3860,N_3553);
nor U4448 (N_4448,N_3754,N_3548);
or U4449 (N_4449,N_3742,N_3860);
and U4450 (N_4450,N_3786,N_3903);
nand U4451 (N_4451,N_3581,N_3963);
or U4452 (N_4452,N_3610,N_3929);
and U4453 (N_4453,N_3873,N_3714);
and U4454 (N_4454,N_3951,N_3866);
nand U4455 (N_4455,N_3927,N_3811);
nand U4456 (N_4456,N_3796,N_3986);
nand U4457 (N_4457,N_3837,N_3706);
nand U4458 (N_4458,N_3807,N_3869);
or U4459 (N_4459,N_3619,N_3678);
and U4460 (N_4460,N_3629,N_3840);
and U4461 (N_4461,N_3983,N_3954);
or U4462 (N_4462,N_3972,N_3991);
nor U4463 (N_4463,N_3950,N_3582);
or U4464 (N_4464,N_3910,N_3767);
nand U4465 (N_4465,N_3529,N_3714);
or U4466 (N_4466,N_3649,N_3674);
and U4467 (N_4467,N_3882,N_3782);
nand U4468 (N_4468,N_3822,N_3671);
nand U4469 (N_4469,N_3926,N_3896);
xnor U4470 (N_4470,N_3829,N_3819);
nor U4471 (N_4471,N_3601,N_3974);
nand U4472 (N_4472,N_3994,N_3629);
nor U4473 (N_4473,N_3931,N_3654);
nand U4474 (N_4474,N_3624,N_3717);
nand U4475 (N_4475,N_3637,N_3556);
xor U4476 (N_4476,N_3596,N_3570);
and U4477 (N_4477,N_3605,N_3986);
nand U4478 (N_4478,N_3652,N_3765);
xor U4479 (N_4479,N_3960,N_3876);
and U4480 (N_4480,N_3945,N_3893);
or U4481 (N_4481,N_3625,N_3745);
nand U4482 (N_4482,N_3557,N_3914);
xnor U4483 (N_4483,N_3705,N_3883);
nor U4484 (N_4484,N_3809,N_3532);
nand U4485 (N_4485,N_3650,N_3947);
nor U4486 (N_4486,N_3579,N_3747);
xnor U4487 (N_4487,N_3961,N_3596);
xor U4488 (N_4488,N_3790,N_3782);
or U4489 (N_4489,N_3828,N_3502);
nand U4490 (N_4490,N_3805,N_3885);
or U4491 (N_4491,N_3933,N_3551);
or U4492 (N_4492,N_3997,N_3803);
nor U4493 (N_4493,N_3578,N_3857);
nor U4494 (N_4494,N_3923,N_3852);
or U4495 (N_4495,N_3747,N_3815);
nand U4496 (N_4496,N_3748,N_3932);
xor U4497 (N_4497,N_3927,N_3677);
and U4498 (N_4498,N_3733,N_3845);
nor U4499 (N_4499,N_3723,N_3620);
and U4500 (N_4500,N_4135,N_4238);
nor U4501 (N_4501,N_4442,N_4226);
nand U4502 (N_4502,N_4185,N_4242);
and U4503 (N_4503,N_4315,N_4471);
xor U4504 (N_4504,N_4396,N_4479);
and U4505 (N_4505,N_4455,N_4175);
and U4506 (N_4506,N_4228,N_4363);
nand U4507 (N_4507,N_4295,N_4461);
and U4508 (N_4508,N_4440,N_4209);
xor U4509 (N_4509,N_4353,N_4148);
nor U4510 (N_4510,N_4111,N_4022);
and U4511 (N_4511,N_4239,N_4345);
nand U4512 (N_4512,N_4052,N_4299);
or U4513 (N_4513,N_4311,N_4445);
nand U4514 (N_4514,N_4280,N_4160);
and U4515 (N_4515,N_4094,N_4014);
and U4516 (N_4516,N_4414,N_4253);
xnor U4517 (N_4517,N_4024,N_4478);
nor U4518 (N_4518,N_4008,N_4459);
nor U4519 (N_4519,N_4051,N_4005);
and U4520 (N_4520,N_4342,N_4402);
nand U4521 (N_4521,N_4172,N_4451);
nor U4522 (N_4522,N_4195,N_4103);
nor U4523 (N_4523,N_4153,N_4317);
nand U4524 (N_4524,N_4448,N_4174);
or U4525 (N_4525,N_4314,N_4494);
or U4526 (N_4526,N_4267,N_4450);
or U4527 (N_4527,N_4208,N_4158);
nand U4528 (N_4528,N_4431,N_4417);
nor U4529 (N_4529,N_4281,N_4370);
and U4530 (N_4530,N_4112,N_4334);
nand U4531 (N_4531,N_4198,N_4132);
nand U4532 (N_4532,N_4040,N_4410);
nor U4533 (N_4533,N_4429,N_4400);
nand U4534 (N_4534,N_4164,N_4145);
nor U4535 (N_4535,N_4187,N_4109);
and U4536 (N_4536,N_4336,N_4197);
or U4537 (N_4537,N_4288,N_4122);
nand U4538 (N_4538,N_4399,N_4229);
nand U4539 (N_4539,N_4064,N_4207);
nand U4540 (N_4540,N_4465,N_4296);
and U4541 (N_4541,N_4035,N_4029);
xnor U4542 (N_4542,N_4154,N_4021);
xor U4543 (N_4543,N_4474,N_4255);
nand U4544 (N_4544,N_4362,N_4234);
nand U4545 (N_4545,N_4201,N_4190);
or U4546 (N_4546,N_4046,N_4216);
nand U4547 (N_4547,N_4110,N_4446);
nor U4548 (N_4548,N_4140,N_4420);
and U4549 (N_4549,N_4276,N_4292);
or U4550 (N_4550,N_4277,N_4230);
xnor U4551 (N_4551,N_4305,N_4074);
or U4552 (N_4552,N_4071,N_4092);
or U4553 (N_4553,N_4133,N_4157);
nor U4554 (N_4554,N_4303,N_4388);
nor U4555 (N_4555,N_4395,N_4224);
or U4556 (N_4556,N_4275,N_4087);
nor U4557 (N_4557,N_4161,N_4423);
nand U4558 (N_4558,N_4047,N_4443);
xor U4559 (N_4559,N_4043,N_4048);
and U4560 (N_4560,N_4285,N_4301);
or U4561 (N_4561,N_4360,N_4181);
or U4562 (N_4562,N_4284,N_4248);
or U4563 (N_4563,N_4086,N_4439);
nor U4564 (N_4564,N_4031,N_4290);
nand U4565 (N_4565,N_4066,N_4485);
nor U4566 (N_4566,N_4119,N_4186);
or U4567 (N_4567,N_4368,N_4204);
nor U4568 (N_4568,N_4020,N_4231);
nor U4569 (N_4569,N_4405,N_4270);
or U4570 (N_4570,N_4467,N_4312);
nor U4571 (N_4571,N_4143,N_4347);
nand U4572 (N_4572,N_4426,N_4348);
xor U4573 (N_4573,N_4412,N_4350);
and U4574 (N_4574,N_4481,N_4010);
and U4575 (N_4575,N_4430,N_4308);
and U4576 (N_4576,N_4105,N_4261);
or U4577 (N_4577,N_4151,N_4404);
nor U4578 (N_4578,N_4482,N_4472);
nor U4579 (N_4579,N_4372,N_4165);
and U4580 (N_4580,N_4265,N_4491);
or U4581 (N_4581,N_4176,N_4406);
and U4582 (N_4582,N_4141,N_4304);
nand U4583 (N_4583,N_4069,N_4468);
or U4584 (N_4584,N_4344,N_4191);
xnor U4585 (N_4585,N_4319,N_4424);
nand U4586 (N_4586,N_4179,N_4089);
or U4587 (N_4587,N_4250,N_4326);
nor U4588 (N_4588,N_4036,N_4337);
or U4589 (N_4589,N_4294,N_4189);
xor U4590 (N_4590,N_4458,N_4203);
nand U4591 (N_4591,N_4058,N_4084);
xnor U4592 (N_4592,N_4477,N_4269);
xnor U4593 (N_4593,N_4329,N_4129);
nand U4594 (N_4594,N_4338,N_4061);
nand U4595 (N_4595,N_4435,N_4114);
nor U4596 (N_4596,N_4335,N_4194);
nor U4597 (N_4597,N_4309,N_4019);
nand U4598 (N_4598,N_4088,N_4480);
and U4599 (N_4599,N_4171,N_4168);
nand U4600 (N_4600,N_4425,N_4015);
nor U4601 (N_4601,N_4398,N_4152);
nor U4602 (N_4602,N_4196,N_4182);
and U4603 (N_4603,N_4016,N_4028);
nor U4604 (N_4604,N_4163,N_4188);
nand U4605 (N_4605,N_4053,N_4466);
nor U4606 (N_4606,N_4123,N_4422);
xnor U4607 (N_4607,N_4386,N_4042);
xor U4608 (N_4608,N_4428,N_4013);
or U4609 (N_4609,N_4436,N_4427);
and U4610 (N_4610,N_4497,N_4221);
or U4611 (N_4611,N_4018,N_4257);
nand U4612 (N_4612,N_4138,N_4392);
nand U4613 (N_4613,N_4038,N_4193);
or U4614 (N_4614,N_4127,N_4246);
nand U4615 (N_4615,N_4441,N_4279);
and U4616 (N_4616,N_4180,N_4322);
nor U4617 (N_4617,N_4159,N_4091);
xor U4618 (N_4618,N_4333,N_4062);
nor U4619 (N_4619,N_4215,N_4050);
nor U4620 (N_4620,N_4413,N_4487);
nand U4621 (N_4621,N_4218,N_4393);
or U4622 (N_4622,N_4098,N_4006);
nand U4623 (N_4623,N_4243,N_4210);
nand U4624 (N_4624,N_4009,N_4155);
or U4625 (N_4625,N_4375,N_4117);
nor U4626 (N_4626,N_4355,N_4104);
and U4627 (N_4627,N_4099,N_4365);
or U4628 (N_4628,N_4244,N_4264);
and U4629 (N_4629,N_4495,N_4356);
nand U4630 (N_4630,N_4034,N_4389);
nor U4631 (N_4631,N_4033,N_4376);
or U4632 (N_4632,N_4225,N_4340);
or U4633 (N_4633,N_4254,N_4409);
nor U4634 (N_4634,N_4093,N_4073);
and U4635 (N_4635,N_4142,N_4444);
or U4636 (N_4636,N_4469,N_4408);
or U4637 (N_4637,N_4004,N_4081);
and U4638 (N_4638,N_4083,N_4027);
and U4639 (N_4639,N_4082,N_4361);
or U4640 (N_4640,N_4212,N_4313);
nor U4641 (N_4641,N_4403,N_4102);
and U4642 (N_4642,N_4354,N_4307);
and U4643 (N_4643,N_4438,N_4045);
and U4644 (N_4644,N_4266,N_4433);
nand U4645 (N_4645,N_4249,N_4382);
and U4646 (N_4646,N_4166,N_4060);
nor U4647 (N_4647,N_4287,N_4121);
xor U4648 (N_4648,N_4156,N_4130);
nand U4649 (N_4649,N_4373,N_4177);
nor U4650 (N_4650,N_4352,N_4377);
nor U4651 (N_4651,N_4057,N_4259);
nor U4652 (N_4652,N_4025,N_4369);
nand U4653 (N_4653,N_4131,N_4067);
xor U4654 (N_4654,N_4456,N_4437);
nor U4655 (N_4655,N_4037,N_4473);
nor U4656 (N_4656,N_4418,N_4359);
or U4657 (N_4657,N_4302,N_4310);
nand U4658 (N_4658,N_4401,N_4273);
and U4659 (N_4659,N_4289,N_4460);
xnor U4660 (N_4660,N_4000,N_4002);
or U4661 (N_4661,N_4080,N_4233);
nand U4662 (N_4662,N_4351,N_4282);
and U4663 (N_4663,N_4330,N_4300);
or U4664 (N_4664,N_4054,N_4007);
nor U4665 (N_4665,N_4371,N_4049);
or U4666 (N_4666,N_4247,N_4268);
or U4667 (N_4667,N_4030,N_4260);
and U4668 (N_4668,N_4490,N_4286);
nand U4669 (N_4669,N_4026,N_4343);
xnor U4670 (N_4670,N_4379,N_4137);
or U4671 (N_4671,N_4380,N_4097);
nand U4672 (N_4672,N_4017,N_4457);
nor U4673 (N_4673,N_4278,N_4100);
or U4674 (N_4674,N_4262,N_4032);
nand U4675 (N_4675,N_4283,N_4486);
nand U4676 (N_4676,N_4381,N_4113);
or U4677 (N_4677,N_4144,N_4011);
xor U4678 (N_4678,N_4124,N_4217);
nor U4679 (N_4679,N_4044,N_4357);
nor U4680 (N_4680,N_4291,N_4251);
nor U4681 (N_4681,N_4331,N_4293);
and U4682 (N_4682,N_4252,N_4075);
and U4683 (N_4683,N_4220,N_4332);
nor U4684 (N_4684,N_4475,N_4419);
and U4685 (N_4685,N_4178,N_4055);
or U4686 (N_4686,N_4076,N_4476);
or U4687 (N_4687,N_4297,N_4235);
nor U4688 (N_4688,N_4241,N_4214);
or U4689 (N_4689,N_4454,N_4449);
nand U4690 (N_4690,N_4432,N_4434);
nand U4691 (N_4691,N_4173,N_4366);
and U4692 (N_4692,N_4390,N_4134);
and U4693 (N_4693,N_4462,N_4072);
or U4694 (N_4694,N_4323,N_4192);
nor U4695 (N_4695,N_4320,N_4183);
nand U4696 (N_4696,N_4120,N_4321);
nor U4697 (N_4697,N_4090,N_4232);
nor U4698 (N_4698,N_4452,N_4391);
nor U4699 (N_4699,N_4063,N_4498);
nor U4700 (N_4700,N_4341,N_4325);
nand U4701 (N_4701,N_4041,N_4106);
xor U4702 (N_4702,N_4318,N_4483);
nor U4703 (N_4703,N_4128,N_4077);
nor U4704 (N_4704,N_4328,N_4306);
nor U4705 (N_4705,N_4079,N_4394);
and U4706 (N_4706,N_4065,N_4378);
xor U4707 (N_4707,N_4492,N_4003);
or U4708 (N_4708,N_4385,N_4167);
nor U4709 (N_4709,N_4096,N_4205);
xnor U4710 (N_4710,N_4384,N_4447);
nor U4711 (N_4711,N_4245,N_4162);
or U4712 (N_4712,N_4339,N_4056);
nor U4713 (N_4713,N_4222,N_4199);
nor U4714 (N_4714,N_4374,N_4346);
nor U4715 (N_4715,N_4263,N_4496);
or U4716 (N_4716,N_4274,N_4316);
nand U4717 (N_4717,N_4411,N_4416);
nand U4718 (N_4718,N_4237,N_4170);
nand U4719 (N_4719,N_4146,N_4211);
and U4720 (N_4720,N_4108,N_4147);
nor U4721 (N_4721,N_4078,N_4085);
nor U4722 (N_4722,N_4407,N_4023);
and U4723 (N_4723,N_4219,N_4240);
nor U4724 (N_4724,N_4126,N_4223);
nand U4725 (N_4725,N_4236,N_4169);
or U4726 (N_4726,N_4101,N_4107);
nor U4727 (N_4727,N_4125,N_4149);
nor U4728 (N_4728,N_4484,N_4001);
or U4729 (N_4729,N_4324,N_4095);
and U4730 (N_4730,N_4364,N_4118);
nor U4731 (N_4731,N_4184,N_4383);
and U4732 (N_4732,N_4464,N_4298);
or U4733 (N_4733,N_4227,N_4453);
nor U4734 (N_4734,N_4421,N_4258);
nand U4735 (N_4735,N_4068,N_4150);
nor U4736 (N_4736,N_4387,N_4271);
nand U4737 (N_4737,N_4349,N_4488);
nor U4738 (N_4738,N_4358,N_4397);
and U4739 (N_4739,N_4202,N_4470);
or U4740 (N_4740,N_4367,N_4206);
or U4741 (N_4741,N_4059,N_4256);
nor U4742 (N_4742,N_4327,N_4136);
and U4743 (N_4743,N_4493,N_4012);
or U4744 (N_4744,N_4070,N_4415);
nand U4745 (N_4745,N_4116,N_4039);
xor U4746 (N_4746,N_4463,N_4489);
xnor U4747 (N_4747,N_4499,N_4139);
nand U4748 (N_4748,N_4115,N_4200);
or U4749 (N_4749,N_4213,N_4272);
nor U4750 (N_4750,N_4184,N_4411);
or U4751 (N_4751,N_4029,N_4444);
nand U4752 (N_4752,N_4022,N_4170);
or U4753 (N_4753,N_4460,N_4300);
xor U4754 (N_4754,N_4098,N_4430);
nor U4755 (N_4755,N_4217,N_4361);
or U4756 (N_4756,N_4070,N_4485);
and U4757 (N_4757,N_4292,N_4396);
or U4758 (N_4758,N_4119,N_4422);
nand U4759 (N_4759,N_4429,N_4130);
and U4760 (N_4760,N_4346,N_4229);
nand U4761 (N_4761,N_4024,N_4302);
nand U4762 (N_4762,N_4330,N_4175);
or U4763 (N_4763,N_4340,N_4421);
nor U4764 (N_4764,N_4160,N_4143);
nor U4765 (N_4765,N_4205,N_4100);
and U4766 (N_4766,N_4011,N_4452);
nor U4767 (N_4767,N_4212,N_4073);
xnor U4768 (N_4768,N_4324,N_4431);
and U4769 (N_4769,N_4130,N_4305);
xnor U4770 (N_4770,N_4450,N_4180);
nand U4771 (N_4771,N_4399,N_4023);
nand U4772 (N_4772,N_4328,N_4464);
or U4773 (N_4773,N_4058,N_4253);
nor U4774 (N_4774,N_4285,N_4368);
nand U4775 (N_4775,N_4032,N_4073);
xor U4776 (N_4776,N_4052,N_4035);
nor U4777 (N_4777,N_4379,N_4142);
and U4778 (N_4778,N_4012,N_4339);
and U4779 (N_4779,N_4247,N_4262);
nor U4780 (N_4780,N_4334,N_4026);
nand U4781 (N_4781,N_4384,N_4215);
nand U4782 (N_4782,N_4264,N_4240);
nand U4783 (N_4783,N_4240,N_4031);
nor U4784 (N_4784,N_4019,N_4080);
or U4785 (N_4785,N_4292,N_4349);
or U4786 (N_4786,N_4391,N_4343);
and U4787 (N_4787,N_4395,N_4139);
and U4788 (N_4788,N_4124,N_4468);
and U4789 (N_4789,N_4438,N_4183);
nand U4790 (N_4790,N_4024,N_4109);
xnor U4791 (N_4791,N_4311,N_4011);
or U4792 (N_4792,N_4292,N_4196);
and U4793 (N_4793,N_4231,N_4334);
nor U4794 (N_4794,N_4224,N_4331);
nand U4795 (N_4795,N_4250,N_4438);
nor U4796 (N_4796,N_4322,N_4476);
and U4797 (N_4797,N_4337,N_4253);
and U4798 (N_4798,N_4003,N_4008);
nor U4799 (N_4799,N_4415,N_4264);
or U4800 (N_4800,N_4191,N_4005);
and U4801 (N_4801,N_4188,N_4381);
and U4802 (N_4802,N_4121,N_4344);
nand U4803 (N_4803,N_4390,N_4259);
nor U4804 (N_4804,N_4494,N_4268);
and U4805 (N_4805,N_4229,N_4343);
xnor U4806 (N_4806,N_4005,N_4479);
nand U4807 (N_4807,N_4040,N_4340);
xor U4808 (N_4808,N_4235,N_4357);
or U4809 (N_4809,N_4280,N_4469);
nor U4810 (N_4810,N_4056,N_4047);
nand U4811 (N_4811,N_4490,N_4365);
nor U4812 (N_4812,N_4113,N_4071);
xor U4813 (N_4813,N_4216,N_4096);
nand U4814 (N_4814,N_4350,N_4121);
or U4815 (N_4815,N_4439,N_4286);
or U4816 (N_4816,N_4087,N_4082);
nand U4817 (N_4817,N_4396,N_4496);
or U4818 (N_4818,N_4126,N_4432);
and U4819 (N_4819,N_4297,N_4414);
nor U4820 (N_4820,N_4397,N_4181);
nand U4821 (N_4821,N_4443,N_4360);
or U4822 (N_4822,N_4392,N_4416);
and U4823 (N_4823,N_4299,N_4022);
or U4824 (N_4824,N_4293,N_4289);
or U4825 (N_4825,N_4497,N_4318);
and U4826 (N_4826,N_4127,N_4453);
nand U4827 (N_4827,N_4158,N_4263);
nand U4828 (N_4828,N_4242,N_4001);
nor U4829 (N_4829,N_4033,N_4480);
nor U4830 (N_4830,N_4262,N_4038);
or U4831 (N_4831,N_4197,N_4379);
or U4832 (N_4832,N_4266,N_4413);
nand U4833 (N_4833,N_4469,N_4098);
nor U4834 (N_4834,N_4020,N_4157);
nor U4835 (N_4835,N_4015,N_4381);
nor U4836 (N_4836,N_4072,N_4424);
nor U4837 (N_4837,N_4365,N_4316);
nand U4838 (N_4838,N_4203,N_4118);
nand U4839 (N_4839,N_4448,N_4012);
nand U4840 (N_4840,N_4090,N_4192);
nor U4841 (N_4841,N_4108,N_4264);
xor U4842 (N_4842,N_4135,N_4232);
and U4843 (N_4843,N_4364,N_4177);
and U4844 (N_4844,N_4299,N_4089);
nor U4845 (N_4845,N_4126,N_4307);
nor U4846 (N_4846,N_4008,N_4022);
or U4847 (N_4847,N_4231,N_4450);
nand U4848 (N_4848,N_4321,N_4401);
nand U4849 (N_4849,N_4300,N_4477);
nand U4850 (N_4850,N_4136,N_4111);
nor U4851 (N_4851,N_4409,N_4076);
or U4852 (N_4852,N_4090,N_4118);
or U4853 (N_4853,N_4114,N_4475);
nor U4854 (N_4854,N_4452,N_4314);
or U4855 (N_4855,N_4304,N_4225);
or U4856 (N_4856,N_4007,N_4499);
nor U4857 (N_4857,N_4037,N_4449);
and U4858 (N_4858,N_4379,N_4347);
xnor U4859 (N_4859,N_4112,N_4255);
and U4860 (N_4860,N_4405,N_4077);
or U4861 (N_4861,N_4120,N_4468);
or U4862 (N_4862,N_4037,N_4234);
nand U4863 (N_4863,N_4462,N_4224);
nand U4864 (N_4864,N_4408,N_4128);
nor U4865 (N_4865,N_4325,N_4411);
nand U4866 (N_4866,N_4462,N_4004);
xnor U4867 (N_4867,N_4028,N_4350);
nand U4868 (N_4868,N_4220,N_4156);
nor U4869 (N_4869,N_4002,N_4206);
nand U4870 (N_4870,N_4354,N_4213);
and U4871 (N_4871,N_4237,N_4197);
or U4872 (N_4872,N_4290,N_4047);
and U4873 (N_4873,N_4060,N_4339);
nand U4874 (N_4874,N_4450,N_4230);
or U4875 (N_4875,N_4225,N_4167);
nand U4876 (N_4876,N_4308,N_4212);
nor U4877 (N_4877,N_4013,N_4101);
or U4878 (N_4878,N_4078,N_4018);
and U4879 (N_4879,N_4387,N_4028);
xor U4880 (N_4880,N_4327,N_4393);
nor U4881 (N_4881,N_4446,N_4107);
nand U4882 (N_4882,N_4074,N_4234);
nand U4883 (N_4883,N_4187,N_4395);
and U4884 (N_4884,N_4382,N_4084);
nand U4885 (N_4885,N_4251,N_4403);
nor U4886 (N_4886,N_4179,N_4494);
and U4887 (N_4887,N_4271,N_4367);
and U4888 (N_4888,N_4218,N_4155);
nor U4889 (N_4889,N_4016,N_4011);
and U4890 (N_4890,N_4315,N_4437);
nor U4891 (N_4891,N_4086,N_4292);
nand U4892 (N_4892,N_4465,N_4197);
nor U4893 (N_4893,N_4407,N_4257);
nand U4894 (N_4894,N_4205,N_4387);
nor U4895 (N_4895,N_4165,N_4099);
or U4896 (N_4896,N_4343,N_4492);
nor U4897 (N_4897,N_4276,N_4194);
nor U4898 (N_4898,N_4121,N_4459);
xor U4899 (N_4899,N_4305,N_4480);
and U4900 (N_4900,N_4412,N_4042);
nor U4901 (N_4901,N_4452,N_4246);
nand U4902 (N_4902,N_4168,N_4488);
nand U4903 (N_4903,N_4455,N_4015);
nor U4904 (N_4904,N_4070,N_4111);
nand U4905 (N_4905,N_4187,N_4047);
or U4906 (N_4906,N_4077,N_4297);
or U4907 (N_4907,N_4204,N_4210);
xor U4908 (N_4908,N_4023,N_4374);
or U4909 (N_4909,N_4060,N_4003);
and U4910 (N_4910,N_4318,N_4258);
nand U4911 (N_4911,N_4003,N_4136);
nor U4912 (N_4912,N_4458,N_4024);
xor U4913 (N_4913,N_4339,N_4488);
nand U4914 (N_4914,N_4143,N_4387);
nor U4915 (N_4915,N_4115,N_4089);
nor U4916 (N_4916,N_4079,N_4031);
nand U4917 (N_4917,N_4445,N_4232);
xor U4918 (N_4918,N_4418,N_4211);
xnor U4919 (N_4919,N_4354,N_4381);
and U4920 (N_4920,N_4343,N_4052);
nor U4921 (N_4921,N_4024,N_4371);
nor U4922 (N_4922,N_4258,N_4174);
nand U4923 (N_4923,N_4355,N_4002);
nor U4924 (N_4924,N_4356,N_4185);
xnor U4925 (N_4925,N_4223,N_4366);
or U4926 (N_4926,N_4198,N_4193);
nor U4927 (N_4927,N_4471,N_4143);
or U4928 (N_4928,N_4072,N_4267);
or U4929 (N_4929,N_4061,N_4194);
nand U4930 (N_4930,N_4446,N_4027);
nand U4931 (N_4931,N_4157,N_4285);
and U4932 (N_4932,N_4150,N_4430);
and U4933 (N_4933,N_4282,N_4045);
and U4934 (N_4934,N_4109,N_4273);
nor U4935 (N_4935,N_4499,N_4493);
nor U4936 (N_4936,N_4307,N_4191);
nand U4937 (N_4937,N_4430,N_4329);
or U4938 (N_4938,N_4292,N_4129);
nand U4939 (N_4939,N_4194,N_4264);
and U4940 (N_4940,N_4355,N_4231);
nor U4941 (N_4941,N_4282,N_4459);
or U4942 (N_4942,N_4269,N_4054);
and U4943 (N_4943,N_4102,N_4449);
nand U4944 (N_4944,N_4491,N_4470);
or U4945 (N_4945,N_4267,N_4388);
and U4946 (N_4946,N_4125,N_4441);
nor U4947 (N_4947,N_4218,N_4342);
or U4948 (N_4948,N_4173,N_4382);
or U4949 (N_4949,N_4123,N_4201);
and U4950 (N_4950,N_4009,N_4066);
nand U4951 (N_4951,N_4499,N_4074);
nand U4952 (N_4952,N_4460,N_4422);
and U4953 (N_4953,N_4120,N_4459);
and U4954 (N_4954,N_4441,N_4494);
and U4955 (N_4955,N_4128,N_4066);
nand U4956 (N_4956,N_4132,N_4183);
or U4957 (N_4957,N_4489,N_4270);
and U4958 (N_4958,N_4304,N_4227);
and U4959 (N_4959,N_4286,N_4200);
or U4960 (N_4960,N_4383,N_4070);
and U4961 (N_4961,N_4177,N_4275);
nor U4962 (N_4962,N_4164,N_4204);
nor U4963 (N_4963,N_4046,N_4470);
nand U4964 (N_4964,N_4107,N_4498);
nand U4965 (N_4965,N_4063,N_4031);
or U4966 (N_4966,N_4251,N_4312);
xor U4967 (N_4967,N_4033,N_4136);
xnor U4968 (N_4968,N_4092,N_4276);
or U4969 (N_4969,N_4046,N_4321);
xor U4970 (N_4970,N_4142,N_4155);
nand U4971 (N_4971,N_4490,N_4380);
or U4972 (N_4972,N_4390,N_4138);
nor U4973 (N_4973,N_4409,N_4209);
nand U4974 (N_4974,N_4201,N_4319);
and U4975 (N_4975,N_4178,N_4436);
or U4976 (N_4976,N_4210,N_4470);
nor U4977 (N_4977,N_4318,N_4341);
nor U4978 (N_4978,N_4092,N_4473);
nand U4979 (N_4979,N_4227,N_4141);
nor U4980 (N_4980,N_4274,N_4183);
and U4981 (N_4981,N_4389,N_4441);
and U4982 (N_4982,N_4481,N_4357);
or U4983 (N_4983,N_4096,N_4446);
nor U4984 (N_4984,N_4186,N_4360);
and U4985 (N_4985,N_4112,N_4450);
and U4986 (N_4986,N_4279,N_4075);
and U4987 (N_4987,N_4336,N_4078);
nand U4988 (N_4988,N_4486,N_4147);
nand U4989 (N_4989,N_4442,N_4231);
or U4990 (N_4990,N_4455,N_4286);
or U4991 (N_4991,N_4354,N_4155);
or U4992 (N_4992,N_4171,N_4052);
nand U4993 (N_4993,N_4294,N_4494);
nand U4994 (N_4994,N_4321,N_4498);
and U4995 (N_4995,N_4256,N_4233);
and U4996 (N_4996,N_4267,N_4175);
or U4997 (N_4997,N_4398,N_4364);
xor U4998 (N_4998,N_4097,N_4107);
or U4999 (N_4999,N_4379,N_4159);
and UO_0 (O_0,N_4604,N_4941);
or UO_1 (O_1,N_4712,N_4779);
nand UO_2 (O_2,N_4553,N_4764);
nor UO_3 (O_3,N_4594,N_4817);
nor UO_4 (O_4,N_4916,N_4533);
nor UO_5 (O_5,N_4707,N_4685);
or UO_6 (O_6,N_4790,N_4726);
and UO_7 (O_7,N_4891,N_4954);
or UO_8 (O_8,N_4780,N_4703);
xor UO_9 (O_9,N_4737,N_4791);
and UO_10 (O_10,N_4918,N_4872);
nor UO_11 (O_11,N_4757,N_4740);
nand UO_12 (O_12,N_4605,N_4635);
nand UO_13 (O_13,N_4501,N_4673);
nand UO_14 (O_14,N_4917,N_4905);
or UO_15 (O_15,N_4567,N_4652);
nand UO_16 (O_16,N_4626,N_4627);
and UO_17 (O_17,N_4769,N_4560);
nor UO_18 (O_18,N_4534,N_4531);
or UO_19 (O_19,N_4702,N_4525);
nand UO_20 (O_20,N_4773,N_4617);
nor UO_21 (O_21,N_4730,N_4692);
and UO_22 (O_22,N_4708,N_4656);
or UO_23 (O_23,N_4913,N_4957);
or UO_24 (O_24,N_4658,N_4888);
and UO_25 (O_25,N_4661,N_4894);
or UO_26 (O_26,N_4969,N_4878);
xor UO_27 (O_27,N_4696,N_4789);
or UO_28 (O_28,N_4674,N_4812);
and UO_29 (O_29,N_4699,N_4928);
or UO_30 (O_30,N_4642,N_4947);
and UO_31 (O_31,N_4630,N_4717);
or UO_32 (O_32,N_4983,N_4677);
nor UO_33 (O_33,N_4749,N_4564);
nand UO_34 (O_34,N_4669,N_4836);
nor UO_35 (O_35,N_4896,N_4752);
xnor UO_36 (O_36,N_4676,N_4710);
and UO_37 (O_37,N_4704,N_4765);
nand UO_38 (O_38,N_4907,N_4644);
and UO_39 (O_39,N_4795,N_4990);
and UO_40 (O_40,N_4964,N_4859);
nand UO_41 (O_41,N_4915,N_4736);
xor UO_42 (O_42,N_4783,N_4648);
and UO_43 (O_43,N_4760,N_4828);
nand UO_44 (O_44,N_4753,N_4970);
and UO_45 (O_45,N_4735,N_4973);
nor UO_46 (O_46,N_4980,N_4680);
nand UO_47 (O_47,N_4848,N_4842);
and UO_48 (O_48,N_4871,N_4716);
nand UO_49 (O_49,N_4517,N_4750);
nor UO_50 (O_50,N_4550,N_4826);
xnor UO_51 (O_51,N_4886,N_4800);
or UO_52 (O_52,N_4953,N_4974);
nor UO_53 (O_53,N_4701,N_4796);
or UO_54 (O_54,N_4759,N_4774);
xnor UO_55 (O_55,N_4602,N_4761);
and UO_56 (O_56,N_4698,N_4833);
nand UO_57 (O_57,N_4768,N_4839);
xnor UO_58 (O_58,N_4874,N_4563);
and UO_59 (O_59,N_4892,N_4925);
and UO_60 (O_60,N_4679,N_4995);
or UO_61 (O_61,N_4709,N_4866);
or UO_62 (O_62,N_4863,N_4511);
and UO_63 (O_63,N_4808,N_4876);
and UO_64 (O_64,N_4621,N_4693);
nand UO_65 (O_65,N_4500,N_4612);
nor UO_66 (O_66,N_4743,N_4898);
xnor UO_67 (O_67,N_4507,N_4725);
xnor UO_68 (O_68,N_4541,N_4547);
or UO_69 (O_69,N_4587,N_4854);
or UO_70 (O_70,N_4792,N_4608);
nand UO_71 (O_71,N_4756,N_4721);
or UO_72 (O_72,N_4598,N_4829);
and UO_73 (O_73,N_4857,N_4771);
nor UO_74 (O_74,N_4806,N_4948);
or UO_75 (O_75,N_4689,N_4720);
or UO_76 (O_76,N_4639,N_4615);
or UO_77 (O_77,N_4975,N_4979);
or UO_78 (O_78,N_4816,N_4610);
and UO_79 (O_79,N_4659,N_4537);
and UO_80 (O_80,N_4629,N_4620);
nand UO_81 (O_81,N_4845,N_4824);
nand UO_82 (O_82,N_4999,N_4906);
and UO_83 (O_83,N_4867,N_4643);
nand UO_84 (O_84,N_4889,N_4847);
xor UO_85 (O_85,N_4784,N_4649);
nor UO_86 (O_86,N_4555,N_4577);
and UO_87 (O_87,N_4711,N_4967);
or UO_88 (O_88,N_4584,N_4846);
or UO_89 (O_89,N_4933,N_4997);
nand UO_90 (O_90,N_4582,N_4840);
nand UO_91 (O_91,N_4573,N_4961);
nor UO_92 (O_92,N_4879,N_4628);
nor UO_93 (O_93,N_4508,N_4744);
xnor UO_94 (O_94,N_4657,N_4922);
nor UO_95 (O_95,N_4927,N_4862);
nor UO_96 (O_96,N_4960,N_4572);
nor UO_97 (O_97,N_4742,N_4820);
nor UO_98 (O_98,N_4580,N_4632);
or UO_99 (O_99,N_4920,N_4908);
or UO_100 (O_100,N_4599,N_4776);
and UO_101 (O_101,N_4959,N_4870);
or UO_102 (O_102,N_4535,N_4601);
and UO_103 (O_103,N_4575,N_4722);
or UO_104 (O_104,N_4664,N_4884);
and UO_105 (O_105,N_4881,N_4516);
or UO_106 (O_106,N_4838,N_4528);
and UO_107 (O_107,N_4931,N_4778);
or UO_108 (O_108,N_4616,N_4714);
nand UO_109 (O_109,N_4849,N_4502);
or UO_110 (O_110,N_4640,N_4772);
nand UO_111 (O_111,N_4825,N_4641);
nor UO_112 (O_112,N_4619,N_4935);
and UO_113 (O_113,N_4586,N_4827);
or UO_114 (O_114,N_4593,N_4631);
nor UO_115 (O_115,N_4688,N_4788);
or UO_116 (O_116,N_4513,N_4561);
and UO_117 (O_117,N_4844,N_4527);
nand UO_118 (O_118,N_4767,N_4545);
xor UO_119 (O_119,N_4650,N_4943);
or UO_120 (O_120,N_4852,N_4793);
and UO_121 (O_121,N_4987,N_4900);
nor UO_122 (O_122,N_4998,N_4532);
nand UO_123 (O_123,N_4625,N_4651);
nor UO_124 (O_124,N_4645,N_4868);
and UO_125 (O_125,N_4942,N_4835);
nor UO_126 (O_126,N_4837,N_4860);
or UO_127 (O_127,N_4682,N_4733);
nand UO_128 (O_128,N_4510,N_4804);
and UO_129 (O_129,N_4924,N_4589);
and UO_130 (O_130,N_4899,N_4951);
nand UO_131 (O_131,N_4934,N_4655);
or UO_132 (O_132,N_4747,N_4543);
or UO_133 (O_133,N_4949,N_4504);
xor UO_134 (O_134,N_4554,N_4890);
nor UO_135 (O_135,N_4850,N_4719);
nor UO_136 (O_136,N_4811,N_4565);
and UO_137 (O_137,N_4962,N_4972);
and UO_138 (O_138,N_4977,N_4869);
or UO_139 (O_139,N_4993,N_4989);
nor UO_140 (O_140,N_4909,N_4996);
and UO_141 (O_141,N_4803,N_4542);
or UO_142 (O_142,N_4591,N_4821);
nand UO_143 (O_143,N_4556,N_4902);
nor UO_144 (O_144,N_4672,N_4579);
nand UO_145 (O_145,N_4777,N_4875);
and UO_146 (O_146,N_4611,N_4819);
nand UO_147 (O_147,N_4536,N_4939);
and UO_148 (O_148,N_4807,N_4665);
nor UO_149 (O_149,N_4706,N_4782);
and UO_150 (O_150,N_4914,N_4624);
nand UO_151 (O_151,N_4938,N_4988);
and UO_152 (O_152,N_4843,N_4901);
or UO_153 (O_153,N_4552,N_4919);
or UO_154 (O_154,N_4603,N_4880);
xor UO_155 (O_155,N_4971,N_4746);
or UO_156 (O_156,N_4540,N_4952);
nand UO_157 (O_157,N_4984,N_4723);
nand UO_158 (O_158,N_4955,N_4945);
xnor UO_159 (O_159,N_4524,N_4690);
nand UO_160 (O_160,N_4815,N_4576);
and UO_161 (O_161,N_4936,N_4530);
nand UO_162 (O_162,N_4570,N_4618);
or UO_163 (O_163,N_4958,N_4566);
or UO_164 (O_164,N_4581,N_4622);
and UO_165 (O_165,N_4520,N_4583);
nand UO_166 (O_166,N_4754,N_4956);
xnor UO_167 (O_167,N_4739,N_4666);
nor UO_168 (O_168,N_4653,N_4623);
nor UO_169 (O_169,N_4663,N_4697);
and UO_170 (O_170,N_4614,N_4683);
or UO_171 (O_171,N_4992,N_4686);
and UO_172 (O_172,N_4841,N_4813);
xnor UO_173 (O_173,N_4763,N_4748);
nand UO_174 (O_174,N_4985,N_4512);
nand UO_175 (O_175,N_4590,N_4882);
nor UO_176 (O_176,N_4910,N_4526);
nor UO_177 (O_177,N_4932,N_4607);
nand UO_178 (O_178,N_4861,N_4687);
nor UO_179 (O_179,N_4731,N_4681);
nand UO_180 (O_180,N_4691,N_4728);
or UO_181 (O_181,N_4718,N_4991);
nand UO_182 (O_182,N_4670,N_4798);
nor UO_183 (O_183,N_4600,N_4660);
nor UO_184 (O_184,N_4794,N_4770);
or UO_185 (O_185,N_4893,N_4781);
nor UO_186 (O_186,N_4865,N_4592);
nand UO_187 (O_187,N_4548,N_4797);
or UO_188 (O_188,N_4732,N_4700);
nor UO_189 (O_189,N_4671,N_4814);
and UO_190 (O_190,N_4810,N_4705);
or UO_191 (O_191,N_4831,N_4544);
nor UO_192 (O_192,N_4982,N_4923);
xor UO_193 (O_193,N_4557,N_4647);
or UO_194 (O_194,N_4522,N_4968);
nor UO_195 (O_195,N_4523,N_4562);
and UO_196 (O_196,N_4911,N_4775);
nor UO_197 (O_197,N_4864,N_4741);
or UO_198 (O_198,N_4823,N_4514);
nand UO_199 (O_199,N_4727,N_4521);
and UO_200 (O_200,N_4937,N_4976);
xor UO_201 (O_201,N_4518,N_4981);
nand UO_202 (O_202,N_4638,N_4802);
nand UO_203 (O_203,N_4904,N_4745);
and UO_204 (O_204,N_4574,N_4529);
and UO_205 (O_205,N_4595,N_4654);
nor UO_206 (O_206,N_4853,N_4832);
nand UO_207 (O_207,N_4978,N_4897);
and UO_208 (O_208,N_4786,N_4950);
nand UO_209 (O_209,N_4636,N_4662);
nand UO_210 (O_210,N_4766,N_4609);
nor UO_211 (O_211,N_4569,N_4559);
or UO_212 (O_212,N_4912,N_4538);
or UO_213 (O_213,N_4503,N_4506);
nor UO_214 (O_214,N_4873,N_4946);
and UO_215 (O_215,N_4637,N_4588);
or UO_216 (O_216,N_4519,N_4965);
nand UO_217 (O_217,N_4578,N_4684);
nor UO_218 (O_218,N_4885,N_4539);
nor UO_219 (O_219,N_4856,N_4613);
nor UO_220 (O_220,N_4877,N_4509);
nand UO_221 (O_221,N_4830,N_4549);
and UO_222 (O_222,N_4738,N_4986);
or UO_223 (O_223,N_4505,N_4675);
or UO_224 (O_224,N_4646,N_4887);
xnor UO_225 (O_225,N_4822,N_4585);
nor UO_226 (O_226,N_4818,N_4963);
or UO_227 (O_227,N_4551,N_4633);
or UO_228 (O_228,N_4558,N_4903);
nor UO_229 (O_229,N_4713,N_4805);
nand UO_230 (O_230,N_4921,N_4929);
or UO_231 (O_231,N_4809,N_4596);
or UO_232 (O_232,N_4724,N_4667);
xnor UO_233 (O_233,N_4966,N_4895);
xor UO_234 (O_234,N_4678,N_4762);
xnor UO_235 (O_235,N_4940,N_4851);
nand UO_236 (O_236,N_4546,N_4568);
xnor UO_237 (O_237,N_4944,N_4755);
nor UO_238 (O_238,N_4930,N_4787);
and UO_239 (O_239,N_4515,N_4734);
nor UO_240 (O_240,N_4855,N_4751);
nor UO_241 (O_241,N_4785,N_4597);
or UO_242 (O_242,N_4799,N_4834);
or UO_243 (O_243,N_4606,N_4883);
or UO_244 (O_244,N_4858,N_4668);
nand UO_245 (O_245,N_4801,N_4758);
nor UO_246 (O_246,N_4571,N_4994);
xnor UO_247 (O_247,N_4634,N_4926);
nand UO_248 (O_248,N_4715,N_4695);
nor UO_249 (O_249,N_4694,N_4729);
nor UO_250 (O_250,N_4891,N_4776);
nand UO_251 (O_251,N_4668,N_4682);
nand UO_252 (O_252,N_4706,N_4808);
nor UO_253 (O_253,N_4616,N_4709);
nand UO_254 (O_254,N_4822,N_4720);
and UO_255 (O_255,N_4756,N_4987);
nand UO_256 (O_256,N_4759,N_4559);
nor UO_257 (O_257,N_4779,N_4965);
and UO_258 (O_258,N_4934,N_4502);
and UO_259 (O_259,N_4808,N_4585);
or UO_260 (O_260,N_4692,N_4599);
and UO_261 (O_261,N_4646,N_4751);
and UO_262 (O_262,N_4924,N_4550);
or UO_263 (O_263,N_4995,N_4885);
xnor UO_264 (O_264,N_4757,N_4707);
nor UO_265 (O_265,N_4539,N_4847);
nor UO_266 (O_266,N_4724,N_4549);
nor UO_267 (O_267,N_4610,N_4990);
and UO_268 (O_268,N_4716,N_4596);
nand UO_269 (O_269,N_4688,N_4779);
nor UO_270 (O_270,N_4775,N_4724);
nand UO_271 (O_271,N_4971,N_4934);
nand UO_272 (O_272,N_4810,N_4861);
and UO_273 (O_273,N_4795,N_4808);
and UO_274 (O_274,N_4749,N_4694);
or UO_275 (O_275,N_4646,N_4731);
nand UO_276 (O_276,N_4931,N_4782);
and UO_277 (O_277,N_4728,N_4697);
nand UO_278 (O_278,N_4729,N_4590);
or UO_279 (O_279,N_4553,N_4657);
and UO_280 (O_280,N_4638,N_4782);
xnor UO_281 (O_281,N_4550,N_4869);
nor UO_282 (O_282,N_4938,N_4864);
nor UO_283 (O_283,N_4891,N_4607);
or UO_284 (O_284,N_4610,N_4983);
or UO_285 (O_285,N_4952,N_4811);
nor UO_286 (O_286,N_4773,N_4833);
nor UO_287 (O_287,N_4955,N_4671);
nand UO_288 (O_288,N_4970,N_4781);
xor UO_289 (O_289,N_4923,N_4651);
or UO_290 (O_290,N_4527,N_4783);
nor UO_291 (O_291,N_4745,N_4666);
nand UO_292 (O_292,N_4837,N_4840);
or UO_293 (O_293,N_4820,N_4931);
nand UO_294 (O_294,N_4902,N_4687);
and UO_295 (O_295,N_4915,N_4602);
nand UO_296 (O_296,N_4626,N_4817);
and UO_297 (O_297,N_4838,N_4834);
nor UO_298 (O_298,N_4963,N_4903);
nor UO_299 (O_299,N_4795,N_4824);
nand UO_300 (O_300,N_4517,N_4911);
nand UO_301 (O_301,N_4816,N_4563);
nand UO_302 (O_302,N_4523,N_4646);
and UO_303 (O_303,N_4690,N_4912);
xnor UO_304 (O_304,N_4626,N_4931);
nand UO_305 (O_305,N_4850,N_4933);
and UO_306 (O_306,N_4750,N_4669);
nand UO_307 (O_307,N_4833,N_4658);
nand UO_308 (O_308,N_4617,N_4777);
nor UO_309 (O_309,N_4808,N_4749);
nand UO_310 (O_310,N_4701,N_4501);
xnor UO_311 (O_311,N_4769,N_4742);
nor UO_312 (O_312,N_4612,N_4698);
xor UO_313 (O_313,N_4690,N_4806);
or UO_314 (O_314,N_4982,N_4555);
or UO_315 (O_315,N_4871,N_4583);
and UO_316 (O_316,N_4994,N_4538);
and UO_317 (O_317,N_4925,N_4968);
or UO_318 (O_318,N_4880,N_4530);
and UO_319 (O_319,N_4959,N_4764);
nor UO_320 (O_320,N_4750,N_4962);
and UO_321 (O_321,N_4914,N_4652);
nand UO_322 (O_322,N_4787,N_4651);
and UO_323 (O_323,N_4668,N_4586);
nand UO_324 (O_324,N_4988,N_4963);
nand UO_325 (O_325,N_4770,N_4590);
or UO_326 (O_326,N_4702,N_4615);
or UO_327 (O_327,N_4671,N_4689);
nand UO_328 (O_328,N_4536,N_4675);
or UO_329 (O_329,N_4553,N_4662);
and UO_330 (O_330,N_4909,N_4906);
nor UO_331 (O_331,N_4833,N_4951);
or UO_332 (O_332,N_4764,N_4801);
nor UO_333 (O_333,N_4593,N_4930);
and UO_334 (O_334,N_4579,N_4554);
or UO_335 (O_335,N_4637,N_4535);
nor UO_336 (O_336,N_4751,N_4621);
nand UO_337 (O_337,N_4699,N_4713);
or UO_338 (O_338,N_4642,N_4650);
or UO_339 (O_339,N_4752,N_4957);
nor UO_340 (O_340,N_4580,N_4699);
nor UO_341 (O_341,N_4605,N_4662);
or UO_342 (O_342,N_4999,N_4837);
and UO_343 (O_343,N_4883,N_4860);
nor UO_344 (O_344,N_4626,N_4693);
nand UO_345 (O_345,N_4972,N_4931);
nand UO_346 (O_346,N_4527,N_4851);
and UO_347 (O_347,N_4596,N_4980);
nand UO_348 (O_348,N_4633,N_4808);
nor UO_349 (O_349,N_4858,N_4582);
nand UO_350 (O_350,N_4551,N_4959);
xor UO_351 (O_351,N_4780,N_4528);
nand UO_352 (O_352,N_4611,N_4728);
xnor UO_353 (O_353,N_4637,N_4819);
xnor UO_354 (O_354,N_4568,N_4569);
nor UO_355 (O_355,N_4794,N_4837);
and UO_356 (O_356,N_4859,N_4785);
and UO_357 (O_357,N_4516,N_4897);
or UO_358 (O_358,N_4530,N_4839);
and UO_359 (O_359,N_4761,N_4956);
or UO_360 (O_360,N_4609,N_4974);
xor UO_361 (O_361,N_4900,N_4797);
nand UO_362 (O_362,N_4818,N_4830);
nor UO_363 (O_363,N_4645,N_4865);
and UO_364 (O_364,N_4517,N_4864);
and UO_365 (O_365,N_4612,N_4950);
nor UO_366 (O_366,N_4710,N_4742);
and UO_367 (O_367,N_4831,N_4595);
nand UO_368 (O_368,N_4502,N_4726);
nand UO_369 (O_369,N_4542,N_4789);
and UO_370 (O_370,N_4952,N_4528);
or UO_371 (O_371,N_4737,N_4898);
or UO_372 (O_372,N_4856,N_4894);
nor UO_373 (O_373,N_4840,N_4547);
nand UO_374 (O_374,N_4948,N_4624);
nand UO_375 (O_375,N_4610,N_4718);
nand UO_376 (O_376,N_4844,N_4912);
and UO_377 (O_377,N_4800,N_4749);
nor UO_378 (O_378,N_4687,N_4626);
or UO_379 (O_379,N_4752,N_4771);
and UO_380 (O_380,N_4538,N_4651);
nor UO_381 (O_381,N_4968,N_4839);
and UO_382 (O_382,N_4529,N_4501);
nor UO_383 (O_383,N_4734,N_4547);
nand UO_384 (O_384,N_4701,N_4936);
or UO_385 (O_385,N_4798,N_4593);
and UO_386 (O_386,N_4813,N_4915);
nand UO_387 (O_387,N_4882,N_4808);
nand UO_388 (O_388,N_4875,N_4961);
xnor UO_389 (O_389,N_4859,N_4898);
nand UO_390 (O_390,N_4643,N_4572);
nand UO_391 (O_391,N_4668,N_4729);
and UO_392 (O_392,N_4968,N_4689);
nor UO_393 (O_393,N_4719,N_4651);
nand UO_394 (O_394,N_4693,N_4511);
or UO_395 (O_395,N_4828,N_4730);
nand UO_396 (O_396,N_4554,N_4652);
nand UO_397 (O_397,N_4505,N_4859);
nand UO_398 (O_398,N_4689,N_4840);
nand UO_399 (O_399,N_4621,N_4913);
nor UO_400 (O_400,N_4576,N_4677);
nor UO_401 (O_401,N_4583,N_4540);
and UO_402 (O_402,N_4941,N_4643);
nand UO_403 (O_403,N_4791,N_4884);
nor UO_404 (O_404,N_4964,N_4929);
nor UO_405 (O_405,N_4761,N_4989);
and UO_406 (O_406,N_4788,N_4699);
nor UO_407 (O_407,N_4629,N_4944);
xor UO_408 (O_408,N_4792,N_4854);
and UO_409 (O_409,N_4766,N_4607);
and UO_410 (O_410,N_4917,N_4872);
xnor UO_411 (O_411,N_4827,N_4837);
nor UO_412 (O_412,N_4965,N_4685);
nand UO_413 (O_413,N_4666,N_4819);
or UO_414 (O_414,N_4748,N_4874);
and UO_415 (O_415,N_4745,N_4810);
nand UO_416 (O_416,N_4669,N_4590);
xnor UO_417 (O_417,N_4713,N_4994);
and UO_418 (O_418,N_4873,N_4674);
or UO_419 (O_419,N_4700,N_4791);
and UO_420 (O_420,N_4833,N_4997);
and UO_421 (O_421,N_4671,N_4989);
or UO_422 (O_422,N_4811,N_4630);
and UO_423 (O_423,N_4654,N_4625);
or UO_424 (O_424,N_4990,N_4759);
or UO_425 (O_425,N_4912,N_4899);
nand UO_426 (O_426,N_4570,N_4720);
or UO_427 (O_427,N_4624,N_4533);
or UO_428 (O_428,N_4623,N_4730);
nor UO_429 (O_429,N_4714,N_4915);
nand UO_430 (O_430,N_4613,N_4547);
nand UO_431 (O_431,N_4555,N_4633);
nand UO_432 (O_432,N_4730,N_4707);
nand UO_433 (O_433,N_4957,N_4631);
xnor UO_434 (O_434,N_4921,N_4547);
nand UO_435 (O_435,N_4639,N_4901);
nand UO_436 (O_436,N_4741,N_4912);
xor UO_437 (O_437,N_4669,N_4614);
nor UO_438 (O_438,N_4558,N_4665);
nand UO_439 (O_439,N_4852,N_4567);
nor UO_440 (O_440,N_4540,N_4969);
or UO_441 (O_441,N_4787,N_4866);
or UO_442 (O_442,N_4895,N_4583);
nand UO_443 (O_443,N_4883,N_4550);
or UO_444 (O_444,N_4561,N_4949);
xnor UO_445 (O_445,N_4502,N_4532);
and UO_446 (O_446,N_4670,N_4535);
nand UO_447 (O_447,N_4855,N_4599);
or UO_448 (O_448,N_4973,N_4613);
and UO_449 (O_449,N_4832,N_4943);
nor UO_450 (O_450,N_4992,N_4673);
nor UO_451 (O_451,N_4892,N_4606);
or UO_452 (O_452,N_4704,N_4899);
nand UO_453 (O_453,N_4584,N_4751);
xor UO_454 (O_454,N_4659,N_4892);
nor UO_455 (O_455,N_4654,N_4665);
xor UO_456 (O_456,N_4569,N_4857);
and UO_457 (O_457,N_4906,N_4976);
and UO_458 (O_458,N_4808,N_4649);
or UO_459 (O_459,N_4936,N_4665);
and UO_460 (O_460,N_4559,N_4562);
nand UO_461 (O_461,N_4625,N_4605);
nand UO_462 (O_462,N_4802,N_4750);
or UO_463 (O_463,N_4614,N_4832);
nand UO_464 (O_464,N_4522,N_4828);
nand UO_465 (O_465,N_4790,N_4835);
nor UO_466 (O_466,N_4876,N_4827);
xnor UO_467 (O_467,N_4967,N_4893);
nand UO_468 (O_468,N_4902,N_4508);
nand UO_469 (O_469,N_4638,N_4741);
and UO_470 (O_470,N_4692,N_4988);
and UO_471 (O_471,N_4683,N_4905);
nor UO_472 (O_472,N_4584,N_4632);
nor UO_473 (O_473,N_4513,N_4886);
and UO_474 (O_474,N_4725,N_4639);
nor UO_475 (O_475,N_4897,N_4573);
and UO_476 (O_476,N_4802,N_4889);
or UO_477 (O_477,N_4573,N_4918);
nor UO_478 (O_478,N_4932,N_4892);
nand UO_479 (O_479,N_4952,N_4598);
or UO_480 (O_480,N_4569,N_4616);
nor UO_481 (O_481,N_4923,N_4586);
nand UO_482 (O_482,N_4902,N_4814);
nand UO_483 (O_483,N_4518,N_4509);
or UO_484 (O_484,N_4947,N_4892);
nand UO_485 (O_485,N_4902,N_4580);
xor UO_486 (O_486,N_4963,N_4823);
nand UO_487 (O_487,N_4988,N_4686);
xnor UO_488 (O_488,N_4588,N_4724);
and UO_489 (O_489,N_4709,N_4527);
and UO_490 (O_490,N_4945,N_4908);
and UO_491 (O_491,N_4991,N_4602);
nand UO_492 (O_492,N_4726,N_4784);
nor UO_493 (O_493,N_4718,N_4852);
and UO_494 (O_494,N_4529,N_4939);
or UO_495 (O_495,N_4995,N_4807);
and UO_496 (O_496,N_4539,N_4767);
nor UO_497 (O_497,N_4792,N_4924);
or UO_498 (O_498,N_4654,N_4579);
nor UO_499 (O_499,N_4988,N_4604);
or UO_500 (O_500,N_4959,N_4822);
nand UO_501 (O_501,N_4543,N_4877);
or UO_502 (O_502,N_4573,N_4991);
nand UO_503 (O_503,N_4899,N_4583);
and UO_504 (O_504,N_4612,N_4630);
and UO_505 (O_505,N_4946,N_4718);
nor UO_506 (O_506,N_4661,N_4632);
nand UO_507 (O_507,N_4950,N_4772);
and UO_508 (O_508,N_4902,N_4810);
xor UO_509 (O_509,N_4500,N_4861);
and UO_510 (O_510,N_4838,N_4881);
or UO_511 (O_511,N_4609,N_4727);
or UO_512 (O_512,N_4608,N_4582);
nor UO_513 (O_513,N_4566,N_4648);
and UO_514 (O_514,N_4680,N_4566);
nor UO_515 (O_515,N_4714,N_4800);
and UO_516 (O_516,N_4514,N_4881);
and UO_517 (O_517,N_4664,N_4965);
or UO_518 (O_518,N_4999,N_4522);
and UO_519 (O_519,N_4596,N_4556);
nor UO_520 (O_520,N_4868,N_4533);
xor UO_521 (O_521,N_4977,N_4901);
nor UO_522 (O_522,N_4663,N_4677);
nand UO_523 (O_523,N_4808,N_4889);
nor UO_524 (O_524,N_4901,N_4535);
nand UO_525 (O_525,N_4707,N_4997);
and UO_526 (O_526,N_4725,N_4938);
nor UO_527 (O_527,N_4807,N_4895);
nor UO_528 (O_528,N_4821,N_4576);
nand UO_529 (O_529,N_4811,N_4878);
and UO_530 (O_530,N_4567,N_4600);
nand UO_531 (O_531,N_4612,N_4687);
nand UO_532 (O_532,N_4825,N_4801);
and UO_533 (O_533,N_4642,N_4552);
or UO_534 (O_534,N_4736,N_4686);
and UO_535 (O_535,N_4983,N_4860);
nor UO_536 (O_536,N_4997,N_4756);
and UO_537 (O_537,N_4910,N_4876);
nor UO_538 (O_538,N_4668,N_4929);
nor UO_539 (O_539,N_4869,N_4752);
nand UO_540 (O_540,N_4980,N_4967);
and UO_541 (O_541,N_4515,N_4907);
nor UO_542 (O_542,N_4798,N_4682);
xor UO_543 (O_543,N_4675,N_4602);
and UO_544 (O_544,N_4829,N_4571);
nand UO_545 (O_545,N_4865,N_4821);
nor UO_546 (O_546,N_4865,N_4662);
and UO_547 (O_547,N_4773,N_4692);
and UO_548 (O_548,N_4930,N_4951);
nand UO_549 (O_549,N_4767,N_4649);
nand UO_550 (O_550,N_4518,N_4508);
xor UO_551 (O_551,N_4637,N_4907);
and UO_552 (O_552,N_4623,N_4593);
and UO_553 (O_553,N_4829,N_4957);
nand UO_554 (O_554,N_4755,N_4766);
and UO_555 (O_555,N_4788,N_4579);
nand UO_556 (O_556,N_4814,N_4920);
nor UO_557 (O_557,N_4924,N_4821);
xnor UO_558 (O_558,N_4603,N_4848);
or UO_559 (O_559,N_4884,N_4868);
and UO_560 (O_560,N_4810,N_4828);
xnor UO_561 (O_561,N_4987,N_4705);
nand UO_562 (O_562,N_4517,N_4642);
xor UO_563 (O_563,N_4985,N_4924);
or UO_564 (O_564,N_4554,N_4929);
and UO_565 (O_565,N_4712,N_4630);
or UO_566 (O_566,N_4886,N_4596);
nor UO_567 (O_567,N_4705,N_4528);
nor UO_568 (O_568,N_4947,N_4780);
or UO_569 (O_569,N_4823,N_4529);
nand UO_570 (O_570,N_4922,N_4929);
nand UO_571 (O_571,N_4718,N_4771);
or UO_572 (O_572,N_4518,N_4608);
or UO_573 (O_573,N_4805,N_4925);
and UO_574 (O_574,N_4845,N_4551);
and UO_575 (O_575,N_4778,N_4877);
or UO_576 (O_576,N_4677,N_4977);
and UO_577 (O_577,N_4571,N_4865);
or UO_578 (O_578,N_4781,N_4849);
nor UO_579 (O_579,N_4916,N_4675);
nor UO_580 (O_580,N_4708,N_4962);
xnor UO_581 (O_581,N_4826,N_4799);
xor UO_582 (O_582,N_4723,N_4694);
nor UO_583 (O_583,N_4762,N_4932);
or UO_584 (O_584,N_4787,N_4921);
xnor UO_585 (O_585,N_4966,N_4720);
nand UO_586 (O_586,N_4727,N_4859);
nand UO_587 (O_587,N_4745,N_4669);
and UO_588 (O_588,N_4587,N_4736);
xnor UO_589 (O_589,N_4769,N_4631);
and UO_590 (O_590,N_4827,N_4564);
nand UO_591 (O_591,N_4869,N_4764);
nor UO_592 (O_592,N_4558,N_4545);
nor UO_593 (O_593,N_4883,N_4535);
and UO_594 (O_594,N_4858,N_4520);
or UO_595 (O_595,N_4793,N_4611);
and UO_596 (O_596,N_4662,N_4539);
and UO_597 (O_597,N_4878,N_4815);
nand UO_598 (O_598,N_4647,N_4823);
and UO_599 (O_599,N_4562,N_4745);
nor UO_600 (O_600,N_4869,N_4656);
or UO_601 (O_601,N_4586,N_4689);
and UO_602 (O_602,N_4626,N_4789);
and UO_603 (O_603,N_4869,N_4792);
nand UO_604 (O_604,N_4567,N_4849);
and UO_605 (O_605,N_4524,N_4886);
and UO_606 (O_606,N_4687,N_4874);
and UO_607 (O_607,N_4730,N_4502);
nor UO_608 (O_608,N_4692,N_4656);
xor UO_609 (O_609,N_4865,N_4788);
or UO_610 (O_610,N_4530,N_4828);
or UO_611 (O_611,N_4980,N_4505);
nor UO_612 (O_612,N_4867,N_4725);
and UO_613 (O_613,N_4615,N_4913);
or UO_614 (O_614,N_4733,N_4539);
nand UO_615 (O_615,N_4852,N_4765);
nor UO_616 (O_616,N_4751,N_4514);
and UO_617 (O_617,N_4591,N_4536);
nor UO_618 (O_618,N_4659,N_4746);
nor UO_619 (O_619,N_4767,N_4630);
or UO_620 (O_620,N_4664,N_4592);
xnor UO_621 (O_621,N_4513,N_4789);
and UO_622 (O_622,N_4744,N_4614);
or UO_623 (O_623,N_4799,N_4944);
nand UO_624 (O_624,N_4591,N_4914);
nand UO_625 (O_625,N_4597,N_4536);
nand UO_626 (O_626,N_4567,N_4584);
nand UO_627 (O_627,N_4630,N_4813);
nor UO_628 (O_628,N_4581,N_4560);
nand UO_629 (O_629,N_4525,N_4582);
xnor UO_630 (O_630,N_4853,N_4651);
nand UO_631 (O_631,N_4612,N_4853);
nand UO_632 (O_632,N_4686,N_4891);
and UO_633 (O_633,N_4632,N_4919);
or UO_634 (O_634,N_4547,N_4612);
or UO_635 (O_635,N_4902,N_4897);
nor UO_636 (O_636,N_4783,N_4915);
nor UO_637 (O_637,N_4897,N_4590);
nor UO_638 (O_638,N_4898,N_4921);
and UO_639 (O_639,N_4697,N_4941);
nor UO_640 (O_640,N_4693,N_4694);
or UO_641 (O_641,N_4635,N_4514);
and UO_642 (O_642,N_4978,N_4650);
or UO_643 (O_643,N_4914,N_4530);
and UO_644 (O_644,N_4727,N_4671);
and UO_645 (O_645,N_4841,N_4806);
or UO_646 (O_646,N_4615,N_4762);
nor UO_647 (O_647,N_4706,N_4680);
nand UO_648 (O_648,N_4909,N_4502);
nand UO_649 (O_649,N_4562,N_4898);
and UO_650 (O_650,N_4935,N_4860);
or UO_651 (O_651,N_4643,N_4994);
xnor UO_652 (O_652,N_4598,N_4523);
or UO_653 (O_653,N_4901,N_4997);
nor UO_654 (O_654,N_4850,N_4888);
or UO_655 (O_655,N_4986,N_4612);
nand UO_656 (O_656,N_4553,N_4701);
nand UO_657 (O_657,N_4574,N_4873);
or UO_658 (O_658,N_4630,N_4636);
or UO_659 (O_659,N_4938,N_4781);
and UO_660 (O_660,N_4586,N_4654);
nor UO_661 (O_661,N_4873,N_4973);
nand UO_662 (O_662,N_4777,N_4697);
or UO_663 (O_663,N_4520,N_4781);
nand UO_664 (O_664,N_4900,N_4808);
nand UO_665 (O_665,N_4923,N_4926);
nand UO_666 (O_666,N_4636,N_4947);
or UO_667 (O_667,N_4541,N_4712);
nor UO_668 (O_668,N_4884,N_4504);
nand UO_669 (O_669,N_4817,N_4787);
xor UO_670 (O_670,N_4519,N_4662);
or UO_671 (O_671,N_4597,N_4629);
or UO_672 (O_672,N_4618,N_4968);
and UO_673 (O_673,N_4794,N_4851);
or UO_674 (O_674,N_4903,N_4508);
and UO_675 (O_675,N_4752,N_4746);
xnor UO_676 (O_676,N_4919,N_4530);
or UO_677 (O_677,N_4949,N_4757);
nand UO_678 (O_678,N_4873,N_4558);
and UO_679 (O_679,N_4695,N_4541);
xnor UO_680 (O_680,N_4881,N_4868);
and UO_681 (O_681,N_4901,N_4728);
and UO_682 (O_682,N_4593,N_4965);
and UO_683 (O_683,N_4718,N_4593);
xnor UO_684 (O_684,N_4882,N_4651);
or UO_685 (O_685,N_4617,N_4907);
nand UO_686 (O_686,N_4749,N_4638);
nor UO_687 (O_687,N_4887,N_4953);
or UO_688 (O_688,N_4626,N_4968);
or UO_689 (O_689,N_4506,N_4750);
nand UO_690 (O_690,N_4773,N_4760);
or UO_691 (O_691,N_4502,N_4754);
nor UO_692 (O_692,N_4817,N_4559);
or UO_693 (O_693,N_4750,N_4702);
xor UO_694 (O_694,N_4923,N_4726);
nand UO_695 (O_695,N_4705,N_4924);
or UO_696 (O_696,N_4697,N_4987);
or UO_697 (O_697,N_4584,N_4843);
and UO_698 (O_698,N_4712,N_4543);
xor UO_699 (O_699,N_4650,N_4557);
nand UO_700 (O_700,N_4687,N_4762);
nand UO_701 (O_701,N_4645,N_4802);
and UO_702 (O_702,N_4641,N_4650);
or UO_703 (O_703,N_4996,N_4653);
and UO_704 (O_704,N_4882,N_4552);
or UO_705 (O_705,N_4623,N_4921);
nand UO_706 (O_706,N_4831,N_4524);
nor UO_707 (O_707,N_4925,N_4766);
or UO_708 (O_708,N_4722,N_4745);
nor UO_709 (O_709,N_4850,N_4874);
nand UO_710 (O_710,N_4855,N_4793);
and UO_711 (O_711,N_4645,N_4801);
and UO_712 (O_712,N_4701,N_4837);
nor UO_713 (O_713,N_4769,N_4763);
and UO_714 (O_714,N_4805,N_4897);
and UO_715 (O_715,N_4724,N_4776);
nor UO_716 (O_716,N_4910,N_4823);
nand UO_717 (O_717,N_4775,N_4676);
nand UO_718 (O_718,N_4994,N_4503);
nor UO_719 (O_719,N_4654,N_4712);
or UO_720 (O_720,N_4662,N_4943);
or UO_721 (O_721,N_4958,N_4983);
and UO_722 (O_722,N_4974,N_4796);
nor UO_723 (O_723,N_4919,N_4577);
and UO_724 (O_724,N_4752,N_4661);
xor UO_725 (O_725,N_4519,N_4895);
nand UO_726 (O_726,N_4908,N_4584);
nor UO_727 (O_727,N_4841,N_4887);
or UO_728 (O_728,N_4682,N_4945);
or UO_729 (O_729,N_4803,N_4962);
nand UO_730 (O_730,N_4739,N_4976);
nor UO_731 (O_731,N_4627,N_4608);
and UO_732 (O_732,N_4643,N_4799);
and UO_733 (O_733,N_4597,N_4796);
and UO_734 (O_734,N_4948,N_4636);
xnor UO_735 (O_735,N_4809,N_4989);
nor UO_736 (O_736,N_4846,N_4757);
nor UO_737 (O_737,N_4655,N_4706);
or UO_738 (O_738,N_4673,N_4927);
or UO_739 (O_739,N_4692,N_4902);
nor UO_740 (O_740,N_4650,N_4965);
nor UO_741 (O_741,N_4896,N_4517);
nor UO_742 (O_742,N_4930,N_4505);
nor UO_743 (O_743,N_4693,N_4671);
nand UO_744 (O_744,N_4776,N_4751);
or UO_745 (O_745,N_4594,N_4505);
nand UO_746 (O_746,N_4536,N_4919);
or UO_747 (O_747,N_4699,N_4771);
and UO_748 (O_748,N_4927,N_4816);
nor UO_749 (O_749,N_4993,N_4755);
and UO_750 (O_750,N_4977,N_4884);
and UO_751 (O_751,N_4928,N_4670);
or UO_752 (O_752,N_4911,N_4871);
nor UO_753 (O_753,N_4807,N_4884);
or UO_754 (O_754,N_4691,N_4913);
and UO_755 (O_755,N_4826,N_4764);
nor UO_756 (O_756,N_4675,N_4872);
and UO_757 (O_757,N_4773,N_4966);
or UO_758 (O_758,N_4782,N_4852);
and UO_759 (O_759,N_4529,N_4954);
xor UO_760 (O_760,N_4564,N_4542);
xor UO_761 (O_761,N_4806,N_4662);
and UO_762 (O_762,N_4601,N_4934);
nand UO_763 (O_763,N_4653,N_4691);
nand UO_764 (O_764,N_4951,N_4921);
nor UO_765 (O_765,N_4613,N_4686);
or UO_766 (O_766,N_4596,N_4723);
and UO_767 (O_767,N_4513,N_4731);
nand UO_768 (O_768,N_4954,N_4661);
nand UO_769 (O_769,N_4571,N_4731);
xnor UO_770 (O_770,N_4763,N_4961);
xor UO_771 (O_771,N_4594,N_4718);
xnor UO_772 (O_772,N_4626,N_4623);
nor UO_773 (O_773,N_4558,N_4876);
nor UO_774 (O_774,N_4604,N_4620);
nor UO_775 (O_775,N_4691,N_4552);
nor UO_776 (O_776,N_4907,N_4566);
or UO_777 (O_777,N_4615,N_4979);
nand UO_778 (O_778,N_4722,N_4859);
nor UO_779 (O_779,N_4715,N_4679);
nand UO_780 (O_780,N_4959,N_4648);
and UO_781 (O_781,N_4904,N_4796);
and UO_782 (O_782,N_4648,N_4814);
and UO_783 (O_783,N_4908,N_4829);
and UO_784 (O_784,N_4840,N_4863);
or UO_785 (O_785,N_4779,N_4843);
nand UO_786 (O_786,N_4947,N_4730);
nor UO_787 (O_787,N_4674,N_4510);
or UO_788 (O_788,N_4543,N_4896);
and UO_789 (O_789,N_4834,N_4738);
nor UO_790 (O_790,N_4612,N_4532);
or UO_791 (O_791,N_4803,N_4605);
and UO_792 (O_792,N_4737,N_4871);
nor UO_793 (O_793,N_4662,N_4775);
nor UO_794 (O_794,N_4857,N_4787);
nor UO_795 (O_795,N_4880,N_4734);
nand UO_796 (O_796,N_4826,N_4615);
or UO_797 (O_797,N_4698,N_4813);
and UO_798 (O_798,N_4657,N_4805);
or UO_799 (O_799,N_4922,N_4857);
or UO_800 (O_800,N_4648,N_4726);
nand UO_801 (O_801,N_4523,N_4803);
nor UO_802 (O_802,N_4987,N_4710);
and UO_803 (O_803,N_4646,N_4500);
nand UO_804 (O_804,N_4759,N_4533);
xnor UO_805 (O_805,N_4664,N_4709);
or UO_806 (O_806,N_4878,N_4564);
nand UO_807 (O_807,N_4912,N_4620);
and UO_808 (O_808,N_4863,N_4652);
nor UO_809 (O_809,N_4541,N_4629);
nand UO_810 (O_810,N_4648,N_4530);
nand UO_811 (O_811,N_4688,N_4724);
or UO_812 (O_812,N_4789,N_4673);
nor UO_813 (O_813,N_4641,N_4537);
and UO_814 (O_814,N_4637,N_4547);
nor UO_815 (O_815,N_4922,N_4966);
nor UO_816 (O_816,N_4582,N_4664);
and UO_817 (O_817,N_4622,N_4750);
nor UO_818 (O_818,N_4562,N_4922);
xnor UO_819 (O_819,N_4833,N_4996);
xor UO_820 (O_820,N_4715,N_4790);
nor UO_821 (O_821,N_4917,N_4804);
nand UO_822 (O_822,N_4759,N_4872);
or UO_823 (O_823,N_4506,N_4534);
xor UO_824 (O_824,N_4601,N_4912);
nor UO_825 (O_825,N_4965,N_4554);
nor UO_826 (O_826,N_4882,N_4624);
xnor UO_827 (O_827,N_4989,N_4745);
xor UO_828 (O_828,N_4595,N_4760);
nand UO_829 (O_829,N_4701,N_4670);
nand UO_830 (O_830,N_4557,N_4958);
nor UO_831 (O_831,N_4950,N_4665);
nor UO_832 (O_832,N_4868,N_4936);
nor UO_833 (O_833,N_4916,N_4732);
or UO_834 (O_834,N_4741,N_4616);
nor UO_835 (O_835,N_4706,N_4752);
nand UO_836 (O_836,N_4857,N_4807);
nor UO_837 (O_837,N_4560,N_4660);
or UO_838 (O_838,N_4649,N_4541);
xor UO_839 (O_839,N_4701,N_4977);
and UO_840 (O_840,N_4601,N_4916);
and UO_841 (O_841,N_4897,N_4860);
nor UO_842 (O_842,N_4584,N_4593);
nor UO_843 (O_843,N_4941,N_4596);
or UO_844 (O_844,N_4541,N_4622);
and UO_845 (O_845,N_4826,N_4628);
nand UO_846 (O_846,N_4695,N_4996);
nor UO_847 (O_847,N_4853,N_4808);
and UO_848 (O_848,N_4531,N_4935);
and UO_849 (O_849,N_4648,N_4504);
and UO_850 (O_850,N_4678,N_4668);
nor UO_851 (O_851,N_4529,N_4749);
nor UO_852 (O_852,N_4635,N_4510);
nand UO_853 (O_853,N_4722,N_4725);
xnor UO_854 (O_854,N_4512,N_4721);
xnor UO_855 (O_855,N_4907,N_4979);
nor UO_856 (O_856,N_4615,N_4557);
nor UO_857 (O_857,N_4609,N_4732);
and UO_858 (O_858,N_4955,N_4612);
and UO_859 (O_859,N_4960,N_4837);
and UO_860 (O_860,N_4884,N_4898);
nor UO_861 (O_861,N_4921,N_4615);
xor UO_862 (O_862,N_4776,N_4764);
nor UO_863 (O_863,N_4901,N_4553);
nor UO_864 (O_864,N_4745,N_4734);
nand UO_865 (O_865,N_4850,N_4667);
nand UO_866 (O_866,N_4538,N_4949);
nor UO_867 (O_867,N_4570,N_4871);
and UO_868 (O_868,N_4500,N_4519);
or UO_869 (O_869,N_4540,N_4899);
and UO_870 (O_870,N_4594,N_4850);
nand UO_871 (O_871,N_4947,N_4928);
and UO_872 (O_872,N_4889,N_4535);
or UO_873 (O_873,N_4877,N_4698);
nor UO_874 (O_874,N_4984,N_4927);
and UO_875 (O_875,N_4944,N_4834);
nor UO_876 (O_876,N_4698,N_4985);
nor UO_877 (O_877,N_4503,N_4610);
and UO_878 (O_878,N_4973,N_4703);
xor UO_879 (O_879,N_4818,N_4670);
and UO_880 (O_880,N_4899,N_4755);
xnor UO_881 (O_881,N_4867,N_4618);
and UO_882 (O_882,N_4561,N_4835);
xnor UO_883 (O_883,N_4684,N_4860);
nand UO_884 (O_884,N_4616,N_4935);
xor UO_885 (O_885,N_4607,N_4830);
nor UO_886 (O_886,N_4789,N_4735);
and UO_887 (O_887,N_4900,N_4778);
and UO_888 (O_888,N_4734,N_4930);
nor UO_889 (O_889,N_4855,N_4965);
nor UO_890 (O_890,N_4547,N_4703);
or UO_891 (O_891,N_4763,N_4730);
or UO_892 (O_892,N_4952,N_4995);
nand UO_893 (O_893,N_4622,N_4988);
or UO_894 (O_894,N_4683,N_4721);
and UO_895 (O_895,N_4742,N_4892);
or UO_896 (O_896,N_4812,N_4820);
nor UO_897 (O_897,N_4745,N_4642);
and UO_898 (O_898,N_4542,N_4525);
and UO_899 (O_899,N_4905,N_4819);
nand UO_900 (O_900,N_4863,N_4651);
and UO_901 (O_901,N_4657,N_4890);
or UO_902 (O_902,N_4576,N_4851);
nor UO_903 (O_903,N_4524,N_4503);
and UO_904 (O_904,N_4736,N_4921);
or UO_905 (O_905,N_4610,N_4979);
nor UO_906 (O_906,N_4689,N_4542);
or UO_907 (O_907,N_4831,N_4561);
nand UO_908 (O_908,N_4665,N_4536);
or UO_909 (O_909,N_4522,N_4512);
nor UO_910 (O_910,N_4812,N_4551);
or UO_911 (O_911,N_4648,N_4878);
nand UO_912 (O_912,N_4660,N_4652);
nor UO_913 (O_913,N_4965,N_4845);
or UO_914 (O_914,N_4579,N_4979);
nor UO_915 (O_915,N_4764,N_4908);
nand UO_916 (O_916,N_4667,N_4593);
nor UO_917 (O_917,N_4570,N_4696);
nor UO_918 (O_918,N_4650,N_4876);
and UO_919 (O_919,N_4638,N_4678);
nor UO_920 (O_920,N_4854,N_4751);
xnor UO_921 (O_921,N_4899,N_4821);
and UO_922 (O_922,N_4688,N_4592);
and UO_923 (O_923,N_4880,N_4713);
or UO_924 (O_924,N_4971,N_4923);
and UO_925 (O_925,N_4824,N_4781);
or UO_926 (O_926,N_4974,N_4904);
or UO_927 (O_927,N_4577,N_4997);
xnor UO_928 (O_928,N_4667,N_4817);
and UO_929 (O_929,N_4544,N_4708);
or UO_930 (O_930,N_4825,N_4741);
nand UO_931 (O_931,N_4991,N_4746);
nand UO_932 (O_932,N_4672,N_4956);
nor UO_933 (O_933,N_4998,N_4997);
nand UO_934 (O_934,N_4885,N_4987);
nor UO_935 (O_935,N_4741,N_4996);
and UO_936 (O_936,N_4993,N_4788);
nor UO_937 (O_937,N_4645,N_4614);
nor UO_938 (O_938,N_4863,N_4548);
nor UO_939 (O_939,N_4755,N_4860);
nor UO_940 (O_940,N_4931,N_4878);
or UO_941 (O_941,N_4758,N_4697);
and UO_942 (O_942,N_4554,N_4721);
and UO_943 (O_943,N_4776,N_4749);
nand UO_944 (O_944,N_4926,N_4831);
and UO_945 (O_945,N_4679,N_4673);
nor UO_946 (O_946,N_4914,N_4707);
or UO_947 (O_947,N_4705,N_4894);
and UO_948 (O_948,N_4787,N_4575);
and UO_949 (O_949,N_4858,N_4846);
or UO_950 (O_950,N_4867,N_4947);
nand UO_951 (O_951,N_4915,N_4922);
nand UO_952 (O_952,N_4775,N_4543);
and UO_953 (O_953,N_4546,N_4693);
nand UO_954 (O_954,N_4627,N_4516);
or UO_955 (O_955,N_4850,N_4880);
xnor UO_956 (O_956,N_4890,N_4627);
or UO_957 (O_957,N_4798,N_4715);
nor UO_958 (O_958,N_4780,N_4546);
nand UO_959 (O_959,N_4591,N_4860);
nor UO_960 (O_960,N_4874,N_4777);
nor UO_961 (O_961,N_4920,N_4854);
xnor UO_962 (O_962,N_4558,N_4598);
and UO_963 (O_963,N_4663,N_4501);
nor UO_964 (O_964,N_4577,N_4671);
nand UO_965 (O_965,N_4712,N_4910);
nand UO_966 (O_966,N_4655,N_4796);
nor UO_967 (O_967,N_4920,N_4603);
or UO_968 (O_968,N_4645,N_4928);
nand UO_969 (O_969,N_4916,N_4611);
or UO_970 (O_970,N_4993,N_4639);
or UO_971 (O_971,N_4693,N_4530);
nor UO_972 (O_972,N_4729,N_4564);
xor UO_973 (O_973,N_4757,N_4737);
and UO_974 (O_974,N_4989,N_4566);
or UO_975 (O_975,N_4835,N_4910);
xnor UO_976 (O_976,N_4709,N_4799);
or UO_977 (O_977,N_4832,N_4640);
nand UO_978 (O_978,N_4563,N_4507);
nor UO_979 (O_979,N_4669,N_4795);
xnor UO_980 (O_980,N_4797,N_4661);
nor UO_981 (O_981,N_4778,N_4621);
nor UO_982 (O_982,N_4615,N_4974);
or UO_983 (O_983,N_4846,N_4562);
nand UO_984 (O_984,N_4853,N_4643);
nand UO_985 (O_985,N_4686,N_4957);
nor UO_986 (O_986,N_4711,N_4993);
xor UO_987 (O_987,N_4944,N_4545);
xnor UO_988 (O_988,N_4508,N_4553);
or UO_989 (O_989,N_4681,N_4773);
xnor UO_990 (O_990,N_4887,N_4860);
xnor UO_991 (O_991,N_4597,N_4574);
nand UO_992 (O_992,N_4793,N_4636);
or UO_993 (O_993,N_4551,N_4761);
nand UO_994 (O_994,N_4731,N_4734);
nand UO_995 (O_995,N_4953,N_4834);
nor UO_996 (O_996,N_4625,N_4921);
and UO_997 (O_997,N_4858,N_4702);
or UO_998 (O_998,N_4732,N_4825);
nand UO_999 (O_999,N_4782,N_4807);
endmodule