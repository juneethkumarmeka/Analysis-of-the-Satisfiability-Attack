module basic_2000_20000_2500_100_levels_10xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
and U0 (N_0,In_786,In_1965);
or U1 (N_1,In_1473,In_1039);
xnor U2 (N_2,In_1657,In_1648);
and U3 (N_3,In_961,In_1942);
or U4 (N_4,In_822,In_1890);
nor U5 (N_5,In_1667,In_1919);
or U6 (N_6,In_1380,In_773);
and U7 (N_7,In_1376,In_559);
or U8 (N_8,In_1018,In_86);
nor U9 (N_9,In_506,In_1501);
or U10 (N_10,In_289,In_1433);
nor U11 (N_11,In_1579,In_1110);
nor U12 (N_12,In_1256,In_1227);
nand U13 (N_13,In_1016,In_988);
xnor U14 (N_14,In_951,In_327);
and U15 (N_15,In_539,In_425);
nor U16 (N_16,In_180,In_771);
and U17 (N_17,In_1645,In_465);
xnor U18 (N_18,In_384,In_639);
nand U19 (N_19,In_386,In_1064);
nor U20 (N_20,In_693,In_8);
xor U21 (N_21,In_1409,In_1818);
or U22 (N_22,In_362,In_1698);
or U23 (N_23,In_1008,In_1998);
xor U24 (N_24,In_39,In_594);
or U25 (N_25,In_1565,In_497);
and U26 (N_26,In_561,In_183);
xor U27 (N_27,In_906,In_462);
nor U28 (N_28,In_1518,In_1617);
nor U29 (N_29,In_983,In_1742);
and U30 (N_30,In_1369,In_1581);
or U31 (N_31,In_1639,In_1594);
nand U32 (N_32,In_356,In_1595);
xor U33 (N_33,In_1245,In_1613);
nor U34 (N_34,In_1306,In_514);
and U35 (N_35,In_1149,In_167);
and U36 (N_36,In_590,In_1566);
or U37 (N_37,In_211,In_1129);
nand U38 (N_38,In_459,In_485);
xor U39 (N_39,In_511,In_214);
and U40 (N_40,In_549,In_1892);
xor U41 (N_41,In_1701,In_1641);
xor U42 (N_42,In_1211,In_1101);
or U43 (N_43,In_1937,In_944);
or U44 (N_44,In_453,In_1628);
nand U45 (N_45,In_133,In_1930);
and U46 (N_46,In_130,In_1050);
and U47 (N_47,In_1378,In_369);
and U48 (N_48,In_1458,In_24);
and U49 (N_49,In_1560,In_629);
xnor U50 (N_50,In_92,In_1157);
nand U51 (N_51,In_168,In_540);
nor U52 (N_52,In_1277,In_1616);
and U53 (N_53,In_1689,In_1598);
xnor U54 (N_54,In_1644,In_292);
and U55 (N_55,In_127,In_603);
and U56 (N_56,In_472,In_575);
xor U57 (N_57,In_1876,In_1454);
or U58 (N_58,In_816,In_253);
xor U59 (N_59,In_1816,In_41);
and U60 (N_60,In_1672,In_1567);
and U61 (N_61,In_656,In_2);
and U62 (N_62,In_813,In_475);
nor U63 (N_63,In_598,In_448);
nor U64 (N_64,In_1106,In_1585);
and U65 (N_65,In_132,In_288);
xor U66 (N_66,In_1195,In_1307);
nand U67 (N_67,In_1449,In_716);
nor U68 (N_68,In_1186,In_1054);
nor U69 (N_69,In_173,In_1949);
or U70 (N_70,In_874,In_703);
xnor U71 (N_71,In_986,In_814);
nor U72 (N_72,In_1122,In_1231);
and U73 (N_73,In_1649,In_1962);
nor U74 (N_74,In_1671,In_522);
xnor U75 (N_75,In_1751,In_121);
nor U76 (N_76,In_1084,In_1547);
xnor U77 (N_77,In_525,In_1483);
nand U78 (N_78,In_1905,In_873);
nor U79 (N_79,In_1274,In_610);
and U80 (N_80,In_935,In_1024);
nor U81 (N_81,In_95,In_1426);
nand U82 (N_82,In_148,In_1944);
nand U83 (N_83,In_701,In_1213);
nor U84 (N_84,In_815,In_1263);
or U85 (N_85,In_116,In_1575);
or U86 (N_86,In_1334,In_838);
xor U87 (N_87,In_1562,In_1988);
nor U88 (N_88,In_1920,In_1446);
nor U89 (N_89,In_574,In_580);
nand U90 (N_90,In_1093,In_1405);
xnor U91 (N_91,In_219,In_182);
nor U92 (N_92,In_1066,In_910);
xnor U93 (N_93,In_223,In_792);
nand U94 (N_94,In_93,In_1552);
or U95 (N_95,In_64,In_1815);
nand U96 (N_96,In_1356,In_978);
xnor U97 (N_97,In_389,In_1831);
xnor U98 (N_98,In_230,In_1134);
or U99 (N_99,In_1499,In_591);
nand U100 (N_100,In_342,In_619);
or U101 (N_101,In_583,In_479);
xnor U102 (N_102,In_1705,In_1512);
nor U103 (N_103,In_1474,In_1296);
and U104 (N_104,In_232,In_663);
xor U105 (N_105,In_55,In_1844);
nor U106 (N_106,In_611,In_99);
or U107 (N_107,In_1264,In_481);
or U108 (N_108,In_1975,In_1957);
and U109 (N_109,In_404,In_1406);
xnor U110 (N_110,In_1208,In_1187);
nand U111 (N_111,In_1428,In_237);
xor U112 (N_112,In_1312,In_1653);
xor U113 (N_113,In_444,In_992);
nor U114 (N_114,In_565,In_482);
nor U115 (N_115,In_772,In_548);
xnor U116 (N_116,In_105,In_934);
nor U117 (N_117,In_1710,In_1519);
xnor U118 (N_118,In_274,In_1488);
nand U119 (N_119,In_904,In_798);
and U120 (N_120,In_541,In_283);
or U121 (N_121,In_9,In_1556);
or U122 (N_122,In_1337,In_242);
or U123 (N_123,In_1315,In_1335);
nand U124 (N_124,In_1496,In_1941);
xnor U125 (N_125,In_1495,In_1765);
or U126 (N_126,In_1222,In_1693);
nor U127 (N_127,In_1058,In_1860);
xor U128 (N_128,In_783,In_1679);
nand U129 (N_129,In_1000,In_1027);
xnor U130 (N_130,In_504,In_1052);
nand U131 (N_131,In_1838,In_284);
or U132 (N_132,In_1713,In_76);
xnor U133 (N_133,In_353,In_449);
nand U134 (N_134,In_907,In_1036);
xnor U135 (N_135,In_708,In_1708);
and U136 (N_136,In_759,In_333);
or U137 (N_137,In_1292,In_733);
and U138 (N_138,In_602,In_421);
nor U139 (N_139,In_849,In_958);
and U140 (N_140,In_722,In_241);
and U141 (N_141,In_700,In_1752);
xnor U142 (N_142,In_311,In_45);
or U143 (N_143,In_394,In_517);
or U144 (N_144,In_98,In_1120);
xor U145 (N_145,In_1533,In_1207);
or U146 (N_146,In_326,In_868);
nand U147 (N_147,In_1075,In_1850);
nor U148 (N_148,In_1619,In_1758);
or U149 (N_149,In_761,In_1869);
or U150 (N_150,In_831,In_802);
nand U151 (N_151,In_347,In_259);
or U152 (N_152,In_252,In_833);
xor U153 (N_153,In_1456,In_1427);
and U154 (N_154,In_1760,In_1469);
nand U155 (N_155,In_756,In_742);
nand U156 (N_156,In_1275,In_1169);
xnor U157 (N_157,In_923,In_885);
nand U158 (N_158,In_1118,In_942);
and U159 (N_159,In_1784,In_212);
nand U160 (N_160,In_1318,In_1285);
nor U161 (N_161,In_1178,In_4);
xnor U162 (N_162,In_431,In_1785);
and U163 (N_163,In_1529,In_1090);
or U164 (N_164,In_736,In_1342);
or U165 (N_165,In_70,In_764);
xor U166 (N_166,In_763,In_271);
and U167 (N_167,In_89,In_898);
nand U168 (N_168,In_258,In_1424);
or U169 (N_169,In_586,In_1339);
xor U170 (N_170,In_398,In_437);
and U171 (N_171,In_186,In_855);
nand U172 (N_172,In_1221,In_1865);
nor U173 (N_173,In_1125,In_280);
nand U174 (N_174,In_999,In_1593);
xor U175 (N_175,In_850,In_1069);
or U176 (N_176,In_385,In_1548);
and U177 (N_177,In_888,In_1726);
nor U178 (N_178,In_1177,In_1254);
xnor U179 (N_179,In_1435,In_618);
xor U180 (N_180,In_1236,In_1210);
nand U181 (N_181,In_1604,In_1421);
nor U182 (N_182,In_170,In_1922);
nor U183 (N_183,In_1534,In_941);
and U184 (N_184,In_946,In_1523);
and U185 (N_185,In_807,In_175);
nor U186 (N_186,In_1078,In_330);
nor U187 (N_187,In_1206,In_1576);
nor U188 (N_188,In_460,In_758);
nor U189 (N_189,In_501,In_102);
xnor U190 (N_190,In_49,In_1111);
nor U191 (N_191,In_1165,In_1270);
or U192 (N_192,In_631,In_1065);
and U193 (N_193,In_892,In_823);
xnor U194 (N_194,In_528,In_1837);
xor U195 (N_195,In_829,In_227);
xor U196 (N_196,In_1080,In_72);
nor U197 (N_197,In_146,In_301);
or U198 (N_198,In_1384,In_126);
and U199 (N_199,In_1026,In_1741);
and U200 (N_200,In_592,N_14);
nor U201 (N_201,N_48,In_1141);
and U202 (N_202,In_1798,In_1035);
xnor U203 (N_203,In_1669,In_336);
nand U204 (N_204,N_158,In_1845);
nor U205 (N_205,In_799,In_1840);
xnor U206 (N_206,In_77,In_363);
xor U207 (N_207,In_243,In_1123);
and U208 (N_208,In_744,In_1773);
nor U209 (N_209,In_1707,In_3);
or U210 (N_210,In_1067,In_1308);
nor U211 (N_211,In_50,N_73);
xor U212 (N_212,In_1717,In_463);
nor U213 (N_213,In_543,In_1163);
xnor U214 (N_214,N_66,In_1743);
or U215 (N_215,N_35,In_1563);
or U216 (N_216,In_1803,In_775);
xor U217 (N_217,In_1722,In_1961);
xor U218 (N_218,In_1047,In_1685);
and U219 (N_219,In_893,In_1891);
and U220 (N_220,In_1045,In_876);
or U221 (N_221,In_265,In_1128);
nand U222 (N_222,N_37,In_1393);
and U223 (N_223,In_204,In_340);
xnor U224 (N_224,N_45,In_662);
and U225 (N_225,In_1351,In_171);
nor U226 (N_226,In_571,In_524);
xnor U227 (N_227,In_1188,In_1746);
or U228 (N_228,In_1172,In_1592);
or U229 (N_229,In_1135,N_185);
xnor U230 (N_230,In_952,In_249);
xor U231 (N_231,In_1468,In_1544);
and U232 (N_232,In_113,In_103);
nor U233 (N_233,N_31,In_659);
nand U234 (N_234,In_323,In_1882);
nor U235 (N_235,In_1699,In_839);
nor U236 (N_236,In_269,In_595);
nand U237 (N_237,In_1521,In_1060);
xnor U238 (N_238,N_106,In_1926);
and U239 (N_239,N_188,In_865);
and U240 (N_240,In_1774,In_203);
or U241 (N_241,In_791,In_526);
or U242 (N_242,In_1167,In_264);
nand U243 (N_243,In_248,In_494);
or U244 (N_244,In_498,In_1102);
nor U245 (N_245,N_174,In_867);
nand U246 (N_246,In_796,In_1681);
nor U247 (N_247,In_1757,In_1680);
and U248 (N_248,In_1257,In_894);
nor U249 (N_249,In_476,In_136);
nand U250 (N_250,In_1301,In_858);
or U251 (N_251,In_557,In_1244);
or U252 (N_252,In_1300,In_877);
and U253 (N_253,N_163,In_1985);
or U254 (N_254,In_674,In_1739);
xor U255 (N_255,In_657,In_234);
nand U256 (N_256,In_332,In_1085);
nor U257 (N_257,In_1728,N_135);
nand U258 (N_258,In_1358,In_1033);
xor U259 (N_259,In_1323,In_1112);
nand U260 (N_260,In_646,In_1146);
nand U261 (N_261,In_529,In_1507);
and U262 (N_262,In_1663,In_606);
or U263 (N_263,In_1833,In_918);
and U264 (N_264,In_1887,N_61);
xor U265 (N_265,N_76,In_1020);
nor U266 (N_266,In_1745,In_1855);
nor U267 (N_267,In_1725,In_1303);
or U268 (N_268,In_1302,In_1161);
xor U269 (N_269,N_175,In_981);
nand U270 (N_270,In_391,In_185);
xor U271 (N_271,In_331,In_836);
xnor U272 (N_272,In_911,In_1956);
or U273 (N_273,In_26,In_527);
nor U274 (N_274,In_218,N_148);
xnor U275 (N_275,In_600,In_668);
nor U276 (N_276,In_1408,In_1530);
xor U277 (N_277,N_177,In_1);
xnor U278 (N_278,In_312,In_480);
nand U279 (N_279,N_179,In_578);
or U280 (N_280,In_544,In_33);
or U281 (N_281,In_715,In_341);
or U282 (N_282,In_35,In_903);
or U283 (N_283,In_1089,N_117);
nand U284 (N_284,In_1968,In_1935);
xor U285 (N_285,In_140,In_1390);
xor U286 (N_286,In_134,In_1202);
nor U287 (N_287,In_1858,N_72);
or U288 (N_288,In_725,In_81);
nor U289 (N_289,In_381,In_17);
or U290 (N_290,N_87,In_1996);
xor U291 (N_291,In_1772,In_620);
or U292 (N_292,In_846,In_360);
or U293 (N_293,In_1776,In_587);
and U294 (N_294,In_1950,In_1911);
xor U295 (N_295,In_469,In_890);
and U296 (N_296,In_54,In_628);
or U297 (N_297,In_1737,In_487);
xor U298 (N_298,In_1383,In_14);
nand U299 (N_299,In_1082,In_1674);
xnor U300 (N_300,In_627,In_1897);
xnor U301 (N_301,In_652,In_1908);
nand U302 (N_302,In_1602,N_9);
xnor U303 (N_303,In_1476,In_660);
xor U304 (N_304,In_1485,In_392);
or U305 (N_305,In_141,In_905);
nor U306 (N_306,N_90,In_435);
xor U307 (N_307,In_1828,In_1761);
xor U308 (N_308,In_782,In_1889);
or U309 (N_309,In_1500,In_427);
and U310 (N_310,In_1666,In_1637);
and U311 (N_311,In_1901,In_1366);
nand U312 (N_312,N_189,In_68);
nor U313 (N_313,In_1370,In_1907);
xnor U314 (N_314,In_1412,In_29);
and U315 (N_315,In_478,In_1931);
xnor U316 (N_316,In_845,In_1219);
nor U317 (N_317,N_25,In_443);
nand U318 (N_318,In_1711,In_1190);
or U319 (N_319,In_23,In_556);
nand U320 (N_320,In_359,In_1197);
or U321 (N_321,In_1088,In_582);
nand U322 (N_322,In_1997,In_69);
xor U323 (N_323,In_1977,In_1888);
and U324 (N_324,In_1736,In_376);
or U325 (N_325,In_1204,In_834);
nor U326 (N_326,N_39,In_339);
and U327 (N_327,In_1801,In_1540);
and U328 (N_328,N_78,In_1531);
xor U329 (N_329,In_290,N_24);
and U330 (N_330,In_569,In_308);
or U331 (N_331,In_1341,In_1175);
nor U332 (N_332,In_672,In_1096);
nor U333 (N_333,In_1431,In_52);
nand U334 (N_334,In_1253,N_5);
or U335 (N_335,In_1750,In_1879);
nor U336 (N_336,In_509,In_1621);
nand U337 (N_337,In_654,In_1392);
nor U338 (N_338,In_704,In_1640);
and U339 (N_339,In_1948,In_929);
nor U340 (N_340,In_1918,In_950);
nand U341 (N_341,In_1768,In_97);
and U342 (N_342,In_1184,In_388);
nor U343 (N_343,In_357,In_785);
nor U344 (N_344,In_938,In_1492);
and U345 (N_345,In_1484,In_1982);
nand U346 (N_346,In_337,In_1422);
xor U347 (N_347,N_115,N_44);
nor U348 (N_348,In_896,In_1294);
xnor U349 (N_349,In_177,In_348);
and U350 (N_350,In_1417,In_1249);
or U351 (N_351,In_1954,In_20);
xor U352 (N_352,In_1987,In_438);
nor U353 (N_353,N_114,In_1255);
xor U354 (N_354,N_125,In_581);
xnor U355 (N_355,In_1524,In_615);
nor U356 (N_356,In_726,N_102);
nor U357 (N_357,In_593,In_365);
and U358 (N_358,N_132,In_1564);
and U359 (N_359,In_419,In_712);
nor U360 (N_360,N_82,In_1781);
xor U361 (N_361,In_181,In_576);
and U362 (N_362,In_1851,In_972);
or U363 (N_363,In_474,In_1029);
nand U364 (N_364,In_1331,In_1241);
and U365 (N_365,In_1043,In_932);
or U366 (N_366,In_139,In_1841);
or U367 (N_367,In_1720,In_144);
nand U368 (N_368,In_1017,In_636);
or U369 (N_369,In_1748,In_432);
nor U370 (N_370,In_364,In_67);
nor U371 (N_371,In_1659,In_770);
xnor U372 (N_372,In_1976,In_299);
xnor U373 (N_373,N_47,In_864);
nand U374 (N_374,In_1445,In_1360);
nor U375 (N_375,In_1098,In_750);
and U376 (N_376,N_130,N_13);
xnor U377 (N_377,In_1668,In_1945);
and U378 (N_378,In_205,In_1001);
nor U379 (N_379,In_881,In_542);
or U380 (N_380,N_26,In_667);
or U381 (N_381,In_1132,In_1557);
or U382 (N_382,In_1654,In_678);
xor U383 (N_383,In_278,In_1636);
nor U384 (N_384,In_466,In_189);
nand U385 (N_385,In_1200,N_169);
and U386 (N_386,In_1543,In_1522);
xor U387 (N_387,In_426,In_781);
xor U388 (N_388,In_1103,In_12);
and U389 (N_389,In_1283,In_1154);
nand U390 (N_390,In_1854,In_1714);
nor U391 (N_391,In_1138,In_1411);
nand U392 (N_392,In_413,In_1401);
nand U393 (N_393,In_1438,N_41);
nor U394 (N_394,In_1343,In_226);
nand U395 (N_395,In_1517,In_1450);
or U396 (N_396,In_1076,In_268);
and U397 (N_397,In_570,In_1041);
nor U398 (N_398,In_1732,In_367);
nor U399 (N_399,In_1754,N_12);
nand U400 (N_400,In_596,In_56);
or U401 (N_401,N_28,In_768);
or U402 (N_402,In_989,N_86);
and U403 (N_403,In_705,In_1839);
nor U404 (N_404,In_42,In_1655);
nor U405 (N_405,In_695,In_1822);
nand U406 (N_406,N_266,In_519);
or U407 (N_407,In_145,In_1808);
xnor U408 (N_408,In_1046,In_505);
and U409 (N_409,N_176,In_307);
xor U410 (N_410,In_1194,In_1142);
nand U411 (N_411,N_136,N_210);
xnor U412 (N_412,In_1282,In_1170);
xor U413 (N_413,In_1248,In_473);
nand U414 (N_414,N_126,In_1497);
xnor U415 (N_415,In_1787,In_953);
xor U416 (N_416,In_719,In_430);
or U417 (N_417,In_1990,In_34);
and U418 (N_418,N_68,In_1441);
nand U419 (N_419,In_879,N_195);
nor U420 (N_420,N_166,In_974);
xnor U421 (N_421,In_1712,In_1400);
and U422 (N_422,N_162,In_739);
or U423 (N_423,In_1180,In_1056);
nand U424 (N_424,In_975,In_638);
nor U425 (N_425,In_224,In_670);
nand U426 (N_426,In_65,In_1226);
nand U427 (N_427,In_614,In_410);
and U428 (N_428,N_374,N_228);
and U429 (N_429,In_442,N_207);
and U430 (N_430,In_1769,N_157);
or U431 (N_431,In_960,N_33);
nor U432 (N_432,In_706,In_1091);
nor U433 (N_433,In_1261,In_1797);
and U434 (N_434,In_1279,In_675);
or U435 (N_435,In_537,In_378);
or U436 (N_436,In_1738,In_375);
xnor U437 (N_437,In_1506,In_1443);
nand U438 (N_438,In_956,N_342);
nand U439 (N_439,N_324,In_63);
xnor U440 (N_440,In_804,In_1032);
or U441 (N_441,In_1903,In_84);
or U442 (N_442,N_367,In_261);
and U443 (N_443,In_1510,In_401);
and U444 (N_444,In_66,In_1656);
and U445 (N_445,In_320,In_538);
nor U446 (N_446,N_302,In_1823);
nor U447 (N_447,N_196,In_315);
xor U448 (N_448,In_1915,In_1265);
nand U449 (N_449,In_1946,In_379);
and U450 (N_450,In_1218,In_1055);
nor U451 (N_451,In_1721,In_397);
or U452 (N_452,In_461,In_980);
and U453 (N_453,In_115,In_1430);
nand U454 (N_454,In_1127,In_1414);
or U455 (N_455,In_352,In_1320);
nor U456 (N_456,In_1799,In_1086);
xor U457 (N_457,In_402,In_1038);
nor U458 (N_458,In_1196,N_53);
and U459 (N_459,N_85,In_1912);
nor U460 (N_460,In_1324,In_1432);
nand U461 (N_461,In_1896,In_1423);
nor U462 (N_462,In_1028,In_495);
or U463 (N_463,In_1842,In_1804);
or U464 (N_464,N_192,N_242);
nand U465 (N_465,In_1921,N_116);
and U466 (N_466,N_149,In_1970);
nand U467 (N_467,N_160,In_1658);
nor U468 (N_468,In_1993,In_1009);
or U469 (N_469,In_302,N_328);
nand U470 (N_470,In_780,N_361);
or U471 (N_471,N_306,In_564);
nand U472 (N_472,In_1386,In_1419);
or U473 (N_473,In_1861,In_811);
nand U474 (N_474,N_161,In_1189);
or U475 (N_475,In_508,N_10);
nor U476 (N_476,In_921,N_3);
and U477 (N_477,In_129,N_164);
and U478 (N_478,N_291,In_553);
and U479 (N_479,In_734,In_669);
xnor U480 (N_480,In_1661,In_545);
and U481 (N_481,In_899,In_1881);
xnor U482 (N_482,In_1355,In_698);
or U483 (N_483,In_1136,In_954);
nor U484 (N_484,N_32,In_1853);
nor U485 (N_485,In_1247,In_1509);
and U486 (N_486,N_131,N_345);
nand U487 (N_487,In_1153,In_1025);
xor U488 (N_488,In_920,In_1416);
or U489 (N_489,In_1623,In_1706);
and U490 (N_490,In_830,N_255);
and U491 (N_491,In_797,In_1928);
nand U492 (N_492,In_1415,In_745);
nor U493 (N_493,In_808,In_206);
nand U494 (N_494,In_1181,N_287);
nand U495 (N_495,In_1591,In_1755);
nor U496 (N_496,In_753,In_1262);
and U497 (N_497,In_1864,In_691);
or U498 (N_498,In_1352,In_1013);
nor U499 (N_499,N_170,N_49);
xor U500 (N_500,N_171,N_301);
or U501 (N_501,In_731,In_88);
or U502 (N_502,N_215,In_1806);
nor U503 (N_503,In_1151,N_263);
xnor U504 (N_504,N_399,N_91);
and U505 (N_505,N_376,N_198);
and U506 (N_506,In_1240,In_990);
and U507 (N_507,In_1087,In_1703);
nand U508 (N_508,In_821,In_1109);
or U509 (N_509,In_354,In_122);
xor U510 (N_510,In_193,N_191);
nor U511 (N_511,In_380,N_84);
xnor U512 (N_512,N_299,In_677);
nor U513 (N_513,In_687,In_1938);
or U514 (N_514,In_1569,In_1482);
nor U515 (N_515,N_145,N_304);
nand U516 (N_516,In_943,In_322);
nand U517 (N_517,In_1243,In_1162);
or U518 (N_518,In_1271,In_1489);
nor U519 (N_519,In_870,In_1981);
nor U520 (N_520,In_1147,N_225);
or U521 (N_521,In_1470,N_57);
and U522 (N_522,In_959,In_872);
or U523 (N_523,N_359,In_1700);
or U524 (N_524,In_1171,N_235);
or U525 (N_525,N_286,In_192);
nor U526 (N_526,In_572,In_917);
or U527 (N_527,N_150,N_75);
nor U528 (N_528,In_61,In_579);
and U529 (N_529,In_229,In_1192);
nand U530 (N_530,In_1568,In_886);
nor U531 (N_531,In_1871,In_651);
nand U532 (N_532,In_1827,In_1381);
nand U533 (N_533,In_90,N_234);
nor U534 (N_534,N_309,N_284);
nor U535 (N_535,In_1173,In_143);
nor U536 (N_536,In_1642,N_303);
or U537 (N_537,In_689,In_1825);
or U538 (N_538,In_1155,N_38);
or U539 (N_539,N_118,In_535);
nand U540 (N_540,N_382,N_314);
or U541 (N_541,In_351,In_533);
nor U542 (N_542,In_1578,N_379);
nor U543 (N_543,N_54,N_258);
nand U544 (N_544,In_1580,In_1479);
or U545 (N_545,N_83,N_273);
or U546 (N_546,In_1004,In_913);
xor U547 (N_547,N_203,In_987);
and U548 (N_548,In_1126,In_1328);
nand U549 (N_549,N_283,In_550);
and U550 (N_550,In_156,In_1440);
nand U551 (N_551,In_1502,N_393);
nor U552 (N_552,N_298,In_163);
nor U553 (N_553,N_190,In_1460);
nand U554 (N_554,In_765,In_247);
xor U555 (N_555,N_270,N_236);
and U556 (N_556,N_40,N_74);
nand U557 (N_557,In_1549,In_933);
nor U558 (N_558,In_945,In_1662);
nor U559 (N_559,N_46,In_1608);
nand U560 (N_560,In_244,N_140);
and U561 (N_561,In_518,In_1425);
and U562 (N_562,In_1373,In_1230);
nor U563 (N_563,In_1777,In_1800);
nand U564 (N_564,In_546,N_267);
or U565 (N_565,In_147,In_1299);
xnor U566 (N_566,In_31,N_364);
or U567 (N_567,In_680,In_1934);
xor U568 (N_568,In_1756,In_1385);
or U569 (N_569,N_56,In_1332);
and U570 (N_570,N_289,In_1363);
nor U571 (N_571,In_1916,In_1525);
and U572 (N_572,In_995,In_415);
xor U573 (N_573,N_172,N_330);
xnor U574 (N_574,In_150,In_101);
nand U575 (N_575,In_377,In_841);
and U576 (N_576,In_1447,N_219);
or U577 (N_577,In_589,In_832);
and U578 (N_578,N_312,In_1322);
or U579 (N_579,In_914,N_18);
nand U580 (N_580,In_623,In_1986);
nor U581 (N_581,N_292,In_1551);
nand U582 (N_582,N_323,In_1228);
or U583 (N_583,N_383,In_107);
nor U584 (N_584,In_729,In_1541);
nor U585 (N_585,In_106,N_15);
nand U586 (N_586,N_372,In_810);
nand U587 (N_587,In_277,N_340);
nand U588 (N_588,In_767,N_127);
and U589 (N_589,N_260,In_1696);
or U590 (N_590,In_1079,In_1491);
and U591 (N_591,In_231,In_1995);
and U592 (N_592,In_1487,In_344);
nand U593 (N_593,In_1902,In_1104);
or U594 (N_594,In_1830,In_1893);
nand U595 (N_595,In_1665,In_702);
nor U596 (N_596,In_1586,In_1607);
or U597 (N_597,In_1597,In_300);
and U598 (N_598,N_347,In_1462);
nor U599 (N_599,In_1716,In_955);
xor U600 (N_600,In_199,N_461);
nand U601 (N_601,N_381,In_85);
xnor U602 (N_602,In_536,In_1609);
xnor U603 (N_603,In_690,In_458);
and U604 (N_604,N_186,In_441);
nand U605 (N_605,In_1437,In_1297);
and U606 (N_606,In_1478,In_174);
and U607 (N_607,N_512,N_421);
nor U608 (N_608,In_1673,In_1448);
nand U609 (N_609,In_1471,In_194);
and U610 (N_610,In_1690,In_1466);
nor U611 (N_611,In_1843,In_1978);
nor U612 (N_612,In_309,In_1786);
xor U613 (N_613,In_801,In_1824);
and U614 (N_614,In_1849,N_478);
and U615 (N_615,In_1418,In_1936);
xnor U616 (N_616,N_253,N_517);
and U617 (N_617,In_730,N_264);
nor U618 (N_618,In_738,N_209);
nor U619 (N_619,In_285,In_686);
and U620 (N_620,In_1821,N_21);
and U621 (N_621,In_225,In_117);
nand U622 (N_622,In_784,N_88);
or U623 (N_623,In_835,N_506);
nor U624 (N_624,In_1513,In_325);
nor U625 (N_625,N_558,In_1252);
nand U626 (N_626,In_5,N_534);
xor U627 (N_627,In_1251,In_926);
and U628 (N_628,In_1814,N_385);
nor U629 (N_629,In_82,In_643);
nor U630 (N_630,In_1338,In_1344);
xnor U631 (N_631,In_221,In_1735);
or U632 (N_632,N_290,In_109);
or U633 (N_633,In_635,In_803);
and U634 (N_634,In_973,In_114);
xnor U635 (N_635,In_688,In_1702);
xor U636 (N_636,N_487,In_1646);
and U637 (N_637,N_450,N_356);
and U638 (N_638,N_245,In_613);
and U639 (N_639,In_1532,N_36);
xnor U640 (N_640,In_1031,N_281);
or U641 (N_641,In_735,In_1546);
and U642 (N_642,In_1852,In_1397);
and U643 (N_643,In_859,In_1611);
or U644 (N_644,In_1862,N_211);
or U645 (N_645,N_378,In_601);
xnor U646 (N_646,N_146,In_1068);
xnor U647 (N_647,N_265,In_1100);
and U648 (N_648,N_541,In_1638);
xor U649 (N_649,In_400,In_1606);
xnor U650 (N_650,In_967,In_1910);
nand U651 (N_651,In_1237,In_228);
nand U652 (N_652,N_261,In_395);
nand U653 (N_653,In_1766,In_439);
nor U654 (N_654,N_562,In_779);
or U655 (N_655,In_510,N_187);
nor U656 (N_656,In_1073,In_568);
xor U657 (N_657,In_1159,In_977);
or U658 (N_658,In_699,In_848);
or U659 (N_659,In_1615,N_69);
and U660 (N_660,N_110,In_692);
nand U661 (N_661,In_776,N_498);
or U662 (N_662,In_1354,In_707);
nand U663 (N_663,In_740,In_1692);
xnor U664 (N_664,In_94,N_423);
nand U665 (N_665,N_30,N_442);
nor U666 (N_666,In_1394,In_21);
nand U667 (N_667,N_441,In_317);
xor U668 (N_668,N_178,N_555);
nor U669 (N_669,In_1365,In_1234);
xnor U670 (N_670,In_456,N_104);
nand U671 (N_671,In_1472,N_470);
xor U672 (N_672,In_1457,In_1969);
nand U673 (N_673,In_1395,In_1764);
xnor U674 (N_674,In_800,In_632);
and U675 (N_675,In_502,In_1511);
or U676 (N_676,In_1992,In_279);
nand U677 (N_677,In_1232,In_1723);
and U678 (N_678,In_184,In_1310);
nor U679 (N_679,N_220,In_1971);
and U680 (N_680,In_1062,In_566);
and U681 (N_681,N_422,N_592);
nand U682 (N_682,In_447,In_516);
and U683 (N_683,In_153,In_1505);
nor U684 (N_684,N_122,N_269);
nor U685 (N_685,N_221,N_499);
or U686 (N_686,In_1536,N_180);
xor U687 (N_687,In_451,In_1242);
nor U688 (N_688,N_34,In_366);
or U689 (N_689,In_1326,In_343);
or U690 (N_690,N_128,In_1883);
nand U691 (N_691,In_1859,In_75);
and U692 (N_692,N_124,N_504);
and U693 (N_693,In_266,N_463);
xnor U694 (N_694,In_0,In_433);
or U695 (N_695,In_1727,In_11);
nor U696 (N_696,In_53,In_197);
xor U697 (N_697,In_87,N_113);
xor U698 (N_698,In_1724,In_338);
xor U699 (N_699,In_216,In_1734);
xor U700 (N_700,In_276,In_19);
xor U701 (N_701,N_476,In_1398);
or U702 (N_702,In_728,In_996);
xor U703 (N_703,In_1618,In_155);
nor U704 (N_704,In_1413,N_459);
or U705 (N_705,N_17,N_333);
nor U706 (N_706,N_204,N_254);
nand U707 (N_707,In_59,In_976);
or U708 (N_708,In_1329,In_1239);
and U709 (N_709,In_1461,In_1116);
or U710 (N_710,N_556,In_673);
xnor U711 (N_711,N_424,In_1224);
nor U712 (N_712,In_1014,In_142);
and U713 (N_713,N_488,N_508);
nand U714 (N_714,In_74,In_1407);
xnor U715 (N_715,In_1137,N_531);
and U716 (N_716,N_71,N_156);
xor U717 (N_717,In_658,In_968);
xor U718 (N_718,N_248,N_233);
nand U719 (N_719,In_1051,N_391);
nor U720 (N_720,N_509,In_684);
and U721 (N_721,N_193,In_1682);
or U722 (N_722,In_166,In_275);
or U723 (N_723,In_1396,N_355);
xnor U724 (N_724,N_0,In_1856);
nand U725 (N_725,In_1225,In_1201);
or U726 (N_726,N_311,N_325);
nor U727 (N_727,In_28,In_1288);
xnor U728 (N_728,In_751,N_216);
nor U729 (N_729,N_444,In_1537);
and U730 (N_730,In_909,N_447);
nand U731 (N_731,In_245,In_1144);
or U732 (N_732,In_966,N_293);
nor U733 (N_733,In_1526,N_503);
nor U734 (N_734,In_282,N_120);
or U735 (N_735,In_250,In_681);
nor U736 (N_736,In_1095,In_1372);
nor U737 (N_737,N_137,In_417);
nor U738 (N_738,In_188,In_13);
nand U739 (N_739,N_365,N_22);
or U740 (N_740,In_1826,In_1108);
xor U741 (N_741,In_857,In_1289);
and U742 (N_742,In_1220,N_147);
nor U743 (N_743,N_213,In_1626);
or U744 (N_744,In_1939,N_237);
nand U745 (N_745,In_1767,N_481);
and U746 (N_746,In_1715,In_1072);
or U747 (N_747,In_210,In_1573);
and U748 (N_748,In_6,In_1927);
and U749 (N_749,N_535,In_666);
or U750 (N_750,N_65,N_285);
nand U751 (N_751,In_1287,N_262);
nand U752 (N_752,In_162,N_390);
nor U753 (N_753,In_151,In_1924);
nand U754 (N_754,N_59,In_774);
or U755 (N_755,In_254,In_812);
nor U756 (N_756,In_422,N_77);
and U757 (N_757,In_110,In_790);
xor U758 (N_758,In_157,In_1217);
xnor U759 (N_759,N_256,In_853);
nor U760 (N_760,In_1269,In_1233);
xor U761 (N_761,In_1003,N_92);
nor U762 (N_762,N_486,In_450);
nand U763 (N_763,N_16,In_314);
or U764 (N_764,N_565,In_947);
and U765 (N_765,In_160,In_1168);
and U766 (N_766,N_452,In_373);
and U767 (N_767,In_1121,N_419);
nor U768 (N_768,In_1316,In_709);
xnor U769 (N_769,N_346,In_239);
nand U770 (N_770,In_1545,N_571);
nand U771 (N_771,N_344,N_396);
nand U772 (N_772,In_1688,N_231);
and U773 (N_773,In_454,In_1333);
nand U774 (N_774,In_71,N_405);
nor U775 (N_775,In_1780,N_407);
nor U776 (N_776,In_622,In_58);
and U777 (N_777,In_1420,In_1362);
or U778 (N_778,In_1298,In_1559);
or U779 (N_779,In_1904,In_1630);
xor U780 (N_780,In_1092,In_676);
or U781 (N_781,In_260,N_249);
xnor U782 (N_782,In_149,N_2);
or U783 (N_783,In_1744,In_1829);
xor U784 (N_784,N_579,In_1164);
and U785 (N_785,In_1281,In_1464);
or U786 (N_786,In_436,In_1191);
nand U787 (N_787,In_1778,In_1747);
and U788 (N_788,In_1346,In_1260);
nand U789 (N_789,In_1807,In_1465);
nand U790 (N_790,In_423,In_1238);
nor U791 (N_791,N_578,In_1273);
nand U792 (N_792,N_257,N_214);
and U793 (N_793,In_547,N_595);
nand U794 (N_794,N_43,In_1913);
or U795 (N_795,N_143,N_308);
xnor U796 (N_796,N_63,In_1367);
xnor U797 (N_797,N_250,In_1885);
and U798 (N_798,In_1779,N_280);
and U799 (N_799,In_1094,N_477);
and U800 (N_800,In_884,In_491);
xnor U801 (N_801,N_704,N_133);
nand U802 (N_802,In_1515,N_655);
xnor U803 (N_803,In_982,N_404);
or U804 (N_804,N_520,N_19);
xnor U805 (N_805,N_268,N_105);
xor U806 (N_806,N_389,N_511);
xnor U807 (N_807,In_915,In_1955);
nand U808 (N_808,In_817,In_1539);
nand U809 (N_809,In_1214,N_725);
nand U810 (N_810,N_496,N_533);
nor U811 (N_811,N_416,In_316);
nor U812 (N_812,N_208,N_337);
xnor U813 (N_813,In_616,N_403);
nor U814 (N_814,N_698,N_569);
or U815 (N_815,N_676,In_805);
nor U816 (N_816,In_1614,In_1809);
nor U817 (N_817,N_451,N_604);
and U818 (N_818,In_655,N_747);
nor U819 (N_819,N_473,In_1660);
nand U820 (N_820,In_138,N_762);
and U821 (N_821,In_1877,In_1775);
and U822 (N_822,In_47,In_57);
or U823 (N_823,In_1387,In_272);
xor U824 (N_824,In_1790,N_11);
xnor U825 (N_825,In_1368,N_627);
xor U826 (N_826,In_1006,N_358);
and U827 (N_827,In_1650,In_1012);
and U828 (N_828,In_1538,N_720);
nor U829 (N_829,In_863,In_1403);
xor U830 (N_830,In_486,In_445);
or U831 (N_831,In_869,N_142);
nand U832 (N_832,In_27,In_1317);
and U833 (N_833,In_1349,In_372);
xnor U834 (N_834,In_1391,N_384);
nor U835 (N_835,In_1357,In_925);
nor U836 (N_836,In_319,In_641);
nand U837 (N_837,In_235,N_501);
nand U838 (N_838,In_1695,N_686);
nand U839 (N_839,N_723,In_1030);
nand U840 (N_840,In_1268,N_550);
xor U841 (N_841,In_747,N_297);
and U842 (N_842,N_609,In_1622);
nor U843 (N_843,In_43,In_1259);
or U844 (N_844,In_1932,In_1049);
and U845 (N_845,N_537,In_965);
nor U846 (N_846,In_724,In_1436);
xor U847 (N_847,N_350,In_48);
nand U848 (N_848,In_1156,N_707);
nand U849 (N_849,N_538,N_776);
nor U850 (N_850,N_714,N_217);
nand U851 (N_851,N_492,In_573);
nor U852 (N_852,N_483,N_402);
nand U853 (N_853,In_624,In_403);
nand U854 (N_854,In_411,In_1835);
nand U855 (N_855,N_329,In_757);
or U856 (N_856,In_1494,N_480);
nor U857 (N_857,N_647,In_60);
nand U858 (N_858,In_374,N_708);
xor U859 (N_859,In_1675,N_413);
or U860 (N_860,N_710,N_729);
nor U861 (N_861,N_200,In_1097);
or U862 (N_862,N_294,In_1124);
nor U863 (N_863,N_240,In_1964);
or U864 (N_864,In_22,In_754);
xnor U865 (N_865,In_645,In_420);
nand U866 (N_866,In_957,In_1074);
nand U867 (N_867,In_303,N_757);
and U868 (N_868,N_584,N_493);
xnor U869 (N_869,In_406,N_521);
nor U870 (N_870,In_73,In_1878);
nand U871 (N_871,In_588,In_1929);
and U872 (N_872,In_187,N_591);
xor U873 (N_873,N_241,In_1010);
and U874 (N_874,In_295,In_296);
and U875 (N_875,In_871,In_112);
or U876 (N_876,N_760,N_202);
nor U877 (N_877,In_1371,In_1477);
or U878 (N_878,N_432,In_489);
and U879 (N_879,N_693,N_756);
or U880 (N_880,N_697,In_196);
nor U881 (N_881,N_320,In_321);
and U882 (N_882,N_799,In_36);
and U883 (N_883,N_653,In_560);
nor U884 (N_884,In_1951,In_1107);
nand U885 (N_885,In_1295,N_152);
xnor U886 (N_886,N_321,In_1527);
and U887 (N_887,N_731,In_1923);
and U888 (N_888,In_1429,In_824);
and U889 (N_889,In_424,N_665);
nor U890 (N_890,N_67,In_697);
nand U891 (N_891,In_748,N_540);
or U892 (N_892,In_608,N_546);
and U893 (N_893,In_979,In_324);
xnor U894 (N_894,In_457,In_329);
or U895 (N_895,N_637,In_434);
xnor U896 (N_896,N_98,N_386);
nor U897 (N_897,N_439,N_80);
nand U898 (N_898,In_1789,N_679);
or U899 (N_899,In_190,In_1788);
or U900 (N_900,N_251,In_1459);
nor U901 (N_901,In_778,In_1810);
nor U902 (N_902,N_572,In_1811);
and U903 (N_903,N_226,N_599);
nor U904 (N_904,In_1185,N_310);
xnor U905 (N_905,N_519,N_518);
nor U906 (N_906,N_636,N_111);
nand U907 (N_907,N_763,In_1909);
nand U908 (N_908,In_607,N_426);
or U909 (N_909,N_109,N_360);
and U910 (N_910,N_522,N_594);
xor U911 (N_911,N_615,In_350);
nor U912 (N_912,In_297,N_617);
nand U913 (N_913,N_339,In_878);
nand U914 (N_914,N_343,N_564);
nor U915 (N_915,In_642,In_931);
xnor U916 (N_916,N_134,N_554);
nor U917 (N_917,N_792,N_689);
or U918 (N_918,N_181,N_789);
nand U919 (N_919,N_277,In_998);
nor U920 (N_920,In_471,N_787);
nand U921 (N_921,In_46,N_456);
and U922 (N_922,N_612,In_1150);
nor U923 (N_923,N_445,In_523);
xor U924 (N_924,In_1350,N_659);
nand U925 (N_925,In_1463,N_772);
nor U926 (N_926,In_1057,N_749);
xor U927 (N_927,N_387,In_1048);
nor U928 (N_928,In_940,N_692);
xor U929 (N_929,N_773,In_335);
and U930 (N_930,In_262,In_1143);
nand U931 (N_931,N_79,In_1439);
xor U932 (N_932,N_648,In_62);
and U933 (N_933,In_1399,N_100);
nand U934 (N_934,In_198,In_1452);
xor U935 (N_935,In_1105,In_334);
or U936 (N_936,In_963,N_683);
xnor U937 (N_937,In_1709,N_640);
and U938 (N_938,N_717,In_217);
and U939 (N_939,N_427,In_1894);
or U940 (N_940,In_1947,In_1374);
nand U941 (N_941,In_664,N_472);
xnor U942 (N_942,In_1099,N_155);
nand U943 (N_943,N_230,N_119);
nor U944 (N_944,In_1794,In_371);
nor U945 (N_945,In_32,N_716);
nand U946 (N_946,N_502,N_410);
or U947 (N_947,In_1683,N_479);
or U948 (N_948,In_900,N_20);
nor U949 (N_949,In_567,In_1691);
xor U950 (N_950,In_1475,N_611);
and U951 (N_951,In_895,In_554);
and U952 (N_952,In_1933,In_852);
or U953 (N_953,In_1131,In_1015);
xnor U954 (N_954,N_701,N_580);
nor U955 (N_955,N_108,In_1011);
and U956 (N_956,In_318,In_1119);
and U957 (N_957,N_23,In_1943);
xnor U958 (N_958,N_682,In_1596);
nor U959 (N_959,In_685,In_159);
and U960 (N_960,N_103,In_1158);
xnor U961 (N_961,In_1874,In_769);
nor U962 (N_962,In_633,In_222);
xor U963 (N_963,In_428,N_745);
and U964 (N_964,In_154,In_794);
or U965 (N_965,N_334,In_393);
or U966 (N_966,N_351,In_1972);
nor U967 (N_967,N_489,In_346);
or U968 (N_968,In_1037,In_1749);
xnor U969 (N_969,In_563,In_1577);
or U970 (N_970,In_1627,N_530);
nand U971 (N_971,N_566,N_768);
nor U972 (N_972,N_94,N_539);
and U973 (N_973,In_1005,N_64);
xnor U974 (N_974,In_1601,In_455);
nor U975 (N_975,In_1520,In_361);
nand U976 (N_976,In_499,In_875);
or U977 (N_977,N_435,In_1834);
nor U978 (N_978,N_643,N_678);
xnor U979 (N_979,N_151,N_770);
or U980 (N_980,N_660,In_1304);
and U981 (N_981,In_1612,In_1979);
xnor U982 (N_982,N_597,In_1719);
xor U983 (N_983,In_842,In_1782);
or U984 (N_984,N_227,N_524);
xnor U985 (N_985,N_700,In_202);
nand U986 (N_986,N_736,In_1820);
nor U987 (N_987,N_778,In_255);
nand U988 (N_988,In_1966,N_680);
xnor U989 (N_989,In_837,N_505);
or U990 (N_990,In_856,In_984);
or U991 (N_991,In_1313,In_1967);
nand U992 (N_992,In_108,N_796);
xor U993 (N_993,In_530,In_1603);
or U994 (N_994,In_1906,N_625);
xnor U995 (N_995,In_1145,In_1199);
nor U996 (N_996,N_475,In_200);
nor U997 (N_997,N_331,In_605);
or U998 (N_998,N_614,In_383);
and U999 (N_999,In_919,N_494);
and U1000 (N_1000,N_870,In_1872);
or U1001 (N_1001,In_263,N_218);
nor U1002 (N_1002,In_104,In_521);
or U1003 (N_1003,N_397,N_905);
xnor U1004 (N_1004,N_585,N_908);
and U1005 (N_1005,N_603,N_6);
or U1006 (N_1006,N_559,N_840);
and U1007 (N_1007,In_795,N_945);
nor U1008 (N_1008,N_243,In_1077);
nand U1009 (N_1009,N_936,In_1633);
nand U1010 (N_1010,N_785,In_1550);
nor U1011 (N_1011,N_601,In_492);
and U1012 (N_1012,In_119,In_634);
or U1013 (N_1013,N_197,In_165);
nor U1014 (N_1014,N_469,N_774);
and U1015 (N_1015,In_1022,N_780);
or U1016 (N_1016,N_942,In_1071);
nand U1017 (N_1017,In_176,In_1960);
and U1018 (N_1018,In_1353,N_417);
xnor U1019 (N_1019,N_750,N_97);
nand U1020 (N_1020,In_1771,N_529);
nand U1021 (N_1021,In_727,In_446);
and U1022 (N_1022,N_600,N_999);
nor U1023 (N_1023,In_158,In_1635);
and U1024 (N_1024,N_952,N_497);
or U1025 (N_1025,N_980,N_851);
and U1026 (N_1026,N_632,N_437);
nand U1027 (N_1027,In_1115,In_720);
nand U1028 (N_1028,In_1817,N_272);
nor U1029 (N_1029,In_172,In_1994);
nand U1030 (N_1030,In_1857,N_639);
and U1031 (N_1031,N_926,N_663);
nand U1032 (N_1032,N_544,In_1983);
nor U1033 (N_1033,N_836,In_1117);
nand U1034 (N_1034,N_878,In_1561);
nand U1035 (N_1035,In_1677,In_1753);
and U1036 (N_1036,N_588,In_647);
or U1037 (N_1037,N_971,In_1733);
nand U1038 (N_1038,N_829,N_631);
xor U1039 (N_1039,N_975,In_1620);
nand U1040 (N_1040,N_60,In_96);
nor U1041 (N_1041,In_1870,In_936);
nor U1042 (N_1042,N_357,N_165);
and U1043 (N_1043,N_930,In_860);
nand U1044 (N_1044,In_653,N_527);
nor U1045 (N_1045,N_841,N_886);
nor U1046 (N_1046,In_939,N_574);
or U1047 (N_1047,In_51,In_1059);
xnor U1048 (N_1048,In_1686,In_1555);
nand U1049 (N_1049,N_622,In_1867);
and U1050 (N_1050,In_1467,In_1223);
and U1051 (N_1051,In_1250,In_1040);
xnor U1052 (N_1052,In_883,N_199);
and U1053 (N_1053,In_520,N_525);
xor U1054 (N_1054,In_1140,N_702);
or U1055 (N_1055,N_978,N_42);
or U1056 (N_1056,N_784,In_1729);
nor U1057 (N_1057,In_732,In_1174);
xnor U1058 (N_1058,N_96,N_551);
nor U1059 (N_1059,N_121,In_1215);
and U1060 (N_1060,N_671,In_1309);
or U1061 (N_1061,In_882,In_840);
nand U1062 (N_1062,In_100,N_786);
xnor U1063 (N_1063,N_336,In_191);
and U1064 (N_1064,N_932,N_316);
or U1065 (N_1065,In_1974,In_298);
or U1066 (N_1066,N_802,In_125);
nor U1067 (N_1067,N_654,N_994);
xnor U1068 (N_1068,N_436,N_917);
nor U1069 (N_1069,N_581,In_1676);
and U1070 (N_1070,N_318,N_380);
xnor U1071 (N_1071,N_395,In_399);
nand U1072 (N_1072,In_1952,N_645);
nand U1073 (N_1073,N_782,N_244);
nor U1074 (N_1074,N_867,N_872);
xor U1075 (N_1075,In_1813,N_852);
nor U1076 (N_1076,In_551,N_788);
and U1077 (N_1077,In_609,N_744);
nor U1078 (N_1078,In_213,In_818);
or U1079 (N_1079,N_326,N_712);
nor U1080 (N_1080,In_755,N_726);
nor U1081 (N_1081,In_496,In_1516);
nand U1082 (N_1082,In_209,N_677);
nand U1083 (N_1083,N_239,N_904);
nor U1084 (N_1084,N_27,N_915);
or U1085 (N_1085,N_471,N_589);
xnor U1086 (N_1086,In_930,N_608);
nand U1087 (N_1087,N_897,N_818);
xor U1088 (N_1088,N_844,N_93);
nand U1089 (N_1089,In_682,N_935);
nor U1090 (N_1090,N_963,N_278);
nor U1091 (N_1091,In_721,In_577);
xnor U1092 (N_1092,N_860,N_687);
xnor U1093 (N_1093,N_881,In_38);
nor U1094 (N_1094,N_401,In_80);
and U1095 (N_1095,N_846,In_1209);
xor U1096 (N_1096,N_993,N_338);
xor U1097 (N_1097,N_138,N_771);
nand U1098 (N_1098,In_1572,N_934);
and U1099 (N_1099,In_358,In_137);
xnor U1100 (N_1100,N_513,N_721);
nand U1101 (N_1101,N_979,In_927);
and U1102 (N_1102,N_467,N_400);
nor U1103 (N_1103,In_1266,In_880);
and U1104 (N_1104,In_1503,In_1070);
nor U1105 (N_1105,In_819,N_370);
xor U1106 (N_1106,In_1678,N_633);
and U1107 (N_1107,In_737,In_7);
and U1108 (N_1108,In_1498,N_862);
or U1109 (N_1109,N_634,In_1442);
nand U1110 (N_1110,N_734,N_570);
nor U1111 (N_1111,N_953,N_949);
nor U1112 (N_1112,In_1176,N_568);
xnor U1113 (N_1113,N_713,In_710);
nand U1114 (N_1114,In_304,N_918);
nor U1115 (N_1115,In_1160,N_532);
nand U1116 (N_1116,In_928,N_879);
and U1117 (N_1117,N_873,In_1917);
nand U1118 (N_1118,N_798,N_940);
nor U1119 (N_1119,N_247,N_662);
nor U1120 (N_1120,N_101,In_1235);
nand U1121 (N_1121,N_182,In_238);
or U1122 (N_1122,In_273,In_908);
or U1123 (N_1123,In_123,N_913);
or U1124 (N_1124,N_613,N_959);
or U1125 (N_1125,In_949,N_900);
and U1126 (N_1126,In_493,N_751);
nand U1127 (N_1127,N_894,In_1480);
nand U1128 (N_1128,In_1361,In_1589);
nor U1129 (N_1129,In_1989,In_440);
nor U1130 (N_1130,In_1796,In_718);
nor U1131 (N_1131,N_411,In_1866);
or U1132 (N_1132,N_373,N_586);
or U1133 (N_1133,In_1340,N_167);
nand U1134 (N_1134,N_990,In_1034);
and U1135 (N_1135,N_812,N_724);
or U1136 (N_1136,In_287,In_111);
or U1137 (N_1137,N_910,N_684);
nor U1138 (N_1138,N_982,N_661);
xnor U1139 (N_1139,In_679,In_281);
nand U1140 (N_1140,N_649,N_629);
nand U1141 (N_1141,N_740,In_828);
nand U1142 (N_1142,N_415,N_808);
nand U1143 (N_1143,N_877,N_992);
nor U1144 (N_1144,In_640,In_306);
xor U1145 (N_1145,In_1311,N_759);
xnor U1146 (N_1146,N_440,N_327);
nand U1147 (N_1147,In_16,In_310);
xnor U1148 (N_1148,In_169,N_956);
or U1149 (N_1149,N_139,In_604);
xor U1150 (N_1150,N_341,N_408);
nor U1151 (N_1151,N_948,N_922);
nor U1152 (N_1152,In_91,In_1280);
or U1153 (N_1153,N_696,In_1327);
xor U1154 (N_1154,N_646,In_597);
nand U1155 (N_1155,In_889,N_375);
and U1156 (N_1156,In_1278,N_628);
xor U1157 (N_1157,N_767,In_683);
xnor U1158 (N_1158,In_468,N_388);
or U1159 (N_1159,N_839,N_722);
and U1160 (N_1160,In_922,N_866);
nor U1161 (N_1161,N_549,In_788);
and U1162 (N_1162,N_154,N_685);
xnor U1163 (N_1163,In_179,N_859);
xnor U1164 (N_1164,In_1684,In_515);
and U1165 (N_1165,In_1863,In_286);
xor U1166 (N_1166,N_583,In_1819);
or U1167 (N_1167,N_307,In_477);
xor U1168 (N_1168,N_414,N_141);
xor U1169 (N_1169,N_939,N_563);
nand U1170 (N_1170,N_995,N_305);
nor U1171 (N_1171,In_648,In_1246);
xor U1172 (N_1172,N_901,In_843);
xor U1173 (N_1173,In_178,N_651);
xor U1174 (N_1174,In_1434,N_409);
xnor U1175 (N_1175,In_806,N_275);
nand U1176 (N_1176,N_791,N_970);
nand U1177 (N_1177,N_658,In_1325);
and U1178 (N_1178,In_10,In_1330);
xnor U1179 (N_1179,In_752,In_1584);
xor U1180 (N_1180,N_966,N_458);
xor U1181 (N_1181,N_392,In_1021);
or U1182 (N_1182,N_500,N_911);
xor U1183 (N_1183,In_993,N_485);
nand U1184 (N_1184,In_1570,In_1847);
or U1185 (N_1185,N_515,N_857);
xor U1186 (N_1186,In_1697,N_944);
nand U1187 (N_1187,N_536,N_434);
and U1188 (N_1188,In_637,N_727);
or U1189 (N_1189,N_468,In_531);
nand U1190 (N_1190,In_490,In_997);
and U1191 (N_1191,N_354,N_793);
and U1192 (N_1192,N_997,In_626);
or U1193 (N_1193,N_987,In_1179);
or U1194 (N_1194,N_875,In_825);
nand U1195 (N_1195,In_1148,In_1590);
xor U1196 (N_1196,N_474,In_270);
nor U1197 (N_1197,In_1583,N_815);
nor U1198 (N_1198,In_1267,N_753);
xnor U1199 (N_1199,N_616,N_955);
and U1200 (N_1200,N_1018,In_1002);
and U1201 (N_1201,In_1664,N_1182);
and U1202 (N_1202,In_1314,N_349);
nor U1203 (N_1203,In_207,In_1846);
nor U1204 (N_1204,N_547,N_835);
and U1205 (N_1205,In_584,In_1587);
xnor U1206 (N_1206,N_1131,In_1553);
and U1207 (N_1207,N_1105,In_1514);
or U1208 (N_1208,In_1321,N_885);
xor U1209 (N_1209,N_55,N_1007);
or U1210 (N_1210,N_1063,N_1138);
or U1211 (N_1211,In_1730,In_854);
xnor U1212 (N_1212,N_668,N_630);
and U1213 (N_1213,In_368,N_925);
nor U1214 (N_1214,In_44,N_831);
or U1215 (N_1215,N_1100,N_962);
and U1216 (N_1216,N_369,N_1162);
or U1217 (N_1217,N_1025,In_1130);
nor U1218 (N_1218,N_967,N_819);
nand U1219 (N_1219,In_1139,N_732);
xnor U1220 (N_1220,In_711,N_842);
xnor U1221 (N_1221,N_274,N_642);
nor U1222 (N_1222,In_713,In_1802);
nand U1223 (N_1223,N_482,In_532);
nand U1224 (N_1224,In_1868,N_123);
nor U1225 (N_1225,N_797,N_1093);
nand U1226 (N_1226,In_1114,N_1167);
or U1227 (N_1227,In_370,N_650);
or U1228 (N_1228,N_983,N_810);
or U1229 (N_1229,In_1535,N_429);
nor U1230 (N_1230,In_1375,N_398);
or U1231 (N_1231,N_607,N_1153);
xor U1232 (N_1232,N_1082,N_880);
and U1233 (N_1233,N_465,In_1848);
nand U1234 (N_1234,N_1145,N_621);
nand U1235 (N_1235,N_1074,In_1083);
xnor U1236 (N_1236,N_95,In_1805);
xor U1237 (N_1237,N_1142,N_998);
and U1238 (N_1238,In_793,N_898);
nand U1239 (N_1239,N_295,N_667);
and U1240 (N_1240,In_1762,N_1031);
and U1241 (N_1241,N_206,N_624);
xor U1242 (N_1242,In_1599,In_1493);
nand U1243 (N_1243,N_838,N_1134);
and U1244 (N_1244,N_593,N_319);
nand U1245 (N_1245,N_1032,In_827);
xor U1246 (N_1246,In_1899,In_1258);
or U1247 (N_1247,In_1382,In_257);
and U1248 (N_1248,N_1071,N_1112);
and U1249 (N_1249,In_1980,N_865);
nand U1250 (N_1250,N_107,N_931);
nand U1251 (N_1251,N_368,N_845);
and U1252 (N_1252,N_794,N_348);
or U1253 (N_1253,N_112,N_752);
and U1254 (N_1254,In_1759,N_813);
and U1255 (N_1255,N_575,In_777);
nand U1256 (N_1256,N_252,In_1634);
or U1257 (N_1257,In_1528,In_1953);
xnor U1258 (N_1258,In_1588,In_766);
nor U1259 (N_1259,N_1101,In_1212);
nand U1260 (N_1260,N_1010,N_1004);
nor U1261 (N_1261,N_626,N_1065);
nand U1262 (N_1262,N_606,N_363);
nor U1263 (N_1263,In_644,N_528);
and U1264 (N_1264,N_656,N_924);
and U1265 (N_1265,In_1670,N_825);
nor U1266 (N_1266,N_464,N_699);
or U1267 (N_1267,N_1015,N_89);
xnor U1268 (N_1268,In_1914,In_1007);
nand U1269 (N_1269,In_1999,N_371);
and U1270 (N_1270,In_1019,N_1125);
and U1271 (N_1271,N_741,In_507);
and U1272 (N_1272,In_1042,N_446);
nand U1273 (N_1273,N_754,N_882);
nor U1274 (N_1274,N_777,N_484);
nor U1275 (N_1275,N_1069,In_233);
and U1276 (N_1276,N_619,N_279);
xnor U1277 (N_1277,N_1196,N_884);
or U1278 (N_1278,N_1039,In_1651);
and U1279 (N_1279,N_864,N_1121);
xor U1280 (N_1280,In_124,N_1132);
nand U1281 (N_1281,N_223,N_1061);
nor U1282 (N_1282,N_454,In_414);
nor U1283 (N_1283,In_962,N_1023);
nor U1284 (N_1284,N_1011,N_981);
xnor U1285 (N_1285,In_1063,In_83);
or U1286 (N_1286,N_510,N_1012);
and U1287 (N_1287,In_418,In_464);
and U1288 (N_1288,N_394,N_803);
nor U1289 (N_1289,N_352,N_801);
nand U1290 (N_1290,In_37,In_534);
nor U1291 (N_1291,N_1050,N_1186);
and U1292 (N_1292,N_1170,N_828);
nor U1293 (N_1293,N_1174,N_830);
nand U1294 (N_1294,N_1139,N_1161);
xor U1295 (N_1295,N_1128,In_1984);
xor U1296 (N_1296,In_1402,In_862);
nor U1297 (N_1297,N_576,N_1175);
nor U1298 (N_1298,N_1127,In_407);
xor U1299 (N_1299,In_789,In_1836);
nand U1300 (N_1300,In_503,N_1195);
nand U1301 (N_1301,In_1053,N_871);
xnor U1302 (N_1302,N_673,N_928);
xor U1303 (N_1303,N_958,In_1791);
or U1304 (N_1304,In_760,In_1198);
nor U1305 (N_1305,N_1197,N_902);
nand U1306 (N_1306,N_706,In_313);
xnor U1307 (N_1307,N_50,N_814);
nand U1308 (N_1308,N_418,In_897);
nand U1309 (N_1309,In_1410,N_834);
xnor U1310 (N_1310,In_396,In_924);
nor U1311 (N_1311,In_1272,N_205);
nor U1312 (N_1312,In_240,In_743);
nand U1313 (N_1313,N_431,In_40);
nor U1314 (N_1314,N_1144,N_672);
or U1315 (N_1315,In_382,N_300);
nand U1316 (N_1316,N_1154,N_694);
nand U1317 (N_1317,N_212,N_1193);
nor U1318 (N_1318,In_1886,N_1083);
and U1319 (N_1319,N_811,N_1044);
and U1320 (N_1320,N_51,N_703);
nand U1321 (N_1321,In_1631,N_1129);
nor U1322 (N_1322,N_1135,N_874);
nand U1323 (N_1323,In_131,N_965);
or U1324 (N_1324,In_1044,In_994);
nor U1325 (N_1325,N_1077,In_484);
and U1326 (N_1326,In_267,In_128);
nor U1327 (N_1327,In_887,N_709);
nor U1328 (N_1328,N_1086,N_735);
nor U1329 (N_1329,In_1652,N_353);
or U1330 (N_1330,N_406,In_1451);
nor U1331 (N_1331,N_448,In_1453);
or U1332 (N_1332,N_542,N_1160);
nor U1333 (N_1333,In_1455,In_1276);
or U1334 (N_1334,N_1187,N_1098);
nor U1335 (N_1335,In_912,N_822);
nand U1336 (N_1336,N_833,N_737);
or U1337 (N_1337,In_1348,In_1113);
and U1338 (N_1338,N_807,N_858);
and U1339 (N_1339,In_866,In_355);
xnor U1340 (N_1340,N_8,N_184);
or U1341 (N_1341,N_991,In_15);
nand U1342 (N_1342,N_577,N_52);
nor U1343 (N_1343,N_850,N_635);
xor U1344 (N_1344,N_1090,In_294);
xor U1345 (N_1345,N_1066,N_1088);
and U1346 (N_1346,N_769,N_923);
xnor U1347 (N_1347,N_288,N_443);
nand U1348 (N_1348,N_823,N_1055);
nand U1349 (N_1349,N_758,N_229);
nand U1350 (N_1350,In_1574,In_1694);
nand U1351 (N_1351,In_470,N_657);
nand U1352 (N_1352,N_947,N_567);
xor U1353 (N_1353,N_514,N_548);
nor U1354 (N_1354,N_711,In_1632);
nor U1355 (N_1355,In_844,N_1111);
xor U1356 (N_1356,In_1925,N_460);
or U1357 (N_1357,N_688,In_1763);
and U1358 (N_1358,N_764,In_1490);
and U1359 (N_1359,N_1084,N_783);
nand U1360 (N_1360,N_1036,N_1097);
or U1361 (N_1361,N_453,N_669);
and U1362 (N_1362,In_500,N_675);
xnor U1363 (N_1363,N_1028,N_99);
xor U1364 (N_1364,In_120,N_1092);
nor U1365 (N_1365,In_555,N_1166);
nor U1366 (N_1366,In_246,In_1873);
and U1367 (N_1367,N_1177,N_1033);
xor U1368 (N_1368,N_430,N_761);
nand U1369 (N_1369,In_1963,N_1080);
nand U1370 (N_1370,In_1347,N_912);
nand U1371 (N_1371,N_1026,In_1958);
and U1372 (N_1372,N_232,N_1118);
nand U1373 (N_1373,In_1291,In_1182);
or U1374 (N_1374,N_1143,N_929);
nor U1375 (N_1375,In_809,N_1173);
and U1376 (N_1376,N_738,In_1205);
nor U1377 (N_1377,In_1345,N_755);
nand U1378 (N_1378,N_920,N_449);
xor U1379 (N_1379,N_1008,N_889);
nor U1380 (N_1380,N_605,N_1024);
nand U1381 (N_1381,N_1062,N_1059);
or U1382 (N_1382,In_746,In_118);
xor U1383 (N_1383,N_1178,N_1001);
or U1384 (N_1384,In_985,In_630);
nand U1385 (N_1385,In_78,N_746);
nor U1386 (N_1386,N_246,N_1096);
nand U1387 (N_1387,N_1009,In_512);
nor U1388 (N_1388,In_1152,N_1176);
nand U1389 (N_1389,N_420,N_1192);
xor U1390 (N_1390,In_1795,N_1183);
nand U1391 (N_1391,In_1554,N_1137);
or U1392 (N_1392,In_18,N_854);
and U1393 (N_1393,N_1140,In_416);
or U1394 (N_1394,N_674,N_62);
nand U1395 (N_1395,In_937,In_847);
nand U1396 (N_1396,In_1359,N_1188);
or U1397 (N_1397,In_717,In_1875);
nor U1398 (N_1398,N_775,N_590);
and U1399 (N_1399,In_1973,In_483);
xnor U1400 (N_1400,N_1230,N_1171);
or U1401 (N_1401,N_1163,N_1022);
or U1402 (N_1402,N_1208,In_412);
nor U1403 (N_1403,In_599,N_1297);
or U1404 (N_1404,In_1290,In_215);
and U1405 (N_1405,N_1087,N_1391);
or U1406 (N_1406,N_1346,In_1133);
and U1407 (N_1407,N_1122,N_462);
nor U1408 (N_1408,N_1159,N_335);
and U1409 (N_1409,N_1343,N_1099);
xor U1410 (N_1410,N_1308,N_1267);
nand U1411 (N_1411,N_428,N_1310);
or U1412 (N_1412,N_691,In_429);
nor U1413 (N_1413,N_941,N_425);
or U1414 (N_1414,N_1328,In_1404);
or U1415 (N_1415,N_1054,N_1048);
xor U1416 (N_1416,In_1793,In_661);
or U1417 (N_1417,N_1189,In_964);
and U1418 (N_1418,N_1253,In_1542);
xnor U1419 (N_1419,N_1042,In_1704);
xor U1420 (N_1420,N_1234,N_1338);
xnor U1421 (N_1421,N_1248,In_1940);
or U1422 (N_1422,N_4,N_1354);
xor U1423 (N_1423,In_612,In_1605);
nand U1424 (N_1424,N_602,N_781);
or U1425 (N_1425,In_916,N_827);
nor U1426 (N_1426,N_1380,In_152);
or U1427 (N_1427,N_888,N_1051);
or U1428 (N_1428,In_1900,N_1114);
nor U1429 (N_1429,N_1325,N_800);
and U1430 (N_1430,In_513,N_1149);
nor U1431 (N_1431,N_984,N_705);
xnor U1432 (N_1432,In_696,In_714);
or U1433 (N_1433,N_1388,N_1116);
nor U1434 (N_1434,N_1034,N_1276);
nor U1435 (N_1435,N_315,In_1571);
and U1436 (N_1436,In_1629,N_526);
xnor U1437 (N_1437,In_1364,In_201);
or U1438 (N_1438,N_1200,In_1229);
nand U1439 (N_1439,N_81,N_806);
or U1440 (N_1440,N_914,N_933);
xnor U1441 (N_1441,In_552,N_1339);
nand U1442 (N_1442,N_623,N_1365);
nand U1443 (N_1443,In_1379,N_1238);
or U1444 (N_1444,N_1222,N_869);
and U1445 (N_1445,N_194,N_985);
nor U1446 (N_1446,N_644,N_1279);
or U1447 (N_1447,N_1043,N_1266);
nand U1448 (N_1448,N_1382,N_1072);
or U1449 (N_1449,N_891,N_1361);
or U1450 (N_1450,N_1249,N_1298);
or U1451 (N_1451,N_438,N_1307);
nand U1452 (N_1452,N_690,N_695);
xnor U1453 (N_1453,N_1203,N_582);
nand U1454 (N_1454,N_29,N_1259);
and U1455 (N_1455,N_1220,N_1284);
nand U1456 (N_1456,In_650,N_820);
nand U1457 (N_1457,N_1201,In_345);
nand U1458 (N_1458,N_282,In_694);
nor U1459 (N_1459,N_144,N_896);
and U1460 (N_1460,In_1081,N_573);
or U1461 (N_1461,N_1299,N_457);
and U1462 (N_1462,N_989,N_950);
or U1463 (N_1463,N_1347,In_1193);
nor U1464 (N_1464,N_1239,N_1359);
xor U1465 (N_1465,In_723,In_901);
nand U1466 (N_1466,N_322,N_893);
nor U1467 (N_1467,N_824,N_715);
and U1468 (N_1468,N_153,In_328);
nor U1469 (N_1469,N_960,N_1060);
or U1470 (N_1470,N_1181,N_1334);
nand U1471 (N_1471,N_1295,N_1030);
and U1472 (N_1472,N_876,N_1037);
nor U1473 (N_1473,N_1076,N_1379);
xnor U1474 (N_1474,N_1095,N_916);
nand U1475 (N_1475,N_1057,N_1387);
and U1476 (N_1476,N_1165,In_861);
nor U1477 (N_1477,N_1212,N_1274);
or U1478 (N_1478,N_961,N_1273);
and U1479 (N_1479,N_1362,In_1504);
or U1480 (N_1480,N_1345,N_718);
or U1481 (N_1481,N_954,N_1104);
or U1482 (N_1482,N_1290,N_1384);
or U1483 (N_1483,N_1094,N_1064);
xnor U1484 (N_1484,In_948,N_183);
nor U1485 (N_1485,N_1102,N_1324);
nand U1486 (N_1486,N_973,N_466);
xor U1487 (N_1487,N_1243,N_1312);
nand U1488 (N_1488,N_1113,N_1352);
nand U1489 (N_1489,N_868,N_366);
nand U1490 (N_1490,N_1306,In_1898);
xnor U1491 (N_1491,N_1315,N_892);
nand U1492 (N_1492,N_1386,N_1395);
nand U1493 (N_1493,N_1247,N_1383);
and U1494 (N_1494,N_837,In_1610);
or U1495 (N_1495,N_1257,N_1035);
nand U1496 (N_1496,N_1258,N_1357);
nor U1497 (N_1497,N_1255,N_1215);
nand U1498 (N_1498,N_1109,In_1319);
or U1499 (N_1499,N_972,N_1302);
and U1500 (N_1500,In_585,N_1377);
or U1501 (N_1501,In_305,N_1252);
and U1502 (N_1502,N_1002,N_1305);
nand U1503 (N_1503,N_1245,N_1376);
nand U1504 (N_1504,N_332,N_259);
nor U1505 (N_1505,N_1353,N_1021);
and U1506 (N_1506,N_804,In_762);
nand U1507 (N_1507,N_1277,N_909);
or U1508 (N_1508,N_821,N_1340);
nand U1509 (N_1509,N_1190,N_1275);
nand U1510 (N_1510,N_1014,N_1320);
and U1511 (N_1511,In_741,In_208);
nor U1512 (N_1512,N_1336,In_1783);
xor U1513 (N_1513,N_1381,In_1731);
and U1514 (N_1514,N_433,In_558);
nand U1515 (N_1515,N_847,N_1363);
or U1516 (N_1516,N_1265,N_490);
xor U1517 (N_1517,N_1244,In_1305);
xnor U1518 (N_1518,N_1120,In_971);
nor U1519 (N_1519,N_1091,N_742);
and U1520 (N_1520,N_1286,N_1146);
nor U1521 (N_1521,N_1214,N_1313);
or U1522 (N_1522,N_739,N_1106);
xnor U1523 (N_1523,In_1481,N_1269);
xnor U1524 (N_1524,N_743,N_843);
xnor U1525 (N_1525,N_817,N_1108);
and U1526 (N_1526,N_1364,N_1256);
nor U1527 (N_1527,N_1329,N_1003);
or U1528 (N_1528,N_1372,N_557);
xor U1529 (N_1529,In_1832,N_1264);
and U1530 (N_1530,N_1281,N_1356);
nor U1531 (N_1531,N_1235,N_1079);
and U1532 (N_1532,N_652,N_1130);
and U1533 (N_1533,N_1303,N_1236);
xor U1534 (N_1534,N_1289,In_1166);
or U1535 (N_1535,N_1184,In_617);
xor U1536 (N_1536,N_1172,N_1210);
nand U1537 (N_1537,N_1242,N_1263);
and U1538 (N_1538,N_1115,N_362);
xor U1539 (N_1539,In_851,N_1394);
or U1540 (N_1540,In_1718,In_1183);
nor U1541 (N_1541,N_1157,N_1399);
xnor U1542 (N_1542,In_671,N_1219);
and U1543 (N_1543,N_1141,N_1355);
or U1544 (N_1544,N_1202,N_1319);
nand U1545 (N_1545,In_293,N_1204);
xnor U1546 (N_1546,N_1217,In_1388);
and U1547 (N_1547,N_937,N_1211);
nand U1548 (N_1548,N_1278,In_1389);
or U1549 (N_1549,N_596,N_766);
or U1550 (N_1550,In_1625,N_826);
xor U1551 (N_1551,In_405,N_1282);
or U1552 (N_1552,N_1368,N_455);
xor U1553 (N_1553,N_1285,N_1369);
nor U1554 (N_1554,N_317,N_1374);
and U1555 (N_1555,N_968,N_377);
or U1556 (N_1556,N_856,N_1147);
xnor U1557 (N_1557,N_1351,N_795);
and U1558 (N_1558,In_665,N_765);
xnor U1559 (N_1559,N_1006,In_621);
or U1560 (N_1560,N_412,N_1333);
xnor U1561 (N_1561,In_1508,In_161);
or U1562 (N_1562,In_1895,N_1078);
nand U1563 (N_1563,N_1268,N_1393);
nand U1564 (N_1564,N_1209,In_562);
and U1565 (N_1565,N_1119,N_1323);
xor U1566 (N_1566,N_561,In_991);
nand U1567 (N_1567,In_409,N_1389);
nor U1568 (N_1568,N_620,N_1085);
or U1569 (N_1569,N_1013,In_891);
or U1570 (N_1570,N_957,In_349);
or U1571 (N_1571,N_1046,In_625);
xor U1572 (N_1572,N_1073,N_238);
xor U1573 (N_1573,N_587,N_748);
and U1574 (N_1574,N_1103,N_1227);
nand U1575 (N_1575,N_168,N_1291);
xor U1576 (N_1576,In_452,N_1123);
and U1577 (N_1577,N_1251,N_1180);
nor U1578 (N_1578,In_30,N_1360);
xnor U1579 (N_1579,N_1335,N_1194);
and U1580 (N_1580,N_1049,N_1371);
nand U1581 (N_1581,In_1624,N_1246);
nand U1582 (N_1582,N_728,N_976);
and U1583 (N_1583,N_1294,N_1136);
xor U1584 (N_1584,N_1124,N_977);
and U1585 (N_1585,N_552,N_809);
nand U1586 (N_1586,N_1027,N_853);
or U1587 (N_1587,N_805,N_1151);
xor U1588 (N_1588,N_1107,N_1332);
xnor U1589 (N_1589,N_1260,N_890);
xor U1590 (N_1590,In_408,N_543);
and U1591 (N_1591,N_618,In_79);
or U1592 (N_1592,N_1327,In_1687);
nor U1593 (N_1593,N_495,N_1378);
nor U1594 (N_1594,N_1126,N_1225);
xor U1595 (N_1595,In_970,N_1396);
nor U1596 (N_1596,N_1341,N_516);
nand U1597 (N_1597,N_1254,N_1272);
xor U1598 (N_1598,N_1179,N_1000);
xor U1599 (N_1599,In_969,In_387);
nor U1600 (N_1600,N_1206,N_1460);
and U1601 (N_1601,N_1317,N_1436);
nand U1602 (N_1602,N_1300,N_1557);
nor U1603 (N_1603,N_1068,N_1053);
nor U1604 (N_1604,N_1520,N_1591);
xor U1605 (N_1605,N_1191,N_271);
nand U1606 (N_1606,N_681,In_1286);
or U1607 (N_1607,N_1567,N_1479);
nor U1608 (N_1608,N_1579,N_1067);
nor U1609 (N_1609,N_1293,N_1458);
and U1610 (N_1610,N_1005,N_296);
xnor U1611 (N_1611,N_1250,N_1198);
or U1612 (N_1612,N_1530,In_1061);
xor U1613 (N_1613,N_491,N_1510);
xor U1614 (N_1614,N_1471,N_887);
nand U1615 (N_1615,N_1472,N_523);
or U1616 (N_1616,N_1508,N_1562);
xor U1617 (N_1617,N_1434,N_1430);
and U1618 (N_1618,N_1311,N_1487);
nand U1619 (N_1619,N_1330,N_1232);
xor U1620 (N_1620,N_1262,N_964);
and U1621 (N_1621,N_1459,N_1029);
nand U1622 (N_1622,In_1770,N_1490);
or U1623 (N_1623,N_1563,N_666);
nor U1624 (N_1624,N_1438,N_1292);
nand U1625 (N_1625,N_173,N_863);
and U1626 (N_1626,N_1500,N_1370);
nor U1627 (N_1627,N_1481,N_1559);
and U1628 (N_1628,N_1469,N_1449);
or U1629 (N_1629,N_553,N_1358);
nor U1630 (N_1630,In_1284,N_276);
and U1631 (N_1631,N_1423,N_1168);
xor U1632 (N_1632,N_1431,N_1491);
nor U1633 (N_1633,N_1477,N_1419);
nor U1634 (N_1634,N_1405,In_1486);
nor U1635 (N_1635,In_291,N_1566);
nand U1636 (N_1636,N_1526,N_1537);
nor U1637 (N_1637,N_1496,N_1505);
and U1638 (N_1638,N_1553,N_1228);
nand U1639 (N_1639,N_664,N_986);
xnor U1640 (N_1640,N_1594,N_1538);
and U1641 (N_1641,N_895,N_1373);
xor U1642 (N_1642,In_1792,N_1081);
nand U1643 (N_1643,N_1482,N_1400);
and U1644 (N_1644,N_1271,N_1571);
nand U1645 (N_1645,N_883,N_222);
and U1646 (N_1646,N_719,N_1385);
nand U1647 (N_1647,N_1462,N_1350);
nand U1648 (N_1648,In_1203,N_1455);
and U1649 (N_1649,N_1463,N_1413);
and U1650 (N_1650,N_951,In_1812);
nor U1651 (N_1651,N_849,N_1052);
nand U1652 (N_1652,N_1038,N_855);
and U1653 (N_1653,N_1390,N_1418);
and U1654 (N_1654,In_135,N_670);
and U1655 (N_1655,N_1420,N_1150);
and U1656 (N_1656,N_1493,N_1040);
xnor U1657 (N_1657,N_1546,N_1583);
or U1658 (N_1658,N_1593,N_1509);
xor U1659 (N_1659,N_1507,N_1445);
or U1660 (N_1660,N_1580,N_969);
xnor U1661 (N_1661,N_1574,N_1539);
nor U1662 (N_1662,N_1429,N_1270);
xnor U1663 (N_1663,N_1047,N_641);
and U1664 (N_1664,N_1322,N_1519);
xnor U1665 (N_1665,In_220,N_1);
nand U1666 (N_1666,In_251,N_1589);
and U1667 (N_1667,N_1494,N_974);
xor U1668 (N_1668,N_1296,N_1522);
or U1669 (N_1669,N_638,N_1527);
and U1670 (N_1670,In_1991,N_1446);
or U1671 (N_1671,N_1576,N_1598);
and U1672 (N_1672,N_1218,N_1544);
nor U1673 (N_1673,N_1221,N_1529);
or U1674 (N_1674,N_1375,N_1440);
nand U1675 (N_1675,N_730,N_1416);
or U1676 (N_1676,N_1473,In_1740);
or U1677 (N_1677,N_919,N_903);
xor U1678 (N_1678,N_1318,N_1058);
and U1679 (N_1679,N_1587,In_25);
and U1680 (N_1680,N_1521,N_1283);
xor U1681 (N_1681,N_1542,N_1524);
nor U1682 (N_1682,N_1569,N_201);
and U1683 (N_1683,N_848,N_1397);
and U1684 (N_1684,N_1582,N_1229);
nand U1685 (N_1685,N_816,N_1443);
and U1686 (N_1686,N_927,N_1503);
xnor U1687 (N_1687,In_390,In_164);
and U1688 (N_1688,N_1550,N_1045);
xnor U1689 (N_1689,N_1422,N_1117);
nor U1690 (N_1690,N_1499,N_1326);
nor U1691 (N_1691,N_1417,N_1536);
or U1692 (N_1692,N_1424,N_1543);
and U1693 (N_1693,N_1485,N_1241);
and U1694 (N_1694,N_1474,N_1467);
nor U1695 (N_1695,N_1599,N_1156);
nand U1696 (N_1696,N_1515,N_1342);
xnor U1697 (N_1697,N_1216,N_1586);
xor U1698 (N_1698,In_820,N_7);
nand U1699 (N_1699,N_906,N_1528);
nor U1700 (N_1700,N_1280,N_1556);
or U1701 (N_1701,N_70,N_1185);
nand U1702 (N_1702,N_1534,N_1089);
and U1703 (N_1703,In_1880,N_1207);
or U1704 (N_1704,N_1056,N_1456);
or U1705 (N_1705,N_1584,N_1497);
and U1706 (N_1706,N_129,In_1293);
nor U1707 (N_1707,N_1017,N_159);
or U1708 (N_1708,N_1560,N_1457);
xnor U1709 (N_1709,N_1435,N_1448);
and U1710 (N_1710,N_907,N_1442);
xnor U1711 (N_1711,N_1401,N_1316);
nand U1712 (N_1712,N_1461,N_1410);
nand U1713 (N_1713,N_1502,N_1041);
nor U1714 (N_1714,N_1439,N_1402);
nand U1715 (N_1715,N_1411,N_1428);
xnor U1716 (N_1716,N_1523,N_1596);
or U1717 (N_1717,N_1578,In_256);
and U1718 (N_1718,N_1452,N_779);
and U1719 (N_1719,N_1555,N_598);
nand U1720 (N_1720,N_1331,N_1447);
xnor U1721 (N_1721,N_1213,N_943);
or U1722 (N_1722,N_1427,In_1023);
and U1723 (N_1723,N_1558,In_649);
or U1724 (N_1724,N_1495,In_1444);
nand U1725 (N_1725,In_1647,N_1415);
nor U1726 (N_1726,N_1464,N_1392);
xnor U1727 (N_1727,N_1349,N_1531);
nand U1728 (N_1728,N_1404,N_1309);
xor U1729 (N_1729,N_1148,N_1561);
nor U1730 (N_1730,N_1240,N_1288);
nor U1731 (N_1731,N_1367,In_236);
or U1732 (N_1732,N_1199,N_1426);
nor U1733 (N_1733,N_1409,N_1226);
xnor U1734 (N_1734,N_1532,N_1070);
or U1735 (N_1735,N_1585,In_787);
nand U1736 (N_1736,N_1506,N_1570);
nor U1737 (N_1737,N_1019,N_224);
or U1738 (N_1738,N_1552,N_1425);
or U1739 (N_1739,N_1450,N_1551);
nand U1740 (N_1740,N_1533,N_1516);
xnor U1741 (N_1741,N_1565,N_610);
xor U1742 (N_1742,N_1169,N_1483);
xnor U1743 (N_1743,N_1398,N_1421);
nor U1744 (N_1744,In_467,N_1261);
and U1745 (N_1745,N_733,N_938);
or U1746 (N_1746,N_1437,N_1133);
nand U1747 (N_1747,N_1453,N_1408);
nand U1748 (N_1748,N_1441,N_1540);
nor U1749 (N_1749,In_749,N_1573);
nand U1750 (N_1750,N_1233,N_507);
nor U1751 (N_1751,In_902,N_1020);
xnor U1752 (N_1752,N_1488,N_1545);
or U1753 (N_1753,N_1468,N_545);
nand U1754 (N_1754,N_1492,N_1433);
xor U1755 (N_1755,In_1336,N_1231);
or U1756 (N_1756,N_1476,N_899);
nor U1757 (N_1757,N_1432,N_1541);
nand U1758 (N_1758,N_996,N_1514);
xor U1759 (N_1759,N_1155,N_1016);
and U1760 (N_1760,N_1554,In_488);
and U1761 (N_1761,N_1512,N_1152);
nor U1762 (N_1762,N_1465,N_861);
nor U1763 (N_1763,N_1592,In_826);
xor U1764 (N_1764,N_1517,N_1321);
xnor U1765 (N_1765,N_1581,N_1470);
xor U1766 (N_1766,In_1377,N_313);
xnor U1767 (N_1767,In_1643,N_1224);
nor U1768 (N_1768,N_1454,N_1475);
nor U1769 (N_1769,N_1489,N_1525);
and U1770 (N_1770,N_1504,N_1511);
or U1771 (N_1771,N_1301,N_1480);
nor U1772 (N_1772,N_1498,N_1590);
or U1773 (N_1773,N_1304,N_1366);
nand U1774 (N_1774,N_1549,N_1572);
nor U1775 (N_1775,N_1597,In_1216);
nor U1776 (N_1776,N_1535,N_1444);
nor U1777 (N_1777,N_1337,N_1414);
xor U1778 (N_1778,N_1158,N_1595);
or U1779 (N_1779,N_1564,N_1223);
and U1780 (N_1780,N_988,N_1164);
nand U1781 (N_1781,N_1478,N_790);
nand U1782 (N_1782,N_1484,N_1577);
and U1783 (N_1783,N_1451,N_921);
xor U1784 (N_1784,N_1407,N_1348);
nor U1785 (N_1785,N_1344,In_1582);
nand U1786 (N_1786,N_946,N_1314);
nor U1787 (N_1787,N_1588,N_1513);
or U1788 (N_1788,In_195,N_1412);
nand U1789 (N_1789,In_1959,In_1558);
xor U1790 (N_1790,N_1568,N_832);
and U1791 (N_1791,N_1406,N_1205);
and U1792 (N_1792,N_1075,N_58);
and U1793 (N_1793,N_1486,N_1518);
nor U1794 (N_1794,N_1403,N_560);
nor U1795 (N_1795,N_1575,In_1884);
and U1796 (N_1796,N_1547,N_1287);
and U1797 (N_1797,N_1237,In_1600);
and U1798 (N_1798,N_1110,N_1466);
or U1799 (N_1799,N_1501,N_1548);
nor U1800 (N_1800,N_1705,N_1794);
xor U1801 (N_1801,N_1735,N_1725);
xor U1802 (N_1802,N_1609,N_1798);
and U1803 (N_1803,N_1619,N_1729);
xor U1804 (N_1804,N_1620,N_1699);
nor U1805 (N_1805,N_1644,N_1704);
and U1806 (N_1806,N_1642,N_1790);
nor U1807 (N_1807,N_1695,N_1721);
or U1808 (N_1808,N_1763,N_1693);
and U1809 (N_1809,N_1740,N_1753);
and U1810 (N_1810,N_1706,N_1750);
nand U1811 (N_1811,N_1643,N_1679);
nor U1812 (N_1812,N_1650,N_1688);
nand U1813 (N_1813,N_1603,N_1662);
or U1814 (N_1814,N_1666,N_1700);
or U1815 (N_1815,N_1655,N_1645);
and U1816 (N_1816,N_1764,N_1604);
or U1817 (N_1817,N_1629,N_1680);
or U1818 (N_1818,N_1727,N_1605);
nand U1819 (N_1819,N_1624,N_1758);
nand U1820 (N_1820,N_1634,N_1775);
nand U1821 (N_1821,N_1777,N_1617);
and U1822 (N_1822,N_1779,N_1610);
and U1823 (N_1823,N_1787,N_1616);
or U1824 (N_1824,N_1697,N_1630);
nand U1825 (N_1825,N_1756,N_1742);
nor U1826 (N_1826,N_1755,N_1622);
or U1827 (N_1827,N_1627,N_1783);
and U1828 (N_1828,N_1771,N_1701);
xor U1829 (N_1829,N_1677,N_1743);
and U1830 (N_1830,N_1639,N_1684);
nand U1831 (N_1831,N_1657,N_1703);
nand U1832 (N_1832,N_1631,N_1691);
nor U1833 (N_1833,N_1646,N_1690);
or U1834 (N_1834,N_1719,N_1683);
xnor U1835 (N_1835,N_1731,N_1702);
or U1836 (N_1836,N_1770,N_1614);
and U1837 (N_1837,N_1602,N_1670);
or U1838 (N_1838,N_1738,N_1789);
nor U1839 (N_1839,N_1728,N_1785);
nand U1840 (N_1840,N_1611,N_1766);
and U1841 (N_1841,N_1724,N_1791);
nor U1842 (N_1842,N_1749,N_1776);
or U1843 (N_1843,N_1754,N_1720);
and U1844 (N_1844,N_1685,N_1759);
nor U1845 (N_1845,N_1711,N_1661);
xnor U1846 (N_1846,N_1793,N_1768);
nor U1847 (N_1847,N_1621,N_1713);
xor U1848 (N_1848,N_1694,N_1736);
or U1849 (N_1849,N_1668,N_1686);
xnor U1850 (N_1850,N_1656,N_1632);
xnor U1851 (N_1851,N_1784,N_1612);
or U1852 (N_1852,N_1652,N_1671);
nor U1853 (N_1853,N_1774,N_1796);
or U1854 (N_1854,N_1633,N_1601);
nor U1855 (N_1855,N_1653,N_1730);
nor U1856 (N_1856,N_1696,N_1752);
xor U1857 (N_1857,N_1741,N_1773);
and U1858 (N_1858,N_1760,N_1682);
and U1859 (N_1859,N_1649,N_1765);
xor U1860 (N_1860,N_1757,N_1663);
xnor U1861 (N_1861,N_1648,N_1709);
nand U1862 (N_1862,N_1669,N_1626);
nor U1863 (N_1863,N_1778,N_1712);
nand U1864 (N_1864,N_1636,N_1795);
xor U1865 (N_1865,N_1715,N_1692);
nor U1866 (N_1866,N_1651,N_1744);
and U1867 (N_1867,N_1673,N_1608);
nand U1868 (N_1868,N_1647,N_1746);
or U1869 (N_1869,N_1618,N_1665);
xor U1870 (N_1870,N_1623,N_1678);
xor U1871 (N_1871,N_1607,N_1710);
nand U1872 (N_1872,N_1726,N_1637);
nand U1873 (N_1873,N_1732,N_1769);
nand U1874 (N_1874,N_1659,N_1792);
and U1875 (N_1875,N_1734,N_1717);
nand U1876 (N_1876,N_1747,N_1733);
nor U1877 (N_1877,N_1672,N_1664);
or U1878 (N_1878,N_1707,N_1788);
and U1879 (N_1879,N_1606,N_1786);
nor U1880 (N_1880,N_1638,N_1772);
xnor U1881 (N_1881,N_1737,N_1675);
nand U1882 (N_1882,N_1654,N_1780);
or U1883 (N_1883,N_1782,N_1723);
xnor U1884 (N_1884,N_1722,N_1640);
nor U1885 (N_1885,N_1745,N_1613);
nor U1886 (N_1886,N_1667,N_1716);
or U1887 (N_1887,N_1698,N_1751);
nand U1888 (N_1888,N_1674,N_1600);
and U1889 (N_1889,N_1689,N_1628);
and U1890 (N_1890,N_1714,N_1708);
nor U1891 (N_1891,N_1718,N_1676);
nor U1892 (N_1892,N_1739,N_1761);
or U1893 (N_1893,N_1658,N_1748);
or U1894 (N_1894,N_1799,N_1797);
and U1895 (N_1895,N_1625,N_1687);
or U1896 (N_1896,N_1762,N_1681);
nand U1897 (N_1897,N_1660,N_1635);
and U1898 (N_1898,N_1641,N_1781);
nand U1899 (N_1899,N_1615,N_1767);
nor U1900 (N_1900,N_1747,N_1721);
or U1901 (N_1901,N_1721,N_1644);
nor U1902 (N_1902,N_1720,N_1722);
nand U1903 (N_1903,N_1677,N_1780);
nand U1904 (N_1904,N_1721,N_1798);
xnor U1905 (N_1905,N_1731,N_1742);
and U1906 (N_1906,N_1744,N_1647);
nand U1907 (N_1907,N_1671,N_1686);
nand U1908 (N_1908,N_1700,N_1613);
or U1909 (N_1909,N_1749,N_1623);
and U1910 (N_1910,N_1784,N_1769);
xnor U1911 (N_1911,N_1666,N_1797);
nand U1912 (N_1912,N_1622,N_1644);
nand U1913 (N_1913,N_1697,N_1664);
or U1914 (N_1914,N_1758,N_1660);
and U1915 (N_1915,N_1667,N_1622);
nand U1916 (N_1916,N_1708,N_1777);
xor U1917 (N_1917,N_1787,N_1711);
and U1918 (N_1918,N_1769,N_1692);
nand U1919 (N_1919,N_1649,N_1729);
or U1920 (N_1920,N_1748,N_1619);
xnor U1921 (N_1921,N_1617,N_1785);
nand U1922 (N_1922,N_1784,N_1602);
nand U1923 (N_1923,N_1659,N_1679);
or U1924 (N_1924,N_1744,N_1687);
nand U1925 (N_1925,N_1749,N_1613);
nor U1926 (N_1926,N_1737,N_1794);
nor U1927 (N_1927,N_1615,N_1635);
and U1928 (N_1928,N_1636,N_1700);
and U1929 (N_1929,N_1735,N_1629);
and U1930 (N_1930,N_1772,N_1618);
nor U1931 (N_1931,N_1638,N_1654);
or U1932 (N_1932,N_1711,N_1775);
and U1933 (N_1933,N_1764,N_1778);
and U1934 (N_1934,N_1790,N_1653);
nor U1935 (N_1935,N_1703,N_1737);
nor U1936 (N_1936,N_1654,N_1757);
xor U1937 (N_1937,N_1601,N_1793);
nor U1938 (N_1938,N_1728,N_1709);
xor U1939 (N_1939,N_1708,N_1745);
nand U1940 (N_1940,N_1721,N_1716);
nor U1941 (N_1941,N_1788,N_1748);
and U1942 (N_1942,N_1655,N_1717);
or U1943 (N_1943,N_1628,N_1608);
nor U1944 (N_1944,N_1779,N_1642);
nor U1945 (N_1945,N_1606,N_1630);
xnor U1946 (N_1946,N_1681,N_1792);
and U1947 (N_1947,N_1787,N_1761);
nor U1948 (N_1948,N_1767,N_1606);
or U1949 (N_1949,N_1670,N_1600);
nand U1950 (N_1950,N_1643,N_1714);
nor U1951 (N_1951,N_1754,N_1742);
and U1952 (N_1952,N_1781,N_1758);
and U1953 (N_1953,N_1736,N_1690);
or U1954 (N_1954,N_1607,N_1756);
or U1955 (N_1955,N_1739,N_1754);
nand U1956 (N_1956,N_1732,N_1645);
xnor U1957 (N_1957,N_1744,N_1730);
nor U1958 (N_1958,N_1738,N_1703);
and U1959 (N_1959,N_1625,N_1727);
xor U1960 (N_1960,N_1770,N_1729);
and U1961 (N_1961,N_1725,N_1660);
and U1962 (N_1962,N_1631,N_1746);
and U1963 (N_1963,N_1683,N_1712);
and U1964 (N_1964,N_1636,N_1634);
xor U1965 (N_1965,N_1665,N_1617);
xor U1966 (N_1966,N_1614,N_1764);
xor U1967 (N_1967,N_1731,N_1666);
nor U1968 (N_1968,N_1740,N_1646);
xnor U1969 (N_1969,N_1763,N_1796);
and U1970 (N_1970,N_1745,N_1698);
nand U1971 (N_1971,N_1657,N_1693);
or U1972 (N_1972,N_1753,N_1713);
nand U1973 (N_1973,N_1748,N_1746);
xor U1974 (N_1974,N_1759,N_1692);
xnor U1975 (N_1975,N_1676,N_1607);
nand U1976 (N_1976,N_1601,N_1752);
nand U1977 (N_1977,N_1642,N_1686);
and U1978 (N_1978,N_1658,N_1791);
or U1979 (N_1979,N_1688,N_1682);
nand U1980 (N_1980,N_1715,N_1650);
or U1981 (N_1981,N_1796,N_1719);
nand U1982 (N_1982,N_1683,N_1639);
xnor U1983 (N_1983,N_1685,N_1787);
nor U1984 (N_1984,N_1679,N_1683);
nand U1985 (N_1985,N_1617,N_1659);
or U1986 (N_1986,N_1621,N_1796);
xor U1987 (N_1987,N_1661,N_1762);
or U1988 (N_1988,N_1625,N_1660);
xor U1989 (N_1989,N_1770,N_1784);
nand U1990 (N_1990,N_1679,N_1784);
xor U1991 (N_1991,N_1786,N_1793);
and U1992 (N_1992,N_1602,N_1758);
nand U1993 (N_1993,N_1680,N_1755);
nor U1994 (N_1994,N_1614,N_1799);
and U1995 (N_1995,N_1753,N_1799);
or U1996 (N_1996,N_1683,N_1695);
or U1997 (N_1997,N_1707,N_1683);
or U1998 (N_1998,N_1692,N_1707);
nand U1999 (N_1999,N_1753,N_1791);
nor U2000 (N_2000,N_1924,N_1818);
nor U2001 (N_2001,N_1954,N_1899);
and U2002 (N_2002,N_1946,N_1896);
xnor U2003 (N_2003,N_1881,N_1996);
or U2004 (N_2004,N_1992,N_1801);
nand U2005 (N_2005,N_1839,N_1858);
or U2006 (N_2006,N_1847,N_1861);
nand U2007 (N_2007,N_1860,N_1935);
or U2008 (N_2008,N_1925,N_1884);
and U2009 (N_2009,N_1857,N_1914);
xnor U2010 (N_2010,N_1800,N_1822);
or U2011 (N_2011,N_1849,N_1909);
nor U2012 (N_2012,N_1886,N_1859);
or U2013 (N_2013,N_1998,N_1983);
nor U2014 (N_2014,N_1916,N_1869);
and U2015 (N_2015,N_1918,N_1961);
nand U2016 (N_2016,N_1811,N_1936);
xnor U2017 (N_2017,N_1862,N_1844);
nand U2018 (N_2018,N_1979,N_1919);
and U2019 (N_2019,N_1870,N_1855);
nor U2020 (N_2020,N_1879,N_1873);
xor U2021 (N_2021,N_1823,N_1981);
nand U2022 (N_2022,N_1955,N_1966);
and U2023 (N_2023,N_1820,N_1923);
xnor U2024 (N_2024,N_1989,N_1851);
xor U2025 (N_2025,N_1980,N_1848);
xor U2026 (N_2026,N_1910,N_1827);
nand U2027 (N_2027,N_1997,N_1937);
and U2028 (N_2028,N_1872,N_1817);
nor U2029 (N_2029,N_1863,N_1991);
xor U2030 (N_2030,N_1803,N_1890);
nor U2031 (N_2031,N_1977,N_1978);
or U2032 (N_2032,N_1846,N_1807);
nand U2033 (N_2033,N_1947,N_1972);
or U2034 (N_2034,N_1994,N_1830);
and U2035 (N_2035,N_1878,N_1831);
or U2036 (N_2036,N_1968,N_1920);
or U2037 (N_2037,N_1926,N_1821);
nand U2038 (N_2038,N_1973,N_1949);
or U2039 (N_2039,N_1845,N_1964);
xor U2040 (N_2040,N_1952,N_1889);
or U2041 (N_2041,N_1934,N_1959);
or U2042 (N_2042,N_1814,N_1834);
nor U2043 (N_2043,N_1852,N_1905);
xnor U2044 (N_2044,N_1948,N_1908);
or U2045 (N_2045,N_1856,N_1880);
nand U2046 (N_2046,N_1885,N_1900);
xor U2047 (N_2047,N_1810,N_1813);
or U2048 (N_2048,N_1999,N_1853);
xnor U2049 (N_2049,N_1805,N_1854);
nand U2050 (N_2050,N_1988,N_1957);
nand U2051 (N_2051,N_1819,N_1891);
xor U2052 (N_2052,N_1887,N_1895);
nand U2053 (N_2053,N_1868,N_1917);
nor U2054 (N_2054,N_1944,N_1963);
or U2055 (N_2055,N_1876,N_1816);
nand U2056 (N_2056,N_1812,N_1833);
nand U2057 (N_2057,N_1930,N_1836);
or U2058 (N_2058,N_1867,N_1967);
or U2059 (N_2059,N_1929,N_1832);
and U2060 (N_2060,N_1874,N_1808);
and U2061 (N_2061,N_1938,N_1829);
nor U2062 (N_2062,N_1941,N_1942);
nor U2063 (N_2063,N_1971,N_1984);
xnor U2064 (N_2064,N_1921,N_1943);
nor U2065 (N_2065,N_1866,N_1898);
nand U2066 (N_2066,N_1939,N_1990);
nand U2067 (N_2067,N_1932,N_1907);
nand U2068 (N_2068,N_1877,N_1986);
nand U2069 (N_2069,N_1806,N_1825);
or U2070 (N_2070,N_1815,N_1842);
or U2071 (N_2071,N_1915,N_1865);
nand U2072 (N_2072,N_1912,N_1951);
or U2073 (N_2073,N_1882,N_1843);
nand U2074 (N_2074,N_1945,N_1970);
xor U2075 (N_2075,N_1883,N_1888);
nand U2076 (N_2076,N_1974,N_1987);
nor U2077 (N_2077,N_1871,N_1841);
nand U2078 (N_2078,N_1904,N_1906);
xnor U2079 (N_2079,N_1953,N_1837);
or U2080 (N_2080,N_1824,N_1903);
and U2081 (N_2081,N_1928,N_1982);
and U2082 (N_2082,N_1913,N_1927);
xor U2083 (N_2083,N_1940,N_1995);
nand U2084 (N_2084,N_1911,N_1864);
or U2085 (N_2085,N_1962,N_1976);
and U2086 (N_2086,N_1840,N_1828);
and U2087 (N_2087,N_1960,N_1956);
xnor U2088 (N_2088,N_1875,N_1950);
or U2089 (N_2089,N_1826,N_1838);
xnor U2090 (N_2090,N_1985,N_1965);
xnor U2091 (N_2091,N_1969,N_1894);
xnor U2092 (N_2092,N_1893,N_1902);
and U2093 (N_2093,N_1922,N_1993);
nor U2094 (N_2094,N_1802,N_1804);
and U2095 (N_2095,N_1892,N_1975);
xor U2096 (N_2096,N_1809,N_1933);
and U2097 (N_2097,N_1897,N_1931);
xnor U2098 (N_2098,N_1901,N_1835);
xor U2099 (N_2099,N_1850,N_1958);
or U2100 (N_2100,N_1846,N_1982);
nor U2101 (N_2101,N_1991,N_1889);
nand U2102 (N_2102,N_1872,N_1971);
nand U2103 (N_2103,N_1815,N_1997);
nor U2104 (N_2104,N_1992,N_1842);
and U2105 (N_2105,N_1874,N_1826);
nor U2106 (N_2106,N_1868,N_1941);
nand U2107 (N_2107,N_1919,N_1860);
nand U2108 (N_2108,N_1861,N_1999);
xor U2109 (N_2109,N_1806,N_1906);
xnor U2110 (N_2110,N_1948,N_1903);
or U2111 (N_2111,N_1838,N_1895);
and U2112 (N_2112,N_1902,N_1959);
xor U2113 (N_2113,N_1894,N_1962);
nor U2114 (N_2114,N_1862,N_1875);
or U2115 (N_2115,N_1804,N_1949);
nand U2116 (N_2116,N_1902,N_1970);
nand U2117 (N_2117,N_1981,N_1949);
or U2118 (N_2118,N_1894,N_1933);
nand U2119 (N_2119,N_1915,N_1868);
xor U2120 (N_2120,N_1841,N_1875);
or U2121 (N_2121,N_1973,N_1943);
and U2122 (N_2122,N_1875,N_1980);
or U2123 (N_2123,N_1895,N_1804);
nand U2124 (N_2124,N_1977,N_1948);
nor U2125 (N_2125,N_1922,N_1894);
and U2126 (N_2126,N_1997,N_1816);
and U2127 (N_2127,N_1887,N_1825);
nand U2128 (N_2128,N_1887,N_1964);
or U2129 (N_2129,N_1970,N_1911);
nor U2130 (N_2130,N_1982,N_1827);
nand U2131 (N_2131,N_1866,N_1807);
nor U2132 (N_2132,N_1934,N_1860);
and U2133 (N_2133,N_1995,N_1876);
xnor U2134 (N_2134,N_1840,N_1910);
xor U2135 (N_2135,N_1895,N_1986);
and U2136 (N_2136,N_1899,N_1890);
nand U2137 (N_2137,N_1813,N_1807);
or U2138 (N_2138,N_1999,N_1888);
or U2139 (N_2139,N_1845,N_1807);
or U2140 (N_2140,N_1953,N_1834);
xnor U2141 (N_2141,N_1996,N_1907);
xnor U2142 (N_2142,N_1984,N_1892);
xor U2143 (N_2143,N_1823,N_1867);
xor U2144 (N_2144,N_1830,N_1978);
and U2145 (N_2145,N_1981,N_1833);
and U2146 (N_2146,N_1861,N_1980);
nor U2147 (N_2147,N_1978,N_1912);
or U2148 (N_2148,N_1922,N_1994);
xnor U2149 (N_2149,N_1856,N_1816);
and U2150 (N_2150,N_1923,N_1977);
xnor U2151 (N_2151,N_1888,N_1966);
nor U2152 (N_2152,N_1871,N_1836);
xor U2153 (N_2153,N_1892,N_1955);
or U2154 (N_2154,N_1890,N_1989);
nor U2155 (N_2155,N_1828,N_1843);
nor U2156 (N_2156,N_1918,N_1800);
and U2157 (N_2157,N_1878,N_1833);
nand U2158 (N_2158,N_1819,N_1958);
or U2159 (N_2159,N_1915,N_1946);
and U2160 (N_2160,N_1951,N_1834);
or U2161 (N_2161,N_1876,N_1806);
and U2162 (N_2162,N_1877,N_1834);
and U2163 (N_2163,N_1957,N_1993);
and U2164 (N_2164,N_1890,N_1868);
nand U2165 (N_2165,N_1993,N_1982);
nand U2166 (N_2166,N_1947,N_1930);
nor U2167 (N_2167,N_1839,N_1899);
or U2168 (N_2168,N_1932,N_1997);
or U2169 (N_2169,N_1826,N_1939);
or U2170 (N_2170,N_1836,N_1983);
xnor U2171 (N_2171,N_1908,N_1828);
nor U2172 (N_2172,N_1852,N_1807);
nand U2173 (N_2173,N_1917,N_1972);
and U2174 (N_2174,N_1916,N_1956);
or U2175 (N_2175,N_1846,N_1895);
nor U2176 (N_2176,N_1867,N_1976);
xnor U2177 (N_2177,N_1969,N_1804);
nor U2178 (N_2178,N_1988,N_1905);
or U2179 (N_2179,N_1845,N_1859);
nand U2180 (N_2180,N_1953,N_1980);
or U2181 (N_2181,N_1878,N_1829);
nor U2182 (N_2182,N_1857,N_1849);
and U2183 (N_2183,N_1922,N_1843);
xor U2184 (N_2184,N_1829,N_1927);
and U2185 (N_2185,N_1910,N_1990);
or U2186 (N_2186,N_1871,N_1966);
or U2187 (N_2187,N_1809,N_1919);
nor U2188 (N_2188,N_1854,N_1943);
nor U2189 (N_2189,N_1999,N_1877);
nor U2190 (N_2190,N_1880,N_1951);
nor U2191 (N_2191,N_1964,N_1862);
or U2192 (N_2192,N_1931,N_1959);
nand U2193 (N_2193,N_1889,N_1940);
nand U2194 (N_2194,N_1967,N_1871);
nand U2195 (N_2195,N_1835,N_1882);
nand U2196 (N_2196,N_1853,N_1958);
or U2197 (N_2197,N_1973,N_1940);
or U2198 (N_2198,N_1910,N_1811);
or U2199 (N_2199,N_1918,N_1936);
nor U2200 (N_2200,N_2156,N_2014);
nand U2201 (N_2201,N_2154,N_2129);
nor U2202 (N_2202,N_2125,N_2009);
or U2203 (N_2203,N_2052,N_2019);
or U2204 (N_2204,N_2101,N_2090);
nand U2205 (N_2205,N_2073,N_2152);
nor U2206 (N_2206,N_2078,N_2170);
xnor U2207 (N_2207,N_2095,N_2040);
and U2208 (N_2208,N_2144,N_2108);
nor U2209 (N_2209,N_2077,N_2146);
and U2210 (N_2210,N_2157,N_2074);
or U2211 (N_2211,N_2091,N_2030);
nand U2212 (N_2212,N_2048,N_2192);
nand U2213 (N_2213,N_2069,N_2173);
and U2214 (N_2214,N_2160,N_2168);
or U2215 (N_2215,N_2049,N_2149);
nor U2216 (N_2216,N_2135,N_2122);
nor U2217 (N_2217,N_2041,N_2183);
xor U2218 (N_2218,N_2169,N_2057);
nor U2219 (N_2219,N_2008,N_2109);
and U2220 (N_2220,N_2116,N_2034);
nand U2221 (N_2221,N_2177,N_2071);
xor U2222 (N_2222,N_2143,N_2191);
and U2223 (N_2223,N_2079,N_2139);
and U2224 (N_2224,N_2059,N_2176);
and U2225 (N_2225,N_2010,N_2188);
nand U2226 (N_2226,N_2136,N_2118);
or U2227 (N_2227,N_2174,N_2134);
or U2228 (N_2228,N_2063,N_2096);
or U2229 (N_2229,N_2054,N_2179);
xor U2230 (N_2230,N_2004,N_2138);
xnor U2231 (N_2231,N_2025,N_2151);
or U2232 (N_2232,N_2092,N_2023);
and U2233 (N_2233,N_2072,N_2158);
xor U2234 (N_2234,N_2032,N_2197);
nand U2235 (N_2235,N_2044,N_2194);
nand U2236 (N_2236,N_2042,N_2015);
or U2237 (N_2237,N_2083,N_2130);
xor U2238 (N_2238,N_2022,N_2126);
nand U2239 (N_2239,N_2045,N_2112);
and U2240 (N_2240,N_2159,N_2120);
and U2241 (N_2241,N_2127,N_2186);
and U2242 (N_2242,N_2180,N_2086);
or U2243 (N_2243,N_2181,N_2142);
and U2244 (N_2244,N_2094,N_2098);
nor U2245 (N_2245,N_2145,N_2141);
nor U2246 (N_2246,N_2187,N_2148);
nor U2247 (N_2247,N_2002,N_2164);
or U2248 (N_2248,N_2161,N_2106);
nor U2249 (N_2249,N_2012,N_2062);
nand U2250 (N_2250,N_2171,N_2036);
xor U2251 (N_2251,N_2113,N_2163);
xnor U2252 (N_2252,N_2123,N_2155);
nand U2253 (N_2253,N_2001,N_2060);
or U2254 (N_2254,N_2137,N_2172);
nand U2255 (N_2255,N_2165,N_2026);
and U2256 (N_2256,N_2190,N_2024);
nor U2257 (N_2257,N_2064,N_2140);
nand U2258 (N_2258,N_2029,N_2153);
xor U2259 (N_2259,N_2018,N_2147);
xnor U2260 (N_2260,N_2035,N_2028);
nand U2261 (N_2261,N_2020,N_2075);
xnor U2262 (N_2262,N_2115,N_2085);
xor U2263 (N_2263,N_2124,N_2082);
nand U2264 (N_2264,N_2076,N_2175);
and U2265 (N_2265,N_2066,N_2110);
nor U2266 (N_2266,N_2097,N_2043);
xnor U2267 (N_2267,N_2102,N_2021);
or U2268 (N_2268,N_2111,N_2117);
and U2269 (N_2269,N_2031,N_2099);
nor U2270 (N_2270,N_2070,N_2055);
nand U2271 (N_2271,N_2038,N_2166);
or U2272 (N_2272,N_2058,N_2119);
or U2273 (N_2273,N_2016,N_2093);
and U2274 (N_2274,N_2162,N_2013);
nand U2275 (N_2275,N_2185,N_2065);
and U2276 (N_2276,N_2103,N_2087);
nor U2277 (N_2277,N_2128,N_2131);
nor U2278 (N_2278,N_2182,N_2017);
xnor U2279 (N_2279,N_2051,N_2189);
xor U2280 (N_2280,N_2105,N_2089);
xnor U2281 (N_2281,N_2100,N_2056);
nand U2282 (N_2282,N_2000,N_2050);
nand U2283 (N_2283,N_2121,N_2053);
and U2284 (N_2284,N_2133,N_2150);
nand U2285 (N_2285,N_2084,N_2037);
or U2286 (N_2286,N_2039,N_2107);
or U2287 (N_2287,N_2199,N_2198);
or U2288 (N_2288,N_2104,N_2033);
nor U2289 (N_2289,N_2067,N_2081);
or U2290 (N_2290,N_2007,N_2193);
xnor U2291 (N_2291,N_2068,N_2003);
xor U2292 (N_2292,N_2005,N_2132);
nor U2293 (N_2293,N_2080,N_2011);
and U2294 (N_2294,N_2061,N_2178);
and U2295 (N_2295,N_2088,N_2196);
and U2296 (N_2296,N_2195,N_2027);
nand U2297 (N_2297,N_2184,N_2006);
xnor U2298 (N_2298,N_2047,N_2167);
xnor U2299 (N_2299,N_2114,N_2046);
nor U2300 (N_2300,N_2187,N_2076);
and U2301 (N_2301,N_2014,N_2143);
and U2302 (N_2302,N_2020,N_2197);
and U2303 (N_2303,N_2081,N_2024);
nand U2304 (N_2304,N_2174,N_2009);
xor U2305 (N_2305,N_2187,N_2120);
nor U2306 (N_2306,N_2024,N_2197);
and U2307 (N_2307,N_2180,N_2013);
or U2308 (N_2308,N_2174,N_2083);
or U2309 (N_2309,N_2198,N_2045);
xor U2310 (N_2310,N_2082,N_2097);
and U2311 (N_2311,N_2001,N_2182);
nor U2312 (N_2312,N_2043,N_2141);
nor U2313 (N_2313,N_2005,N_2131);
xor U2314 (N_2314,N_2186,N_2048);
nand U2315 (N_2315,N_2039,N_2101);
and U2316 (N_2316,N_2122,N_2134);
and U2317 (N_2317,N_2134,N_2192);
or U2318 (N_2318,N_2029,N_2121);
nand U2319 (N_2319,N_2172,N_2035);
nand U2320 (N_2320,N_2074,N_2160);
xor U2321 (N_2321,N_2118,N_2025);
xnor U2322 (N_2322,N_2052,N_2158);
nor U2323 (N_2323,N_2158,N_2007);
nand U2324 (N_2324,N_2103,N_2080);
xnor U2325 (N_2325,N_2090,N_2130);
nand U2326 (N_2326,N_2039,N_2158);
nand U2327 (N_2327,N_2046,N_2061);
nor U2328 (N_2328,N_2189,N_2108);
nand U2329 (N_2329,N_2152,N_2008);
nand U2330 (N_2330,N_2016,N_2033);
or U2331 (N_2331,N_2137,N_2125);
or U2332 (N_2332,N_2041,N_2085);
and U2333 (N_2333,N_2115,N_2017);
nand U2334 (N_2334,N_2063,N_2014);
or U2335 (N_2335,N_2075,N_2066);
xnor U2336 (N_2336,N_2069,N_2197);
xor U2337 (N_2337,N_2164,N_2138);
and U2338 (N_2338,N_2193,N_2084);
xnor U2339 (N_2339,N_2034,N_2058);
or U2340 (N_2340,N_2044,N_2063);
nor U2341 (N_2341,N_2108,N_2124);
and U2342 (N_2342,N_2035,N_2021);
and U2343 (N_2343,N_2049,N_2158);
and U2344 (N_2344,N_2024,N_2139);
nand U2345 (N_2345,N_2144,N_2129);
or U2346 (N_2346,N_2137,N_2138);
nand U2347 (N_2347,N_2055,N_2107);
nor U2348 (N_2348,N_2058,N_2101);
xnor U2349 (N_2349,N_2173,N_2049);
xnor U2350 (N_2350,N_2072,N_2150);
nor U2351 (N_2351,N_2031,N_2018);
and U2352 (N_2352,N_2011,N_2005);
xor U2353 (N_2353,N_2074,N_2178);
and U2354 (N_2354,N_2146,N_2041);
nor U2355 (N_2355,N_2053,N_2097);
nand U2356 (N_2356,N_2142,N_2178);
or U2357 (N_2357,N_2065,N_2059);
nand U2358 (N_2358,N_2112,N_2061);
or U2359 (N_2359,N_2084,N_2050);
nor U2360 (N_2360,N_2015,N_2079);
xnor U2361 (N_2361,N_2197,N_2007);
xor U2362 (N_2362,N_2044,N_2052);
nor U2363 (N_2363,N_2082,N_2065);
xnor U2364 (N_2364,N_2151,N_2164);
nor U2365 (N_2365,N_2172,N_2079);
nand U2366 (N_2366,N_2184,N_2175);
and U2367 (N_2367,N_2027,N_2183);
xor U2368 (N_2368,N_2066,N_2109);
or U2369 (N_2369,N_2122,N_2007);
nor U2370 (N_2370,N_2031,N_2022);
nor U2371 (N_2371,N_2113,N_2134);
or U2372 (N_2372,N_2177,N_2031);
nand U2373 (N_2373,N_2053,N_2083);
xor U2374 (N_2374,N_2014,N_2000);
and U2375 (N_2375,N_2176,N_2086);
nor U2376 (N_2376,N_2196,N_2069);
xor U2377 (N_2377,N_2013,N_2137);
xnor U2378 (N_2378,N_2100,N_2113);
xor U2379 (N_2379,N_2003,N_2164);
nor U2380 (N_2380,N_2012,N_2189);
nand U2381 (N_2381,N_2082,N_2128);
nor U2382 (N_2382,N_2062,N_2176);
nor U2383 (N_2383,N_2146,N_2090);
xnor U2384 (N_2384,N_2147,N_2110);
and U2385 (N_2385,N_2055,N_2174);
or U2386 (N_2386,N_2176,N_2105);
nand U2387 (N_2387,N_2019,N_2079);
nor U2388 (N_2388,N_2158,N_2128);
nor U2389 (N_2389,N_2036,N_2178);
xor U2390 (N_2390,N_2041,N_2023);
or U2391 (N_2391,N_2108,N_2198);
nand U2392 (N_2392,N_2113,N_2101);
or U2393 (N_2393,N_2026,N_2010);
nand U2394 (N_2394,N_2079,N_2098);
or U2395 (N_2395,N_2163,N_2072);
or U2396 (N_2396,N_2023,N_2175);
nand U2397 (N_2397,N_2048,N_2098);
nor U2398 (N_2398,N_2023,N_2125);
xnor U2399 (N_2399,N_2178,N_2044);
nor U2400 (N_2400,N_2363,N_2225);
and U2401 (N_2401,N_2377,N_2354);
nor U2402 (N_2402,N_2235,N_2381);
or U2403 (N_2403,N_2229,N_2378);
or U2404 (N_2404,N_2216,N_2215);
xor U2405 (N_2405,N_2246,N_2355);
xor U2406 (N_2406,N_2301,N_2226);
or U2407 (N_2407,N_2283,N_2277);
nand U2408 (N_2408,N_2324,N_2273);
xnor U2409 (N_2409,N_2268,N_2334);
nand U2410 (N_2410,N_2349,N_2389);
xnor U2411 (N_2411,N_2206,N_2285);
nor U2412 (N_2412,N_2234,N_2364);
and U2413 (N_2413,N_2244,N_2238);
nor U2414 (N_2414,N_2331,N_2221);
nor U2415 (N_2415,N_2306,N_2272);
and U2416 (N_2416,N_2232,N_2298);
nand U2417 (N_2417,N_2304,N_2311);
xnor U2418 (N_2418,N_2382,N_2371);
nor U2419 (N_2419,N_2274,N_2386);
xnor U2420 (N_2420,N_2217,N_2295);
and U2421 (N_2421,N_2394,N_2322);
nand U2422 (N_2422,N_2296,N_2200);
nand U2423 (N_2423,N_2271,N_2224);
nor U2424 (N_2424,N_2258,N_2208);
xor U2425 (N_2425,N_2280,N_2313);
and U2426 (N_2426,N_2310,N_2275);
and U2427 (N_2427,N_2319,N_2211);
or U2428 (N_2428,N_2305,N_2372);
nor U2429 (N_2429,N_2312,N_2250);
xnor U2430 (N_2430,N_2366,N_2395);
nand U2431 (N_2431,N_2264,N_2332);
nand U2432 (N_2432,N_2262,N_2210);
and U2433 (N_2433,N_2257,N_2228);
nor U2434 (N_2434,N_2352,N_2202);
nand U2435 (N_2435,N_2241,N_2237);
xnor U2436 (N_2436,N_2397,N_2392);
nand U2437 (N_2437,N_2353,N_2203);
xor U2438 (N_2438,N_2270,N_2309);
xor U2439 (N_2439,N_2279,N_2209);
nand U2440 (N_2440,N_2287,N_2205);
nand U2441 (N_2441,N_2333,N_2370);
nand U2442 (N_2442,N_2359,N_2335);
and U2443 (N_2443,N_2385,N_2391);
nand U2444 (N_2444,N_2214,N_2259);
and U2445 (N_2445,N_2323,N_2218);
nand U2446 (N_2446,N_2297,N_2294);
and U2447 (N_2447,N_2346,N_2360);
or U2448 (N_2448,N_2384,N_2222);
and U2449 (N_2449,N_2236,N_2293);
nor U2450 (N_2450,N_2343,N_2252);
and U2451 (N_2451,N_2338,N_2329);
xnor U2452 (N_2452,N_2248,N_2340);
nor U2453 (N_2453,N_2336,N_2373);
nand U2454 (N_2454,N_2266,N_2227);
or U2455 (N_2455,N_2263,N_2289);
and U2456 (N_2456,N_2220,N_2302);
xor U2457 (N_2457,N_2219,N_2253);
nor U2458 (N_2458,N_2230,N_2328);
xor U2459 (N_2459,N_2251,N_2292);
nor U2460 (N_2460,N_2369,N_2278);
and U2461 (N_2461,N_2314,N_2291);
or U2462 (N_2462,N_2325,N_2288);
or U2463 (N_2463,N_2256,N_2357);
nor U2464 (N_2464,N_2327,N_2265);
or U2465 (N_2465,N_2269,N_2290);
nand U2466 (N_2466,N_2342,N_2339);
xor U2467 (N_2467,N_2337,N_2380);
nor U2468 (N_2468,N_2233,N_2347);
and U2469 (N_2469,N_2223,N_2242);
nand U2470 (N_2470,N_2390,N_2308);
nand U2471 (N_2471,N_2383,N_2345);
and U2472 (N_2472,N_2368,N_2320);
nor U2473 (N_2473,N_2286,N_2261);
xnor U2474 (N_2474,N_2387,N_2321);
and U2475 (N_2475,N_2361,N_2303);
xor U2476 (N_2476,N_2276,N_2300);
or U2477 (N_2477,N_2240,N_2375);
xor U2478 (N_2478,N_2398,N_2358);
xor U2479 (N_2479,N_2362,N_2254);
xnor U2480 (N_2480,N_2316,N_2284);
nor U2481 (N_2481,N_2330,N_2213);
and U2482 (N_2482,N_2318,N_2212);
xor U2483 (N_2483,N_2374,N_2245);
xnor U2484 (N_2484,N_2396,N_2239);
nor U2485 (N_2485,N_2367,N_2393);
or U2486 (N_2486,N_2243,N_2341);
nand U2487 (N_2487,N_2260,N_2365);
or U2488 (N_2488,N_2231,N_2201);
nor U2489 (N_2489,N_2207,N_2351);
or U2490 (N_2490,N_2315,N_2348);
xor U2491 (N_2491,N_2299,N_2204);
or U2492 (N_2492,N_2379,N_2350);
and U2493 (N_2493,N_2267,N_2388);
xnor U2494 (N_2494,N_2255,N_2281);
nor U2495 (N_2495,N_2326,N_2249);
or U2496 (N_2496,N_2307,N_2247);
or U2497 (N_2497,N_2282,N_2399);
nand U2498 (N_2498,N_2356,N_2344);
or U2499 (N_2499,N_2317,N_2376);
or U2500 (N_2500,N_2255,N_2261);
and U2501 (N_2501,N_2374,N_2270);
and U2502 (N_2502,N_2284,N_2300);
nor U2503 (N_2503,N_2364,N_2380);
xnor U2504 (N_2504,N_2351,N_2217);
or U2505 (N_2505,N_2237,N_2398);
and U2506 (N_2506,N_2212,N_2383);
nand U2507 (N_2507,N_2308,N_2248);
xor U2508 (N_2508,N_2348,N_2339);
and U2509 (N_2509,N_2388,N_2256);
xnor U2510 (N_2510,N_2253,N_2236);
and U2511 (N_2511,N_2329,N_2378);
and U2512 (N_2512,N_2287,N_2297);
or U2513 (N_2513,N_2226,N_2390);
nand U2514 (N_2514,N_2388,N_2329);
nor U2515 (N_2515,N_2381,N_2393);
or U2516 (N_2516,N_2398,N_2212);
or U2517 (N_2517,N_2387,N_2368);
nor U2518 (N_2518,N_2351,N_2379);
nor U2519 (N_2519,N_2342,N_2284);
and U2520 (N_2520,N_2391,N_2375);
and U2521 (N_2521,N_2386,N_2384);
xor U2522 (N_2522,N_2331,N_2380);
and U2523 (N_2523,N_2227,N_2361);
xor U2524 (N_2524,N_2338,N_2284);
or U2525 (N_2525,N_2255,N_2301);
xor U2526 (N_2526,N_2224,N_2251);
nor U2527 (N_2527,N_2271,N_2376);
nand U2528 (N_2528,N_2297,N_2304);
xor U2529 (N_2529,N_2209,N_2203);
or U2530 (N_2530,N_2237,N_2385);
nand U2531 (N_2531,N_2364,N_2209);
or U2532 (N_2532,N_2396,N_2254);
nor U2533 (N_2533,N_2310,N_2348);
or U2534 (N_2534,N_2303,N_2214);
nor U2535 (N_2535,N_2395,N_2343);
nand U2536 (N_2536,N_2210,N_2249);
nor U2537 (N_2537,N_2354,N_2378);
xor U2538 (N_2538,N_2340,N_2321);
nor U2539 (N_2539,N_2209,N_2349);
or U2540 (N_2540,N_2319,N_2242);
nand U2541 (N_2541,N_2341,N_2220);
or U2542 (N_2542,N_2388,N_2360);
nand U2543 (N_2543,N_2356,N_2392);
and U2544 (N_2544,N_2320,N_2296);
xnor U2545 (N_2545,N_2388,N_2304);
nor U2546 (N_2546,N_2221,N_2211);
and U2547 (N_2547,N_2357,N_2266);
nor U2548 (N_2548,N_2285,N_2293);
nor U2549 (N_2549,N_2330,N_2377);
xnor U2550 (N_2550,N_2287,N_2317);
or U2551 (N_2551,N_2270,N_2378);
xor U2552 (N_2552,N_2321,N_2227);
nor U2553 (N_2553,N_2367,N_2377);
nor U2554 (N_2554,N_2257,N_2277);
nand U2555 (N_2555,N_2363,N_2266);
nor U2556 (N_2556,N_2360,N_2210);
nand U2557 (N_2557,N_2320,N_2244);
xnor U2558 (N_2558,N_2301,N_2361);
nand U2559 (N_2559,N_2370,N_2283);
xnor U2560 (N_2560,N_2327,N_2336);
or U2561 (N_2561,N_2256,N_2274);
and U2562 (N_2562,N_2373,N_2287);
nand U2563 (N_2563,N_2252,N_2239);
or U2564 (N_2564,N_2304,N_2318);
or U2565 (N_2565,N_2399,N_2372);
and U2566 (N_2566,N_2358,N_2345);
or U2567 (N_2567,N_2238,N_2362);
nand U2568 (N_2568,N_2290,N_2260);
and U2569 (N_2569,N_2288,N_2368);
and U2570 (N_2570,N_2222,N_2262);
xnor U2571 (N_2571,N_2243,N_2221);
or U2572 (N_2572,N_2261,N_2377);
nand U2573 (N_2573,N_2378,N_2243);
nand U2574 (N_2574,N_2271,N_2331);
or U2575 (N_2575,N_2267,N_2308);
xor U2576 (N_2576,N_2362,N_2310);
nand U2577 (N_2577,N_2289,N_2275);
or U2578 (N_2578,N_2270,N_2240);
xnor U2579 (N_2579,N_2387,N_2303);
nand U2580 (N_2580,N_2343,N_2368);
xor U2581 (N_2581,N_2291,N_2302);
and U2582 (N_2582,N_2221,N_2386);
xnor U2583 (N_2583,N_2223,N_2317);
xnor U2584 (N_2584,N_2310,N_2301);
nor U2585 (N_2585,N_2349,N_2323);
or U2586 (N_2586,N_2367,N_2395);
or U2587 (N_2587,N_2312,N_2325);
or U2588 (N_2588,N_2282,N_2269);
nor U2589 (N_2589,N_2292,N_2268);
or U2590 (N_2590,N_2394,N_2202);
xnor U2591 (N_2591,N_2372,N_2286);
nand U2592 (N_2592,N_2297,N_2291);
nor U2593 (N_2593,N_2371,N_2300);
nor U2594 (N_2594,N_2309,N_2212);
nor U2595 (N_2595,N_2221,N_2337);
nor U2596 (N_2596,N_2363,N_2257);
nand U2597 (N_2597,N_2367,N_2311);
nand U2598 (N_2598,N_2334,N_2284);
and U2599 (N_2599,N_2286,N_2270);
xor U2600 (N_2600,N_2545,N_2560);
or U2601 (N_2601,N_2446,N_2430);
nor U2602 (N_2602,N_2599,N_2436);
xnor U2603 (N_2603,N_2571,N_2403);
nand U2604 (N_2604,N_2514,N_2416);
nor U2605 (N_2605,N_2561,N_2562);
and U2606 (N_2606,N_2517,N_2563);
xnor U2607 (N_2607,N_2508,N_2434);
nand U2608 (N_2608,N_2598,N_2455);
nor U2609 (N_2609,N_2539,N_2490);
nand U2610 (N_2610,N_2529,N_2590);
and U2611 (N_2611,N_2537,N_2462);
xor U2612 (N_2612,N_2536,N_2445);
and U2613 (N_2613,N_2484,N_2573);
xor U2614 (N_2614,N_2465,N_2415);
and U2615 (N_2615,N_2466,N_2477);
and U2616 (N_2616,N_2404,N_2450);
and U2617 (N_2617,N_2593,N_2554);
nand U2618 (N_2618,N_2471,N_2497);
xnor U2619 (N_2619,N_2424,N_2583);
xor U2620 (N_2620,N_2475,N_2582);
or U2621 (N_2621,N_2505,N_2542);
or U2622 (N_2622,N_2578,N_2486);
nor U2623 (N_2623,N_2451,N_2531);
nand U2624 (N_2624,N_2534,N_2487);
and U2625 (N_2625,N_2572,N_2511);
nand U2626 (N_2626,N_2480,N_2589);
nand U2627 (N_2627,N_2488,N_2453);
and U2628 (N_2628,N_2557,N_2525);
xor U2629 (N_2629,N_2584,N_2526);
nand U2630 (N_2630,N_2425,N_2500);
nand U2631 (N_2631,N_2570,N_2524);
and U2632 (N_2632,N_2577,N_2468);
nand U2633 (N_2633,N_2550,N_2555);
or U2634 (N_2634,N_2489,N_2421);
nor U2635 (N_2635,N_2454,N_2540);
or U2636 (N_2636,N_2433,N_2512);
nor U2637 (N_2637,N_2469,N_2513);
or U2638 (N_2638,N_2479,N_2410);
and U2639 (N_2639,N_2429,N_2470);
nand U2640 (N_2640,N_2478,N_2442);
xor U2641 (N_2641,N_2543,N_2575);
nor U2642 (N_2642,N_2413,N_2595);
or U2643 (N_2643,N_2435,N_2432);
nor U2644 (N_2644,N_2581,N_2426);
and U2645 (N_2645,N_2585,N_2541);
xor U2646 (N_2646,N_2499,N_2519);
and U2647 (N_2647,N_2516,N_2548);
and U2648 (N_2648,N_2461,N_2501);
and U2649 (N_2649,N_2552,N_2408);
and U2650 (N_2650,N_2483,N_2456);
nor U2651 (N_2651,N_2522,N_2579);
nor U2652 (N_2652,N_2460,N_2472);
xnor U2653 (N_2653,N_2504,N_2444);
xor U2654 (N_2654,N_2503,N_2564);
nor U2655 (N_2655,N_2439,N_2464);
or U2656 (N_2656,N_2457,N_2482);
nand U2657 (N_2657,N_2586,N_2515);
and U2658 (N_2658,N_2414,N_2588);
nor U2659 (N_2659,N_2574,N_2565);
and U2660 (N_2660,N_2447,N_2509);
nand U2661 (N_2661,N_2594,N_2474);
and U2662 (N_2662,N_2449,N_2441);
nand U2663 (N_2663,N_2507,N_2559);
and U2664 (N_2664,N_2587,N_2544);
nand U2665 (N_2665,N_2580,N_2418);
xor U2666 (N_2666,N_2530,N_2576);
nor U2667 (N_2667,N_2440,N_2431);
xnor U2668 (N_2668,N_2496,N_2420);
or U2669 (N_2669,N_2506,N_2538);
nor U2670 (N_2670,N_2568,N_2467);
and U2671 (N_2671,N_2405,N_2528);
nor U2672 (N_2672,N_2402,N_2553);
xor U2673 (N_2673,N_2411,N_2492);
xnor U2674 (N_2674,N_2566,N_2494);
nor U2675 (N_2675,N_2567,N_2422);
nor U2676 (N_2676,N_2556,N_2448);
nand U2677 (N_2677,N_2401,N_2532);
nor U2678 (N_2678,N_2452,N_2438);
and U2679 (N_2679,N_2510,N_2407);
and U2680 (N_2680,N_2521,N_2591);
xnor U2681 (N_2681,N_2428,N_2409);
nand U2682 (N_2682,N_2535,N_2527);
nor U2683 (N_2683,N_2592,N_2596);
or U2684 (N_2684,N_2558,N_2495);
nand U2685 (N_2685,N_2476,N_2459);
nor U2686 (N_2686,N_2502,N_2518);
xnor U2687 (N_2687,N_2400,N_2437);
xnor U2688 (N_2688,N_2463,N_2443);
nor U2689 (N_2689,N_2481,N_2458);
and U2690 (N_2690,N_2549,N_2427);
and U2691 (N_2691,N_2569,N_2419);
xnor U2692 (N_2692,N_2417,N_2406);
xor U2693 (N_2693,N_2533,N_2473);
nor U2694 (N_2694,N_2547,N_2520);
nand U2695 (N_2695,N_2597,N_2412);
nor U2696 (N_2696,N_2523,N_2485);
nor U2697 (N_2697,N_2551,N_2546);
or U2698 (N_2698,N_2423,N_2498);
and U2699 (N_2699,N_2493,N_2491);
nand U2700 (N_2700,N_2413,N_2580);
nand U2701 (N_2701,N_2574,N_2538);
or U2702 (N_2702,N_2442,N_2422);
xor U2703 (N_2703,N_2599,N_2487);
or U2704 (N_2704,N_2495,N_2530);
and U2705 (N_2705,N_2561,N_2557);
nor U2706 (N_2706,N_2570,N_2582);
or U2707 (N_2707,N_2532,N_2567);
xor U2708 (N_2708,N_2432,N_2400);
nor U2709 (N_2709,N_2538,N_2588);
nand U2710 (N_2710,N_2524,N_2487);
nand U2711 (N_2711,N_2511,N_2414);
and U2712 (N_2712,N_2504,N_2511);
nor U2713 (N_2713,N_2524,N_2466);
nor U2714 (N_2714,N_2502,N_2475);
or U2715 (N_2715,N_2588,N_2469);
nor U2716 (N_2716,N_2565,N_2429);
or U2717 (N_2717,N_2407,N_2431);
and U2718 (N_2718,N_2547,N_2480);
and U2719 (N_2719,N_2585,N_2431);
or U2720 (N_2720,N_2426,N_2434);
or U2721 (N_2721,N_2502,N_2468);
and U2722 (N_2722,N_2442,N_2514);
xor U2723 (N_2723,N_2432,N_2410);
and U2724 (N_2724,N_2489,N_2574);
nand U2725 (N_2725,N_2424,N_2574);
nand U2726 (N_2726,N_2453,N_2575);
nor U2727 (N_2727,N_2444,N_2414);
xnor U2728 (N_2728,N_2586,N_2525);
nor U2729 (N_2729,N_2555,N_2467);
and U2730 (N_2730,N_2483,N_2505);
and U2731 (N_2731,N_2541,N_2592);
or U2732 (N_2732,N_2491,N_2588);
xor U2733 (N_2733,N_2551,N_2508);
and U2734 (N_2734,N_2588,N_2592);
xor U2735 (N_2735,N_2441,N_2580);
xnor U2736 (N_2736,N_2470,N_2449);
nor U2737 (N_2737,N_2538,N_2459);
xnor U2738 (N_2738,N_2546,N_2515);
xor U2739 (N_2739,N_2422,N_2406);
xnor U2740 (N_2740,N_2483,N_2508);
xor U2741 (N_2741,N_2556,N_2548);
or U2742 (N_2742,N_2456,N_2410);
and U2743 (N_2743,N_2459,N_2411);
or U2744 (N_2744,N_2413,N_2545);
xor U2745 (N_2745,N_2584,N_2479);
nand U2746 (N_2746,N_2521,N_2485);
nor U2747 (N_2747,N_2554,N_2493);
or U2748 (N_2748,N_2498,N_2583);
nand U2749 (N_2749,N_2536,N_2431);
nor U2750 (N_2750,N_2522,N_2488);
nand U2751 (N_2751,N_2536,N_2507);
nor U2752 (N_2752,N_2507,N_2552);
and U2753 (N_2753,N_2427,N_2491);
or U2754 (N_2754,N_2433,N_2407);
or U2755 (N_2755,N_2416,N_2453);
or U2756 (N_2756,N_2484,N_2490);
nand U2757 (N_2757,N_2492,N_2403);
and U2758 (N_2758,N_2496,N_2411);
xor U2759 (N_2759,N_2435,N_2536);
nand U2760 (N_2760,N_2524,N_2585);
xnor U2761 (N_2761,N_2489,N_2416);
nor U2762 (N_2762,N_2516,N_2463);
nand U2763 (N_2763,N_2524,N_2593);
nor U2764 (N_2764,N_2588,N_2584);
and U2765 (N_2765,N_2502,N_2541);
nand U2766 (N_2766,N_2550,N_2403);
xor U2767 (N_2767,N_2464,N_2460);
xnor U2768 (N_2768,N_2453,N_2478);
and U2769 (N_2769,N_2594,N_2568);
nor U2770 (N_2770,N_2500,N_2597);
xnor U2771 (N_2771,N_2492,N_2500);
xnor U2772 (N_2772,N_2447,N_2557);
xnor U2773 (N_2773,N_2556,N_2402);
nor U2774 (N_2774,N_2591,N_2580);
and U2775 (N_2775,N_2443,N_2497);
xor U2776 (N_2776,N_2507,N_2529);
nand U2777 (N_2777,N_2525,N_2400);
or U2778 (N_2778,N_2479,N_2443);
xor U2779 (N_2779,N_2594,N_2443);
xnor U2780 (N_2780,N_2483,N_2470);
or U2781 (N_2781,N_2431,N_2492);
nand U2782 (N_2782,N_2419,N_2470);
nor U2783 (N_2783,N_2470,N_2473);
nor U2784 (N_2784,N_2417,N_2469);
or U2785 (N_2785,N_2409,N_2534);
nor U2786 (N_2786,N_2506,N_2534);
nand U2787 (N_2787,N_2436,N_2469);
nor U2788 (N_2788,N_2573,N_2532);
nand U2789 (N_2789,N_2573,N_2498);
and U2790 (N_2790,N_2471,N_2520);
or U2791 (N_2791,N_2439,N_2450);
nand U2792 (N_2792,N_2573,N_2490);
nor U2793 (N_2793,N_2542,N_2529);
and U2794 (N_2794,N_2591,N_2582);
and U2795 (N_2795,N_2571,N_2560);
nor U2796 (N_2796,N_2469,N_2418);
and U2797 (N_2797,N_2431,N_2497);
xor U2798 (N_2798,N_2532,N_2575);
and U2799 (N_2799,N_2561,N_2560);
nor U2800 (N_2800,N_2662,N_2785);
nand U2801 (N_2801,N_2631,N_2646);
xnor U2802 (N_2802,N_2652,N_2738);
xor U2803 (N_2803,N_2676,N_2601);
nor U2804 (N_2804,N_2718,N_2656);
nor U2805 (N_2805,N_2786,N_2782);
nand U2806 (N_2806,N_2695,N_2666);
nand U2807 (N_2807,N_2637,N_2690);
xnor U2808 (N_2808,N_2745,N_2746);
nor U2809 (N_2809,N_2748,N_2697);
nor U2810 (N_2810,N_2723,N_2649);
nand U2811 (N_2811,N_2759,N_2667);
nand U2812 (N_2812,N_2750,N_2756);
xnor U2813 (N_2813,N_2642,N_2682);
nor U2814 (N_2814,N_2657,N_2633);
nor U2815 (N_2815,N_2626,N_2623);
xor U2816 (N_2816,N_2728,N_2770);
xor U2817 (N_2817,N_2635,N_2651);
nor U2818 (N_2818,N_2634,N_2689);
and U2819 (N_2819,N_2619,N_2778);
nand U2820 (N_2820,N_2669,N_2769);
and U2821 (N_2821,N_2730,N_2688);
nor U2822 (N_2822,N_2789,N_2740);
xnor U2823 (N_2823,N_2773,N_2654);
nor U2824 (N_2824,N_2610,N_2727);
or U2825 (N_2825,N_2641,N_2638);
nor U2826 (N_2826,N_2620,N_2713);
nand U2827 (N_2827,N_2603,N_2677);
nor U2828 (N_2828,N_2614,N_2604);
nand U2829 (N_2829,N_2643,N_2671);
xor U2830 (N_2830,N_2665,N_2679);
xnor U2831 (N_2831,N_2729,N_2771);
xor U2832 (N_2832,N_2644,N_2606);
or U2833 (N_2833,N_2650,N_2717);
nand U2834 (N_2834,N_2684,N_2777);
or U2835 (N_2835,N_2749,N_2744);
nand U2836 (N_2836,N_2758,N_2668);
xor U2837 (N_2837,N_2701,N_2658);
and U2838 (N_2838,N_2732,N_2797);
nand U2839 (N_2839,N_2780,N_2743);
or U2840 (N_2840,N_2704,N_2790);
nor U2841 (N_2841,N_2618,N_2703);
and U2842 (N_2842,N_2622,N_2757);
and U2843 (N_2843,N_2678,N_2653);
xor U2844 (N_2844,N_2673,N_2766);
nor U2845 (N_2845,N_2664,N_2764);
and U2846 (N_2846,N_2742,N_2788);
nand U2847 (N_2847,N_2632,N_2624);
nand U2848 (N_2848,N_2661,N_2726);
nor U2849 (N_2849,N_2627,N_2600);
and U2850 (N_2850,N_2692,N_2612);
or U2851 (N_2851,N_2609,N_2733);
or U2852 (N_2852,N_2663,N_2613);
nand U2853 (N_2853,N_2615,N_2629);
or U2854 (N_2854,N_2795,N_2747);
or U2855 (N_2855,N_2783,N_2720);
and U2856 (N_2856,N_2693,N_2716);
or U2857 (N_2857,N_2608,N_2779);
and U2858 (N_2858,N_2791,N_2731);
nand U2859 (N_2859,N_2696,N_2705);
and U2860 (N_2860,N_2799,N_2762);
nand U2861 (N_2861,N_2640,N_2672);
xnor U2862 (N_2862,N_2772,N_2605);
nand U2863 (N_2863,N_2784,N_2711);
nand U2864 (N_2864,N_2755,N_2694);
and U2865 (N_2865,N_2630,N_2787);
nor U2866 (N_2866,N_2700,N_2685);
nor U2867 (N_2867,N_2602,N_2683);
nor U2868 (N_2868,N_2794,N_2781);
or U2869 (N_2869,N_2774,N_2765);
nor U2870 (N_2870,N_2735,N_2681);
or U2871 (N_2871,N_2708,N_2763);
xnor U2872 (N_2872,N_2709,N_2776);
or U2873 (N_2873,N_2691,N_2686);
xor U2874 (N_2874,N_2739,N_2674);
and U2875 (N_2875,N_2734,N_2760);
nor U2876 (N_2876,N_2725,N_2645);
and U2877 (N_2877,N_2761,N_2655);
and U2878 (N_2878,N_2792,N_2660);
nand U2879 (N_2879,N_2753,N_2706);
or U2880 (N_2880,N_2798,N_2714);
nand U2881 (N_2881,N_2675,N_2767);
xnor U2882 (N_2882,N_2710,N_2616);
nor U2883 (N_2883,N_2699,N_2722);
nor U2884 (N_2884,N_2715,N_2719);
and U2885 (N_2885,N_2768,N_2737);
and U2886 (N_2886,N_2680,N_2702);
or U2887 (N_2887,N_2611,N_2636);
nand U2888 (N_2888,N_2741,N_2775);
and U2889 (N_2889,N_2621,N_2639);
nand U2890 (N_2890,N_2712,N_2707);
nor U2891 (N_2891,N_2751,N_2625);
nand U2892 (N_2892,N_2687,N_2736);
nor U2893 (N_2893,N_2670,N_2793);
and U2894 (N_2894,N_2648,N_2659);
or U2895 (N_2895,N_2617,N_2796);
nor U2896 (N_2896,N_2647,N_2754);
xor U2897 (N_2897,N_2607,N_2628);
xnor U2898 (N_2898,N_2752,N_2698);
and U2899 (N_2899,N_2724,N_2721);
xnor U2900 (N_2900,N_2761,N_2686);
xnor U2901 (N_2901,N_2715,N_2638);
nor U2902 (N_2902,N_2742,N_2669);
nor U2903 (N_2903,N_2682,N_2655);
xor U2904 (N_2904,N_2699,N_2639);
nand U2905 (N_2905,N_2718,N_2695);
or U2906 (N_2906,N_2706,N_2617);
and U2907 (N_2907,N_2791,N_2636);
and U2908 (N_2908,N_2601,N_2617);
and U2909 (N_2909,N_2672,N_2737);
xnor U2910 (N_2910,N_2653,N_2790);
nand U2911 (N_2911,N_2664,N_2792);
xnor U2912 (N_2912,N_2731,N_2661);
and U2913 (N_2913,N_2649,N_2712);
or U2914 (N_2914,N_2695,N_2697);
or U2915 (N_2915,N_2668,N_2793);
and U2916 (N_2916,N_2706,N_2672);
xor U2917 (N_2917,N_2643,N_2778);
or U2918 (N_2918,N_2678,N_2788);
and U2919 (N_2919,N_2753,N_2633);
nand U2920 (N_2920,N_2623,N_2617);
and U2921 (N_2921,N_2680,N_2771);
nor U2922 (N_2922,N_2655,N_2602);
or U2923 (N_2923,N_2778,N_2729);
xnor U2924 (N_2924,N_2678,N_2736);
or U2925 (N_2925,N_2622,N_2793);
and U2926 (N_2926,N_2612,N_2713);
or U2927 (N_2927,N_2614,N_2761);
nor U2928 (N_2928,N_2770,N_2700);
nor U2929 (N_2929,N_2722,N_2681);
nand U2930 (N_2930,N_2632,N_2772);
nand U2931 (N_2931,N_2706,N_2787);
nand U2932 (N_2932,N_2647,N_2697);
nor U2933 (N_2933,N_2620,N_2769);
xor U2934 (N_2934,N_2683,N_2779);
nor U2935 (N_2935,N_2772,N_2651);
nor U2936 (N_2936,N_2718,N_2670);
nand U2937 (N_2937,N_2764,N_2661);
nand U2938 (N_2938,N_2694,N_2726);
and U2939 (N_2939,N_2779,N_2696);
nor U2940 (N_2940,N_2799,N_2606);
or U2941 (N_2941,N_2608,N_2760);
xnor U2942 (N_2942,N_2613,N_2752);
xnor U2943 (N_2943,N_2641,N_2757);
nand U2944 (N_2944,N_2784,N_2795);
nand U2945 (N_2945,N_2780,N_2611);
or U2946 (N_2946,N_2778,N_2686);
nand U2947 (N_2947,N_2736,N_2619);
nor U2948 (N_2948,N_2694,N_2696);
nor U2949 (N_2949,N_2791,N_2703);
or U2950 (N_2950,N_2792,N_2784);
and U2951 (N_2951,N_2645,N_2734);
nor U2952 (N_2952,N_2628,N_2605);
nor U2953 (N_2953,N_2730,N_2687);
or U2954 (N_2954,N_2787,N_2767);
nand U2955 (N_2955,N_2751,N_2648);
nor U2956 (N_2956,N_2727,N_2765);
or U2957 (N_2957,N_2735,N_2632);
nor U2958 (N_2958,N_2728,N_2655);
and U2959 (N_2959,N_2682,N_2746);
nand U2960 (N_2960,N_2647,N_2725);
xor U2961 (N_2961,N_2644,N_2767);
or U2962 (N_2962,N_2761,N_2728);
nor U2963 (N_2963,N_2638,N_2698);
xnor U2964 (N_2964,N_2683,N_2747);
and U2965 (N_2965,N_2724,N_2780);
nor U2966 (N_2966,N_2603,N_2621);
xor U2967 (N_2967,N_2682,N_2630);
nor U2968 (N_2968,N_2642,N_2760);
xor U2969 (N_2969,N_2629,N_2749);
nor U2970 (N_2970,N_2677,N_2743);
and U2971 (N_2971,N_2646,N_2639);
nor U2972 (N_2972,N_2655,N_2722);
nand U2973 (N_2973,N_2604,N_2615);
xnor U2974 (N_2974,N_2683,N_2739);
xor U2975 (N_2975,N_2656,N_2634);
xnor U2976 (N_2976,N_2735,N_2614);
xnor U2977 (N_2977,N_2728,N_2733);
nor U2978 (N_2978,N_2611,N_2627);
and U2979 (N_2979,N_2612,N_2716);
nand U2980 (N_2980,N_2738,N_2625);
and U2981 (N_2981,N_2716,N_2655);
nor U2982 (N_2982,N_2655,N_2648);
nor U2983 (N_2983,N_2610,N_2666);
and U2984 (N_2984,N_2701,N_2686);
or U2985 (N_2985,N_2680,N_2693);
and U2986 (N_2986,N_2608,N_2747);
or U2987 (N_2987,N_2729,N_2739);
nor U2988 (N_2988,N_2666,N_2659);
or U2989 (N_2989,N_2657,N_2687);
xnor U2990 (N_2990,N_2777,N_2778);
nand U2991 (N_2991,N_2627,N_2749);
or U2992 (N_2992,N_2687,N_2659);
and U2993 (N_2993,N_2606,N_2642);
xor U2994 (N_2994,N_2624,N_2681);
xor U2995 (N_2995,N_2741,N_2601);
xor U2996 (N_2996,N_2725,N_2631);
nor U2997 (N_2997,N_2732,N_2714);
xnor U2998 (N_2998,N_2636,N_2661);
and U2999 (N_2999,N_2609,N_2688);
nand U3000 (N_3000,N_2928,N_2936);
nor U3001 (N_3001,N_2893,N_2950);
nor U3002 (N_3002,N_2981,N_2926);
nor U3003 (N_3003,N_2863,N_2998);
nor U3004 (N_3004,N_2839,N_2959);
or U3005 (N_3005,N_2967,N_2983);
nand U3006 (N_3006,N_2917,N_2963);
xor U3007 (N_3007,N_2804,N_2809);
nand U3008 (N_3008,N_2855,N_2988);
nor U3009 (N_3009,N_2901,N_2817);
and U3010 (N_3010,N_2908,N_2831);
xor U3011 (N_3011,N_2826,N_2848);
and U3012 (N_3012,N_2896,N_2820);
nor U3013 (N_3013,N_2949,N_2915);
xor U3014 (N_3014,N_2866,N_2997);
or U3015 (N_3015,N_2887,N_2843);
xnor U3016 (N_3016,N_2904,N_2822);
xor U3017 (N_3017,N_2937,N_2869);
xor U3018 (N_3018,N_2911,N_2986);
or U3019 (N_3019,N_2883,N_2847);
xor U3020 (N_3020,N_2953,N_2973);
nand U3021 (N_3021,N_2801,N_2881);
nor U3022 (N_3022,N_2990,N_2941);
nor U3023 (N_3023,N_2871,N_2832);
xnor U3024 (N_3024,N_2955,N_2849);
and U3025 (N_3025,N_2920,N_2823);
xor U3026 (N_3026,N_2877,N_2886);
and U3027 (N_3027,N_2902,N_2929);
xnor U3028 (N_3028,N_2912,N_2961);
nand U3029 (N_3029,N_2837,N_2840);
xnor U3030 (N_3030,N_2897,N_2982);
xor U3031 (N_3031,N_2819,N_2977);
and U3032 (N_3032,N_2878,N_2813);
and U3033 (N_3033,N_2800,N_2931);
nand U3034 (N_3034,N_2939,N_2900);
xor U3035 (N_3035,N_2923,N_2924);
nor U3036 (N_3036,N_2879,N_2960);
nor U3037 (N_3037,N_2815,N_2838);
nand U3038 (N_3038,N_2818,N_2814);
xnor U3039 (N_3039,N_2962,N_2864);
nor U3040 (N_3040,N_2940,N_2805);
and U3041 (N_3041,N_2991,N_2892);
or U3042 (N_3042,N_2907,N_2957);
or U3043 (N_3043,N_2899,N_2905);
and U3044 (N_3044,N_2968,N_2859);
nand U3045 (N_3045,N_2946,N_2942);
nor U3046 (N_3046,N_2860,N_2965);
and U3047 (N_3047,N_2857,N_2974);
or U3048 (N_3048,N_2827,N_2874);
nor U3049 (N_3049,N_2922,N_2943);
nand U3050 (N_3050,N_2807,N_2992);
xnor U3051 (N_3051,N_2803,N_2811);
nand U3052 (N_3052,N_2952,N_2964);
and U3053 (N_3053,N_2858,N_2845);
or U3054 (N_3054,N_2872,N_2828);
or U3055 (N_3055,N_2970,N_2945);
or U3056 (N_3056,N_2966,N_2935);
or U3057 (N_3057,N_2850,N_2889);
xnor U3058 (N_3058,N_2898,N_2993);
nor U3059 (N_3059,N_2994,N_2853);
xnor U3060 (N_3060,N_2979,N_2999);
and U3061 (N_3061,N_2851,N_2916);
and U3062 (N_3062,N_2969,N_2852);
or U3063 (N_3063,N_2958,N_2895);
nand U3064 (N_3064,N_2802,N_2972);
nand U3065 (N_3065,N_2821,N_2885);
xor U3066 (N_3066,N_2861,N_2989);
xor U3067 (N_3067,N_2862,N_2996);
or U3068 (N_3068,N_2875,N_2906);
nand U3069 (N_3069,N_2956,N_2867);
nand U3070 (N_3070,N_2835,N_2921);
and U3071 (N_3071,N_2980,N_2919);
or U3072 (N_3072,N_2825,N_2985);
xnor U3073 (N_3073,N_2913,N_2951);
nand U3074 (N_3074,N_2903,N_2918);
nand U3075 (N_3075,N_2933,N_2865);
xnor U3076 (N_3076,N_2909,N_2870);
nand U3077 (N_3077,N_2995,N_2925);
or U3078 (N_3078,N_2944,N_2934);
xor U3079 (N_3079,N_2868,N_2971);
or U3080 (N_3080,N_2856,N_2938);
or U3081 (N_3081,N_2842,N_2954);
and U3082 (N_3082,N_2884,N_2890);
nand U3083 (N_3083,N_2836,N_2978);
and U3084 (N_3084,N_2829,N_2833);
or U3085 (N_3085,N_2806,N_2930);
and U3086 (N_3086,N_2987,N_2846);
xor U3087 (N_3087,N_2854,N_2876);
or U3088 (N_3088,N_2844,N_2824);
xor U3089 (N_3089,N_2891,N_2834);
nor U3090 (N_3090,N_2888,N_2873);
xnor U3091 (N_3091,N_2947,N_2910);
xor U3092 (N_3092,N_2816,N_2812);
nor U3093 (N_3093,N_2948,N_2810);
or U3094 (N_3094,N_2976,N_2932);
and U3095 (N_3095,N_2975,N_2914);
xnor U3096 (N_3096,N_2927,N_2880);
and U3097 (N_3097,N_2808,N_2830);
or U3098 (N_3098,N_2984,N_2841);
or U3099 (N_3099,N_2894,N_2882);
or U3100 (N_3100,N_2846,N_2959);
nor U3101 (N_3101,N_2912,N_2875);
nand U3102 (N_3102,N_2946,N_2871);
and U3103 (N_3103,N_2942,N_2808);
or U3104 (N_3104,N_2874,N_2956);
xnor U3105 (N_3105,N_2909,N_2990);
xnor U3106 (N_3106,N_2827,N_2922);
and U3107 (N_3107,N_2921,N_2825);
and U3108 (N_3108,N_2842,N_2864);
nor U3109 (N_3109,N_2948,N_2854);
or U3110 (N_3110,N_2816,N_2891);
nor U3111 (N_3111,N_2979,N_2892);
and U3112 (N_3112,N_2955,N_2900);
and U3113 (N_3113,N_2988,N_2920);
xnor U3114 (N_3114,N_2926,N_2895);
nand U3115 (N_3115,N_2990,N_2868);
or U3116 (N_3116,N_2869,N_2803);
xnor U3117 (N_3117,N_2831,N_2954);
or U3118 (N_3118,N_2891,N_2999);
nor U3119 (N_3119,N_2903,N_2902);
and U3120 (N_3120,N_2902,N_2841);
or U3121 (N_3121,N_2827,N_2889);
xnor U3122 (N_3122,N_2888,N_2945);
nor U3123 (N_3123,N_2927,N_2827);
or U3124 (N_3124,N_2851,N_2824);
or U3125 (N_3125,N_2903,N_2977);
or U3126 (N_3126,N_2961,N_2939);
or U3127 (N_3127,N_2937,N_2876);
or U3128 (N_3128,N_2830,N_2996);
nor U3129 (N_3129,N_2999,N_2993);
xor U3130 (N_3130,N_2968,N_2893);
nor U3131 (N_3131,N_2868,N_2950);
or U3132 (N_3132,N_2996,N_2815);
nor U3133 (N_3133,N_2826,N_2832);
nor U3134 (N_3134,N_2953,N_2820);
or U3135 (N_3135,N_2859,N_2971);
and U3136 (N_3136,N_2947,N_2852);
or U3137 (N_3137,N_2975,N_2895);
nor U3138 (N_3138,N_2894,N_2872);
or U3139 (N_3139,N_2815,N_2895);
nor U3140 (N_3140,N_2833,N_2893);
nand U3141 (N_3141,N_2952,N_2925);
and U3142 (N_3142,N_2948,N_2885);
nor U3143 (N_3143,N_2813,N_2843);
or U3144 (N_3144,N_2900,N_2934);
nor U3145 (N_3145,N_2835,N_2917);
nand U3146 (N_3146,N_2965,N_2934);
nor U3147 (N_3147,N_2923,N_2893);
xnor U3148 (N_3148,N_2852,N_2972);
nand U3149 (N_3149,N_2991,N_2839);
or U3150 (N_3150,N_2935,N_2893);
nor U3151 (N_3151,N_2826,N_2925);
or U3152 (N_3152,N_2890,N_2905);
nor U3153 (N_3153,N_2957,N_2983);
and U3154 (N_3154,N_2919,N_2959);
nor U3155 (N_3155,N_2893,N_2825);
nor U3156 (N_3156,N_2934,N_2882);
or U3157 (N_3157,N_2874,N_2962);
xor U3158 (N_3158,N_2867,N_2986);
and U3159 (N_3159,N_2845,N_2883);
nand U3160 (N_3160,N_2925,N_2905);
or U3161 (N_3161,N_2937,N_2885);
and U3162 (N_3162,N_2898,N_2897);
nand U3163 (N_3163,N_2932,N_2928);
xor U3164 (N_3164,N_2894,N_2949);
xnor U3165 (N_3165,N_2976,N_2853);
xnor U3166 (N_3166,N_2859,N_2977);
nand U3167 (N_3167,N_2981,N_2912);
nand U3168 (N_3168,N_2824,N_2836);
or U3169 (N_3169,N_2993,N_2946);
xnor U3170 (N_3170,N_2852,N_2992);
or U3171 (N_3171,N_2912,N_2913);
nor U3172 (N_3172,N_2926,N_2940);
nor U3173 (N_3173,N_2942,N_2884);
and U3174 (N_3174,N_2930,N_2941);
and U3175 (N_3175,N_2909,N_2837);
or U3176 (N_3176,N_2870,N_2872);
nor U3177 (N_3177,N_2955,N_2984);
or U3178 (N_3178,N_2942,N_2931);
nor U3179 (N_3179,N_2848,N_2834);
nor U3180 (N_3180,N_2931,N_2939);
nor U3181 (N_3181,N_2866,N_2905);
xor U3182 (N_3182,N_2844,N_2890);
nand U3183 (N_3183,N_2899,N_2989);
and U3184 (N_3184,N_2884,N_2866);
xnor U3185 (N_3185,N_2842,N_2859);
xor U3186 (N_3186,N_2851,N_2892);
xor U3187 (N_3187,N_2991,N_2832);
and U3188 (N_3188,N_2977,N_2929);
and U3189 (N_3189,N_2884,N_2886);
nand U3190 (N_3190,N_2993,N_2860);
and U3191 (N_3191,N_2911,N_2839);
nor U3192 (N_3192,N_2889,N_2996);
nor U3193 (N_3193,N_2934,N_2820);
nor U3194 (N_3194,N_2964,N_2859);
xnor U3195 (N_3195,N_2995,N_2979);
or U3196 (N_3196,N_2982,N_2934);
nand U3197 (N_3197,N_2929,N_2894);
or U3198 (N_3198,N_2825,N_2850);
nor U3199 (N_3199,N_2918,N_2882);
and U3200 (N_3200,N_3032,N_3121);
nand U3201 (N_3201,N_3075,N_3153);
nor U3202 (N_3202,N_3004,N_3174);
xor U3203 (N_3203,N_3160,N_3193);
and U3204 (N_3204,N_3099,N_3014);
xnor U3205 (N_3205,N_3183,N_3085);
nand U3206 (N_3206,N_3078,N_3176);
or U3207 (N_3207,N_3198,N_3158);
xnor U3208 (N_3208,N_3175,N_3053);
xor U3209 (N_3209,N_3019,N_3043);
nor U3210 (N_3210,N_3033,N_3129);
or U3211 (N_3211,N_3161,N_3050);
or U3212 (N_3212,N_3197,N_3196);
or U3213 (N_3213,N_3144,N_3170);
nor U3214 (N_3214,N_3165,N_3127);
or U3215 (N_3215,N_3178,N_3172);
nor U3216 (N_3216,N_3061,N_3066);
and U3217 (N_3217,N_3086,N_3022);
or U3218 (N_3218,N_3133,N_3159);
nand U3219 (N_3219,N_3194,N_3115);
nor U3220 (N_3220,N_3134,N_3108);
nor U3221 (N_3221,N_3013,N_3171);
xor U3222 (N_3222,N_3017,N_3025);
nand U3223 (N_3223,N_3179,N_3168);
nor U3224 (N_3224,N_3040,N_3024);
nand U3225 (N_3225,N_3111,N_3096);
xnor U3226 (N_3226,N_3021,N_3109);
and U3227 (N_3227,N_3138,N_3152);
or U3228 (N_3228,N_3114,N_3047);
and U3229 (N_3229,N_3026,N_3195);
nor U3230 (N_3230,N_3154,N_3052);
or U3231 (N_3231,N_3180,N_3141);
nand U3232 (N_3232,N_3039,N_3177);
and U3233 (N_3233,N_3199,N_3117);
and U3234 (N_3234,N_3136,N_3166);
xnor U3235 (N_3235,N_3035,N_3103);
and U3236 (N_3236,N_3132,N_3023);
nor U3237 (N_3237,N_3167,N_3130);
and U3238 (N_3238,N_3087,N_3045);
nand U3239 (N_3239,N_3143,N_3191);
and U3240 (N_3240,N_3092,N_3020);
xnor U3241 (N_3241,N_3034,N_3037);
xor U3242 (N_3242,N_3018,N_3041);
nand U3243 (N_3243,N_3173,N_3006);
nor U3244 (N_3244,N_3122,N_3135);
or U3245 (N_3245,N_3084,N_3169);
and U3246 (N_3246,N_3104,N_3003);
nor U3247 (N_3247,N_3031,N_3091);
or U3248 (N_3248,N_3123,N_3067);
nor U3249 (N_3249,N_3089,N_3106);
xnor U3250 (N_3250,N_3151,N_3070);
and U3251 (N_3251,N_3181,N_3016);
or U3252 (N_3252,N_3137,N_3128);
nor U3253 (N_3253,N_3057,N_3101);
nand U3254 (N_3254,N_3028,N_3188);
and U3255 (N_3255,N_3190,N_3098);
or U3256 (N_3256,N_3094,N_3063);
xnor U3257 (N_3257,N_3119,N_3097);
nand U3258 (N_3258,N_3008,N_3069);
xor U3259 (N_3259,N_3120,N_3146);
nand U3260 (N_3260,N_3163,N_3187);
xor U3261 (N_3261,N_3015,N_3142);
nor U3262 (N_3262,N_3083,N_3048);
nand U3263 (N_3263,N_3095,N_3077);
or U3264 (N_3264,N_3079,N_3002);
nand U3265 (N_3265,N_3059,N_3071);
or U3266 (N_3266,N_3124,N_3001);
xor U3267 (N_3267,N_3065,N_3007);
and U3268 (N_3268,N_3185,N_3005);
and U3269 (N_3269,N_3076,N_3062);
nor U3270 (N_3270,N_3036,N_3147);
and U3271 (N_3271,N_3182,N_3010);
or U3272 (N_3272,N_3030,N_3046);
and U3273 (N_3273,N_3038,N_3110);
nand U3274 (N_3274,N_3060,N_3054);
or U3275 (N_3275,N_3162,N_3150);
or U3276 (N_3276,N_3157,N_3029);
nand U3277 (N_3277,N_3100,N_3042);
and U3278 (N_3278,N_3105,N_3189);
and U3279 (N_3279,N_3051,N_3072);
nor U3280 (N_3280,N_3080,N_3184);
nor U3281 (N_3281,N_3068,N_3156);
nand U3282 (N_3282,N_3140,N_3145);
or U3283 (N_3283,N_3139,N_3125);
nor U3284 (N_3284,N_3148,N_3107);
xor U3285 (N_3285,N_3000,N_3073);
and U3286 (N_3286,N_3102,N_3164);
or U3287 (N_3287,N_3044,N_3064);
nor U3288 (N_3288,N_3088,N_3192);
or U3289 (N_3289,N_3093,N_3113);
and U3290 (N_3290,N_3118,N_3012);
and U3291 (N_3291,N_3149,N_3056);
nor U3292 (N_3292,N_3081,N_3126);
nand U3293 (N_3293,N_3049,N_3112);
or U3294 (N_3294,N_3011,N_3131);
nor U3295 (N_3295,N_3082,N_3186);
xor U3296 (N_3296,N_3009,N_3116);
nor U3297 (N_3297,N_3055,N_3027);
and U3298 (N_3298,N_3058,N_3090);
and U3299 (N_3299,N_3155,N_3074);
nand U3300 (N_3300,N_3103,N_3131);
and U3301 (N_3301,N_3040,N_3095);
nor U3302 (N_3302,N_3130,N_3195);
nor U3303 (N_3303,N_3184,N_3004);
xor U3304 (N_3304,N_3105,N_3003);
nor U3305 (N_3305,N_3112,N_3098);
nand U3306 (N_3306,N_3124,N_3071);
nor U3307 (N_3307,N_3069,N_3198);
or U3308 (N_3308,N_3145,N_3062);
or U3309 (N_3309,N_3060,N_3061);
nand U3310 (N_3310,N_3177,N_3110);
nor U3311 (N_3311,N_3177,N_3151);
nor U3312 (N_3312,N_3197,N_3185);
xor U3313 (N_3313,N_3074,N_3101);
nor U3314 (N_3314,N_3046,N_3002);
or U3315 (N_3315,N_3108,N_3115);
xnor U3316 (N_3316,N_3037,N_3195);
and U3317 (N_3317,N_3154,N_3033);
xnor U3318 (N_3318,N_3182,N_3092);
xor U3319 (N_3319,N_3166,N_3090);
nand U3320 (N_3320,N_3090,N_3085);
nand U3321 (N_3321,N_3129,N_3108);
and U3322 (N_3322,N_3000,N_3026);
nor U3323 (N_3323,N_3170,N_3094);
xnor U3324 (N_3324,N_3054,N_3088);
or U3325 (N_3325,N_3043,N_3013);
nand U3326 (N_3326,N_3140,N_3166);
or U3327 (N_3327,N_3025,N_3190);
nor U3328 (N_3328,N_3140,N_3079);
nand U3329 (N_3329,N_3093,N_3057);
or U3330 (N_3330,N_3058,N_3019);
or U3331 (N_3331,N_3071,N_3185);
nor U3332 (N_3332,N_3159,N_3079);
and U3333 (N_3333,N_3033,N_3182);
or U3334 (N_3334,N_3129,N_3043);
nor U3335 (N_3335,N_3135,N_3164);
nand U3336 (N_3336,N_3131,N_3186);
and U3337 (N_3337,N_3098,N_3142);
xor U3338 (N_3338,N_3070,N_3107);
or U3339 (N_3339,N_3077,N_3061);
and U3340 (N_3340,N_3059,N_3082);
xor U3341 (N_3341,N_3020,N_3183);
and U3342 (N_3342,N_3023,N_3194);
nor U3343 (N_3343,N_3013,N_3140);
nor U3344 (N_3344,N_3014,N_3140);
nor U3345 (N_3345,N_3029,N_3102);
xnor U3346 (N_3346,N_3122,N_3127);
or U3347 (N_3347,N_3062,N_3121);
and U3348 (N_3348,N_3001,N_3041);
nor U3349 (N_3349,N_3105,N_3085);
and U3350 (N_3350,N_3149,N_3150);
xnor U3351 (N_3351,N_3177,N_3161);
nor U3352 (N_3352,N_3035,N_3040);
nor U3353 (N_3353,N_3118,N_3015);
and U3354 (N_3354,N_3133,N_3148);
or U3355 (N_3355,N_3092,N_3105);
or U3356 (N_3356,N_3137,N_3036);
and U3357 (N_3357,N_3011,N_3054);
or U3358 (N_3358,N_3166,N_3027);
and U3359 (N_3359,N_3049,N_3145);
nor U3360 (N_3360,N_3106,N_3134);
and U3361 (N_3361,N_3018,N_3062);
and U3362 (N_3362,N_3076,N_3174);
nand U3363 (N_3363,N_3175,N_3052);
and U3364 (N_3364,N_3088,N_3160);
nor U3365 (N_3365,N_3041,N_3085);
and U3366 (N_3366,N_3085,N_3143);
or U3367 (N_3367,N_3015,N_3080);
nand U3368 (N_3368,N_3156,N_3136);
nor U3369 (N_3369,N_3023,N_3035);
nor U3370 (N_3370,N_3092,N_3111);
or U3371 (N_3371,N_3066,N_3174);
or U3372 (N_3372,N_3100,N_3075);
xor U3373 (N_3373,N_3153,N_3000);
nand U3374 (N_3374,N_3132,N_3024);
and U3375 (N_3375,N_3138,N_3039);
or U3376 (N_3376,N_3074,N_3113);
or U3377 (N_3377,N_3174,N_3050);
xor U3378 (N_3378,N_3010,N_3116);
nand U3379 (N_3379,N_3020,N_3058);
nor U3380 (N_3380,N_3095,N_3131);
nand U3381 (N_3381,N_3141,N_3132);
nor U3382 (N_3382,N_3129,N_3127);
and U3383 (N_3383,N_3046,N_3182);
nand U3384 (N_3384,N_3076,N_3065);
xnor U3385 (N_3385,N_3134,N_3017);
or U3386 (N_3386,N_3172,N_3190);
xor U3387 (N_3387,N_3094,N_3071);
nand U3388 (N_3388,N_3097,N_3007);
and U3389 (N_3389,N_3144,N_3063);
nand U3390 (N_3390,N_3123,N_3137);
or U3391 (N_3391,N_3142,N_3150);
nand U3392 (N_3392,N_3076,N_3129);
nand U3393 (N_3393,N_3141,N_3070);
or U3394 (N_3394,N_3099,N_3114);
nand U3395 (N_3395,N_3115,N_3098);
xor U3396 (N_3396,N_3128,N_3086);
or U3397 (N_3397,N_3013,N_3121);
nor U3398 (N_3398,N_3165,N_3171);
nor U3399 (N_3399,N_3103,N_3189);
and U3400 (N_3400,N_3259,N_3328);
nor U3401 (N_3401,N_3201,N_3223);
and U3402 (N_3402,N_3204,N_3233);
xor U3403 (N_3403,N_3388,N_3254);
or U3404 (N_3404,N_3271,N_3247);
nand U3405 (N_3405,N_3322,N_3319);
and U3406 (N_3406,N_3318,N_3206);
xnor U3407 (N_3407,N_3297,N_3225);
nand U3408 (N_3408,N_3220,N_3250);
or U3409 (N_3409,N_3324,N_3380);
and U3410 (N_3410,N_3272,N_3392);
nor U3411 (N_3411,N_3292,N_3373);
nand U3412 (N_3412,N_3384,N_3228);
nor U3413 (N_3413,N_3245,N_3365);
and U3414 (N_3414,N_3263,N_3231);
or U3415 (N_3415,N_3289,N_3266);
xor U3416 (N_3416,N_3218,N_3371);
or U3417 (N_3417,N_3200,N_3309);
nand U3418 (N_3418,N_3213,N_3284);
nand U3419 (N_3419,N_3312,N_3367);
xor U3420 (N_3420,N_3255,N_3298);
xor U3421 (N_3421,N_3379,N_3376);
or U3422 (N_3422,N_3336,N_3208);
xnor U3423 (N_3423,N_3258,N_3333);
and U3424 (N_3424,N_3214,N_3252);
nor U3425 (N_3425,N_3342,N_3345);
and U3426 (N_3426,N_3275,N_3381);
and U3427 (N_3427,N_3207,N_3224);
xor U3428 (N_3428,N_3209,N_3375);
xor U3429 (N_3429,N_3279,N_3339);
or U3430 (N_3430,N_3317,N_3326);
xor U3431 (N_3431,N_3248,N_3349);
nor U3432 (N_3432,N_3321,N_3203);
nor U3433 (N_3433,N_3305,N_3205);
xor U3434 (N_3434,N_3315,N_3308);
or U3435 (N_3435,N_3210,N_3390);
nand U3436 (N_3436,N_3249,N_3219);
nand U3437 (N_3437,N_3285,N_3242);
xnor U3438 (N_3438,N_3368,N_3341);
nor U3439 (N_3439,N_3230,N_3359);
nand U3440 (N_3440,N_3378,N_3391);
nor U3441 (N_3441,N_3399,N_3251);
nand U3442 (N_3442,N_3240,N_3291);
and U3443 (N_3443,N_3356,N_3314);
and U3444 (N_3444,N_3243,N_3229);
xnor U3445 (N_3445,N_3282,N_3277);
nor U3446 (N_3446,N_3307,N_3236);
xor U3447 (N_3447,N_3262,N_3238);
nand U3448 (N_3448,N_3395,N_3267);
nand U3449 (N_3449,N_3363,N_3302);
nor U3450 (N_3450,N_3222,N_3329);
xor U3451 (N_3451,N_3348,N_3202);
and U3452 (N_3452,N_3288,N_3332);
xnor U3453 (N_3453,N_3234,N_3389);
or U3454 (N_3454,N_3337,N_3352);
nand U3455 (N_3455,N_3331,N_3360);
xnor U3456 (N_3456,N_3343,N_3320);
nor U3457 (N_3457,N_3217,N_3265);
xnor U3458 (N_3458,N_3276,N_3301);
nand U3459 (N_3459,N_3283,N_3215);
or U3460 (N_3460,N_3344,N_3280);
and U3461 (N_3461,N_3237,N_3323);
and U3462 (N_3462,N_3299,N_3216);
xor U3463 (N_3463,N_3221,N_3346);
nand U3464 (N_3464,N_3294,N_3244);
xnor U3465 (N_3465,N_3261,N_3246);
nand U3466 (N_3466,N_3287,N_3311);
or U3467 (N_3467,N_3316,N_3327);
xor U3468 (N_3468,N_3382,N_3330);
or U3469 (N_3469,N_3286,N_3269);
nor U3470 (N_3470,N_3232,N_3334);
xor U3471 (N_3471,N_3295,N_3370);
and U3472 (N_3472,N_3303,N_3354);
xnor U3473 (N_3473,N_3335,N_3353);
xor U3474 (N_3474,N_3385,N_3227);
nor U3475 (N_3475,N_3351,N_3383);
nand U3476 (N_3476,N_3257,N_3355);
or U3477 (N_3477,N_3274,N_3212);
nand U3478 (N_3478,N_3369,N_3296);
or U3479 (N_3479,N_3226,N_3304);
nor U3480 (N_3480,N_3347,N_3270);
nand U3481 (N_3481,N_3393,N_3387);
xnor U3482 (N_3482,N_3361,N_3397);
or U3483 (N_3483,N_3372,N_3256);
nand U3484 (N_3484,N_3362,N_3357);
or U3485 (N_3485,N_3264,N_3310);
nand U3486 (N_3486,N_3313,N_3300);
xor U3487 (N_3487,N_3374,N_3235);
xor U3488 (N_3488,N_3396,N_3350);
or U3489 (N_3489,N_3293,N_3325);
or U3490 (N_3490,N_3241,N_3306);
and U3491 (N_3491,N_3290,N_3268);
and U3492 (N_3492,N_3398,N_3366);
nand U3493 (N_3493,N_3278,N_3281);
nor U3494 (N_3494,N_3364,N_3358);
and U3495 (N_3495,N_3273,N_3253);
or U3496 (N_3496,N_3211,N_3394);
and U3497 (N_3497,N_3239,N_3377);
nand U3498 (N_3498,N_3338,N_3260);
nand U3499 (N_3499,N_3386,N_3340);
xnor U3500 (N_3500,N_3251,N_3253);
or U3501 (N_3501,N_3356,N_3334);
xor U3502 (N_3502,N_3246,N_3204);
nor U3503 (N_3503,N_3232,N_3276);
and U3504 (N_3504,N_3317,N_3322);
nand U3505 (N_3505,N_3232,N_3216);
or U3506 (N_3506,N_3221,N_3386);
nor U3507 (N_3507,N_3381,N_3204);
nor U3508 (N_3508,N_3380,N_3275);
xnor U3509 (N_3509,N_3227,N_3352);
and U3510 (N_3510,N_3360,N_3217);
nand U3511 (N_3511,N_3292,N_3270);
xnor U3512 (N_3512,N_3321,N_3207);
nand U3513 (N_3513,N_3355,N_3363);
nand U3514 (N_3514,N_3232,N_3230);
nor U3515 (N_3515,N_3389,N_3284);
nand U3516 (N_3516,N_3363,N_3306);
nor U3517 (N_3517,N_3272,N_3304);
nand U3518 (N_3518,N_3276,N_3302);
or U3519 (N_3519,N_3398,N_3307);
and U3520 (N_3520,N_3314,N_3381);
or U3521 (N_3521,N_3275,N_3347);
or U3522 (N_3522,N_3329,N_3203);
nand U3523 (N_3523,N_3226,N_3391);
xor U3524 (N_3524,N_3305,N_3243);
and U3525 (N_3525,N_3393,N_3288);
nor U3526 (N_3526,N_3257,N_3241);
xor U3527 (N_3527,N_3220,N_3218);
or U3528 (N_3528,N_3287,N_3205);
xnor U3529 (N_3529,N_3286,N_3264);
and U3530 (N_3530,N_3300,N_3377);
xnor U3531 (N_3531,N_3280,N_3358);
xnor U3532 (N_3532,N_3362,N_3306);
xor U3533 (N_3533,N_3201,N_3379);
and U3534 (N_3534,N_3307,N_3293);
and U3535 (N_3535,N_3357,N_3220);
or U3536 (N_3536,N_3396,N_3263);
and U3537 (N_3537,N_3386,N_3277);
xor U3538 (N_3538,N_3219,N_3230);
nor U3539 (N_3539,N_3300,N_3306);
nand U3540 (N_3540,N_3219,N_3335);
xnor U3541 (N_3541,N_3247,N_3234);
or U3542 (N_3542,N_3347,N_3385);
nor U3543 (N_3543,N_3398,N_3255);
and U3544 (N_3544,N_3286,N_3381);
or U3545 (N_3545,N_3297,N_3230);
nand U3546 (N_3546,N_3318,N_3225);
xnor U3547 (N_3547,N_3309,N_3385);
xor U3548 (N_3548,N_3217,N_3297);
nor U3549 (N_3549,N_3339,N_3387);
or U3550 (N_3550,N_3208,N_3203);
or U3551 (N_3551,N_3278,N_3231);
or U3552 (N_3552,N_3383,N_3311);
xnor U3553 (N_3553,N_3303,N_3231);
xor U3554 (N_3554,N_3355,N_3331);
nor U3555 (N_3555,N_3317,N_3341);
and U3556 (N_3556,N_3222,N_3356);
nand U3557 (N_3557,N_3300,N_3378);
xor U3558 (N_3558,N_3223,N_3358);
nor U3559 (N_3559,N_3272,N_3238);
nor U3560 (N_3560,N_3313,N_3240);
xor U3561 (N_3561,N_3321,N_3293);
nor U3562 (N_3562,N_3355,N_3273);
or U3563 (N_3563,N_3246,N_3304);
or U3564 (N_3564,N_3362,N_3325);
xor U3565 (N_3565,N_3330,N_3362);
or U3566 (N_3566,N_3205,N_3394);
nand U3567 (N_3567,N_3209,N_3243);
and U3568 (N_3568,N_3316,N_3312);
nand U3569 (N_3569,N_3385,N_3265);
or U3570 (N_3570,N_3268,N_3383);
or U3571 (N_3571,N_3269,N_3276);
nand U3572 (N_3572,N_3309,N_3210);
and U3573 (N_3573,N_3204,N_3276);
or U3574 (N_3574,N_3204,N_3327);
nor U3575 (N_3575,N_3337,N_3321);
nand U3576 (N_3576,N_3298,N_3289);
or U3577 (N_3577,N_3215,N_3356);
or U3578 (N_3578,N_3337,N_3361);
xor U3579 (N_3579,N_3280,N_3200);
nand U3580 (N_3580,N_3312,N_3215);
or U3581 (N_3581,N_3206,N_3202);
xor U3582 (N_3582,N_3270,N_3253);
nor U3583 (N_3583,N_3348,N_3246);
nand U3584 (N_3584,N_3396,N_3287);
and U3585 (N_3585,N_3254,N_3256);
or U3586 (N_3586,N_3244,N_3367);
nand U3587 (N_3587,N_3265,N_3290);
xnor U3588 (N_3588,N_3298,N_3310);
nor U3589 (N_3589,N_3205,N_3254);
xor U3590 (N_3590,N_3358,N_3227);
xnor U3591 (N_3591,N_3209,N_3306);
or U3592 (N_3592,N_3375,N_3265);
xnor U3593 (N_3593,N_3232,N_3223);
or U3594 (N_3594,N_3309,N_3330);
nand U3595 (N_3595,N_3264,N_3241);
xor U3596 (N_3596,N_3311,N_3230);
and U3597 (N_3597,N_3391,N_3302);
nor U3598 (N_3598,N_3268,N_3328);
nor U3599 (N_3599,N_3288,N_3230);
or U3600 (N_3600,N_3419,N_3493);
xnor U3601 (N_3601,N_3583,N_3438);
and U3602 (N_3602,N_3514,N_3418);
or U3603 (N_3603,N_3406,N_3451);
or U3604 (N_3604,N_3504,N_3554);
xor U3605 (N_3605,N_3586,N_3528);
or U3606 (N_3606,N_3549,N_3596);
xnor U3607 (N_3607,N_3575,N_3413);
or U3608 (N_3608,N_3574,N_3559);
nand U3609 (N_3609,N_3436,N_3466);
nand U3610 (N_3610,N_3547,N_3478);
or U3611 (N_3611,N_3459,N_3538);
xor U3612 (N_3612,N_3472,N_3485);
or U3613 (N_3613,N_3446,N_3563);
or U3614 (N_3614,N_3512,N_3543);
nor U3615 (N_3615,N_3507,N_3524);
xor U3616 (N_3616,N_3502,N_3428);
nand U3617 (N_3617,N_3498,N_3531);
and U3618 (N_3618,N_3542,N_3598);
and U3619 (N_3619,N_3470,N_3500);
and U3620 (N_3620,N_3577,N_3407);
or U3621 (N_3621,N_3537,N_3469);
xor U3622 (N_3622,N_3536,N_3511);
nand U3623 (N_3623,N_3440,N_3402);
or U3624 (N_3624,N_3488,N_3495);
nand U3625 (N_3625,N_3425,N_3517);
or U3626 (N_3626,N_3423,N_3473);
nand U3627 (N_3627,N_3442,N_3494);
xor U3628 (N_3628,N_3471,N_3565);
nor U3629 (N_3629,N_3429,N_3403);
nor U3630 (N_3630,N_3573,N_3439);
nand U3631 (N_3631,N_3427,N_3450);
or U3632 (N_3632,N_3441,N_3580);
nor U3633 (N_3633,N_3545,N_3550);
nor U3634 (N_3634,N_3530,N_3465);
and U3635 (N_3635,N_3510,N_3490);
nor U3636 (N_3636,N_3467,N_3477);
xor U3637 (N_3637,N_3454,N_3457);
or U3638 (N_3638,N_3408,N_3509);
xnor U3639 (N_3639,N_3569,N_3434);
nor U3640 (N_3640,N_3597,N_3489);
and U3641 (N_3641,N_3560,N_3513);
or U3642 (N_3642,N_3404,N_3480);
or U3643 (N_3643,N_3525,N_3458);
nand U3644 (N_3644,N_3519,N_3435);
xor U3645 (N_3645,N_3593,N_3420);
nand U3646 (N_3646,N_3595,N_3572);
xor U3647 (N_3647,N_3579,N_3400);
and U3648 (N_3648,N_3452,N_3431);
nand U3649 (N_3649,N_3557,N_3476);
nor U3650 (N_3650,N_3437,N_3540);
nor U3651 (N_3651,N_3468,N_3496);
xnor U3652 (N_3652,N_3492,N_3430);
nand U3653 (N_3653,N_3416,N_3412);
nor U3654 (N_3654,N_3456,N_3571);
or U3655 (N_3655,N_3432,N_3567);
xor U3656 (N_3656,N_3516,N_3591);
or U3657 (N_3657,N_3523,N_3405);
nand U3658 (N_3658,N_3534,N_3551);
nor U3659 (N_3659,N_3558,N_3535);
or U3660 (N_3660,N_3556,N_3529);
or U3661 (N_3661,N_3564,N_3422);
or U3662 (N_3662,N_3548,N_3479);
and U3663 (N_3663,N_3594,N_3462);
or U3664 (N_3664,N_3444,N_3409);
and U3665 (N_3665,N_3464,N_3562);
nor U3666 (N_3666,N_3590,N_3463);
xor U3667 (N_3667,N_3526,N_3426);
nor U3668 (N_3668,N_3508,N_3578);
or U3669 (N_3669,N_3497,N_3455);
and U3670 (N_3670,N_3566,N_3448);
or U3671 (N_3671,N_3414,N_3453);
xor U3672 (N_3672,N_3424,N_3587);
nor U3673 (N_3673,N_3585,N_3532);
and U3674 (N_3674,N_3553,N_3410);
or U3675 (N_3675,N_3544,N_3445);
or U3676 (N_3676,N_3487,N_3433);
nand U3677 (N_3677,N_3539,N_3501);
nand U3678 (N_3678,N_3527,N_3491);
nand U3679 (N_3679,N_3484,N_3460);
nor U3680 (N_3680,N_3499,N_3576);
nand U3681 (N_3681,N_3599,N_3584);
or U3682 (N_3682,N_3515,N_3582);
nor U3683 (N_3683,N_3555,N_3483);
or U3684 (N_3684,N_3447,N_3592);
nor U3685 (N_3685,N_3533,N_3552);
nor U3686 (N_3686,N_3561,N_3570);
nand U3687 (N_3687,N_3443,N_3401);
or U3688 (N_3688,N_3581,N_3475);
nor U3689 (N_3689,N_3449,N_3486);
or U3690 (N_3690,N_3568,N_3518);
xor U3691 (N_3691,N_3506,N_3505);
and U3692 (N_3692,N_3411,N_3481);
or U3693 (N_3693,N_3503,N_3474);
nand U3694 (N_3694,N_3546,N_3541);
nand U3695 (N_3695,N_3415,N_3421);
and U3696 (N_3696,N_3482,N_3521);
xor U3697 (N_3697,N_3417,N_3522);
xnor U3698 (N_3698,N_3520,N_3588);
or U3699 (N_3699,N_3589,N_3461);
nand U3700 (N_3700,N_3562,N_3574);
and U3701 (N_3701,N_3411,N_3424);
nor U3702 (N_3702,N_3516,N_3533);
nor U3703 (N_3703,N_3502,N_3450);
and U3704 (N_3704,N_3488,N_3532);
nand U3705 (N_3705,N_3433,N_3522);
nand U3706 (N_3706,N_3419,N_3408);
xor U3707 (N_3707,N_3560,N_3454);
or U3708 (N_3708,N_3495,N_3562);
or U3709 (N_3709,N_3590,N_3555);
xnor U3710 (N_3710,N_3572,N_3432);
or U3711 (N_3711,N_3530,N_3543);
or U3712 (N_3712,N_3547,N_3564);
and U3713 (N_3713,N_3400,N_3428);
and U3714 (N_3714,N_3426,N_3584);
xnor U3715 (N_3715,N_3412,N_3470);
or U3716 (N_3716,N_3478,N_3480);
nand U3717 (N_3717,N_3517,N_3491);
xor U3718 (N_3718,N_3464,N_3486);
nand U3719 (N_3719,N_3530,N_3401);
nand U3720 (N_3720,N_3422,N_3566);
xnor U3721 (N_3721,N_3462,N_3458);
xor U3722 (N_3722,N_3564,N_3510);
xnor U3723 (N_3723,N_3558,N_3406);
xor U3724 (N_3724,N_3493,N_3569);
or U3725 (N_3725,N_3520,N_3420);
nor U3726 (N_3726,N_3438,N_3435);
nor U3727 (N_3727,N_3523,N_3514);
nand U3728 (N_3728,N_3563,N_3414);
nand U3729 (N_3729,N_3541,N_3583);
xnor U3730 (N_3730,N_3450,N_3522);
and U3731 (N_3731,N_3595,N_3574);
nor U3732 (N_3732,N_3495,N_3591);
or U3733 (N_3733,N_3476,N_3431);
nor U3734 (N_3734,N_3489,N_3529);
nor U3735 (N_3735,N_3517,N_3594);
and U3736 (N_3736,N_3462,N_3419);
or U3737 (N_3737,N_3506,N_3568);
nand U3738 (N_3738,N_3520,N_3567);
xnor U3739 (N_3739,N_3472,N_3413);
nand U3740 (N_3740,N_3548,N_3480);
nand U3741 (N_3741,N_3437,N_3543);
xnor U3742 (N_3742,N_3578,N_3541);
nand U3743 (N_3743,N_3523,N_3486);
or U3744 (N_3744,N_3400,N_3486);
or U3745 (N_3745,N_3490,N_3479);
or U3746 (N_3746,N_3401,N_3584);
nor U3747 (N_3747,N_3471,N_3532);
nor U3748 (N_3748,N_3460,N_3578);
or U3749 (N_3749,N_3523,N_3512);
nand U3750 (N_3750,N_3510,N_3492);
and U3751 (N_3751,N_3576,N_3485);
nor U3752 (N_3752,N_3504,N_3522);
nor U3753 (N_3753,N_3446,N_3552);
xnor U3754 (N_3754,N_3575,N_3581);
or U3755 (N_3755,N_3487,N_3512);
and U3756 (N_3756,N_3576,N_3476);
or U3757 (N_3757,N_3521,N_3548);
xnor U3758 (N_3758,N_3486,N_3424);
nand U3759 (N_3759,N_3592,N_3478);
or U3760 (N_3760,N_3513,N_3515);
or U3761 (N_3761,N_3457,N_3514);
xor U3762 (N_3762,N_3512,N_3518);
and U3763 (N_3763,N_3475,N_3454);
nor U3764 (N_3764,N_3534,N_3597);
xnor U3765 (N_3765,N_3442,N_3499);
nand U3766 (N_3766,N_3552,N_3469);
or U3767 (N_3767,N_3404,N_3401);
xor U3768 (N_3768,N_3449,N_3579);
nor U3769 (N_3769,N_3468,N_3400);
nand U3770 (N_3770,N_3537,N_3593);
or U3771 (N_3771,N_3411,N_3596);
xnor U3772 (N_3772,N_3466,N_3529);
and U3773 (N_3773,N_3501,N_3403);
nand U3774 (N_3774,N_3551,N_3425);
nor U3775 (N_3775,N_3442,N_3465);
nor U3776 (N_3776,N_3483,N_3553);
nor U3777 (N_3777,N_3471,N_3570);
and U3778 (N_3778,N_3550,N_3585);
nand U3779 (N_3779,N_3515,N_3507);
nor U3780 (N_3780,N_3538,N_3580);
nand U3781 (N_3781,N_3421,N_3436);
and U3782 (N_3782,N_3463,N_3530);
xor U3783 (N_3783,N_3459,N_3550);
nor U3784 (N_3784,N_3425,N_3536);
nand U3785 (N_3785,N_3530,N_3528);
xor U3786 (N_3786,N_3459,N_3535);
and U3787 (N_3787,N_3503,N_3424);
xnor U3788 (N_3788,N_3423,N_3558);
or U3789 (N_3789,N_3587,N_3400);
nand U3790 (N_3790,N_3536,N_3401);
nor U3791 (N_3791,N_3431,N_3467);
nand U3792 (N_3792,N_3515,N_3420);
or U3793 (N_3793,N_3408,N_3460);
nand U3794 (N_3794,N_3573,N_3580);
or U3795 (N_3795,N_3404,N_3461);
nor U3796 (N_3796,N_3509,N_3544);
nand U3797 (N_3797,N_3471,N_3428);
xor U3798 (N_3798,N_3580,N_3489);
or U3799 (N_3799,N_3480,N_3535);
xor U3800 (N_3800,N_3717,N_3650);
or U3801 (N_3801,N_3793,N_3643);
xor U3802 (N_3802,N_3774,N_3699);
nand U3803 (N_3803,N_3614,N_3683);
xor U3804 (N_3804,N_3630,N_3675);
or U3805 (N_3805,N_3606,N_3746);
nand U3806 (N_3806,N_3637,N_3732);
or U3807 (N_3807,N_3751,N_3693);
and U3808 (N_3808,N_3765,N_3784);
or U3809 (N_3809,N_3604,N_3674);
nor U3810 (N_3810,N_3678,N_3617);
or U3811 (N_3811,N_3785,N_3748);
and U3812 (N_3812,N_3640,N_3691);
nor U3813 (N_3813,N_3631,N_3777);
or U3814 (N_3814,N_3641,N_3649);
and U3815 (N_3815,N_3670,N_3638);
or U3816 (N_3816,N_3610,N_3627);
nor U3817 (N_3817,N_3710,N_3706);
or U3818 (N_3818,N_3620,N_3787);
and U3819 (N_3819,N_3716,N_3718);
or U3820 (N_3820,N_3734,N_3753);
xnor U3821 (N_3821,N_3619,N_3736);
nor U3822 (N_3822,N_3731,N_3665);
and U3823 (N_3823,N_3618,N_3671);
nor U3824 (N_3824,N_3708,N_3611);
nand U3825 (N_3825,N_3729,N_3696);
xor U3826 (N_3826,N_3791,N_3714);
xnor U3827 (N_3827,N_3612,N_3603);
nand U3828 (N_3828,N_3656,N_3642);
nand U3829 (N_3829,N_3616,N_3752);
or U3830 (N_3830,N_3712,N_3795);
xor U3831 (N_3831,N_3715,N_3644);
or U3832 (N_3832,N_3609,N_3763);
or U3833 (N_3833,N_3738,N_3628);
or U3834 (N_3834,N_3781,N_3672);
nand U3835 (N_3835,N_3632,N_3663);
or U3836 (N_3836,N_3747,N_3694);
nor U3837 (N_3837,N_3759,N_3709);
or U3838 (N_3838,N_3662,N_3705);
xor U3839 (N_3839,N_3745,N_3739);
nor U3840 (N_3840,N_3756,N_3703);
and U3841 (N_3841,N_3783,N_3666);
and U3842 (N_3842,N_3677,N_3761);
xor U3843 (N_3843,N_3668,N_3647);
or U3844 (N_3844,N_3687,N_3764);
or U3845 (N_3845,N_3776,N_3689);
xnor U3846 (N_3846,N_3725,N_3797);
nor U3847 (N_3847,N_3772,N_3702);
and U3848 (N_3848,N_3704,N_3646);
or U3849 (N_3849,N_3779,N_3654);
nand U3850 (N_3850,N_3684,N_3770);
nor U3851 (N_3851,N_3664,N_3790);
xor U3852 (N_3852,N_3771,N_3697);
and U3853 (N_3853,N_3636,N_3648);
xor U3854 (N_3854,N_3608,N_3722);
xor U3855 (N_3855,N_3707,N_3645);
xor U3856 (N_3856,N_3629,N_3701);
or U3857 (N_3857,N_3723,N_3667);
or U3858 (N_3858,N_3624,N_3639);
or U3859 (N_3859,N_3773,N_3615);
xnor U3860 (N_3860,N_3623,N_3653);
nand U3861 (N_3861,N_3726,N_3735);
and U3862 (N_3862,N_3767,N_3601);
or U3863 (N_3863,N_3760,N_3741);
xor U3864 (N_3864,N_3762,N_3657);
xnor U3865 (N_3865,N_3690,N_3676);
nor U3866 (N_3866,N_3652,N_3799);
nor U3867 (N_3867,N_3733,N_3655);
and U3868 (N_3868,N_3659,N_3755);
nand U3869 (N_3869,N_3788,N_3768);
and U3870 (N_3870,N_3782,N_3794);
xnor U3871 (N_3871,N_3658,N_3721);
xnor U3872 (N_3872,N_3730,N_3713);
nand U3873 (N_3873,N_3673,N_3724);
and U3874 (N_3874,N_3698,N_3622);
nand U3875 (N_3875,N_3719,N_3625);
nor U3876 (N_3876,N_3681,N_3786);
nand U3877 (N_3877,N_3633,N_3749);
nand U3878 (N_3878,N_3743,N_3780);
nor U3879 (N_3879,N_3792,N_3685);
nand U3880 (N_3880,N_3635,N_3740);
nor U3881 (N_3881,N_3798,N_3742);
xor U3882 (N_3882,N_3682,N_3789);
xor U3883 (N_3883,N_3728,N_3679);
and U3884 (N_3884,N_3692,N_3778);
or U3885 (N_3885,N_3626,N_3661);
or U3886 (N_3886,N_3769,N_3700);
nor U3887 (N_3887,N_3669,N_3775);
nand U3888 (N_3888,N_3727,N_3607);
nor U3889 (N_3889,N_3680,N_3754);
or U3890 (N_3890,N_3602,N_3600);
and U3891 (N_3891,N_3758,N_3605);
nor U3892 (N_3892,N_3796,N_3660);
and U3893 (N_3893,N_3621,N_3757);
nor U3894 (N_3894,N_3613,N_3695);
nand U3895 (N_3895,N_3737,N_3766);
and U3896 (N_3896,N_3720,N_3750);
nand U3897 (N_3897,N_3688,N_3651);
and U3898 (N_3898,N_3711,N_3686);
nor U3899 (N_3899,N_3634,N_3744);
nor U3900 (N_3900,N_3771,N_3767);
nor U3901 (N_3901,N_3761,N_3645);
xnor U3902 (N_3902,N_3723,N_3701);
and U3903 (N_3903,N_3730,N_3702);
or U3904 (N_3904,N_3647,N_3695);
or U3905 (N_3905,N_3664,N_3785);
nor U3906 (N_3906,N_3762,N_3620);
and U3907 (N_3907,N_3693,N_3719);
xnor U3908 (N_3908,N_3758,N_3639);
nor U3909 (N_3909,N_3646,N_3643);
or U3910 (N_3910,N_3766,N_3603);
and U3911 (N_3911,N_3627,N_3752);
nand U3912 (N_3912,N_3752,N_3704);
nand U3913 (N_3913,N_3692,N_3785);
or U3914 (N_3914,N_3723,N_3779);
nand U3915 (N_3915,N_3657,N_3767);
and U3916 (N_3916,N_3615,N_3667);
nand U3917 (N_3917,N_3679,N_3663);
and U3918 (N_3918,N_3651,N_3666);
and U3919 (N_3919,N_3605,N_3629);
or U3920 (N_3920,N_3760,N_3663);
nor U3921 (N_3921,N_3788,N_3743);
nand U3922 (N_3922,N_3774,N_3656);
nor U3923 (N_3923,N_3789,N_3775);
and U3924 (N_3924,N_3633,N_3688);
xor U3925 (N_3925,N_3715,N_3655);
and U3926 (N_3926,N_3756,N_3679);
or U3927 (N_3927,N_3756,N_3617);
or U3928 (N_3928,N_3798,N_3660);
nand U3929 (N_3929,N_3705,N_3636);
xor U3930 (N_3930,N_3608,N_3730);
and U3931 (N_3931,N_3612,N_3704);
and U3932 (N_3932,N_3738,N_3627);
xnor U3933 (N_3933,N_3620,N_3779);
nand U3934 (N_3934,N_3654,N_3672);
or U3935 (N_3935,N_3612,N_3629);
nand U3936 (N_3936,N_3657,N_3688);
xor U3937 (N_3937,N_3660,N_3749);
nand U3938 (N_3938,N_3654,N_3665);
nor U3939 (N_3939,N_3704,N_3685);
xnor U3940 (N_3940,N_3664,N_3707);
xor U3941 (N_3941,N_3664,N_3612);
and U3942 (N_3942,N_3766,N_3669);
and U3943 (N_3943,N_3602,N_3677);
or U3944 (N_3944,N_3670,N_3768);
nand U3945 (N_3945,N_3675,N_3733);
nand U3946 (N_3946,N_3620,N_3770);
or U3947 (N_3947,N_3741,N_3748);
nor U3948 (N_3948,N_3615,N_3775);
and U3949 (N_3949,N_3783,N_3608);
and U3950 (N_3950,N_3654,N_3700);
nor U3951 (N_3951,N_3770,N_3601);
xor U3952 (N_3952,N_3783,N_3619);
nand U3953 (N_3953,N_3784,N_3608);
nor U3954 (N_3954,N_3619,N_3766);
and U3955 (N_3955,N_3719,N_3685);
xnor U3956 (N_3956,N_3607,N_3629);
or U3957 (N_3957,N_3765,N_3790);
and U3958 (N_3958,N_3734,N_3729);
xor U3959 (N_3959,N_3635,N_3679);
nor U3960 (N_3960,N_3775,N_3630);
and U3961 (N_3961,N_3772,N_3703);
nand U3962 (N_3962,N_3762,N_3664);
nor U3963 (N_3963,N_3713,N_3604);
nand U3964 (N_3964,N_3650,N_3625);
xnor U3965 (N_3965,N_3664,N_3709);
nor U3966 (N_3966,N_3726,N_3687);
nand U3967 (N_3967,N_3647,N_3721);
or U3968 (N_3968,N_3773,N_3662);
nand U3969 (N_3969,N_3631,N_3662);
nand U3970 (N_3970,N_3738,N_3695);
nor U3971 (N_3971,N_3792,N_3736);
and U3972 (N_3972,N_3761,N_3652);
xor U3973 (N_3973,N_3668,N_3696);
xnor U3974 (N_3974,N_3608,N_3733);
nor U3975 (N_3975,N_3795,N_3605);
or U3976 (N_3976,N_3637,N_3616);
and U3977 (N_3977,N_3740,N_3642);
nand U3978 (N_3978,N_3749,N_3617);
nand U3979 (N_3979,N_3634,N_3719);
and U3980 (N_3980,N_3746,N_3776);
nand U3981 (N_3981,N_3649,N_3780);
nor U3982 (N_3982,N_3704,N_3629);
nand U3983 (N_3983,N_3706,N_3769);
nand U3984 (N_3984,N_3721,N_3741);
nand U3985 (N_3985,N_3792,N_3710);
and U3986 (N_3986,N_3792,N_3659);
or U3987 (N_3987,N_3756,N_3670);
or U3988 (N_3988,N_3794,N_3783);
xnor U3989 (N_3989,N_3659,N_3673);
nand U3990 (N_3990,N_3764,N_3785);
nand U3991 (N_3991,N_3722,N_3786);
nand U3992 (N_3992,N_3649,N_3788);
nor U3993 (N_3993,N_3707,N_3712);
nor U3994 (N_3994,N_3787,N_3676);
xor U3995 (N_3995,N_3704,N_3682);
or U3996 (N_3996,N_3695,N_3606);
nor U3997 (N_3997,N_3651,N_3616);
or U3998 (N_3998,N_3751,N_3606);
and U3999 (N_3999,N_3621,N_3663);
xnor U4000 (N_4000,N_3979,N_3803);
or U4001 (N_4001,N_3832,N_3956);
xor U4002 (N_4002,N_3865,N_3823);
xor U4003 (N_4003,N_3961,N_3836);
nand U4004 (N_4004,N_3895,N_3872);
nor U4005 (N_4005,N_3971,N_3863);
or U4006 (N_4006,N_3871,N_3985);
nand U4007 (N_4007,N_3842,N_3897);
xor U4008 (N_4008,N_3870,N_3957);
and U4009 (N_4009,N_3876,N_3964);
xnor U4010 (N_4010,N_3954,N_3918);
nand U4011 (N_4011,N_3931,N_3883);
nand U4012 (N_4012,N_3910,N_3952);
and U4013 (N_4013,N_3982,N_3824);
nand U4014 (N_4014,N_3840,N_3846);
nand U4015 (N_4015,N_3990,N_3942);
or U4016 (N_4016,N_3830,N_3955);
nor U4017 (N_4017,N_3810,N_3940);
and U4018 (N_4018,N_3906,N_3953);
and U4019 (N_4019,N_3959,N_3843);
and U4020 (N_4020,N_3914,N_3888);
xor U4021 (N_4021,N_3907,N_3977);
or U4022 (N_4022,N_3894,N_3978);
nand U4023 (N_4023,N_3908,N_3904);
nand U4024 (N_4024,N_3944,N_3868);
nor U4025 (N_4025,N_3885,N_3976);
nor U4026 (N_4026,N_3975,N_3889);
and U4027 (N_4027,N_3951,N_3828);
xor U4028 (N_4028,N_3972,N_3877);
or U4029 (N_4029,N_3852,N_3800);
nand U4030 (N_4030,N_3847,N_3815);
and U4031 (N_4031,N_3802,N_3822);
and U4032 (N_4032,N_3835,N_3821);
xor U4033 (N_4033,N_3893,N_3921);
nor U4034 (N_4034,N_3996,N_3864);
xor U4035 (N_4035,N_3991,N_3986);
and U4036 (N_4036,N_3860,N_3820);
or U4037 (N_4037,N_3981,N_3958);
nor U4038 (N_4038,N_3929,N_3880);
and U4039 (N_4039,N_3933,N_3818);
or U4040 (N_4040,N_3930,N_3999);
or U4041 (N_4041,N_3941,N_3817);
and U4042 (N_4042,N_3816,N_3851);
or U4043 (N_4043,N_3943,N_3899);
and U4044 (N_4044,N_3838,N_3915);
xnor U4045 (N_4045,N_3960,N_3890);
and U4046 (N_4046,N_3968,N_3973);
nand U4047 (N_4047,N_3917,N_3989);
or U4048 (N_4048,N_3903,N_3934);
nor U4049 (N_4049,N_3855,N_3969);
xnor U4050 (N_4050,N_3994,N_3833);
nor U4051 (N_4051,N_3873,N_3927);
xnor U4052 (N_4052,N_3850,N_3984);
or U4053 (N_4053,N_3965,N_3862);
or U4054 (N_4054,N_3966,N_3809);
nor U4055 (N_4055,N_3928,N_3892);
nand U4056 (N_4056,N_3920,N_3839);
nor U4057 (N_4057,N_3900,N_3980);
nand U4058 (N_4058,N_3845,N_3861);
nor U4059 (N_4059,N_3879,N_3806);
and U4060 (N_4060,N_3932,N_3801);
nor U4061 (N_4061,N_3948,N_3884);
and U4062 (N_4062,N_3938,N_3997);
and U4063 (N_4063,N_3913,N_3878);
xnor U4064 (N_4064,N_3831,N_3826);
nand U4065 (N_4065,N_3808,N_3812);
and U4066 (N_4066,N_3924,N_3858);
nor U4067 (N_4067,N_3967,N_3939);
nand U4068 (N_4068,N_3891,N_3912);
nor U4069 (N_4069,N_3827,N_3995);
or U4070 (N_4070,N_3935,N_3902);
or U4071 (N_4071,N_3882,N_3983);
nor U4072 (N_4072,N_3841,N_3998);
nor U4073 (N_4073,N_3992,N_3814);
nor U4074 (N_4074,N_3911,N_3962);
and U4075 (N_4075,N_3813,N_3898);
or U4076 (N_4076,N_3947,N_3926);
and U4077 (N_4077,N_3993,N_3849);
xnor U4078 (N_4078,N_3805,N_3937);
nor U4079 (N_4079,N_3874,N_3854);
or U4080 (N_4080,N_3844,N_3804);
or U4081 (N_4081,N_3909,N_3881);
xor U4082 (N_4082,N_3936,N_3988);
xnor U4083 (N_4083,N_3922,N_3974);
nand U4084 (N_4084,N_3825,N_3896);
or U4085 (N_4085,N_3857,N_3859);
and U4086 (N_4086,N_3869,N_3925);
nor U4087 (N_4087,N_3887,N_3950);
xnor U4088 (N_4088,N_3875,N_3949);
xnor U4089 (N_4089,N_3819,N_3853);
or U4090 (N_4090,N_3946,N_3837);
nand U4091 (N_4091,N_3963,N_3970);
and U4092 (N_4092,N_3905,N_3886);
and U4093 (N_4093,N_3867,N_3856);
nor U4094 (N_4094,N_3829,N_3811);
or U4095 (N_4095,N_3916,N_3848);
nand U4096 (N_4096,N_3834,N_3807);
nand U4097 (N_4097,N_3945,N_3919);
xnor U4098 (N_4098,N_3923,N_3866);
or U4099 (N_4099,N_3901,N_3987);
and U4100 (N_4100,N_3907,N_3952);
xor U4101 (N_4101,N_3857,N_3956);
or U4102 (N_4102,N_3845,N_3844);
nand U4103 (N_4103,N_3823,N_3996);
nand U4104 (N_4104,N_3827,N_3874);
nand U4105 (N_4105,N_3931,N_3835);
xor U4106 (N_4106,N_3839,N_3821);
nand U4107 (N_4107,N_3941,N_3990);
xor U4108 (N_4108,N_3967,N_3801);
and U4109 (N_4109,N_3835,N_3852);
xnor U4110 (N_4110,N_3978,N_3835);
nor U4111 (N_4111,N_3873,N_3918);
xnor U4112 (N_4112,N_3865,N_3977);
nor U4113 (N_4113,N_3977,N_3891);
nor U4114 (N_4114,N_3819,N_3928);
nand U4115 (N_4115,N_3875,N_3962);
nor U4116 (N_4116,N_3984,N_3972);
and U4117 (N_4117,N_3998,N_3915);
or U4118 (N_4118,N_3855,N_3891);
xnor U4119 (N_4119,N_3867,N_3810);
nor U4120 (N_4120,N_3975,N_3873);
nor U4121 (N_4121,N_3942,N_3917);
and U4122 (N_4122,N_3807,N_3918);
or U4123 (N_4123,N_3971,N_3825);
nand U4124 (N_4124,N_3843,N_3835);
nor U4125 (N_4125,N_3817,N_3880);
nand U4126 (N_4126,N_3848,N_3874);
xor U4127 (N_4127,N_3980,N_3816);
and U4128 (N_4128,N_3981,N_3948);
nor U4129 (N_4129,N_3869,N_3852);
xnor U4130 (N_4130,N_3934,N_3991);
xnor U4131 (N_4131,N_3812,N_3801);
or U4132 (N_4132,N_3983,N_3930);
and U4133 (N_4133,N_3893,N_3959);
and U4134 (N_4134,N_3892,N_3950);
or U4135 (N_4135,N_3874,N_3882);
or U4136 (N_4136,N_3828,N_3981);
nand U4137 (N_4137,N_3856,N_3866);
or U4138 (N_4138,N_3932,N_3952);
nor U4139 (N_4139,N_3864,N_3801);
xnor U4140 (N_4140,N_3853,N_3907);
nand U4141 (N_4141,N_3913,N_3866);
nor U4142 (N_4142,N_3835,N_3982);
or U4143 (N_4143,N_3842,N_3849);
xnor U4144 (N_4144,N_3928,N_3809);
nor U4145 (N_4145,N_3985,N_3823);
and U4146 (N_4146,N_3950,N_3987);
nand U4147 (N_4147,N_3972,N_3988);
xnor U4148 (N_4148,N_3883,N_3863);
nand U4149 (N_4149,N_3885,N_3817);
or U4150 (N_4150,N_3930,N_3895);
and U4151 (N_4151,N_3862,N_3898);
nor U4152 (N_4152,N_3985,N_3976);
or U4153 (N_4153,N_3808,N_3909);
nand U4154 (N_4154,N_3847,N_3939);
or U4155 (N_4155,N_3958,N_3969);
or U4156 (N_4156,N_3895,N_3881);
nor U4157 (N_4157,N_3995,N_3903);
nor U4158 (N_4158,N_3822,N_3954);
and U4159 (N_4159,N_3893,N_3837);
and U4160 (N_4160,N_3909,N_3812);
xor U4161 (N_4161,N_3916,N_3865);
xnor U4162 (N_4162,N_3850,N_3920);
nand U4163 (N_4163,N_3998,N_3936);
xnor U4164 (N_4164,N_3857,N_3825);
nand U4165 (N_4165,N_3979,N_3817);
nand U4166 (N_4166,N_3917,N_3813);
and U4167 (N_4167,N_3845,N_3821);
nor U4168 (N_4168,N_3800,N_3838);
or U4169 (N_4169,N_3929,N_3830);
xnor U4170 (N_4170,N_3804,N_3850);
nand U4171 (N_4171,N_3907,N_3962);
and U4172 (N_4172,N_3953,N_3838);
xor U4173 (N_4173,N_3883,N_3946);
xor U4174 (N_4174,N_3974,N_3808);
and U4175 (N_4175,N_3828,N_3841);
nor U4176 (N_4176,N_3816,N_3847);
xnor U4177 (N_4177,N_3961,N_3889);
nand U4178 (N_4178,N_3881,N_3897);
or U4179 (N_4179,N_3952,N_3942);
or U4180 (N_4180,N_3876,N_3946);
and U4181 (N_4181,N_3892,N_3940);
xor U4182 (N_4182,N_3999,N_3891);
or U4183 (N_4183,N_3895,N_3812);
xor U4184 (N_4184,N_3987,N_3937);
nor U4185 (N_4185,N_3970,N_3944);
and U4186 (N_4186,N_3828,N_3931);
and U4187 (N_4187,N_3833,N_3843);
xor U4188 (N_4188,N_3967,N_3981);
or U4189 (N_4189,N_3838,N_3836);
and U4190 (N_4190,N_3932,N_3935);
or U4191 (N_4191,N_3915,N_3972);
and U4192 (N_4192,N_3830,N_3875);
nor U4193 (N_4193,N_3863,N_3949);
or U4194 (N_4194,N_3945,N_3865);
nand U4195 (N_4195,N_3996,N_3887);
and U4196 (N_4196,N_3955,N_3861);
xor U4197 (N_4197,N_3980,N_3975);
and U4198 (N_4198,N_3961,N_3843);
nor U4199 (N_4199,N_3865,N_3942);
nand U4200 (N_4200,N_4022,N_4077);
nor U4201 (N_4201,N_4154,N_4126);
or U4202 (N_4202,N_4108,N_4132);
nand U4203 (N_4203,N_4041,N_4046);
and U4204 (N_4204,N_4009,N_4111);
nor U4205 (N_4205,N_4191,N_4002);
and U4206 (N_4206,N_4184,N_4113);
xnor U4207 (N_4207,N_4166,N_4155);
or U4208 (N_4208,N_4019,N_4138);
nand U4209 (N_4209,N_4016,N_4035);
nor U4210 (N_4210,N_4068,N_4038);
xor U4211 (N_4211,N_4027,N_4193);
xnor U4212 (N_4212,N_4144,N_4040);
or U4213 (N_4213,N_4175,N_4171);
or U4214 (N_4214,N_4042,N_4092);
or U4215 (N_4215,N_4026,N_4010);
or U4216 (N_4216,N_4051,N_4061);
nor U4217 (N_4217,N_4099,N_4018);
xor U4218 (N_4218,N_4090,N_4196);
nand U4219 (N_4219,N_4140,N_4112);
xnor U4220 (N_4220,N_4178,N_4174);
nor U4221 (N_4221,N_4074,N_4122);
xnor U4222 (N_4222,N_4105,N_4199);
xor U4223 (N_4223,N_4078,N_4153);
nor U4224 (N_4224,N_4001,N_4192);
or U4225 (N_4225,N_4062,N_4173);
xor U4226 (N_4226,N_4063,N_4005);
nor U4227 (N_4227,N_4120,N_4034);
xnor U4228 (N_4228,N_4057,N_4043);
or U4229 (N_4229,N_4011,N_4124);
and U4230 (N_4230,N_4020,N_4080);
or U4231 (N_4231,N_4064,N_4006);
xor U4232 (N_4232,N_4045,N_4013);
nand U4233 (N_4233,N_4036,N_4150);
xnor U4234 (N_4234,N_4170,N_4181);
and U4235 (N_4235,N_4141,N_4121);
xor U4236 (N_4236,N_4176,N_4130);
and U4237 (N_4237,N_4033,N_4028);
nor U4238 (N_4238,N_4156,N_4101);
and U4239 (N_4239,N_4125,N_4084);
or U4240 (N_4240,N_4085,N_4071);
nor U4241 (N_4241,N_4169,N_4116);
xor U4242 (N_4242,N_4148,N_4008);
xor U4243 (N_4243,N_4044,N_4098);
nand U4244 (N_4244,N_4052,N_4159);
and U4245 (N_4245,N_4152,N_4114);
and U4246 (N_4246,N_4056,N_4082);
nor U4247 (N_4247,N_4086,N_4023);
or U4248 (N_4248,N_4160,N_4190);
nand U4249 (N_4249,N_4142,N_4177);
nand U4250 (N_4250,N_4146,N_4048);
nand U4251 (N_4251,N_4197,N_4164);
nor U4252 (N_4252,N_4198,N_4089);
xnor U4253 (N_4253,N_4187,N_4032);
nand U4254 (N_4254,N_4151,N_4093);
nor U4255 (N_4255,N_4054,N_4070);
or U4256 (N_4256,N_4115,N_4157);
or U4257 (N_4257,N_4096,N_4119);
nand U4258 (N_4258,N_4188,N_4147);
xor U4259 (N_4259,N_4004,N_4185);
xnor U4260 (N_4260,N_4129,N_4037);
or U4261 (N_4261,N_4088,N_4059);
nand U4262 (N_4262,N_4072,N_4110);
or U4263 (N_4263,N_4118,N_4106);
nor U4264 (N_4264,N_4149,N_4183);
nand U4265 (N_4265,N_4135,N_4097);
or U4266 (N_4266,N_4029,N_4047);
or U4267 (N_4267,N_4179,N_4075);
xor U4268 (N_4268,N_4014,N_4102);
or U4269 (N_4269,N_4058,N_4131);
or U4270 (N_4270,N_4065,N_4060);
nor U4271 (N_4271,N_4133,N_4031);
xor U4272 (N_4272,N_4145,N_4158);
nand U4273 (N_4273,N_4073,N_4134);
nor U4274 (N_4274,N_4087,N_4039);
or U4275 (N_4275,N_4021,N_4000);
nor U4276 (N_4276,N_4189,N_4163);
and U4277 (N_4277,N_4007,N_4172);
nor U4278 (N_4278,N_4117,N_4017);
nand U4279 (N_4279,N_4012,N_4100);
or U4280 (N_4280,N_4186,N_4103);
xnor U4281 (N_4281,N_4024,N_4182);
nand U4282 (N_4282,N_4180,N_4194);
nand U4283 (N_4283,N_4109,N_4076);
nor U4284 (N_4284,N_4049,N_4094);
or U4285 (N_4285,N_4168,N_4050);
nor U4286 (N_4286,N_4136,N_4161);
nor U4287 (N_4287,N_4123,N_4053);
xnor U4288 (N_4288,N_4137,N_4066);
or U4289 (N_4289,N_4079,N_4095);
nor U4290 (N_4290,N_4055,N_4195);
nand U4291 (N_4291,N_4081,N_4003);
nand U4292 (N_4292,N_4127,N_4083);
and U4293 (N_4293,N_4025,N_4165);
and U4294 (N_4294,N_4069,N_4067);
and U4295 (N_4295,N_4091,N_4015);
or U4296 (N_4296,N_4030,N_4162);
and U4297 (N_4297,N_4107,N_4128);
nand U4298 (N_4298,N_4139,N_4167);
or U4299 (N_4299,N_4143,N_4104);
nand U4300 (N_4300,N_4022,N_4016);
nor U4301 (N_4301,N_4129,N_4141);
or U4302 (N_4302,N_4128,N_4075);
and U4303 (N_4303,N_4094,N_4033);
nor U4304 (N_4304,N_4196,N_4127);
nor U4305 (N_4305,N_4184,N_4069);
nor U4306 (N_4306,N_4022,N_4179);
nand U4307 (N_4307,N_4099,N_4095);
or U4308 (N_4308,N_4032,N_4108);
nand U4309 (N_4309,N_4042,N_4186);
and U4310 (N_4310,N_4089,N_4038);
xnor U4311 (N_4311,N_4002,N_4062);
or U4312 (N_4312,N_4112,N_4191);
nor U4313 (N_4313,N_4189,N_4085);
nand U4314 (N_4314,N_4055,N_4113);
nand U4315 (N_4315,N_4089,N_4154);
xnor U4316 (N_4316,N_4050,N_4124);
and U4317 (N_4317,N_4151,N_4173);
and U4318 (N_4318,N_4111,N_4103);
nor U4319 (N_4319,N_4184,N_4140);
xor U4320 (N_4320,N_4029,N_4006);
nor U4321 (N_4321,N_4199,N_4163);
and U4322 (N_4322,N_4154,N_4052);
xnor U4323 (N_4323,N_4169,N_4132);
xor U4324 (N_4324,N_4032,N_4048);
xor U4325 (N_4325,N_4009,N_4118);
nand U4326 (N_4326,N_4149,N_4098);
xnor U4327 (N_4327,N_4014,N_4137);
nor U4328 (N_4328,N_4009,N_4008);
xor U4329 (N_4329,N_4030,N_4164);
xnor U4330 (N_4330,N_4173,N_4150);
nand U4331 (N_4331,N_4021,N_4146);
or U4332 (N_4332,N_4083,N_4124);
nand U4333 (N_4333,N_4142,N_4110);
or U4334 (N_4334,N_4195,N_4073);
nand U4335 (N_4335,N_4196,N_4103);
or U4336 (N_4336,N_4105,N_4050);
or U4337 (N_4337,N_4143,N_4124);
xor U4338 (N_4338,N_4175,N_4069);
or U4339 (N_4339,N_4189,N_4140);
and U4340 (N_4340,N_4064,N_4012);
xor U4341 (N_4341,N_4015,N_4036);
nor U4342 (N_4342,N_4155,N_4135);
nand U4343 (N_4343,N_4140,N_4125);
and U4344 (N_4344,N_4076,N_4158);
and U4345 (N_4345,N_4094,N_4140);
xnor U4346 (N_4346,N_4164,N_4171);
and U4347 (N_4347,N_4177,N_4000);
nand U4348 (N_4348,N_4158,N_4000);
or U4349 (N_4349,N_4074,N_4117);
and U4350 (N_4350,N_4080,N_4125);
and U4351 (N_4351,N_4151,N_4062);
nor U4352 (N_4352,N_4104,N_4082);
or U4353 (N_4353,N_4107,N_4131);
or U4354 (N_4354,N_4030,N_4095);
xnor U4355 (N_4355,N_4079,N_4136);
nor U4356 (N_4356,N_4054,N_4130);
or U4357 (N_4357,N_4065,N_4174);
nor U4358 (N_4358,N_4006,N_4108);
and U4359 (N_4359,N_4152,N_4053);
nor U4360 (N_4360,N_4055,N_4030);
and U4361 (N_4361,N_4051,N_4094);
nand U4362 (N_4362,N_4076,N_4095);
nor U4363 (N_4363,N_4123,N_4019);
nand U4364 (N_4364,N_4038,N_4003);
and U4365 (N_4365,N_4141,N_4018);
xor U4366 (N_4366,N_4097,N_4055);
and U4367 (N_4367,N_4003,N_4138);
nand U4368 (N_4368,N_4165,N_4089);
and U4369 (N_4369,N_4072,N_4173);
nor U4370 (N_4370,N_4137,N_4112);
and U4371 (N_4371,N_4091,N_4040);
nor U4372 (N_4372,N_4058,N_4010);
nand U4373 (N_4373,N_4118,N_4016);
nor U4374 (N_4374,N_4133,N_4169);
nand U4375 (N_4375,N_4156,N_4066);
or U4376 (N_4376,N_4041,N_4154);
nand U4377 (N_4377,N_4193,N_4103);
and U4378 (N_4378,N_4095,N_4070);
and U4379 (N_4379,N_4009,N_4080);
nor U4380 (N_4380,N_4081,N_4062);
or U4381 (N_4381,N_4057,N_4078);
nand U4382 (N_4382,N_4021,N_4086);
nor U4383 (N_4383,N_4060,N_4006);
and U4384 (N_4384,N_4004,N_4043);
and U4385 (N_4385,N_4016,N_4190);
nand U4386 (N_4386,N_4193,N_4083);
nor U4387 (N_4387,N_4062,N_4078);
nor U4388 (N_4388,N_4046,N_4126);
nand U4389 (N_4389,N_4189,N_4077);
nand U4390 (N_4390,N_4105,N_4027);
xnor U4391 (N_4391,N_4048,N_4111);
xnor U4392 (N_4392,N_4131,N_4171);
nor U4393 (N_4393,N_4125,N_4028);
xnor U4394 (N_4394,N_4007,N_4109);
and U4395 (N_4395,N_4087,N_4096);
xnor U4396 (N_4396,N_4128,N_4119);
xnor U4397 (N_4397,N_4104,N_4087);
xnor U4398 (N_4398,N_4140,N_4107);
xnor U4399 (N_4399,N_4082,N_4185);
nor U4400 (N_4400,N_4378,N_4219);
nor U4401 (N_4401,N_4286,N_4223);
nand U4402 (N_4402,N_4247,N_4369);
or U4403 (N_4403,N_4208,N_4243);
and U4404 (N_4404,N_4248,N_4245);
or U4405 (N_4405,N_4314,N_4298);
nor U4406 (N_4406,N_4250,N_4399);
nand U4407 (N_4407,N_4278,N_4391);
nor U4408 (N_4408,N_4255,N_4239);
nand U4409 (N_4409,N_4336,N_4319);
xnor U4410 (N_4410,N_4232,N_4218);
and U4411 (N_4411,N_4241,N_4386);
or U4412 (N_4412,N_4394,N_4200);
or U4413 (N_4413,N_4383,N_4290);
and U4414 (N_4414,N_4261,N_4252);
nand U4415 (N_4415,N_4274,N_4367);
nand U4416 (N_4416,N_4393,N_4253);
nor U4417 (N_4417,N_4307,N_4375);
nand U4418 (N_4418,N_4352,N_4339);
nand U4419 (N_4419,N_4364,N_4311);
xnor U4420 (N_4420,N_4348,N_4272);
nor U4421 (N_4421,N_4287,N_4216);
nand U4422 (N_4422,N_4318,N_4275);
nor U4423 (N_4423,N_4358,N_4396);
and U4424 (N_4424,N_4395,N_4237);
xnor U4425 (N_4425,N_4342,N_4266);
and U4426 (N_4426,N_4257,N_4256);
xnor U4427 (N_4427,N_4310,N_4203);
or U4428 (N_4428,N_4202,N_4335);
nor U4429 (N_4429,N_4331,N_4337);
nand U4430 (N_4430,N_4224,N_4258);
nor U4431 (N_4431,N_4388,N_4326);
and U4432 (N_4432,N_4284,N_4236);
nand U4433 (N_4433,N_4238,N_4276);
or U4434 (N_4434,N_4327,N_4301);
and U4435 (N_4435,N_4332,N_4281);
or U4436 (N_4436,N_4270,N_4366);
or U4437 (N_4437,N_4347,N_4268);
and U4438 (N_4438,N_4242,N_4246);
xor U4439 (N_4439,N_4338,N_4211);
nand U4440 (N_4440,N_4225,N_4244);
nand U4441 (N_4441,N_4215,N_4315);
or U4442 (N_4442,N_4341,N_4385);
or U4443 (N_4443,N_4285,N_4325);
xor U4444 (N_4444,N_4259,N_4212);
nand U4445 (N_4445,N_4296,N_4260);
or U4446 (N_4446,N_4373,N_4220);
nor U4447 (N_4447,N_4350,N_4390);
xnor U4448 (N_4448,N_4322,N_4230);
or U4449 (N_4449,N_4271,N_4324);
xor U4450 (N_4450,N_4262,N_4309);
xor U4451 (N_4451,N_4300,N_4283);
nor U4452 (N_4452,N_4345,N_4392);
nor U4453 (N_4453,N_4360,N_4289);
nor U4454 (N_4454,N_4376,N_4240);
xor U4455 (N_4455,N_4389,N_4294);
nand U4456 (N_4456,N_4277,N_4288);
xnor U4457 (N_4457,N_4353,N_4302);
xor U4458 (N_4458,N_4233,N_4282);
xor U4459 (N_4459,N_4306,N_4303);
nor U4460 (N_4460,N_4299,N_4228);
or U4461 (N_4461,N_4354,N_4265);
and U4462 (N_4462,N_4205,N_4214);
or U4463 (N_4463,N_4361,N_4201);
xnor U4464 (N_4464,N_4397,N_4351);
nand U4465 (N_4465,N_4280,N_4297);
xnor U4466 (N_4466,N_4359,N_4363);
xor U4467 (N_4467,N_4209,N_4356);
xor U4468 (N_4468,N_4382,N_4380);
xnor U4469 (N_4469,N_4372,N_4206);
xor U4470 (N_4470,N_4334,N_4330);
xor U4471 (N_4471,N_4362,N_4304);
nor U4472 (N_4472,N_4316,N_4387);
xnor U4473 (N_4473,N_4371,N_4217);
nand U4474 (N_4474,N_4210,N_4221);
nor U4475 (N_4475,N_4235,N_4229);
xor U4476 (N_4476,N_4207,N_4254);
nand U4477 (N_4477,N_4312,N_4222);
and U4478 (N_4478,N_4291,N_4370);
or U4479 (N_4479,N_4346,N_4398);
nand U4480 (N_4480,N_4295,N_4377);
or U4481 (N_4481,N_4251,N_4343);
and U4482 (N_4482,N_4357,N_4213);
or U4483 (N_4483,N_4349,N_4333);
nor U4484 (N_4484,N_4263,N_4273);
xor U4485 (N_4485,N_4355,N_4231);
xor U4486 (N_4486,N_4379,N_4293);
and U4487 (N_4487,N_4320,N_4323);
or U4488 (N_4488,N_4329,N_4384);
xnor U4489 (N_4489,N_4269,N_4279);
nand U4490 (N_4490,N_4317,N_4305);
and U4491 (N_4491,N_4344,N_4226);
nor U4492 (N_4492,N_4321,N_4313);
nand U4493 (N_4493,N_4227,N_4381);
or U4494 (N_4494,N_4374,N_4204);
or U4495 (N_4495,N_4267,N_4340);
nor U4496 (N_4496,N_4328,N_4234);
xor U4497 (N_4497,N_4249,N_4368);
nor U4498 (N_4498,N_4264,N_4292);
xnor U4499 (N_4499,N_4365,N_4308);
nand U4500 (N_4500,N_4278,N_4283);
xor U4501 (N_4501,N_4303,N_4384);
xor U4502 (N_4502,N_4251,N_4305);
and U4503 (N_4503,N_4249,N_4211);
nor U4504 (N_4504,N_4274,N_4384);
or U4505 (N_4505,N_4246,N_4316);
and U4506 (N_4506,N_4323,N_4381);
xor U4507 (N_4507,N_4221,N_4249);
xor U4508 (N_4508,N_4265,N_4211);
nor U4509 (N_4509,N_4362,N_4391);
or U4510 (N_4510,N_4370,N_4232);
xor U4511 (N_4511,N_4246,N_4345);
nand U4512 (N_4512,N_4360,N_4291);
or U4513 (N_4513,N_4269,N_4212);
nand U4514 (N_4514,N_4309,N_4329);
xnor U4515 (N_4515,N_4225,N_4341);
xnor U4516 (N_4516,N_4309,N_4210);
and U4517 (N_4517,N_4353,N_4343);
and U4518 (N_4518,N_4250,N_4237);
nor U4519 (N_4519,N_4275,N_4287);
nor U4520 (N_4520,N_4288,N_4314);
or U4521 (N_4521,N_4354,N_4370);
and U4522 (N_4522,N_4274,N_4288);
nor U4523 (N_4523,N_4228,N_4239);
nor U4524 (N_4524,N_4397,N_4288);
or U4525 (N_4525,N_4285,N_4397);
and U4526 (N_4526,N_4344,N_4217);
and U4527 (N_4527,N_4241,N_4265);
or U4528 (N_4528,N_4307,N_4206);
nand U4529 (N_4529,N_4321,N_4253);
nand U4530 (N_4530,N_4283,N_4335);
nand U4531 (N_4531,N_4252,N_4200);
nor U4532 (N_4532,N_4340,N_4318);
or U4533 (N_4533,N_4353,N_4360);
or U4534 (N_4534,N_4202,N_4365);
or U4535 (N_4535,N_4278,N_4330);
nor U4536 (N_4536,N_4347,N_4221);
or U4537 (N_4537,N_4250,N_4214);
nor U4538 (N_4538,N_4295,N_4358);
nand U4539 (N_4539,N_4230,N_4262);
xor U4540 (N_4540,N_4345,N_4307);
nand U4541 (N_4541,N_4215,N_4240);
xor U4542 (N_4542,N_4228,N_4256);
xnor U4543 (N_4543,N_4213,N_4236);
xor U4544 (N_4544,N_4312,N_4347);
and U4545 (N_4545,N_4261,N_4324);
nand U4546 (N_4546,N_4364,N_4397);
and U4547 (N_4547,N_4252,N_4242);
or U4548 (N_4548,N_4349,N_4375);
and U4549 (N_4549,N_4245,N_4227);
nand U4550 (N_4550,N_4332,N_4299);
nor U4551 (N_4551,N_4210,N_4326);
nor U4552 (N_4552,N_4289,N_4242);
xor U4553 (N_4553,N_4382,N_4233);
or U4554 (N_4554,N_4319,N_4323);
or U4555 (N_4555,N_4284,N_4363);
nand U4556 (N_4556,N_4221,N_4398);
or U4557 (N_4557,N_4232,N_4369);
nor U4558 (N_4558,N_4389,N_4255);
xor U4559 (N_4559,N_4369,N_4283);
nor U4560 (N_4560,N_4384,N_4304);
or U4561 (N_4561,N_4363,N_4289);
xor U4562 (N_4562,N_4300,N_4209);
xnor U4563 (N_4563,N_4351,N_4207);
nor U4564 (N_4564,N_4310,N_4277);
and U4565 (N_4565,N_4277,N_4390);
xor U4566 (N_4566,N_4251,N_4344);
nand U4567 (N_4567,N_4236,N_4381);
nor U4568 (N_4568,N_4371,N_4364);
or U4569 (N_4569,N_4280,N_4254);
and U4570 (N_4570,N_4269,N_4222);
nand U4571 (N_4571,N_4226,N_4278);
xor U4572 (N_4572,N_4372,N_4356);
nor U4573 (N_4573,N_4393,N_4262);
nor U4574 (N_4574,N_4261,N_4336);
nand U4575 (N_4575,N_4285,N_4395);
nand U4576 (N_4576,N_4363,N_4261);
and U4577 (N_4577,N_4243,N_4351);
nor U4578 (N_4578,N_4222,N_4226);
or U4579 (N_4579,N_4222,N_4274);
and U4580 (N_4580,N_4308,N_4360);
xor U4581 (N_4581,N_4399,N_4321);
nand U4582 (N_4582,N_4291,N_4387);
nor U4583 (N_4583,N_4389,N_4291);
or U4584 (N_4584,N_4270,N_4343);
xnor U4585 (N_4585,N_4220,N_4207);
nand U4586 (N_4586,N_4276,N_4368);
xor U4587 (N_4587,N_4250,N_4391);
nor U4588 (N_4588,N_4372,N_4231);
nor U4589 (N_4589,N_4201,N_4266);
xor U4590 (N_4590,N_4294,N_4324);
nor U4591 (N_4591,N_4385,N_4222);
nor U4592 (N_4592,N_4323,N_4372);
nor U4593 (N_4593,N_4388,N_4237);
nor U4594 (N_4594,N_4371,N_4277);
nor U4595 (N_4595,N_4261,N_4271);
or U4596 (N_4596,N_4254,N_4261);
xor U4597 (N_4597,N_4270,N_4282);
or U4598 (N_4598,N_4223,N_4376);
and U4599 (N_4599,N_4380,N_4336);
nor U4600 (N_4600,N_4468,N_4495);
and U4601 (N_4601,N_4485,N_4409);
or U4602 (N_4602,N_4505,N_4474);
nor U4603 (N_4603,N_4530,N_4430);
and U4604 (N_4604,N_4547,N_4550);
and U4605 (N_4605,N_4467,N_4540);
and U4606 (N_4606,N_4515,N_4438);
and U4607 (N_4607,N_4426,N_4479);
xor U4608 (N_4608,N_4507,N_4434);
nor U4609 (N_4609,N_4439,N_4535);
and U4610 (N_4610,N_4444,N_4517);
or U4611 (N_4611,N_4597,N_4504);
xor U4612 (N_4612,N_4579,N_4451);
nor U4613 (N_4613,N_4522,N_4442);
and U4614 (N_4614,N_4556,N_4538);
or U4615 (N_4615,N_4454,N_4459);
and U4616 (N_4616,N_4576,N_4491);
nand U4617 (N_4617,N_4445,N_4494);
and U4618 (N_4618,N_4584,N_4411);
or U4619 (N_4619,N_4518,N_4562);
xnor U4620 (N_4620,N_4524,N_4588);
nor U4621 (N_4621,N_4460,N_4493);
and U4622 (N_4622,N_4596,N_4432);
xnor U4623 (N_4623,N_4441,N_4574);
xor U4624 (N_4624,N_4590,N_4404);
or U4625 (N_4625,N_4589,N_4570);
or U4626 (N_4626,N_4553,N_4421);
or U4627 (N_4627,N_4528,N_4497);
or U4628 (N_4628,N_4583,N_4422);
xnor U4629 (N_4629,N_4448,N_4400);
xnor U4630 (N_4630,N_4465,N_4566);
nor U4631 (N_4631,N_4402,N_4527);
or U4632 (N_4632,N_4464,N_4561);
nand U4633 (N_4633,N_4471,N_4489);
nand U4634 (N_4634,N_4514,N_4548);
and U4635 (N_4635,N_4578,N_4593);
nor U4636 (N_4636,N_4539,N_4506);
and U4637 (N_4637,N_4551,N_4473);
xnor U4638 (N_4638,N_4478,N_4557);
nor U4639 (N_4639,N_4418,N_4552);
and U4640 (N_4640,N_4568,N_4487);
or U4641 (N_4641,N_4424,N_4536);
and U4642 (N_4642,N_4427,N_4577);
or U4643 (N_4643,N_4449,N_4499);
nor U4644 (N_4644,N_4521,N_4523);
or U4645 (N_4645,N_4470,N_4525);
nor U4646 (N_4646,N_4598,N_4433);
or U4647 (N_4647,N_4435,N_4575);
xnor U4648 (N_4648,N_4437,N_4549);
or U4649 (N_4649,N_4476,N_4417);
nand U4650 (N_4650,N_4520,N_4469);
and U4651 (N_4651,N_4516,N_4453);
or U4652 (N_4652,N_4452,N_4484);
or U4653 (N_4653,N_4581,N_4455);
and U4654 (N_4654,N_4486,N_4554);
nand U4655 (N_4655,N_4429,N_4480);
nand U4656 (N_4656,N_4563,N_4415);
nand U4657 (N_4657,N_4545,N_4475);
nand U4658 (N_4658,N_4501,N_4423);
or U4659 (N_4659,N_4477,N_4502);
or U4660 (N_4660,N_4412,N_4447);
xnor U4661 (N_4661,N_4463,N_4407);
or U4662 (N_4662,N_4503,N_4466);
xor U4663 (N_4663,N_4414,N_4537);
xor U4664 (N_4664,N_4496,N_4595);
and U4665 (N_4665,N_4519,N_4458);
or U4666 (N_4666,N_4416,N_4567);
nor U4667 (N_4667,N_4419,N_4559);
nor U4668 (N_4668,N_4587,N_4532);
xnor U4669 (N_4669,N_4436,N_4586);
or U4670 (N_4670,N_4420,N_4462);
xor U4671 (N_4671,N_4443,N_4599);
nor U4672 (N_4672,N_4513,N_4500);
nand U4673 (N_4673,N_4572,N_4582);
xnor U4674 (N_4674,N_4533,N_4403);
xnor U4675 (N_4675,N_4565,N_4406);
nand U4676 (N_4676,N_4425,N_4543);
xnor U4677 (N_4677,N_4405,N_4541);
nor U4678 (N_4678,N_4510,N_4401);
nand U4679 (N_4679,N_4591,N_4534);
nor U4680 (N_4680,N_4457,N_4555);
nand U4681 (N_4681,N_4529,N_4490);
and U4682 (N_4682,N_4526,N_4488);
nor U4683 (N_4683,N_4580,N_4450);
xor U4684 (N_4684,N_4410,N_4571);
and U4685 (N_4685,N_4511,N_4512);
nand U4686 (N_4686,N_4508,N_4542);
nor U4687 (N_4687,N_4592,N_4456);
and U4688 (N_4688,N_4569,N_4413);
nand U4689 (N_4689,N_4558,N_4546);
or U4690 (N_4690,N_4472,N_4461);
and U4691 (N_4691,N_4531,N_4492);
and U4692 (N_4692,N_4594,N_4483);
and U4693 (N_4693,N_4573,N_4481);
and U4694 (N_4694,N_4431,N_4428);
xor U4695 (N_4695,N_4509,N_4446);
and U4696 (N_4696,N_4560,N_4440);
nor U4697 (N_4697,N_4585,N_4408);
or U4698 (N_4698,N_4544,N_4498);
and U4699 (N_4699,N_4564,N_4482);
or U4700 (N_4700,N_4425,N_4453);
and U4701 (N_4701,N_4495,N_4474);
nor U4702 (N_4702,N_4532,N_4549);
nand U4703 (N_4703,N_4581,N_4461);
nand U4704 (N_4704,N_4496,N_4431);
xor U4705 (N_4705,N_4543,N_4542);
nand U4706 (N_4706,N_4466,N_4485);
nand U4707 (N_4707,N_4510,N_4576);
or U4708 (N_4708,N_4412,N_4522);
xnor U4709 (N_4709,N_4563,N_4566);
or U4710 (N_4710,N_4528,N_4571);
and U4711 (N_4711,N_4441,N_4517);
or U4712 (N_4712,N_4493,N_4534);
or U4713 (N_4713,N_4430,N_4447);
xor U4714 (N_4714,N_4564,N_4459);
nand U4715 (N_4715,N_4572,N_4437);
or U4716 (N_4716,N_4567,N_4593);
or U4717 (N_4717,N_4509,N_4447);
and U4718 (N_4718,N_4583,N_4539);
or U4719 (N_4719,N_4572,N_4555);
xor U4720 (N_4720,N_4573,N_4469);
and U4721 (N_4721,N_4446,N_4536);
nor U4722 (N_4722,N_4533,N_4418);
nand U4723 (N_4723,N_4595,N_4472);
or U4724 (N_4724,N_4483,N_4497);
nor U4725 (N_4725,N_4527,N_4543);
and U4726 (N_4726,N_4465,N_4436);
nor U4727 (N_4727,N_4451,N_4495);
and U4728 (N_4728,N_4477,N_4521);
and U4729 (N_4729,N_4528,N_4471);
and U4730 (N_4730,N_4404,N_4435);
or U4731 (N_4731,N_4568,N_4566);
nor U4732 (N_4732,N_4530,N_4437);
and U4733 (N_4733,N_4405,N_4558);
nand U4734 (N_4734,N_4533,N_4508);
nor U4735 (N_4735,N_4569,N_4567);
or U4736 (N_4736,N_4482,N_4474);
and U4737 (N_4737,N_4589,N_4564);
nor U4738 (N_4738,N_4466,N_4464);
xnor U4739 (N_4739,N_4577,N_4448);
and U4740 (N_4740,N_4574,N_4531);
or U4741 (N_4741,N_4502,N_4561);
xor U4742 (N_4742,N_4438,N_4415);
nand U4743 (N_4743,N_4517,N_4481);
nor U4744 (N_4744,N_4503,N_4570);
nand U4745 (N_4745,N_4569,N_4417);
or U4746 (N_4746,N_4559,N_4583);
nand U4747 (N_4747,N_4587,N_4518);
or U4748 (N_4748,N_4553,N_4526);
nor U4749 (N_4749,N_4513,N_4424);
nand U4750 (N_4750,N_4423,N_4459);
xnor U4751 (N_4751,N_4540,N_4542);
and U4752 (N_4752,N_4540,N_4476);
xnor U4753 (N_4753,N_4415,N_4453);
and U4754 (N_4754,N_4584,N_4599);
xnor U4755 (N_4755,N_4544,N_4451);
nand U4756 (N_4756,N_4468,N_4492);
xnor U4757 (N_4757,N_4476,N_4429);
xor U4758 (N_4758,N_4585,N_4507);
or U4759 (N_4759,N_4588,N_4523);
and U4760 (N_4760,N_4546,N_4511);
nor U4761 (N_4761,N_4574,N_4533);
and U4762 (N_4762,N_4527,N_4500);
or U4763 (N_4763,N_4464,N_4590);
or U4764 (N_4764,N_4422,N_4573);
or U4765 (N_4765,N_4566,N_4580);
and U4766 (N_4766,N_4420,N_4526);
or U4767 (N_4767,N_4558,N_4409);
nand U4768 (N_4768,N_4466,N_4454);
nand U4769 (N_4769,N_4561,N_4406);
and U4770 (N_4770,N_4522,N_4549);
or U4771 (N_4771,N_4577,N_4419);
or U4772 (N_4772,N_4566,N_4457);
and U4773 (N_4773,N_4496,N_4531);
nor U4774 (N_4774,N_4553,N_4541);
or U4775 (N_4775,N_4561,N_4549);
and U4776 (N_4776,N_4421,N_4499);
nand U4777 (N_4777,N_4408,N_4492);
nor U4778 (N_4778,N_4533,N_4419);
and U4779 (N_4779,N_4471,N_4588);
nand U4780 (N_4780,N_4581,N_4570);
xor U4781 (N_4781,N_4486,N_4588);
and U4782 (N_4782,N_4471,N_4590);
or U4783 (N_4783,N_4431,N_4487);
or U4784 (N_4784,N_4470,N_4496);
nor U4785 (N_4785,N_4557,N_4509);
nor U4786 (N_4786,N_4418,N_4577);
nand U4787 (N_4787,N_4490,N_4566);
nor U4788 (N_4788,N_4486,N_4522);
xor U4789 (N_4789,N_4490,N_4570);
and U4790 (N_4790,N_4487,N_4409);
nor U4791 (N_4791,N_4419,N_4441);
nor U4792 (N_4792,N_4401,N_4536);
nor U4793 (N_4793,N_4587,N_4410);
xor U4794 (N_4794,N_4424,N_4505);
nand U4795 (N_4795,N_4543,N_4405);
nand U4796 (N_4796,N_4550,N_4468);
xor U4797 (N_4797,N_4502,N_4447);
and U4798 (N_4798,N_4520,N_4526);
xor U4799 (N_4799,N_4502,N_4480);
nand U4800 (N_4800,N_4789,N_4676);
nor U4801 (N_4801,N_4716,N_4626);
nor U4802 (N_4802,N_4675,N_4639);
xnor U4803 (N_4803,N_4660,N_4745);
xnor U4804 (N_4804,N_4774,N_4711);
and U4805 (N_4805,N_4667,N_4687);
nand U4806 (N_4806,N_4738,N_4621);
and U4807 (N_4807,N_4693,N_4771);
xor U4808 (N_4808,N_4627,N_4638);
nor U4809 (N_4809,N_4733,N_4763);
and U4810 (N_4810,N_4723,N_4715);
and U4811 (N_4811,N_4632,N_4788);
nor U4812 (N_4812,N_4799,N_4757);
or U4813 (N_4813,N_4739,N_4682);
xor U4814 (N_4814,N_4721,N_4790);
xnor U4815 (N_4815,N_4641,N_4755);
nor U4816 (N_4816,N_4686,N_4635);
xnor U4817 (N_4817,N_4615,N_4713);
xnor U4818 (N_4818,N_4701,N_4668);
nand U4819 (N_4819,N_4724,N_4764);
and U4820 (N_4820,N_4732,N_4729);
nor U4821 (N_4821,N_4749,N_4797);
xor U4822 (N_4822,N_4703,N_4760);
nand U4823 (N_4823,N_4636,N_4623);
nor U4824 (N_4824,N_4658,N_4787);
and U4825 (N_4825,N_4700,N_4674);
xor U4826 (N_4826,N_4785,N_4718);
nand U4827 (N_4827,N_4734,N_4654);
and U4828 (N_4828,N_4694,N_4720);
nor U4829 (N_4829,N_4747,N_4756);
and U4830 (N_4830,N_4746,N_4618);
or U4831 (N_4831,N_4620,N_4696);
and U4832 (N_4832,N_4689,N_4792);
nor U4833 (N_4833,N_4672,N_4791);
nand U4834 (N_4834,N_4653,N_4614);
or U4835 (N_4835,N_4648,N_4657);
and U4836 (N_4836,N_4731,N_4619);
and U4837 (N_4837,N_4735,N_4697);
xnor U4838 (N_4838,N_4767,N_4656);
and U4839 (N_4839,N_4659,N_4690);
nand U4840 (N_4840,N_4795,N_4630);
xor U4841 (N_4841,N_4766,N_4642);
xnor U4842 (N_4842,N_4714,N_4742);
or U4843 (N_4843,N_4691,N_4605);
xnor U4844 (N_4844,N_4768,N_4751);
or U4845 (N_4845,N_4706,N_4699);
xnor U4846 (N_4846,N_4611,N_4727);
and U4847 (N_4847,N_4683,N_4625);
nor U4848 (N_4848,N_4779,N_4728);
nor U4849 (N_4849,N_4786,N_4695);
nand U4850 (N_4850,N_4651,N_4707);
xor U4851 (N_4851,N_4750,N_4784);
or U4852 (N_4852,N_4730,N_4783);
xnor U4853 (N_4853,N_4773,N_4743);
nand U4854 (N_4854,N_4705,N_4796);
nor U4855 (N_4855,N_4669,N_4606);
and U4856 (N_4856,N_4617,N_4794);
nand U4857 (N_4857,N_4652,N_4793);
nor U4858 (N_4858,N_4765,N_4717);
nand U4859 (N_4859,N_4628,N_4612);
nor U4860 (N_4860,N_4604,N_4744);
nor U4861 (N_4861,N_4702,N_4666);
nand U4862 (N_4862,N_4671,N_4780);
and U4863 (N_4863,N_4762,N_4608);
and U4864 (N_4864,N_4778,N_4692);
or U4865 (N_4865,N_4775,N_4709);
xor U4866 (N_4866,N_4631,N_4610);
nand U4867 (N_4867,N_4600,N_4679);
nor U4868 (N_4868,N_4748,N_4722);
nor U4869 (N_4869,N_4754,N_4646);
nand U4870 (N_4870,N_4725,N_4650);
or U4871 (N_4871,N_4673,N_4737);
nand U4872 (N_4872,N_4678,N_4740);
xnor U4873 (N_4873,N_4704,N_4770);
nor U4874 (N_4874,N_4645,N_4640);
and U4875 (N_4875,N_4649,N_4607);
nor U4876 (N_4876,N_4655,N_4634);
and U4877 (N_4877,N_4609,N_4633);
nand U4878 (N_4878,N_4719,N_4664);
and U4879 (N_4879,N_4681,N_4613);
or U4880 (N_4880,N_4684,N_4708);
or U4881 (N_4881,N_4644,N_4753);
and U4882 (N_4882,N_4680,N_4798);
and U4883 (N_4883,N_4759,N_4643);
nand U4884 (N_4884,N_4688,N_4698);
xnor U4885 (N_4885,N_4647,N_4781);
and U4886 (N_4886,N_4670,N_4710);
xor U4887 (N_4887,N_4741,N_4776);
nor U4888 (N_4888,N_4712,N_4663);
nand U4889 (N_4889,N_4622,N_4677);
nor U4890 (N_4890,N_4661,N_4602);
and U4891 (N_4891,N_4782,N_4736);
nand U4892 (N_4892,N_4761,N_4616);
or U4893 (N_4893,N_4601,N_4685);
xnor U4894 (N_4894,N_4772,N_4777);
xnor U4895 (N_4895,N_4624,N_4637);
and U4896 (N_4896,N_4665,N_4752);
and U4897 (N_4897,N_4769,N_4662);
and U4898 (N_4898,N_4758,N_4629);
and U4899 (N_4899,N_4603,N_4726);
xnor U4900 (N_4900,N_4611,N_4661);
xnor U4901 (N_4901,N_4612,N_4690);
xnor U4902 (N_4902,N_4680,N_4659);
and U4903 (N_4903,N_4655,N_4642);
and U4904 (N_4904,N_4697,N_4673);
or U4905 (N_4905,N_4793,N_4762);
xor U4906 (N_4906,N_4650,N_4773);
xor U4907 (N_4907,N_4749,N_4704);
xnor U4908 (N_4908,N_4677,N_4730);
nor U4909 (N_4909,N_4748,N_4686);
nand U4910 (N_4910,N_4652,N_4770);
nand U4911 (N_4911,N_4648,N_4741);
nor U4912 (N_4912,N_4670,N_4742);
nor U4913 (N_4913,N_4681,N_4607);
nor U4914 (N_4914,N_4659,N_4753);
nand U4915 (N_4915,N_4778,N_4707);
nor U4916 (N_4916,N_4605,N_4656);
nand U4917 (N_4917,N_4749,N_4700);
nor U4918 (N_4918,N_4605,N_4741);
nand U4919 (N_4919,N_4654,N_4742);
xor U4920 (N_4920,N_4679,N_4609);
and U4921 (N_4921,N_4716,N_4732);
nor U4922 (N_4922,N_4730,N_4695);
xor U4923 (N_4923,N_4624,N_4634);
nand U4924 (N_4924,N_4735,N_4722);
nor U4925 (N_4925,N_4622,N_4646);
or U4926 (N_4926,N_4600,N_4650);
nand U4927 (N_4927,N_4649,N_4708);
or U4928 (N_4928,N_4799,N_4745);
and U4929 (N_4929,N_4610,N_4705);
or U4930 (N_4930,N_4601,N_4650);
or U4931 (N_4931,N_4702,N_4676);
xnor U4932 (N_4932,N_4624,N_4726);
xnor U4933 (N_4933,N_4609,N_4739);
nand U4934 (N_4934,N_4696,N_4704);
nor U4935 (N_4935,N_4762,N_4767);
xor U4936 (N_4936,N_4760,N_4734);
and U4937 (N_4937,N_4741,N_4736);
xor U4938 (N_4938,N_4622,N_4674);
xor U4939 (N_4939,N_4759,N_4762);
nor U4940 (N_4940,N_4791,N_4660);
nor U4941 (N_4941,N_4798,N_4632);
or U4942 (N_4942,N_4731,N_4772);
nor U4943 (N_4943,N_4663,N_4623);
nand U4944 (N_4944,N_4731,N_4696);
nor U4945 (N_4945,N_4741,N_4608);
nand U4946 (N_4946,N_4653,N_4602);
nand U4947 (N_4947,N_4773,N_4748);
nor U4948 (N_4948,N_4717,N_4649);
xor U4949 (N_4949,N_4654,N_4700);
nor U4950 (N_4950,N_4725,N_4695);
or U4951 (N_4951,N_4635,N_4701);
and U4952 (N_4952,N_4747,N_4770);
nor U4953 (N_4953,N_4706,N_4658);
nand U4954 (N_4954,N_4767,N_4634);
nand U4955 (N_4955,N_4793,N_4632);
nor U4956 (N_4956,N_4718,N_4780);
or U4957 (N_4957,N_4683,N_4778);
or U4958 (N_4958,N_4678,N_4682);
and U4959 (N_4959,N_4796,N_4665);
and U4960 (N_4960,N_4669,N_4726);
or U4961 (N_4961,N_4710,N_4734);
nand U4962 (N_4962,N_4613,N_4733);
or U4963 (N_4963,N_4651,N_4770);
nor U4964 (N_4964,N_4662,N_4768);
nand U4965 (N_4965,N_4619,N_4770);
nand U4966 (N_4966,N_4711,N_4754);
and U4967 (N_4967,N_4741,N_4712);
xnor U4968 (N_4968,N_4728,N_4714);
nor U4969 (N_4969,N_4637,N_4775);
xnor U4970 (N_4970,N_4737,N_4629);
nand U4971 (N_4971,N_4782,N_4772);
and U4972 (N_4972,N_4794,N_4783);
nor U4973 (N_4973,N_4750,N_4666);
nor U4974 (N_4974,N_4668,N_4631);
nand U4975 (N_4975,N_4669,N_4764);
nand U4976 (N_4976,N_4778,N_4741);
xor U4977 (N_4977,N_4630,N_4794);
and U4978 (N_4978,N_4619,N_4777);
and U4979 (N_4979,N_4707,N_4722);
and U4980 (N_4980,N_4754,N_4793);
or U4981 (N_4981,N_4608,N_4656);
and U4982 (N_4982,N_4687,N_4675);
nand U4983 (N_4983,N_4641,N_4685);
nand U4984 (N_4984,N_4759,N_4607);
or U4985 (N_4985,N_4781,N_4778);
nor U4986 (N_4986,N_4748,N_4689);
and U4987 (N_4987,N_4689,N_4683);
xor U4988 (N_4988,N_4775,N_4741);
nand U4989 (N_4989,N_4754,N_4760);
nand U4990 (N_4990,N_4767,N_4626);
and U4991 (N_4991,N_4720,N_4602);
nand U4992 (N_4992,N_4705,N_4618);
nor U4993 (N_4993,N_4784,N_4672);
xnor U4994 (N_4994,N_4765,N_4631);
or U4995 (N_4995,N_4632,N_4639);
nor U4996 (N_4996,N_4705,N_4640);
nor U4997 (N_4997,N_4733,N_4649);
and U4998 (N_4998,N_4674,N_4792);
nor U4999 (N_4999,N_4625,N_4752);
xor U5000 (N_5000,N_4926,N_4958);
nand U5001 (N_5001,N_4876,N_4910);
nor U5002 (N_5002,N_4839,N_4811);
xor U5003 (N_5003,N_4827,N_4945);
xor U5004 (N_5004,N_4805,N_4814);
xor U5005 (N_5005,N_4897,N_4823);
nor U5006 (N_5006,N_4912,N_4903);
nand U5007 (N_5007,N_4937,N_4930);
nor U5008 (N_5008,N_4806,N_4851);
nor U5009 (N_5009,N_4885,N_4880);
nor U5010 (N_5010,N_4883,N_4801);
and U5011 (N_5011,N_4884,N_4950);
or U5012 (N_5012,N_4855,N_4964);
nor U5013 (N_5013,N_4981,N_4828);
or U5014 (N_5014,N_4970,N_4902);
nor U5015 (N_5015,N_4918,N_4800);
and U5016 (N_5016,N_4980,N_4860);
or U5017 (N_5017,N_4908,N_4988);
xor U5018 (N_5018,N_4810,N_4931);
and U5019 (N_5019,N_4871,N_4946);
nand U5020 (N_5020,N_4812,N_4972);
nand U5021 (N_5021,N_4909,N_4922);
xor U5022 (N_5022,N_4889,N_4847);
and U5023 (N_5023,N_4953,N_4863);
and U5024 (N_5024,N_4968,N_4916);
nand U5025 (N_5025,N_4923,N_4928);
or U5026 (N_5026,N_4874,N_4818);
nand U5027 (N_5027,N_4940,N_4804);
nor U5028 (N_5028,N_4987,N_4846);
nor U5029 (N_5029,N_4878,N_4997);
xor U5030 (N_5030,N_4813,N_4948);
xor U5031 (N_5031,N_4963,N_4886);
nand U5032 (N_5032,N_4951,N_4919);
xor U5033 (N_5033,N_4973,N_4906);
nand U5034 (N_5034,N_4840,N_4891);
nand U5035 (N_5035,N_4843,N_4947);
or U5036 (N_5036,N_4977,N_4957);
or U5037 (N_5037,N_4830,N_4857);
nor U5038 (N_5038,N_4899,N_4868);
and U5039 (N_5039,N_4821,N_4954);
xor U5040 (N_5040,N_4925,N_4905);
nor U5041 (N_5041,N_4959,N_4960);
or U5042 (N_5042,N_4861,N_4802);
or U5043 (N_5043,N_4869,N_4845);
nand U5044 (N_5044,N_4835,N_4882);
nand U5045 (N_5045,N_4849,N_4978);
nand U5046 (N_5046,N_4924,N_4894);
nor U5047 (N_5047,N_4854,N_4865);
or U5048 (N_5048,N_4967,N_4850);
xnor U5049 (N_5049,N_4842,N_4979);
or U5050 (N_5050,N_4832,N_4862);
nor U5051 (N_5051,N_4971,N_4826);
xnor U5052 (N_5052,N_4819,N_4833);
nor U5053 (N_5053,N_4962,N_4927);
or U5054 (N_5054,N_4848,N_4994);
or U5055 (N_5055,N_4838,N_4983);
nor U5056 (N_5056,N_4870,N_4895);
and U5057 (N_5057,N_4932,N_4866);
nand U5058 (N_5058,N_4935,N_4993);
and U5059 (N_5059,N_4995,N_4991);
and U5060 (N_5060,N_4820,N_4888);
xnor U5061 (N_5061,N_4803,N_4969);
nor U5062 (N_5062,N_4816,N_4952);
nor U5063 (N_5063,N_4896,N_4873);
nor U5064 (N_5064,N_4900,N_4809);
nor U5065 (N_5065,N_4966,N_4841);
nand U5066 (N_5066,N_4893,N_4859);
xor U5067 (N_5067,N_4929,N_4834);
nand U5068 (N_5068,N_4877,N_4998);
or U5069 (N_5069,N_4934,N_4907);
xor U5070 (N_5070,N_4824,N_4949);
xor U5071 (N_5071,N_4999,N_4996);
and U5072 (N_5072,N_4887,N_4892);
or U5073 (N_5073,N_4990,N_4875);
or U5074 (N_5074,N_4941,N_4881);
and U5075 (N_5075,N_4879,N_4984);
or U5076 (N_5076,N_4982,N_4808);
xor U5077 (N_5077,N_4939,N_4975);
nand U5078 (N_5078,N_4852,N_4933);
nor U5079 (N_5079,N_4974,N_4858);
and U5080 (N_5080,N_4901,N_4822);
and U5081 (N_5081,N_4936,N_4965);
nand U5082 (N_5082,N_4917,N_4829);
xnor U5083 (N_5083,N_4921,N_4844);
nand U5084 (N_5084,N_4986,N_4943);
nor U5085 (N_5085,N_4992,N_4898);
and U5086 (N_5086,N_4904,N_4837);
nand U5087 (N_5087,N_4961,N_4864);
nand U5088 (N_5088,N_4867,N_4911);
xnor U5089 (N_5089,N_4914,N_4944);
or U5090 (N_5090,N_4836,N_4890);
or U5091 (N_5091,N_4831,N_4853);
and U5092 (N_5092,N_4938,N_4807);
nor U5093 (N_5093,N_4817,N_4856);
xnor U5094 (N_5094,N_4956,N_4976);
nor U5095 (N_5095,N_4985,N_4915);
and U5096 (N_5096,N_4815,N_4920);
nor U5097 (N_5097,N_4825,N_4942);
nand U5098 (N_5098,N_4955,N_4872);
xnor U5099 (N_5099,N_4913,N_4989);
nor U5100 (N_5100,N_4943,N_4833);
and U5101 (N_5101,N_4810,N_4952);
nand U5102 (N_5102,N_4909,N_4864);
or U5103 (N_5103,N_4921,N_4992);
nor U5104 (N_5104,N_4985,N_4979);
or U5105 (N_5105,N_4952,N_4849);
nand U5106 (N_5106,N_4912,N_4810);
xor U5107 (N_5107,N_4998,N_4869);
nor U5108 (N_5108,N_4956,N_4870);
and U5109 (N_5109,N_4879,N_4961);
nor U5110 (N_5110,N_4921,N_4954);
and U5111 (N_5111,N_4989,N_4901);
or U5112 (N_5112,N_4812,N_4892);
and U5113 (N_5113,N_4892,N_4811);
nand U5114 (N_5114,N_4810,N_4934);
or U5115 (N_5115,N_4909,N_4990);
nor U5116 (N_5116,N_4919,N_4926);
and U5117 (N_5117,N_4818,N_4944);
and U5118 (N_5118,N_4910,N_4967);
and U5119 (N_5119,N_4854,N_4828);
and U5120 (N_5120,N_4892,N_4925);
nor U5121 (N_5121,N_4958,N_4881);
or U5122 (N_5122,N_4989,N_4835);
or U5123 (N_5123,N_4892,N_4870);
and U5124 (N_5124,N_4844,N_4938);
nand U5125 (N_5125,N_4834,N_4985);
nand U5126 (N_5126,N_4859,N_4868);
nand U5127 (N_5127,N_4981,N_4894);
and U5128 (N_5128,N_4808,N_4905);
nand U5129 (N_5129,N_4922,N_4941);
or U5130 (N_5130,N_4829,N_4876);
nor U5131 (N_5131,N_4831,N_4874);
or U5132 (N_5132,N_4838,N_4853);
nand U5133 (N_5133,N_4901,N_4903);
nand U5134 (N_5134,N_4925,N_4819);
nor U5135 (N_5135,N_4978,N_4953);
and U5136 (N_5136,N_4991,N_4892);
xor U5137 (N_5137,N_4835,N_4957);
nor U5138 (N_5138,N_4814,N_4943);
nand U5139 (N_5139,N_4823,N_4962);
nor U5140 (N_5140,N_4867,N_4848);
and U5141 (N_5141,N_4855,N_4896);
and U5142 (N_5142,N_4894,N_4897);
or U5143 (N_5143,N_4992,N_4887);
nand U5144 (N_5144,N_4920,N_4824);
or U5145 (N_5145,N_4981,N_4810);
nor U5146 (N_5146,N_4969,N_4927);
nor U5147 (N_5147,N_4852,N_4844);
nand U5148 (N_5148,N_4852,N_4872);
nand U5149 (N_5149,N_4933,N_4909);
and U5150 (N_5150,N_4828,N_4886);
and U5151 (N_5151,N_4978,N_4811);
or U5152 (N_5152,N_4949,N_4979);
xor U5153 (N_5153,N_4825,N_4914);
and U5154 (N_5154,N_4817,N_4893);
nor U5155 (N_5155,N_4943,N_4825);
nand U5156 (N_5156,N_4941,N_4952);
or U5157 (N_5157,N_4827,N_4801);
and U5158 (N_5158,N_4854,N_4856);
and U5159 (N_5159,N_4886,N_4949);
nand U5160 (N_5160,N_4897,N_4926);
xor U5161 (N_5161,N_4858,N_4904);
or U5162 (N_5162,N_4969,N_4866);
or U5163 (N_5163,N_4951,N_4920);
and U5164 (N_5164,N_4946,N_4863);
and U5165 (N_5165,N_4986,N_4848);
nor U5166 (N_5166,N_4852,N_4960);
nor U5167 (N_5167,N_4852,N_4953);
xnor U5168 (N_5168,N_4849,N_4801);
xor U5169 (N_5169,N_4883,N_4827);
nand U5170 (N_5170,N_4881,N_4888);
or U5171 (N_5171,N_4981,N_4888);
xor U5172 (N_5172,N_4955,N_4982);
xnor U5173 (N_5173,N_4854,N_4972);
or U5174 (N_5174,N_4947,N_4948);
nand U5175 (N_5175,N_4820,N_4985);
nand U5176 (N_5176,N_4852,N_4848);
xor U5177 (N_5177,N_4921,N_4922);
and U5178 (N_5178,N_4902,N_4952);
nand U5179 (N_5179,N_4878,N_4922);
and U5180 (N_5180,N_4871,N_4823);
nand U5181 (N_5181,N_4839,N_4848);
or U5182 (N_5182,N_4961,N_4959);
nor U5183 (N_5183,N_4899,N_4805);
xor U5184 (N_5184,N_4909,N_4960);
and U5185 (N_5185,N_4975,N_4842);
xnor U5186 (N_5186,N_4870,N_4852);
and U5187 (N_5187,N_4988,N_4911);
nor U5188 (N_5188,N_4838,N_4943);
nor U5189 (N_5189,N_4874,N_4825);
nand U5190 (N_5190,N_4833,N_4904);
xor U5191 (N_5191,N_4904,N_4873);
nand U5192 (N_5192,N_4936,N_4861);
xor U5193 (N_5193,N_4887,N_4924);
nand U5194 (N_5194,N_4911,N_4908);
and U5195 (N_5195,N_4879,N_4919);
or U5196 (N_5196,N_4863,N_4835);
and U5197 (N_5197,N_4896,N_4823);
and U5198 (N_5198,N_4990,N_4854);
nor U5199 (N_5199,N_4824,N_4968);
or U5200 (N_5200,N_5068,N_5184);
xor U5201 (N_5201,N_5090,N_5175);
nor U5202 (N_5202,N_5057,N_5069);
or U5203 (N_5203,N_5018,N_5092);
nor U5204 (N_5204,N_5152,N_5136);
nand U5205 (N_5205,N_5168,N_5038);
or U5206 (N_5206,N_5170,N_5169);
xnor U5207 (N_5207,N_5197,N_5122);
nor U5208 (N_5208,N_5005,N_5118);
and U5209 (N_5209,N_5104,N_5107);
xnor U5210 (N_5210,N_5027,N_5139);
nand U5211 (N_5211,N_5129,N_5051);
xnor U5212 (N_5212,N_5185,N_5064);
and U5213 (N_5213,N_5074,N_5199);
or U5214 (N_5214,N_5110,N_5101);
nor U5215 (N_5215,N_5191,N_5126);
nor U5216 (N_5216,N_5077,N_5164);
nand U5217 (N_5217,N_5010,N_5017);
xor U5218 (N_5218,N_5054,N_5020);
xor U5219 (N_5219,N_5148,N_5145);
nand U5220 (N_5220,N_5186,N_5016);
and U5221 (N_5221,N_5040,N_5179);
nor U5222 (N_5222,N_5008,N_5174);
or U5223 (N_5223,N_5082,N_5162);
or U5224 (N_5224,N_5177,N_5056);
or U5225 (N_5225,N_5006,N_5099);
and U5226 (N_5226,N_5131,N_5198);
or U5227 (N_5227,N_5055,N_5161);
nor U5228 (N_5228,N_5045,N_5085);
nand U5229 (N_5229,N_5146,N_5048);
or U5230 (N_5230,N_5115,N_5156);
and U5231 (N_5231,N_5030,N_5111);
and U5232 (N_5232,N_5067,N_5021);
or U5233 (N_5233,N_5154,N_5182);
or U5234 (N_5234,N_5071,N_5044);
nor U5235 (N_5235,N_5142,N_5163);
xor U5236 (N_5236,N_5172,N_5034);
nor U5237 (N_5237,N_5187,N_5060);
nor U5238 (N_5238,N_5087,N_5072);
or U5239 (N_5239,N_5094,N_5171);
and U5240 (N_5240,N_5007,N_5102);
and U5241 (N_5241,N_5108,N_5037);
nand U5242 (N_5242,N_5141,N_5181);
nand U5243 (N_5243,N_5011,N_5091);
and U5244 (N_5244,N_5123,N_5157);
nand U5245 (N_5245,N_5004,N_5003);
or U5246 (N_5246,N_5116,N_5119);
xor U5247 (N_5247,N_5079,N_5046);
and U5248 (N_5248,N_5032,N_5132);
nor U5249 (N_5249,N_5137,N_5150);
nand U5250 (N_5250,N_5023,N_5196);
nand U5251 (N_5251,N_5155,N_5176);
and U5252 (N_5252,N_5124,N_5173);
nor U5253 (N_5253,N_5138,N_5000);
nand U5254 (N_5254,N_5001,N_5167);
xor U5255 (N_5255,N_5042,N_5058);
xor U5256 (N_5256,N_5089,N_5193);
xor U5257 (N_5257,N_5151,N_5097);
and U5258 (N_5258,N_5002,N_5195);
nand U5259 (N_5259,N_5061,N_5066);
nand U5260 (N_5260,N_5052,N_5120);
xor U5261 (N_5261,N_5062,N_5105);
nor U5262 (N_5262,N_5043,N_5117);
nand U5263 (N_5263,N_5028,N_5096);
or U5264 (N_5264,N_5147,N_5047);
nor U5265 (N_5265,N_5053,N_5070);
nor U5266 (N_5266,N_5026,N_5063);
nand U5267 (N_5267,N_5165,N_5153);
xnor U5268 (N_5268,N_5050,N_5113);
nand U5269 (N_5269,N_5081,N_5095);
nand U5270 (N_5270,N_5036,N_5149);
or U5271 (N_5271,N_5029,N_5015);
xor U5272 (N_5272,N_5073,N_5166);
and U5273 (N_5273,N_5121,N_5024);
xnor U5274 (N_5274,N_5013,N_5035);
and U5275 (N_5275,N_5180,N_5178);
and U5276 (N_5276,N_5109,N_5093);
nand U5277 (N_5277,N_5134,N_5049);
nand U5278 (N_5278,N_5088,N_5098);
nor U5279 (N_5279,N_5112,N_5194);
xnor U5280 (N_5280,N_5128,N_5012);
and U5281 (N_5281,N_5133,N_5103);
xnor U5282 (N_5282,N_5183,N_5084);
nor U5283 (N_5283,N_5059,N_5076);
or U5284 (N_5284,N_5159,N_5014);
nand U5285 (N_5285,N_5160,N_5078);
nand U5286 (N_5286,N_5190,N_5031);
or U5287 (N_5287,N_5143,N_5158);
and U5288 (N_5288,N_5075,N_5033);
and U5289 (N_5289,N_5125,N_5009);
nor U5290 (N_5290,N_5106,N_5022);
xnor U5291 (N_5291,N_5189,N_5140);
nor U5292 (N_5292,N_5127,N_5114);
and U5293 (N_5293,N_5025,N_5039);
nand U5294 (N_5294,N_5192,N_5100);
and U5295 (N_5295,N_5086,N_5130);
or U5296 (N_5296,N_5041,N_5019);
nor U5297 (N_5297,N_5065,N_5083);
and U5298 (N_5298,N_5144,N_5135);
nor U5299 (N_5299,N_5080,N_5188);
nor U5300 (N_5300,N_5119,N_5039);
xor U5301 (N_5301,N_5163,N_5053);
or U5302 (N_5302,N_5054,N_5024);
or U5303 (N_5303,N_5160,N_5118);
or U5304 (N_5304,N_5124,N_5089);
and U5305 (N_5305,N_5060,N_5165);
nand U5306 (N_5306,N_5139,N_5182);
xor U5307 (N_5307,N_5120,N_5094);
or U5308 (N_5308,N_5195,N_5045);
nand U5309 (N_5309,N_5038,N_5010);
nand U5310 (N_5310,N_5181,N_5194);
nand U5311 (N_5311,N_5166,N_5120);
or U5312 (N_5312,N_5181,N_5045);
nand U5313 (N_5313,N_5142,N_5012);
nor U5314 (N_5314,N_5065,N_5149);
nand U5315 (N_5315,N_5135,N_5055);
and U5316 (N_5316,N_5083,N_5045);
or U5317 (N_5317,N_5063,N_5097);
nand U5318 (N_5318,N_5068,N_5077);
nor U5319 (N_5319,N_5075,N_5108);
and U5320 (N_5320,N_5024,N_5119);
nand U5321 (N_5321,N_5008,N_5184);
nand U5322 (N_5322,N_5113,N_5179);
and U5323 (N_5323,N_5127,N_5011);
nand U5324 (N_5324,N_5059,N_5146);
and U5325 (N_5325,N_5041,N_5045);
xnor U5326 (N_5326,N_5110,N_5006);
nand U5327 (N_5327,N_5129,N_5180);
nand U5328 (N_5328,N_5057,N_5175);
and U5329 (N_5329,N_5045,N_5081);
nand U5330 (N_5330,N_5140,N_5132);
or U5331 (N_5331,N_5087,N_5075);
nand U5332 (N_5332,N_5102,N_5123);
nand U5333 (N_5333,N_5160,N_5068);
nand U5334 (N_5334,N_5180,N_5010);
xor U5335 (N_5335,N_5190,N_5033);
nand U5336 (N_5336,N_5175,N_5124);
and U5337 (N_5337,N_5129,N_5123);
or U5338 (N_5338,N_5146,N_5115);
and U5339 (N_5339,N_5072,N_5146);
and U5340 (N_5340,N_5018,N_5061);
nand U5341 (N_5341,N_5037,N_5148);
xnor U5342 (N_5342,N_5151,N_5080);
nor U5343 (N_5343,N_5181,N_5174);
nand U5344 (N_5344,N_5034,N_5124);
xor U5345 (N_5345,N_5110,N_5015);
nor U5346 (N_5346,N_5128,N_5004);
xnor U5347 (N_5347,N_5041,N_5082);
nand U5348 (N_5348,N_5142,N_5152);
xor U5349 (N_5349,N_5139,N_5189);
or U5350 (N_5350,N_5059,N_5096);
nand U5351 (N_5351,N_5065,N_5139);
xor U5352 (N_5352,N_5174,N_5146);
nor U5353 (N_5353,N_5196,N_5032);
and U5354 (N_5354,N_5132,N_5165);
or U5355 (N_5355,N_5070,N_5160);
or U5356 (N_5356,N_5087,N_5028);
nor U5357 (N_5357,N_5072,N_5038);
or U5358 (N_5358,N_5188,N_5127);
or U5359 (N_5359,N_5169,N_5023);
nor U5360 (N_5360,N_5033,N_5048);
xor U5361 (N_5361,N_5117,N_5045);
or U5362 (N_5362,N_5141,N_5114);
nand U5363 (N_5363,N_5071,N_5183);
nand U5364 (N_5364,N_5023,N_5093);
or U5365 (N_5365,N_5150,N_5107);
and U5366 (N_5366,N_5102,N_5128);
xor U5367 (N_5367,N_5041,N_5022);
and U5368 (N_5368,N_5030,N_5057);
nor U5369 (N_5369,N_5183,N_5123);
and U5370 (N_5370,N_5162,N_5077);
and U5371 (N_5371,N_5086,N_5005);
nand U5372 (N_5372,N_5074,N_5148);
nor U5373 (N_5373,N_5026,N_5040);
or U5374 (N_5374,N_5123,N_5125);
nor U5375 (N_5375,N_5188,N_5136);
or U5376 (N_5376,N_5171,N_5055);
nand U5377 (N_5377,N_5199,N_5072);
or U5378 (N_5378,N_5041,N_5035);
and U5379 (N_5379,N_5162,N_5165);
nand U5380 (N_5380,N_5020,N_5081);
nor U5381 (N_5381,N_5023,N_5072);
xor U5382 (N_5382,N_5118,N_5125);
and U5383 (N_5383,N_5197,N_5177);
xor U5384 (N_5384,N_5057,N_5028);
nand U5385 (N_5385,N_5140,N_5126);
nor U5386 (N_5386,N_5025,N_5043);
xnor U5387 (N_5387,N_5005,N_5006);
and U5388 (N_5388,N_5032,N_5113);
nand U5389 (N_5389,N_5019,N_5150);
or U5390 (N_5390,N_5096,N_5054);
or U5391 (N_5391,N_5001,N_5015);
xor U5392 (N_5392,N_5005,N_5047);
nand U5393 (N_5393,N_5007,N_5172);
or U5394 (N_5394,N_5041,N_5011);
or U5395 (N_5395,N_5057,N_5039);
or U5396 (N_5396,N_5132,N_5196);
and U5397 (N_5397,N_5093,N_5020);
nor U5398 (N_5398,N_5089,N_5186);
or U5399 (N_5399,N_5024,N_5143);
or U5400 (N_5400,N_5326,N_5239);
and U5401 (N_5401,N_5270,N_5219);
nand U5402 (N_5402,N_5359,N_5381);
and U5403 (N_5403,N_5266,N_5319);
nand U5404 (N_5404,N_5230,N_5389);
xor U5405 (N_5405,N_5399,N_5333);
nand U5406 (N_5406,N_5334,N_5235);
xnor U5407 (N_5407,N_5224,N_5371);
nor U5408 (N_5408,N_5363,N_5383);
xnor U5409 (N_5409,N_5338,N_5375);
and U5410 (N_5410,N_5216,N_5376);
nor U5411 (N_5411,N_5308,N_5227);
nand U5412 (N_5412,N_5233,N_5397);
and U5413 (N_5413,N_5382,N_5264);
or U5414 (N_5414,N_5242,N_5274);
nand U5415 (N_5415,N_5342,N_5365);
nand U5416 (N_5416,N_5206,N_5325);
or U5417 (N_5417,N_5317,N_5355);
xor U5418 (N_5418,N_5335,N_5340);
and U5419 (N_5419,N_5214,N_5241);
and U5420 (N_5420,N_5314,N_5370);
xnor U5421 (N_5421,N_5352,N_5278);
or U5422 (N_5422,N_5294,N_5210);
and U5423 (N_5423,N_5276,N_5395);
or U5424 (N_5424,N_5373,N_5313);
xnor U5425 (N_5425,N_5282,N_5258);
or U5426 (N_5426,N_5257,N_5215);
and U5427 (N_5427,N_5288,N_5372);
xnor U5428 (N_5428,N_5348,N_5318);
xor U5429 (N_5429,N_5267,N_5298);
nor U5430 (N_5430,N_5273,N_5386);
xor U5431 (N_5431,N_5320,N_5240);
and U5432 (N_5432,N_5204,N_5262);
or U5433 (N_5433,N_5337,N_5339);
or U5434 (N_5434,N_5279,N_5329);
xnor U5435 (N_5435,N_5226,N_5377);
and U5436 (N_5436,N_5366,N_5350);
or U5437 (N_5437,N_5272,N_5300);
and U5438 (N_5438,N_5379,N_5302);
or U5439 (N_5439,N_5311,N_5238);
or U5440 (N_5440,N_5292,N_5207);
and U5441 (N_5441,N_5220,N_5346);
or U5442 (N_5442,N_5263,N_5307);
xnor U5443 (N_5443,N_5269,N_5255);
nor U5444 (N_5444,N_5261,N_5286);
or U5445 (N_5445,N_5331,N_5237);
nand U5446 (N_5446,N_5327,N_5232);
nand U5447 (N_5447,N_5354,N_5349);
or U5448 (N_5448,N_5378,N_5396);
xnor U5449 (N_5449,N_5211,N_5218);
nor U5450 (N_5450,N_5243,N_5336);
xnor U5451 (N_5451,N_5205,N_5287);
nor U5452 (N_5452,N_5361,N_5385);
or U5453 (N_5453,N_5347,N_5223);
nor U5454 (N_5454,N_5344,N_5275);
nand U5455 (N_5455,N_5290,N_5222);
nor U5456 (N_5456,N_5203,N_5280);
nand U5457 (N_5457,N_5393,N_5316);
nor U5458 (N_5458,N_5217,N_5252);
or U5459 (N_5459,N_5388,N_5341);
nand U5460 (N_5460,N_5281,N_5312);
and U5461 (N_5461,N_5229,N_5249);
nand U5462 (N_5462,N_5209,N_5343);
nor U5463 (N_5463,N_5291,N_5380);
nor U5464 (N_5464,N_5353,N_5293);
xnor U5465 (N_5465,N_5356,N_5283);
and U5466 (N_5466,N_5387,N_5303);
nor U5467 (N_5467,N_5390,N_5248);
nor U5468 (N_5468,N_5323,N_5328);
nand U5469 (N_5469,N_5299,N_5332);
nand U5470 (N_5470,N_5367,N_5260);
nand U5471 (N_5471,N_5244,N_5256);
and U5472 (N_5472,N_5271,N_5247);
nor U5473 (N_5473,N_5322,N_5268);
or U5474 (N_5474,N_5259,N_5236);
or U5475 (N_5475,N_5345,N_5285);
and U5476 (N_5476,N_5357,N_5362);
xor U5477 (N_5477,N_5277,N_5351);
or U5478 (N_5478,N_5394,N_5213);
and U5479 (N_5479,N_5368,N_5289);
or U5480 (N_5480,N_5212,N_5310);
and U5481 (N_5481,N_5360,N_5225);
xor U5482 (N_5482,N_5228,N_5231);
xor U5483 (N_5483,N_5324,N_5221);
nor U5484 (N_5484,N_5330,N_5246);
nand U5485 (N_5485,N_5296,N_5305);
xor U5486 (N_5486,N_5392,N_5301);
and U5487 (N_5487,N_5254,N_5297);
nor U5488 (N_5488,N_5265,N_5201);
xnor U5489 (N_5489,N_5306,N_5369);
and U5490 (N_5490,N_5321,N_5358);
nor U5491 (N_5491,N_5295,N_5315);
xor U5492 (N_5492,N_5304,N_5253);
xor U5493 (N_5493,N_5309,N_5391);
nand U5494 (N_5494,N_5284,N_5384);
nor U5495 (N_5495,N_5200,N_5398);
xor U5496 (N_5496,N_5202,N_5245);
nor U5497 (N_5497,N_5374,N_5234);
and U5498 (N_5498,N_5251,N_5208);
or U5499 (N_5499,N_5250,N_5364);
nand U5500 (N_5500,N_5201,N_5395);
or U5501 (N_5501,N_5298,N_5290);
and U5502 (N_5502,N_5289,N_5398);
xnor U5503 (N_5503,N_5292,N_5374);
xnor U5504 (N_5504,N_5317,N_5323);
xnor U5505 (N_5505,N_5388,N_5255);
and U5506 (N_5506,N_5280,N_5253);
and U5507 (N_5507,N_5210,N_5232);
and U5508 (N_5508,N_5232,N_5251);
nand U5509 (N_5509,N_5283,N_5303);
nand U5510 (N_5510,N_5212,N_5332);
nand U5511 (N_5511,N_5384,N_5274);
and U5512 (N_5512,N_5285,N_5235);
xnor U5513 (N_5513,N_5275,N_5287);
and U5514 (N_5514,N_5367,N_5256);
or U5515 (N_5515,N_5341,N_5333);
nor U5516 (N_5516,N_5331,N_5219);
or U5517 (N_5517,N_5245,N_5216);
or U5518 (N_5518,N_5263,N_5265);
or U5519 (N_5519,N_5260,N_5290);
or U5520 (N_5520,N_5385,N_5208);
xnor U5521 (N_5521,N_5275,N_5242);
xnor U5522 (N_5522,N_5261,N_5313);
nand U5523 (N_5523,N_5338,N_5224);
nand U5524 (N_5524,N_5272,N_5378);
and U5525 (N_5525,N_5207,N_5261);
and U5526 (N_5526,N_5357,N_5327);
xor U5527 (N_5527,N_5244,N_5294);
xnor U5528 (N_5528,N_5318,N_5225);
nor U5529 (N_5529,N_5211,N_5368);
and U5530 (N_5530,N_5399,N_5335);
nor U5531 (N_5531,N_5346,N_5393);
nand U5532 (N_5532,N_5396,N_5254);
xor U5533 (N_5533,N_5257,N_5310);
nor U5534 (N_5534,N_5315,N_5379);
or U5535 (N_5535,N_5388,N_5317);
xnor U5536 (N_5536,N_5258,N_5343);
nand U5537 (N_5537,N_5336,N_5294);
and U5538 (N_5538,N_5223,N_5241);
nor U5539 (N_5539,N_5333,N_5394);
xor U5540 (N_5540,N_5283,N_5325);
nand U5541 (N_5541,N_5342,N_5396);
and U5542 (N_5542,N_5385,N_5221);
nand U5543 (N_5543,N_5350,N_5268);
nor U5544 (N_5544,N_5359,N_5312);
or U5545 (N_5545,N_5330,N_5255);
nor U5546 (N_5546,N_5278,N_5337);
and U5547 (N_5547,N_5394,N_5250);
and U5548 (N_5548,N_5378,N_5329);
or U5549 (N_5549,N_5208,N_5396);
and U5550 (N_5550,N_5347,N_5267);
xor U5551 (N_5551,N_5211,N_5243);
or U5552 (N_5552,N_5213,N_5210);
nor U5553 (N_5553,N_5343,N_5295);
xor U5554 (N_5554,N_5281,N_5383);
nand U5555 (N_5555,N_5250,N_5332);
and U5556 (N_5556,N_5356,N_5260);
or U5557 (N_5557,N_5313,N_5391);
nand U5558 (N_5558,N_5397,N_5375);
and U5559 (N_5559,N_5337,N_5314);
nand U5560 (N_5560,N_5385,N_5384);
nor U5561 (N_5561,N_5399,N_5256);
nor U5562 (N_5562,N_5341,N_5395);
nor U5563 (N_5563,N_5230,N_5317);
nand U5564 (N_5564,N_5229,N_5375);
and U5565 (N_5565,N_5373,N_5240);
nor U5566 (N_5566,N_5327,N_5309);
nand U5567 (N_5567,N_5238,N_5363);
or U5568 (N_5568,N_5325,N_5279);
nor U5569 (N_5569,N_5239,N_5224);
xnor U5570 (N_5570,N_5283,N_5328);
or U5571 (N_5571,N_5348,N_5256);
nor U5572 (N_5572,N_5314,N_5299);
or U5573 (N_5573,N_5376,N_5271);
xnor U5574 (N_5574,N_5290,N_5253);
nand U5575 (N_5575,N_5332,N_5353);
nor U5576 (N_5576,N_5210,N_5330);
and U5577 (N_5577,N_5297,N_5377);
xnor U5578 (N_5578,N_5338,N_5237);
nand U5579 (N_5579,N_5289,N_5230);
or U5580 (N_5580,N_5328,N_5343);
nand U5581 (N_5581,N_5295,N_5259);
or U5582 (N_5582,N_5275,N_5229);
or U5583 (N_5583,N_5396,N_5322);
nor U5584 (N_5584,N_5329,N_5337);
nor U5585 (N_5585,N_5293,N_5369);
or U5586 (N_5586,N_5284,N_5364);
xor U5587 (N_5587,N_5331,N_5217);
nor U5588 (N_5588,N_5372,N_5373);
or U5589 (N_5589,N_5265,N_5398);
nand U5590 (N_5590,N_5383,N_5201);
xnor U5591 (N_5591,N_5244,N_5327);
xnor U5592 (N_5592,N_5299,N_5334);
nor U5593 (N_5593,N_5261,N_5237);
and U5594 (N_5594,N_5340,N_5268);
nor U5595 (N_5595,N_5279,N_5373);
or U5596 (N_5596,N_5248,N_5219);
nand U5597 (N_5597,N_5351,N_5356);
or U5598 (N_5598,N_5364,N_5203);
xor U5599 (N_5599,N_5223,N_5341);
and U5600 (N_5600,N_5487,N_5452);
and U5601 (N_5601,N_5471,N_5538);
nand U5602 (N_5602,N_5596,N_5533);
or U5603 (N_5603,N_5551,N_5453);
and U5604 (N_5604,N_5427,N_5440);
or U5605 (N_5605,N_5567,N_5485);
and U5606 (N_5606,N_5597,N_5511);
xor U5607 (N_5607,N_5474,N_5508);
and U5608 (N_5608,N_5585,N_5575);
xnor U5609 (N_5609,N_5531,N_5528);
xor U5610 (N_5610,N_5592,N_5483);
or U5611 (N_5611,N_5515,N_5490);
and U5612 (N_5612,N_5498,N_5543);
xor U5613 (N_5613,N_5430,N_5507);
xnor U5614 (N_5614,N_5496,N_5488);
nor U5615 (N_5615,N_5569,N_5524);
nor U5616 (N_5616,N_5595,N_5449);
xor U5617 (N_5617,N_5432,N_5428);
nand U5618 (N_5618,N_5505,N_5421);
and U5619 (N_5619,N_5426,N_5541);
nor U5620 (N_5620,N_5502,N_5521);
nor U5621 (N_5621,N_5557,N_5436);
nand U5622 (N_5622,N_5469,N_5423);
nand U5623 (N_5623,N_5580,N_5562);
nand U5624 (N_5624,N_5573,N_5413);
nand U5625 (N_5625,N_5410,N_5500);
and U5626 (N_5626,N_5402,N_5493);
nand U5627 (N_5627,N_5547,N_5462);
xnor U5628 (N_5628,N_5518,N_5486);
nor U5629 (N_5629,N_5470,N_5442);
nand U5630 (N_5630,N_5571,N_5527);
nor U5631 (N_5631,N_5459,N_5454);
nor U5632 (N_5632,N_5472,N_5499);
and U5633 (N_5633,N_5534,N_5460);
xnor U5634 (N_5634,N_5549,N_5420);
and U5635 (N_5635,N_5482,N_5444);
xor U5636 (N_5636,N_5552,N_5503);
nand U5637 (N_5637,N_5583,N_5455);
nor U5638 (N_5638,N_5556,N_5407);
and U5639 (N_5639,N_5591,N_5588);
or U5640 (N_5640,N_5526,N_5548);
nand U5641 (N_5641,N_5418,N_5555);
nor U5642 (N_5642,N_5559,N_5582);
nand U5643 (N_5643,N_5450,N_5491);
xnor U5644 (N_5644,N_5476,N_5540);
xnor U5645 (N_5645,N_5512,N_5593);
nor U5646 (N_5646,N_5401,N_5536);
and U5647 (N_5647,N_5404,N_5479);
nor U5648 (N_5648,N_5566,N_5544);
and U5649 (N_5649,N_5523,N_5473);
and U5650 (N_5650,N_5519,N_5599);
nand U5651 (N_5651,N_5461,N_5587);
nor U5652 (N_5652,N_5445,N_5522);
or U5653 (N_5653,N_5513,N_5537);
xor U5654 (N_5654,N_5561,N_5400);
and U5655 (N_5655,N_5589,N_5532);
xnor U5656 (N_5656,N_5466,N_5530);
nor U5657 (N_5657,N_5412,N_5446);
or U5658 (N_5658,N_5458,N_5542);
nor U5659 (N_5659,N_5563,N_5572);
nand U5660 (N_5660,N_5405,N_5424);
xnor U5661 (N_5661,N_5516,N_5489);
nand U5662 (N_5662,N_5517,N_5484);
and U5663 (N_5663,N_5558,N_5584);
and U5664 (N_5664,N_5550,N_5409);
xor U5665 (N_5665,N_5594,N_5497);
or U5666 (N_5666,N_5429,N_5431);
or U5667 (N_5667,N_5577,N_5457);
or U5668 (N_5668,N_5448,N_5415);
nand U5669 (N_5669,N_5411,N_5579);
and U5670 (N_5670,N_5414,N_5475);
nand U5671 (N_5671,N_5564,N_5465);
nor U5672 (N_5672,N_5529,N_5539);
nand U5673 (N_5673,N_5416,N_5438);
and U5674 (N_5674,N_5560,N_5525);
and U5675 (N_5675,N_5422,N_5477);
nand U5676 (N_5676,N_5494,N_5514);
and U5677 (N_5677,N_5510,N_5439);
nand U5678 (N_5678,N_5492,N_5403);
nor U5679 (N_5679,N_5481,N_5435);
nand U5680 (N_5680,N_5419,N_5447);
xor U5681 (N_5681,N_5408,N_5554);
xor U5682 (N_5682,N_5535,N_5520);
nand U5683 (N_5683,N_5598,N_5576);
and U5684 (N_5684,N_5586,N_5478);
nor U5685 (N_5685,N_5506,N_5495);
and U5686 (N_5686,N_5553,N_5467);
and U5687 (N_5687,N_5425,N_5574);
nand U5688 (N_5688,N_5504,N_5568);
nand U5689 (N_5689,N_5406,N_5437);
and U5690 (N_5690,N_5451,N_5578);
xor U5691 (N_5691,N_5463,N_5546);
xor U5692 (N_5692,N_5501,N_5417);
or U5693 (N_5693,N_5443,N_5590);
and U5694 (N_5694,N_5581,N_5456);
and U5695 (N_5695,N_5509,N_5480);
and U5696 (N_5696,N_5468,N_5570);
nand U5697 (N_5697,N_5433,N_5434);
nand U5698 (N_5698,N_5464,N_5565);
or U5699 (N_5699,N_5441,N_5545);
and U5700 (N_5700,N_5434,N_5563);
nor U5701 (N_5701,N_5559,N_5466);
or U5702 (N_5702,N_5407,N_5589);
and U5703 (N_5703,N_5527,N_5542);
nand U5704 (N_5704,N_5584,N_5549);
nand U5705 (N_5705,N_5422,N_5441);
xnor U5706 (N_5706,N_5496,N_5526);
or U5707 (N_5707,N_5476,N_5575);
xor U5708 (N_5708,N_5431,N_5554);
nor U5709 (N_5709,N_5515,N_5414);
and U5710 (N_5710,N_5529,N_5523);
and U5711 (N_5711,N_5484,N_5465);
nor U5712 (N_5712,N_5400,N_5458);
xnor U5713 (N_5713,N_5440,N_5510);
xor U5714 (N_5714,N_5414,N_5498);
nand U5715 (N_5715,N_5473,N_5489);
xor U5716 (N_5716,N_5422,N_5471);
nand U5717 (N_5717,N_5425,N_5597);
or U5718 (N_5718,N_5481,N_5508);
or U5719 (N_5719,N_5512,N_5582);
or U5720 (N_5720,N_5470,N_5467);
xor U5721 (N_5721,N_5544,N_5578);
or U5722 (N_5722,N_5565,N_5562);
and U5723 (N_5723,N_5449,N_5521);
xnor U5724 (N_5724,N_5504,N_5485);
and U5725 (N_5725,N_5404,N_5581);
and U5726 (N_5726,N_5591,N_5491);
nor U5727 (N_5727,N_5404,N_5510);
and U5728 (N_5728,N_5460,N_5470);
xor U5729 (N_5729,N_5586,N_5402);
nor U5730 (N_5730,N_5480,N_5497);
nor U5731 (N_5731,N_5579,N_5444);
nor U5732 (N_5732,N_5442,N_5569);
and U5733 (N_5733,N_5582,N_5444);
and U5734 (N_5734,N_5498,N_5442);
and U5735 (N_5735,N_5494,N_5418);
xor U5736 (N_5736,N_5459,N_5529);
nor U5737 (N_5737,N_5433,N_5474);
nor U5738 (N_5738,N_5590,N_5448);
and U5739 (N_5739,N_5417,N_5433);
nor U5740 (N_5740,N_5546,N_5508);
or U5741 (N_5741,N_5412,N_5473);
nand U5742 (N_5742,N_5570,N_5578);
nor U5743 (N_5743,N_5503,N_5517);
or U5744 (N_5744,N_5404,N_5587);
and U5745 (N_5745,N_5575,N_5423);
xor U5746 (N_5746,N_5478,N_5438);
xor U5747 (N_5747,N_5420,N_5401);
xor U5748 (N_5748,N_5582,N_5581);
or U5749 (N_5749,N_5436,N_5563);
nand U5750 (N_5750,N_5577,N_5585);
or U5751 (N_5751,N_5471,N_5569);
nor U5752 (N_5752,N_5448,N_5551);
and U5753 (N_5753,N_5521,N_5443);
or U5754 (N_5754,N_5428,N_5418);
or U5755 (N_5755,N_5548,N_5459);
nand U5756 (N_5756,N_5530,N_5588);
nor U5757 (N_5757,N_5590,N_5575);
or U5758 (N_5758,N_5438,N_5556);
and U5759 (N_5759,N_5543,N_5546);
and U5760 (N_5760,N_5541,N_5498);
xor U5761 (N_5761,N_5457,N_5595);
nand U5762 (N_5762,N_5424,N_5460);
nand U5763 (N_5763,N_5510,N_5575);
and U5764 (N_5764,N_5433,N_5554);
xnor U5765 (N_5765,N_5521,N_5596);
or U5766 (N_5766,N_5491,N_5549);
or U5767 (N_5767,N_5574,N_5515);
nand U5768 (N_5768,N_5569,N_5505);
and U5769 (N_5769,N_5560,N_5588);
or U5770 (N_5770,N_5519,N_5533);
nand U5771 (N_5771,N_5482,N_5537);
xor U5772 (N_5772,N_5527,N_5578);
or U5773 (N_5773,N_5447,N_5450);
or U5774 (N_5774,N_5547,N_5467);
and U5775 (N_5775,N_5532,N_5586);
nor U5776 (N_5776,N_5582,N_5579);
nor U5777 (N_5777,N_5425,N_5450);
and U5778 (N_5778,N_5537,N_5523);
xor U5779 (N_5779,N_5527,N_5458);
nand U5780 (N_5780,N_5501,N_5592);
xnor U5781 (N_5781,N_5429,N_5579);
xnor U5782 (N_5782,N_5512,N_5452);
xnor U5783 (N_5783,N_5433,N_5524);
nand U5784 (N_5784,N_5444,N_5471);
nand U5785 (N_5785,N_5440,N_5559);
nor U5786 (N_5786,N_5479,N_5527);
or U5787 (N_5787,N_5431,N_5561);
nor U5788 (N_5788,N_5412,N_5507);
or U5789 (N_5789,N_5487,N_5490);
xnor U5790 (N_5790,N_5532,N_5598);
or U5791 (N_5791,N_5520,N_5541);
xnor U5792 (N_5792,N_5556,N_5405);
and U5793 (N_5793,N_5585,N_5586);
or U5794 (N_5794,N_5573,N_5457);
or U5795 (N_5795,N_5585,N_5456);
and U5796 (N_5796,N_5451,N_5530);
nand U5797 (N_5797,N_5484,N_5499);
nor U5798 (N_5798,N_5519,N_5583);
or U5799 (N_5799,N_5592,N_5424);
or U5800 (N_5800,N_5755,N_5600);
or U5801 (N_5801,N_5640,N_5642);
and U5802 (N_5802,N_5713,N_5638);
or U5803 (N_5803,N_5610,N_5679);
nand U5804 (N_5804,N_5792,N_5765);
or U5805 (N_5805,N_5677,N_5795);
nand U5806 (N_5806,N_5668,N_5714);
or U5807 (N_5807,N_5673,N_5750);
xnor U5808 (N_5808,N_5774,N_5617);
and U5809 (N_5809,N_5698,N_5696);
xor U5810 (N_5810,N_5629,N_5747);
or U5811 (N_5811,N_5781,N_5704);
nor U5812 (N_5812,N_5633,N_5631);
and U5813 (N_5813,N_5691,N_5794);
nand U5814 (N_5814,N_5606,N_5743);
xnor U5815 (N_5815,N_5670,N_5685);
nor U5816 (N_5816,N_5654,N_5793);
nor U5817 (N_5817,N_5707,N_5660);
or U5818 (N_5818,N_5632,N_5614);
nand U5819 (N_5819,N_5760,N_5784);
and U5820 (N_5820,N_5608,N_5788);
xor U5821 (N_5821,N_5653,N_5643);
or U5822 (N_5822,N_5720,N_5761);
nand U5823 (N_5823,N_5607,N_5627);
or U5824 (N_5824,N_5729,N_5712);
xnor U5825 (N_5825,N_5796,N_5611);
nand U5826 (N_5826,N_5605,N_5733);
or U5827 (N_5827,N_5757,N_5635);
nor U5828 (N_5828,N_5694,N_5728);
xnor U5829 (N_5829,N_5613,N_5647);
nor U5830 (N_5830,N_5651,N_5766);
nand U5831 (N_5831,N_5775,N_5697);
and U5832 (N_5832,N_5648,N_5620);
nand U5833 (N_5833,N_5721,N_5604);
xor U5834 (N_5834,N_5759,N_5674);
xor U5835 (N_5835,N_5767,N_5780);
nand U5836 (N_5836,N_5734,N_5739);
nand U5837 (N_5837,N_5783,N_5754);
nand U5838 (N_5838,N_5601,N_5602);
nor U5839 (N_5839,N_5661,N_5778);
or U5840 (N_5840,N_5786,N_5634);
nand U5841 (N_5841,N_5692,N_5715);
nor U5842 (N_5842,N_5756,N_5687);
xor U5843 (N_5843,N_5763,N_5693);
or U5844 (N_5844,N_5652,N_5650);
or U5845 (N_5845,N_5625,N_5737);
nor U5846 (N_5846,N_5742,N_5695);
and U5847 (N_5847,N_5748,N_5686);
nor U5848 (N_5848,N_5680,N_5669);
or U5849 (N_5849,N_5645,N_5641);
and U5850 (N_5850,N_5787,N_5624);
or U5851 (N_5851,N_5785,N_5615);
nand U5852 (N_5852,N_5740,N_5744);
and U5853 (N_5853,N_5749,N_5789);
and U5854 (N_5854,N_5738,N_5639);
nand U5855 (N_5855,N_5776,N_5609);
nand U5856 (N_5856,N_5730,N_5665);
nor U5857 (N_5857,N_5798,N_5736);
xor U5858 (N_5858,N_5758,N_5701);
and U5859 (N_5859,N_5671,N_5727);
nand U5860 (N_5860,N_5618,N_5675);
nand U5861 (N_5861,N_5710,N_5658);
or U5862 (N_5862,N_5626,N_5644);
or U5863 (N_5863,N_5630,N_5772);
and U5864 (N_5864,N_5782,N_5731);
xnor U5865 (N_5865,N_5699,N_5623);
and U5866 (N_5866,N_5619,N_5657);
or U5867 (N_5867,N_5797,N_5649);
xor U5868 (N_5868,N_5735,N_5666);
nor U5869 (N_5869,N_5708,N_5636);
or U5870 (N_5870,N_5700,N_5779);
nor U5871 (N_5871,N_5732,N_5664);
nand U5872 (N_5872,N_5777,N_5616);
xnor U5873 (N_5873,N_5722,N_5790);
nor U5874 (N_5874,N_5655,N_5706);
or U5875 (N_5875,N_5746,N_5667);
xnor U5876 (N_5876,N_5702,N_5689);
nor U5877 (N_5877,N_5711,N_5684);
and U5878 (N_5878,N_5764,N_5716);
or U5879 (N_5879,N_5769,N_5672);
nand U5880 (N_5880,N_5718,N_5603);
and U5881 (N_5881,N_5621,N_5725);
or U5882 (N_5882,N_5724,N_5709);
nand U5883 (N_5883,N_5703,N_5683);
xnor U5884 (N_5884,N_5646,N_5705);
xor U5885 (N_5885,N_5799,N_5771);
xnor U5886 (N_5886,N_5762,N_5768);
nor U5887 (N_5887,N_5637,N_5622);
or U5888 (N_5888,N_5659,N_5753);
and U5889 (N_5889,N_5745,N_5773);
or U5890 (N_5890,N_5752,N_5628);
and U5891 (N_5891,N_5682,N_5676);
xor U5892 (N_5892,N_5726,N_5741);
nor U5893 (N_5893,N_5662,N_5690);
nor U5894 (N_5894,N_5770,N_5688);
xor U5895 (N_5895,N_5681,N_5791);
nand U5896 (N_5896,N_5723,N_5751);
nor U5897 (N_5897,N_5678,N_5717);
nand U5898 (N_5898,N_5663,N_5656);
xor U5899 (N_5899,N_5612,N_5719);
or U5900 (N_5900,N_5653,N_5714);
xnor U5901 (N_5901,N_5736,N_5754);
and U5902 (N_5902,N_5646,N_5676);
nand U5903 (N_5903,N_5714,N_5739);
nand U5904 (N_5904,N_5735,N_5782);
nor U5905 (N_5905,N_5743,N_5663);
nor U5906 (N_5906,N_5662,N_5735);
nand U5907 (N_5907,N_5798,N_5745);
or U5908 (N_5908,N_5694,N_5778);
or U5909 (N_5909,N_5667,N_5617);
nand U5910 (N_5910,N_5753,N_5660);
nand U5911 (N_5911,N_5758,N_5746);
or U5912 (N_5912,N_5777,N_5627);
nor U5913 (N_5913,N_5763,N_5701);
nor U5914 (N_5914,N_5778,N_5605);
and U5915 (N_5915,N_5674,N_5688);
and U5916 (N_5916,N_5656,N_5792);
nor U5917 (N_5917,N_5762,N_5654);
and U5918 (N_5918,N_5692,N_5734);
xnor U5919 (N_5919,N_5678,N_5723);
or U5920 (N_5920,N_5628,N_5713);
and U5921 (N_5921,N_5773,N_5613);
nor U5922 (N_5922,N_5692,N_5642);
and U5923 (N_5923,N_5706,N_5747);
or U5924 (N_5924,N_5796,N_5772);
nor U5925 (N_5925,N_5609,N_5769);
nand U5926 (N_5926,N_5684,N_5778);
or U5927 (N_5927,N_5602,N_5627);
nand U5928 (N_5928,N_5660,N_5667);
nor U5929 (N_5929,N_5708,N_5724);
nor U5930 (N_5930,N_5630,N_5649);
or U5931 (N_5931,N_5630,N_5631);
xor U5932 (N_5932,N_5724,N_5702);
nand U5933 (N_5933,N_5632,N_5755);
or U5934 (N_5934,N_5762,N_5740);
or U5935 (N_5935,N_5621,N_5627);
nand U5936 (N_5936,N_5708,N_5607);
or U5937 (N_5937,N_5701,N_5605);
xor U5938 (N_5938,N_5695,N_5668);
and U5939 (N_5939,N_5773,N_5659);
nand U5940 (N_5940,N_5663,N_5617);
xor U5941 (N_5941,N_5665,N_5739);
and U5942 (N_5942,N_5661,N_5712);
nor U5943 (N_5943,N_5758,N_5600);
nor U5944 (N_5944,N_5677,N_5603);
nor U5945 (N_5945,N_5699,N_5622);
or U5946 (N_5946,N_5736,N_5766);
and U5947 (N_5947,N_5731,N_5719);
or U5948 (N_5948,N_5721,N_5642);
or U5949 (N_5949,N_5683,N_5644);
or U5950 (N_5950,N_5766,N_5632);
and U5951 (N_5951,N_5683,N_5695);
nor U5952 (N_5952,N_5655,N_5788);
and U5953 (N_5953,N_5654,N_5789);
nor U5954 (N_5954,N_5635,N_5625);
or U5955 (N_5955,N_5686,N_5765);
and U5956 (N_5956,N_5796,N_5613);
or U5957 (N_5957,N_5664,N_5628);
nand U5958 (N_5958,N_5758,N_5627);
and U5959 (N_5959,N_5729,N_5670);
xor U5960 (N_5960,N_5723,N_5702);
and U5961 (N_5961,N_5646,N_5615);
nand U5962 (N_5962,N_5606,N_5738);
or U5963 (N_5963,N_5753,N_5766);
or U5964 (N_5964,N_5637,N_5721);
nor U5965 (N_5965,N_5698,N_5618);
nor U5966 (N_5966,N_5689,N_5672);
nand U5967 (N_5967,N_5619,N_5678);
and U5968 (N_5968,N_5600,N_5651);
nand U5969 (N_5969,N_5797,N_5720);
or U5970 (N_5970,N_5634,N_5699);
nor U5971 (N_5971,N_5602,N_5669);
nor U5972 (N_5972,N_5676,N_5641);
nand U5973 (N_5973,N_5648,N_5766);
nand U5974 (N_5974,N_5681,N_5672);
and U5975 (N_5975,N_5606,N_5796);
nand U5976 (N_5976,N_5780,N_5612);
nand U5977 (N_5977,N_5671,N_5711);
xnor U5978 (N_5978,N_5618,N_5646);
nand U5979 (N_5979,N_5732,N_5752);
xnor U5980 (N_5980,N_5626,N_5761);
or U5981 (N_5981,N_5783,N_5607);
nand U5982 (N_5982,N_5681,N_5661);
and U5983 (N_5983,N_5780,N_5779);
and U5984 (N_5984,N_5628,N_5762);
nor U5985 (N_5985,N_5673,N_5725);
nor U5986 (N_5986,N_5792,N_5732);
and U5987 (N_5987,N_5659,N_5699);
xnor U5988 (N_5988,N_5662,N_5650);
or U5989 (N_5989,N_5631,N_5692);
xor U5990 (N_5990,N_5680,N_5657);
nor U5991 (N_5991,N_5777,N_5608);
or U5992 (N_5992,N_5616,N_5692);
xor U5993 (N_5993,N_5623,N_5701);
nor U5994 (N_5994,N_5623,N_5674);
xor U5995 (N_5995,N_5750,N_5755);
and U5996 (N_5996,N_5713,N_5615);
xnor U5997 (N_5997,N_5708,N_5694);
nand U5998 (N_5998,N_5758,N_5742);
or U5999 (N_5999,N_5717,N_5738);
and U6000 (N_6000,N_5942,N_5820);
nor U6001 (N_6001,N_5803,N_5932);
or U6002 (N_6002,N_5986,N_5938);
or U6003 (N_6003,N_5821,N_5949);
and U6004 (N_6004,N_5880,N_5846);
or U6005 (N_6005,N_5983,N_5886);
and U6006 (N_6006,N_5895,N_5967);
nor U6007 (N_6007,N_5940,N_5947);
xnor U6008 (N_6008,N_5988,N_5975);
xor U6009 (N_6009,N_5999,N_5931);
nor U6010 (N_6010,N_5995,N_5875);
or U6011 (N_6011,N_5815,N_5876);
nand U6012 (N_6012,N_5869,N_5836);
nand U6013 (N_6013,N_5851,N_5955);
nor U6014 (N_6014,N_5837,N_5963);
nand U6015 (N_6015,N_5933,N_5897);
xnor U6016 (N_6016,N_5968,N_5984);
nand U6017 (N_6017,N_5900,N_5874);
nand U6018 (N_6018,N_5921,N_5887);
and U6019 (N_6019,N_5996,N_5832);
xnor U6020 (N_6020,N_5926,N_5970);
and U6021 (N_6021,N_5861,N_5878);
and U6022 (N_6022,N_5866,N_5884);
nor U6023 (N_6023,N_5953,N_5948);
xor U6024 (N_6024,N_5960,N_5989);
nor U6025 (N_6025,N_5936,N_5980);
and U6026 (N_6026,N_5828,N_5864);
or U6027 (N_6027,N_5808,N_5981);
xnor U6028 (N_6028,N_5863,N_5993);
xor U6029 (N_6029,N_5838,N_5951);
or U6030 (N_6030,N_5823,N_5817);
or U6031 (N_6031,N_5859,N_5892);
and U6032 (N_6032,N_5841,N_5829);
nand U6033 (N_6033,N_5872,N_5814);
and U6034 (N_6034,N_5908,N_5957);
or U6035 (N_6035,N_5972,N_5910);
nor U6036 (N_6036,N_5925,N_5944);
nor U6037 (N_6037,N_5894,N_5802);
nand U6038 (N_6038,N_5896,N_5881);
nand U6039 (N_6039,N_5825,N_5819);
and U6040 (N_6040,N_5840,N_5907);
or U6041 (N_6041,N_5835,N_5915);
or U6042 (N_6042,N_5992,N_5853);
xor U6043 (N_6043,N_5974,N_5826);
nor U6044 (N_6044,N_5816,N_5801);
nand U6045 (N_6045,N_5843,N_5800);
nand U6046 (N_6046,N_5950,N_5918);
nand U6047 (N_6047,N_5935,N_5810);
or U6048 (N_6048,N_5994,N_5804);
nor U6049 (N_6049,N_5877,N_5952);
xnor U6050 (N_6050,N_5901,N_5807);
nand U6051 (N_6051,N_5844,N_5871);
xnor U6052 (N_6052,N_5973,N_5987);
and U6053 (N_6053,N_5873,N_5812);
and U6054 (N_6054,N_5862,N_5834);
or U6055 (N_6055,N_5852,N_5839);
and U6056 (N_6056,N_5905,N_5958);
nor U6057 (N_6057,N_5976,N_5930);
nor U6058 (N_6058,N_5911,N_5856);
and U6059 (N_6059,N_5906,N_5961);
nand U6060 (N_6060,N_5858,N_5854);
nand U6061 (N_6061,N_5865,N_5912);
nand U6062 (N_6062,N_5870,N_5927);
or U6063 (N_6063,N_5822,N_5937);
xor U6064 (N_6064,N_5917,N_5833);
nor U6065 (N_6065,N_5850,N_5998);
nand U6066 (N_6066,N_5965,N_5885);
nand U6067 (N_6067,N_5818,N_5997);
or U6068 (N_6068,N_5923,N_5929);
xor U6069 (N_6069,N_5831,N_5978);
nand U6070 (N_6070,N_5943,N_5824);
xnor U6071 (N_6071,N_5919,N_5945);
nand U6072 (N_6072,N_5946,N_5888);
nand U6073 (N_6073,N_5860,N_5916);
nor U6074 (N_6074,N_5879,N_5849);
nand U6075 (N_6075,N_5966,N_5848);
nand U6076 (N_6076,N_5845,N_5893);
xor U6077 (N_6077,N_5939,N_5954);
nor U6078 (N_6078,N_5928,N_5934);
nand U6079 (N_6079,N_5982,N_5842);
and U6080 (N_6080,N_5979,N_5898);
xor U6081 (N_6081,N_5867,N_5902);
xor U6082 (N_6082,N_5985,N_5969);
or U6083 (N_6083,N_5890,N_5920);
or U6084 (N_6084,N_5991,N_5956);
nor U6085 (N_6085,N_5847,N_5809);
or U6086 (N_6086,N_5914,N_5990);
or U6087 (N_6087,N_5962,N_5806);
or U6088 (N_6088,N_5813,N_5805);
nand U6089 (N_6089,N_5855,N_5959);
or U6090 (N_6090,N_5941,N_5883);
xor U6091 (N_6091,N_5811,N_5977);
nor U6092 (N_6092,N_5868,N_5882);
nor U6093 (N_6093,N_5899,N_5889);
or U6094 (N_6094,N_5904,N_5857);
or U6095 (N_6095,N_5913,N_5909);
nor U6096 (N_6096,N_5964,N_5891);
and U6097 (N_6097,N_5971,N_5924);
nor U6098 (N_6098,N_5830,N_5903);
and U6099 (N_6099,N_5922,N_5827);
xor U6100 (N_6100,N_5817,N_5835);
and U6101 (N_6101,N_5926,N_5875);
and U6102 (N_6102,N_5842,N_5954);
and U6103 (N_6103,N_5874,N_5821);
nor U6104 (N_6104,N_5980,N_5821);
or U6105 (N_6105,N_5990,N_5801);
and U6106 (N_6106,N_5802,N_5993);
xor U6107 (N_6107,N_5982,N_5931);
nand U6108 (N_6108,N_5828,N_5942);
or U6109 (N_6109,N_5919,N_5938);
nand U6110 (N_6110,N_5841,N_5946);
xnor U6111 (N_6111,N_5819,N_5896);
xor U6112 (N_6112,N_5930,N_5895);
nor U6113 (N_6113,N_5883,N_5925);
nor U6114 (N_6114,N_5821,N_5897);
nor U6115 (N_6115,N_5803,N_5824);
or U6116 (N_6116,N_5883,N_5830);
or U6117 (N_6117,N_5952,N_5806);
and U6118 (N_6118,N_5848,N_5932);
nand U6119 (N_6119,N_5893,N_5849);
nor U6120 (N_6120,N_5856,N_5953);
xnor U6121 (N_6121,N_5937,N_5854);
nand U6122 (N_6122,N_5939,N_5838);
nor U6123 (N_6123,N_5915,N_5853);
or U6124 (N_6124,N_5866,N_5989);
nor U6125 (N_6125,N_5838,N_5829);
or U6126 (N_6126,N_5836,N_5942);
nor U6127 (N_6127,N_5860,N_5819);
nand U6128 (N_6128,N_5999,N_5900);
or U6129 (N_6129,N_5994,N_5894);
and U6130 (N_6130,N_5934,N_5848);
nand U6131 (N_6131,N_5972,N_5922);
nand U6132 (N_6132,N_5910,N_5807);
or U6133 (N_6133,N_5996,N_5995);
and U6134 (N_6134,N_5967,N_5844);
nor U6135 (N_6135,N_5955,N_5803);
or U6136 (N_6136,N_5898,N_5875);
nor U6137 (N_6137,N_5928,N_5916);
or U6138 (N_6138,N_5921,N_5915);
and U6139 (N_6139,N_5810,N_5909);
xnor U6140 (N_6140,N_5968,N_5878);
xnor U6141 (N_6141,N_5892,N_5815);
and U6142 (N_6142,N_5801,N_5888);
and U6143 (N_6143,N_5917,N_5866);
nor U6144 (N_6144,N_5982,N_5950);
nor U6145 (N_6145,N_5873,N_5955);
and U6146 (N_6146,N_5965,N_5884);
nand U6147 (N_6147,N_5912,N_5848);
nand U6148 (N_6148,N_5821,N_5855);
nor U6149 (N_6149,N_5817,N_5916);
nor U6150 (N_6150,N_5902,N_5811);
and U6151 (N_6151,N_5863,N_5828);
or U6152 (N_6152,N_5868,N_5806);
nor U6153 (N_6153,N_5947,N_5886);
nand U6154 (N_6154,N_5919,N_5904);
and U6155 (N_6155,N_5853,N_5938);
nand U6156 (N_6156,N_5936,N_5839);
and U6157 (N_6157,N_5985,N_5871);
or U6158 (N_6158,N_5891,N_5816);
or U6159 (N_6159,N_5808,N_5885);
nor U6160 (N_6160,N_5925,N_5978);
nor U6161 (N_6161,N_5883,N_5886);
nand U6162 (N_6162,N_5924,N_5811);
and U6163 (N_6163,N_5904,N_5863);
and U6164 (N_6164,N_5897,N_5946);
xnor U6165 (N_6165,N_5892,N_5853);
xnor U6166 (N_6166,N_5983,N_5849);
nand U6167 (N_6167,N_5831,N_5847);
or U6168 (N_6168,N_5838,N_5869);
nand U6169 (N_6169,N_5926,N_5985);
xor U6170 (N_6170,N_5898,N_5944);
and U6171 (N_6171,N_5874,N_5979);
nand U6172 (N_6172,N_5880,N_5936);
nand U6173 (N_6173,N_5959,N_5988);
xor U6174 (N_6174,N_5818,N_5956);
nand U6175 (N_6175,N_5850,N_5936);
nor U6176 (N_6176,N_5807,N_5977);
or U6177 (N_6177,N_5871,N_5957);
nor U6178 (N_6178,N_5953,N_5947);
and U6179 (N_6179,N_5969,N_5925);
nor U6180 (N_6180,N_5899,N_5961);
nor U6181 (N_6181,N_5866,N_5977);
nand U6182 (N_6182,N_5956,N_5977);
nand U6183 (N_6183,N_5897,N_5998);
nand U6184 (N_6184,N_5884,N_5995);
nand U6185 (N_6185,N_5965,N_5807);
xor U6186 (N_6186,N_5852,N_5891);
nand U6187 (N_6187,N_5920,N_5967);
or U6188 (N_6188,N_5805,N_5875);
nand U6189 (N_6189,N_5816,N_5998);
or U6190 (N_6190,N_5859,N_5959);
xor U6191 (N_6191,N_5978,N_5999);
nor U6192 (N_6192,N_5891,N_5899);
and U6193 (N_6193,N_5923,N_5965);
and U6194 (N_6194,N_5822,N_5992);
xnor U6195 (N_6195,N_5924,N_5830);
xnor U6196 (N_6196,N_5804,N_5902);
nor U6197 (N_6197,N_5981,N_5911);
or U6198 (N_6198,N_5958,N_5972);
and U6199 (N_6199,N_5890,N_5914);
nor U6200 (N_6200,N_6083,N_6033);
nand U6201 (N_6201,N_6099,N_6055);
xnor U6202 (N_6202,N_6092,N_6176);
nor U6203 (N_6203,N_6103,N_6028);
and U6204 (N_6204,N_6021,N_6008);
nand U6205 (N_6205,N_6041,N_6047);
and U6206 (N_6206,N_6091,N_6090);
nor U6207 (N_6207,N_6130,N_6076);
and U6208 (N_6208,N_6114,N_6012);
or U6209 (N_6209,N_6072,N_6175);
or U6210 (N_6210,N_6115,N_6146);
nand U6211 (N_6211,N_6081,N_6117);
and U6212 (N_6212,N_6185,N_6144);
xnor U6213 (N_6213,N_6181,N_6166);
xnor U6214 (N_6214,N_6156,N_6109);
nand U6215 (N_6215,N_6174,N_6095);
nor U6216 (N_6216,N_6140,N_6048);
or U6217 (N_6217,N_6105,N_6085);
or U6218 (N_6218,N_6006,N_6122);
nand U6219 (N_6219,N_6043,N_6116);
and U6220 (N_6220,N_6193,N_6158);
and U6221 (N_6221,N_6194,N_6100);
nor U6222 (N_6222,N_6017,N_6135);
nor U6223 (N_6223,N_6057,N_6183);
or U6224 (N_6224,N_6142,N_6179);
and U6225 (N_6225,N_6066,N_6037);
nand U6226 (N_6226,N_6040,N_6123);
or U6227 (N_6227,N_6065,N_6190);
nor U6228 (N_6228,N_6010,N_6042);
and U6229 (N_6229,N_6056,N_6199);
xnor U6230 (N_6230,N_6112,N_6126);
nor U6231 (N_6231,N_6016,N_6075);
nor U6232 (N_6232,N_6071,N_6108);
nor U6233 (N_6233,N_6074,N_6138);
and U6234 (N_6234,N_6080,N_6162);
and U6235 (N_6235,N_6184,N_6155);
and U6236 (N_6236,N_6059,N_6125);
nand U6237 (N_6237,N_6002,N_6068);
nor U6238 (N_6238,N_6195,N_6198);
and U6239 (N_6239,N_6004,N_6061);
or U6240 (N_6240,N_6035,N_6089);
nand U6241 (N_6241,N_6029,N_6069);
or U6242 (N_6242,N_6157,N_6128);
nand U6243 (N_6243,N_6054,N_6171);
nor U6244 (N_6244,N_6143,N_6024);
nor U6245 (N_6245,N_6079,N_6014);
nand U6246 (N_6246,N_6177,N_6187);
nand U6247 (N_6247,N_6088,N_6032);
nor U6248 (N_6248,N_6005,N_6182);
or U6249 (N_6249,N_6051,N_6159);
nor U6250 (N_6250,N_6107,N_6023);
or U6251 (N_6251,N_6036,N_6082);
nand U6252 (N_6252,N_6149,N_6173);
xnor U6253 (N_6253,N_6087,N_6077);
xnor U6254 (N_6254,N_6009,N_6104);
nor U6255 (N_6255,N_6191,N_6015);
or U6256 (N_6256,N_6011,N_6169);
nand U6257 (N_6257,N_6164,N_6063);
nor U6258 (N_6258,N_6038,N_6102);
xnor U6259 (N_6259,N_6013,N_6027);
nor U6260 (N_6260,N_6148,N_6058);
nand U6261 (N_6261,N_6073,N_6129);
or U6262 (N_6262,N_6007,N_6049);
and U6263 (N_6263,N_6031,N_6165);
and U6264 (N_6264,N_6101,N_6044);
nand U6265 (N_6265,N_6163,N_6139);
nor U6266 (N_6266,N_6180,N_6018);
nand U6267 (N_6267,N_6094,N_6168);
xnor U6268 (N_6268,N_6111,N_6045);
xor U6269 (N_6269,N_6192,N_6064);
nor U6270 (N_6270,N_6060,N_6046);
and U6271 (N_6271,N_6106,N_6084);
nor U6272 (N_6272,N_6134,N_6019);
nand U6273 (N_6273,N_6154,N_6152);
xor U6274 (N_6274,N_6003,N_6132);
nor U6275 (N_6275,N_6025,N_6062);
nor U6276 (N_6276,N_6160,N_6196);
or U6277 (N_6277,N_6098,N_6186);
xor U6278 (N_6278,N_6189,N_6030);
xnor U6279 (N_6279,N_6039,N_6151);
and U6280 (N_6280,N_6120,N_6086);
xor U6281 (N_6281,N_6118,N_6110);
xor U6282 (N_6282,N_6167,N_6124);
nor U6283 (N_6283,N_6053,N_6178);
xor U6284 (N_6284,N_6093,N_6113);
and U6285 (N_6285,N_6150,N_6161);
nand U6286 (N_6286,N_6121,N_6188);
nand U6287 (N_6287,N_6001,N_6078);
xnor U6288 (N_6288,N_6000,N_6197);
and U6289 (N_6289,N_6145,N_6127);
nor U6290 (N_6290,N_6137,N_6026);
nand U6291 (N_6291,N_6172,N_6020);
or U6292 (N_6292,N_6141,N_6070);
or U6293 (N_6293,N_6119,N_6097);
and U6294 (N_6294,N_6147,N_6096);
nor U6295 (N_6295,N_6133,N_6153);
xnor U6296 (N_6296,N_6067,N_6050);
and U6297 (N_6297,N_6170,N_6131);
and U6298 (N_6298,N_6034,N_6022);
and U6299 (N_6299,N_6136,N_6052);
or U6300 (N_6300,N_6072,N_6108);
and U6301 (N_6301,N_6161,N_6156);
nor U6302 (N_6302,N_6011,N_6101);
and U6303 (N_6303,N_6071,N_6024);
or U6304 (N_6304,N_6030,N_6101);
xor U6305 (N_6305,N_6183,N_6180);
and U6306 (N_6306,N_6044,N_6068);
nand U6307 (N_6307,N_6105,N_6042);
nand U6308 (N_6308,N_6156,N_6003);
nor U6309 (N_6309,N_6047,N_6074);
or U6310 (N_6310,N_6192,N_6180);
or U6311 (N_6311,N_6050,N_6157);
xnor U6312 (N_6312,N_6116,N_6077);
nor U6313 (N_6313,N_6195,N_6177);
xnor U6314 (N_6314,N_6022,N_6172);
nor U6315 (N_6315,N_6090,N_6127);
or U6316 (N_6316,N_6188,N_6153);
xnor U6317 (N_6317,N_6059,N_6096);
or U6318 (N_6318,N_6033,N_6191);
and U6319 (N_6319,N_6030,N_6071);
nor U6320 (N_6320,N_6023,N_6102);
or U6321 (N_6321,N_6077,N_6096);
nor U6322 (N_6322,N_6115,N_6164);
nor U6323 (N_6323,N_6052,N_6106);
and U6324 (N_6324,N_6092,N_6023);
xor U6325 (N_6325,N_6056,N_6152);
or U6326 (N_6326,N_6087,N_6133);
and U6327 (N_6327,N_6067,N_6128);
nand U6328 (N_6328,N_6123,N_6048);
nand U6329 (N_6329,N_6198,N_6131);
or U6330 (N_6330,N_6168,N_6107);
and U6331 (N_6331,N_6089,N_6196);
and U6332 (N_6332,N_6157,N_6012);
xor U6333 (N_6333,N_6121,N_6070);
or U6334 (N_6334,N_6185,N_6122);
or U6335 (N_6335,N_6005,N_6022);
or U6336 (N_6336,N_6159,N_6196);
nand U6337 (N_6337,N_6008,N_6112);
xor U6338 (N_6338,N_6096,N_6186);
xnor U6339 (N_6339,N_6176,N_6175);
or U6340 (N_6340,N_6033,N_6037);
and U6341 (N_6341,N_6152,N_6158);
nand U6342 (N_6342,N_6004,N_6094);
nor U6343 (N_6343,N_6019,N_6081);
nor U6344 (N_6344,N_6163,N_6020);
or U6345 (N_6345,N_6038,N_6074);
or U6346 (N_6346,N_6137,N_6046);
xor U6347 (N_6347,N_6034,N_6173);
nand U6348 (N_6348,N_6153,N_6103);
xnor U6349 (N_6349,N_6109,N_6041);
or U6350 (N_6350,N_6002,N_6056);
or U6351 (N_6351,N_6084,N_6154);
or U6352 (N_6352,N_6064,N_6131);
nand U6353 (N_6353,N_6054,N_6168);
nor U6354 (N_6354,N_6137,N_6078);
xnor U6355 (N_6355,N_6053,N_6033);
or U6356 (N_6356,N_6138,N_6062);
nand U6357 (N_6357,N_6111,N_6118);
xor U6358 (N_6358,N_6099,N_6165);
or U6359 (N_6359,N_6115,N_6159);
nand U6360 (N_6360,N_6106,N_6140);
or U6361 (N_6361,N_6191,N_6101);
nand U6362 (N_6362,N_6143,N_6182);
nor U6363 (N_6363,N_6102,N_6179);
xnor U6364 (N_6364,N_6156,N_6147);
xor U6365 (N_6365,N_6073,N_6174);
and U6366 (N_6366,N_6027,N_6083);
and U6367 (N_6367,N_6163,N_6152);
and U6368 (N_6368,N_6107,N_6105);
nand U6369 (N_6369,N_6169,N_6083);
or U6370 (N_6370,N_6136,N_6074);
and U6371 (N_6371,N_6015,N_6112);
nor U6372 (N_6372,N_6066,N_6108);
or U6373 (N_6373,N_6058,N_6056);
xor U6374 (N_6374,N_6032,N_6189);
nand U6375 (N_6375,N_6195,N_6024);
xnor U6376 (N_6376,N_6023,N_6078);
or U6377 (N_6377,N_6151,N_6061);
nand U6378 (N_6378,N_6169,N_6102);
nor U6379 (N_6379,N_6004,N_6032);
nor U6380 (N_6380,N_6163,N_6023);
or U6381 (N_6381,N_6028,N_6013);
xor U6382 (N_6382,N_6008,N_6140);
and U6383 (N_6383,N_6170,N_6171);
and U6384 (N_6384,N_6171,N_6094);
or U6385 (N_6385,N_6126,N_6056);
nor U6386 (N_6386,N_6152,N_6036);
and U6387 (N_6387,N_6189,N_6038);
nand U6388 (N_6388,N_6119,N_6059);
nand U6389 (N_6389,N_6127,N_6108);
nand U6390 (N_6390,N_6081,N_6002);
or U6391 (N_6391,N_6012,N_6043);
and U6392 (N_6392,N_6077,N_6054);
xnor U6393 (N_6393,N_6029,N_6137);
nand U6394 (N_6394,N_6125,N_6048);
nor U6395 (N_6395,N_6069,N_6101);
and U6396 (N_6396,N_6042,N_6135);
xor U6397 (N_6397,N_6166,N_6040);
and U6398 (N_6398,N_6104,N_6148);
and U6399 (N_6399,N_6069,N_6145);
xor U6400 (N_6400,N_6283,N_6299);
xor U6401 (N_6401,N_6254,N_6211);
and U6402 (N_6402,N_6257,N_6262);
nand U6403 (N_6403,N_6301,N_6365);
nand U6404 (N_6404,N_6368,N_6291);
nor U6405 (N_6405,N_6286,N_6242);
or U6406 (N_6406,N_6247,N_6230);
or U6407 (N_6407,N_6349,N_6369);
nor U6408 (N_6408,N_6295,N_6231);
xor U6409 (N_6409,N_6285,N_6320);
nand U6410 (N_6410,N_6215,N_6228);
or U6411 (N_6411,N_6281,N_6225);
nand U6412 (N_6412,N_6219,N_6212);
nor U6413 (N_6413,N_6278,N_6246);
and U6414 (N_6414,N_6364,N_6352);
nor U6415 (N_6415,N_6380,N_6378);
or U6416 (N_6416,N_6294,N_6233);
nor U6417 (N_6417,N_6213,N_6298);
or U6418 (N_6418,N_6336,N_6297);
nor U6419 (N_6419,N_6379,N_6326);
or U6420 (N_6420,N_6385,N_6355);
and U6421 (N_6421,N_6389,N_6370);
or U6422 (N_6422,N_6248,N_6358);
or U6423 (N_6423,N_6338,N_6396);
and U6424 (N_6424,N_6393,N_6284);
nor U6425 (N_6425,N_6333,N_6209);
or U6426 (N_6426,N_6207,N_6204);
xor U6427 (N_6427,N_6328,N_6245);
nor U6428 (N_6428,N_6282,N_6392);
or U6429 (N_6429,N_6322,N_6305);
xor U6430 (N_6430,N_6376,N_6271);
xnor U6431 (N_6431,N_6201,N_6388);
nand U6432 (N_6432,N_6210,N_6224);
nand U6433 (N_6433,N_6335,N_6239);
xor U6434 (N_6434,N_6311,N_6258);
and U6435 (N_6435,N_6243,N_6289);
xnor U6436 (N_6436,N_6259,N_6309);
or U6437 (N_6437,N_6202,N_6325);
and U6438 (N_6438,N_6268,N_6218);
xnor U6439 (N_6439,N_6316,N_6321);
nand U6440 (N_6440,N_6237,N_6390);
or U6441 (N_6441,N_6312,N_6354);
nor U6442 (N_6442,N_6363,N_6252);
or U6443 (N_6443,N_6310,N_6366);
xor U6444 (N_6444,N_6220,N_6275);
and U6445 (N_6445,N_6357,N_6266);
and U6446 (N_6446,N_6250,N_6342);
or U6447 (N_6447,N_6300,N_6323);
xnor U6448 (N_6448,N_6223,N_6375);
nand U6449 (N_6449,N_6332,N_6399);
nor U6450 (N_6450,N_6315,N_6350);
xnor U6451 (N_6451,N_6339,N_6361);
and U6452 (N_6452,N_6234,N_6372);
nand U6453 (N_6453,N_6255,N_6217);
or U6454 (N_6454,N_6308,N_6253);
and U6455 (N_6455,N_6249,N_6270);
nand U6456 (N_6456,N_6344,N_6306);
xnor U6457 (N_6457,N_6373,N_6334);
nor U6458 (N_6458,N_6324,N_6203);
and U6459 (N_6459,N_6235,N_6327);
nor U6460 (N_6460,N_6331,N_6329);
nor U6461 (N_6461,N_6341,N_6314);
xnor U6462 (N_6462,N_6229,N_6232);
nor U6463 (N_6463,N_6387,N_6391);
and U6464 (N_6464,N_6359,N_6345);
nand U6465 (N_6465,N_6296,N_6280);
and U6466 (N_6466,N_6276,N_6353);
xor U6467 (N_6467,N_6360,N_6302);
xnor U6468 (N_6468,N_6371,N_6265);
and U6469 (N_6469,N_6227,N_6240);
and U6470 (N_6470,N_6290,N_6304);
or U6471 (N_6471,N_6288,N_6381);
nand U6472 (N_6472,N_6395,N_6398);
nand U6473 (N_6473,N_6293,N_6362);
xnor U6474 (N_6474,N_6330,N_6251);
and U6475 (N_6475,N_6317,N_6356);
xor U6476 (N_6476,N_6244,N_6241);
nor U6477 (N_6477,N_6337,N_6307);
xor U6478 (N_6478,N_6384,N_6263);
xor U6479 (N_6479,N_6397,N_6216);
or U6480 (N_6480,N_6319,N_6292);
and U6481 (N_6481,N_6269,N_6222);
or U6482 (N_6482,N_6238,N_6382);
or U6483 (N_6483,N_6206,N_6340);
nand U6484 (N_6484,N_6214,N_6303);
nand U6485 (N_6485,N_6374,N_6272);
xor U6486 (N_6486,N_6256,N_6261);
and U6487 (N_6487,N_6273,N_6394);
and U6488 (N_6488,N_6351,N_6386);
nand U6489 (N_6489,N_6208,N_6260);
xnor U6490 (N_6490,N_6377,N_6205);
nor U6491 (N_6491,N_6348,N_6226);
or U6492 (N_6492,N_6346,N_6267);
nand U6493 (N_6493,N_6200,N_6383);
or U6494 (N_6494,N_6279,N_6343);
xor U6495 (N_6495,N_6367,N_6264);
and U6496 (N_6496,N_6347,N_6236);
nand U6497 (N_6497,N_6287,N_6313);
and U6498 (N_6498,N_6221,N_6274);
or U6499 (N_6499,N_6277,N_6318);
or U6500 (N_6500,N_6367,N_6209);
or U6501 (N_6501,N_6296,N_6367);
and U6502 (N_6502,N_6252,N_6356);
nor U6503 (N_6503,N_6312,N_6202);
xnor U6504 (N_6504,N_6332,N_6281);
nand U6505 (N_6505,N_6372,N_6239);
nand U6506 (N_6506,N_6252,N_6376);
nor U6507 (N_6507,N_6389,N_6322);
xor U6508 (N_6508,N_6231,N_6292);
nor U6509 (N_6509,N_6304,N_6303);
or U6510 (N_6510,N_6217,N_6306);
nor U6511 (N_6511,N_6225,N_6262);
or U6512 (N_6512,N_6298,N_6225);
nor U6513 (N_6513,N_6359,N_6291);
nor U6514 (N_6514,N_6294,N_6346);
nor U6515 (N_6515,N_6328,N_6211);
nor U6516 (N_6516,N_6372,N_6241);
xnor U6517 (N_6517,N_6356,N_6215);
xnor U6518 (N_6518,N_6213,N_6327);
xnor U6519 (N_6519,N_6382,N_6267);
nand U6520 (N_6520,N_6274,N_6344);
and U6521 (N_6521,N_6206,N_6375);
xor U6522 (N_6522,N_6274,N_6363);
or U6523 (N_6523,N_6320,N_6396);
xor U6524 (N_6524,N_6389,N_6330);
xnor U6525 (N_6525,N_6231,N_6357);
xor U6526 (N_6526,N_6299,N_6384);
nand U6527 (N_6527,N_6380,N_6318);
nand U6528 (N_6528,N_6252,N_6305);
nand U6529 (N_6529,N_6213,N_6349);
nand U6530 (N_6530,N_6276,N_6366);
nand U6531 (N_6531,N_6213,N_6332);
xor U6532 (N_6532,N_6206,N_6395);
nand U6533 (N_6533,N_6243,N_6237);
or U6534 (N_6534,N_6223,N_6351);
and U6535 (N_6535,N_6291,N_6248);
xnor U6536 (N_6536,N_6294,N_6343);
and U6537 (N_6537,N_6253,N_6204);
or U6538 (N_6538,N_6268,N_6349);
nand U6539 (N_6539,N_6273,N_6354);
xor U6540 (N_6540,N_6290,N_6203);
xnor U6541 (N_6541,N_6202,N_6223);
xnor U6542 (N_6542,N_6234,N_6253);
and U6543 (N_6543,N_6202,N_6200);
and U6544 (N_6544,N_6396,N_6341);
nand U6545 (N_6545,N_6395,N_6262);
and U6546 (N_6546,N_6203,N_6202);
nor U6547 (N_6547,N_6362,N_6358);
nand U6548 (N_6548,N_6327,N_6322);
nor U6549 (N_6549,N_6235,N_6381);
nor U6550 (N_6550,N_6343,N_6233);
nor U6551 (N_6551,N_6305,N_6361);
nor U6552 (N_6552,N_6333,N_6283);
or U6553 (N_6553,N_6393,N_6232);
nor U6554 (N_6554,N_6243,N_6255);
and U6555 (N_6555,N_6236,N_6359);
and U6556 (N_6556,N_6290,N_6359);
nor U6557 (N_6557,N_6254,N_6210);
or U6558 (N_6558,N_6231,N_6358);
and U6559 (N_6559,N_6244,N_6257);
nor U6560 (N_6560,N_6373,N_6340);
or U6561 (N_6561,N_6275,N_6236);
or U6562 (N_6562,N_6393,N_6377);
xor U6563 (N_6563,N_6309,N_6277);
nand U6564 (N_6564,N_6386,N_6213);
nand U6565 (N_6565,N_6338,N_6258);
nand U6566 (N_6566,N_6310,N_6202);
nor U6567 (N_6567,N_6247,N_6369);
and U6568 (N_6568,N_6374,N_6226);
xnor U6569 (N_6569,N_6300,N_6274);
or U6570 (N_6570,N_6225,N_6305);
xnor U6571 (N_6571,N_6289,N_6206);
nor U6572 (N_6572,N_6374,N_6326);
or U6573 (N_6573,N_6289,N_6216);
nor U6574 (N_6574,N_6271,N_6358);
or U6575 (N_6575,N_6300,N_6321);
xnor U6576 (N_6576,N_6326,N_6249);
and U6577 (N_6577,N_6340,N_6236);
or U6578 (N_6578,N_6304,N_6224);
or U6579 (N_6579,N_6353,N_6211);
or U6580 (N_6580,N_6367,N_6253);
nand U6581 (N_6581,N_6201,N_6390);
or U6582 (N_6582,N_6229,N_6333);
xnor U6583 (N_6583,N_6216,N_6288);
xnor U6584 (N_6584,N_6205,N_6381);
and U6585 (N_6585,N_6218,N_6329);
or U6586 (N_6586,N_6255,N_6394);
nor U6587 (N_6587,N_6242,N_6243);
or U6588 (N_6588,N_6218,N_6291);
nand U6589 (N_6589,N_6217,N_6250);
or U6590 (N_6590,N_6280,N_6362);
nand U6591 (N_6591,N_6396,N_6273);
nor U6592 (N_6592,N_6288,N_6252);
or U6593 (N_6593,N_6248,N_6237);
nand U6594 (N_6594,N_6236,N_6313);
nand U6595 (N_6595,N_6247,N_6324);
nor U6596 (N_6596,N_6200,N_6261);
and U6597 (N_6597,N_6285,N_6231);
and U6598 (N_6598,N_6374,N_6308);
nand U6599 (N_6599,N_6341,N_6259);
and U6600 (N_6600,N_6496,N_6461);
xnor U6601 (N_6601,N_6446,N_6534);
and U6602 (N_6602,N_6441,N_6532);
xnor U6603 (N_6603,N_6445,N_6504);
xnor U6604 (N_6604,N_6573,N_6512);
xor U6605 (N_6605,N_6481,N_6550);
nor U6606 (N_6606,N_6588,N_6572);
xnor U6607 (N_6607,N_6569,N_6505);
nor U6608 (N_6608,N_6564,N_6474);
xor U6609 (N_6609,N_6570,N_6423);
and U6610 (N_6610,N_6462,N_6459);
xor U6611 (N_6611,N_6475,N_6428);
xor U6612 (N_6612,N_6530,N_6528);
or U6613 (N_6613,N_6408,N_6400);
and U6614 (N_6614,N_6472,N_6576);
nor U6615 (N_6615,N_6574,N_6566);
nor U6616 (N_6616,N_6458,N_6582);
nand U6617 (N_6617,N_6490,N_6448);
and U6618 (N_6618,N_6430,N_6575);
nor U6619 (N_6619,N_6546,N_6467);
xnor U6620 (N_6620,N_6452,N_6523);
nand U6621 (N_6621,N_6488,N_6536);
nor U6622 (N_6622,N_6509,N_6561);
nor U6623 (N_6623,N_6513,N_6497);
nor U6624 (N_6624,N_6439,N_6544);
or U6625 (N_6625,N_6501,N_6495);
nor U6626 (N_6626,N_6436,N_6421);
and U6627 (N_6627,N_6487,N_6471);
and U6628 (N_6628,N_6407,N_6485);
and U6629 (N_6629,N_6547,N_6560);
xor U6630 (N_6630,N_6577,N_6466);
nor U6631 (N_6631,N_6537,N_6585);
xnor U6632 (N_6632,N_6579,N_6420);
nand U6633 (N_6633,N_6508,N_6522);
and U6634 (N_6634,N_6412,N_6568);
nor U6635 (N_6635,N_6533,N_6514);
or U6636 (N_6636,N_6595,N_6404);
or U6637 (N_6637,N_6593,N_6596);
nand U6638 (N_6638,N_6415,N_6493);
or U6639 (N_6639,N_6525,N_6469);
or U6640 (N_6640,N_6411,N_6492);
nor U6641 (N_6641,N_6431,N_6507);
xnor U6642 (N_6642,N_6498,N_6451);
nor U6643 (N_6643,N_6516,N_6456);
nor U6644 (N_6644,N_6586,N_6535);
nand U6645 (N_6645,N_6410,N_6597);
and U6646 (N_6646,N_6491,N_6552);
or U6647 (N_6647,N_6540,N_6539);
or U6648 (N_6648,N_6524,N_6417);
or U6649 (N_6649,N_6418,N_6478);
or U6650 (N_6650,N_6480,N_6506);
and U6651 (N_6651,N_6494,N_6444);
nor U6652 (N_6652,N_6482,N_6538);
and U6653 (N_6653,N_6580,N_6425);
xor U6654 (N_6654,N_6435,N_6434);
xnor U6655 (N_6655,N_6521,N_6542);
or U6656 (N_6656,N_6598,N_6565);
or U6657 (N_6657,N_6587,N_6571);
xor U6658 (N_6658,N_6432,N_6527);
or U6659 (N_6659,N_6479,N_6548);
and U6660 (N_6660,N_6454,N_6515);
nand U6661 (N_6661,N_6558,N_6510);
nor U6662 (N_6662,N_6464,N_6594);
and U6663 (N_6663,N_6402,N_6465);
nor U6664 (N_6664,N_6406,N_6589);
or U6665 (N_6665,N_6419,N_6405);
nor U6666 (N_6666,N_6557,N_6590);
nor U6667 (N_6667,N_6483,N_6486);
nand U6668 (N_6668,N_6545,N_6442);
nor U6669 (N_6669,N_6567,N_6519);
nor U6670 (N_6670,N_6457,N_6551);
or U6671 (N_6671,N_6424,N_6591);
nor U6672 (N_6672,N_6447,N_6460);
or U6673 (N_6673,N_6592,N_6581);
nand U6674 (N_6674,N_6518,N_6543);
nand U6675 (N_6675,N_6450,N_6531);
xnor U6676 (N_6676,N_6541,N_6453);
xor U6677 (N_6677,N_6529,N_6455);
and U6678 (N_6678,N_6555,N_6429);
or U6679 (N_6679,N_6440,N_6584);
xor U6680 (N_6680,N_6437,N_6463);
and U6681 (N_6681,N_6489,N_6401);
xor U6682 (N_6682,N_6438,N_6416);
and U6683 (N_6683,N_6553,N_6520);
or U6684 (N_6684,N_6426,N_6500);
or U6685 (N_6685,N_6559,N_6477);
nand U6686 (N_6686,N_6409,N_6403);
or U6687 (N_6687,N_6468,N_6422);
nand U6688 (N_6688,N_6503,N_6517);
or U6689 (N_6689,N_6583,N_6578);
and U6690 (N_6690,N_6511,N_6413);
xnor U6691 (N_6691,N_6470,N_6549);
xor U6692 (N_6692,N_6433,N_6484);
or U6693 (N_6693,N_6449,N_6476);
xor U6694 (N_6694,N_6414,N_6563);
and U6695 (N_6695,N_6562,N_6499);
nand U6696 (N_6696,N_6502,N_6443);
xor U6697 (N_6697,N_6556,N_6473);
xnor U6698 (N_6698,N_6427,N_6599);
or U6699 (N_6699,N_6554,N_6526);
and U6700 (N_6700,N_6481,N_6575);
xor U6701 (N_6701,N_6431,N_6516);
xnor U6702 (N_6702,N_6592,N_6447);
nand U6703 (N_6703,N_6494,N_6534);
and U6704 (N_6704,N_6546,N_6524);
nor U6705 (N_6705,N_6577,N_6494);
and U6706 (N_6706,N_6565,N_6529);
and U6707 (N_6707,N_6592,N_6570);
nand U6708 (N_6708,N_6404,N_6437);
or U6709 (N_6709,N_6438,N_6582);
xnor U6710 (N_6710,N_6459,N_6439);
xnor U6711 (N_6711,N_6550,N_6448);
and U6712 (N_6712,N_6552,N_6544);
or U6713 (N_6713,N_6492,N_6559);
or U6714 (N_6714,N_6505,N_6498);
or U6715 (N_6715,N_6401,N_6436);
nand U6716 (N_6716,N_6594,N_6406);
nor U6717 (N_6717,N_6475,N_6457);
or U6718 (N_6718,N_6537,N_6533);
xor U6719 (N_6719,N_6543,N_6479);
nand U6720 (N_6720,N_6597,N_6459);
and U6721 (N_6721,N_6526,N_6585);
and U6722 (N_6722,N_6414,N_6493);
nand U6723 (N_6723,N_6475,N_6537);
or U6724 (N_6724,N_6584,N_6446);
xnor U6725 (N_6725,N_6547,N_6584);
or U6726 (N_6726,N_6518,N_6513);
xor U6727 (N_6727,N_6570,N_6543);
xor U6728 (N_6728,N_6422,N_6589);
nand U6729 (N_6729,N_6536,N_6429);
xnor U6730 (N_6730,N_6590,N_6561);
nand U6731 (N_6731,N_6414,N_6497);
nor U6732 (N_6732,N_6447,N_6508);
and U6733 (N_6733,N_6547,N_6447);
or U6734 (N_6734,N_6542,N_6594);
or U6735 (N_6735,N_6495,N_6454);
nand U6736 (N_6736,N_6508,N_6424);
xnor U6737 (N_6737,N_6594,N_6418);
xnor U6738 (N_6738,N_6527,N_6486);
nand U6739 (N_6739,N_6450,N_6498);
or U6740 (N_6740,N_6443,N_6460);
or U6741 (N_6741,N_6570,N_6502);
and U6742 (N_6742,N_6414,N_6492);
nor U6743 (N_6743,N_6484,N_6535);
nand U6744 (N_6744,N_6548,N_6584);
and U6745 (N_6745,N_6489,N_6576);
or U6746 (N_6746,N_6437,N_6571);
xnor U6747 (N_6747,N_6542,N_6404);
or U6748 (N_6748,N_6535,N_6466);
and U6749 (N_6749,N_6567,N_6537);
xor U6750 (N_6750,N_6596,N_6472);
nor U6751 (N_6751,N_6424,N_6496);
nor U6752 (N_6752,N_6440,N_6481);
nand U6753 (N_6753,N_6428,N_6406);
nor U6754 (N_6754,N_6518,N_6583);
or U6755 (N_6755,N_6485,N_6444);
xnor U6756 (N_6756,N_6502,N_6455);
nand U6757 (N_6757,N_6429,N_6570);
and U6758 (N_6758,N_6509,N_6430);
and U6759 (N_6759,N_6411,N_6521);
nor U6760 (N_6760,N_6457,N_6543);
xnor U6761 (N_6761,N_6584,N_6538);
nor U6762 (N_6762,N_6472,N_6529);
xor U6763 (N_6763,N_6408,N_6491);
or U6764 (N_6764,N_6499,N_6568);
nand U6765 (N_6765,N_6586,N_6563);
nand U6766 (N_6766,N_6551,N_6552);
nor U6767 (N_6767,N_6435,N_6471);
xor U6768 (N_6768,N_6556,N_6446);
and U6769 (N_6769,N_6465,N_6543);
nand U6770 (N_6770,N_6404,N_6510);
or U6771 (N_6771,N_6461,N_6445);
nor U6772 (N_6772,N_6502,N_6558);
and U6773 (N_6773,N_6401,N_6586);
nand U6774 (N_6774,N_6480,N_6502);
or U6775 (N_6775,N_6509,N_6467);
nor U6776 (N_6776,N_6427,N_6566);
nand U6777 (N_6777,N_6558,N_6595);
and U6778 (N_6778,N_6417,N_6511);
xor U6779 (N_6779,N_6404,N_6468);
and U6780 (N_6780,N_6490,N_6598);
and U6781 (N_6781,N_6520,N_6452);
xnor U6782 (N_6782,N_6458,N_6490);
xnor U6783 (N_6783,N_6428,N_6436);
and U6784 (N_6784,N_6544,N_6498);
nand U6785 (N_6785,N_6572,N_6472);
or U6786 (N_6786,N_6440,N_6593);
nor U6787 (N_6787,N_6590,N_6455);
and U6788 (N_6788,N_6566,N_6569);
nor U6789 (N_6789,N_6442,N_6424);
nor U6790 (N_6790,N_6496,N_6596);
nand U6791 (N_6791,N_6411,N_6528);
and U6792 (N_6792,N_6454,N_6594);
and U6793 (N_6793,N_6463,N_6451);
or U6794 (N_6794,N_6567,N_6517);
or U6795 (N_6795,N_6506,N_6561);
and U6796 (N_6796,N_6426,N_6538);
xnor U6797 (N_6797,N_6486,N_6549);
or U6798 (N_6798,N_6595,N_6505);
and U6799 (N_6799,N_6438,N_6524);
and U6800 (N_6800,N_6728,N_6770);
and U6801 (N_6801,N_6704,N_6723);
nand U6802 (N_6802,N_6603,N_6715);
xor U6803 (N_6803,N_6610,N_6739);
xor U6804 (N_6804,N_6626,N_6689);
nor U6805 (N_6805,N_6780,N_6729);
and U6806 (N_6806,N_6787,N_6743);
nor U6807 (N_6807,N_6751,N_6662);
and U6808 (N_6808,N_6684,N_6675);
nand U6809 (N_6809,N_6660,N_6763);
and U6810 (N_6810,N_6627,N_6771);
nand U6811 (N_6811,N_6734,N_6764);
xor U6812 (N_6812,N_6732,N_6676);
and U6813 (N_6813,N_6776,N_6657);
or U6814 (N_6814,N_6719,N_6693);
nor U6815 (N_6815,N_6744,N_6621);
nor U6816 (N_6816,N_6637,N_6775);
nand U6817 (N_6817,N_6714,N_6712);
and U6818 (N_6818,N_6685,N_6761);
xnor U6819 (N_6819,N_6798,N_6613);
xor U6820 (N_6820,N_6773,N_6651);
xnor U6821 (N_6821,N_6717,N_6654);
nand U6822 (N_6822,N_6788,N_6791);
nand U6823 (N_6823,N_6768,N_6674);
and U6824 (N_6824,N_6686,N_6725);
xnor U6825 (N_6825,N_6633,N_6606);
xnor U6826 (N_6826,N_6741,N_6797);
xnor U6827 (N_6827,N_6647,N_6671);
and U6828 (N_6828,N_6778,N_6696);
xor U6829 (N_6829,N_6716,N_6783);
nor U6830 (N_6830,N_6666,N_6668);
nor U6831 (N_6831,N_6672,N_6615);
nor U6832 (N_6832,N_6738,N_6635);
or U6833 (N_6833,N_6740,N_6745);
nand U6834 (N_6834,N_6694,N_6638);
nor U6835 (N_6835,N_6653,N_6730);
nand U6836 (N_6836,N_6752,N_6681);
nor U6837 (N_6837,N_6656,N_6750);
nand U6838 (N_6838,N_6644,N_6746);
xor U6839 (N_6839,N_6659,N_6619);
nor U6840 (N_6840,N_6616,N_6697);
or U6841 (N_6841,N_6756,N_6663);
nand U6842 (N_6842,N_6604,N_6785);
and U6843 (N_6843,N_6683,N_6782);
nor U6844 (N_6844,N_6630,N_6688);
or U6845 (N_6845,N_6608,N_6641);
and U6846 (N_6846,N_6648,N_6677);
or U6847 (N_6847,N_6735,N_6699);
xnor U6848 (N_6848,N_6720,N_6607);
and U6849 (N_6849,N_6624,N_6792);
nor U6850 (N_6850,N_6611,N_6731);
and U6851 (N_6851,N_6636,N_6755);
nand U6852 (N_6852,N_6758,N_6767);
nor U6853 (N_6853,N_6760,N_6625);
xor U6854 (N_6854,N_6747,N_6678);
nor U6855 (N_6855,N_6667,N_6779);
xnor U6856 (N_6856,N_6799,N_6661);
nand U6857 (N_6857,N_6742,N_6679);
nor U6858 (N_6858,N_6658,N_6777);
and U6859 (N_6859,N_6759,N_6701);
xor U6860 (N_6860,N_6706,N_6774);
xor U6861 (N_6861,N_6794,N_6665);
nand U6862 (N_6862,N_6722,N_6650);
nand U6863 (N_6863,N_6602,N_6691);
or U6864 (N_6864,N_6727,N_6737);
nor U6865 (N_6865,N_6707,N_6772);
nand U6866 (N_6866,N_6762,N_6639);
nand U6867 (N_6867,N_6784,N_6605);
or U6868 (N_6868,N_6631,N_6640);
or U6869 (N_6869,N_6645,N_6664);
nand U6870 (N_6870,N_6692,N_6702);
and U6871 (N_6871,N_6623,N_6700);
nor U6872 (N_6872,N_6690,N_6786);
xnor U6873 (N_6873,N_6670,N_6673);
or U6874 (N_6874,N_6749,N_6753);
nor U6875 (N_6875,N_6680,N_6682);
nor U6876 (N_6876,N_6687,N_6726);
nor U6877 (N_6877,N_6622,N_6614);
xnor U6878 (N_6878,N_6609,N_6793);
xor U6879 (N_6879,N_6620,N_6748);
nand U6880 (N_6880,N_6646,N_6669);
nor U6881 (N_6881,N_6769,N_6710);
xor U6882 (N_6882,N_6757,N_6618);
or U6883 (N_6883,N_6789,N_6754);
xor U6884 (N_6884,N_6632,N_6766);
nand U6885 (N_6885,N_6709,N_6617);
nand U6886 (N_6886,N_6711,N_6698);
nor U6887 (N_6887,N_6652,N_6629);
xor U6888 (N_6888,N_6695,N_6649);
nand U6889 (N_6889,N_6601,N_6655);
xor U6890 (N_6890,N_6713,N_6705);
nor U6891 (N_6891,N_6721,N_6628);
or U6892 (N_6892,N_6718,N_6708);
or U6893 (N_6893,N_6733,N_6736);
nand U6894 (N_6894,N_6600,N_6643);
or U6895 (N_6895,N_6612,N_6642);
xnor U6896 (N_6896,N_6724,N_6796);
or U6897 (N_6897,N_6634,N_6781);
and U6898 (N_6898,N_6790,N_6765);
nor U6899 (N_6899,N_6795,N_6703);
nand U6900 (N_6900,N_6746,N_6775);
xor U6901 (N_6901,N_6691,N_6751);
xor U6902 (N_6902,N_6773,N_6670);
xnor U6903 (N_6903,N_6621,N_6746);
or U6904 (N_6904,N_6688,N_6671);
or U6905 (N_6905,N_6684,N_6673);
or U6906 (N_6906,N_6770,N_6649);
or U6907 (N_6907,N_6788,N_6789);
nand U6908 (N_6908,N_6683,N_6744);
nor U6909 (N_6909,N_6692,N_6716);
nor U6910 (N_6910,N_6723,N_6644);
nor U6911 (N_6911,N_6748,N_6731);
nand U6912 (N_6912,N_6653,N_6796);
and U6913 (N_6913,N_6647,N_6634);
or U6914 (N_6914,N_6691,N_6607);
xnor U6915 (N_6915,N_6734,N_6747);
and U6916 (N_6916,N_6785,N_6786);
or U6917 (N_6917,N_6711,N_6710);
nand U6918 (N_6918,N_6669,N_6715);
or U6919 (N_6919,N_6742,N_6707);
nand U6920 (N_6920,N_6684,N_6722);
nand U6921 (N_6921,N_6603,N_6749);
xnor U6922 (N_6922,N_6690,N_6735);
and U6923 (N_6923,N_6667,N_6634);
or U6924 (N_6924,N_6627,N_6625);
nor U6925 (N_6925,N_6681,N_6793);
or U6926 (N_6926,N_6701,N_6627);
nand U6927 (N_6927,N_6624,N_6799);
nor U6928 (N_6928,N_6788,N_6652);
and U6929 (N_6929,N_6770,N_6724);
and U6930 (N_6930,N_6787,N_6605);
or U6931 (N_6931,N_6772,N_6709);
and U6932 (N_6932,N_6625,N_6649);
or U6933 (N_6933,N_6764,N_6629);
nand U6934 (N_6934,N_6711,N_6728);
nand U6935 (N_6935,N_6795,N_6638);
or U6936 (N_6936,N_6639,N_6653);
nand U6937 (N_6937,N_6791,N_6637);
and U6938 (N_6938,N_6730,N_6721);
or U6939 (N_6939,N_6691,N_6720);
xnor U6940 (N_6940,N_6704,N_6661);
and U6941 (N_6941,N_6632,N_6793);
nor U6942 (N_6942,N_6666,N_6663);
nor U6943 (N_6943,N_6679,N_6703);
and U6944 (N_6944,N_6766,N_6741);
nand U6945 (N_6945,N_6779,N_6600);
nand U6946 (N_6946,N_6666,N_6657);
nor U6947 (N_6947,N_6767,N_6675);
and U6948 (N_6948,N_6668,N_6640);
or U6949 (N_6949,N_6741,N_6750);
or U6950 (N_6950,N_6788,N_6710);
nor U6951 (N_6951,N_6625,N_6662);
and U6952 (N_6952,N_6634,N_6612);
nand U6953 (N_6953,N_6626,N_6713);
xor U6954 (N_6954,N_6691,N_6768);
nand U6955 (N_6955,N_6602,N_6743);
nand U6956 (N_6956,N_6790,N_6758);
xor U6957 (N_6957,N_6746,N_6790);
nand U6958 (N_6958,N_6758,N_6784);
and U6959 (N_6959,N_6645,N_6667);
and U6960 (N_6960,N_6610,N_6771);
or U6961 (N_6961,N_6638,N_6753);
or U6962 (N_6962,N_6784,N_6636);
nor U6963 (N_6963,N_6706,N_6744);
and U6964 (N_6964,N_6614,N_6767);
nor U6965 (N_6965,N_6720,N_6692);
and U6966 (N_6966,N_6767,N_6780);
or U6967 (N_6967,N_6781,N_6641);
or U6968 (N_6968,N_6756,N_6641);
nand U6969 (N_6969,N_6621,N_6649);
xnor U6970 (N_6970,N_6768,N_6785);
nor U6971 (N_6971,N_6617,N_6773);
and U6972 (N_6972,N_6678,N_6702);
xnor U6973 (N_6973,N_6677,N_6675);
nand U6974 (N_6974,N_6705,N_6770);
or U6975 (N_6975,N_6789,N_6729);
nand U6976 (N_6976,N_6683,N_6650);
and U6977 (N_6977,N_6662,N_6776);
and U6978 (N_6978,N_6747,N_6693);
and U6979 (N_6979,N_6774,N_6714);
nand U6980 (N_6980,N_6689,N_6765);
nor U6981 (N_6981,N_6673,N_6722);
nand U6982 (N_6982,N_6708,N_6618);
nor U6983 (N_6983,N_6762,N_6710);
or U6984 (N_6984,N_6608,N_6776);
nand U6985 (N_6985,N_6763,N_6665);
nor U6986 (N_6986,N_6611,N_6671);
xor U6987 (N_6987,N_6602,N_6687);
xnor U6988 (N_6988,N_6714,N_6775);
and U6989 (N_6989,N_6783,N_6705);
or U6990 (N_6990,N_6763,N_6750);
or U6991 (N_6991,N_6707,N_6709);
and U6992 (N_6992,N_6733,N_6767);
nor U6993 (N_6993,N_6607,N_6690);
nand U6994 (N_6994,N_6662,N_6709);
or U6995 (N_6995,N_6750,N_6753);
and U6996 (N_6996,N_6639,N_6743);
nor U6997 (N_6997,N_6702,N_6737);
and U6998 (N_6998,N_6736,N_6776);
xor U6999 (N_6999,N_6783,N_6789);
nand U7000 (N_7000,N_6895,N_6894);
nand U7001 (N_7001,N_6846,N_6928);
and U7002 (N_7002,N_6879,N_6955);
nand U7003 (N_7003,N_6976,N_6810);
xnor U7004 (N_7004,N_6917,N_6864);
and U7005 (N_7005,N_6890,N_6885);
nand U7006 (N_7006,N_6823,N_6907);
nor U7007 (N_7007,N_6912,N_6877);
xor U7008 (N_7008,N_6868,N_6874);
and U7009 (N_7009,N_6978,N_6816);
or U7010 (N_7010,N_6909,N_6977);
and U7011 (N_7011,N_6880,N_6971);
nor U7012 (N_7012,N_6830,N_6944);
and U7013 (N_7013,N_6964,N_6819);
nand U7014 (N_7014,N_6925,N_6916);
xnor U7015 (N_7015,N_6870,N_6869);
nor U7016 (N_7016,N_6815,N_6800);
xor U7017 (N_7017,N_6973,N_6833);
nand U7018 (N_7018,N_6991,N_6886);
or U7019 (N_7019,N_6999,N_6838);
nand U7020 (N_7020,N_6935,N_6959);
xor U7021 (N_7021,N_6901,N_6872);
xnor U7022 (N_7022,N_6835,N_6862);
nand U7023 (N_7023,N_6926,N_6986);
xnor U7024 (N_7024,N_6807,N_6873);
nand U7025 (N_7025,N_6858,N_6836);
or U7026 (N_7026,N_6803,N_6826);
xor U7027 (N_7027,N_6906,N_6859);
nand U7028 (N_7028,N_6996,N_6941);
or U7029 (N_7029,N_6811,N_6972);
or U7030 (N_7030,N_6965,N_6841);
nor U7031 (N_7031,N_6905,N_6997);
and U7032 (N_7032,N_6929,N_6855);
nor U7033 (N_7033,N_6891,N_6911);
and U7034 (N_7034,N_6847,N_6831);
and U7035 (N_7035,N_6913,N_6957);
nand U7036 (N_7036,N_6994,N_6893);
xnor U7037 (N_7037,N_6834,N_6939);
and U7038 (N_7038,N_6936,N_6837);
nand U7039 (N_7039,N_6854,N_6861);
xor U7040 (N_7040,N_6923,N_6952);
or U7041 (N_7041,N_6853,N_6949);
and U7042 (N_7042,N_6863,N_6947);
nand U7043 (N_7043,N_6984,N_6968);
or U7044 (N_7044,N_6801,N_6943);
nor U7045 (N_7045,N_6993,N_6808);
or U7046 (N_7046,N_6942,N_6856);
or U7047 (N_7047,N_6883,N_6975);
xor U7048 (N_7048,N_6843,N_6933);
or U7049 (N_7049,N_6802,N_6962);
nor U7050 (N_7050,N_6848,N_6974);
nand U7051 (N_7051,N_6828,N_6887);
and U7052 (N_7052,N_6966,N_6951);
xor U7053 (N_7053,N_6983,N_6931);
xor U7054 (N_7054,N_6938,N_6845);
and U7055 (N_7055,N_6940,N_6820);
or U7056 (N_7056,N_6960,N_6813);
or U7057 (N_7057,N_6981,N_6982);
nor U7058 (N_7058,N_6995,N_6967);
nand U7059 (N_7059,N_6932,N_6956);
or U7060 (N_7060,N_6998,N_6878);
or U7061 (N_7061,N_6817,N_6988);
xor U7062 (N_7062,N_6866,N_6897);
nor U7063 (N_7063,N_6839,N_6822);
xor U7064 (N_7064,N_6805,N_6934);
and U7065 (N_7065,N_6946,N_6892);
or U7066 (N_7066,N_6829,N_6904);
xor U7067 (N_7067,N_6899,N_6961);
nand U7068 (N_7068,N_6958,N_6871);
nor U7069 (N_7069,N_6865,N_6881);
xnor U7070 (N_7070,N_6985,N_6804);
nand U7071 (N_7071,N_6806,N_6954);
or U7072 (N_7072,N_6824,N_6930);
and U7073 (N_7073,N_6849,N_6884);
or U7074 (N_7074,N_6857,N_6896);
nand U7075 (N_7075,N_6852,N_6851);
xnor U7076 (N_7076,N_6987,N_6827);
nand U7077 (N_7077,N_6888,N_6840);
xnor U7078 (N_7078,N_6914,N_6922);
nor U7079 (N_7079,N_6910,N_6950);
or U7080 (N_7080,N_6969,N_6860);
or U7081 (N_7081,N_6963,N_6809);
xor U7082 (N_7082,N_6920,N_6903);
nand U7083 (N_7083,N_6919,N_6867);
nand U7084 (N_7084,N_6915,N_6908);
or U7085 (N_7085,N_6818,N_6924);
or U7086 (N_7086,N_6900,N_6918);
or U7087 (N_7087,N_6825,N_6812);
and U7088 (N_7088,N_6990,N_6821);
nor U7089 (N_7089,N_6927,N_6876);
nor U7090 (N_7090,N_6832,N_6844);
nand U7091 (N_7091,N_6875,N_6889);
or U7092 (N_7092,N_6989,N_6937);
nor U7093 (N_7093,N_6814,N_6902);
or U7094 (N_7094,N_6948,N_6980);
nand U7095 (N_7095,N_6850,N_6898);
xor U7096 (N_7096,N_6921,N_6953);
xor U7097 (N_7097,N_6882,N_6945);
or U7098 (N_7098,N_6970,N_6992);
or U7099 (N_7099,N_6979,N_6842);
or U7100 (N_7100,N_6802,N_6876);
nand U7101 (N_7101,N_6849,N_6886);
and U7102 (N_7102,N_6887,N_6899);
nor U7103 (N_7103,N_6939,N_6807);
or U7104 (N_7104,N_6965,N_6983);
nand U7105 (N_7105,N_6902,N_6867);
or U7106 (N_7106,N_6909,N_6937);
xor U7107 (N_7107,N_6900,N_6922);
or U7108 (N_7108,N_6805,N_6900);
nand U7109 (N_7109,N_6803,N_6862);
and U7110 (N_7110,N_6985,N_6932);
nand U7111 (N_7111,N_6868,N_6864);
xnor U7112 (N_7112,N_6974,N_6830);
or U7113 (N_7113,N_6966,N_6842);
nand U7114 (N_7114,N_6941,N_6987);
nor U7115 (N_7115,N_6846,N_6977);
nor U7116 (N_7116,N_6946,N_6995);
nand U7117 (N_7117,N_6858,N_6956);
nor U7118 (N_7118,N_6865,N_6830);
xor U7119 (N_7119,N_6954,N_6953);
nand U7120 (N_7120,N_6852,N_6951);
nor U7121 (N_7121,N_6833,N_6937);
or U7122 (N_7122,N_6820,N_6840);
nand U7123 (N_7123,N_6938,N_6985);
xnor U7124 (N_7124,N_6920,N_6868);
or U7125 (N_7125,N_6898,N_6833);
nor U7126 (N_7126,N_6915,N_6940);
or U7127 (N_7127,N_6943,N_6900);
or U7128 (N_7128,N_6917,N_6863);
or U7129 (N_7129,N_6958,N_6876);
or U7130 (N_7130,N_6923,N_6847);
xor U7131 (N_7131,N_6968,N_6956);
xnor U7132 (N_7132,N_6982,N_6976);
nor U7133 (N_7133,N_6854,N_6996);
nand U7134 (N_7134,N_6909,N_6919);
or U7135 (N_7135,N_6984,N_6864);
or U7136 (N_7136,N_6857,N_6817);
nor U7137 (N_7137,N_6802,N_6946);
xnor U7138 (N_7138,N_6807,N_6911);
xor U7139 (N_7139,N_6847,N_6996);
and U7140 (N_7140,N_6937,N_6838);
xor U7141 (N_7141,N_6861,N_6824);
nor U7142 (N_7142,N_6998,N_6896);
or U7143 (N_7143,N_6834,N_6940);
nand U7144 (N_7144,N_6860,N_6875);
nor U7145 (N_7145,N_6894,N_6886);
xnor U7146 (N_7146,N_6924,N_6800);
xor U7147 (N_7147,N_6897,N_6813);
xor U7148 (N_7148,N_6930,N_6945);
and U7149 (N_7149,N_6940,N_6833);
and U7150 (N_7150,N_6985,N_6861);
or U7151 (N_7151,N_6805,N_6907);
nand U7152 (N_7152,N_6890,N_6820);
and U7153 (N_7153,N_6999,N_6934);
nand U7154 (N_7154,N_6823,N_6874);
nor U7155 (N_7155,N_6868,N_6862);
nand U7156 (N_7156,N_6955,N_6939);
and U7157 (N_7157,N_6837,N_6873);
and U7158 (N_7158,N_6902,N_6860);
and U7159 (N_7159,N_6980,N_6882);
and U7160 (N_7160,N_6868,N_6905);
or U7161 (N_7161,N_6970,N_6937);
nand U7162 (N_7162,N_6997,N_6957);
nor U7163 (N_7163,N_6840,N_6812);
or U7164 (N_7164,N_6871,N_6996);
nor U7165 (N_7165,N_6937,N_6998);
xnor U7166 (N_7166,N_6917,N_6812);
xor U7167 (N_7167,N_6855,N_6940);
and U7168 (N_7168,N_6884,N_6944);
xnor U7169 (N_7169,N_6910,N_6848);
and U7170 (N_7170,N_6932,N_6971);
nor U7171 (N_7171,N_6932,N_6901);
nor U7172 (N_7172,N_6915,N_6911);
nor U7173 (N_7173,N_6807,N_6982);
nand U7174 (N_7174,N_6837,N_6908);
xor U7175 (N_7175,N_6983,N_6918);
and U7176 (N_7176,N_6976,N_6944);
nor U7177 (N_7177,N_6847,N_6820);
xor U7178 (N_7178,N_6908,N_6949);
or U7179 (N_7179,N_6957,N_6845);
nand U7180 (N_7180,N_6869,N_6927);
or U7181 (N_7181,N_6910,N_6865);
nor U7182 (N_7182,N_6994,N_6957);
nand U7183 (N_7183,N_6858,N_6894);
and U7184 (N_7184,N_6897,N_6983);
or U7185 (N_7185,N_6806,N_6888);
and U7186 (N_7186,N_6887,N_6855);
and U7187 (N_7187,N_6859,N_6984);
and U7188 (N_7188,N_6860,N_6995);
xnor U7189 (N_7189,N_6940,N_6893);
and U7190 (N_7190,N_6904,N_6948);
nor U7191 (N_7191,N_6830,N_6883);
xnor U7192 (N_7192,N_6847,N_6876);
xor U7193 (N_7193,N_6922,N_6933);
nor U7194 (N_7194,N_6853,N_6928);
or U7195 (N_7195,N_6810,N_6887);
or U7196 (N_7196,N_6980,N_6905);
xor U7197 (N_7197,N_6870,N_6940);
nand U7198 (N_7198,N_6892,N_6974);
xor U7199 (N_7199,N_6828,N_6977);
xor U7200 (N_7200,N_7083,N_7181);
or U7201 (N_7201,N_7058,N_7177);
and U7202 (N_7202,N_7105,N_7130);
nand U7203 (N_7203,N_7072,N_7149);
xor U7204 (N_7204,N_7097,N_7123);
nor U7205 (N_7205,N_7001,N_7169);
and U7206 (N_7206,N_7088,N_7156);
and U7207 (N_7207,N_7170,N_7028);
nor U7208 (N_7208,N_7055,N_7132);
and U7209 (N_7209,N_7128,N_7068);
nand U7210 (N_7210,N_7092,N_7114);
nor U7211 (N_7211,N_7095,N_7066);
nor U7212 (N_7212,N_7047,N_7020);
or U7213 (N_7213,N_7137,N_7133);
or U7214 (N_7214,N_7065,N_7050);
xnor U7215 (N_7215,N_7005,N_7030);
or U7216 (N_7216,N_7184,N_7015);
xnor U7217 (N_7217,N_7051,N_7178);
and U7218 (N_7218,N_7032,N_7194);
xnor U7219 (N_7219,N_7035,N_7148);
nor U7220 (N_7220,N_7037,N_7183);
and U7221 (N_7221,N_7111,N_7163);
and U7222 (N_7222,N_7182,N_7011);
nor U7223 (N_7223,N_7171,N_7094);
nand U7224 (N_7224,N_7027,N_7091);
and U7225 (N_7225,N_7101,N_7014);
nor U7226 (N_7226,N_7048,N_7098);
xor U7227 (N_7227,N_7074,N_7168);
nor U7228 (N_7228,N_7008,N_7036);
nand U7229 (N_7229,N_7108,N_7045);
and U7230 (N_7230,N_7084,N_7164);
nor U7231 (N_7231,N_7131,N_7023);
xnor U7232 (N_7232,N_7039,N_7140);
xor U7233 (N_7233,N_7021,N_7063);
nor U7234 (N_7234,N_7079,N_7107);
and U7235 (N_7235,N_7087,N_7049);
nand U7236 (N_7236,N_7176,N_7024);
and U7237 (N_7237,N_7004,N_7086);
or U7238 (N_7238,N_7031,N_7112);
and U7239 (N_7239,N_7025,N_7198);
xor U7240 (N_7240,N_7003,N_7090);
xor U7241 (N_7241,N_7126,N_7153);
nor U7242 (N_7242,N_7010,N_7017);
xnor U7243 (N_7243,N_7062,N_7147);
nand U7244 (N_7244,N_7012,N_7061);
nor U7245 (N_7245,N_7002,N_7117);
and U7246 (N_7246,N_7059,N_7155);
and U7247 (N_7247,N_7009,N_7110);
or U7248 (N_7248,N_7071,N_7185);
or U7249 (N_7249,N_7172,N_7154);
nor U7250 (N_7250,N_7007,N_7077);
nand U7251 (N_7251,N_7122,N_7158);
nor U7252 (N_7252,N_7139,N_7040);
and U7253 (N_7253,N_7142,N_7165);
xor U7254 (N_7254,N_7161,N_7076);
nand U7255 (N_7255,N_7118,N_7042);
xor U7256 (N_7256,N_7067,N_7034);
xor U7257 (N_7257,N_7016,N_7179);
and U7258 (N_7258,N_7113,N_7053);
xor U7259 (N_7259,N_7054,N_7186);
and U7260 (N_7260,N_7115,N_7173);
xor U7261 (N_7261,N_7109,N_7138);
nor U7262 (N_7262,N_7057,N_7141);
or U7263 (N_7263,N_7104,N_7196);
xor U7264 (N_7264,N_7174,N_7099);
or U7265 (N_7265,N_7160,N_7199);
or U7266 (N_7266,N_7124,N_7082);
nand U7267 (N_7267,N_7145,N_7081);
or U7268 (N_7268,N_7120,N_7166);
nor U7269 (N_7269,N_7106,N_7075);
and U7270 (N_7270,N_7080,N_7070);
nor U7271 (N_7271,N_7006,N_7085);
nand U7272 (N_7272,N_7078,N_7000);
nor U7273 (N_7273,N_7193,N_7038);
or U7274 (N_7274,N_7100,N_7102);
xnor U7275 (N_7275,N_7056,N_7129);
or U7276 (N_7276,N_7119,N_7069);
or U7277 (N_7277,N_7022,N_7144);
nand U7278 (N_7278,N_7180,N_7135);
nand U7279 (N_7279,N_7162,N_7064);
and U7280 (N_7280,N_7041,N_7134);
and U7281 (N_7281,N_7018,N_7060);
and U7282 (N_7282,N_7052,N_7096);
and U7283 (N_7283,N_7192,N_7151);
nor U7284 (N_7284,N_7191,N_7073);
or U7285 (N_7285,N_7188,N_7197);
nor U7286 (N_7286,N_7019,N_7033);
nand U7287 (N_7287,N_7195,N_7143);
or U7288 (N_7288,N_7146,N_7013);
or U7289 (N_7289,N_7026,N_7190);
and U7290 (N_7290,N_7152,N_7159);
and U7291 (N_7291,N_7093,N_7150);
or U7292 (N_7292,N_7121,N_7157);
nor U7293 (N_7293,N_7189,N_7127);
or U7294 (N_7294,N_7116,N_7043);
xor U7295 (N_7295,N_7167,N_7044);
nand U7296 (N_7296,N_7029,N_7046);
or U7297 (N_7297,N_7136,N_7103);
and U7298 (N_7298,N_7125,N_7175);
and U7299 (N_7299,N_7089,N_7187);
nand U7300 (N_7300,N_7073,N_7087);
or U7301 (N_7301,N_7081,N_7016);
xnor U7302 (N_7302,N_7064,N_7018);
or U7303 (N_7303,N_7076,N_7106);
or U7304 (N_7304,N_7163,N_7113);
nor U7305 (N_7305,N_7009,N_7145);
xnor U7306 (N_7306,N_7043,N_7004);
or U7307 (N_7307,N_7174,N_7155);
nand U7308 (N_7308,N_7134,N_7047);
nand U7309 (N_7309,N_7001,N_7065);
or U7310 (N_7310,N_7125,N_7154);
xnor U7311 (N_7311,N_7184,N_7155);
nand U7312 (N_7312,N_7118,N_7113);
or U7313 (N_7313,N_7080,N_7177);
nor U7314 (N_7314,N_7075,N_7049);
xor U7315 (N_7315,N_7016,N_7155);
and U7316 (N_7316,N_7176,N_7101);
or U7317 (N_7317,N_7182,N_7122);
xor U7318 (N_7318,N_7096,N_7093);
nand U7319 (N_7319,N_7054,N_7067);
xnor U7320 (N_7320,N_7035,N_7104);
nor U7321 (N_7321,N_7040,N_7165);
nand U7322 (N_7322,N_7147,N_7109);
or U7323 (N_7323,N_7169,N_7008);
nand U7324 (N_7324,N_7177,N_7119);
nand U7325 (N_7325,N_7147,N_7087);
and U7326 (N_7326,N_7081,N_7070);
xnor U7327 (N_7327,N_7168,N_7116);
and U7328 (N_7328,N_7188,N_7038);
xor U7329 (N_7329,N_7176,N_7153);
nand U7330 (N_7330,N_7195,N_7105);
or U7331 (N_7331,N_7120,N_7159);
and U7332 (N_7332,N_7143,N_7059);
and U7333 (N_7333,N_7129,N_7150);
nor U7334 (N_7334,N_7107,N_7001);
and U7335 (N_7335,N_7017,N_7189);
nor U7336 (N_7336,N_7006,N_7186);
nor U7337 (N_7337,N_7191,N_7104);
and U7338 (N_7338,N_7062,N_7153);
xor U7339 (N_7339,N_7046,N_7035);
nand U7340 (N_7340,N_7059,N_7005);
and U7341 (N_7341,N_7179,N_7028);
or U7342 (N_7342,N_7193,N_7049);
xnor U7343 (N_7343,N_7162,N_7021);
and U7344 (N_7344,N_7135,N_7146);
or U7345 (N_7345,N_7023,N_7025);
nand U7346 (N_7346,N_7044,N_7004);
xor U7347 (N_7347,N_7188,N_7168);
and U7348 (N_7348,N_7011,N_7140);
or U7349 (N_7349,N_7171,N_7053);
nand U7350 (N_7350,N_7194,N_7057);
nor U7351 (N_7351,N_7137,N_7125);
nand U7352 (N_7352,N_7018,N_7006);
and U7353 (N_7353,N_7036,N_7086);
or U7354 (N_7354,N_7129,N_7122);
and U7355 (N_7355,N_7114,N_7110);
and U7356 (N_7356,N_7065,N_7165);
and U7357 (N_7357,N_7109,N_7091);
xnor U7358 (N_7358,N_7105,N_7028);
nand U7359 (N_7359,N_7113,N_7137);
xor U7360 (N_7360,N_7192,N_7193);
and U7361 (N_7361,N_7029,N_7128);
nand U7362 (N_7362,N_7067,N_7001);
xnor U7363 (N_7363,N_7003,N_7123);
or U7364 (N_7364,N_7107,N_7155);
nand U7365 (N_7365,N_7129,N_7141);
nand U7366 (N_7366,N_7141,N_7006);
nor U7367 (N_7367,N_7037,N_7088);
or U7368 (N_7368,N_7123,N_7160);
xnor U7369 (N_7369,N_7016,N_7102);
and U7370 (N_7370,N_7073,N_7027);
and U7371 (N_7371,N_7045,N_7052);
xor U7372 (N_7372,N_7075,N_7174);
nand U7373 (N_7373,N_7040,N_7155);
xor U7374 (N_7374,N_7098,N_7097);
or U7375 (N_7375,N_7002,N_7077);
and U7376 (N_7376,N_7151,N_7098);
or U7377 (N_7377,N_7161,N_7115);
nand U7378 (N_7378,N_7199,N_7052);
or U7379 (N_7379,N_7069,N_7094);
nand U7380 (N_7380,N_7102,N_7101);
nor U7381 (N_7381,N_7051,N_7086);
nand U7382 (N_7382,N_7195,N_7199);
xnor U7383 (N_7383,N_7070,N_7091);
nand U7384 (N_7384,N_7034,N_7036);
nand U7385 (N_7385,N_7153,N_7189);
xnor U7386 (N_7386,N_7140,N_7156);
nor U7387 (N_7387,N_7026,N_7142);
or U7388 (N_7388,N_7015,N_7028);
or U7389 (N_7389,N_7078,N_7156);
xor U7390 (N_7390,N_7074,N_7051);
nand U7391 (N_7391,N_7030,N_7189);
and U7392 (N_7392,N_7075,N_7138);
nand U7393 (N_7393,N_7140,N_7026);
and U7394 (N_7394,N_7048,N_7121);
or U7395 (N_7395,N_7174,N_7012);
nor U7396 (N_7396,N_7159,N_7184);
nand U7397 (N_7397,N_7127,N_7060);
xnor U7398 (N_7398,N_7130,N_7031);
nand U7399 (N_7399,N_7038,N_7158);
and U7400 (N_7400,N_7258,N_7273);
or U7401 (N_7401,N_7354,N_7341);
xor U7402 (N_7402,N_7272,N_7377);
nand U7403 (N_7403,N_7386,N_7374);
and U7404 (N_7404,N_7360,N_7389);
xor U7405 (N_7405,N_7245,N_7305);
and U7406 (N_7406,N_7234,N_7286);
nand U7407 (N_7407,N_7280,N_7214);
nand U7408 (N_7408,N_7224,N_7356);
and U7409 (N_7409,N_7366,N_7253);
or U7410 (N_7410,N_7205,N_7269);
nand U7411 (N_7411,N_7319,N_7327);
nand U7412 (N_7412,N_7352,N_7202);
nor U7413 (N_7413,N_7378,N_7304);
nand U7414 (N_7414,N_7333,N_7302);
or U7415 (N_7415,N_7266,N_7331);
and U7416 (N_7416,N_7287,N_7242);
nand U7417 (N_7417,N_7313,N_7271);
nand U7418 (N_7418,N_7220,N_7387);
nor U7419 (N_7419,N_7330,N_7209);
or U7420 (N_7420,N_7316,N_7328);
nor U7421 (N_7421,N_7268,N_7215);
or U7422 (N_7422,N_7345,N_7390);
nand U7423 (N_7423,N_7257,N_7281);
nor U7424 (N_7424,N_7226,N_7284);
nand U7425 (N_7425,N_7288,N_7325);
or U7426 (N_7426,N_7218,N_7381);
xnor U7427 (N_7427,N_7329,N_7376);
or U7428 (N_7428,N_7221,N_7332);
xor U7429 (N_7429,N_7346,N_7296);
xor U7430 (N_7430,N_7267,N_7339);
and U7431 (N_7431,N_7206,N_7203);
xor U7432 (N_7432,N_7223,N_7278);
xor U7433 (N_7433,N_7247,N_7303);
nand U7434 (N_7434,N_7357,N_7398);
and U7435 (N_7435,N_7320,N_7300);
and U7436 (N_7436,N_7384,N_7365);
or U7437 (N_7437,N_7229,N_7363);
or U7438 (N_7438,N_7235,N_7350);
nor U7439 (N_7439,N_7219,N_7348);
nor U7440 (N_7440,N_7236,N_7369);
or U7441 (N_7441,N_7317,N_7222);
nand U7442 (N_7442,N_7298,N_7250);
nand U7443 (N_7443,N_7394,N_7241);
nand U7444 (N_7444,N_7263,N_7260);
nand U7445 (N_7445,N_7204,N_7309);
xnor U7446 (N_7446,N_7393,N_7334);
or U7447 (N_7447,N_7255,N_7395);
nor U7448 (N_7448,N_7212,N_7290);
xor U7449 (N_7449,N_7385,N_7252);
nor U7450 (N_7450,N_7326,N_7311);
xnor U7451 (N_7451,N_7307,N_7349);
and U7452 (N_7452,N_7340,N_7210);
and U7453 (N_7453,N_7392,N_7337);
nand U7454 (N_7454,N_7367,N_7279);
nor U7455 (N_7455,N_7399,N_7379);
nand U7456 (N_7456,N_7383,N_7373);
nand U7457 (N_7457,N_7238,N_7239);
nand U7458 (N_7458,N_7347,N_7342);
nor U7459 (N_7459,N_7361,N_7291);
or U7460 (N_7460,N_7324,N_7217);
or U7461 (N_7461,N_7225,N_7201);
xnor U7462 (N_7462,N_7382,N_7227);
xor U7463 (N_7463,N_7276,N_7297);
nand U7464 (N_7464,N_7270,N_7256);
nand U7465 (N_7465,N_7230,N_7254);
xnor U7466 (N_7466,N_7207,N_7293);
xnor U7467 (N_7467,N_7295,N_7338);
nor U7468 (N_7468,N_7240,N_7244);
or U7469 (N_7469,N_7380,N_7371);
and U7470 (N_7470,N_7248,N_7310);
nand U7471 (N_7471,N_7322,N_7368);
and U7472 (N_7472,N_7355,N_7233);
xor U7473 (N_7473,N_7249,N_7312);
or U7474 (N_7474,N_7274,N_7283);
and U7475 (N_7475,N_7216,N_7251);
nand U7476 (N_7476,N_7397,N_7344);
xor U7477 (N_7477,N_7246,N_7264);
and U7478 (N_7478,N_7375,N_7299);
nand U7479 (N_7479,N_7358,N_7237);
and U7480 (N_7480,N_7208,N_7275);
nand U7481 (N_7481,N_7335,N_7343);
nand U7482 (N_7482,N_7213,N_7314);
nand U7483 (N_7483,N_7372,N_7370);
nand U7484 (N_7484,N_7211,N_7323);
and U7485 (N_7485,N_7289,N_7294);
nand U7486 (N_7486,N_7364,N_7228);
nand U7487 (N_7487,N_7318,N_7353);
and U7488 (N_7488,N_7277,N_7265);
xor U7489 (N_7489,N_7243,N_7259);
and U7490 (N_7490,N_7396,N_7262);
nand U7491 (N_7491,N_7362,N_7351);
or U7492 (N_7492,N_7308,N_7306);
and U7493 (N_7493,N_7321,N_7391);
and U7494 (N_7494,N_7200,N_7285);
xnor U7495 (N_7495,N_7282,N_7388);
xor U7496 (N_7496,N_7261,N_7231);
nand U7497 (N_7497,N_7292,N_7359);
nand U7498 (N_7498,N_7301,N_7336);
or U7499 (N_7499,N_7315,N_7232);
nor U7500 (N_7500,N_7208,N_7360);
nand U7501 (N_7501,N_7317,N_7293);
or U7502 (N_7502,N_7394,N_7239);
nand U7503 (N_7503,N_7334,N_7224);
xor U7504 (N_7504,N_7270,N_7375);
and U7505 (N_7505,N_7377,N_7352);
and U7506 (N_7506,N_7358,N_7377);
xor U7507 (N_7507,N_7346,N_7267);
xor U7508 (N_7508,N_7270,N_7268);
nor U7509 (N_7509,N_7322,N_7394);
xor U7510 (N_7510,N_7345,N_7327);
nor U7511 (N_7511,N_7390,N_7272);
and U7512 (N_7512,N_7217,N_7373);
nor U7513 (N_7513,N_7300,N_7330);
nand U7514 (N_7514,N_7383,N_7231);
and U7515 (N_7515,N_7203,N_7369);
or U7516 (N_7516,N_7316,N_7232);
or U7517 (N_7517,N_7242,N_7221);
xor U7518 (N_7518,N_7264,N_7329);
nor U7519 (N_7519,N_7225,N_7266);
or U7520 (N_7520,N_7280,N_7282);
or U7521 (N_7521,N_7301,N_7362);
or U7522 (N_7522,N_7260,N_7317);
and U7523 (N_7523,N_7266,N_7385);
nand U7524 (N_7524,N_7274,N_7333);
nand U7525 (N_7525,N_7239,N_7261);
xor U7526 (N_7526,N_7340,N_7391);
nand U7527 (N_7527,N_7303,N_7257);
nand U7528 (N_7528,N_7382,N_7225);
xor U7529 (N_7529,N_7285,N_7367);
nand U7530 (N_7530,N_7346,N_7297);
and U7531 (N_7531,N_7223,N_7222);
nand U7532 (N_7532,N_7395,N_7215);
xor U7533 (N_7533,N_7279,N_7305);
xor U7534 (N_7534,N_7243,N_7361);
and U7535 (N_7535,N_7280,N_7242);
xnor U7536 (N_7536,N_7391,N_7342);
nand U7537 (N_7537,N_7320,N_7305);
and U7538 (N_7538,N_7316,N_7247);
or U7539 (N_7539,N_7224,N_7365);
nor U7540 (N_7540,N_7223,N_7296);
nor U7541 (N_7541,N_7244,N_7303);
xnor U7542 (N_7542,N_7327,N_7322);
or U7543 (N_7543,N_7313,N_7296);
nor U7544 (N_7544,N_7320,N_7286);
or U7545 (N_7545,N_7366,N_7316);
nor U7546 (N_7546,N_7292,N_7396);
and U7547 (N_7547,N_7210,N_7317);
nor U7548 (N_7548,N_7292,N_7270);
or U7549 (N_7549,N_7294,N_7324);
or U7550 (N_7550,N_7317,N_7307);
xnor U7551 (N_7551,N_7304,N_7263);
nor U7552 (N_7552,N_7226,N_7277);
and U7553 (N_7553,N_7309,N_7280);
and U7554 (N_7554,N_7367,N_7287);
nand U7555 (N_7555,N_7372,N_7330);
xor U7556 (N_7556,N_7303,N_7398);
nor U7557 (N_7557,N_7327,N_7381);
nand U7558 (N_7558,N_7323,N_7256);
or U7559 (N_7559,N_7321,N_7263);
nand U7560 (N_7560,N_7273,N_7212);
and U7561 (N_7561,N_7294,N_7233);
xnor U7562 (N_7562,N_7338,N_7209);
nor U7563 (N_7563,N_7299,N_7257);
xnor U7564 (N_7564,N_7284,N_7315);
or U7565 (N_7565,N_7228,N_7239);
or U7566 (N_7566,N_7208,N_7398);
nand U7567 (N_7567,N_7264,N_7348);
or U7568 (N_7568,N_7329,N_7323);
nand U7569 (N_7569,N_7316,N_7341);
nor U7570 (N_7570,N_7347,N_7260);
or U7571 (N_7571,N_7354,N_7302);
xor U7572 (N_7572,N_7281,N_7245);
or U7573 (N_7573,N_7386,N_7274);
and U7574 (N_7574,N_7393,N_7213);
nand U7575 (N_7575,N_7358,N_7372);
nand U7576 (N_7576,N_7237,N_7282);
nand U7577 (N_7577,N_7332,N_7273);
xnor U7578 (N_7578,N_7324,N_7341);
nor U7579 (N_7579,N_7227,N_7211);
or U7580 (N_7580,N_7275,N_7271);
and U7581 (N_7581,N_7375,N_7305);
nor U7582 (N_7582,N_7200,N_7338);
nand U7583 (N_7583,N_7348,N_7284);
and U7584 (N_7584,N_7220,N_7348);
xor U7585 (N_7585,N_7205,N_7385);
and U7586 (N_7586,N_7354,N_7266);
xor U7587 (N_7587,N_7230,N_7233);
and U7588 (N_7588,N_7242,N_7258);
nand U7589 (N_7589,N_7200,N_7264);
or U7590 (N_7590,N_7208,N_7355);
nand U7591 (N_7591,N_7286,N_7200);
xor U7592 (N_7592,N_7246,N_7292);
xor U7593 (N_7593,N_7376,N_7312);
nand U7594 (N_7594,N_7241,N_7357);
xor U7595 (N_7595,N_7286,N_7248);
xnor U7596 (N_7596,N_7355,N_7302);
or U7597 (N_7597,N_7293,N_7339);
or U7598 (N_7598,N_7212,N_7395);
nor U7599 (N_7599,N_7265,N_7335);
nand U7600 (N_7600,N_7409,N_7404);
nor U7601 (N_7601,N_7583,N_7589);
nor U7602 (N_7602,N_7521,N_7435);
nand U7603 (N_7603,N_7503,N_7405);
nor U7604 (N_7604,N_7483,N_7509);
nand U7605 (N_7605,N_7574,N_7438);
xor U7606 (N_7606,N_7570,N_7577);
or U7607 (N_7607,N_7587,N_7530);
or U7608 (N_7608,N_7416,N_7507);
nor U7609 (N_7609,N_7452,N_7519);
nor U7610 (N_7610,N_7440,N_7415);
and U7611 (N_7611,N_7550,N_7543);
xnor U7612 (N_7612,N_7517,N_7460);
or U7613 (N_7613,N_7418,N_7508);
xor U7614 (N_7614,N_7564,N_7485);
or U7615 (N_7615,N_7513,N_7496);
or U7616 (N_7616,N_7477,N_7497);
nand U7617 (N_7617,N_7518,N_7437);
nor U7618 (N_7618,N_7400,N_7420);
and U7619 (N_7619,N_7585,N_7489);
nor U7620 (N_7620,N_7599,N_7545);
and U7621 (N_7621,N_7598,N_7449);
nand U7622 (N_7622,N_7554,N_7504);
nor U7623 (N_7623,N_7582,N_7520);
nor U7624 (N_7624,N_7514,N_7568);
nor U7625 (N_7625,N_7590,N_7484);
or U7626 (N_7626,N_7524,N_7469);
and U7627 (N_7627,N_7542,N_7558);
nor U7628 (N_7628,N_7562,N_7546);
or U7629 (N_7629,N_7412,N_7492);
nor U7630 (N_7630,N_7549,N_7476);
and U7631 (N_7631,N_7436,N_7414);
xnor U7632 (N_7632,N_7426,N_7559);
xor U7633 (N_7633,N_7433,N_7527);
nand U7634 (N_7634,N_7486,N_7548);
nor U7635 (N_7635,N_7547,N_7472);
xor U7636 (N_7636,N_7540,N_7493);
nor U7637 (N_7637,N_7471,N_7499);
and U7638 (N_7638,N_7417,N_7466);
or U7639 (N_7639,N_7584,N_7528);
nand U7640 (N_7640,N_7555,N_7579);
nor U7641 (N_7641,N_7478,N_7432);
nand U7642 (N_7642,N_7408,N_7423);
nor U7643 (N_7643,N_7595,N_7488);
nor U7644 (N_7644,N_7557,N_7475);
nand U7645 (N_7645,N_7410,N_7479);
and U7646 (N_7646,N_7441,N_7516);
nand U7647 (N_7647,N_7451,N_7586);
xnor U7648 (N_7648,N_7462,N_7551);
xnor U7649 (N_7649,N_7526,N_7544);
xor U7650 (N_7650,N_7459,N_7463);
nand U7651 (N_7651,N_7500,N_7455);
or U7652 (N_7652,N_7443,N_7580);
nand U7653 (N_7653,N_7474,N_7538);
nand U7654 (N_7654,N_7402,N_7422);
nor U7655 (N_7655,N_7413,N_7439);
nor U7656 (N_7656,N_7591,N_7470);
and U7657 (N_7657,N_7597,N_7575);
or U7658 (N_7658,N_7446,N_7461);
nand U7659 (N_7659,N_7487,N_7531);
xnor U7660 (N_7660,N_7468,N_7578);
xnor U7661 (N_7661,N_7573,N_7525);
and U7662 (N_7662,N_7532,N_7406);
nand U7663 (N_7663,N_7522,N_7529);
nor U7664 (N_7664,N_7510,N_7491);
and U7665 (N_7665,N_7553,N_7450);
xnor U7666 (N_7666,N_7481,N_7502);
and U7667 (N_7667,N_7565,N_7447);
xor U7668 (N_7668,N_7403,N_7566);
xnor U7669 (N_7669,N_7572,N_7465);
or U7670 (N_7670,N_7464,N_7560);
nand U7671 (N_7671,N_7596,N_7511);
xnor U7672 (N_7672,N_7505,N_7430);
nor U7673 (N_7673,N_7458,N_7567);
nor U7674 (N_7674,N_7494,N_7424);
or U7675 (N_7675,N_7482,N_7429);
or U7676 (N_7676,N_7563,N_7495);
and U7677 (N_7677,N_7523,N_7541);
and U7678 (N_7678,N_7581,N_7490);
xnor U7679 (N_7679,N_7407,N_7556);
and U7680 (N_7680,N_7534,N_7576);
or U7681 (N_7681,N_7498,N_7533);
nand U7682 (N_7682,N_7431,N_7593);
and U7683 (N_7683,N_7536,N_7448);
nor U7684 (N_7684,N_7453,N_7539);
nor U7685 (N_7685,N_7480,N_7442);
nor U7686 (N_7686,N_7515,N_7457);
nor U7687 (N_7687,N_7537,N_7425);
or U7688 (N_7688,N_7552,N_7506);
or U7689 (N_7689,N_7401,N_7419);
and U7690 (N_7690,N_7512,N_7473);
nand U7691 (N_7691,N_7428,N_7571);
nor U7692 (N_7692,N_7561,N_7592);
and U7693 (N_7693,N_7411,N_7467);
nand U7694 (N_7694,N_7421,N_7454);
xnor U7695 (N_7695,N_7445,N_7427);
nor U7696 (N_7696,N_7569,N_7501);
xnor U7697 (N_7697,N_7594,N_7456);
and U7698 (N_7698,N_7444,N_7535);
and U7699 (N_7699,N_7434,N_7588);
xor U7700 (N_7700,N_7543,N_7428);
nand U7701 (N_7701,N_7505,N_7482);
nand U7702 (N_7702,N_7508,N_7557);
or U7703 (N_7703,N_7496,N_7523);
xnor U7704 (N_7704,N_7482,N_7493);
nand U7705 (N_7705,N_7568,N_7441);
and U7706 (N_7706,N_7528,N_7579);
xnor U7707 (N_7707,N_7572,N_7495);
nand U7708 (N_7708,N_7594,N_7517);
or U7709 (N_7709,N_7494,N_7522);
nand U7710 (N_7710,N_7589,N_7471);
nor U7711 (N_7711,N_7422,N_7575);
and U7712 (N_7712,N_7529,N_7506);
or U7713 (N_7713,N_7541,N_7511);
xor U7714 (N_7714,N_7441,N_7519);
nor U7715 (N_7715,N_7591,N_7499);
nand U7716 (N_7716,N_7447,N_7550);
nor U7717 (N_7717,N_7583,N_7573);
and U7718 (N_7718,N_7572,N_7496);
nor U7719 (N_7719,N_7490,N_7510);
nor U7720 (N_7720,N_7578,N_7532);
or U7721 (N_7721,N_7481,N_7519);
or U7722 (N_7722,N_7469,N_7593);
nand U7723 (N_7723,N_7472,N_7464);
xor U7724 (N_7724,N_7476,N_7592);
and U7725 (N_7725,N_7541,N_7439);
xor U7726 (N_7726,N_7497,N_7462);
xor U7727 (N_7727,N_7575,N_7428);
or U7728 (N_7728,N_7540,N_7448);
nand U7729 (N_7729,N_7579,N_7529);
and U7730 (N_7730,N_7495,N_7467);
xor U7731 (N_7731,N_7460,N_7457);
nor U7732 (N_7732,N_7591,N_7589);
nor U7733 (N_7733,N_7505,N_7477);
nor U7734 (N_7734,N_7569,N_7440);
nand U7735 (N_7735,N_7582,N_7490);
xnor U7736 (N_7736,N_7538,N_7528);
nand U7737 (N_7737,N_7599,N_7461);
nand U7738 (N_7738,N_7559,N_7473);
nor U7739 (N_7739,N_7474,N_7565);
xor U7740 (N_7740,N_7519,N_7520);
nor U7741 (N_7741,N_7513,N_7526);
xnor U7742 (N_7742,N_7407,N_7533);
xnor U7743 (N_7743,N_7497,N_7421);
nor U7744 (N_7744,N_7585,N_7598);
xnor U7745 (N_7745,N_7476,N_7432);
nand U7746 (N_7746,N_7552,N_7559);
nand U7747 (N_7747,N_7567,N_7526);
nand U7748 (N_7748,N_7514,N_7482);
nand U7749 (N_7749,N_7590,N_7468);
or U7750 (N_7750,N_7434,N_7492);
xor U7751 (N_7751,N_7533,N_7494);
nand U7752 (N_7752,N_7455,N_7507);
nor U7753 (N_7753,N_7597,N_7421);
and U7754 (N_7754,N_7573,N_7432);
nor U7755 (N_7755,N_7404,N_7511);
and U7756 (N_7756,N_7412,N_7505);
or U7757 (N_7757,N_7482,N_7556);
nand U7758 (N_7758,N_7405,N_7504);
nor U7759 (N_7759,N_7557,N_7583);
xnor U7760 (N_7760,N_7586,N_7587);
or U7761 (N_7761,N_7511,N_7583);
nand U7762 (N_7762,N_7585,N_7531);
or U7763 (N_7763,N_7581,N_7598);
nor U7764 (N_7764,N_7430,N_7408);
and U7765 (N_7765,N_7456,N_7552);
and U7766 (N_7766,N_7586,N_7561);
and U7767 (N_7767,N_7489,N_7499);
and U7768 (N_7768,N_7538,N_7420);
nand U7769 (N_7769,N_7578,N_7459);
nor U7770 (N_7770,N_7596,N_7487);
and U7771 (N_7771,N_7557,N_7556);
xnor U7772 (N_7772,N_7590,N_7505);
xnor U7773 (N_7773,N_7474,N_7594);
and U7774 (N_7774,N_7566,N_7589);
and U7775 (N_7775,N_7441,N_7533);
xor U7776 (N_7776,N_7506,N_7407);
and U7777 (N_7777,N_7444,N_7401);
nand U7778 (N_7778,N_7551,N_7471);
or U7779 (N_7779,N_7487,N_7567);
nand U7780 (N_7780,N_7574,N_7545);
and U7781 (N_7781,N_7402,N_7462);
nand U7782 (N_7782,N_7434,N_7535);
nor U7783 (N_7783,N_7504,N_7424);
xor U7784 (N_7784,N_7487,N_7574);
or U7785 (N_7785,N_7408,N_7445);
or U7786 (N_7786,N_7528,N_7557);
and U7787 (N_7787,N_7537,N_7458);
nor U7788 (N_7788,N_7590,N_7425);
xnor U7789 (N_7789,N_7412,N_7460);
xor U7790 (N_7790,N_7450,N_7581);
or U7791 (N_7791,N_7575,N_7524);
nand U7792 (N_7792,N_7403,N_7441);
or U7793 (N_7793,N_7426,N_7429);
xnor U7794 (N_7794,N_7463,N_7477);
or U7795 (N_7795,N_7573,N_7426);
xnor U7796 (N_7796,N_7512,N_7510);
and U7797 (N_7797,N_7436,N_7551);
or U7798 (N_7798,N_7451,N_7488);
nor U7799 (N_7799,N_7436,N_7475);
nand U7800 (N_7800,N_7777,N_7627);
and U7801 (N_7801,N_7671,N_7719);
and U7802 (N_7802,N_7607,N_7672);
and U7803 (N_7803,N_7731,N_7623);
xnor U7804 (N_7804,N_7609,N_7765);
or U7805 (N_7805,N_7668,N_7673);
nand U7806 (N_7806,N_7649,N_7628);
nor U7807 (N_7807,N_7794,N_7782);
nand U7808 (N_7808,N_7652,N_7648);
nand U7809 (N_7809,N_7694,N_7662);
nor U7810 (N_7810,N_7769,N_7746);
and U7811 (N_7811,N_7644,N_7634);
and U7812 (N_7812,N_7772,N_7733);
and U7813 (N_7813,N_7748,N_7760);
and U7814 (N_7814,N_7755,N_7636);
nor U7815 (N_7815,N_7653,N_7656);
nand U7816 (N_7816,N_7764,N_7758);
nor U7817 (N_7817,N_7783,N_7768);
and U7818 (N_7818,N_7657,N_7693);
nor U7819 (N_7819,N_7602,N_7788);
and U7820 (N_7820,N_7659,N_7647);
nor U7821 (N_7821,N_7727,N_7745);
and U7822 (N_7822,N_7626,N_7631);
nor U7823 (N_7823,N_7744,N_7650);
nor U7824 (N_7824,N_7669,N_7775);
nor U7825 (N_7825,N_7606,N_7698);
and U7826 (N_7826,N_7722,N_7785);
and U7827 (N_7827,N_7739,N_7793);
and U7828 (N_7828,N_7608,N_7786);
or U7829 (N_7829,N_7685,N_7618);
and U7830 (N_7830,N_7735,N_7633);
and U7831 (N_7831,N_7701,N_7614);
nor U7832 (N_7832,N_7663,N_7730);
nand U7833 (N_7833,N_7741,N_7717);
and U7834 (N_7834,N_7686,N_7610);
or U7835 (N_7835,N_7665,N_7705);
xor U7836 (N_7836,N_7674,N_7661);
nand U7837 (N_7837,N_7711,N_7639);
or U7838 (N_7838,N_7664,N_7754);
nor U7839 (N_7839,N_7729,N_7790);
or U7840 (N_7840,N_7638,N_7750);
or U7841 (N_7841,N_7751,N_7767);
or U7842 (N_7842,N_7688,N_7712);
nor U7843 (N_7843,N_7797,N_7718);
nand U7844 (N_7844,N_7704,N_7703);
and U7845 (N_7845,N_7655,N_7660);
or U7846 (N_7846,N_7742,N_7714);
nor U7847 (N_7847,N_7779,N_7678);
or U7848 (N_7848,N_7734,N_7799);
and U7849 (N_7849,N_7696,N_7620);
or U7850 (N_7850,N_7612,N_7747);
nor U7851 (N_7851,N_7773,N_7738);
or U7852 (N_7852,N_7736,N_7687);
xor U7853 (N_7853,N_7654,N_7667);
nor U7854 (N_7854,N_7713,N_7737);
xor U7855 (N_7855,N_7680,N_7640);
xor U7856 (N_7856,N_7684,N_7621);
nand U7857 (N_7857,N_7726,N_7642);
and U7858 (N_7858,N_7635,N_7616);
xnor U7859 (N_7859,N_7641,N_7749);
xor U7860 (N_7860,N_7702,N_7677);
or U7861 (N_7861,N_7622,N_7781);
xor U7862 (N_7862,N_7697,N_7708);
xnor U7863 (N_7863,N_7700,N_7699);
nand U7864 (N_7864,N_7690,N_7695);
and U7865 (N_7865,N_7796,N_7604);
or U7866 (N_7866,N_7691,N_7784);
nor U7867 (N_7867,N_7721,N_7689);
nand U7868 (N_7868,N_7629,N_7753);
nor U7869 (N_7869,N_7715,N_7752);
or U7870 (N_7870,N_7724,N_7603);
xnor U7871 (N_7871,N_7666,N_7798);
or U7872 (N_7872,N_7676,N_7658);
xor U7873 (N_7873,N_7732,N_7716);
nand U7874 (N_7874,N_7759,N_7625);
or U7875 (N_7875,N_7770,N_7619);
xnor U7876 (N_7876,N_7624,N_7709);
and U7877 (N_7877,N_7675,N_7723);
nor U7878 (N_7878,N_7651,N_7681);
and U7879 (N_7879,N_7761,N_7789);
xnor U7880 (N_7880,N_7632,N_7740);
and U7881 (N_7881,N_7646,N_7787);
nand U7882 (N_7882,N_7728,N_7743);
and U7883 (N_7883,N_7778,N_7601);
nor U7884 (N_7884,N_7615,N_7780);
and U7885 (N_7885,N_7643,N_7766);
nor U7886 (N_7886,N_7683,N_7771);
or U7887 (N_7887,N_7630,N_7757);
nor U7888 (N_7888,N_7605,N_7611);
or U7889 (N_7889,N_7613,N_7791);
nand U7890 (N_7890,N_7795,N_7774);
or U7891 (N_7891,N_7600,N_7725);
and U7892 (N_7892,N_7645,N_7710);
xnor U7893 (N_7893,N_7776,N_7692);
xnor U7894 (N_7894,N_7707,N_7720);
nor U7895 (N_7895,N_7670,N_7617);
xor U7896 (N_7896,N_7682,N_7637);
or U7897 (N_7897,N_7792,N_7762);
or U7898 (N_7898,N_7679,N_7763);
nor U7899 (N_7899,N_7756,N_7706);
xnor U7900 (N_7900,N_7629,N_7602);
xor U7901 (N_7901,N_7624,N_7724);
xor U7902 (N_7902,N_7690,N_7777);
nor U7903 (N_7903,N_7707,N_7714);
nor U7904 (N_7904,N_7769,N_7788);
and U7905 (N_7905,N_7735,N_7631);
nor U7906 (N_7906,N_7655,N_7798);
xor U7907 (N_7907,N_7738,N_7707);
xnor U7908 (N_7908,N_7669,N_7609);
nor U7909 (N_7909,N_7626,N_7654);
nand U7910 (N_7910,N_7787,N_7675);
xor U7911 (N_7911,N_7739,N_7715);
nand U7912 (N_7912,N_7633,N_7649);
or U7913 (N_7913,N_7656,N_7604);
nor U7914 (N_7914,N_7704,N_7673);
or U7915 (N_7915,N_7673,N_7785);
and U7916 (N_7916,N_7776,N_7786);
nor U7917 (N_7917,N_7654,N_7738);
nand U7918 (N_7918,N_7743,N_7730);
nand U7919 (N_7919,N_7760,N_7787);
and U7920 (N_7920,N_7743,N_7721);
and U7921 (N_7921,N_7721,N_7724);
xnor U7922 (N_7922,N_7660,N_7760);
nor U7923 (N_7923,N_7796,N_7799);
xnor U7924 (N_7924,N_7611,N_7706);
nand U7925 (N_7925,N_7735,N_7626);
nor U7926 (N_7926,N_7789,N_7720);
xnor U7927 (N_7927,N_7610,N_7722);
xnor U7928 (N_7928,N_7655,N_7736);
and U7929 (N_7929,N_7699,N_7604);
nor U7930 (N_7930,N_7778,N_7679);
xnor U7931 (N_7931,N_7671,N_7656);
nor U7932 (N_7932,N_7666,N_7691);
and U7933 (N_7933,N_7668,N_7782);
nor U7934 (N_7934,N_7723,N_7787);
and U7935 (N_7935,N_7739,N_7782);
nand U7936 (N_7936,N_7630,N_7615);
nand U7937 (N_7937,N_7701,N_7691);
and U7938 (N_7938,N_7731,N_7791);
xnor U7939 (N_7939,N_7784,N_7663);
nor U7940 (N_7940,N_7677,N_7637);
nand U7941 (N_7941,N_7664,N_7715);
nand U7942 (N_7942,N_7630,N_7609);
nand U7943 (N_7943,N_7676,N_7645);
nand U7944 (N_7944,N_7639,N_7736);
xor U7945 (N_7945,N_7616,N_7623);
and U7946 (N_7946,N_7765,N_7688);
and U7947 (N_7947,N_7774,N_7681);
xor U7948 (N_7948,N_7751,N_7762);
nand U7949 (N_7949,N_7678,N_7783);
nand U7950 (N_7950,N_7622,N_7705);
xnor U7951 (N_7951,N_7653,N_7632);
nand U7952 (N_7952,N_7790,N_7695);
nor U7953 (N_7953,N_7709,N_7716);
or U7954 (N_7954,N_7749,N_7680);
nand U7955 (N_7955,N_7731,N_7679);
nor U7956 (N_7956,N_7725,N_7779);
nand U7957 (N_7957,N_7619,N_7794);
or U7958 (N_7958,N_7687,N_7733);
xor U7959 (N_7959,N_7788,N_7635);
xor U7960 (N_7960,N_7603,N_7752);
and U7961 (N_7961,N_7667,N_7642);
xor U7962 (N_7962,N_7748,N_7794);
and U7963 (N_7963,N_7612,N_7693);
and U7964 (N_7964,N_7677,N_7762);
and U7965 (N_7965,N_7630,N_7633);
and U7966 (N_7966,N_7622,N_7770);
nand U7967 (N_7967,N_7743,N_7733);
nand U7968 (N_7968,N_7750,N_7698);
and U7969 (N_7969,N_7787,N_7680);
and U7970 (N_7970,N_7635,N_7760);
xnor U7971 (N_7971,N_7629,N_7784);
xor U7972 (N_7972,N_7703,N_7689);
and U7973 (N_7973,N_7786,N_7679);
or U7974 (N_7974,N_7624,N_7641);
nand U7975 (N_7975,N_7608,N_7643);
xor U7976 (N_7976,N_7688,N_7785);
nand U7977 (N_7977,N_7668,N_7655);
and U7978 (N_7978,N_7699,N_7697);
nand U7979 (N_7979,N_7760,N_7630);
nand U7980 (N_7980,N_7621,N_7655);
and U7981 (N_7981,N_7744,N_7661);
nor U7982 (N_7982,N_7791,N_7752);
or U7983 (N_7983,N_7624,N_7797);
nor U7984 (N_7984,N_7606,N_7640);
and U7985 (N_7985,N_7686,N_7626);
and U7986 (N_7986,N_7739,N_7662);
and U7987 (N_7987,N_7608,N_7686);
nand U7988 (N_7988,N_7787,N_7713);
nand U7989 (N_7989,N_7619,N_7640);
and U7990 (N_7990,N_7775,N_7684);
nand U7991 (N_7991,N_7648,N_7698);
xor U7992 (N_7992,N_7669,N_7618);
or U7993 (N_7993,N_7764,N_7778);
xnor U7994 (N_7994,N_7745,N_7611);
nand U7995 (N_7995,N_7756,N_7641);
xnor U7996 (N_7996,N_7703,N_7786);
nand U7997 (N_7997,N_7713,N_7609);
or U7998 (N_7998,N_7649,N_7733);
xor U7999 (N_7999,N_7776,N_7616);
and U8000 (N_8000,N_7909,N_7871);
nor U8001 (N_8001,N_7885,N_7968);
or U8002 (N_8002,N_7981,N_7878);
nor U8003 (N_8003,N_7858,N_7944);
or U8004 (N_8004,N_7856,N_7945);
nor U8005 (N_8005,N_7894,N_7836);
nand U8006 (N_8006,N_7838,N_7879);
and U8007 (N_8007,N_7905,N_7870);
or U8008 (N_8008,N_7946,N_7817);
xnor U8009 (N_8009,N_7962,N_7986);
nor U8010 (N_8010,N_7803,N_7854);
xnor U8011 (N_8011,N_7896,N_7855);
and U8012 (N_8012,N_7847,N_7957);
nor U8013 (N_8013,N_7943,N_7900);
and U8014 (N_8014,N_7910,N_7874);
or U8015 (N_8015,N_7851,N_7906);
nor U8016 (N_8016,N_7974,N_7973);
nor U8017 (N_8017,N_7930,N_7891);
nand U8018 (N_8018,N_7996,N_7800);
and U8019 (N_8019,N_7915,N_7970);
nor U8020 (N_8020,N_7809,N_7921);
or U8021 (N_8021,N_7967,N_7966);
nor U8022 (N_8022,N_7977,N_7883);
and U8023 (N_8023,N_7826,N_7865);
nor U8024 (N_8024,N_7824,N_7994);
and U8025 (N_8025,N_7857,N_7927);
and U8026 (N_8026,N_7807,N_7842);
nor U8027 (N_8027,N_7805,N_7984);
xnor U8028 (N_8028,N_7983,N_7848);
xor U8029 (N_8029,N_7814,N_7908);
xnor U8030 (N_8030,N_7890,N_7822);
nor U8031 (N_8031,N_7999,N_7845);
nand U8032 (N_8032,N_7956,N_7887);
nor U8033 (N_8033,N_7825,N_7960);
nor U8034 (N_8034,N_7922,N_7835);
nand U8035 (N_8035,N_7931,N_7837);
or U8036 (N_8036,N_7976,N_7849);
xor U8037 (N_8037,N_7911,N_7925);
xnor U8038 (N_8038,N_7989,N_7802);
xor U8039 (N_8039,N_7827,N_7889);
nor U8040 (N_8040,N_7859,N_7954);
nand U8041 (N_8041,N_7917,N_7852);
nand U8042 (N_8042,N_7939,N_7808);
or U8043 (N_8043,N_7951,N_7846);
and U8044 (N_8044,N_7961,N_7913);
xor U8045 (N_8045,N_7868,N_7903);
or U8046 (N_8046,N_7963,N_7926);
nor U8047 (N_8047,N_7923,N_7801);
and U8048 (N_8048,N_7950,N_7810);
xor U8049 (N_8049,N_7937,N_7928);
nor U8050 (N_8050,N_7830,N_7948);
xor U8051 (N_8051,N_7895,N_7947);
and U8052 (N_8052,N_7843,N_7916);
xnor U8053 (N_8053,N_7952,N_7893);
or U8054 (N_8054,N_7959,N_7853);
xnor U8055 (N_8055,N_7812,N_7936);
and U8056 (N_8056,N_7990,N_7932);
nand U8057 (N_8057,N_7933,N_7978);
nor U8058 (N_8058,N_7877,N_7819);
xor U8059 (N_8059,N_7969,N_7949);
or U8060 (N_8060,N_7840,N_7876);
or U8061 (N_8061,N_7940,N_7832);
nand U8062 (N_8062,N_7864,N_7875);
and U8063 (N_8063,N_7839,N_7964);
nor U8064 (N_8064,N_7834,N_7899);
nand U8065 (N_8065,N_7831,N_7958);
nor U8066 (N_8066,N_7892,N_7955);
or U8067 (N_8067,N_7924,N_7881);
nor U8068 (N_8068,N_7841,N_7844);
nand U8069 (N_8069,N_7888,N_7993);
xor U8070 (N_8070,N_7897,N_7995);
nand U8071 (N_8071,N_7863,N_7998);
or U8072 (N_8072,N_7965,N_7997);
xnor U8073 (N_8073,N_7882,N_7971);
nor U8074 (N_8074,N_7804,N_7980);
nand U8075 (N_8075,N_7828,N_7866);
nand U8076 (N_8076,N_7907,N_7918);
and U8077 (N_8077,N_7813,N_7873);
or U8078 (N_8078,N_7942,N_7823);
nand U8079 (N_8079,N_7901,N_7985);
xnor U8080 (N_8080,N_7982,N_7867);
nand U8081 (N_8081,N_7816,N_7860);
or U8082 (N_8082,N_7934,N_7912);
or U8083 (N_8083,N_7861,N_7938);
and U8084 (N_8084,N_7902,N_7818);
or U8085 (N_8085,N_7806,N_7988);
and U8086 (N_8086,N_7975,N_7920);
and U8087 (N_8087,N_7898,N_7991);
and U8088 (N_8088,N_7919,N_7884);
or U8089 (N_8089,N_7821,N_7904);
nor U8090 (N_8090,N_7880,N_7869);
nand U8091 (N_8091,N_7929,N_7829);
or U8092 (N_8092,N_7815,N_7811);
or U8093 (N_8093,N_7914,N_7953);
nand U8094 (N_8094,N_7862,N_7979);
nor U8095 (N_8095,N_7987,N_7833);
nor U8096 (N_8096,N_7850,N_7820);
or U8097 (N_8097,N_7872,N_7972);
or U8098 (N_8098,N_7886,N_7941);
nand U8099 (N_8099,N_7992,N_7935);
and U8100 (N_8100,N_7963,N_7886);
nand U8101 (N_8101,N_7908,N_7955);
or U8102 (N_8102,N_7927,N_7972);
or U8103 (N_8103,N_7872,N_7922);
or U8104 (N_8104,N_7959,N_7914);
and U8105 (N_8105,N_7952,N_7902);
or U8106 (N_8106,N_7978,N_7974);
nor U8107 (N_8107,N_7809,N_7834);
xnor U8108 (N_8108,N_7908,N_7949);
and U8109 (N_8109,N_7863,N_7854);
and U8110 (N_8110,N_7947,N_7863);
and U8111 (N_8111,N_7875,N_7869);
xnor U8112 (N_8112,N_7846,N_7965);
xnor U8113 (N_8113,N_7861,N_7982);
xnor U8114 (N_8114,N_7811,N_7870);
or U8115 (N_8115,N_7856,N_7828);
nor U8116 (N_8116,N_7921,N_7810);
xor U8117 (N_8117,N_7894,N_7818);
or U8118 (N_8118,N_7884,N_7945);
or U8119 (N_8119,N_7961,N_7805);
or U8120 (N_8120,N_7941,N_7983);
xnor U8121 (N_8121,N_7893,N_7825);
nor U8122 (N_8122,N_7866,N_7820);
nor U8123 (N_8123,N_7958,N_7981);
xor U8124 (N_8124,N_7848,N_7885);
nor U8125 (N_8125,N_7804,N_7892);
or U8126 (N_8126,N_7960,N_7853);
nor U8127 (N_8127,N_7805,N_7931);
xnor U8128 (N_8128,N_7987,N_7910);
and U8129 (N_8129,N_7918,N_7947);
nor U8130 (N_8130,N_7818,N_7813);
xnor U8131 (N_8131,N_7922,N_7886);
or U8132 (N_8132,N_7957,N_7811);
nand U8133 (N_8133,N_7860,N_7961);
nor U8134 (N_8134,N_7938,N_7993);
and U8135 (N_8135,N_7955,N_7819);
nand U8136 (N_8136,N_7808,N_7977);
or U8137 (N_8137,N_7935,N_7963);
or U8138 (N_8138,N_7858,N_7970);
and U8139 (N_8139,N_7858,N_7855);
nor U8140 (N_8140,N_7988,N_7823);
nor U8141 (N_8141,N_7941,N_7889);
xor U8142 (N_8142,N_7807,N_7844);
or U8143 (N_8143,N_7999,N_7925);
or U8144 (N_8144,N_7872,N_7803);
or U8145 (N_8145,N_7817,N_7970);
or U8146 (N_8146,N_7894,N_7976);
xnor U8147 (N_8147,N_7953,N_7938);
and U8148 (N_8148,N_7876,N_7802);
nand U8149 (N_8149,N_7808,N_7959);
nand U8150 (N_8150,N_7830,N_7862);
nor U8151 (N_8151,N_7885,N_7855);
nor U8152 (N_8152,N_7975,N_7897);
or U8153 (N_8153,N_7883,N_7884);
and U8154 (N_8154,N_7884,N_7984);
nand U8155 (N_8155,N_7908,N_7962);
nor U8156 (N_8156,N_7878,N_7912);
and U8157 (N_8157,N_7926,N_7946);
and U8158 (N_8158,N_7883,N_7834);
or U8159 (N_8159,N_7959,N_7909);
or U8160 (N_8160,N_7874,N_7891);
xor U8161 (N_8161,N_7998,N_7945);
or U8162 (N_8162,N_7899,N_7972);
or U8163 (N_8163,N_7945,N_7960);
nand U8164 (N_8164,N_7815,N_7904);
and U8165 (N_8165,N_7865,N_7808);
nor U8166 (N_8166,N_7843,N_7945);
or U8167 (N_8167,N_7849,N_7813);
and U8168 (N_8168,N_7890,N_7999);
nand U8169 (N_8169,N_7992,N_7965);
or U8170 (N_8170,N_7937,N_7864);
nand U8171 (N_8171,N_7805,N_7987);
or U8172 (N_8172,N_7942,N_7817);
xor U8173 (N_8173,N_7871,N_7868);
and U8174 (N_8174,N_7810,N_7932);
and U8175 (N_8175,N_7940,N_7904);
nand U8176 (N_8176,N_7821,N_7988);
and U8177 (N_8177,N_7864,N_7920);
or U8178 (N_8178,N_7927,N_7964);
or U8179 (N_8179,N_7813,N_7814);
xor U8180 (N_8180,N_7856,N_7998);
and U8181 (N_8181,N_7916,N_7835);
nor U8182 (N_8182,N_7845,N_7880);
or U8183 (N_8183,N_7871,N_7980);
and U8184 (N_8184,N_7948,N_7942);
and U8185 (N_8185,N_7822,N_7808);
nor U8186 (N_8186,N_7941,N_7813);
xor U8187 (N_8187,N_7865,N_7937);
or U8188 (N_8188,N_7973,N_7854);
or U8189 (N_8189,N_7860,N_7825);
nor U8190 (N_8190,N_7867,N_7994);
nand U8191 (N_8191,N_7873,N_7884);
xor U8192 (N_8192,N_7976,N_7897);
or U8193 (N_8193,N_7928,N_7970);
or U8194 (N_8194,N_7923,N_7990);
or U8195 (N_8195,N_7933,N_7809);
nand U8196 (N_8196,N_7818,N_7897);
xnor U8197 (N_8197,N_7934,N_7894);
and U8198 (N_8198,N_7896,N_7846);
and U8199 (N_8199,N_7881,N_7944);
nand U8200 (N_8200,N_8142,N_8153);
nor U8201 (N_8201,N_8161,N_8192);
nor U8202 (N_8202,N_8120,N_8118);
and U8203 (N_8203,N_8176,N_8149);
xnor U8204 (N_8204,N_8177,N_8012);
nor U8205 (N_8205,N_8171,N_8003);
nand U8206 (N_8206,N_8134,N_8129);
and U8207 (N_8207,N_8045,N_8019);
and U8208 (N_8208,N_8108,N_8007);
and U8209 (N_8209,N_8035,N_8094);
nor U8210 (N_8210,N_8160,N_8029);
xnor U8211 (N_8211,N_8135,N_8180);
nand U8212 (N_8212,N_8126,N_8158);
nor U8213 (N_8213,N_8167,N_8106);
nand U8214 (N_8214,N_8086,N_8021);
and U8215 (N_8215,N_8138,N_8119);
xnor U8216 (N_8216,N_8146,N_8066);
and U8217 (N_8217,N_8165,N_8091);
and U8218 (N_8218,N_8057,N_8162);
xor U8219 (N_8219,N_8103,N_8078);
xnor U8220 (N_8220,N_8175,N_8048);
nor U8221 (N_8221,N_8133,N_8122);
nand U8222 (N_8222,N_8024,N_8111);
and U8223 (N_8223,N_8184,N_8069);
or U8224 (N_8224,N_8156,N_8101);
nand U8225 (N_8225,N_8185,N_8014);
xor U8226 (N_8226,N_8198,N_8015);
or U8227 (N_8227,N_8168,N_8063);
and U8228 (N_8228,N_8163,N_8102);
or U8229 (N_8229,N_8052,N_8188);
or U8230 (N_8230,N_8089,N_8056);
or U8231 (N_8231,N_8082,N_8186);
nand U8232 (N_8232,N_8125,N_8193);
xor U8233 (N_8233,N_8020,N_8178);
and U8234 (N_8234,N_8050,N_8047);
and U8235 (N_8235,N_8055,N_8154);
or U8236 (N_8236,N_8009,N_8110);
nand U8237 (N_8237,N_8034,N_8013);
nand U8238 (N_8238,N_8004,N_8017);
and U8239 (N_8239,N_8025,N_8073);
or U8240 (N_8240,N_8005,N_8112);
nand U8241 (N_8241,N_8145,N_8059);
nand U8242 (N_8242,N_8010,N_8183);
or U8243 (N_8243,N_8137,N_8113);
or U8244 (N_8244,N_8051,N_8194);
or U8245 (N_8245,N_8100,N_8088);
nand U8246 (N_8246,N_8011,N_8084);
and U8247 (N_8247,N_8123,N_8182);
xnor U8248 (N_8248,N_8130,N_8109);
nor U8249 (N_8249,N_8097,N_8022);
and U8250 (N_8250,N_8117,N_8199);
nor U8251 (N_8251,N_8053,N_8040);
nand U8252 (N_8252,N_8061,N_8077);
or U8253 (N_8253,N_8174,N_8043);
xor U8254 (N_8254,N_8038,N_8008);
nor U8255 (N_8255,N_8189,N_8187);
and U8256 (N_8256,N_8087,N_8002);
nor U8257 (N_8257,N_8042,N_8152);
or U8258 (N_8258,N_8181,N_8131);
and U8259 (N_8259,N_8070,N_8068);
and U8260 (N_8260,N_8169,N_8143);
xnor U8261 (N_8261,N_8058,N_8046);
nand U8262 (N_8262,N_8132,N_8067);
nand U8263 (N_8263,N_8157,N_8018);
xnor U8264 (N_8264,N_8166,N_8054);
xnor U8265 (N_8265,N_8027,N_8136);
xor U8266 (N_8266,N_8060,N_8036);
xor U8267 (N_8267,N_8096,N_8032);
or U8268 (N_8268,N_8028,N_8000);
or U8269 (N_8269,N_8093,N_8075);
nor U8270 (N_8270,N_8127,N_8172);
or U8271 (N_8271,N_8006,N_8116);
nor U8272 (N_8272,N_8124,N_8033);
nand U8273 (N_8273,N_8071,N_8115);
nand U8274 (N_8274,N_8105,N_8148);
or U8275 (N_8275,N_8121,N_8173);
and U8276 (N_8276,N_8023,N_8114);
and U8277 (N_8277,N_8140,N_8065);
nor U8278 (N_8278,N_8044,N_8076);
nor U8279 (N_8279,N_8141,N_8090);
or U8280 (N_8280,N_8095,N_8179);
nand U8281 (N_8281,N_8197,N_8037);
nand U8282 (N_8282,N_8079,N_8195);
and U8283 (N_8283,N_8098,N_8190);
xor U8284 (N_8284,N_8170,N_8026);
or U8285 (N_8285,N_8016,N_8062);
xor U8286 (N_8286,N_8196,N_8039);
and U8287 (N_8287,N_8151,N_8064);
nand U8288 (N_8288,N_8001,N_8159);
xor U8289 (N_8289,N_8072,N_8139);
or U8290 (N_8290,N_8107,N_8099);
and U8291 (N_8291,N_8074,N_8031);
nand U8292 (N_8292,N_8041,N_8147);
and U8293 (N_8293,N_8144,N_8049);
or U8294 (N_8294,N_8030,N_8092);
nor U8295 (N_8295,N_8104,N_8150);
nor U8296 (N_8296,N_8081,N_8128);
and U8297 (N_8297,N_8080,N_8155);
nand U8298 (N_8298,N_8083,N_8085);
or U8299 (N_8299,N_8164,N_8191);
nor U8300 (N_8300,N_8073,N_8146);
xnor U8301 (N_8301,N_8049,N_8125);
xor U8302 (N_8302,N_8184,N_8084);
or U8303 (N_8303,N_8017,N_8091);
and U8304 (N_8304,N_8136,N_8175);
and U8305 (N_8305,N_8035,N_8041);
xnor U8306 (N_8306,N_8048,N_8057);
nand U8307 (N_8307,N_8192,N_8136);
xor U8308 (N_8308,N_8007,N_8027);
nand U8309 (N_8309,N_8081,N_8162);
and U8310 (N_8310,N_8055,N_8123);
nor U8311 (N_8311,N_8085,N_8111);
or U8312 (N_8312,N_8091,N_8056);
nand U8313 (N_8313,N_8104,N_8179);
nor U8314 (N_8314,N_8112,N_8067);
nand U8315 (N_8315,N_8036,N_8084);
xnor U8316 (N_8316,N_8000,N_8113);
xor U8317 (N_8317,N_8100,N_8057);
nor U8318 (N_8318,N_8119,N_8143);
xnor U8319 (N_8319,N_8008,N_8195);
xnor U8320 (N_8320,N_8168,N_8138);
or U8321 (N_8321,N_8050,N_8186);
nand U8322 (N_8322,N_8004,N_8028);
nor U8323 (N_8323,N_8117,N_8078);
xor U8324 (N_8324,N_8019,N_8137);
nor U8325 (N_8325,N_8133,N_8083);
or U8326 (N_8326,N_8173,N_8108);
and U8327 (N_8327,N_8194,N_8146);
or U8328 (N_8328,N_8016,N_8042);
or U8329 (N_8329,N_8105,N_8081);
xor U8330 (N_8330,N_8130,N_8062);
nor U8331 (N_8331,N_8082,N_8133);
and U8332 (N_8332,N_8142,N_8020);
nand U8333 (N_8333,N_8074,N_8024);
nand U8334 (N_8334,N_8004,N_8019);
or U8335 (N_8335,N_8171,N_8009);
xor U8336 (N_8336,N_8143,N_8125);
nor U8337 (N_8337,N_8112,N_8184);
nand U8338 (N_8338,N_8110,N_8042);
nor U8339 (N_8339,N_8054,N_8125);
nor U8340 (N_8340,N_8019,N_8026);
or U8341 (N_8341,N_8104,N_8115);
and U8342 (N_8342,N_8113,N_8124);
and U8343 (N_8343,N_8040,N_8179);
or U8344 (N_8344,N_8192,N_8150);
xor U8345 (N_8345,N_8070,N_8042);
nor U8346 (N_8346,N_8034,N_8025);
nor U8347 (N_8347,N_8079,N_8025);
or U8348 (N_8348,N_8001,N_8062);
xnor U8349 (N_8349,N_8032,N_8061);
nor U8350 (N_8350,N_8094,N_8030);
nand U8351 (N_8351,N_8119,N_8186);
and U8352 (N_8352,N_8129,N_8021);
nand U8353 (N_8353,N_8020,N_8032);
xor U8354 (N_8354,N_8193,N_8127);
nand U8355 (N_8355,N_8113,N_8041);
nor U8356 (N_8356,N_8150,N_8081);
or U8357 (N_8357,N_8148,N_8079);
nand U8358 (N_8358,N_8135,N_8119);
nand U8359 (N_8359,N_8059,N_8076);
xnor U8360 (N_8360,N_8144,N_8198);
xnor U8361 (N_8361,N_8154,N_8090);
and U8362 (N_8362,N_8086,N_8157);
xnor U8363 (N_8363,N_8174,N_8037);
xor U8364 (N_8364,N_8027,N_8177);
or U8365 (N_8365,N_8150,N_8023);
and U8366 (N_8366,N_8138,N_8096);
nor U8367 (N_8367,N_8175,N_8095);
nor U8368 (N_8368,N_8046,N_8024);
nor U8369 (N_8369,N_8160,N_8102);
xnor U8370 (N_8370,N_8055,N_8164);
nor U8371 (N_8371,N_8073,N_8086);
nand U8372 (N_8372,N_8089,N_8190);
nor U8373 (N_8373,N_8127,N_8144);
xor U8374 (N_8374,N_8009,N_8077);
or U8375 (N_8375,N_8113,N_8052);
nand U8376 (N_8376,N_8105,N_8035);
nand U8377 (N_8377,N_8118,N_8129);
or U8378 (N_8378,N_8119,N_8036);
and U8379 (N_8379,N_8129,N_8037);
nor U8380 (N_8380,N_8185,N_8091);
and U8381 (N_8381,N_8144,N_8092);
nor U8382 (N_8382,N_8037,N_8156);
and U8383 (N_8383,N_8129,N_8002);
nor U8384 (N_8384,N_8113,N_8185);
nor U8385 (N_8385,N_8014,N_8072);
or U8386 (N_8386,N_8166,N_8127);
or U8387 (N_8387,N_8007,N_8079);
nand U8388 (N_8388,N_8066,N_8025);
nor U8389 (N_8389,N_8092,N_8168);
and U8390 (N_8390,N_8095,N_8114);
and U8391 (N_8391,N_8023,N_8047);
nor U8392 (N_8392,N_8045,N_8168);
nor U8393 (N_8393,N_8093,N_8147);
nor U8394 (N_8394,N_8028,N_8091);
nand U8395 (N_8395,N_8149,N_8185);
nor U8396 (N_8396,N_8007,N_8136);
nand U8397 (N_8397,N_8159,N_8153);
xnor U8398 (N_8398,N_8095,N_8149);
nand U8399 (N_8399,N_8124,N_8199);
nor U8400 (N_8400,N_8380,N_8237);
or U8401 (N_8401,N_8269,N_8200);
or U8402 (N_8402,N_8372,N_8240);
xor U8403 (N_8403,N_8394,N_8228);
and U8404 (N_8404,N_8259,N_8229);
and U8405 (N_8405,N_8387,N_8360);
nand U8406 (N_8406,N_8310,N_8381);
or U8407 (N_8407,N_8329,N_8388);
xor U8408 (N_8408,N_8221,N_8249);
or U8409 (N_8409,N_8293,N_8317);
nand U8410 (N_8410,N_8333,N_8377);
nor U8411 (N_8411,N_8267,N_8276);
nor U8412 (N_8412,N_8318,N_8211);
and U8413 (N_8413,N_8322,N_8358);
xnor U8414 (N_8414,N_8367,N_8206);
and U8415 (N_8415,N_8218,N_8216);
and U8416 (N_8416,N_8363,N_8224);
nor U8417 (N_8417,N_8342,N_8369);
and U8418 (N_8418,N_8327,N_8390);
xnor U8419 (N_8419,N_8371,N_8303);
or U8420 (N_8420,N_8316,N_8313);
nand U8421 (N_8421,N_8279,N_8320);
and U8422 (N_8422,N_8202,N_8278);
nor U8423 (N_8423,N_8384,N_8323);
or U8424 (N_8424,N_8338,N_8283);
nand U8425 (N_8425,N_8289,N_8212);
nor U8426 (N_8426,N_8235,N_8298);
xor U8427 (N_8427,N_8335,N_8217);
xnor U8428 (N_8428,N_8359,N_8364);
and U8429 (N_8429,N_8232,N_8311);
nor U8430 (N_8430,N_8356,N_8348);
or U8431 (N_8431,N_8376,N_8399);
and U8432 (N_8432,N_8368,N_8365);
or U8433 (N_8433,N_8350,N_8246);
or U8434 (N_8434,N_8287,N_8393);
or U8435 (N_8435,N_8203,N_8351);
nand U8436 (N_8436,N_8354,N_8282);
and U8437 (N_8437,N_8286,N_8334);
and U8438 (N_8438,N_8361,N_8225);
or U8439 (N_8439,N_8392,N_8331);
or U8440 (N_8440,N_8397,N_8352);
nor U8441 (N_8441,N_8250,N_8209);
nand U8442 (N_8442,N_8280,N_8353);
and U8443 (N_8443,N_8288,N_8332);
and U8444 (N_8444,N_8213,N_8328);
nand U8445 (N_8445,N_8346,N_8260);
xor U8446 (N_8446,N_8270,N_8277);
nand U8447 (N_8447,N_8349,N_8239);
or U8448 (N_8448,N_8336,N_8324);
or U8449 (N_8449,N_8247,N_8355);
nand U8450 (N_8450,N_8344,N_8208);
xor U8451 (N_8451,N_8326,N_8304);
nand U8452 (N_8452,N_8366,N_8396);
or U8453 (N_8453,N_8220,N_8274);
nand U8454 (N_8454,N_8297,N_8243);
nor U8455 (N_8455,N_8256,N_8284);
or U8456 (N_8456,N_8315,N_8251);
nand U8457 (N_8457,N_8308,N_8378);
nand U8458 (N_8458,N_8252,N_8374);
nor U8459 (N_8459,N_8242,N_8345);
and U8460 (N_8460,N_8226,N_8253);
nor U8461 (N_8461,N_8291,N_8385);
or U8462 (N_8462,N_8244,N_8292);
xor U8463 (N_8463,N_8210,N_8307);
nand U8464 (N_8464,N_8330,N_8296);
nand U8465 (N_8465,N_8238,N_8357);
nor U8466 (N_8466,N_8362,N_8261);
nand U8467 (N_8467,N_8214,N_8248);
xnor U8468 (N_8468,N_8343,N_8271);
nor U8469 (N_8469,N_8285,N_8379);
or U8470 (N_8470,N_8236,N_8272);
nand U8471 (N_8471,N_8231,N_8268);
and U8472 (N_8472,N_8312,N_8201);
or U8473 (N_8473,N_8255,N_8337);
nand U8474 (N_8474,N_8340,N_8264);
xnor U8475 (N_8475,N_8223,N_8227);
or U8476 (N_8476,N_8383,N_8300);
nand U8477 (N_8477,N_8205,N_8302);
xnor U8478 (N_8478,N_8265,N_8222);
or U8479 (N_8479,N_8266,N_8299);
or U8480 (N_8480,N_8281,N_8230);
nand U8481 (N_8481,N_8319,N_8321);
and U8482 (N_8482,N_8395,N_8241);
or U8483 (N_8483,N_8207,N_8306);
nor U8484 (N_8484,N_8262,N_8204);
nand U8485 (N_8485,N_8234,N_8295);
or U8486 (N_8486,N_8294,N_8391);
or U8487 (N_8487,N_8382,N_8301);
or U8488 (N_8488,N_8258,N_8290);
nor U8489 (N_8489,N_8305,N_8341);
nor U8490 (N_8490,N_8245,N_8375);
xor U8491 (N_8491,N_8309,N_8273);
xnor U8492 (N_8492,N_8263,N_8373);
and U8493 (N_8493,N_8389,N_8347);
and U8494 (N_8494,N_8215,N_8233);
nand U8495 (N_8495,N_8398,N_8275);
nor U8496 (N_8496,N_8339,N_8325);
and U8497 (N_8497,N_8254,N_8257);
xnor U8498 (N_8498,N_8219,N_8314);
and U8499 (N_8499,N_8386,N_8370);
nand U8500 (N_8500,N_8210,N_8241);
nand U8501 (N_8501,N_8349,N_8332);
nand U8502 (N_8502,N_8358,N_8209);
xnor U8503 (N_8503,N_8383,N_8396);
nand U8504 (N_8504,N_8311,N_8389);
nand U8505 (N_8505,N_8377,N_8349);
or U8506 (N_8506,N_8259,N_8220);
nand U8507 (N_8507,N_8308,N_8385);
and U8508 (N_8508,N_8289,N_8209);
xnor U8509 (N_8509,N_8241,N_8311);
or U8510 (N_8510,N_8269,N_8239);
or U8511 (N_8511,N_8286,N_8271);
or U8512 (N_8512,N_8324,N_8257);
nor U8513 (N_8513,N_8309,N_8365);
or U8514 (N_8514,N_8217,N_8237);
or U8515 (N_8515,N_8366,N_8330);
xnor U8516 (N_8516,N_8282,N_8200);
or U8517 (N_8517,N_8372,N_8321);
nand U8518 (N_8518,N_8354,N_8285);
nor U8519 (N_8519,N_8339,N_8370);
nand U8520 (N_8520,N_8325,N_8220);
nor U8521 (N_8521,N_8216,N_8324);
nor U8522 (N_8522,N_8277,N_8299);
or U8523 (N_8523,N_8343,N_8252);
xor U8524 (N_8524,N_8233,N_8394);
nand U8525 (N_8525,N_8288,N_8250);
xor U8526 (N_8526,N_8381,N_8290);
and U8527 (N_8527,N_8364,N_8241);
and U8528 (N_8528,N_8278,N_8317);
or U8529 (N_8529,N_8268,N_8308);
or U8530 (N_8530,N_8310,N_8380);
xor U8531 (N_8531,N_8390,N_8340);
or U8532 (N_8532,N_8396,N_8288);
nor U8533 (N_8533,N_8291,N_8221);
and U8534 (N_8534,N_8358,N_8275);
nand U8535 (N_8535,N_8212,N_8335);
xor U8536 (N_8536,N_8223,N_8277);
or U8537 (N_8537,N_8221,N_8338);
and U8538 (N_8538,N_8202,N_8387);
xnor U8539 (N_8539,N_8207,N_8261);
or U8540 (N_8540,N_8347,N_8248);
nand U8541 (N_8541,N_8373,N_8374);
nor U8542 (N_8542,N_8210,N_8213);
and U8543 (N_8543,N_8251,N_8289);
and U8544 (N_8544,N_8269,N_8207);
nor U8545 (N_8545,N_8293,N_8259);
or U8546 (N_8546,N_8370,N_8344);
xnor U8547 (N_8547,N_8316,N_8368);
nand U8548 (N_8548,N_8238,N_8219);
and U8549 (N_8549,N_8291,N_8293);
or U8550 (N_8550,N_8399,N_8286);
xnor U8551 (N_8551,N_8334,N_8209);
xor U8552 (N_8552,N_8348,N_8385);
nor U8553 (N_8553,N_8268,N_8395);
xor U8554 (N_8554,N_8232,N_8354);
xor U8555 (N_8555,N_8272,N_8306);
xnor U8556 (N_8556,N_8391,N_8317);
nand U8557 (N_8557,N_8286,N_8323);
nand U8558 (N_8558,N_8251,N_8325);
or U8559 (N_8559,N_8332,N_8374);
nor U8560 (N_8560,N_8269,N_8352);
nor U8561 (N_8561,N_8381,N_8245);
nor U8562 (N_8562,N_8339,N_8231);
nor U8563 (N_8563,N_8333,N_8223);
and U8564 (N_8564,N_8389,N_8256);
or U8565 (N_8565,N_8272,N_8344);
and U8566 (N_8566,N_8313,N_8346);
xnor U8567 (N_8567,N_8321,N_8259);
and U8568 (N_8568,N_8330,N_8298);
or U8569 (N_8569,N_8268,N_8267);
and U8570 (N_8570,N_8378,N_8375);
or U8571 (N_8571,N_8233,N_8382);
and U8572 (N_8572,N_8372,N_8220);
and U8573 (N_8573,N_8366,N_8221);
nor U8574 (N_8574,N_8333,N_8317);
or U8575 (N_8575,N_8285,N_8338);
nand U8576 (N_8576,N_8216,N_8380);
nor U8577 (N_8577,N_8260,N_8280);
or U8578 (N_8578,N_8266,N_8268);
or U8579 (N_8579,N_8269,N_8278);
and U8580 (N_8580,N_8299,N_8269);
nand U8581 (N_8581,N_8239,N_8281);
nor U8582 (N_8582,N_8297,N_8321);
nor U8583 (N_8583,N_8226,N_8359);
and U8584 (N_8584,N_8293,N_8338);
nand U8585 (N_8585,N_8278,N_8370);
and U8586 (N_8586,N_8262,N_8256);
nand U8587 (N_8587,N_8276,N_8382);
nand U8588 (N_8588,N_8305,N_8349);
nor U8589 (N_8589,N_8303,N_8307);
or U8590 (N_8590,N_8362,N_8266);
nand U8591 (N_8591,N_8206,N_8256);
or U8592 (N_8592,N_8299,N_8387);
nor U8593 (N_8593,N_8304,N_8354);
and U8594 (N_8594,N_8330,N_8204);
and U8595 (N_8595,N_8265,N_8298);
nand U8596 (N_8596,N_8280,N_8227);
or U8597 (N_8597,N_8225,N_8322);
nand U8598 (N_8598,N_8288,N_8326);
nor U8599 (N_8599,N_8221,N_8353);
nor U8600 (N_8600,N_8444,N_8487);
nand U8601 (N_8601,N_8562,N_8573);
and U8602 (N_8602,N_8599,N_8466);
xnor U8603 (N_8603,N_8489,N_8531);
nand U8604 (N_8604,N_8417,N_8585);
nand U8605 (N_8605,N_8414,N_8557);
xor U8606 (N_8606,N_8513,N_8432);
nor U8607 (N_8607,N_8482,N_8518);
nand U8608 (N_8608,N_8552,N_8581);
and U8609 (N_8609,N_8413,N_8535);
and U8610 (N_8610,N_8462,N_8500);
xor U8611 (N_8611,N_8403,N_8407);
nand U8612 (N_8612,N_8577,N_8586);
nand U8613 (N_8613,N_8426,N_8437);
nor U8614 (N_8614,N_8598,N_8569);
or U8615 (N_8615,N_8570,N_8497);
nand U8616 (N_8616,N_8507,N_8543);
or U8617 (N_8617,N_8425,N_8430);
or U8618 (N_8618,N_8514,N_8431);
and U8619 (N_8619,N_8511,N_8589);
or U8620 (N_8620,N_8578,N_8405);
or U8621 (N_8621,N_8490,N_8546);
or U8622 (N_8622,N_8434,N_8449);
or U8623 (N_8623,N_8406,N_8421);
and U8624 (N_8624,N_8488,N_8538);
nand U8625 (N_8625,N_8478,N_8472);
nand U8626 (N_8626,N_8540,N_8469);
xnor U8627 (N_8627,N_8465,N_8526);
nand U8628 (N_8628,N_8503,N_8592);
or U8629 (N_8629,N_8452,N_8549);
or U8630 (N_8630,N_8456,N_8420);
nand U8631 (N_8631,N_8555,N_8568);
nand U8632 (N_8632,N_8429,N_8499);
and U8633 (N_8633,N_8587,N_8433);
nor U8634 (N_8634,N_8508,N_8556);
or U8635 (N_8635,N_8485,N_8590);
or U8636 (N_8636,N_8537,N_8484);
or U8637 (N_8637,N_8498,N_8550);
and U8638 (N_8638,N_8491,N_8460);
and U8639 (N_8639,N_8439,N_8442);
nor U8640 (N_8640,N_8523,N_8560);
and U8641 (N_8641,N_8527,N_8551);
nand U8642 (N_8642,N_8582,N_8597);
and U8643 (N_8643,N_8558,N_8509);
and U8644 (N_8644,N_8541,N_8544);
and U8645 (N_8645,N_8576,N_8445);
and U8646 (N_8646,N_8505,N_8580);
nand U8647 (N_8647,N_8436,N_8474);
nor U8648 (N_8648,N_8402,N_8440);
and U8649 (N_8649,N_8567,N_8565);
nand U8650 (N_8650,N_8423,N_8554);
and U8651 (N_8651,N_8563,N_8506);
or U8652 (N_8652,N_8447,N_8476);
nor U8653 (N_8653,N_8453,N_8411);
or U8654 (N_8654,N_8424,N_8532);
nor U8655 (N_8655,N_8441,N_8528);
nand U8656 (N_8656,N_8483,N_8404);
nor U8657 (N_8657,N_8545,N_8448);
xnor U8658 (N_8658,N_8593,N_8418);
and U8659 (N_8659,N_8400,N_8517);
xnor U8660 (N_8660,N_8471,N_8553);
xnor U8661 (N_8661,N_8416,N_8521);
and U8662 (N_8662,N_8461,N_8409);
and U8663 (N_8663,N_8559,N_8480);
xnor U8664 (N_8664,N_8533,N_8579);
nand U8665 (N_8665,N_8548,N_8492);
nand U8666 (N_8666,N_8455,N_8494);
nand U8667 (N_8667,N_8464,N_8561);
or U8668 (N_8668,N_8501,N_8486);
or U8669 (N_8669,N_8584,N_8596);
nand U8670 (N_8670,N_8525,N_8519);
xor U8671 (N_8671,N_8470,N_8401);
or U8672 (N_8672,N_8529,N_8427);
and U8673 (N_8673,N_8534,N_8536);
nor U8674 (N_8674,N_8571,N_8502);
and U8675 (N_8675,N_8473,N_8419);
nand U8676 (N_8676,N_8564,N_8458);
xor U8677 (N_8677,N_8463,N_8422);
and U8678 (N_8678,N_8495,N_8583);
and U8679 (N_8679,N_8594,N_8591);
and U8680 (N_8680,N_8415,N_8443);
nand U8681 (N_8681,N_8410,N_8504);
or U8682 (N_8682,N_8438,N_8435);
nor U8683 (N_8683,N_8539,N_8459);
or U8684 (N_8684,N_8510,N_8454);
nand U8685 (N_8685,N_8468,N_8574);
and U8686 (N_8686,N_8477,N_8515);
nand U8687 (N_8687,N_8408,N_8595);
nor U8688 (N_8688,N_8566,N_8512);
nor U8689 (N_8689,N_8520,N_8457);
or U8690 (N_8690,N_8446,N_8450);
or U8691 (N_8691,N_8547,N_8588);
xnor U8692 (N_8692,N_8530,N_8524);
xor U8693 (N_8693,N_8493,N_8542);
nor U8694 (N_8694,N_8481,N_8516);
and U8695 (N_8695,N_8572,N_8496);
or U8696 (N_8696,N_8412,N_8522);
nand U8697 (N_8697,N_8467,N_8428);
nor U8698 (N_8698,N_8479,N_8475);
xnor U8699 (N_8699,N_8451,N_8575);
and U8700 (N_8700,N_8509,N_8429);
or U8701 (N_8701,N_8485,N_8574);
nor U8702 (N_8702,N_8559,N_8529);
nor U8703 (N_8703,N_8402,N_8400);
nor U8704 (N_8704,N_8430,N_8560);
nor U8705 (N_8705,N_8443,N_8465);
nor U8706 (N_8706,N_8513,N_8584);
nor U8707 (N_8707,N_8458,N_8482);
nand U8708 (N_8708,N_8569,N_8423);
nand U8709 (N_8709,N_8540,N_8501);
xnor U8710 (N_8710,N_8517,N_8417);
or U8711 (N_8711,N_8448,N_8585);
xor U8712 (N_8712,N_8480,N_8483);
or U8713 (N_8713,N_8467,N_8584);
nor U8714 (N_8714,N_8532,N_8480);
nor U8715 (N_8715,N_8425,N_8404);
and U8716 (N_8716,N_8444,N_8579);
and U8717 (N_8717,N_8498,N_8421);
or U8718 (N_8718,N_8547,N_8486);
and U8719 (N_8719,N_8459,N_8578);
and U8720 (N_8720,N_8549,N_8447);
xor U8721 (N_8721,N_8534,N_8572);
xor U8722 (N_8722,N_8534,N_8532);
nor U8723 (N_8723,N_8490,N_8462);
or U8724 (N_8724,N_8561,N_8546);
and U8725 (N_8725,N_8485,N_8540);
xnor U8726 (N_8726,N_8594,N_8522);
and U8727 (N_8727,N_8556,N_8550);
xnor U8728 (N_8728,N_8538,N_8487);
xor U8729 (N_8729,N_8554,N_8472);
xnor U8730 (N_8730,N_8583,N_8483);
and U8731 (N_8731,N_8405,N_8582);
and U8732 (N_8732,N_8499,N_8512);
nand U8733 (N_8733,N_8567,N_8400);
nor U8734 (N_8734,N_8467,N_8571);
or U8735 (N_8735,N_8552,N_8442);
nand U8736 (N_8736,N_8413,N_8593);
or U8737 (N_8737,N_8407,N_8543);
nor U8738 (N_8738,N_8452,N_8471);
nor U8739 (N_8739,N_8539,N_8464);
and U8740 (N_8740,N_8558,N_8511);
nand U8741 (N_8741,N_8524,N_8593);
xor U8742 (N_8742,N_8596,N_8446);
nand U8743 (N_8743,N_8419,N_8487);
and U8744 (N_8744,N_8441,N_8598);
nor U8745 (N_8745,N_8533,N_8527);
or U8746 (N_8746,N_8411,N_8532);
and U8747 (N_8747,N_8470,N_8412);
and U8748 (N_8748,N_8508,N_8484);
nand U8749 (N_8749,N_8422,N_8447);
xor U8750 (N_8750,N_8428,N_8481);
and U8751 (N_8751,N_8506,N_8540);
xnor U8752 (N_8752,N_8425,N_8446);
nand U8753 (N_8753,N_8475,N_8486);
nand U8754 (N_8754,N_8584,N_8588);
nor U8755 (N_8755,N_8531,N_8400);
or U8756 (N_8756,N_8571,N_8511);
nor U8757 (N_8757,N_8480,N_8535);
and U8758 (N_8758,N_8428,N_8477);
and U8759 (N_8759,N_8517,N_8529);
xnor U8760 (N_8760,N_8450,N_8570);
or U8761 (N_8761,N_8504,N_8558);
nand U8762 (N_8762,N_8477,N_8561);
xnor U8763 (N_8763,N_8487,N_8434);
xnor U8764 (N_8764,N_8400,N_8491);
nand U8765 (N_8765,N_8553,N_8584);
xnor U8766 (N_8766,N_8554,N_8534);
and U8767 (N_8767,N_8516,N_8424);
or U8768 (N_8768,N_8452,N_8466);
and U8769 (N_8769,N_8456,N_8467);
or U8770 (N_8770,N_8490,N_8480);
nor U8771 (N_8771,N_8405,N_8469);
nand U8772 (N_8772,N_8439,N_8451);
xnor U8773 (N_8773,N_8585,N_8582);
and U8774 (N_8774,N_8523,N_8463);
nor U8775 (N_8775,N_8590,N_8584);
and U8776 (N_8776,N_8540,N_8427);
nor U8777 (N_8777,N_8451,N_8483);
or U8778 (N_8778,N_8527,N_8534);
or U8779 (N_8779,N_8499,N_8505);
or U8780 (N_8780,N_8539,N_8599);
xor U8781 (N_8781,N_8595,N_8466);
and U8782 (N_8782,N_8423,N_8565);
or U8783 (N_8783,N_8530,N_8539);
nor U8784 (N_8784,N_8490,N_8475);
nor U8785 (N_8785,N_8594,N_8534);
or U8786 (N_8786,N_8503,N_8541);
xnor U8787 (N_8787,N_8442,N_8479);
nand U8788 (N_8788,N_8476,N_8453);
xnor U8789 (N_8789,N_8555,N_8486);
nor U8790 (N_8790,N_8532,N_8576);
nand U8791 (N_8791,N_8520,N_8468);
and U8792 (N_8792,N_8549,N_8568);
or U8793 (N_8793,N_8496,N_8521);
nand U8794 (N_8794,N_8426,N_8453);
or U8795 (N_8795,N_8577,N_8571);
or U8796 (N_8796,N_8499,N_8581);
and U8797 (N_8797,N_8492,N_8469);
or U8798 (N_8798,N_8442,N_8411);
and U8799 (N_8799,N_8462,N_8461);
and U8800 (N_8800,N_8673,N_8739);
nor U8801 (N_8801,N_8605,N_8670);
or U8802 (N_8802,N_8731,N_8793);
nand U8803 (N_8803,N_8666,N_8720);
or U8804 (N_8804,N_8736,N_8622);
nand U8805 (N_8805,N_8613,N_8697);
or U8806 (N_8806,N_8600,N_8692);
nor U8807 (N_8807,N_8758,N_8761);
or U8808 (N_8808,N_8752,N_8764);
nand U8809 (N_8809,N_8616,N_8661);
nand U8810 (N_8810,N_8647,N_8745);
xnor U8811 (N_8811,N_8615,N_8729);
and U8812 (N_8812,N_8783,N_8672);
nand U8813 (N_8813,N_8728,N_8723);
nand U8814 (N_8814,N_8707,N_8799);
xor U8815 (N_8815,N_8791,N_8663);
nor U8816 (N_8816,N_8669,N_8769);
nand U8817 (N_8817,N_8607,N_8631);
nand U8818 (N_8818,N_8696,N_8685);
nor U8819 (N_8819,N_8637,N_8733);
xor U8820 (N_8820,N_8694,N_8727);
and U8821 (N_8821,N_8762,N_8742);
nand U8822 (N_8822,N_8650,N_8784);
or U8823 (N_8823,N_8687,N_8734);
xor U8824 (N_8824,N_8725,N_8660);
xor U8825 (N_8825,N_8747,N_8618);
nor U8826 (N_8826,N_8610,N_8743);
nand U8827 (N_8827,N_8778,N_8676);
or U8828 (N_8828,N_8681,N_8744);
nand U8829 (N_8829,N_8726,N_8780);
nor U8830 (N_8830,N_8656,N_8732);
or U8831 (N_8831,N_8754,N_8710);
or U8832 (N_8832,N_8738,N_8782);
and U8833 (N_8833,N_8774,N_8621);
nand U8834 (N_8834,N_8716,N_8679);
nand U8835 (N_8835,N_8722,N_8649);
and U8836 (N_8836,N_8604,N_8737);
or U8837 (N_8837,N_8624,N_8628);
nor U8838 (N_8838,N_8794,N_8682);
nor U8839 (N_8839,N_8635,N_8639);
or U8840 (N_8840,N_8705,N_8788);
or U8841 (N_8841,N_8662,N_8627);
nand U8842 (N_8842,N_8792,N_8735);
nor U8843 (N_8843,N_8766,N_8689);
xor U8844 (N_8844,N_8638,N_8702);
nor U8845 (N_8845,N_8773,N_8648);
xnor U8846 (N_8846,N_8797,N_8675);
or U8847 (N_8847,N_8630,N_8760);
nand U8848 (N_8848,N_8636,N_8677);
or U8849 (N_8849,N_8659,N_8775);
nor U8850 (N_8850,N_8645,N_8688);
nor U8851 (N_8851,N_8763,N_8750);
nand U8852 (N_8852,N_8704,N_8686);
xor U8853 (N_8853,N_8796,N_8608);
nor U8854 (N_8854,N_8785,N_8641);
nand U8855 (N_8855,N_8644,N_8714);
or U8856 (N_8856,N_8625,N_8700);
xnor U8857 (N_8857,N_8632,N_8768);
xnor U8858 (N_8858,N_8711,N_8602);
xnor U8859 (N_8859,N_8620,N_8718);
or U8860 (N_8860,N_8695,N_8671);
nand U8861 (N_8861,N_8614,N_8642);
nor U8862 (N_8862,N_8756,N_8798);
or U8863 (N_8863,N_8717,N_8629);
or U8864 (N_8864,N_8612,N_8703);
nor U8865 (N_8865,N_8651,N_8643);
or U8866 (N_8866,N_8684,N_8713);
xor U8867 (N_8867,N_8789,N_8668);
or U8868 (N_8868,N_8701,N_8748);
or U8869 (N_8869,N_8683,N_8776);
nor U8870 (N_8870,N_8712,N_8779);
xor U8871 (N_8871,N_8772,N_8657);
or U8872 (N_8872,N_8740,N_8787);
nand U8873 (N_8873,N_8652,N_8640);
nor U8874 (N_8874,N_8653,N_8757);
or U8875 (N_8875,N_8795,N_8746);
nor U8876 (N_8876,N_8724,N_8658);
nand U8877 (N_8877,N_8655,N_8665);
xnor U8878 (N_8878,N_8617,N_8606);
xor U8879 (N_8879,N_8759,N_8634);
xnor U8880 (N_8880,N_8646,N_8715);
or U8881 (N_8881,N_8693,N_8730);
or U8882 (N_8882,N_8633,N_8708);
or U8883 (N_8883,N_8664,N_8751);
or U8884 (N_8884,N_8786,N_8749);
xnor U8885 (N_8885,N_8690,N_8699);
nand U8886 (N_8886,N_8667,N_8706);
xnor U8887 (N_8887,N_8765,N_8623);
or U8888 (N_8888,N_8626,N_8709);
or U8889 (N_8889,N_8680,N_8721);
and U8890 (N_8890,N_8678,N_8619);
nand U8891 (N_8891,N_8767,N_8609);
xor U8892 (N_8892,N_8753,N_8654);
xnor U8893 (N_8893,N_8698,N_8601);
xnor U8894 (N_8894,N_8781,N_8603);
nor U8895 (N_8895,N_8755,N_8691);
xnor U8896 (N_8896,N_8790,N_8741);
xnor U8897 (N_8897,N_8770,N_8719);
or U8898 (N_8898,N_8771,N_8674);
and U8899 (N_8899,N_8777,N_8611);
or U8900 (N_8900,N_8621,N_8616);
xor U8901 (N_8901,N_8652,N_8753);
nor U8902 (N_8902,N_8675,N_8763);
xnor U8903 (N_8903,N_8791,N_8648);
nand U8904 (N_8904,N_8650,N_8638);
and U8905 (N_8905,N_8790,N_8673);
nor U8906 (N_8906,N_8769,N_8663);
or U8907 (N_8907,N_8711,N_8688);
nand U8908 (N_8908,N_8786,N_8748);
xnor U8909 (N_8909,N_8602,N_8657);
xnor U8910 (N_8910,N_8759,N_8728);
xor U8911 (N_8911,N_8703,N_8631);
nand U8912 (N_8912,N_8685,N_8782);
nor U8913 (N_8913,N_8620,N_8749);
nand U8914 (N_8914,N_8629,N_8735);
or U8915 (N_8915,N_8770,N_8747);
nand U8916 (N_8916,N_8764,N_8746);
or U8917 (N_8917,N_8674,N_8668);
xor U8918 (N_8918,N_8770,N_8635);
nand U8919 (N_8919,N_8752,N_8602);
xor U8920 (N_8920,N_8798,N_8750);
xnor U8921 (N_8921,N_8607,N_8696);
nand U8922 (N_8922,N_8724,N_8728);
or U8923 (N_8923,N_8634,N_8726);
nand U8924 (N_8924,N_8609,N_8694);
nand U8925 (N_8925,N_8772,N_8698);
and U8926 (N_8926,N_8785,N_8754);
or U8927 (N_8927,N_8736,N_8678);
nor U8928 (N_8928,N_8657,N_8775);
and U8929 (N_8929,N_8730,N_8661);
and U8930 (N_8930,N_8602,N_8764);
nand U8931 (N_8931,N_8671,N_8785);
and U8932 (N_8932,N_8731,N_8759);
or U8933 (N_8933,N_8674,N_8655);
and U8934 (N_8934,N_8621,N_8700);
nor U8935 (N_8935,N_8628,N_8743);
or U8936 (N_8936,N_8687,N_8740);
xnor U8937 (N_8937,N_8647,N_8668);
or U8938 (N_8938,N_8779,N_8719);
nand U8939 (N_8939,N_8764,N_8674);
nand U8940 (N_8940,N_8635,N_8678);
nor U8941 (N_8941,N_8694,N_8691);
or U8942 (N_8942,N_8618,N_8641);
and U8943 (N_8943,N_8644,N_8604);
xnor U8944 (N_8944,N_8699,N_8684);
nor U8945 (N_8945,N_8756,N_8753);
nor U8946 (N_8946,N_8783,N_8640);
nand U8947 (N_8947,N_8794,N_8603);
and U8948 (N_8948,N_8641,N_8615);
or U8949 (N_8949,N_8675,N_8738);
xor U8950 (N_8950,N_8787,N_8647);
and U8951 (N_8951,N_8654,N_8691);
or U8952 (N_8952,N_8680,N_8700);
nor U8953 (N_8953,N_8752,N_8695);
or U8954 (N_8954,N_8613,N_8687);
or U8955 (N_8955,N_8673,N_8610);
and U8956 (N_8956,N_8747,N_8781);
nand U8957 (N_8957,N_8776,N_8717);
xor U8958 (N_8958,N_8752,N_8625);
xnor U8959 (N_8959,N_8668,N_8634);
or U8960 (N_8960,N_8618,N_8710);
or U8961 (N_8961,N_8651,N_8780);
and U8962 (N_8962,N_8603,N_8744);
nand U8963 (N_8963,N_8740,N_8762);
xor U8964 (N_8964,N_8750,N_8666);
nor U8965 (N_8965,N_8755,N_8644);
nand U8966 (N_8966,N_8743,N_8726);
or U8967 (N_8967,N_8729,N_8779);
nor U8968 (N_8968,N_8683,N_8653);
xnor U8969 (N_8969,N_8617,N_8781);
and U8970 (N_8970,N_8778,N_8785);
or U8971 (N_8971,N_8607,N_8688);
nand U8972 (N_8972,N_8711,N_8600);
and U8973 (N_8973,N_8676,N_8733);
or U8974 (N_8974,N_8740,N_8665);
xnor U8975 (N_8975,N_8732,N_8680);
nand U8976 (N_8976,N_8624,N_8722);
nand U8977 (N_8977,N_8660,N_8635);
or U8978 (N_8978,N_8748,N_8643);
xnor U8979 (N_8979,N_8737,N_8622);
and U8980 (N_8980,N_8610,N_8755);
nor U8981 (N_8981,N_8754,N_8656);
and U8982 (N_8982,N_8643,N_8714);
xor U8983 (N_8983,N_8618,N_8616);
nand U8984 (N_8984,N_8631,N_8760);
and U8985 (N_8985,N_8620,N_8615);
nor U8986 (N_8986,N_8795,N_8754);
or U8987 (N_8987,N_8675,N_8646);
xnor U8988 (N_8988,N_8763,N_8658);
and U8989 (N_8989,N_8705,N_8701);
nand U8990 (N_8990,N_8718,N_8746);
nor U8991 (N_8991,N_8674,N_8770);
and U8992 (N_8992,N_8629,N_8622);
and U8993 (N_8993,N_8745,N_8751);
xnor U8994 (N_8994,N_8778,N_8700);
or U8995 (N_8995,N_8728,N_8789);
and U8996 (N_8996,N_8643,N_8609);
nand U8997 (N_8997,N_8755,N_8637);
or U8998 (N_8998,N_8607,N_8729);
and U8999 (N_8999,N_8687,N_8768);
nor U9000 (N_9000,N_8824,N_8856);
xnor U9001 (N_9001,N_8850,N_8876);
xor U9002 (N_9002,N_8842,N_8955);
xnor U9003 (N_9003,N_8880,N_8898);
nor U9004 (N_9004,N_8970,N_8813);
nand U9005 (N_9005,N_8940,N_8860);
or U9006 (N_9006,N_8868,N_8874);
nor U9007 (N_9007,N_8869,N_8957);
nor U9008 (N_9008,N_8812,N_8895);
or U9009 (N_9009,N_8924,N_8975);
xor U9010 (N_9010,N_8831,N_8980);
nand U9011 (N_9011,N_8901,N_8804);
xnor U9012 (N_9012,N_8973,N_8990);
or U9013 (N_9013,N_8949,N_8841);
nand U9014 (N_9014,N_8838,N_8912);
xnor U9015 (N_9015,N_8892,N_8821);
and U9016 (N_9016,N_8968,N_8918);
nand U9017 (N_9017,N_8861,N_8986);
nand U9018 (N_9018,N_8997,N_8839);
nor U9019 (N_9019,N_8849,N_8829);
and U9020 (N_9020,N_8891,N_8884);
xnor U9021 (N_9021,N_8988,N_8864);
nor U9022 (N_9022,N_8843,N_8858);
or U9023 (N_9023,N_8866,N_8826);
xor U9024 (N_9024,N_8832,N_8886);
or U9025 (N_9025,N_8919,N_8888);
xnor U9026 (N_9026,N_8974,N_8966);
xor U9027 (N_9027,N_8930,N_8904);
or U9028 (N_9028,N_8983,N_8854);
and U9029 (N_9029,N_8873,N_8865);
nor U9030 (N_9030,N_8808,N_8967);
xor U9031 (N_9031,N_8942,N_8945);
xor U9032 (N_9032,N_8987,N_8885);
nand U9033 (N_9033,N_8846,N_8943);
and U9034 (N_9034,N_8897,N_8837);
or U9035 (N_9035,N_8823,N_8879);
nand U9036 (N_9036,N_8972,N_8996);
xnor U9037 (N_9037,N_8999,N_8969);
nor U9038 (N_9038,N_8902,N_8925);
or U9039 (N_9039,N_8870,N_8907);
or U9040 (N_9040,N_8903,N_8931);
nor U9041 (N_9041,N_8862,N_8852);
nand U9042 (N_9042,N_8828,N_8887);
and U9043 (N_9043,N_8857,N_8899);
nor U9044 (N_9044,N_8917,N_8819);
nor U9045 (N_9045,N_8953,N_8991);
or U9046 (N_9046,N_8995,N_8989);
nand U9047 (N_9047,N_8805,N_8913);
or U9048 (N_9048,N_8905,N_8994);
or U9049 (N_9049,N_8802,N_8954);
nand U9050 (N_9050,N_8937,N_8948);
and U9051 (N_9051,N_8863,N_8810);
nor U9052 (N_9052,N_8911,N_8836);
or U9053 (N_9053,N_8883,N_8827);
or U9054 (N_9054,N_8906,N_8801);
nand U9055 (N_9055,N_8803,N_8908);
and U9056 (N_9056,N_8951,N_8878);
and U9057 (N_9057,N_8992,N_8978);
xnor U9058 (N_9058,N_8914,N_8835);
xnor U9059 (N_9059,N_8882,N_8981);
and U9060 (N_9060,N_8960,N_8872);
nor U9061 (N_9061,N_8933,N_8946);
nor U9062 (N_9062,N_8890,N_8947);
xnor U9063 (N_9063,N_8847,N_8815);
or U9064 (N_9064,N_8859,N_8923);
nor U9065 (N_9065,N_8932,N_8964);
nor U9066 (N_9066,N_8845,N_8928);
nand U9067 (N_9067,N_8977,N_8825);
nor U9068 (N_9068,N_8920,N_8929);
xor U9069 (N_9069,N_8922,N_8984);
nand U9070 (N_9070,N_8935,N_8822);
or U9071 (N_9071,N_8963,N_8851);
xnor U9072 (N_9072,N_8962,N_8806);
and U9073 (N_9073,N_8959,N_8848);
nor U9074 (N_9074,N_8910,N_8915);
nor U9075 (N_9075,N_8844,N_8976);
nand U9076 (N_9076,N_8900,N_8971);
xor U9077 (N_9077,N_8867,N_8871);
xnor U9078 (N_9078,N_8958,N_8820);
xor U9079 (N_9079,N_8853,N_8855);
nor U9080 (N_9080,N_8833,N_8926);
and U9081 (N_9081,N_8840,N_8965);
or U9082 (N_9082,N_8961,N_8800);
nor U9083 (N_9083,N_8881,N_8894);
xor U9084 (N_9084,N_8936,N_8950);
or U9085 (N_9085,N_8877,N_8921);
nor U9086 (N_9086,N_8939,N_8982);
nor U9087 (N_9087,N_8944,N_8993);
nand U9088 (N_9088,N_8811,N_8875);
or U9089 (N_9089,N_8893,N_8809);
nor U9090 (N_9090,N_8938,N_8889);
nand U9091 (N_9091,N_8979,N_8916);
nand U9092 (N_9092,N_8817,N_8952);
and U9093 (N_9093,N_8896,N_8934);
nand U9094 (N_9094,N_8998,N_8941);
or U9095 (N_9095,N_8834,N_8956);
xor U9096 (N_9096,N_8807,N_8830);
nand U9097 (N_9097,N_8909,N_8814);
nand U9098 (N_9098,N_8816,N_8818);
and U9099 (N_9099,N_8985,N_8927);
or U9100 (N_9100,N_8815,N_8938);
or U9101 (N_9101,N_8966,N_8803);
nand U9102 (N_9102,N_8871,N_8885);
and U9103 (N_9103,N_8971,N_8941);
or U9104 (N_9104,N_8876,N_8940);
and U9105 (N_9105,N_8879,N_8988);
or U9106 (N_9106,N_8884,N_8971);
or U9107 (N_9107,N_8971,N_8878);
or U9108 (N_9108,N_8918,N_8976);
or U9109 (N_9109,N_8875,N_8825);
and U9110 (N_9110,N_8884,N_8859);
xnor U9111 (N_9111,N_8907,N_8815);
nor U9112 (N_9112,N_8975,N_8840);
nor U9113 (N_9113,N_8876,N_8823);
and U9114 (N_9114,N_8822,N_8910);
or U9115 (N_9115,N_8860,N_8975);
or U9116 (N_9116,N_8885,N_8807);
or U9117 (N_9117,N_8956,N_8992);
nor U9118 (N_9118,N_8993,N_8819);
and U9119 (N_9119,N_8802,N_8959);
and U9120 (N_9120,N_8954,N_8889);
nor U9121 (N_9121,N_8832,N_8816);
nand U9122 (N_9122,N_8861,N_8867);
xor U9123 (N_9123,N_8886,N_8928);
nor U9124 (N_9124,N_8909,N_8956);
nand U9125 (N_9125,N_8817,N_8860);
nand U9126 (N_9126,N_8841,N_8921);
xor U9127 (N_9127,N_8952,N_8862);
and U9128 (N_9128,N_8859,N_8928);
nor U9129 (N_9129,N_8933,N_8867);
and U9130 (N_9130,N_8952,N_8860);
and U9131 (N_9131,N_8809,N_8912);
nand U9132 (N_9132,N_8823,N_8861);
and U9133 (N_9133,N_8944,N_8896);
and U9134 (N_9134,N_8996,N_8925);
xnor U9135 (N_9135,N_8882,N_8956);
xor U9136 (N_9136,N_8873,N_8899);
or U9137 (N_9137,N_8944,N_8943);
nand U9138 (N_9138,N_8837,N_8999);
nor U9139 (N_9139,N_8930,N_8851);
nor U9140 (N_9140,N_8969,N_8949);
and U9141 (N_9141,N_8904,N_8931);
or U9142 (N_9142,N_8946,N_8989);
or U9143 (N_9143,N_8917,N_8857);
xnor U9144 (N_9144,N_8834,N_8899);
nand U9145 (N_9145,N_8884,N_8946);
xor U9146 (N_9146,N_8883,N_8905);
or U9147 (N_9147,N_8905,N_8858);
nand U9148 (N_9148,N_8873,N_8992);
xor U9149 (N_9149,N_8865,N_8925);
and U9150 (N_9150,N_8933,N_8930);
nand U9151 (N_9151,N_8858,N_8944);
nand U9152 (N_9152,N_8834,N_8949);
nand U9153 (N_9153,N_8970,N_8939);
or U9154 (N_9154,N_8882,N_8859);
nand U9155 (N_9155,N_8881,N_8955);
xnor U9156 (N_9156,N_8849,N_8867);
xnor U9157 (N_9157,N_8802,N_8981);
xor U9158 (N_9158,N_8925,N_8848);
nand U9159 (N_9159,N_8973,N_8858);
nor U9160 (N_9160,N_8826,N_8869);
nand U9161 (N_9161,N_8989,N_8932);
xnor U9162 (N_9162,N_8920,N_8845);
xnor U9163 (N_9163,N_8807,N_8888);
nand U9164 (N_9164,N_8870,N_8904);
nor U9165 (N_9165,N_8973,N_8929);
nor U9166 (N_9166,N_8879,N_8911);
or U9167 (N_9167,N_8830,N_8818);
xor U9168 (N_9168,N_8966,N_8891);
and U9169 (N_9169,N_8903,N_8823);
nand U9170 (N_9170,N_8863,N_8974);
nor U9171 (N_9171,N_8858,N_8820);
and U9172 (N_9172,N_8854,N_8828);
xor U9173 (N_9173,N_8908,N_8834);
or U9174 (N_9174,N_8806,N_8824);
and U9175 (N_9175,N_8832,N_8842);
xor U9176 (N_9176,N_8896,N_8997);
and U9177 (N_9177,N_8827,N_8841);
nor U9178 (N_9178,N_8911,N_8964);
nand U9179 (N_9179,N_8951,N_8930);
nand U9180 (N_9180,N_8896,N_8839);
or U9181 (N_9181,N_8966,N_8960);
and U9182 (N_9182,N_8955,N_8911);
nand U9183 (N_9183,N_8844,N_8885);
or U9184 (N_9184,N_8979,N_8953);
nand U9185 (N_9185,N_8819,N_8960);
xnor U9186 (N_9186,N_8868,N_8826);
and U9187 (N_9187,N_8969,N_8871);
and U9188 (N_9188,N_8992,N_8878);
or U9189 (N_9189,N_8908,N_8828);
and U9190 (N_9190,N_8937,N_8956);
nor U9191 (N_9191,N_8827,N_8866);
nor U9192 (N_9192,N_8920,N_8927);
nand U9193 (N_9193,N_8933,N_8915);
and U9194 (N_9194,N_8956,N_8847);
xnor U9195 (N_9195,N_8837,N_8874);
xor U9196 (N_9196,N_8996,N_8881);
and U9197 (N_9197,N_8945,N_8899);
xor U9198 (N_9198,N_8845,N_8948);
or U9199 (N_9199,N_8813,N_8814);
nor U9200 (N_9200,N_9028,N_9162);
or U9201 (N_9201,N_9055,N_9159);
nand U9202 (N_9202,N_9094,N_9047);
xnor U9203 (N_9203,N_9146,N_9073);
xnor U9204 (N_9204,N_9113,N_9134);
or U9205 (N_9205,N_9096,N_9154);
nand U9206 (N_9206,N_9107,N_9187);
nor U9207 (N_9207,N_9046,N_9072);
nor U9208 (N_9208,N_9034,N_9130);
xor U9209 (N_9209,N_9036,N_9156);
or U9210 (N_9210,N_9062,N_9075);
or U9211 (N_9211,N_9139,N_9179);
and U9212 (N_9212,N_9189,N_9033);
nor U9213 (N_9213,N_9083,N_9129);
xnor U9214 (N_9214,N_9043,N_9005);
or U9215 (N_9215,N_9110,N_9131);
and U9216 (N_9216,N_9050,N_9085);
and U9217 (N_9217,N_9059,N_9174);
nand U9218 (N_9218,N_9183,N_9144);
nand U9219 (N_9219,N_9126,N_9063);
nand U9220 (N_9220,N_9192,N_9120);
xnor U9221 (N_9221,N_9054,N_9136);
and U9222 (N_9222,N_9012,N_9127);
nor U9223 (N_9223,N_9084,N_9178);
nor U9224 (N_9224,N_9194,N_9066);
or U9225 (N_9225,N_9061,N_9020);
or U9226 (N_9226,N_9170,N_9089);
xnor U9227 (N_9227,N_9048,N_9041);
and U9228 (N_9228,N_9155,N_9071);
nor U9229 (N_9229,N_9070,N_9079);
xnor U9230 (N_9230,N_9024,N_9090);
and U9231 (N_9231,N_9147,N_9039);
xnor U9232 (N_9232,N_9140,N_9015);
nor U9233 (N_9233,N_9091,N_9006);
nand U9234 (N_9234,N_9175,N_9009);
nor U9235 (N_9235,N_9186,N_9037);
and U9236 (N_9236,N_9151,N_9188);
nor U9237 (N_9237,N_9051,N_9132);
nor U9238 (N_9238,N_9171,N_9038);
or U9239 (N_9239,N_9088,N_9095);
nand U9240 (N_9240,N_9023,N_9143);
nand U9241 (N_9241,N_9082,N_9161);
or U9242 (N_9242,N_9040,N_9123);
or U9243 (N_9243,N_9199,N_9030);
and U9244 (N_9244,N_9137,N_9153);
and U9245 (N_9245,N_9013,N_9001);
nor U9246 (N_9246,N_9022,N_9058);
nand U9247 (N_9247,N_9027,N_9198);
nor U9248 (N_9248,N_9152,N_9053);
nor U9249 (N_9249,N_9108,N_9104);
xnor U9250 (N_9250,N_9057,N_9182);
xor U9251 (N_9251,N_9169,N_9010);
or U9252 (N_9252,N_9031,N_9026);
nor U9253 (N_9253,N_9135,N_9087);
and U9254 (N_9254,N_9018,N_9068);
nor U9255 (N_9255,N_9021,N_9165);
and U9256 (N_9256,N_9035,N_9029);
nor U9257 (N_9257,N_9017,N_9111);
and U9258 (N_9258,N_9177,N_9116);
nor U9259 (N_9259,N_9185,N_9060);
nand U9260 (N_9260,N_9124,N_9045);
nand U9261 (N_9261,N_9157,N_9191);
nor U9262 (N_9262,N_9007,N_9133);
xor U9263 (N_9263,N_9196,N_9121);
xnor U9264 (N_9264,N_9158,N_9000);
nand U9265 (N_9265,N_9014,N_9052);
and U9266 (N_9266,N_9172,N_9002);
nand U9267 (N_9267,N_9067,N_9180);
or U9268 (N_9268,N_9142,N_9019);
xnor U9269 (N_9269,N_9106,N_9049);
xnor U9270 (N_9270,N_9117,N_9118);
nand U9271 (N_9271,N_9197,N_9016);
nor U9272 (N_9272,N_9069,N_9109);
or U9273 (N_9273,N_9077,N_9150);
or U9274 (N_9274,N_9065,N_9099);
nor U9275 (N_9275,N_9148,N_9093);
and U9276 (N_9276,N_9115,N_9044);
nor U9277 (N_9277,N_9004,N_9122);
nand U9278 (N_9278,N_9074,N_9101);
nand U9279 (N_9279,N_9056,N_9160);
xor U9280 (N_9280,N_9167,N_9176);
or U9281 (N_9281,N_9173,N_9190);
nor U9282 (N_9282,N_9092,N_9098);
nand U9283 (N_9283,N_9081,N_9080);
or U9284 (N_9284,N_9078,N_9103);
nand U9285 (N_9285,N_9112,N_9138);
and U9286 (N_9286,N_9168,N_9195);
or U9287 (N_9287,N_9149,N_9145);
and U9288 (N_9288,N_9119,N_9128);
nor U9289 (N_9289,N_9008,N_9163);
xor U9290 (N_9290,N_9011,N_9076);
and U9291 (N_9291,N_9086,N_9064);
or U9292 (N_9292,N_9166,N_9193);
or U9293 (N_9293,N_9032,N_9025);
xor U9294 (N_9294,N_9097,N_9102);
xor U9295 (N_9295,N_9141,N_9100);
nand U9296 (N_9296,N_9164,N_9125);
xor U9297 (N_9297,N_9114,N_9181);
and U9298 (N_9298,N_9184,N_9105);
or U9299 (N_9299,N_9003,N_9042);
or U9300 (N_9300,N_9047,N_9012);
xnor U9301 (N_9301,N_9041,N_9036);
nand U9302 (N_9302,N_9080,N_9103);
nor U9303 (N_9303,N_9154,N_9198);
nand U9304 (N_9304,N_9091,N_9158);
or U9305 (N_9305,N_9136,N_9170);
nor U9306 (N_9306,N_9161,N_9014);
nor U9307 (N_9307,N_9065,N_9009);
nand U9308 (N_9308,N_9002,N_9048);
or U9309 (N_9309,N_9012,N_9106);
or U9310 (N_9310,N_9073,N_9157);
or U9311 (N_9311,N_9152,N_9039);
or U9312 (N_9312,N_9028,N_9053);
nand U9313 (N_9313,N_9133,N_9039);
xor U9314 (N_9314,N_9043,N_9054);
nand U9315 (N_9315,N_9082,N_9094);
nand U9316 (N_9316,N_9033,N_9058);
nand U9317 (N_9317,N_9095,N_9025);
or U9318 (N_9318,N_9167,N_9158);
and U9319 (N_9319,N_9102,N_9010);
nor U9320 (N_9320,N_9185,N_9161);
nand U9321 (N_9321,N_9020,N_9028);
xnor U9322 (N_9322,N_9047,N_9028);
nor U9323 (N_9323,N_9169,N_9152);
nor U9324 (N_9324,N_9181,N_9107);
and U9325 (N_9325,N_9054,N_9080);
nand U9326 (N_9326,N_9156,N_9117);
nor U9327 (N_9327,N_9123,N_9073);
nor U9328 (N_9328,N_9028,N_9113);
nand U9329 (N_9329,N_9003,N_9023);
xnor U9330 (N_9330,N_9131,N_9003);
nor U9331 (N_9331,N_9193,N_9126);
nand U9332 (N_9332,N_9139,N_9021);
and U9333 (N_9333,N_9154,N_9120);
and U9334 (N_9334,N_9066,N_9076);
xnor U9335 (N_9335,N_9096,N_9055);
or U9336 (N_9336,N_9129,N_9124);
xnor U9337 (N_9337,N_9110,N_9079);
xnor U9338 (N_9338,N_9099,N_9019);
xor U9339 (N_9339,N_9126,N_9060);
nand U9340 (N_9340,N_9092,N_9113);
nor U9341 (N_9341,N_9077,N_9168);
and U9342 (N_9342,N_9145,N_9129);
xor U9343 (N_9343,N_9087,N_9055);
and U9344 (N_9344,N_9174,N_9116);
or U9345 (N_9345,N_9076,N_9170);
and U9346 (N_9346,N_9088,N_9128);
or U9347 (N_9347,N_9096,N_9121);
nor U9348 (N_9348,N_9066,N_9195);
or U9349 (N_9349,N_9181,N_9105);
or U9350 (N_9350,N_9065,N_9168);
or U9351 (N_9351,N_9062,N_9164);
and U9352 (N_9352,N_9132,N_9159);
nand U9353 (N_9353,N_9127,N_9049);
xnor U9354 (N_9354,N_9111,N_9104);
xnor U9355 (N_9355,N_9106,N_9176);
nand U9356 (N_9356,N_9023,N_9198);
nor U9357 (N_9357,N_9005,N_9134);
nor U9358 (N_9358,N_9132,N_9098);
and U9359 (N_9359,N_9036,N_9063);
and U9360 (N_9360,N_9100,N_9058);
or U9361 (N_9361,N_9118,N_9197);
and U9362 (N_9362,N_9058,N_9004);
or U9363 (N_9363,N_9158,N_9046);
nor U9364 (N_9364,N_9198,N_9001);
xnor U9365 (N_9365,N_9120,N_9041);
or U9366 (N_9366,N_9014,N_9143);
or U9367 (N_9367,N_9133,N_9157);
nor U9368 (N_9368,N_9154,N_9014);
xnor U9369 (N_9369,N_9073,N_9012);
xnor U9370 (N_9370,N_9116,N_9070);
nand U9371 (N_9371,N_9111,N_9091);
nor U9372 (N_9372,N_9182,N_9122);
nor U9373 (N_9373,N_9127,N_9073);
or U9374 (N_9374,N_9106,N_9080);
nor U9375 (N_9375,N_9099,N_9058);
or U9376 (N_9376,N_9142,N_9198);
or U9377 (N_9377,N_9160,N_9110);
and U9378 (N_9378,N_9095,N_9173);
nor U9379 (N_9379,N_9180,N_9120);
and U9380 (N_9380,N_9001,N_9151);
and U9381 (N_9381,N_9134,N_9067);
nand U9382 (N_9382,N_9037,N_9056);
nor U9383 (N_9383,N_9087,N_9086);
or U9384 (N_9384,N_9126,N_9089);
nor U9385 (N_9385,N_9098,N_9130);
nor U9386 (N_9386,N_9050,N_9064);
nor U9387 (N_9387,N_9101,N_9137);
and U9388 (N_9388,N_9111,N_9037);
and U9389 (N_9389,N_9044,N_9091);
nor U9390 (N_9390,N_9087,N_9172);
nor U9391 (N_9391,N_9080,N_9038);
or U9392 (N_9392,N_9149,N_9029);
nor U9393 (N_9393,N_9000,N_9145);
and U9394 (N_9394,N_9044,N_9198);
or U9395 (N_9395,N_9007,N_9175);
xor U9396 (N_9396,N_9178,N_9060);
nand U9397 (N_9397,N_9043,N_9094);
or U9398 (N_9398,N_9166,N_9039);
xor U9399 (N_9399,N_9038,N_9060);
or U9400 (N_9400,N_9376,N_9358);
and U9401 (N_9401,N_9309,N_9315);
and U9402 (N_9402,N_9226,N_9232);
and U9403 (N_9403,N_9246,N_9386);
nor U9404 (N_9404,N_9342,N_9330);
and U9405 (N_9405,N_9324,N_9366);
nand U9406 (N_9406,N_9201,N_9258);
or U9407 (N_9407,N_9387,N_9294);
xnor U9408 (N_9408,N_9397,N_9394);
xnor U9409 (N_9409,N_9235,N_9254);
nand U9410 (N_9410,N_9299,N_9250);
and U9411 (N_9411,N_9349,N_9352);
nor U9412 (N_9412,N_9367,N_9273);
nor U9413 (N_9413,N_9283,N_9312);
nor U9414 (N_9414,N_9219,N_9346);
nor U9415 (N_9415,N_9372,N_9248);
nand U9416 (N_9416,N_9302,N_9236);
and U9417 (N_9417,N_9378,N_9337);
or U9418 (N_9418,N_9396,N_9295);
xnor U9419 (N_9419,N_9204,N_9325);
nand U9420 (N_9420,N_9365,N_9284);
nand U9421 (N_9421,N_9213,N_9368);
and U9422 (N_9422,N_9261,N_9275);
and U9423 (N_9423,N_9209,N_9215);
xnor U9424 (N_9424,N_9227,N_9390);
or U9425 (N_9425,N_9357,N_9313);
xnor U9426 (N_9426,N_9267,N_9255);
or U9427 (N_9427,N_9266,N_9286);
nor U9428 (N_9428,N_9289,N_9272);
and U9429 (N_9429,N_9340,N_9208);
xnor U9430 (N_9430,N_9389,N_9280);
or U9431 (N_9431,N_9356,N_9343);
nor U9432 (N_9432,N_9217,N_9382);
nand U9433 (N_9433,N_9228,N_9203);
and U9434 (N_9434,N_9323,N_9224);
xor U9435 (N_9435,N_9344,N_9296);
xnor U9436 (N_9436,N_9355,N_9263);
nand U9437 (N_9437,N_9395,N_9301);
or U9438 (N_9438,N_9300,N_9205);
xor U9439 (N_9439,N_9305,N_9212);
or U9440 (N_9440,N_9316,N_9384);
and U9441 (N_9441,N_9370,N_9265);
xor U9442 (N_9442,N_9334,N_9270);
and U9443 (N_9443,N_9262,N_9335);
nor U9444 (N_9444,N_9223,N_9363);
or U9445 (N_9445,N_9380,N_9233);
xnor U9446 (N_9446,N_9249,N_9242);
nor U9447 (N_9447,N_9285,N_9381);
or U9448 (N_9448,N_9293,N_9359);
xor U9449 (N_9449,N_9225,N_9239);
nand U9450 (N_9450,N_9351,N_9327);
and U9451 (N_9451,N_9276,N_9211);
xor U9452 (N_9452,N_9328,N_9392);
nand U9453 (N_9453,N_9338,N_9256);
xor U9454 (N_9454,N_9383,N_9311);
xnor U9455 (N_9455,N_9206,N_9279);
or U9456 (N_9456,N_9281,N_9398);
or U9457 (N_9457,N_9234,N_9336);
nor U9458 (N_9458,N_9287,N_9310);
xor U9459 (N_9459,N_9391,N_9371);
nand U9460 (N_9460,N_9321,N_9210);
xor U9461 (N_9461,N_9218,N_9216);
and U9462 (N_9462,N_9319,N_9241);
and U9463 (N_9463,N_9220,N_9307);
xnor U9464 (N_9464,N_9345,N_9317);
nand U9465 (N_9465,N_9332,N_9347);
and U9466 (N_9466,N_9229,N_9329);
nand U9467 (N_9467,N_9251,N_9306);
or U9468 (N_9468,N_9354,N_9377);
nand U9469 (N_9469,N_9257,N_9290);
nor U9470 (N_9470,N_9320,N_9399);
or U9471 (N_9471,N_9314,N_9388);
nand U9472 (N_9472,N_9231,N_9348);
xor U9473 (N_9473,N_9341,N_9361);
xor U9474 (N_9474,N_9364,N_9373);
xor U9475 (N_9475,N_9331,N_9339);
or U9476 (N_9476,N_9259,N_9214);
and U9477 (N_9477,N_9202,N_9303);
and U9478 (N_9478,N_9304,N_9369);
and U9479 (N_9479,N_9260,N_9385);
nand U9480 (N_9480,N_9222,N_9238);
and U9481 (N_9481,N_9230,N_9292);
nor U9482 (N_9482,N_9288,N_9221);
and U9483 (N_9483,N_9200,N_9333);
nand U9484 (N_9484,N_9298,N_9297);
xnor U9485 (N_9485,N_9247,N_9264);
xnor U9486 (N_9486,N_9291,N_9393);
nand U9487 (N_9487,N_9326,N_9237);
nand U9488 (N_9488,N_9207,N_9243);
xnor U9489 (N_9489,N_9379,N_9271);
xnor U9490 (N_9490,N_9277,N_9253);
nand U9491 (N_9491,N_9240,N_9374);
or U9492 (N_9492,N_9278,N_9274);
xor U9493 (N_9493,N_9244,N_9353);
and U9494 (N_9494,N_9375,N_9282);
xnor U9495 (N_9495,N_9268,N_9308);
nand U9496 (N_9496,N_9350,N_9269);
nor U9497 (N_9497,N_9322,N_9360);
and U9498 (N_9498,N_9318,N_9245);
and U9499 (N_9499,N_9362,N_9252);
and U9500 (N_9500,N_9282,N_9363);
nand U9501 (N_9501,N_9232,N_9392);
nand U9502 (N_9502,N_9232,N_9220);
nand U9503 (N_9503,N_9363,N_9232);
or U9504 (N_9504,N_9321,N_9362);
and U9505 (N_9505,N_9389,N_9203);
and U9506 (N_9506,N_9209,N_9204);
and U9507 (N_9507,N_9207,N_9202);
nand U9508 (N_9508,N_9277,N_9300);
nor U9509 (N_9509,N_9265,N_9346);
or U9510 (N_9510,N_9219,N_9393);
nand U9511 (N_9511,N_9359,N_9201);
or U9512 (N_9512,N_9381,N_9297);
or U9513 (N_9513,N_9273,N_9302);
and U9514 (N_9514,N_9265,N_9247);
and U9515 (N_9515,N_9309,N_9389);
and U9516 (N_9516,N_9259,N_9322);
and U9517 (N_9517,N_9293,N_9334);
nor U9518 (N_9518,N_9258,N_9202);
and U9519 (N_9519,N_9213,N_9322);
xor U9520 (N_9520,N_9238,N_9293);
and U9521 (N_9521,N_9209,N_9318);
nand U9522 (N_9522,N_9323,N_9218);
and U9523 (N_9523,N_9250,N_9323);
xor U9524 (N_9524,N_9280,N_9298);
nand U9525 (N_9525,N_9355,N_9246);
nor U9526 (N_9526,N_9293,N_9259);
nor U9527 (N_9527,N_9339,N_9343);
xor U9528 (N_9528,N_9261,N_9387);
nor U9529 (N_9529,N_9204,N_9231);
nor U9530 (N_9530,N_9296,N_9387);
nand U9531 (N_9531,N_9354,N_9348);
nor U9532 (N_9532,N_9393,N_9208);
or U9533 (N_9533,N_9284,N_9362);
xor U9534 (N_9534,N_9355,N_9366);
xor U9535 (N_9535,N_9372,N_9322);
nor U9536 (N_9536,N_9359,N_9315);
nor U9537 (N_9537,N_9378,N_9229);
nor U9538 (N_9538,N_9357,N_9321);
nor U9539 (N_9539,N_9370,N_9218);
or U9540 (N_9540,N_9346,N_9284);
or U9541 (N_9541,N_9296,N_9214);
or U9542 (N_9542,N_9379,N_9218);
xor U9543 (N_9543,N_9231,N_9394);
and U9544 (N_9544,N_9323,N_9378);
xnor U9545 (N_9545,N_9301,N_9204);
nand U9546 (N_9546,N_9290,N_9320);
or U9547 (N_9547,N_9253,N_9269);
and U9548 (N_9548,N_9357,N_9392);
nor U9549 (N_9549,N_9277,N_9295);
nor U9550 (N_9550,N_9209,N_9287);
nor U9551 (N_9551,N_9386,N_9363);
and U9552 (N_9552,N_9382,N_9390);
xnor U9553 (N_9553,N_9289,N_9299);
or U9554 (N_9554,N_9265,N_9368);
nor U9555 (N_9555,N_9262,N_9363);
or U9556 (N_9556,N_9316,N_9256);
or U9557 (N_9557,N_9269,N_9255);
nand U9558 (N_9558,N_9348,N_9253);
or U9559 (N_9559,N_9219,N_9358);
nor U9560 (N_9560,N_9294,N_9279);
xnor U9561 (N_9561,N_9364,N_9339);
nand U9562 (N_9562,N_9337,N_9393);
nor U9563 (N_9563,N_9213,N_9239);
nand U9564 (N_9564,N_9211,N_9378);
nand U9565 (N_9565,N_9239,N_9369);
or U9566 (N_9566,N_9281,N_9294);
or U9567 (N_9567,N_9375,N_9293);
nor U9568 (N_9568,N_9281,N_9300);
or U9569 (N_9569,N_9398,N_9222);
and U9570 (N_9570,N_9232,N_9321);
xor U9571 (N_9571,N_9295,N_9370);
nand U9572 (N_9572,N_9237,N_9361);
and U9573 (N_9573,N_9340,N_9317);
nand U9574 (N_9574,N_9315,N_9327);
nand U9575 (N_9575,N_9339,N_9266);
xor U9576 (N_9576,N_9347,N_9338);
or U9577 (N_9577,N_9200,N_9336);
and U9578 (N_9578,N_9233,N_9249);
or U9579 (N_9579,N_9379,N_9340);
and U9580 (N_9580,N_9280,N_9366);
xnor U9581 (N_9581,N_9334,N_9397);
xnor U9582 (N_9582,N_9337,N_9379);
nor U9583 (N_9583,N_9219,N_9308);
and U9584 (N_9584,N_9243,N_9324);
and U9585 (N_9585,N_9303,N_9273);
or U9586 (N_9586,N_9350,N_9291);
xnor U9587 (N_9587,N_9256,N_9301);
nor U9588 (N_9588,N_9325,N_9363);
xor U9589 (N_9589,N_9252,N_9220);
xnor U9590 (N_9590,N_9260,N_9312);
and U9591 (N_9591,N_9335,N_9270);
nand U9592 (N_9592,N_9275,N_9223);
nand U9593 (N_9593,N_9356,N_9257);
or U9594 (N_9594,N_9275,N_9252);
nand U9595 (N_9595,N_9207,N_9270);
xnor U9596 (N_9596,N_9258,N_9311);
nand U9597 (N_9597,N_9336,N_9215);
and U9598 (N_9598,N_9243,N_9395);
nor U9599 (N_9599,N_9213,N_9214);
nand U9600 (N_9600,N_9459,N_9420);
or U9601 (N_9601,N_9467,N_9429);
xor U9602 (N_9602,N_9503,N_9578);
nand U9603 (N_9603,N_9403,N_9589);
xnor U9604 (N_9604,N_9480,N_9411);
xnor U9605 (N_9605,N_9547,N_9434);
nor U9606 (N_9606,N_9495,N_9442);
nor U9607 (N_9607,N_9409,N_9516);
nor U9608 (N_9608,N_9583,N_9494);
nand U9609 (N_9609,N_9458,N_9577);
nand U9610 (N_9610,N_9407,N_9457);
or U9611 (N_9611,N_9533,N_9576);
xnor U9612 (N_9612,N_9437,N_9497);
or U9613 (N_9613,N_9505,N_9594);
nor U9614 (N_9614,N_9562,N_9596);
nor U9615 (N_9615,N_9511,N_9490);
or U9616 (N_9616,N_9502,N_9479);
nor U9617 (N_9617,N_9460,N_9537);
xor U9618 (N_9618,N_9529,N_9572);
nand U9619 (N_9619,N_9451,N_9421);
and U9620 (N_9620,N_9474,N_9462);
nor U9621 (N_9621,N_9419,N_9546);
nor U9622 (N_9622,N_9402,N_9415);
nand U9623 (N_9623,N_9477,N_9426);
and U9624 (N_9624,N_9565,N_9591);
and U9625 (N_9625,N_9581,N_9564);
or U9626 (N_9626,N_9584,N_9585);
and U9627 (N_9627,N_9416,N_9456);
nand U9628 (N_9628,N_9553,N_9555);
and U9629 (N_9629,N_9463,N_9573);
or U9630 (N_9630,N_9549,N_9580);
xnor U9631 (N_9631,N_9515,N_9417);
xnor U9632 (N_9632,N_9520,N_9466);
or U9633 (N_9633,N_9539,N_9544);
nand U9634 (N_9634,N_9513,N_9540);
nor U9635 (N_9635,N_9561,N_9405);
xnor U9636 (N_9636,N_9563,N_9569);
or U9637 (N_9637,N_9512,N_9438);
nand U9638 (N_9638,N_9430,N_9567);
or U9639 (N_9639,N_9439,N_9414);
nor U9640 (N_9640,N_9510,N_9541);
nand U9641 (N_9641,N_9597,N_9550);
or U9642 (N_9642,N_9444,N_9493);
nand U9643 (N_9643,N_9506,N_9508);
or U9644 (N_9644,N_9556,N_9445);
xnor U9645 (N_9645,N_9514,N_9598);
nor U9646 (N_9646,N_9424,N_9518);
nor U9647 (N_9647,N_9436,N_9412);
nor U9648 (N_9648,N_9486,N_9566);
or U9649 (N_9649,N_9453,N_9452);
nor U9650 (N_9650,N_9408,N_9532);
and U9651 (N_9651,N_9473,N_9568);
nand U9652 (N_9652,N_9454,N_9545);
nand U9653 (N_9653,N_9491,N_9446);
or U9654 (N_9654,N_9593,N_9534);
and U9655 (N_9655,N_9588,N_9410);
nor U9656 (N_9656,N_9504,N_9423);
and U9657 (N_9657,N_9482,N_9440);
nor U9658 (N_9658,N_9527,N_9400);
xor U9659 (N_9659,N_9554,N_9575);
nand U9660 (N_9660,N_9425,N_9447);
or U9661 (N_9661,N_9431,N_9464);
xnor U9662 (N_9662,N_9489,N_9485);
nand U9663 (N_9663,N_9579,N_9559);
xnor U9664 (N_9664,N_9468,N_9432);
xnor U9665 (N_9665,N_9465,N_9528);
nand U9666 (N_9666,N_9543,N_9481);
and U9667 (N_9667,N_9449,N_9476);
nor U9668 (N_9668,N_9418,N_9441);
nor U9669 (N_9669,N_9443,N_9492);
nand U9670 (N_9670,N_9524,N_9587);
xor U9671 (N_9671,N_9519,N_9517);
nor U9672 (N_9672,N_9496,N_9570);
or U9673 (N_9673,N_9586,N_9499);
xor U9674 (N_9674,N_9448,N_9590);
nor U9675 (N_9675,N_9557,N_9428);
nand U9676 (N_9676,N_9535,N_9560);
nand U9677 (N_9677,N_9469,N_9475);
or U9678 (N_9678,N_9530,N_9435);
nand U9679 (N_9679,N_9487,N_9536);
or U9680 (N_9680,N_9470,N_9531);
and U9681 (N_9681,N_9522,N_9433);
or U9682 (N_9682,N_9526,N_9472);
nand U9683 (N_9683,N_9542,N_9422);
nor U9684 (N_9684,N_9404,N_9406);
nand U9685 (N_9685,N_9461,N_9484);
nor U9686 (N_9686,N_9551,N_9509);
nor U9687 (N_9687,N_9455,N_9488);
xor U9688 (N_9688,N_9558,N_9401);
nor U9689 (N_9689,N_9582,N_9574);
or U9690 (N_9690,N_9592,N_9450);
xor U9691 (N_9691,N_9548,N_9498);
or U9692 (N_9692,N_9525,N_9521);
nor U9693 (N_9693,N_9500,N_9471);
xnor U9694 (N_9694,N_9538,N_9501);
xor U9695 (N_9695,N_9478,N_9523);
and U9696 (N_9696,N_9427,N_9599);
and U9697 (N_9697,N_9483,N_9552);
nor U9698 (N_9698,N_9595,N_9413);
or U9699 (N_9699,N_9507,N_9571);
or U9700 (N_9700,N_9541,N_9580);
or U9701 (N_9701,N_9436,N_9521);
and U9702 (N_9702,N_9419,N_9486);
nand U9703 (N_9703,N_9486,N_9442);
nand U9704 (N_9704,N_9437,N_9448);
and U9705 (N_9705,N_9453,N_9512);
nand U9706 (N_9706,N_9590,N_9518);
or U9707 (N_9707,N_9547,N_9577);
xor U9708 (N_9708,N_9480,N_9554);
or U9709 (N_9709,N_9594,N_9445);
nor U9710 (N_9710,N_9531,N_9573);
nor U9711 (N_9711,N_9497,N_9402);
nor U9712 (N_9712,N_9549,N_9586);
nor U9713 (N_9713,N_9439,N_9424);
or U9714 (N_9714,N_9498,N_9465);
or U9715 (N_9715,N_9420,N_9554);
nor U9716 (N_9716,N_9427,N_9583);
nand U9717 (N_9717,N_9537,N_9481);
xor U9718 (N_9718,N_9434,N_9463);
xnor U9719 (N_9719,N_9516,N_9541);
or U9720 (N_9720,N_9429,N_9418);
or U9721 (N_9721,N_9500,N_9503);
nor U9722 (N_9722,N_9594,N_9589);
nor U9723 (N_9723,N_9520,N_9562);
nor U9724 (N_9724,N_9470,N_9453);
nor U9725 (N_9725,N_9584,N_9552);
nand U9726 (N_9726,N_9576,N_9451);
nand U9727 (N_9727,N_9506,N_9464);
xor U9728 (N_9728,N_9554,N_9464);
and U9729 (N_9729,N_9475,N_9412);
xnor U9730 (N_9730,N_9465,N_9407);
xor U9731 (N_9731,N_9553,N_9455);
nand U9732 (N_9732,N_9438,N_9434);
xor U9733 (N_9733,N_9538,N_9540);
nand U9734 (N_9734,N_9578,N_9597);
or U9735 (N_9735,N_9468,N_9404);
xor U9736 (N_9736,N_9568,N_9525);
nor U9737 (N_9737,N_9404,N_9580);
or U9738 (N_9738,N_9473,N_9520);
nand U9739 (N_9739,N_9493,N_9516);
or U9740 (N_9740,N_9495,N_9440);
or U9741 (N_9741,N_9493,N_9456);
xor U9742 (N_9742,N_9404,N_9411);
nor U9743 (N_9743,N_9404,N_9444);
xnor U9744 (N_9744,N_9409,N_9462);
or U9745 (N_9745,N_9430,N_9572);
xor U9746 (N_9746,N_9591,N_9574);
nor U9747 (N_9747,N_9508,N_9428);
xor U9748 (N_9748,N_9456,N_9417);
nand U9749 (N_9749,N_9510,N_9434);
or U9750 (N_9750,N_9456,N_9450);
nand U9751 (N_9751,N_9441,N_9577);
and U9752 (N_9752,N_9587,N_9527);
nand U9753 (N_9753,N_9422,N_9531);
nand U9754 (N_9754,N_9402,N_9579);
xor U9755 (N_9755,N_9599,N_9573);
xnor U9756 (N_9756,N_9472,N_9520);
and U9757 (N_9757,N_9547,N_9485);
and U9758 (N_9758,N_9481,N_9521);
nand U9759 (N_9759,N_9498,N_9441);
nor U9760 (N_9760,N_9427,N_9582);
nand U9761 (N_9761,N_9459,N_9520);
nand U9762 (N_9762,N_9560,N_9470);
nand U9763 (N_9763,N_9483,N_9476);
nor U9764 (N_9764,N_9561,N_9473);
nor U9765 (N_9765,N_9559,N_9448);
or U9766 (N_9766,N_9594,N_9559);
nand U9767 (N_9767,N_9401,N_9417);
and U9768 (N_9768,N_9496,N_9443);
and U9769 (N_9769,N_9471,N_9442);
or U9770 (N_9770,N_9587,N_9493);
nand U9771 (N_9771,N_9446,N_9468);
or U9772 (N_9772,N_9475,N_9431);
and U9773 (N_9773,N_9469,N_9493);
nand U9774 (N_9774,N_9568,N_9412);
and U9775 (N_9775,N_9452,N_9560);
nand U9776 (N_9776,N_9571,N_9547);
and U9777 (N_9777,N_9406,N_9440);
or U9778 (N_9778,N_9503,N_9521);
or U9779 (N_9779,N_9471,N_9412);
nor U9780 (N_9780,N_9406,N_9518);
nand U9781 (N_9781,N_9494,N_9414);
nor U9782 (N_9782,N_9571,N_9492);
xor U9783 (N_9783,N_9538,N_9541);
or U9784 (N_9784,N_9562,N_9484);
xor U9785 (N_9785,N_9452,N_9481);
xor U9786 (N_9786,N_9490,N_9556);
and U9787 (N_9787,N_9470,N_9547);
or U9788 (N_9788,N_9451,N_9419);
nor U9789 (N_9789,N_9485,N_9554);
nand U9790 (N_9790,N_9495,N_9422);
xor U9791 (N_9791,N_9458,N_9521);
nand U9792 (N_9792,N_9534,N_9547);
or U9793 (N_9793,N_9484,N_9421);
xnor U9794 (N_9794,N_9592,N_9426);
or U9795 (N_9795,N_9545,N_9522);
nor U9796 (N_9796,N_9426,N_9492);
or U9797 (N_9797,N_9402,N_9575);
or U9798 (N_9798,N_9525,N_9401);
nor U9799 (N_9799,N_9520,N_9485);
and U9800 (N_9800,N_9723,N_9657);
nand U9801 (N_9801,N_9763,N_9786);
nor U9802 (N_9802,N_9677,N_9619);
nor U9803 (N_9803,N_9616,N_9693);
nor U9804 (N_9804,N_9758,N_9714);
or U9805 (N_9805,N_9740,N_9697);
xnor U9806 (N_9806,N_9748,N_9671);
nor U9807 (N_9807,N_9743,N_9759);
and U9808 (N_9808,N_9682,N_9708);
nand U9809 (N_9809,N_9673,N_9711);
or U9810 (N_9810,N_9684,N_9600);
and U9811 (N_9811,N_9615,N_9627);
and U9812 (N_9812,N_9610,N_9744);
xnor U9813 (N_9813,N_9783,N_9674);
nand U9814 (N_9814,N_9655,N_9733);
and U9815 (N_9815,N_9781,N_9672);
xnor U9816 (N_9816,N_9742,N_9643);
nand U9817 (N_9817,N_9730,N_9716);
nor U9818 (N_9818,N_9611,N_9628);
or U9819 (N_9819,N_9698,N_9754);
xor U9820 (N_9820,N_9686,N_9602);
and U9821 (N_9821,N_9727,N_9666);
xnor U9822 (N_9822,N_9683,N_9669);
nor U9823 (N_9823,N_9623,N_9646);
xor U9824 (N_9824,N_9606,N_9788);
nand U9825 (N_9825,N_9654,N_9648);
nor U9826 (N_9826,N_9775,N_9726);
xnor U9827 (N_9827,N_9787,N_9649);
nor U9828 (N_9828,N_9722,N_9713);
nor U9829 (N_9829,N_9629,N_9718);
and U9830 (N_9830,N_9650,N_9706);
nand U9831 (N_9831,N_9753,N_9661);
and U9832 (N_9832,N_9784,N_9729);
xnor U9833 (N_9833,N_9645,N_9685);
nand U9834 (N_9834,N_9792,N_9717);
nor U9835 (N_9835,N_9774,N_9641);
and U9836 (N_9836,N_9769,N_9656);
nor U9837 (N_9837,N_9695,N_9764);
xor U9838 (N_9838,N_9705,N_9622);
xnor U9839 (N_9839,N_9636,N_9620);
nand U9840 (N_9840,N_9724,N_9728);
xor U9841 (N_9841,N_9704,N_9618);
nand U9842 (N_9842,N_9752,N_9687);
or U9843 (N_9843,N_9689,N_9780);
and U9844 (N_9844,N_9731,N_9751);
xnor U9845 (N_9845,N_9710,N_9696);
nand U9846 (N_9846,N_9608,N_9678);
and U9847 (N_9847,N_9789,N_9798);
and U9848 (N_9848,N_9675,N_9624);
xnor U9849 (N_9849,N_9778,N_9761);
and U9850 (N_9850,N_9719,N_9664);
nor U9851 (N_9851,N_9612,N_9692);
nor U9852 (N_9852,N_9614,N_9796);
or U9853 (N_9853,N_9736,N_9663);
nor U9854 (N_9854,N_9756,N_9715);
nand U9855 (N_9855,N_9662,N_9734);
nor U9856 (N_9856,N_9737,N_9735);
nor U9857 (N_9857,N_9691,N_9746);
nand U9858 (N_9858,N_9621,N_9631);
or U9859 (N_9859,N_9762,N_9720);
nand U9860 (N_9860,N_9745,N_9694);
nand U9861 (N_9861,N_9772,N_9630);
nor U9862 (N_9862,N_9676,N_9680);
and U9863 (N_9863,N_9799,N_9760);
nand U9864 (N_9864,N_9603,N_9604);
nand U9865 (N_9865,N_9770,N_9750);
nor U9866 (N_9866,N_9709,N_9681);
xor U9867 (N_9867,N_9773,N_9639);
nor U9868 (N_9868,N_9640,N_9642);
and U9869 (N_9869,N_9647,N_9660);
nor U9870 (N_9870,N_9679,N_9749);
and U9871 (N_9871,N_9757,N_9794);
nand U9872 (N_9872,N_9795,N_9791);
nand U9873 (N_9873,N_9651,N_9617);
nor U9874 (N_9874,N_9703,N_9644);
or U9875 (N_9875,N_9702,N_9785);
nor U9876 (N_9876,N_9632,N_9739);
xnor U9877 (N_9877,N_9605,N_9699);
xor U9878 (N_9878,N_9667,N_9653);
and U9879 (N_9879,N_9793,N_9637);
nand U9880 (N_9880,N_9765,N_9609);
or U9881 (N_9881,N_9652,N_9707);
xnor U9882 (N_9882,N_9638,N_9601);
nor U9883 (N_9883,N_9782,N_9670);
xor U9884 (N_9884,N_9790,N_9658);
nand U9885 (N_9885,N_9777,N_9607);
nand U9886 (N_9886,N_9797,N_9712);
or U9887 (N_9887,N_9625,N_9688);
and U9888 (N_9888,N_9766,N_9665);
nand U9889 (N_9889,N_9725,N_9767);
nor U9890 (N_9890,N_9721,N_9741);
nand U9891 (N_9891,N_9613,N_9768);
or U9892 (N_9892,N_9700,N_9771);
and U9893 (N_9893,N_9659,N_9779);
nor U9894 (N_9894,N_9668,N_9738);
or U9895 (N_9895,N_9732,N_9634);
nand U9896 (N_9896,N_9626,N_9690);
or U9897 (N_9897,N_9776,N_9633);
or U9898 (N_9898,N_9635,N_9701);
nor U9899 (N_9899,N_9755,N_9747);
nor U9900 (N_9900,N_9686,N_9717);
xnor U9901 (N_9901,N_9671,N_9689);
or U9902 (N_9902,N_9657,N_9634);
and U9903 (N_9903,N_9740,N_9656);
or U9904 (N_9904,N_9650,N_9636);
nand U9905 (N_9905,N_9768,N_9734);
nor U9906 (N_9906,N_9678,N_9756);
or U9907 (N_9907,N_9613,N_9724);
and U9908 (N_9908,N_9740,N_9659);
xor U9909 (N_9909,N_9674,N_9616);
xnor U9910 (N_9910,N_9625,N_9716);
nor U9911 (N_9911,N_9612,N_9786);
nand U9912 (N_9912,N_9681,N_9631);
nor U9913 (N_9913,N_9708,N_9647);
nand U9914 (N_9914,N_9701,N_9611);
nand U9915 (N_9915,N_9641,N_9792);
and U9916 (N_9916,N_9667,N_9779);
xnor U9917 (N_9917,N_9685,N_9774);
nand U9918 (N_9918,N_9612,N_9690);
nand U9919 (N_9919,N_9748,N_9606);
nor U9920 (N_9920,N_9638,N_9714);
and U9921 (N_9921,N_9614,N_9639);
xor U9922 (N_9922,N_9708,N_9641);
xor U9923 (N_9923,N_9739,N_9631);
xor U9924 (N_9924,N_9792,N_9653);
or U9925 (N_9925,N_9641,N_9685);
and U9926 (N_9926,N_9762,N_9649);
nand U9927 (N_9927,N_9701,N_9784);
or U9928 (N_9928,N_9603,N_9798);
xor U9929 (N_9929,N_9706,N_9705);
nor U9930 (N_9930,N_9788,N_9683);
xnor U9931 (N_9931,N_9701,N_9642);
or U9932 (N_9932,N_9657,N_9769);
and U9933 (N_9933,N_9689,N_9799);
nor U9934 (N_9934,N_9741,N_9618);
nand U9935 (N_9935,N_9654,N_9687);
and U9936 (N_9936,N_9721,N_9706);
nor U9937 (N_9937,N_9740,N_9683);
or U9938 (N_9938,N_9630,N_9771);
or U9939 (N_9939,N_9649,N_9777);
nor U9940 (N_9940,N_9738,N_9732);
nor U9941 (N_9941,N_9775,N_9790);
and U9942 (N_9942,N_9629,N_9655);
xor U9943 (N_9943,N_9792,N_9659);
nand U9944 (N_9944,N_9651,N_9748);
nand U9945 (N_9945,N_9777,N_9720);
and U9946 (N_9946,N_9611,N_9732);
nor U9947 (N_9947,N_9707,N_9628);
nand U9948 (N_9948,N_9781,N_9713);
nor U9949 (N_9949,N_9638,N_9692);
nor U9950 (N_9950,N_9796,N_9771);
and U9951 (N_9951,N_9649,N_9680);
and U9952 (N_9952,N_9619,N_9797);
nand U9953 (N_9953,N_9675,N_9606);
or U9954 (N_9954,N_9661,N_9791);
xor U9955 (N_9955,N_9746,N_9723);
or U9956 (N_9956,N_9721,N_9758);
and U9957 (N_9957,N_9707,N_9656);
and U9958 (N_9958,N_9746,N_9766);
xnor U9959 (N_9959,N_9744,N_9728);
and U9960 (N_9960,N_9751,N_9756);
nor U9961 (N_9961,N_9788,N_9740);
nor U9962 (N_9962,N_9706,N_9730);
nor U9963 (N_9963,N_9696,N_9655);
xor U9964 (N_9964,N_9734,N_9674);
and U9965 (N_9965,N_9701,N_9751);
nor U9966 (N_9966,N_9709,N_9794);
or U9967 (N_9967,N_9780,N_9716);
nor U9968 (N_9968,N_9786,N_9634);
nor U9969 (N_9969,N_9674,N_9646);
nor U9970 (N_9970,N_9681,N_9785);
xor U9971 (N_9971,N_9743,N_9690);
or U9972 (N_9972,N_9622,N_9652);
or U9973 (N_9973,N_9792,N_9795);
nor U9974 (N_9974,N_9631,N_9689);
and U9975 (N_9975,N_9654,N_9665);
or U9976 (N_9976,N_9691,N_9611);
nand U9977 (N_9977,N_9796,N_9648);
nand U9978 (N_9978,N_9780,N_9792);
nand U9979 (N_9979,N_9662,N_9655);
xor U9980 (N_9980,N_9669,N_9751);
and U9981 (N_9981,N_9658,N_9723);
nor U9982 (N_9982,N_9712,N_9650);
xor U9983 (N_9983,N_9667,N_9780);
xnor U9984 (N_9984,N_9616,N_9704);
xnor U9985 (N_9985,N_9730,N_9755);
xor U9986 (N_9986,N_9773,N_9795);
and U9987 (N_9987,N_9630,N_9640);
and U9988 (N_9988,N_9753,N_9630);
nor U9989 (N_9989,N_9623,N_9752);
nand U9990 (N_9990,N_9705,N_9730);
and U9991 (N_9991,N_9684,N_9754);
xnor U9992 (N_9992,N_9605,N_9647);
and U9993 (N_9993,N_9622,N_9749);
nor U9994 (N_9994,N_9714,N_9717);
xnor U9995 (N_9995,N_9783,N_9606);
and U9996 (N_9996,N_9659,N_9688);
nor U9997 (N_9997,N_9630,N_9768);
nand U9998 (N_9998,N_9758,N_9717);
xor U9999 (N_9999,N_9716,N_9704);
or U10000 (N_10000,N_9878,N_9948);
and U10001 (N_10001,N_9831,N_9992);
xor U10002 (N_10002,N_9898,N_9904);
nand U10003 (N_10003,N_9834,N_9850);
xor U10004 (N_10004,N_9931,N_9823);
and U10005 (N_10005,N_9891,N_9937);
and U10006 (N_10006,N_9844,N_9859);
nor U10007 (N_10007,N_9828,N_9856);
and U10008 (N_10008,N_9887,N_9955);
nor U10009 (N_10009,N_9886,N_9813);
nor U10010 (N_10010,N_9996,N_9968);
nand U10011 (N_10011,N_9936,N_9854);
nand U10012 (N_10012,N_9929,N_9991);
and U10013 (N_10013,N_9877,N_9910);
xor U10014 (N_10014,N_9956,N_9922);
or U10015 (N_10015,N_9837,N_9868);
nor U10016 (N_10016,N_9804,N_9880);
nor U10017 (N_10017,N_9918,N_9864);
nand U10018 (N_10018,N_9935,N_9920);
nand U10019 (N_10019,N_9836,N_9940);
and U10020 (N_10020,N_9999,N_9954);
or U10021 (N_10021,N_9815,N_9913);
nor U10022 (N_10022,N_9841,N_9966);
xnor U10023 (N_10023,N_9874,N_9973);
and U10024 (N_10024,N_9852,N_9958);
nor U10025 (N_10025,N_9811,N_9893);
and U10026 (N_10026,N_9847,N_9860);
and U10027 (N_10027,N_9826,N_9977);
or U10028 (N_10028,N_9916,N_9986);
or U10029 (N_10029,N_9812,N_9923);
or U10030 (N_10030,N_9978,N_9981);
and U10031 (N_10031,N_9928,N_9907);
or U10032 (N_10032,N_9985,N_9930);
nand U10033 (N_10033,N_9901,N_9875);
and U10034 (N_10034,N_9820,N_9855);
and U10035 (N_10035,N_9803,N_9863);
nor U10036 (N_10036,N_9818,N_9833);
nor U10037 (N_10037,N_9805,N_9869);
xnor U10038 (N_10038,N_9896,N_9962);
nor U10039 (N_10039,N_9848,N_9824);
or U10040 (N_10040,N_9881,N_9885);
nand U10041 (N_10041,N_9957,N_9870);
and U10042 (N_10042,N_9861,N_9819);
nor U10043 (N_10043,N_9921,N_9959);
and U10044 (N_10044,N_9932,N_9899);
xnor U10045 (N_10045,N_9865,N_9914);
nor U10046 (N_10046,N_9909,N_9845);
or U10047 (N_10047,N_9912,N_9942);
nor U10048 (N_10048,N_9822,N_9843);
nor U10049 (N_10049,N_9884,N_9984);
or U10050 (N_10050,N_9969,N_9998);
or U10051 (N_10051,N_9926,N_9933);
or U10052 (N_10052,N_9924,N_9816);
xnor U10053 (N_10053,N_9989,N_9943);
nor U10054 (N_10054,N_9947,N_9892);
and U10055 (N_10055,N_9906,N_9801);
or U10056 (N_10056,N_9853,N_9876);
and U10057 (N_10057,N_9849,N_9951);
or U10058 (N_10058,N_9953,N_9964);
and U10059 (N_10059,N_9990,N_9939);
or U10060 (N_10060,N_9871,N_9825);
and U10061 (N_10061,N_9872,N_9975);
xnor U10062 (N_10062,N_9900,N_9915);
nand U10063 (N_10063,N_9846,N_9817);
xor U10064 (N_10064,N_9895,N_9919);
and U10065 (N_10065,N_9889,N_9808);
and U10066 (N_10066,N_9821,N_9945);
or U10067 (N_10067,N_9938,N_9961);
nand U10068 (N_10068,N_9888,N_9806);
xor U10069 (N_10069,N_9979,N_9829);
nor U10070 (N_10070,N_9995,N_9967);
nand U10071 (N_10071,N_9927,N_9827);
nand U10072 (N_10072,N_9832,N_9840);
or U10073 (N_10073,N_9988,N_9835);
nor U10074 (N_10074,N_9862,N_9934);
nand U10075 (N_10075,N_9987,N_9842);
xor U10076 (N_10076,N_9903,N_9949);
or U10077 (N_10077,N_9946,N_9917);
nand U10078 (N_10078,N_9976,N_9897);
and U10079 (N_10079,N_9965,N_9950);
and U10080 (N_10080,N_9980,N_9857);
or U10081 (N_10081,N_9866,N_9858);
nor U10082 (N_10082,N_9807,N_9944);
xor U10083 (N_10083,N_9941,N_9802);
nor U10084 (N_10084,N_9963,N_9993);
and U10085 (N_10085,N_9960,N_9970);
and U10086 (N_10086,N_9971,N_9982);
nor U10087 (N_10087,N_9908,N_9873);
nand U10088 (N_10088,N_9890,N_9879);
nor U10089 (N_10089,N_9905,N_9882);
nor U10090 (N_10090,N_9810,N_9838);
or U10091 (N_10091,N_9997,N_9809);
nor U10092 (N_10092,N_9851,N_9839);
nor U10093 (N_10093,N_9883,N_9983);
nor U10094 (N_10094,N_9972,N_9994);
nor U10095 (N_10095,N_9814,N_9800);
xnor U10096 (N_10096,N_9925,N_9830);
or U10097 (N_10097,N_9952,N_9974);
xor U10098 (N_10098,N_9894,N_9911);
nand U10099 (N_10099,N_9902,N_9867);
xnor U10100 (N_10100,N_9849,N_9818);
nand U10101 (N_10101,N_9946,N_9848);
xnor U10102 (N_10102,N_9815,N_9801);
or U10103 (N_10103,N_9936,N_9939);
xnor U10104 (N_10104,N_9902,N_9811);
nor U10105 (N_10105,N_9848,N_9852);
xor U10106 (N_10106,N_9948,N_9928);
nand U10107 (N_10107,N_9863,N_9921);
nor U10108 (N_10108,N_9908,N_9843);
xor U10109 (N_10109,N_9907,N_9961);
nand U10110 (N_10110,N_9811,N_9942);
nor U10111 (N_10111,N_9886,N_9857);
or U10112 (N_10112,N_9877,N_9878);
xnor U10113 (N_10113,N_9827,N_9940);
xnor U10114 (N_10114,N_9848,N_9923);
and U10115 (N_10115,N_9895,N_9804);
or U10116 (N_10116,N_9940,N_9838);
nor U10117 (N_10117,N_9873,N_9879);
nor U10118 (N_10118,N_9907,N_9962);
nand U10119 (N_10119,N_9942,N_9872);
nor U10120 (N_10120,N_9891,N_9838);
xor U10121 (N_10121,N_9802,N_9990);
or U10122 (N_10122,N_9818,N_9943);
xor U10123 (N_10123,N_9896,N_9800);
nor U10124 (N_10124,N_9815,N_9969);
nor U10125 (N_10125,N_9970,N_9984);
nand U10126 (N_10126,N_9977,N_9939);
nor U10127 (N_10127,N_9965,N_9910);
nand U10128 (N_10128,N_9936,N_9886);
or U10129 (N_10129,N_9946,N_9949);
or U10130 (N_10130,N_9892,N_9926);
or U10131 (N_10131,N_9862,N_9930);
and U10132 (N_10132,N_9813,N_9838);
nor U10133 (N_10133,N_9874,N_9841);
nand U10134 (N_10134,N_9891,N_9870);
nor U10135 (N_10135,N_9839,N_9931);
and U10136 (N_10136,N_9885,N_9973);
nand U10137 (N_10137,N_9877,N_9977);
nor U10138 (N_10138,N_9878,N_9828);
or U10139 (N_10139,N_9988,N_9974);
or U10140 (N_10140,N_9828,N_9844);
xnor U10141 (N_10141,N_9843,N_9943);
xnor U10142 (N_10142,N_9851,N_9823);
and U10143 (N_10143,N_9843,N_9825);
nor U10144 (N_10144,N_9927,N_9845);
nor U10145 (N_10145,N_9900,N_9827);
or U10146 (N_10146,N_9846,N_9878);
or U10147 (N_10147,N_9849,N_9979);
nand U10148 (N_10148,N_9970,N_9910);
nor U10149 (N_10149,N_9979,N_9957);
nand U10150 (N_10150,N_9956,N_9839);
nand U10151 (N_10151,N_9873,N_9961);
or U10152 (N_10152,N_9813,N_9979);
nand U10153 (N_10153,N_9805,N_9823);
xnor U10154 (N_10154,N_9891,N_9999);
or U10155 (N_10155,N_9872,N_9844);
and U10156 (N_10156,N_9810,N_9801);
nor U10157 (N_10157,N_9865,N_9964);
nor U10158 (N_10158,N_9886,N_9883);
nand U10159 (N_10159,N_9954,N_9989);
nor U10160 (N_10160,N_9836,N_9902);
nand U10161 (N_10161,N_9953,N_9880);
and U10162 (N_10162,N_9984,N_9831);
and U10163 (N_10163,N_9940,N_9935);
or U10164 (N_10164,N_9934,N_9956);
nor U10165 (N_10165,N_9849,N_9966);
nand U10166 (N_10166,N_9951,N_9981);
or U10167 (N_10167,N_9972,N_9954);
or U10168 (N_10168,N_9812,N_9924);
nor U10169 (N_10169,N_9851,N_9965);
xor U10170 (N_10170,N_9873,N_9904);
nor U10171 (N_10171,N_9852,N_9956);
xor U10172 (N_10172,N_9874,N_9963);
and U10173 (N_10173,N_9816,N_9913);
nand U10174 (N_10174,N_9881,N_9969);
or U10175 (N_10175,N_9937,N_9856);
and U10176 (N_10176,N_9803,N_9909);
nor U10177 (N_10177,N_9915,N_9928);
and U10178 (N_10178,N_9807,N_9947);
and U10179 (N_10179,N_9905,N_9945);
or U10180 (N_10180,N_9939,N_9805);
and U10181 (N_10181,N_9994,N_9999);
xnor U10182 (N_10182,N_9986,N_9993);
nand U10183 (N_10183,N_9995,N_9890);
xor U10184 (N_10184,N_9827,N_9976);
xor U10185 (N_10185,N_9863,N_9830);
nor U10186 (N_10186,N_9993,N_9887);
nand U10187 (N_10187,N_9813,N_9959);
and U10188 (N_10188,N_9990,N_9916);
nand U10189 (N_10189,N_9846,N_9887);
xnor U10190 (N_10190,N_9944,N_9875);
xor U10191 (N_10191,N_9954,N_9979);
and U10192 (N_10192,N_9818,N_9933);
or U10193 (N_10193,N_9927,N_9960);
nand U10194 (N_10194,N_9895,N_9853);
and U10195 (N_10195,N_9845,N_9837);
and U10196 (N_10196,N_9940,N_9823);
xnor U10197 (N_10197,N_9834,N_9857);
or U10198 (N_10198,N_9891,N_9878);
and U10199 (N_10199,N_9969,N_9812);
or U10200 (N_10200,N_10060,N_10146);
and U10201 (N_10201,N_10173,N_10107);
and U10202 (N_10202,N_10027,N_10064);
xnor U10203 (N_10203,N_10048,N_10078);
and U10204 (N_10204,N_10136,N_10114);
nor U10205 (N_10205,N_10163,N_10036);
or U10206 (N_10206,N_10162,N_10089);
nand U10207 (N_10207,N_10132,N_10122);
xor U10208 (N_10208,N_10196,N_10123);
nand U10209 (N_10209,N_10033,N_10138);
or U10210 (N_10210,N_10002,N_10135);
nand U10211 (N_10211,N_10096,N_10017);
xor U10212 (N_10212,N_10149,N_10130);
xnor U10213 (N_10213,N_10056,N_10053);
xnor U10214 (N_10214,N_10043,N_10026);
xor U10215 (N_10215,N_10194,N_10145);
or U10216 (N_10216,N_10186,N_10118);
nor U10217 (N_10217,N_10023,N_10137);
nand U10218 (N_10218,N_10192,N_10021);
nor U10219 (N_10219,N_10166,N_10083);
and U10220 (N_10220,N_10158,N_10030);
xnor U10221 (N_10221,N_10087,N_10115);
nor U10222 (N_10222,N_10046,N_10108);
nor U10223 (N_10223,N_10010,N_10032);
or U10224 (N_10224,N_10045,N_10151);
or U10225 (N_10225,N_10024,N_10015);
nor U10226 (N_10226,N_10003,N_10019);
and U10227 (N_10227,N_10116,N_10040);
or U10228 (N_10228,N_10093,N_10117);
xor U10229 (N_10229,N_10148,N_10172);
or U10230 (N_10230,N_10178,N_10041);
nand U10231 (N_10231,N_10066,N_10126);
or U10232 (N_10232,N_10052,N_10165);
nor U10233 (N_10233,N_10081,N_10020);
nor U10234 (N_10234,N_10014,N_10197);
xor U10235 (N_10235,N_10198,N_10098);
and U10236 (N_10236,N_10125,N_10062);
xor U10237 (N_10237,N_10028,N_10049);
or U10238 (N_10238,N_10059,N_10067);
nor U10239 (N_10239,N_10101,N_10057);
nand U10240 (N_10240,N_10072,N_10119);
or U10241 (N_10241,N_10000,N_10035);
xor U10242 (N_10242,N_10073,N_10168);
nor U10243 (N_10243,N_10169,N_10183);
and U10244 (N_10244,N_10063,N_10140);
and U10245 (N_10245,N_10167,N_10009);
and U10246 (N_10246,N_10055,N_10004);
nor U10247 (N_10247,N_10187,N_10179);
nand U10248 (N_10248,N_10005,N_10121);
or U10249 (N_10249,N_10124,N_10171);
nor U10250 (N_10250,N_10180,N_10177);
nor U10251 (N_10251,N_10037,N_10071);
or U10252 (N_10252,N_10085,N_10088);
or U10253 (N_10253,N_10007,N_10082);
or U10254 (N_10254,N_10157,N_10142);
or U10255 (N_10255,N_10141,N_10022);
nand U10256 (N_10256,N_10075,N_10025);
and U10257 (N_10257,N_10099,N_10133);
xnor U10258 (N_10258,N_10008,N_10068);
or U10259 (N_10259,N_10012,N_10150);
xnor U10260 (N_10260,N_10013,N_10164);
and U10261 (N_10261,N_10170,N_10105);
or U10262 (N_10262,N_10160,N_10065);
and U10263 (N_10263,N_10079,N_10104);
and U10264 (N_10264,N_10070,N_10190);
or U10265 (N_10265,N_10016,N_10097);
xor U10266 (N_10266,N_10129,N_10143);
nand U10267 (N_10267,N_10039,N_10018);
or U10268 (N_10268,N_10131,N_10086);
and U10269 (N_10269,N_10011,N_10175);
and U10270 (N_10270,N_10113,N_10161);
nor U10271 (N_10271,N_10184,N_10195);
nand U10272 (N_10272,N_10061,N_10102);
xor U10273 (N_10273,N_10069,N_10159);
xor U10274 (N_10274,N_10174,N_10006);
and U10275 (N_10275,N_10127,N_10154);
and U10276 (N_10276,N_10090,N_10095);
and U10277 (N_10277,N_10139,N_10029);
xnor U10278 (N_10278,N_10176,N_10074);
and U10279 (N_10279,N_10189,N_10054);
xor U10280 (N_10280,N_10038,N_10134);
or U10281 (N_10281,N_10120,N_10084);
nor U10282 (N_10282,N_10076,N_10044);
xor U10283 (N_10283,N_10153,N_10047);
nor U10284 (N_10284,N_10128,N_10185);
or U10285 (N_10285,N_10077,N_10144);
and U10286 (N_10286,N_10034,N_10103);
xor U10287 (N_10287,N_10188,N_10091);
xnor U10288 (N_10288,N_10109,N_10080);
or U10289 (N_10289,N_10182,N_10191);
and U10290 (N_10290,N_10051,N_10199);
xnor U10291 (N_10291,N_10155,N_10001);
or U10292 (N_10292,N_10110,N_10181);
and U10293 (N_10293,N_10156,N_10152);
xnor U10294 (N_10294,N_10094,N_10112);
xnor U10295 (N_10295,N_10100,N_10042);
or U10296 (N_10296,N_10147,N_10050);
and U10297 (N_10297,N_10106,N_10111);
or U10298 (N_10298,N_10058,N_10031);
and U10299 (N_10299,N_10092,N_10193);
and U10300 (N_10300,N_10122,N_10151);
and U10301 (N_10301,N_10083,N_10181);
or U10302 (N_10302,N_10124,N_10079);
nand U10303 (N_10303,N_10064,N_10029);
xnor U10304 (N_10304,N_10186,N_10173);
or U10305 (N_10305,N_10129,N_10079);
nand U10306 (N_10306,N_10198,N_10074);
or U10307 (N_10307,N_10052,N_10039);
nand U10308 (N_10308,N_10175,N_10191);
xor U10309 (N_10309,N_10055,N_10001);
nand U10310 (N_10310,N_10187,N_10063);
or U10311 (N_10311,N_10194,N_10009);
xnor U10312 (N_10312,N_10055,N_10030);
xnor U10313 (N_10313,N_10034,N_10080);
xor U10314 (N_10314,N_10038,N_10055);
nand U10315 (N_10315,N_10039,N_10138);
nor U10316 (N_10316,N_10063,N_10065);
and U10317 (N_10317,N_10173,N_10160);
nor U10318 (N_10318,N_10168,N_10031);
or U10319 (N_10319,N_10192,N_10072);
xnor U10320 (N_10320,N_10168,N_10003);
nor U10321 (N_10321,N_10086,N_10097);
xnor U10322 (N_10322,N_10043,N_10046);
and U10323 (N_10323,N_10089,N_10166);
and U10324 (N_10324,N_10122,N_10044);
or U10325 (N_10325,N_10193,N_10051);
nor U10326 (N_10326,N_10191,N_10133);
xnor U10327 (N_10327,N_10085,N_10017);
nor U10328 (N_10328,N_10087,N_10159);
xor U10329 (N_10329,N_10168,N_10177);
and U10330 (N_10330,N_10087,N_10022);
nor U10331 (N_10331,N_10123,N_10195);
or U10332 (N_10332,N_10047,N_10090);
nor U10333 (N_10333,N_10006,N_10199);
xor U10334 (N_10334,N_10053,N_10129);
nand U10335 (N_10335,N_10114,N_10085);
xnor U10336 (N_10336,N_10067,N_10002);
nor U10337 (N_10337,N_10054,N_10073);
or U10338 (N_10338,N_10180,N_10189);
nor U10339 (N_10339,N_10190,N_10136);
nand U10340 (N_10340,N_10009,N_10163);
nor U10341 (N_10341,N_10078,N_10186);
nor U10342 (N_10342,N_10032,N_10118);
and U10343 (N_10343,N_10049,N_10001);
xor U10344 (N_10344,N_10091,N_10174);
nor U10345 (N_10345,N_10191,N_10072);
xor U10346 (N_10346,N_10178,N_10056);
and U10347 (N_10347,N_10123,N_10011);
or U10348 (N_10348,N_10152,N_10194);
and U10349 (N_10349,N_10141,N_10180);
nand U10350 (N_10350,N_10168,N_10035);
nor U10351 (N_10351,N_10082,N_10018);
nor U10352 (N_10352,N_10061,N_10138);
nor U10353 (N_10353,N_10107,N_10017);
nor U10354 (N_10354,N_10152,N_10024);
nor U10355 (N_10355,N_10029,N_10021);
and U10356 (N_10356,N_10154,N_10026);
xor U10357 (N_10357,N_10160,N_10198);
xor U10358 (N_10358,N_10149,N_10020);
and U10359 (N_10359,N_10047,N_10026);
nand U10360 (N_10360,N_10175,N_10127);
xor U10361 (N_10361,N_10074,N_10075);
nand U10362 (N_10362,N_10037,N_10026);
and U10363 (N_10363,N_10031,N_10196);
xnor U10364 (N_10364,N_10161,N_10080);
xnor U10365 (N_10365,N_10104,N_10147);
xor U10366 (N_10366,N_10169,N_10086);
xnor U10367 (N_10367,N_10138,N_10136);
or U10368 (N_10368,N_10138,N_10128);
nor U10369 (N_10369,N_10072,N_10089);
and U10370 (N_10370,N_10025,N_10128);
and U10371 (N_10371,N_10145,N_10106);
xnor U10372 (N_10372,N_10044,N_10104);
and U10373 (N_10373,N_10061,N_10110);
nand U10374 (N_10374,N_10076,N_10196);
nand U10375 (N_10375,N_10182,N_10164);
and U10376 (N_10376,N_10032,N_10042);
nor U10377 (N_10377,N_10006,N_10197);
xnor U10378 (N_10378,N_10068,N_10019);
xnor U10379 (N_10379,N_10060,N_10105);
xnor U10380 (N_10380,N_10061,N_10127);
or U10381 (N_10381,N_10069,N_10002);
or U10382 (N_10382,N_10036,N_10164);
and U10383 (N_10383,N_10152,N_10071);
nor U10384 (N_10384,N_10087,N_10168);
and U10385 (N_10385,N_10029,N_10057);
nor U10386 (N_10386,N_10135,N_10073);
or U10387 (N_10387,N_10128,N_10196);
or U10388 (N_10388,N_10154,N_10077);
xnor U10389 (N_10389,N_10074,N_10013);
or U10390 (N_10390,N_10067,N_10091);
nor U10391 (N_10391,N_10071,N_10019);
or U10392 (N_10392,N_10186,N_10000);
nor U10393 (N_10393,N_10189,N_10153);
and U10394 (N_10394,N_10163,N_10080);
nor U10395 (N_10395,N_10052,N_10057);
or U10396 (N_10396,N_10038,N_10045);
nand U10397 (N_10397,N_10018,N_10139);
xnor U10398 (N_10398,N_10025,N_10023);
xnor U10399 (N_10399,N_10018,N_10074);
xnor U10400 (N_10400,N_10209,N_10308);
xnor U10401 (N_10401,N_10398,N_10325);
and U10402 (N_10402,N_10371,N_10377);
xnor U10403 (N_10403,N_10284,N_10347);
nor U10404 (N_10404,N_10217,N_10262);
nand U10405 (N_10405,N_10296,N_10357);
or U10406 (N_10406,N_10240,N_10206);
nor U10407 (N_10407,N_10245,N_10310);
nor U10408 (N_10408,N_10250,N_10231);
or U10409 (N_10409,N_10225,N_10266);
and U10410 (N_10410,N_10214,N_10312);
xor U10411 (N_10411,N_10317,N_10280);
nand U10412 (N_10412,N_10211,N_10331);
nor U10413 (N_10413,N_10332,N_10324);
and U10414 (N_10414,N_10311,N_10239);
or U10415 (N_10415,N_10374,N_10322);
xnor U10416 (N_10416,N_10323,N_10368);
nor U10417 (N_10417,N_10227,N_10259);
nand U10418 (N_10418,N_10335,N_10223);
xor U10419 (N_10419,N_10226,N_10346);
xnor U10420 (N_10420,N_10359,N_10285);
nand U10421 (N_10421,N_10229,N_10261);
and U10422 (N_10422,N_10307,N_10385);
and U10423 (N_10423,N_10265,N_10330);
nand U10424 (N_10424,N_10337,N_10329);
nand U10425 (N_10425,N_10276,N_10349);
nand U10426 (N_10426,N_10201,N_10222);
nor U10427 (N_10427,N_10388,N_10339);
xor U10428 (N_10428,N_10275,N_10355);
or U10429 (N_10429,N_10288,N_10313);
or U10430 (N_10430,N_10294,N_10251);
or U10431 (N_10431,N_10302,N_10375);
or U10432 (N_10432,N_10356,N_10394);
nor U10433 (N_10433,N_10381,N_10309);
nor U10434 (N_10434,N_10213,N_10242);
or U10435 (N_10435,N_10272,N_10352);
or U10436 (N_10436,N_10334,N_10342);
or U10437 (N_10437,N_10292,N_10344);
nand U10438 (N_10438,N_10220,N_10278);
nand U10439 (N_10439,N_10348,N_10293);
nor U10440 (N_10440,N_10271,N_10380);
nand U10441 (N_10441,N_10301,N_10267);
nor U10442 (N_10442,N_10389,N_10345);
nand U10443 (N_10443,N_10364,N_10353);
and U10444 (N_10444,N_10274,N_10290);
and U10445 (N_10445,N_10260,N_10319);
xnor U10446 (N_10446,N_10306,N_10314);
nor U10447 (N_10447,N_10338,N_10282);
or U10448 (N_10448,N_10383,N_10295);
and U10449 (N_10449,N_10254,N_10249);
nor U10450 (N_10450,N_10237,N_10273);
xnor U10451 (N_10451,N_10246,N_10283);
or U10452 (N_10452,N_10287,N_10263);
nor U10453 (N_10453,N_10219,N_10256);
nor U10454 (N_10454,N_10304,N_10387);
nand U10455 (N_10455,N_10233,N_10247);
or U10456 (N_10456,N_10243,N_10315);
nand U10457 (N_10457,N_10361,N_10351);
nor U10458 (N_10458,N_10257,N_10396);
nand U10459 (N_10459,N_10269,N_10232);
nand U10460 (N_10460,N_10203,N_10221);
nor U10461 (N_10461,N_10224,N_10299);
nor U10462 (N_10462,N_10321,N_10391);
and U10463 (N_10463,N_10297,N_10370);
xor U10464 (N_10464,N_10358,N_10390);
nor U10465 (N_10465,N_10316,N_10258);
and U10466 (N_10466,N_10270,N_10363);
and U10467 (N_10467,N_10382,N_10320);
or U10468 (N_10468,N_10204,N_10212);
xnor U10469 (N_10469,N_10255,N_10291);
or U10470 (N_10470,N_10379,N_10215);
nor U10471 (N_10471,N_10367,N_10289);
or U10472 (N_10472,N_10340,N_10399);
or U10473 (N_10473,N_10241,N_10360);
or U10474 (N_10474,N_10298,N_10264);
nand U10475 (N_10475,N_10362,N_10397);
nand U10476 (N_10476,N_10328,N_10218);
xor U10477 (N_10477,N_10279,N_10210);
or U10478 (N_10478,N_10392,N_10286);
or U10479 (N_10479,N_10318,N_10253);
nand U10480 (N_10480,N_10277,N_10234);
nor U10481 (N_10481,N_10305,N_10235);
nand U10482 (N_10482,N_10200,N_10216);
or U10483 (N_10483,N_10207,N_10372);
or U10484 (N_10484,N_10393,N_10303);
xor U10485 (N_10485,N_10350,N_10244);
xor U10486 (N_10486,N_10327,N_10384);
xnor U10487 (N_10487,N_10366,N_10230);
and U10488 (N_10488,N_10268,N_10365);
and U10489 (N_10489,N_10373,N_10228);
nand U10490 (N_10490,N_10341,N_10252);
nor U10491 (N_10491,N_10202,N_10208);
and U10492 (N_10492,N_10238,N_10378);
nand U10493 (N_10493,N_10354,N_10386);
xor U10494 (N_10494,N_10333,N_10205);
or U10495 (N_10495,N_10369,N_10343);
nor U10496 (N_10496,N_10281,N_10326);
and U10497 (N_10497,N_10300,N_10395);
and U10498 (N_10498,N_10336,N_10376);
xnor U10499 (N_10499,N_10248,N_10236);
xor U10500 (N_10500,N_10233,N_10356);
xnor U10501 (N_10501,N_10351,N_10332);
and U10502 (N_10502,N_10305,N_10218);
xnor U10503 (N_10503,N_10302,N_10362);
and U10504 (N_10504,N_10335,N_10282);
nand U10505 (N_10505,N_10303,N_10376);
xor U10506 (N_10506,N_10221,N_10211);
nand U10507 (N_10507,N_10217,N_10340);
and U10508 (N_10508,N_10249,N_10369);
xnor U10509 (N_10509,N_10364,N_10238);
and U10510 (N_10510,N_10207,N_10213);
xnor U10511 (N_10511,N_10367,N_10266);
nand U10512 (N_10512,N_10332,N_10399);
nand U10513 (N_10513,N_10262,N_10306);
or U10514 (N_10514,N_10393,N_10334);
nand U10515 (N_10515,N_10382,N_10298);
or U10516 (N_10516,N_10319,N_10245);
xnor U10517 (N_10517,N_10212,N_10322);
nor U10518 (N_10518,N_10305,N_10219);
xor U10519 (N_10519,N_10250,N_10380);
xnor U10520 (N_10520,N_10351,N_10245);
and U10521 (N_10521,N_10307,N_10359);
nor U10522 (N_10522,N_10281,N_10258);
nand U10523 (N_10523,N_10258,N_10312);
nand U10524 (N_10524,N_10273,N_10200);
nor U10525 (N_10525,N_10236,N_10395);
xnor U10526 (N_10526,N_10377,N_10247);
or U10527 (N_10527,N_10243,N_10267);
xor U10528 (N_10528,N_10289,N_10377);
nor U10529 (N_10529,N_10292,N_10224);
nor U10530 (N_10530,N_10238,N_10354);
or U10531 (N_10531,N_10213,N_10348);
nand U10532 (N_10532,N_10356,N_10362);
nor U10533 (N_10533,N_10229,N_10323);
nand U10534 (N_10534,N_10283,N_10220);
nand U10535 (N_10535,N_10387,N_10315);
or U10536 (N_10536,N_10310,N_10225);
or U10537 (N_10537,N_10324,N_10252);
xor U10538 (N_10538,N_10348,N_10325);
nand U10539 (N_10539,N_10353,N_10256);
or U10540 (N_10540,N_10394,N_10225);
nand U10541 (N_10541,N_10267,N_10302);
or U10542 (N_10542,N_10333,N_10209);
nor U10543 (N_10543,N_10235,N_10224);
or U10544 (N_10544,N_10399,N_10226);
nand U10545 (N_10545,N_10300,N_10386);
and U10546 (N_10546,N_10319,N_10332);
or U10547 (N_10547,N_10340,N_10240);
nor U10548 (N_10548,N_10244,N_10246);
and U10549 (N_10549,N_10373,N_10382);
nor U10550 (N_10550,N_10274,N_10321);
and U10551 (N_10551,N_10396,N_10351);
nand U10552 (N_10552,N_10370,N_10272);
nor U10553 (N_10553,N_10342,N_10354);
nand U10554 (N_10554,N_10214,N_10240);
xnor U10555 (N_10555,N_10285,N_10346);
or U10556 (N_10556,N_10204,N_10273);
nand U10557 (N_10557,N_10227,N_10224);
or U10558 (N_10558,N_10202,N_10207);
or U10559 (N_10559,N_10214,N_10222);
and U10560 (N_10560,N_10273,N_10369);
xor U10561 (N_10561,N_10255,N_10376);
nor U10562 (N_10562,N_10393,N_10354);
nor U10563 (N_10563,N_10224,N_10225);
xnor U10564 (N_10564,N_10324,N_10350);
xnor U10565 (N_10565,N_10394,N_10318);
nor U10566 (N_10566,N_10225,N_10392);
and U10567 (N_10567,N_10314,N_10235);
nor U10568 (N_10568,N_10375,N_10204);
or U10569 (N_10569,N_10379,N_10203);
xor U10570 (N_10570,N_10220,N_10230);
xor U10571 (N_10571,N_10246,N_10383);
or U10572 (N_10572,N_10261,N_10331);
or U10573 (N_10573,N_10389,N_10300);
nor U10574 (N_10574,N_10295,N_10223);
or U10575 (N_10575,N_10398,N_10326);
xor U10576 (N_10576,N_10331,N_10208);
nand U10577 (N_10577,N_10327,N_10320);
nand U10578 (N_10578,N_10256,N_10341);
nor U10579 (N_10579,N_10387,N_10229);
or U10580 (N_10580,N_10252,N_10369);
and U10581 (N_10581,N_10365,N_10261);
or U10582 (N_10582,N_10326,N_10360);
nor U10583 (N_10583,N_10365,N_10234);
xnor U10584 (N_10584,N_10398,N_10263);
xnor U10585 (N_10585,N_10259,N_10313);
or U10586 (N_10586,N_10234,N_10395);
nor U10587 (N_10587,N_10306,N_10380);
or U10588 (N_10588,N_10380,N_10260);
xor U10589 (N_10589,N_10276,N_10230);
xor U10590 (N_10590,N_10394,N_10320);
and U10591 (N_10591,N_10264,N_10238);
nor U10592 (N_10592,N_10218,N_10399);
xor U10593 (N_10593,N_10215,N_10224);
or U10594 (N_10594,N_10221,N_10238);
and U10595 (N_10595,N_10257,N_10385);
or U10596 (N_10596,N_10349,N_10260);
nor U10597 (N_10597,N_10272,N_10338);
nand U10598 (N_10598,N_10247,N_10266);
or U10599 (N_10599,N_10209,N_10321);
nand U10600 (N_10600,N_10497,N_10593);
or U10601 (N_10601,N_10558,N_10437);
nand U10602 (N_10602,N_10580,N_10546);
xnor U10603 (N_10603,N_10518,N_10404);
nand U10604 (N_10604,N_10428,N_10464);
nor U10605 (N_10605,N_10566,N_10587);
xnor U10606 (N_10606,N_10554,N_10448);
xnor U10607 (N_10607,N_10533,N_10576);
xor U10608 (N_10608,N_10571,N_10457);
or U10609 (N_10609,N_10569,N_10541);
xor U10610 (N_10610,N_10543,N_10458);
and U10611 (N_10611,N_10570,N_10461);
nand U10612 (N_10612,N_10473,N_10577);
nand U10613 (N_10613,N_10534,N_10421);
or U10614 (N_10614,N_10503,N_10438);
or U10615 (N_10615,N_10504,N_10487);
nand U10616 (N_10616,N_10500,N_10424);
nor U10617 (N_10617,N_10526,N_10462);
or U10618 (N_10618,N_10405,N_10557);
and U10619 (N_10619,N_10446,N_10562);
xnor U10620 (N_10620,N_10559,N_10548);
and U10621 (N_10621,N_10444,N_10535);
or U10622 (N_10622,N_10422,N_10555);
nor U10623 (N_10623,N_10590,N_10493);
nor U10624 (N_10624,N_10469,N_10476);
nor U10625 (N_10625,N_10494,N_10578);
xnor U10626 (N_10626,N_10435,N_10478);
xor U10627 (N_10627,N_10521,N_10505);
and U10628 (N_10628,N_10407,N_10412);
nor U10629 (N_10629,N_10452,N_10402);
or U10630 (N_10630,N_10418,N_10517);
xor U10631 (N_10631,N_10551,N_10550);
and U10632 (N_10632,N_10575,N_10519);
or U10633 (N_10633,N_10544,N_10479);
nor U10634 (N_10634,N_10513,N_10455);
nor U10635 (N_10635,N_10465,N_10463);
or U10636 (N_10636,N_10403,N_10467);
xor U10637 (N_10637,N_10483,N_10434);
nor U10638 (N_10638,N_10433,N_10573);
or U10639 (N_10639,N_10511,N_10415);
nor U10640 (N_10640,N_10549,N_10529);
or U10641 (N_10641,N_10498,N_10472);
nor U10642 (N_10642,N_10409,N_10481);
or U10643 (N_10643,N_10413,N_10419);
or U10644 (N_10644,N_10508,N_10515);
nand U10645 (N_10645,N_10430,N_10471);
xnor U10646 (N_10646,N_10441,N_10445);
xor U10647 (N_10647,N_10443,N_10496);
or U10648 (N_10648,N_10583,N_10432);
xnor U10649 (N_10649,N_10522,N_10524);
and U10650 (N_10650,N_10540,N_10482);
xor U10651 (N_10651,N_10574,N_10568);
nand U10652 (N_10652,N_10523,N_10506);
nand U10653 (N_10653,N_10596,N_10449);
xor U10654 (N_10654,N_10561,N_10408);
xnor U10655 (N_10655,N_10563,N_10490);
or U10656 (N_10656,N_10410,N_10456);
nand U10657 (N_10657,N_10588,N_10507);
nand U10658 (N_10658,N_10488,N_10556);
xor U10659 (N_10659,N_10470,N_10436);
xnor U10660 (N_10660,N_10466,N_10547);
and U10661 (N_10661,N_10589,N_10429);
and U10662 (N_10662,N_10401,N_10538);
nand U10663 (N_10663,N_10509,N_10599);
and U10664 (N_10664,N_10485,N_10579);
xnor U10665 (N_10665,N_10423,N_10501);
and U10666 (N_10666,N_10442,N_10420);
nor U10667 (N_10667,N_10595,N_10460);
xnor U10668 (N_10668,N_10451,N_10565);
nor U10669 (N_10669,N_10597,N_10416);
nor U10670 (N_10670,N_10499,N_10581);
nand U10671 (N_10671,N_10453,N_10427);
and U10672 (N_10672,N_10447,N_10425);
nand U10673 (N_10673,N_10525,N_10553);
xor U10674 (N_10674,N_10530,N_10531);
and U10675 (N_10675,N_10492,N_10572);
nor U10676 (N_10676,N_10585,N_10439);
nor U10677 (N_10677,N_10468,N_10520);
or U10678 (N_10678,N_10510,N_10414);
or U10679 (N_10679,N_10539,N_10564);
and U10680 (N_10680,N_10454,N_10459);
nor U10681 (N_10681,N_10560,N_10516);
and U10682 (N_10682,N_10489,N_10591);
xnor U10683 (N_10683,N_10584,N_10502);
or U10684 (N_10684,N_10532,N_10528);
xnor U10685 (N_10685,N_10495,N_10545);
nor U10686 (N_10686,N_10474,N_10431);
and U10687 (N_10687,N_10598,N_10411);
xor U10688 (N_10688,N_10594,N_10475);
or U10689 (N_10689,N_10586,N_10542);
or U10690 (N_10690,N_10512,N_10537);
xnor U10691 (N_10691,N_10592,N_10582);
nor U10692 (N_10692,N_10486,N_10514);
nor U10693 (N_10693,N_10527,N_10450);
nor U10694 (N_10694,N_10400,N_10491);
xnor U10695 (N_10695,N_10567,N_10536);
nor U10696 (N_10696,N_10440,N_10406);
nor U10697 (N_10697,N_10417,N_10484);
nor U10698 (N_10698,N_10480,N_10477);
or U10699 (N_10699,N_10552,N_10426);
nor U10700 (N_10700,N_10581,N_10580);
nand U10701 (N_10701,N_10405,N_10528);
nand U10702 (N_10702,N_10507,N_10568);
and U10703 (N_10703,N_10436,N_10454);
and U10704 (N_10704,N_10431,N_10508);
xor U10705 (N_10705,N_10504,N_10543);
nor U10706 (N_10706,N_10526,N_10562);
nand U10707 (N_10707,N_10414,N_10537);
nor U10708 (N_10708,N_10547,N_10578);
or U10709 (N_10709,N_10458,N_10524);
xnor U10710 (N_10710,N_10576,N_10592);
and U10711 (N_10711,N_10459,N_10407);
xor U10712 (N_10712,N_10510,N_10576);
and U10713 (N_10713,N_10570,N_10438);
nand U10714 (N_10714,N_10477,N_10568);
nand U10715 (N_10715,N_10485,N_10551);
xor U10716 (N_10716,N_10519,N_10426);
or U10717 (N_10717,N_10496,N_10550);
or U10718 (N_10718,N_10457,N_10452);
xor U10719 (N_10719,N_10509,N_10436);
and U10720 (N_10720,N_10577,N_10470);
xor U10721 (N_10721,N_10455,N_10491);
xor U10722 (N_10722,N_10515,N_10528);
and U10723 (N_10723,N_10410,N_10526);
nor U10724 (N_10724,N_10468,N_10516);
nor U10725 (N_10725,N_10470,N_10432);
or U10726 (N_10726,N_10552,N_10428);
nand U10727 (N_10727,N_10545,N_10549);
xnor U10728 (N_10728,N_10569,N_10487);
or U10729 (N_10729,N_10526,N_10525);
nor U10730 (N_10730,N_10536,N_10465);
xnor U10731 (N_10731,N_10558,N_10469);
or U10732 (N_10732,N_10586,N_10498);
nand U10733 (N_10733,N_10507,N_10520);
or U10734 (N_10734,N_10444,N_10503);
or U10735 (N_10735,N_10585,N_10563);
nor U10736 (N_10736,N_10524,N_10454);
or U10737 (N_10737,N_10410,N_10423);
or U10738 (N_10738,N_10431,N_10475);
nor U10739 (N_10739,N_10476,N_10504);
nand U10740 (N_10740,N_10442,N_10431);
nand U10741 (N_10741,N_10522,N_10535);
and U10742 (N_10742,N_10531,N_10570);
or U10743 (N_10743,N_10405,N_10583);
or U10744 (N_10744,N_10437,N_10477);
or U10745 (N_10745,N_10590,N_10466);
and U10746 (N_10746,N_10495,N_10412);
or U10747 (N_10747,N_10536,N_10480);
xor U10748 (N_10748,N_10511,N_10469);
nor U10749 (N_10749,N_10442,N_10411);
nand U10750 (N_10750,N_10555,N_10524);
xnor U10751 (N_10751,N_10409,N_10594);
or U10752 (N_10752,N_10567,N_10500);
nor U10753 (N_10753,N_10434,N_10580);
nand U10754 (N_10754,N_10514,N_10530);
nor U10755 (N_10755,N_10597,N_10572);
or U10756 (N_10756,N_10425,N_10407);
nand U10757 (N_10757,N_10526,N_10570);
or U10758 (N_10758,N_10502,N_10412);
nor U10759 (N_10759,N_10456,N_10593);
and U10760 (N_10760,N_10412,N_10588);
or U10761 (N_10761,N_10410,N_10467);
xor U10762 (N_10762,N_10498,N_10402);
nor U10763 (N_10763,N_10598,N_10413);
nand U10764 (N_10764,N_10591,N_10592);
xnor U10765 (N_10765,N_10564,N_10429);
or U10766 (N_10766,N_10567,N_10583);
nand U10767 (N_10767,N_10580,N_10567);
or U10768 (N_10768,N_10483,N_10466);
and U10769 (N_10769,N_10424,N_10596);
or U10770 (N_10770,N_10458,N_10404);
nor U10771 (N_10771,N_10467,N_10418);
and U10772 (N_10772,N_10552,N_10451);
xor U10773 (N_10773,N_10596,N_10538);
xor U10774 (N_10774,N_10546,N_10440);
or U10775 (N_10775,N_10498,N_10473);
and U10776 (N_10776,N_10459,N_10415);
and U10777 (N_10777,N_10405,N_10541);
or U10778 (N_10778,N_10582,N_10531);
nand U10779 (N_10779,N_10591,N_10531);
nand U10780 (N_10780,N_10594,N_10478);
or U10781 (N_10781,N_10433,N_10567);
and U10782 (N_10782,N_10585,N_10530);
nor U10783 (N_10783,N_10486,N_10517);
xor U10784 (N_10784,N_10553,N_10480);
or U10785 (N_10785,N_10552,N_10473);
nor U10786 (N_10786,N_10518,N_10480);
or U10787 (N_10787,N_10599,N_10445);
or U10788 (N_10788,N_10500,N_10515);
and U10789 (N_10789,N_10579,N_10494);
nand U10790 (N_10790,N_10463,N_10525);
nand U10791 (N_10791,N_10581,N_10406);
nand U10792 (N_10792,N_10504,N_10579);
nand U10793 (N_10793,N_10473,N_10561);
or U10794 (N_10794,N_10414,N_10593);
nor U10795 (N_10795,N_10567,N_10539);
nor U10796 (N_10796,N_10444,N_10460);
nor U10797 (N_10797,N_10540,N_10515);
and U10798 (N_10798,N_10483,N_10556);
nand U10799 (N_10799,N_10513,N_10453);
or U10800 (N_10800,N_10733,N_10706);
nor U10801 (N_10801,N_10723,N_10720);
xnor U10802 (N_10802,N_10680,N_10788);
and U10803 (N_10803,N_10747,N_10745);
or U10804 (N_10804,N_10644,N_10697);
nor U10805 (N_10805,N_10634,N_10728);
or U10806 (N_10806,N_10732,N_10712);
xnor U10807 (N_10807,N_10770,N_10662);
and U10808 (N_10808,N_10762,N_10650);
nor U10809 (N_10809,N_10795,N_10725);
nor U10810 (N_10810,N_10798,N_10763);
nand U10811 (N_10811,N_10666,N_10628);
xor U10812 (N_10812,N_10738,N_10799);
and U10813 (N_10813,N_10699,N_10619);
and U10814 (N_10814,N_10754,N_10794);
and U10815 (N_10815,N_10711,N_10748);
nor U10816 (N_10816,N_10627,N_10753);
nor U10817 (N_10817,N_10740,N_10615);
xnor U10818 (N_10818,N_10769,N_10651);
or U10819 (N_10819,N_10672,N_10792);
or U10820 (N_10820,N_10750,N_10622);
nand U10821 (N_10821,N_10756,N_10760);
or U10822 (N_10822,N_10677,N_10653);
nor U10823 (N_10823,N_10759,N_10621);
or U10824 (N_10824,N_10718,N_10772);
nand U10825 (N_10825,N_10702,N_10601);
nor U10826 (N_10826,N_10708,N_10613);
and U10827 (N_10827,N_10624,N_10746);
and U10828 (N_10828,N_10700,N_10668);
and U10829 (N_10829,N_10657,N_10771);
xnor U10830 (N_10830,N_10638,N_10695);
nand U10831 (N_10831,N_10710,N_10678);
or U10832 (N_10832,N_10658,N_10682);
nor U10833 (N_10833,N_10781,N_10761);
or U10834 (N_10834,N_10609,N_10716);
nor U10835 (N_10835,N_10780,N_10612);
and U10836 (N_10836,N_10715,N_10656);
and U10837 (N_10837,N_10630,N_10793);
nand U10838 (N_10838,N_10623,N_10783);
nor U10839 (N_10839,N_10643,N_10669);
nand U10840 (N_10840,N_10734,N_10703);
and U10841 (N_10841,N_10757,N_10641);
and U10842 (N_10842,N_10721,N_10696);
nor U10843 (N_10843,N_10743,N_10691);
nand U10844 (N_10844,N_10661,N_10778);
and U10845 (N_10845,N_10637,N_10646);
or U10846 (N_10846,N_10704,N_10776);
nor U10847 (N_10847,N_10633,N_10797);
or U10848 (N_10848,N_10726,N_10654);
xor U10849 (N_10849,N_10614,N_10603);
nand U10850 (N_10850,N_10705,N_10735);
xnor U10851 (N_10851,N_10629,N_10602);
or U10852 (N_10852,N_10681,N_10667);
xnor U10853 (N_10853,N_10786,N_10604);
or U10854 (N_10854,N_10683,N_10722);
nor U10855 (N_10855,N_10736,N_10664);
nand U10856 (N_10856,N_10719,N_10782);
nor U10857 (N_10857,N_10766,N_10655);
xnor U10858 (N_10858,N_10777,N_10767);
nand U10859 (N_10859,N_10671,N_10730);
or U10860 (N_10860,N_10775,N_10694);
or U10861 (N_10861,N_10616,N_10779);
nand U10862 (N_10862,N_10687,N_10749);
nor U10863 (N_10863,N_10625,N_10685);
and U10864 (N_10864,N_10618,N_10635);
xnor U10865 (N_10865,N_10773,N_10688);
xnor U10866 (N_10866,N_10751,N_10676);
nor U10867 (N_10867,N_10605,N_10673);
xor U10868 (N_10868,N_10639,N_10692);
and U10869 (N_10869,N_10758,N_10665);
xnor U10870 (N_10870,N_10600,N_10689);
xnor U10871 (N_10871,N_10713,N_10724);
nand U10872 (N_10872,N_10606,N_10659);
and U10873 (N_10873,N_10737,N_10729);
nand U10874 (N_10874,N_10774,N_10701);
xor U10875 (N_10875,N_10789,N_10631);
or U10876 (N_10876,N_10607,N_10647);
nor U10877 (N_10877,N_10610,N_10707);
xnor U10878 (N_10878,N_10690,N_10611);
nor U10879 (N_10879,N_10674,N_10660);
and U10880 (N_10880,N_10741,N_10709);
or U10881 (N_10881,N_10620,N_10632);
nand U10882 (N_10882,N_10755,N_10768);
nand U10883 (N_10883,N_10608,N_10765);
or U10884 (N_10884,N_10640,N_10791);
or U10885 (N_10885,N_10714,N_10790);
and U10886 (N_10886,N_10649,N_10670);
nor U10887 (N_10887,N_10739,N_10698);
or U10888 (N_10888,N_10686,N_10663);
xnor U10889 (N_10889,N_10675,N_10679);
nand U10890 (N_10890,N_10693,N_10648);
nor U10891 (N_10891,N_10636,N_10642);
xor U10892 (N_10892,N_10626,N_10764);
and U10893 (N_10893,N_10785,N_10784);
and U10894 (N_10894,N_10652,N_10742);
xnor U10895 (N_10895,N_10796,N_10744);
nor U10896 (N_10896,N_10717,N_10617);
nor U10897 (N_10897,N_10645,N_10787);
xor U10898 (N_10898,N_10727,N_10684);
nor U10899 (N_10899,N_10752,N_10731);
and U10900 (N_10900,N_10730,N_10746);
and U10901 (N_10901,N_10687,N_10651);
xor U10902 (N_10902,N_10658,N_10622);
or U10903 (N_10903,N_10691,N_10733);
or U10904 (N_10904,N_10783,N_10687);
nor U10905 (N_10905,N_10725,N_10624);
and U10906 (N_10906,N_10678,N_10711);
nand U10907 (N_10907,N_10601,N_10675);
and U10908 (N_10908,N_10794,N_10762);
nor U10909 (N_10909,N_10794,N_10757);
or U10910 (N_10910,N_10623,N_10661);
nand U10911 (N_10911,N_10712,N_10674);
or U10912 (N_10912,N_10651,N_10792);
nor U10913 (N_10913,N_10719,N_10699);
nor U10914 (N_10914,N_10665,N_10781);
and U10915 (N_10915,N_10765,N_10612);
and U10916 (N_10916,N_10792,N_10745);
xor U10917 (N_10917,N_10666,N_10670);
xnor U10918 (N_10918,N_10621,N_10723);
and U10919 (N_10919,N_10761,N_10667);
and U10920 (N_10920,N_10775,N_10763);
nand U10921 (N_10921,N_10689,N_10722);
and U10922 (N_10922,N_10676,N_10622);
or U10923 (N_10923,N_10755,N_10793);
and U10924 (N_10924,N_10618,N_10612);
nand U10925 (N_10925,N_10797,N_10715);
and U10926 (N_10926,N_10709,N_10748);
nor U10927 (N_10927,N_10688,N_10737);
xor U10928 (N_10928,N_10610,N_10755);
and U10929 (N_10929,N_10709,N_10771);
xor U10930 (N_10930,N_10764,N_10745);
or U10931 (N_10931,N_10642,N_10631);
nor U10932 (N_10932,N_10740,N_10674);
or U10933 (N_10933,N_10694,N_10716);
nor U10934 (N_10934,N_10697,N_10631);
nor U10935 (N_10935,N_10740,N_10760);
nor U10936 (N_10936,N_10695,N_10618);
and U10937 (N_10937,N_10693,N_10701);
xnor U10938 (N_10938,N_10691,N_10721);
or U10939 (N_10939,N_10771,N_10670);
nor U10940 (N_10940,N_10627,N_10799);
nor U10941 (N_10941,N_10692,N_10753);
nand U10942 (N_10942,N_10600,N_10743);
nor U10943 (N_10943,N_10754,N_10625);
nand U10944 (N_10944,N_10651,N_10765);
nand U10945 (N_10945,N_10732,N_10704);
nor U10946 (N_10946,N_10716,N_10710);
or U10947 (N_10947,N_10642,N_10661);
and U10948 (N_10948,N_10708,N_10712);
nor U10949 (N_10949,N_10743,N_10709);
nand U10950 (N_10950,N_10759,N_10676);
and U10951 (N_10951,N_10785,N_10761);
nor U10952 (N_10952,N_10691,N_10630);
xnor U10953 (N_10953,N_10730,N_10642);
nor U10954 (N_10954,N_10780,N_10684);
or U10955 (N_10955,N_10654,N_10784);
or U10956 (N_10956,N_10625,N_10628);
or U10957 (N_10957,N_10721,N_10760);
and U10958 (N_10958,N_10602,N_10674);
or U10959 (N_10959,N_10659,N_10760);
and U10960 (N_10960,N_10760,N_10769);
xor U10961 (N_10961,N_10688,N_10763);
or U10962 (N_10962,N_10739,N_10606);
nand U10963 (N_10963,N_10605,N_10796);
xor U10964 (N_10964,N_10774,N_10712);
and U10965 (N_10965,N_10607,N_10657);
or U10966 (N_10966,N_10726,N_10730);
and U10967 (N_10967,N_10684,N_10700);
and U10968 (N_10968,N_10784,N_10731);
nor U10969 (N_10969,N_10743,N_10721);
xnor U10970 (N_10970,N_10726,N_10602);
and U10971 (N_10971,N_10702,N_10692);
xor U10972 (N_10972,N_10657,N_10787);
xnor U10973 (N_10973,N_10663,N_10654);
nand U10974 (N_10974,N_10651,N_10602);
nand U10975 (N_10975,N_10657,N_10731);
or U10976 (N_10976,N_10776,N_10672);
nand U10977 (N_10977,N_10649,N_10673);
or U10978 (N_10978,N_10736,N_10711);
xor U10979 (N_10979,N_10636,N_10798);
nor U10980 (N_10980,N_10680,N_10703);
xor U10981 (N_10981,N_10788,N_10662);
xnor U10982 (N_10982,N_10655,N_10770);
xor U10983 (N_10983,N_10776,N_10765);
or U10984 (N_10984,N_10759,N_10614);
nand U10985 (N_10985,N_10617,N_10618);
nand U10986 (N_10986,N_10602,N_10658);
and U10987 (N_10987,N_10724,N_10793);
xnor U10988 (N_10988,N_10784,N_10732);
nand U10989 (N_10989,N_10686,N_10748);
and U10990 (N_10990,N_10735,N_10608);
or U10991 (N_10991,N_10645,N_10610);
nand U10992 (N_10992,N_10737,N_10739);
and U10993 (N_10993,N_10679,N_10760);
nor U10994 (N_10994,N_10723,N_10618);
or U10995 (N_10995,N_10799,N_10764);
nand U10996 (N_10996,N_10606,N_10759);
nor U10997 (N_10997,N_10607,N_10654);
xor U10998 (N_10998,N_10780,N_10785);
xnor U10999 (N_10999,N_10752,N_10644);
and U11000 (N_11000,N_10995,N_10899);
nand U11001 (N_11001,N_10841,N_10906);
xor U11002 (N_11002,N_10832,N_10850);
xor U11003 (N_11003,N_10986,N_10955);
nand U11004 (N_11004,N_10957,N_10867);
and U11005 (N_11005,N_10944,N_10990);
nand U11006 (N_11006,N_10814,N_10881);
or U11007 (N_11007,N_10868,N_10828);
nor U11008 (N_11008,N_10985,N_10908);
nand U11009 (N_11009,N_10831,N_10958);
xnor U11010 (N_11010,N_10921,N_10945);
nand U11011 (N_11011,N_10970,N_10893);
and U11012 (N_11012,N_10938,N_10894);
nand U11013 (N_11013,N_10956,N_10964);
xor U11014 (N_11014,N_10960,N_10910);
nand U11015 (N_11015,N_10837,N_10948);
nand U11016 (N_11016,N_10816,N_10890);
nand U11017 (N_11017,N_10805,N_10822);
and U11018 (N_11018,N_10982,N_10834);
nand U11019 (N_11019,N_10809,N_10838);
nand U11020 (N_11020,N_10847,N_10917);
xor U11021 (N_11021,N_10929,N_10999);
nand U11022 (N_11022,N_10974,N_10839);
or U11023 (N_11023,N_10933,N_10876);
nor U11024 (N_11024,N_10873,N_10994);
or U11025 (N_11025,N_10940,N_10845);
and U11026 (N_11026,N_10951,N_10934);
nor U11027 (N_11027,N_10806,N_10820);
nand U11028 (N_11028,N_10861,N_10930);
nand U11029 (N_11029,N_10836,N_10898);
or U11030 (N_11030,N_10833,N_10927);
nand U11031 (N_11031,N_10878,N_10924);
nor U11032 (N_11032,N_10907,N_10966);
xor U11033 (N_11033,N_10961,N_10991);
or U11034 (N_11034,N_10928,N_10942);
xor U11035 (N_11035,N_10920,N_10926);
nand U11036 (N_11036,N_10988,N_10801);
and U11037 (N_11037,N_10952,N_10973);
xnor U11038 (N_11038,N_10887,N_10932);
nor U11039 (N_11039,N_10849,N_10853);
nor U11040 (N_11040,N_10891,N_10923);
and U11041 (N_11041,N_10998,N_10824);
nor U11042 (N_11042,N_10830,N_10874);
and U11043 (N_11043,N_10871,N_10968);
xor U11044 (N_11044,N_10912,N_10866);
or U11045 (N_11045,N_10901,N_10877);
xor U11046 (N_11046,N_10855,N_10807);
or U11047 (N_11047,N_10872,N_10935);
nor U11048 (N_11048,N_10902,N_10984);
nor U11049 (N_11049,N_10802,N_10888);
nand U11050 (N_11050,N_10827,N_10804);
nor U11051 (N_11051,N_10953,N_10875);
and U11052 (N_11052,N_10884,N_10880);
or U11053 (N_11053,N_10865,N_10900);
or U11054 (N_11054,N_10949,N_10925);
and U11055 (N_11055,N_10862,N_10829);
nor U11056 (N_11056,N_10840,N_10800);
nand U11057 (N_11057,N_10978,N_10863);
or U11058 (N_11058,N_10821,N_10914);
nand U11059 (N_11059,N_10971,N_10922);
nand U11060 (N_11060,N_10864,N_10818);
nand U11061 (N_11061,N_10980,N_10859);
nor U11062 (N_11062,N_10936,N_10857);
nand U11063 (N_11063,N_10883,N_10911);
nor U11064 (N_11064,N_10909,N_10989);
nand U11065 (N_11065,N_10886,N_10993);
or U11066 (N_11066,N_10916,N_10941);
or U11067 (N_11067,N_10903,N_10889);
or U11068 (N_11068,N_10896,N_10969);
xor U11069 (N_11069,N_10915,N_10846);
nor U11070 (N_11070,N_10870,N_10882);
and U11071 (N_11071,N_10848,N_10858);
nor U11072 (N_11072,N_10904,N_10972);
nand U11073 (N_11073,N_10962,N_10996);
and U11074 (N_11074,N_10892,N_10918);
xnor U11075 (N_11075,N_10856,N_10967);
and U11076 (N_11076,N_10987,N_10819);
nor U11077 (N_11077,N_10812,N_10815);
nand U11078 (N_11078,N_10913,N_10869);
xor U11079 (N_11079,N_10947,N_10808);
and U11080 (N_11080,N_10842,N_10897);
and U11081 (N_11081,N_10979,N_10997);
xnor U11082 (N_11082,N_10854,N_10977);
xnor U11083 (N_11083,N_10826,N_10844);
nand U11084 (N_11084,N_10843,N_10817);
and U11085 (N_11085,N_10992,N_10976);
nor U11086 (N_11086,N_10803,N_10813);
xnor U11087 (N_11087,N_10860,N_10905);
nand U11088 (N_11088,N_10835,N_10983);
or U11089 (N_11089,N_10937,N_10950);
xor U11090 (N_11090,N_10879,N_10981);
or U11091 (N_11091,N_10943,N_10825);
xor U11092 (N_11092,N_10851,N_10954);
nor U11093 (N_11093,N_10885,N_10895);
or U11094 (N_11094,N_10823,N_10963);
nand U11095 (N_11095,N_10810,N_10946);
and U11096 (N_11096,N_10965,N_10975);
nor U11097 (N_11097,N_10959,N_10852);
nand U11098 (N_11098,N_10919,N_10811);
xnor U11099 (N_11099,N_10931,N_10939);
or U11100 (N_11100,N_10926,N_10969);
nor U11101 (N_11101,N_10967,N_10862);
or U11102 (N_11102,N_10922,N_10991);
and U11103 (N_11103,N_10959,N_10978);
nor U11104 (N_11104,N_10812,N_10967);
xor U11105 (N_11105,N_10952,N_10985);
nand U11106 (N_11106,N_10877,N_10881);
nand U11107 (N_11107,N_10888,N_10818);
nand U11108 (N_11108,N_10883,N_10948);
nand U11109 (N_11109,N_10849,N_10883);
nand U11110 (N_11110,N_10977,N_10997);
nand U11111 (N_11111,N_10891,N_10983);
and U11112 (N_11112,N_10886,N_10905);
or U11113 (N_11113,N_10968,N_10808);
nor U11114 (N_11114,N_10960,N_10956);
nor U11115 (N_11115,N_10945,N_10966);
nor U11116 (N_11116,N_10818,N_10899);
nor U11117 (N_11117,N_10854,N_10953);
xor U11118 (N_11118,N_10844,N_10907);
and U11119 (N_11119,N_10966,N_10860);
nand U11120 (N_11120,N_10998,N_10930);
or U11121 (N_11121,N_10911,N_10945);
or U11122 (N_11122,N_10983,N_10884);
or U11123 (N_11123,N_10960,N_10894);
nand U11124 (N_11124,N_10926,N_10943);
nand U11125 (N_11125,N_10977,N_10949);
or U11126 (N_11126,N_10957,N_10886);
or U11127 (N_11127,N_10956,N_10955);
or U11128 (N_11128,N_10918,N_10801);
and U11129 (N_11129,N_10826,N_10901);
or U11130 (N_11130,N_10802,N_10815);
nor U11131 (N_11131,N_10922,N_10821);
and U11132 (N_11132,N_10808,N_10833);
xnor U11133 (N_11133,N_10804,N_10859);
and U11134 (N_11134,N_10851,N_10914);
and U11135 (N_11135,N_10923,N_10974);
and U11136 (N_11136,N_10949,N_10944);
xor U11137 (N_11137,N_10813,N_10810);
nor U11138 (N_11138,N_10945,N_10861);
or U11139 (N_11139,N_10997,N_10957);
and U11140 (N_11140,N_10857,N_10824);
nor U11141 (N_11141,N_10877,N_10807);
nor U11142 (N_11142,N_10843,N_10931);
xor U11143 (N_11143,N_10910,N_10904);
xnor U11144 (N_11144,N_10992,N_10928);
nor U11145 (N_11145,N_10972,N_10991);
xnor U11146 (N_11146,N_10864,N_10961);
and U11147 (N_11147,N_10891,N_10973);
and U11148 (N_11148,N_10944,N_10810);
xor U11149 (N_11149,N_10917,N_10871);
nor U11150 (N_11150,N_10955,N_10944);
nand U11151 (N_11151,N_10952,N_10877);
nor U11152 (N_11152,N_10871,N_10958);
xnor U11153 (N_11153,N_10975,N_10931);
nand U11154 (N_11154,N_10921,N_10804);
nand U11155 (N_11155,N_10956,N_10876);
and U11156 (N_11156,N_10932,N_10815);
or U11157 (N_11157,N_10936,N_10852);
nor U11158 (N_11158,N_10944,N_10961);
nor U11159 (N_11159,N_10872,N_10886);
and U11160 (N_11160,N_10858,N_10939);
nor U11161 (N_11161,N_10886,N_10843);
nand U11162 (N_11162,N_10939,N_10977);
xnor U11163 (N_11163,N_10917,N_10941);
or U11164 (N_11164,N_10806,N_10894);
or U11165 (N_11165,N_10929,N_10851);
nor U11166 (N_11166,N_10821,N_10867);
nand U11167 (N_11167,N_10850,N_10929);
or U11168 (N_11168,N_10992,N_10810);
nor U11169 (N_11169,N_10813,N_10999);
nor U11170 (N_11170,N_10803,N_10848);
or U11171 (N_11171,N_10918,N_10986);
nor U11172 (N_11172,N_10887,N_10845);
or U11173 (N_11173,N_10931,N_10984);
xor U11174 (N_11174,N_10837,N_10973);
and U11175 (N_11175,N_10888,N_10814);
xnor U11176 (N_11176,N_10829,N_10845);
nor U11177 (N_11177,N_10991,N_10916);
nor U11178 (N_11178,N_10932,N_10893);
and U11179 (N_11179,N_10805,N_10811);
or U11180 (N_11180,N_10859,N_10916);
and U11181 (N_11181,N_10908,N_10975);
and U11182 (N_11182,N_10945,N_10845);
and U11183 (N_11183,N_10908,N_10984);
and U11184 (N_11184,N_10933,N_10950);
xor U11185 (N_11185,N_10936,N_10894);
nor U11186 (N_11186,N_10927,N_10908);
or U11187 (N_11187,N_10922,N_10892);
or U11188 (N_11188,N_10844,N_10938);
xnor U11189 (N_11189,N_10957,N_10830);
and U11190 (N_11190,N_10954,N_10849);
xnor U11191 (N_11191,N_10824,N_10832);
xnor U11192 (N_11192,N_10912,N_10833);
or U11193 (N_11193,N_10862,N_10972);
or U11194 (N_11194,N_10843,N_10939);
xor U11195 (N_11195,N_10830,N_10812);
nor U11196 (N_11196,N_10919,N_10996);
or U11197 (N_11197,N_10990,N_10813);
nor U11198 (N_11198,N_10895,N_10957);
nand U11199 (N_11199,N_10842,N_10899);
or U11200 (N_11200,N_11100,N_11143);
or U11201 (N_11201,N_11175,N_11128);
xor U11202 (N_11202,N_11088,N_11033);
and U11203 (N_11203,N_11045,N_11115);
xor U11204 (N_11204,N_11192,N_11073);
nor U11205 (N_11205,N_11164,N_11172);
nand U11206 (N_11206,N_11180,N_11022);
nand U11207 (N_11207,N_11184,N_11080);
xor U11208 (N_11208,N_11044,N_11144);
nand U11209 (N_11209,N_11104,N_11125);
or U11210 (N_11210,N_11032,N_11089);
nor U11211 (N_11211,N_11159,N_11136);
nor U11212 (N_11212,N_11038,N_11004);
or U11213 (N_11213,N_11047,N_11106);
nand U11214 (N_11214,N_11151,N_11096);
and U11215 (N_11215,N_11034,N_11024);
nand U11216 (N_11216,N_11086,N_11085);
or U11217 (N_11217,N_11193,N_11176);
nand U11218 (N_11218,N_11148,N_11134);
nand U11219 (N_11219,N_11036,N_11035);
nor U11220 (N_11220,N_11025,N_11083);
nand U11221 (N_11221,N_11195,N_11166);
xor U11222 (N_11222,N_11087,N_11040);
xnor U11223 (N_11223,N_11050,N_11152);
nand U11224 (N_11224,N_11124,N_11116);
and U11225 (N_11225,N_11093,N_11140);
xnor U11226 (N_11226,N_11133,N_11163);
nor U11227 (N_11227,N_11101,N_11103);
nand U11228 (N_11228,N_11186,N_11170);
or U11229 (N_11229,N_11005,N_11183);
xnor U11230 (N_11230,N_11006,N_11196);
nor U11231 (N_11231,N_11135,N_11127);
and U11232 (N_11232,N_11132,N_11185);
and U11233 (N_11233,N_11191,N_11165);
and U11234 (N_11234,N_11173,N_11149);
or U11235 (N_11235,N_11002,N_11008);
and U11236 (N_11236,N_11131,N_11137);
or U11237 (N_11237,N_11190,N_11070);
and U11238 (N_11238,N_11039,N_11054);
nor U11239 (N_11239,N_11154,N_11189);
and U11240 (N_11240,N_11015,N_11065);
nand U11241 (N_11241,N_11042,N_11120);
or U11242 (N_11242,N_11078,N_11119);
or U11243 (N_11243,N_11082,N_11059);
xor U11244 (N_11244,N_11112,N_11097);
or U11245 (N_11245,N_11056,N_11066);
nor U11246 (N_11246,N_11197,N_11198);
or U11247 (N_11247,N_11026,N_11153);
xnor U11248 (N_11248,N_11155,N_11156);
nor U11249 (N_11249,N_11023,N_11074);
xnor U11250 (N_11250,N_11064,N_11011);
xnor U11251 (N_11251,N_11061,N_11091);
or U11252 (N_11252,N_11010,N_11142);
nand U11253 (N_11253,N_11123,N_11177);
and U11254 (N_11254,N_11053,N_11157);
xnor U11255 (N_11255,N_11020,N_11090);
and U11256 (N_11256,N_11094,N_11147);
and U11257 (N_11257,N_11138,N_11145);
nor U11258 (N_11258,N_11076,N_11063);
xor U11259 (N_11259,N_11055,N_11079);
or U11260 (N_11260,N_11129,N_11069);
xnor U11261 (N_11261,N_11046,N_11108);
or U11262 (N_11262,N_11169,N_11058);
xnor U11263 (N_11263,N_11187,N_11048);
nor U11264 (N_11264,N_11111,N_11081);
xnor U11265 (N_11265,N_11113,N_11077);
xnor U11266 (N_11266,N_11049,N_11084);
xnor U11267 (N_11267,N_11167,N_11099);
or U11268 (N_11268,N_11030,N_11109);
nor U11269 (N_11269,N_11095,N_11179);
nor U11270 (N_11270,N_11027,N_11107);
nand U11271 (N_11271,N_11150,N_11003);
nand U11272 (N_11272,N_11071,N_11199);
nand U11273 (N_11273,N_11013,N_11188);
or U11274 (N_11274,N_11052,N_11075);
or U11275 (N_11275,N_11067,N_11021);
or U11276 (N_11276,N_11029,N_11181);
and U11277 (N_11277,N_11037,N_11068);
nor U11278 (N_11278,N_11174,N_11018);
or U11279 (N_11279,N_11194,N_11126);
nand U11280 (N_11280,N_11171,N_11017);
nor U11281 (N_11281,N_11105,N_11146);
nand U11282 (N_11282,N_11016,N_11012);
nor U11283 (N_11283,N_11031,N_11168);
nand U11284 (N_11284,N_11110,N_11009);
nand U11285 (N_11285,N_11139,N_11072);
xor U11286 (N_11286,N_11019,N_11014);
or U11287 (N_11287,N_11114,N_11182);
xnor U11288 (N_11288,N_11007,N_11162);
nand U11289 (N_11289,N_11028,N_11160);
nor U11290 (N_11290,N_11051,N_11178);
xnor U11291 (N_11291,N_11098,N_11057);
and U11292 (N_11292,N_11158,N_11000);
xor U11293 (N_11293,N_11001,N_11121);
xor U11294 (N_11294,N_11092,N_11118);
nand U11295 (N_11295,N_11102,N_11161);
nor U11296 (N_11296,N_11043,N_11141);
nand U11297 (N_11297,N_11117,N_11060);
nand U11298 (N_11298,N_11041,N_11130);
or U11299 (N_11299,N_11062,N_11122);
xor U11300 (N_11300,N_11145,N_11096);
nand U11301 (N_11301,N_11079,N_11011);
nand U11302 (N_11302,N_11135,N_11046);
xnor U11303 (N_11303,N_11113,N_11104);
nand U11304 (N_11304,N_11180,N_11136);
or U11305 (N_11305,N_11053,N_11181);
and U11306 (N_11306,N_11182,N_11189);
and U11307 (N_11307,N_11169,N_11149);
xnor U11308 (N_11308,N_11100,N_11003);
nor U11309 (N_11309,N_11141,N_11158);
xnor U11310 (N_11310,N_11172,N_11126);
xnor U11311 (N_11311,N_11182,N_11193);
and U11312 (N_11312,N_11046,N_11091);
and U11313 (N_11313,N_11100,N_11196);
xor U11314 (N_11314,N_11078,N_11188);
xnor U11315 (N_11315,N_11034,N_11096);
or U11316 (N_11316,N_11008,N_11163);
nor U11317 (N_11317,N_11038,N_11130);
nand U11318 (N_11318,N_11051,N_11023);
or U11319 (N_11319,N_11166,N_11126);
nor U11320 (N_11320,N_11005,N_11009);
or U11321 (N_11321,N_11189,N_11190);
or U11322 (N_11322,N_11088,N_11130);
nor U11323 (N_11323,N_11064,N_11146);
xor U11324 (N_11324,N_11128,N_11187);
or U11325 (N_11325,N_11000,N_11155);
nand U11326 (N_11326,N_11173,N_11074);
or U11327 (N_11327,N_11162,N_11125);
xor U11328 (N_11328,N_11103,N_11181);
or U11329 (N_11329,N_11042,N_11044);
xnor U11330 (N_11330,N_11183,N_11129);
or U11331 (N_11331,N_11041,N_11056);
or U11332 (N_11332,N_11020,N_11016);
or U11333 (N_11333,N_11196,N_11040);
or U11334 (N_11334,N_11123,N_11188);
and U11335 (N_11335,N_11128,N_11037);
or U11336 (N_11336,N_11104,N_11139);
or U11337 (N_11337,N_11169,N_11098);
xor U11338 (N_11338,N_11099,N_11024);
nand U11339 (N_11339,N_11142,N_11196);
nor U11340 (N_11340,N_11193,N_11188);
nor U11341 (N_11341,N_11087,N_11106);
nor U11342 (N_11342,N_11003,N_11084);
nor U11343 (N_11343,N_11185,N_11152);
nand U11344 (N_11344,N_11189,N_11076);
nand U11345 (N_11345,N_11122,N_11019);
and U11346 (N_11346,N_11153,N_11148);
and U11347 (N_11347,N_11065,N_11069);
and U11348 (N_11348,N_11113,N_11128);
nand U11349 (N_11349,N_11115,N_11076);
nand U11350 (N_11350,N_11103,N_11136);
and U11351 (N_11351,N_11187,N_11084);
nor U11352 (N_11352,N_11184,N_11090);
nand U11353 (N_11353,N_11133,N_11140);
or U11354 (N_11354,N_11016,N_11004);
xnor U11355 (N_11355,N_11094,N_11123);
or U11356 (N_11356,N_11006,N_11111);
nor U11357 (N_11357,N_11089,N_11041);
or U11358 (N_11358,N_11175,N_11095);
nand U11359 (N_11359,N_11169,N_11039);
nand U11360 (N_11360,N_11190,N_11125);
or U11361 (N_11361,N_11188,N_11199);
nand U11362 (N_11362,N_11194,N_11179);
xnor U11363 (N_11363,N_11129,N_11192);
nor U11364 (N_11364,N_11040,N_11049);
nor U11365 (N_11365,N_11089,N_11028);
xor U11366 (N_11366,N_11008,N_11095);
or U11367 (N_11367,N_11086,N_11048);
nor U11368 (N_11368,N_11121,N_11019);
nand U11369 (N_11369,N_11142,N_11104);
nor U11370 (N_11370,N_11021,N_11000);
or U11371 (N_11371,N_11138,N_11194);
or U11372 (N_11372,N_11148,N_11149);
nand U11373 (N_11373,N_11090,N_11039);
nand U11374 (N_11374,N_11137,N_11048);
nor U11375 (N_11375,N_11150,N_11073);
nand U11376 (N_11376,N_11149,N_11139);
nand U11377 (N_11377,N_11171,N_11109);
and U11378 (N_11378,N_11173,N_11142);
and U11379 (N_11379,N_11186,N_11153);
or U11380 (N_11380,N_11182,N_11159);
nand U11381 (N_11381,N_11195,N_11168);
xnor U11382 (N_11382,N_11170,N_11125);
nor U11383 (N_11383,N_11198,N_11135);
nand U11384 (N_11384,N_11048,N_11176);
or U11385 (N_11385,N_11089,N_11100);
xnor U11386 (N_11386,N_11142,N_11091);
or U11387 (N_11387,N_11013,N_11041);
xnor U11388 (N_11388,N_11097,N_11039);
nand U11389 (N_11389,N_11150,N_11052);
nor U11390 (N_11390,N_11177,N_11174);
xnor U11391 (N_11391,N_11130,N_11036);
xnor U11392 (N_11392,N_11076,N_11057);
nor U11393 (N_11393,N_11114,N_11015);
and U11394 (N_11394,N_11182,N_11151);
xor U11395 (N_11395,N_11050,N_11070);
nor U11396 (N_11396,N_11195,N_11130);
nor U11397 (N_11397,N_11021,N_11127);
nor U11398 (N_11398,N_11000,N_11121);
and U11399 (N_11399,N_11062,N_11152);
xnor U11400 (N_11400,N_11283,N_11353);
nand U11401 (N_11401,N_11364,N_11248);
nor U11402 (N_11402,N_11337,N_11201);
and U11403 (N_11403,N_11340,N_11384);
xor U11404 (N_11404,N_11275,N_11318);
xor U11405 (N_11405,N_11385,N_11391);
and U11406 (N_11406,N_11257,N_11269);
nor U11407 (N_11407,N_11284,N_11222);
nor U11408 (N_11408,N_11224,N_11276);
or U11409 (N_11409,N_11311,N_11388);
nor U11410 (N_11410,N_11328,N_11220);
or U11411 (N_11411,N_11301,N_11254);
xnor U11412 (N_11412,N_11300,N_11377);
and U11413 (N_11413,N_11305,N_11249);
and U11414 (N_11414,N_11374,N_11346);
xor U11415 (N_11415,N_11329,N_11314);
nor U11416 (N_11416,N_11218,N_11237);
and U11417 (N_11417,N_11217,N_11270);
xnor U11418 (N_11418,N_11280,N_11351);
and U11419 (N_11419,N_11345,N_11312);
xnor U11420 (N_11420,N_11332,N_11245);
xnor U11421 (N_11421,N_11211,N_11371);
nand U11422 (N_11422,N_11278,N_11358);
xor U11423 (N_11423,N_11227,N_11341);
xnor U11424 (N_11424,N_11365,N_11297);
or U11425 (N_11425,N_11212,N_11376);
xor U11426 (N_11426,N_11336,N_11285);
and U11427 (N_11427,N_11363,N_11286);
nand U11428 (N_11428,N_11348,N_11251);
nor U11429 (N_11429,N_11309,N_11206);
nand U11430 (N_11430,N_11308,N_11261);
or U11431 (N_11431,N_11343,N_11277);
xnor U11432 (N_11432,N_11317,N_11321);
xor U11433 (N_11433,N_11272,N_11273);
nor U11434 (N_11434,N_11387,N_11253);
and U11435 (N_11435,N_11294,N_11350);
or U11436 (N_11436,N_11303,N_11219);
and U11437 (N_11437,N_11356,N_11307);
xnor U11438 (N_11438,N_11203,N_11306);
and U11439 (N_11439,N_11247,N_11352);
or U11440 (N_11440,N_11240,N_11349);
or U11441 (N_11441,N_11373,N_11271);
or U11442 (N_11442,N_11221,N_11234);
or U11443 (N_11443,N_11210,N_11357);
or U11444 (N_11444,N_11265,N_11209);
and U11445 (N_11445,N_11204,N_11231);
and U11446 (N_11446,N_11292,N_11327);
xor U11447 (N_11447,N_11389,N_11287);
nor U11448 (N_11448,N_11255,N_11347);
nand U11449 (N_11449,N_11200,N_11335);
or U11450 (N_11450,N_11323,N_11302);
and U11451 (N_11451,N_11394,N_11208);
nor U11452 (N_11452,N_11214,N_11263);
xor U11453 (N_11453,N_11225,N_11246);
or U11454 (N_11454,N_11291,N_11322);
and U11455 (N_11455,N_11393,N_11370);
nand U11456 (N_11456,N_11315,N_11250);
nor U11457 (N_11457,N_11252,N_11216);
nand U11458 (N_11458,N_11354,N_11330);
or U11459 (N_11459,N_11397,N_11367);
xnor U11460 (N_11460,N_11360,N_11230);
nor U11461 (N_11461,N_11372,N_11238);
xnor U11462 (N_11462,N_11264,N_11399);
nand U11463 (N_11463,N_11375,N_11256);
nand U11464 (N_11464,N_11266,N_11205);
nor U11465 (N_11465,N_11244,N_11344);
or U11466 (N_11466,N_11369,N_11299);
nand U11467 (N_11467,N_11362,N_11355);
nor U11468 (N_11468,N_11223,N_11368);
and U11469 (N_11469,N_11268,N_11331);
nand U11470 (N_11470,N_11282,N_11281);
xnor U11471 (N_11471,N_11274,N_11279);
nor U11472 (N_11472,N_11359,N_11235);
or U11473 (N_11473,N_11324,N_11380);
nor U11474 (N_11474,N_11334,N_11293);
xor U11475 (N_11475,N_11361,N_11242);
xor U11476 (N_11476,N_11239,N_11383);
xor U11477 (N_11477,N_11288,N_11241);
nor U11478 (N_11478,N_11326,N_11366);
nor U11479 (N_11479,N_11298,N_11207);
nor U11480 (N_11480,N_11313,N_11316);
xor U11481 (N_11481,N_11333,N_11392);
nor U11482 (N_11482,N_11226,N_11396);
nor U11483 (N_11483,N_11296,N_11382);
nand U11484 (N_11484,N_11325,N_11228);
nor U11485 (N_11485,N_11378,N_11379);
nor U11486 (N_11486,N_11342,N_11229);
or U11487 (N_11487,N_11319,N_11258);
nand U11488 (N_11488,N_11215,N_11202);
nand U11489 (N_11489,N_11338,N_11213);
and U11490 (N_11490,N_11295,N_11320);
xor U11491 (N_11491,N_11289,N_11310);
xor U11492 (N_11492,N_11386,N_11339);
nand U11493 (N_11493,N_11290,N_11232);
and U11494 (N_11494,N_11304,N_11398);
nand U11495 (N_11495,N_11262,N_11233);
or U11496 (N_11496,N_11395,N_11260);
nor U11497 (N_11497,N_11236,N_11243);
nor U11498 (N_11498,N_11390,N_11381);
nand U11499 (N_11499,N_11259,N_11267);
nor U11500 (N_11500,N_11386,N_11240);
or U11501 (N_11501,N_11345,N_11375);
or U11502 (N_11502,N_11271,N_11278);
nand U11503 (N_11503,N_11295,N_11213);
nand U11504 (N_11504,N_11289,N_11365);
nand U11505 (N_11505,N_11389,N_11398);
and U11506 (N_11506,N_11393,N_11318);
nor U11507 (N_11507,N_11282,N_11333);
or U11508 (N_11508,N_11324,N_11260);
or U11509 (N_11509,N_11357,N_11391);
nand U11510 (N_11510,N_11399,N_11281);
xnor U11511 (N_11511,N_11369,N_11202);
xnor U11512 (N_11512,N_11373,N_11242);
xnor U11513 (N_11513,N_11305,N_11369);
or U11514 (N_11514,N_11325,N_11233);
or U11515 (N_11515,N_11352,N_11308);
xor U11516 (N_11516,N_11321,N_11231);
nand U11517 (N_11517,N_11333,N_11349);
or U11518 (N_11518,N_11320,N_11273);
xor U11519 (N_11519,N_11283,N_11392);
nor U11520 (N_11520,N_11372,N_11260);
nor U11521 (N_11521,N_11272,N_11200);
and U11522 (N_11522,N_11243,N_11216);
and U11523 (N_11523,N_11296,N_11249);
and U11524 (N_11524,N_11203,N_11391);
and U11525 (N_11525,N_11237,N_11315);
or U11526 (N_11526,N_11393,N_11233);
xnor U11527 (N_11527,N_11295,N_11315);
nand U11528 (N_11528,N_11371,N_11376);
nor U11529 (N_11529,N_11327,N_11372);
or U11530 (N_11530,N_11277,N_11349);
or U11531 (N_11531,N_11276,N_11282);
or U11532 (N_11532,N_11350,N_11244);
nor U11533 (N_11533,N_11220,N_11284);
or U11534 (N_11534,N_11287,N_11289);
or U11535 (N_11535,N_11284,N_11260);
nand U11536 (N_11536,N_11257,N_11383);
xor U11537 (N_11537,N_11222,N_11294);
nor U11538 (N_11538,N_11366,N_11346);
and U11539 (N_11539,N_11387,N_11270);
and U11540 (N_11540,N_11337,N_11231);
or U11541 (N_11541,N_11309,N_11343);
or U11542 (N_11542,N_11354,N_11226);
xnor U11543 (N_11543,N_11384,N_11241);
and U11544 (N_11544,N_11256,N_11206);
nor U11545 (N_11545,N_11379,N_11236);
and U11546 (N_11546,N_11207,N_11275);
nand U11547 (N_11547,N_11201,N_11208);
and U11548 (N_11548,N_11237,N_11253);
or U11549 (N_11549,N_11337,N_11381);
nor U11550 (N_11550,N_11239,N_11350);
xor U11551 (N_11551,N_11384,N_11363);
and U11552 (N_11552,N_11298,N_11284);
nand U11553 (N_11553,N_11327,N_11307);
or U11554 (N_11554,N_11254,N_11221);
xor U11555 (N_11555,N_11224,N_11262);
nand U11556 (N_11556,N_11251,N_11244);
xor U11557 (N_11557,N_11319,N_11375);
nor U11558 (N_11558,N_11367,N_11324);
nor U11559 (N_11559,N_11202,N_11268);
and U11560 (N_11560,N_11275,N_11356);
or U11561 (N_11561,N_11366,N_11242);
nor U11562 (N_11562,N_11379,N_11227);
xor U11563 (N_11563,N_11286,N_11295);
xnor U11564 (N_11564,N_11225,N_11316);
or U11565 (N_11565,N_11226,N_11281);
nand U11566 (N_11566,N_11244,N_11259);
nand U11567 (N_11567,N_11258,N_11219);
xor U11568 (N_11568,N_11293,N_11312);
nor U11569 (N_11569,N_11357,N_11209);
or U11570 (N_11570,N_11389,N_11339);
nand U11571 (N_11571,N_11341,N_11252);
and U11572 (N_11572,N_11319,N_11394);
nor U11573 (N_11573,N_11313,N_11261);
nand U11574 (N_11574,N_11356,N_11214);
or U11575 (N_11575,N_11301,N_11212);
nand U11576 (N_11576,N_11382,N_11323);
xnor U11577 (N_11577,N_11221,N_11204);
and U11578 (N_11578,N_11399,N_11326);
nor U11579 (N_11579,N_11288,N_11203);
nor U11580 (N_11580,N_11251,N_11322);
and U11581 (N_11581,N_11351,N_11219);
nor U11582 (N_11582,N_11329,N_11330);
and U11583 (N_11583,N_11300,N_11372);
nor U11584 (N_11584,N_11374,N_11315);
or U11585 (N_11585,N_11225,N_11249);
xor U11586 (N_11586,N_11359,N_11201);
or U11587 (N_11587,N_11261,N_11373);
or U11588 (N_11588,N_11257,N_11302);
or U11589 (N_11589,N_11372,N_11352);
and U11590 (N_11590,N_11273,N_11378);
or U11591 (N_11591,N_11343,N_11237);
xnor U11592 (N_11592,N_11375,N_11309);
and U11593 (N_11593,N_11385,N_11314);
nand U11594 (N_11594,N_11252,N_11389);
xor U11595 (N_11595,N_11396,N_11219);
and U11596 (N_11596,N_11392,N_11251);
or U11597 (N_11597,N_11384,N_11301);
xor U11598 (N_11598,N_11278,N_11353);
nor U11599 (N_11599,N_11269,N_11253);
nand U11600 (N_11600,N_11417,N_11493);
and U11601 (N_11601,N_11535,N_11447);
nand U11602 (N_11602,N_11555,N_11483);
and U11603 (N_11603,N_11484,N_11542);
xnor U11604 (N_11604,N_11440,N_11441);
xnor U11605 (N_11605,N_11463,N_11402);
and U11606 (N_11606,N_11582,N_11599);
and U11607 (N_11607,N_11517,N_11414);
xnor U11608 (N_11608,N_11587,N_11504);
nor U11609 (N_11609,N_11506,N_11468);
nand U11610 (N_11610,N_11435,N_11460);
xnor U11611 (N_11611,N_11481,N_11411);
nand U11612 (N_11612,N_11586,N_11433);
nor U11613 (N_11613,N_11462,N_11475);
xor U11614 (N_11614,N_11561,N_11482);
xnor U11615 (N_11615,N_11540,N_11422);
nand U11616 (N_11616,N_11522,N_11449);
and U11617 (N_11617,N_11568,N_11434);
or U11618 (N_11618,N_11425,N_11486);
xnor U11619 (N_11619,N_11472,N_11490);
nor U11620 (N_11620,N_11569,N_11471);
nand U11621 (N_11621,N_11442,N_11461);
or U11622 (N_11622,N_11576,N_11458);
xnor U11623 (N_11623,N_11403,N_11562);
xor U11624 (N_11624,N_11480,N_11575);
nor U11625 (N_11625,N_11456,N_11531);
nor U11626 (N_11626,N_11571,N_11572);
xor U11627 (N_11627,N_11554,N_11598);
and U11628 (N_11628,N_11501,N_11439);
xor U11629 (N_11629,N_11583,N_11548);
nor U11630 (N_11630,N_11436,N_11426);
nor U11631 (N_11631,N_11451,N_11512);
xor U11632 (N_11632,N_11528,N_11541);
and U11633 (N_11633,N_11450,N_11574);
nor U11634 (N_11634,N_11525,N_11401);
nand U11635 (N_11635,N_11419,N_11565);
nor U11636 (N_11636,N_11534,N_11563);
and U11637 (N_11637,N_11487,N_11592);
and U11638 (N_11638,N_11597,N_11552);
or U11639 (N_11639,N_11473,N_11577);
xor U11640 (N_11640,N_11416,N_11474);
nand U11641 (N_11641,N_11438,N_11524);
xor U11642 (N_11642,N_11467,N_11537);
xor U11643 (N_11643,N_11544,N_11500);
nand U11644 (N_11644,N_11545,N_11551);
xor U11645 (N_11645,N_11459,N_11591);
xor U11646 (N_11646,N_11497,N_11594);
xor U11647 (N_11647,N_11520,N_11590);
nor U11648 (N_11648,N_11432,N_11503);
xnor U11649 (N_11649,N_11408,N_11530);
nand U11650 (N_11650,N_11496,N_11515);
or U11651 (N_11651,N_11557,N_11498);
xnor U11652 (N_11652,N_11499,N_11404);
or U11653 (N_11653,N_11469,N_11412);
nand U11654 (N_11654,N_11550,N_11448);
or U11655 (N_11655,N_11585,N_11532);
or U11656 (N_11656,N_11479,N_11464);
or U11657 (N_11657,N_11477,N_11521);
nor U11658 (N_11658,N_11478,N_11547);
nor U11659 (N_11659,N_11589,N_11507);
nand U11660 (N_11660,N_11445,N_11579);
and U11661 (N_11661,N_11409,N_11424);
and U11662 (N_11662,N_11457,N_11446);
or U11663 (N_11663,N_11470,N_11526);
xnor U11664 (N_11664,N_11529,N_11533);
nor U11665 (N_11665,N_11553,N_11508);
xor U11666 (N_11666,N_11514,N_11431);
or U11667 (N_11667,N_11567,N_11410);
nor U11668 (N_11668,N_11420,N_11581);
nand U11669 (N_11669,N_11538,N_11418);
nor U11670 (N_11670,N_11427,N_11564);
xor U11671 (N_11671,N_11546,N_11465);
or U11672 (N_11672,N_11489,N_11492);
nand U11673 (N_11673,N_11406,N_11556);
nand U11674 (N_11674,N_11573,N_11516);
xnor U11675 (N_11675,N_11518,N_11527);
xor U11676 (N_11676,N_11566,N_11536);
nor U11677 (N_11677,N_11519,N_11570);
or U11678 (N_11678,N_11588,N_11491);
nor U11679 (N_11679,N_11495,N_11596);
nand U11680 (N_11680,N_11454,N_11452);
and U11681 (N_11681,N_11549,N_11421);
or U11682 (N_11682,N_11488,N_11415);
and U11683 (N_11683,N_11580,N_11558);
xor U11684 (N_11684,N_11510,N_11578);
nand U11685 (N_11685,N_11485,N_11523);
nor U11686 (N_11686,N_11429,N_11466);
or U11687 (N_11687,N_11444,N_11511);
or U11688 (N_11688,N_11584,N_11593);
or U11689 (N_11689,N_11423,N_11455);
nand U11690 (N_11690,N_11437,N_11560);
and U11691 (N_11691,N_11428,N_11494);
or U11692 (N_11692,N_11400,N_11513);
or U11693 (N_11693,N_11505,N_11509);
xor U11694 (N_11694,N_11502,N_11430);
and U11695 (N_11695,N_11543,N_11476);
or U11696 (N_11696,N_11559,N_11405);
nand U11697 (N_11697,N_11539,N_11413);
nand U11698 (N_11698,N_11443,N_11407);
nor U11699 (N_11699,N_11453,N_11595);
nor U11700 (N_11700,N_11481,N_11499);
and U11701 (N_11701,N_11449,N_11483);
xnor U11702 (N_11702,N_11490,N_11530);
or U11703 (N_11703,N_11471,N_11472);
and U11704 (N_11704,N_11400,N_11569);
nand U11705 (N_11705,N_11585,N_11492);
or U11706 (N_11706,N_11473,N_11509);
nand U11707 (N_11707,N_11599,N_11580);
or U11708 (N_11708,N_11548,N_11434);
and U11709 (N_11709,N_11457,N_11415);
nand U11710 (N_11710,N_11505,N_11502);
nand U11711 (N_11711,N_11559,N_11586);
xor U11712 (N_11712,N_11506,N_11536);
xnor U11713 (N_11713,N_11521,N_11519);
nor U11714 (N_11714,N_11425,N_11574);
xnor U11715 (N_11715,N_11508,N_11402);
nor U11716 (N_11716,N_11510,N_11545);
nor U11717 (N_11717,N_11473,N_11576);
nor U11718 (N_11718,N_11561,N_11440);
nor U11719 (N_11719,N_11556,N_11506);
nor U11720 (N_11720,N_11407,N_11583);
nor U11721 (N_11721,N_11405,N_11498);
and U11722 (N_11722,N_11554,N_11555);
nor U11723 (N_11723,N_11554,N_11575);
or U11724 (N_11724,N_11577,N_11446);
nand U11725 (N_11725,N_11411,N_11534);
nor U11726 (N_11726,N_11512,N_11561);
xnor U11727 (N_11727,N_11563,N_11544);
or U11728 (N_11728,N_11443,N_11576);
nor U11729 (N_11729,N_11460,N_11592);
nand U11730 (N_11730,N_11513,N_11557);
or U11731 (N_11731,N_11451,N_11478);
and U11732 (N_11732,N_11575,N_11427);
xor U11733 (N_11733,N_11453,N_11566);
and U11734 (N_11734,N_11400,N_11503);
xnor U11735 (N_11735,N_11541,N_11473);
or U11736 (N_11736,N_11594,N_11491);
xnor U11737 (N_11737,N_11533,N_11460);
and U11738 (N_11738,N_11547,N_11529);
xnor U11739 (N_11739,N_11538,N_11485);
nand U11740 (N_11740,N_11469,N_11581);
nand U11741 (N_11741,N_11532,N_11470);
nor U11742 (N_11742,N_11599,N_11475);
and U11743 (N_11743,N_11420,N_11563);
xor U11744 (N_11744,N_11487,N_11483);
and U11745 (N_11745,N_11443,N_11587);
xnor U11746 (N_11746,N_11486,N_11418);
nor U11747 (N_11747,N_11426,N_11401);
or U11748 (N_11748,N_11590,N_11422);
or U11749 (N_11749,N_11543,N_11581);
nand U11750 (N_11750,N_11528,N_11446);
nand U11751 (N_11751,N_11513,N_11434);
xor U11752 (N_11752,N_11405,N_11538);
xnor U11753 (N_11753,N_11489,N_11591);
or U11754 (N_11754,N_11558,N_11492);
xnor U11755 (N_11755,N_11417,N_11533);
nand U11756 (N_11756,N_11529,N_11460);
xnor U11757 (N_11757,N_11511,N_11474);
and U11758 (N_11758,N_11541,N_11420);
nand U11759 (N_11759,N_11442,N_11574);
nor U11760 (N_11760,N_11588,N_11553);
and U11761 (N_11761,N_11497,N_11534);
nor U11762 (N_11762,N_11555,N_11567);
nand U11763 (N_11763,N_11509,N_11496);
nor U11764 (N_11764,N_11521,N_11475);
and U11765 (N_11765,N_11459,N_11587);
nor U11766 (N_11766,N_11472,N_11580);
and U11767 (N_11767,N_11565,N_11524);
xor U11768 (N_11768,N_11458,N_11523);
nand U11769 (N_11769,N_11509,N_11493);
and U11770 (N_11770,N_11551,N_11403);
xor U11771 (N_11771,N_11578,N_11574);
nand U11772 (N_11772,N_11413,N_11443);
nand U11773 (N_11773,N_11451,N_11502);
nor U11774 (N_11774,N_11467,N_11501);
or U11775 (N_11775,N_11401,N_11555);
and U11776 (N_11776,N_11408,N_11499);
xor U11777 (N_11777,N_11440,N_11562);
or U11778 (N_11778,N_11435,N_11451);
and U11779 (N_11779,N_11462,N_11548);
nor U11780 (N_11780,N_11579,N_11524);
nor U11781 (N_11781,N_11572,N_11511);
nor U11782 (N_11782,N_11418,N_11592);
or U11783 (N_11783,N_11433,N_11454);
nor U11784 (N_11784,N_11595,N_11418);
or U11785 (N_11785,N_11460,N_11572);
nor U11786 (N_11786,N_11408,N_11585);
or U11787 (N_11787,N_11584,N_11500);
xnor U11788 (N_11788,N_11562,N_11531);
nand U11789 (N_11789,N_11482,N_11411);
or U11790 (N_11790,N_11597,N_11531);
or U11791 (N_11791,N_11534,N_11504);
or U11792 (N_11792,N_11403,N_11496);
nand U11793 (N_11793,N_11410,N_11413);
nor U11794 (N_11794,N_11520,N_11420);
nor U11795 (N_11795,N_11528,N_11449);
nor U11796 (N_11796,N_11574,N_11466);
or U11797 (N_11797,N_11574,N_11502);
xor U11798 (N_11798,N_11539,N_11584);
and U11799 (N_11799,N_11563,N_11467);
xor U11800 (N_11800,N_11625,N_11719);
nand U11801 (N_11801,N_11658,N_11712);
nand U11802 (N_11802,N_11656,N_11709);
xnor U11803 (N_11803,N_11617,N_11711);
nor U11804 (N_11804,N_11665,N_11681);
nand U11805 (N_11805,N_11687,N_11798);
and U11806 (N_11806,N_11660,N_11771);
and U11807 (N_11807,N_11701,N_11782);
or U11808 (N_11808,N_11764,N_11708);
or U11809 (N_11809,N_11723,N_11653);
or U11810 (N_11810,N_11671,N_11763);
and U11811 (N_11811,N_11794,N_11652);
nand U11812 (N_11812,N_11759,N_11788);
or U11813 (N_11813,N_11781,N_11715);
nand U11814 (N_11814,N_11699,N_11783);
xor U11815 (N_11815,N_11669,N_11655);
and U11816 (N_11816,N_11734,N_11741);
or U11817 (N_11817,N_11694,N_11647);
nor U11818 (N_11818,N_11608,N_11718);
and U11819 (N_11819,N_11722,N_11620);
xor U11820 (N_11820,N_11789,N_11686);
and U11821 (N_11821,N_11720,N_11728);
or U11822 (N_11822,N_11676,N_11683);
nand U11823 (N_11823,N_11744,N_11774);
xnor U11824 (N_11824,N_11677,N_11706);
nor U11825 (N_11825,N_11614,N_11631);
xor U11826 (N_11826,N_11639,N_11606);
nor U11827 (N_11827,N_11662,N_11746);
or U11828 (N_11828,N_11799,N_11635);
xor U11829 (N_11829,N_11648,N_11766);
nand U11830 (N_11830,N_11700,N_11748);
xnor U11831 (N_11831,N_11650,N_11791);
and U11832 (N_11832,N_11775,N_11679);
or U11833 (N_11833,N_11634,N_11772);
xor U11834 (N_11834,N_11790,N_11754);
xor U11835 (N_11835,N_11616,N_11695);
or U11836 (N_11836,N_11736,N_11738);
and U11837 (N_11837,N_11601,N_11777);
nor U11838 (N_11838,N_11664,N_11675);
or U11839 (N_11839,N_11666,N_11716);
or U11840 (N_11840,N_11770,N_11795);
nor U11841 (N_11841,N_11621,N_11640);
and U11842 (N_11842,N_11613,N_11615);
nand U11843 (N_11843,N_11690,N_11727);
nand U11844 (N_11844,N_11678,N_11619);
xnor U11845 (N_11845,N_11724,N_11729);
and U11846 (N_11846,N_11731,N_11630);
nand U11847 (N_11847,N_11644,N_11604);
or U11848 (N_11848,N_11760,N_11674);
or U11849 (N_11849,N_11735,N_11793);
xor U11850 (N_11850,N_11638,N_11673);
nor U11851 (N_11851,N_11628,N_11624);
or U11852 (N_11852,N_11663,N_11607);
xor U11853 (N_11853,N_11784,N_11717);
and U11854 (N_11854,N_11626,N_11762);
and U11855 (N_11855,N_11618,N_11725);
nor U11856 (N_11856,N_11726,N_11642);
or U11857 (N_11857,N_11761,N_11713);
nor U11858 (N_11858,N_11750,N_11749);
or U11859 (N_11859,N_11751,N_11691);
or U11860 (N_11860,N_11636,N_11797);
nand U11861 (N_11861,N_11767,N_11792);
xor U11862 (N_11862,N_11629,N_11747);
and U11863 (N_11863,N_11769,N_11609);
and U11864 (N_11864,N_11633,N_11742);
or U11865 (N_11865,N_11623,N_11646);
or U11866 (N_11866,N_11680,N_11707);
or U11867 (N_11867,N_11600,N_11670);
and U11868 (N_11868,N_11697,N_11737);
nor U11869 (N_11869,N_11704,N_11649);
and U11870 (N_11870,N_11721,N_11796);
and U11871 (N_11871,N_11661,N_11732);
xor U11872 (N_11872,N_11710,N_11672);
nor U11873 (N_11873,N_11730,N_11705);
nand U11874 (N_11874,N_11692,N_11756);
nor U11875 (N_11875,N_11645,N_11698);
and U11876 (N_11876,N_11702,N_11602);
nand U11877 (N_11877,N_11776,N_11780);
nor U11878 (N_11878,N_11714,N_11752);
xnor U11879 (N_11879,N_11622,N_11657);
or U11880 (N_11880,N_11693,N_11632);
or U11881 (N_11881,N_11753,N_11740);
and U11882 (N_11882,N_11733,N_11641);
nand U11883 (N_11883,N_11745,N_11605);
nor U11884 (N_11884,N_11685,N_11703);
xnor U11885 (N_11885,N_11758,N_11659);
nor U11886 (N_11886,N_11787,N_11643);
xor U11887 (N_11887,N_11773,N_11757);
or U11888 (N_11888,N_11603,N_11689);
nand U11889 (N_11889,N_11637,N_11779);
nand U11890 (N_11890,N_11682,N_11765);
nand U11891 (N_11891,N_11610,N_11786);
nand U11892 (N_11892,N_11612,N_11668);
nand U11893 (N_11893,N_11688,N_11755);
or U11894 (N_11894,N_11696,N_11739);
nand U11895 (N_11895,N_11768,N_11627);
nor U11896 (N_11896,N_11778,N_11667);
and U11897 (N_11897,N_11651,N_11654);
nor U11898 (N_11898,N_11684,N_11611);
and U11899 (N_11899,N_11743,N_11785);
xor U11900 (N_11900,N_11623,N_11687);
nor U11901 (N_11901,N_11677,N_11739);
nand U11902 (N_11902,N_11761,N_11744);
xnor U11903 (N_11903,N_11784,N_11751);
and U11904 (N_11904,N_11785,N_11792);
nand U11905 (N_11905,N_11653,N_11684);
nand U11906 (N_11906,N_11635,N_11730);
and U11907 (N_11907,N_11733,N_11644);
nor U11908 (N_11908,N_11658,N_11652);
and U11909 (N_11909,N_11653,N_11668);
xnor U11910 (N_11910,N_11629,N_11642);
nand U11911 (N_11911,N_11713,N_11700);
nand U11912 (N_11912,N_11649,N_11740);
nand U11913 (N_11913,N_11610,N_11760);
and U11914 (N_11914,N_11612,N_11795);
and U11915 (N_11915,N_11679,N_11697);
nand U11916 (N_11916,N_11688,N_11662);
or U11917 (N_11917,N_11611,N_11632);
or U11918 (N_11918,N_11783,N_11787);
or U11919 (N_11919,N_11625,N_11630);
xor U11920 (N_11920,N_11775,N_11672);
and U11921 (N_11921,N_11605,N_11725);
and U11922 (N_11922,N_11682,N_11766);
xor U11923 (N_11923,N_11622,N_11642);
nor U11924 (N_11924,N_11680,N_11742);
nor U11925 (N_11925,N_11665,N_11642);
or U11926 (N_11926,N_11696,N_11744);
and U11927 (N_11927,N_11671,N_11773);
xnor U11928 (N_11928,N_11744,N_11777);
xnor U11929 (N_11929,N_11641,N_11742);
or U11930 (N_11930,N_11716,N_11682);
nand U11931 (N_11931,N_11601,N_11609);
and U11932 (N_11932,N_11746,N_11638);
nand U11933 (N_11933,N_11683,N_11708);
nand U11934 (N_11934,N_11707,N_11742);
xnor U11935 (N_11935,N_11796,N_11675);
nor U11936 (N_11936,N_11618,N_11799);
nand U11937 (N_11937,N_11621,N_11795);
and U11938 (N_11938,N_11722,N_11716);
or U11939 (N_11939,N_11639,N_11764);
nor U11940 (N_11940,N_11756,N_11780);
nor U11941 (N_11941,N_11672,N_11652);
nor U11942 (N_11942,N_11769,N_11790);
and U11943 (N_11943,N_11693,N_11791);
nor U11944 (N_11944,N_11709,N_11757);
and U11945 (N_11945,N_11647,N_11734);
nor U11946 (N_11946,N_11683,N_11726);
nand U11947 (N_11947,N_11682,N_11733);
and U11948 (N_11948,N_11783,N_11754);
and U11949 (N_11949,N_11700,N_11655);
xor U11950 (N_11950,N_11727,N_11780);
xnor U11951 (N_11951,N_11752,N_11701);
nand U11952 (N_11952,N_11708,N_11613);
xor U11953 (N_11953,N_11736,N_11623);
nor U11954 (N_11954,N_11651,N_11630);
nor U11955 (N_11955,N_11689,N_11736);
nor U11956 (N_11956,N_11794,N_11651);
xor U11957 (N_11957,N_11737,N_11650);
or U11958 (N_11958,N_11768,N_11764);
nand U11959 (N_11959,N_11617,N_11730);
or U11960 (N_11960,N_11797,N_11616);
nor U11961 (N_11961,N_11637,N_11602);
nand U11962 (N_11962,N_11777,N_11673);
and U11963 (N_11963,N_11619,N_11659);
and U11964 (N_11964,N_11630,N_11648);
xor U11965 (N_11965,N_11786,N_11648);
and U11966 (N_11966,N_11740,N_11659);
and U11967 (N_11967,N_11659,N_11759);
or U11968 (N_11968,N_11687,N_11711);
and U11969 (N_11969,N_11797,N_11659);
or U11970 (N_11970,N_11636,N_11640);
nand U11971 (N_11971,N_11797,N_11795);
and U11972 (N_11972,N_11789,N_11724);
xnor U11973 (N_11973,N_11602,N_11789);
and U11974 (N_11974,N_11670,N_11734);
nand U11975 (N_11975,N_11763,N_11786);
nand U11976 (N_11976,N_11743,N_11697);
or U11977 (N_11977,N_11665,N_11679);
and U11978 (N_11978,N_11702,N_11785);
or U11979 (N_11979,N_11660,N_11683);
or U11980 (N_11980,N_11617,N_11793);
and U11981 (N_11981,N_11646,N_11733);
and U11982 (N_11982,N_11779,N_11787);
and U11983 (N_11983,N_11629,N_11792);
and U11984 (N_11984,N_11783,N_11789);
nand U11985 (N_11985,N_11651,N_11754);
nand U11986 (N_11986,N_11756,N_11784);
or U11987 (N_11987,N_11708,N_11654);
or U11988 (N_11988,N_11708,N_11727);
nand U11989 (N_11989,N_11696,N_11771);
xnor U11990 (N_11990,N_11782,N_11762);
xnor U11991 (N_11991,N_11614,N_11703);
nor U11992 (N_11992,N_11763,N_11622);
nor U11993 (N_11993,N_11689,N_11625);
xnor U11994 (N_11994,N_11759,N_11656);
or U11995 (N_11995,N_11766,N_11730);
or U11996 (N_11996,N_11753,N_11710);
nand U11997 (N_11997,N_11795,N_11630);
nand U11998 (N_11998,N_11768,N_11736);
or U11999 (N_11999,N_11609,N_11694);
and U12000 (N_12000,N_11885,N_11862);
xor U12001 (N_12001,N_11854,N_11838);
nand U12002 (N_12002,N_11959,N_11839);
or U12003 (N_12003,N_11999,N_11895);
nor U12004 (N_12004,N_11948,N_11971);
nand U12005 (N_12005,N_11863,N_11917);
nor U12006 (N_12006,N_11932,N_11820);
nand U12007 (N_12007,N_11991,N_11855);
nand U12008 (N_12008,N_11870,N_11931);
xor U12009 (N_12009,N_11918,N_11802);
nor U12010 (N_12010,N_11837,N_11925);
or U12011 (N_12011,N_11850,N_11866);
nand U12012 (N_12012,N_11849,N_11842);
xor U12013 (N_12013,N_11894,N_11889);
nand U12014 (N_12014,N_11886,N_11983);
nand U12015 (N_12015,N_11934,N_11800);
or U12016 (N_12016,N_11815,N_11804);
xor U12017 (N_12017,N_11969,N_11845);
xor U12018 (N_12018,N_11919,N_11888);
nor U12019 (N_12019,N_11953,N_11909);
xor U12020 (N_12020,N_11887,N_11935);
nand U12021 (N_12021,N_11973,N_11806);
and U12022 (N_12022,N_11975,N_11989);
and U12023 (N_12023,N_11981,N_11957);
and U12024 (N_12024,N_11988,N_11883);
nand U12025 (N_12025,N_11924,N_11923);
nor U12026 (N_12026,N_11902,N_11961);
and U12027 (N_12027,N_11930,N_11907);
nor U12028 (N_12028,N_11995,N_11891);
xor U12029 (N_12029,N_11821,N_11834);
xor U12030 (N_12030,N_11950,N_11805);
or U12031 (N_12031,N_11952,N_11828);
xnor U12032 (N_12032,N_11819,N_11979);
nand U12033 (N_12033,N_11847,N_11940);
xnor U12034 (N_12034,N_11899,N_11947);
nor U12035 (N_12035,N_11808,N_11914);
nand U12036 (N_12036,N_11915,N_11865);
nor U12037 (N_12037,N_11943,N_11916);
xnor U12038 (N_12038,N_11929,N_11853);
xnor U12039 (N_12039,N_11811,N_11985);
nor U12040 (N_12040,N_11910,N_11938);
and U12041 (N_12041,N_11872,N_11864);
nor U12042 (N_12042,N_11913,N_11968);
and U12043 (N_12043,N_11990,N_11951);
nor U12044 (N_12044,N_11927,N_11826);
xnor U12045 (N_12045,N_11976,N_11861);
and U12046 (N_12046,N_11807,N_11956);
xor U12047 (N_12047,N_11904,N_11936);
or U12048 (N_12048,N_11876,N_11949);
or U12049 (N_12049,N_11978,N_11986);
nor U12050 (N_12050,N_11884,N_11848);
nand U12051 (N_12051,N_11954,N_11997);
xor U12052 (N_12052,N_11896,N_11869);
xor U12053 (N_12053,N_11880,N_11830);
and U12054 (N_12054,N_11857,N_11825);
nand U12055 (N_12055,N_11814,N_11926);
nand U12056 (N_12056,N_11852,N_11882);
and U12057 (N_12057,N_11942,N_11960);
and U12058 (N_12058,N_11832,N_11875);
xnor U12059 (N_12059,N_11858,N_11900);
xnor U12060 (N_12060,N_11937,N_11977);
and U12061 (N_12061,N_11987,N_11881);
nand U12062 (N_12062,N_11836,N_11996);
and U12063 (N_12063,N_11809,N_11967);
xnor U12064 (N_12064,N_11812,N_11803);
nand U12065 (N_12065,N_11966,N_11972);
and U12066 (N_12066,N_11906,N_11851);
xor U12067 (N_12067,N_11958,N_11993);
nand U12068 (N_12068,N_11982,N_11903);
nand U12069 (N_12069,N_11817,N_11928);
nand U12070 (N_12070,N_11879,N_11874);
xor U12071 (N_12071,N_11898,N_11846);
nand U12072 (N_12072,N_11843,N_11871);
nand U12073 (N_12073,N_11827,N_11856);
or U12074 (N_12074,N_11939,N_11829);
and U12075 (N_12075,N_11860,N_11922);
xnor U12076 (N_12076,N_11908,N_11920);
nor U12077 (N_12077,N_11974,N_11810);
nor U12078 (N_12078,N_11962,N_11844);
or U12079 (N_12079,N_11941,N_11831);
nor U12080 (N_12080,N_11998,N_11893);
xor U12081 (N_12081,N_11801,N_11859);
and U12082 (N_12082,N_11873,N_11822);
nand U12083 (N_12083,N_11984,N_11877);
nor U12084 (N_12084,N_11933,N_11867);
nand U12085 (N_12085,N_11911,N_11992);
nor U12086 (N_12086,N_11868,N_11813);
and U12087 (N_12087,N_11841,N_11945);
and U12088 (N_12088,N_11816,N_11824);
and U12089 (N_12089,N_11835,N_11955);
and U12090 (N_12090,N_11921,N_11912);
nand U12091 (N_12091,N_11963,N_11892);
nor U12092 (N_12092,N_11994,N_11878);
and U12093 (N_12093,N_11897,N_11840);
nor U12094 (N_12094,N_11901,N_11905);
xnor U12095 (N_12095,N_11946,N_11818);
nor U12096 (N_12096,N_11823,N_11964);
nand U12097 (N_12097,N_11890,N_11965);
or U12098 (N_12098,N_11970,N_11980);
xor U12099 (N_12099,N_11833,N_11944);
nand U12100 (N_12100,N_11921,N_11989);
xor U12101 (N_12101,N_11804,N_11896);
xor U12102 (N_12102,N_11958,N_11994);
nand U12103 (N_12103,N_11958,N_11855);
nor U12104 (N_12104,N_11911,N_11873);
xnor U12105 (N_12105,N_11867,N_11903);
nand U12106 (N_12106,N_11848,N_11937);
or U12107 (N_12107,N_11866,N_11870);
and U12108 (N_12108,N_11932,N_11945);
xor U12109 (N_12109,N_11991,N_11865);
xnor U12110 (N_12110,N_11985,N_11909);
and U12111 (N_12111,N_11826,N_11963);
nand U12112 (N_12112,N_11833,N_11931);
nor U12113 (N_12113,N_11987,N_11891);
nand U12114 (N_12114,N_11923,N_11903);
or U12115 (N_12115,N_11962,N_11875);
nor U12116 (N_12116,N_11918,N_11866);
nand U12117 (N_12117,N_11804,N_11836);
nand U12118 (N_12118,N_11824,N_11940);
or U12119 (N_12119,N_11980,N_11874);
and U12120 (N_12120,N_11941,N_11870);
or U12121 (N_12121,N_11903,N_11871);
xor U12122 (N_12122,N_11871,N_11850);
or U12123 (N_12123,N_11930,N_11886);
nor U12124 (N_12124,N_11810,N_11899);
nor U12125 (N_12125,N_11895,N_11923);
and U12126 (N_12126,N_11820,N_11807);
xor U12127 (N_12127,N_11936,N_11909);
or U12128 (N_12128,N_11982,N_11895);
and U12129 (N_12129,N_11855,N_11972);
xor U12130 (N_12130,N_11919,N_11959);
and U12131 (N_12131,N_11828,N_11976);
nand U12132 (N_12132,N_11964,N_11992);
or U12133 (N_12133,N_11831,N_11837);
xnor U12134 (N_12134,N_11928,N_11814);
and U12135 (N_12135,N_11950,N_11809);
xnor U12136 (N_12136,N_11811,N_11913);
nand U12137 (N_12137,N_11992,N_11851);
or U12138 (N_12138,N_11807,N_11963);
or U12139 (N_12139,N_11996,N_11972);
or U12140 (N_12140,N_11876,N_11941);
or U12141 (N_12141,N_11885,N_11882);
and U12142 (N_12142,N_11836,N_11905);
nor U12143 (N_12143,N_11830,N_11857);
xor U12144 (N_12144,N_11834,N_11936);
nor U12145 (N_12145,N_11849,N_11912);
nand U12146 (N_12146,N_11909,N_11902);
or U12147 (N_12147,N_11810,N_11919);
nand U12148 (N_12148,N_11868,N_11866);
nor U12149 (N_12149,N_11858,N_11972);
or U12150 (N_12150,N_11921,N_11814);
and U12151 (N_12151,N_11801,N_11985);
xor U12152 (N_12152,N_11865,N_11957);
or U12153 (N_12153,N_11954,N_11941);
and U12154 (N_12154,N_11809,N_11989);
nor U12155 (N_12155,N_11959,N_11933);
and U12156 (N_12156,N_11891,N_11984);
or U12157 (N_12157,N_11885,N_11812);
and U12158 (N_12158,N_11927,N_11961);
or U12159 (N_12159,N_11862,N_11868);
xnor U12160 (N_12160,N_11916,N_11867);
xor U12161 (N_12161,N_11809,N_11858);
nand U12162 (N_12162,N_11889,N_11823);
nand U12163 (N_12163,N_11821,N_11885);
xnor U12164 (N_12164,N_11878,N_11904);
or U12165 (N_12165,N_11940,N_11878);
or U12166 (N_12166,N_11905,N_11923);
xnor U12167 (N_12167,N_11961,N_11911);
nor U12168 (N_12168,N_11954,N_11824);
nor U12169 (N_12169,N_11928,N_11995);
xor U12170 (N_12170,N_11968,N_11938);
xnor U12171 (N_12171,N_11813,N_11863);
or U12172 (N_12172,N_11913,N_11972);
or U12173 (N_12173,N_11892,N_11954);
nor U12174 (N_12174,N_11865,N_11989);
xor U12175 (N_12175,N_11833,N_11986);
xnor U12176 (N_12176,N_11805,N_11874);
and U12177 (N_12177,N_11966,N_11881);
xnor U12178 (N_12178,N_11941,N_11813);
nor U12179 (N_12179,N_11834,N_11906);
xor U12180 (N_12180,N_11860,N_11808);
nor U12181 (N_12181,N_11954,N_11904);
nor U12182 (N_12182,N_11880,N_11894);
xnor U12183 (N_12183,N_11981,N_11898);
or U12184 (N_12184,N_11939,N_11990);
nor U12185 (N_12185,N_11919,N_11821);
nor U12186 (N_12186,N_11874,N_11925);
nand U12187 (N_12187,N_11938,N_11906);
and U12188 (N_12188,N_11876,N_11868);
and U12189 (N_12189,N_11818,N_11847);
xnor U12190 (N_12190,N_11825,N_11962);
and U12191 (N_12191,N_11848,N_11949);
xor U12192 (N_12192,N_11895,N_11802);
and U12193 (N_12193,N_11970,N_11858);
nand U12194 (N_12194,N_11918,N_11898);
or U12195 (N_12195,N_11826,N_11906);
nand U12196 (N_12196,N_11949,N_11979);
nor U12197 (N_12197,N_11896,N_11875);
and U12198 (N_12198,N_11887,N_11973);
nor U12199 (N_12199,N_11965,N_11805);
and U12200 (N_12200,N_12013,N_12109);
and U12201 (N_12201,N_12103,N_12006);
xor U12202 (N_12202,N_12180,N_12140);
nor U12203 (N_12203,N_12134,N_12070);
xor U12204 (N_12204,N_12104,N_12038);
nor U12205 (N_12205,N_12082,N_12099);
nor U12206 (N_12206,N_12065,N_12007);
nor U12207 (N_12207,N_12021,N_12019);
nand U12208 (N_12208,N_12121,N_12044);
and U12209 (N_12209,N_12122,N_12048);
and U12210 (N_12210,N_12031,N_12067);
and U12211 (N_12211,N_12075,N_12128);
nor U12212 (N_12212,N_12085,N_12097);
nor U12213 (N_12213,N_12023,N_12039);
nand U12214 (N_12214,N_12174,N_12105);
nor U12215 (N_12215,N_12094,N_12059);
nand U12216 (N_12216,N_12111,N_12107);
xnor U12217 (N_12217,N_12143,N_12139);
nor U12218 (N_12218,N_12197,N_12000);
nand U12219 (N_12219,N_12110,N_12062);
or U12220 (N_12220,N_12163,N_12171);
nand U12221 (N_12221,N_12133,N_12046);
or U12222 (N_12222,N_12170,N_12068);
and U12223 (N_12223,N_12159,N_12074);
xor U12224 (N_12224,N_12035,N_12173);
nand U12225 (N_12225,N_12151,N_12029);
xor U12226 (N_12226,N_12020,N_12145);
nand U12227 (N_12227,N_12098,N_12177);
and U12228 (N_12228,N_12175,N_12096);
or U12229 (N_12229,N_12108,N_12005);
or U12230 (N_12230,N_12189,N_12022);
nor U12231 (N_12231,N_12192,N_12193);
and U12232 (N_12232,N_12057,N_12066);
xnor U12233 (N_12233,N_12084,N_12041);
nand U12234 (N_12234,N_12149,N_12072);
and U12235 (N_12235,N_12116,N_12036);
and U12236 (N_12236,N_12091,N_12119);
nand U12237 (N_12237,N_12001,N_12188);
nand U12238 (N_12238,N_12186,N_12079);
or U12239 (N_12239,N_12078,N_12167);
or U12240 (N_12240,N_12049,N_12069);
nand U12241 (N_12241,N_12073,N_12040);
nand U12242 (N_12242,N_12126,N_12131);
xor U12243 (N_12243,N_12172,N_12009);
xnor U12244 (N_12244,N_12125,N_12194);
nand U12245 (N_12245,N_12028,N_12165);
or U12246 (N_12246,N_12004,N_12014);
or U12247 (N_12247,N_12127,N_12156);
xnor U12248 (N_12248,N_12042,N_12010);
xnor U12249 (N_12249,N_12034,N_12088);
or U12250 (N_12250,N_12015,N_12083);
nand U12251 (N_12251,N_12148,N_12132);
xor U12252 (N_12252,N_12179,N_12168);
or U12253 (N_12253,N_12053,N_12118);
and U12254 (N_12254,N_12064,N_12137);
nor U12255 (N_12255,N_12011,N_12050);
nor U12256 (N_12256,N_12155,N_12037);
and U12257 (N_12257,N_12076,N_12164);
nor U12258 (N_12258,N_12135,N_12112);
nor U12259 (N_12259,N_12113,N_12181);
and U12260 (N_12260,N_12101,N_12061);
nor U12261 (N_12261,N_12086,N_12056);
nand U12262 (N_12262,N_12003,N_12185);
xor U12263 (N_12263,N_12152,N_12195);
nor U12264 (N_12264,N_12154,N_12160);
xnor U12265 (N_12265,N_12198,N_12123);
nand U12266 (N_12266,N_12115,N_12055);
and U12267 (N_12267,N_12077,N_12147);
nand U12268 (N_12268,N_12161,N_12138);
nor U12269 (N_12269,N_12045,N_12183);
nor U12270 (N_12270,N_12129,N_12063);
nor U12271 (N_12271,N_12169,N_12178);
xor U12272 (N_12272,N_12018,N_12047);
nand U12273 (N_12273,N_12157,N_12054);
nand U12274 (N_12274,N_12002,N_12024);
nand U12275 (N_12275,N_12136,N_12124);
or U12276 (N_12276,N_12058,N_12196);
and U12277 (N_12277,N_12026,N_12080);
xnor U12278 (N_12278,N_12093,N_12184);
xnor U12279 (N_12279,N_12117,N_12027);
xnor U12280 (N_12280,N_12141,N_12017);
or U12281 (N_12281,N_12142,N_12052);
nand U12282 (N_12282,N_12102,N_12095);
nor U12283 (N_12283,N_12162,N_12051);
nand U12284 (N_12284,N_12130,N_12012);
and U12285 (N_12285,N_12025,N_12106);
nand U12286 (N_12286,N_12182,N_12199);
and U12287 (N_12287,N_12090,N_12191);
or U12288 (N_12288,N_12146,N_12071);
xor U12289 (N_12289,N_12089,N_12016);
nor U12290 (N_12290,N_12030,N_12166);
xnor U12291 (N_12291,N_12120,N_12153);
nor U12292 (N_12292,N_12060,N_12158);
and U12293 (N_12293,N_12087,N_12033);
or U12294 (N_12294,N_12150,N_12081);
xnor U12295 (N_12295,N_12100,N_12144);
or U12296 (N_12296,N_12092,N_12114);
nor U12297 (N_12297,N_12032,N_12008);
and U12298 (N_12298,N_12190,N_12187);
and U12299 (N_12299,N_12043,N_12176);
xor U12300 (N_12300,N_12035,N_12105);
nor U12301 (N_12301,N_12067,N_12058);
or U12302 (N_12302,N_12152,N_12117);
or U12303 (N_12303,N_12104,N_12067);
and U12304 (N_12304,N_12105,N_12145);
and U12305 (N_12305,N_12148,N_12092);
nor U12306 (N_12306,N_12087,N_12088);
and U12307 (N_12307,N_12185,N_12050);
xnor U12308 (N_12308,N_12142,N_12177);
nor U12309 (N_12309,N_12093,N_12104);
xnor U12310 (N_12310,N_12155,N_12184);
or U12311 (N_12311,N_12022,N_12069);
nor U12312 (N_12312,N_12107,N_12181);
nand U12313 (N_12313,N_12183,N_12040);
nor U12314 (N_12314,N_12000,N_12165);
nor U12315 (N_12315,N_12036,N_12181);
nor U12316 (N_12316,N_12024,N_12115);
xor U12317 (N_12317,N_12118,N_12132);
nor U12318 (N_12318,N_12026,N_12162);
nor U12319 (N_12319,N_12124,N_12107);
and U12320 (N_12320,N_12008,N_12124);
or U12321 (N_12321,N_12139,N_12011);
xnor U12322 (N_12322,N_12010,N_12159);
and U12323 (N_12323,N_12006,N_12073);
nor U12324 (N_12324,N_12138,N_12034);
nor U12325 (N_12325,N_12075,N_12181);
and U12326 (N_12326,N_12185,N_12169);
and U12327 (N_12327,N_12145,N_12086);
or U12328 (N_12328,N_12015,N_12081);
nor U12329 (N_12329,N_12132,N_12196);
xor U12330 (N_12330,N_12000,N_12051);
or U12331 (N_12331,N_12094,N_12004);
nor U12332 (N_12332,N_12047,N_12108);
xnor U12333 (N_12333,N_12124,N_12064);
or U12334 (N_12334,N_12026,N_12076);
and U12335 (N_12335,N_12079,N_12089);
or U12336 (N_12336,N_12171,N_12022);
xor U12337 (N_12337,N_12056,N_12007);
nand U12338 (N_12338,N_12151,N_12005);
nand U12339 (N_12339,N_12198,N_12056);
xnor U12340 (N_12340,N_12116,N_12163);
xnor U12341 (N_12341,N_12024,N_12123);
and U12342 (N_12342,N_12020,N_12024);
xor U12343 (N_12343,N_12069,N_12029);
or U12344 (N_12344,N_12034,N_12115);
nor U12345 (N_12345,N_12057,N_12095);
xnor U12346 (N_12346,N_12041,N_12055);
xor U12347 (N_12347,N_12196,N_12117);
xor U12348 (N_12348,N_12074,N_12023);
nor U12349 (N_12349,N_12129,N_12083);
xor U12350 (N_12350,N_12048,N_12176);
xor U12351 (N_12351,N_12190,N_12024);
and U12352 (N_12352,N_12107,N_12095);
nand U12353 (N_12353,N_12151,N_12198);
and U12354 (N_12354,N_12169,N_12122);
or U12355 (N_12355,N_12199,N_12155);
and U12356 (N_12356,N_12055,N_12139);
nand U12357 (N_12357,N_12130,N_12194);
and U12358 (N_12358,N_12075,N_12172);
xnor U12359 (N_12359,N_12033,N_12146);
nor U12360 (N_12360,N_12011,N_12160);
xnor U12361 (N_12361,N_12190,N_12128);
nand U12362 (N_12362,N_12188,N_12126);
xnor U12363 (N_12363,N_12109,N_12055);
nor U12364 (N_12364,N_12194,N_12008);
xor U12365 (N_12365,N_12145,N_12136);
nand U12366 (N_12366,N_12062,N_12014);
nand U12367 (N_12367,N_12101,N_12168);
nor U12368 (N_12368,N_12086,N_12198);
and U12369 (N_12369,N_12095,N_12019);
xnor U12370 (N_12370,N_12043,N_12036);
xor U12371 (N_12371,N_12175,N_12016);
and U12372 (N_12372,N_12197,N_12083);
nand U12373 (N_12373,N_12116,N_12169);
nand U12374 (N_12374,N_12166,N_12095);
and U12375 (N_12375,N_12116,N_12176);
and U12376 (N_12376,N_12116,N_12026);
or U12377 (N_12377,N_12116,N_12197);
nor U12378 (N_12378,N_12012,N_12054);
xor U12379 (N_12379,N_12119,N_12138);
nand U12380 (N_12380,N_12179,N_12076);
xnor U12381 (N_12381,N_12031,N_12149);
or U12382 (N_12382,N_12064,N_12050);
xnor U12383 (N_12383,N_12042,N_12155);
nor U12384 (N_12384,N_12137,N_12030);
nor U12385 (N_12385,N_12177,N_12045);
xnor U12386 (N_12386,N_12077,N_12100);
nor U12387 (N_12387,N_12055,N_12008);
and U12388 (N_12388,N_12036,N_12017);
or U12389 (N_12389,N_12186,N_12041);
xor U12390 (N_12390,N_12159,N_12078);
xor U12391 (N_12391,N_12049,N_12123);
and U12392 (N_12392,N_12006,N_12152);
xnor U12393 (N_12393,N_12147,N_12171);
nand U12394 (N_12394,N_12173,N_12130);
nor U12395 (N_12395,N_12184,N_12182);
nand U12396 (N_12396,N_12158,N_12154);
xnor U12397 (N_12397,N_12035,N_12050);
xor U12398 (N_12398,N_12032,N_12136);
nor U12399 (N_12399,N_12100,N_12003);
xor U12400 (N_12400,N_12215,N_12337);
xor U12401 (N_12401,N_12387,N_12383);
xor U12402 (N_12402,N_12250,N_12245);
xnor U12403 (N_12403,N_12377,N_12283);
xor U12404 (N_12404,N_12395,N_12207);
xnor U12405 (N_12405,N_12299,N_12224);
xor U12406 (N_12406,N_12346,N_12246);
or U12407 (N_12407,N_12364,N_12225);
xnor U12408 (N_12408,N_12307,N_12220);
nand U12409 (N_12409,N_12233,N_12301);
or U12410 (N_12410,N_12267,N_12338);
or U12411 (N_12411,N_12238,N_12232);
nand U12412 (N_12412,N_12200,N_12239);
and U12413 (N_12413,N_12334,N_12317);
nand U12414 (N_12414,N_12252,N_12302);
nand U12415 (N_12415,N_12336,N_12234);
nand U12416 (N_12416,N_12362,N_12290);
nand U12417 (N_12417,N_12343,N_12274);
nor U12418 (N_12418,N_12376,N_12341);
nor U12419 (N_12419,N_12359,N_12351);
xor U12420 (N_12420,N_12356,N_12329);
nand U12421 (N_12421,N_12260,N_12325);
xor U12422 (N_12422,N_12349,N_12357);
nand U12423 (N_12423,N_12235,N_12320);
or U12424 (N_12424,N_12229,N_12298);
nor U12425 (N_12425,N_12399,N_12253);
nand U12426 (N_12426,N_12282,N_12292);
xnor U12427 (N_12427,N_12396,N_12308);
nor U12428 (N_12428,N_12261,N_12248);
or U12429 (N_12429,N_12321,N_12210);
and U12430 (N_12430,N_12392,N_12216);
xnor U12431 (N_12431,N_12398,N_12284);
and U12432 (N_12432,N_12312,N_12353);
nand U12433 (N_12433,N_12240,N_12319);
nand U12434 (N_12434,N_12300,N_12222);
nor U12435 (N_12435,N_12213,N_12231);
nor U12436 (N_12436,N_12350,N_12297);
or U12437 (N_12437,N_12388,N_12258);
nand U12438 (N_12438,N_12397,N_12286);
nand U12439 (N_12439,N_12244,N_12326);
nand U12440 (N_12440,N_12281,N_12278);
and U12441 (N_12441,N_12324,N_12344);
nand U12442 (N_12442,N_12269,N_12360);
nor U12443 (N_12443,N_12389,N_12202);
nand U12444 (N_12444,N_12294,N_12348);
nor U12445 (N_12445,N_12276,N_12355);
nor U12446 (N_12446,N_12205,N_12272);
or U12447 (N_12447,N_12279,N_12322);
nor U12448 (N_12448,N_12306,N_12211);
nand U12449 (N_12449,N_12365,N_12331);
nor U12450 (N_12450,N_12374,N_12369);
nor U12451 (N_12451,N_12333,N_12393);
xor U12452 (N_12452,N_12358,N_12247);
or U12453 (N_12453,N_12316,N_12288);
nor U12454 (N_12454,N_12370,N_12271);
or U12455 (N_12455,N_12277,N_12296);
and U12456 (N_12456,N_12226,N_12372);
and U12457 (N_12457,N_12382,N_12262);
xor U12458 (N_12458,N_12380,N_12264);
xnor U12459 (N_12459,N_12209,N_12265);
and U12460 (N_12460,N_12270,N_12318);
or U12461 (N_12461,N_12304,N_12295);
xor U12462 (N_12462,N_12375,N_12381);
xor U12463 (N_12463,N_12259,N_12352);
or U12464 (N_12464,N_12219,N_12257);
or U12465 (N_12465,N_12354,N_12243);
nor U12466 (N_12466,N_12371,N_12367);
and U12467 (N_12467,N_12221,N_12228);
nand U12468 (N_12468,N_12218,N_12201);
xnor U12469 (N_12469,N_12291,N_12214);
xor U12470 (N_12470,N_12315,N_12368);
and U12471 (N_12471,N_12390,N_12242);
xnor U12472 (N_12472,N_12386,N_12285);
nand U12473 (N_12473,N_12251,N_12223);
xnor U12474 (N_12474,N_12342,N_12335);
nand U12475 (N_12475,N_12293,N_12206);
xnor U12476 (N_12476,N_12266,N_12384);
or U12477 (N_12477,N_12204,N_12328);
or U12478 (N_12478,N_12263,N_12311);
xor U12479 (N_12479,N_12254,N_12237);
or U12480 (N_12480,N_12273,N_12217);
or U12481 (N_12481,N_12391,N_12363);
xor U12482 (N_12482,N_12268,N_12345);
or U12483 (N_12483,N_12255,N_12378);
and U12484 (N_12484,N_12256,N_12289);
nor U12485 (N_12485,N_12385,N_12394);
or U12486 (N_12486,N_12323,N_12203);
xor U12487 (N_12487,N_12275,N_12332);
xnor U12488 (N_12488,N_12339,N_12280);
or U12489 (N_12489,N_12366,N_12309);
xnor U12490 (N_12490,N_12305,N_12373);
or U12491 (N_12491,N_12340,N_12379);
nor U12492 (N_12492,N_12249,N_12327);
nor U12493 (N_12493,N_12230,N_12208);
or U12494 (N_12494,N_12227,N_12361);
nor U12495 (N_12495,N_12287,N_12347);
nor U12496 (N_12496,N_12330,N_12303);
xnor U12497 (N_12497,N_12314,N_12212);
nand U12498 (N_12498,N_12236,N_12313);
and U12499 (N_12499,N_12241,N_12310);
nor U12500 (N_12500,N_12208,N_12234);
nor U12501 (N_12501,N_12380,N_12292);
or U12502 (N_12502,N_12226,N_12357);
nor U12503 (N_12503,N_12375,N_12300);
nor U12504 (N_12504,N_12288,N_12224);
nor U12505 (N_12505,N_12380,N_12243);
xnor U12506 (N_12506,N_12274,N_12214);
or U12507 (N_12507,N_12369,N_12302);
xor U12508 (N_12508,N_12370,N_12244);
or U12509 (N_12509,N_12354,N_12286);
or U12510 (N_12510,N_12284,N_12377);
xor U12511 (N_12511,N_12216,N_12286);
or U12512 (N_12512,N_12248,N_12280);
and U12513 (N_12513,N_12216,N_12346);
xnor U12514 (N_12514,N_12227,N_12332);
or U12515 (N_12515,N_12332,N_12246);
nor U12516 (N_12516,N_12251,N_12336);
nand U12517 (N_12517,N_12249,N_12220);
or U12518 (N_12518,N_12227,N_12306);
and U12519 (N_12519,N_12301,N_12280);
and U12520 (N_12520,N_12394,N_12261);
nor U12521 (N_12521,N_12300,N_12337);
or U12522 (N_12522,N_12285,N_12372);
nor U12523 (N_12523,N_12262,N_12395);
nor U12524 (N_12524,N_12323,N_12245);
nand U12525 (N_12525,N_12256,N_12362);
xor U12526 (N_12526,N_12314,N_12203);
nand U12527 (N_12527,N_12250,N_12376);
and U12528 (N_12528,N_12396,N_12210);
xnor U12529 (N_12529,N_12217,N_12296);
nor U12530 (N_12530,N_12287,N_12211);
xnor U12531 (N_12531,N_12203,N_12313);
and U12532 (N_12532,N_12239,N_12346);
nor U12533 (N_12533,N_12279,N_12272);
xor U12534 (N_12534,N_12316,N_12385);
or U12535 (N_12535,N_12281,N_12220);
or U12536 (N_12536,N_12279,N_12385);
or U12537 (N_12537,N_12391,N_12267);
nand U12538 (N_12538,N_12362,N_12321);
or U12539 (N_12539,N_12393,N_12278);
or U12540 (N_12540,N_12319,N_12304);
and U12541 (N_12541,N_12252,N_12241);
nand U12542 (N_12542,N_12359,N_12271);
or U12543 (N_12543,N_12255,N_12207);
or U12544 (N_12544,N_12359,N_12304);
or U12545 (N_12545,N_12272,N_12347);
nor U12546 (N_12546,N_12385,N_12370);
nand U12547 (N_12547,N_12297,N_12311);
nor U12548 (N_12548,N_12230,N_12327);
xor U12549 (N_12549,N_12324,N_12332);
or U12550 (N_12550,N_12236,N_12322);
nand U12551 (N_12551,N_12398,N_12266);
xor U12552 (N_12552,N_12390,N_12272);
nor U12553 (N_12553,N_12340,N_12281);
or U12554 (N_12554,N_12221,N_12341);
xnor U12555 (N_12555,N_12253,N_12321);
nor U12556 (N_12556,N_12377,N_12384);
xnor U12557 (N_12557,N_12289,N_12359);
and U12558 (N_12558,N_12370,N_12374);
or U12559 (N_12559,N_12386,N_12287);
nand U12560 (N_12560,N_12370,N_12234);
and U12561 (N_12561,N_12205,N_12374);
nand U12562 (N_12562,N_12398,N_12274);
nand U12563 (N_12563,N_12241,N_12213);
nor U12564 (N_12564,N_12281,N_12218);
xnor U12565 (N_12565,N_12340,N_12204);
nand U12566 (N_12566,N_12237,N_12225);
xnor U12567 (N_12567,N_12348,N_12238);
xor U12568 (N_12568,N_12388,N_12329);
nand U12569 (N_12569,N_12343,N_12396);
or U12570 (N_12570,N_12236,N_12278);
and U12571 (N_12571,N_12370,N_12227);
or U12572 (N_12572,N_12233,N_12217);
or U12573 (N_12573,N_12285,N_12384);
and U12574 (N_12574,N_12319,N_12233);
xor U12575 (N_12575,N_12374,N_12227);
nor U12576 (N_12576,N_12337,N_12270);
nand U12577 (N_12577,N_12202,N_12368);
xor U12578 (N_12578,N_12245,N_12385);
and U12579 (N_12579,N_12255,N_12231);
nor U12580 (N_12580,N_12243,N_12269);
xnor U12581 (N_12581,N_12347,N_12392);
nor U12582 (N_12582,N_12311,N_12266);
xor U12583 (N_12583,N_12224,N_12398);
and U12584 (N_12584,N_12204,N_12338);
nand U12585 (N_12585,N_12267,N_12251);
nor U12586 (N_12586,N_12259,N_12273);
and U12587 (N_12587,N_12204,N_12226);
and U12588 (N_12588,N_12328,N_12322);
and U12589 (N_12589,N_12238,N_12265);
or U12590 (N_12590,N_12386,N_12309);
xnor U12591 (N_12591,N_12304,N_12325);
nor U12592 (N_12592,N_12211,N_12282);
nand U12593 (N_12593,N_12292,N_12319);
nand U12594 (N_12594,N_12212,N_12313);
nand U12595 (N_12595,N_12207,N_12388);
nand U12596 (N_12596,N_12360,N_12276);
nand U12597 (N_12597,N_12334,N_12273);
xnor U12598 (N_12598,N_12294,N_12221);
nor U12599 (N_12599,N_12256,N_12395);
or U12600 (N_12600,N_12587,N_12413);
or U12601 (N_12601,N_12513,N_12585);
or U12602 (N_12602,N_12477,N_12417);
xnor U12603 (N_12603,N_12459,N_12435);
or U12604 (N_12604,N_12568,N_12570);
nor U12605 (N_12605,N_12541,N_12569);
or U12606 (N_12606,N_12474,N_12412);
and U12607 (N_12607,N_12420,N_12497);
or U12608 (N_12608,N_12532,N_12437);
and U12609 (N_12609,N_12489,N_12466);
and U12610 (N_12610,N_12400,N_12451);
nand U12611 (N_12611,N_12411,N_12582);
or U12612 (N_12612,N_12523,N_12554);
and U12613 (N_12613,N_12555,N_12482);
nand U12614 (N_12614,N_12567,N_12594);
xor U12615 (N_12615,N_12467,N_12551);
and U12616 (N_12616,N_12572,N_12552);
nand U12617 (N_12617,N_12476,N_12506);
nand U12618 (N_12618,N_12422,N_12447);
or U12619 (N_12619,N_12470,N_12531);
nand U12620 (N_12620,N_12425,N_12414);
or U12621 (N_12621,N_12516,N_12596);
nor U12622 (N_12622,N_12574,N_12591);
and U12623 (N_12623,N_12561,N_12548);
and U12624 (N_12624,N_12547,N_12500);
nand U12625 (N_12625,N_12529,N_12403);
nor U12626 (N_12626,N_12521,N_12431);
nor U12627 (N_12627,N_12540,N_12433);
nor U12628 (N_12628,N_12571,N_12441);
or U12629 (N_12629,N_12498,N_12449);
xor U12630 (N_12630,N_12592,N_12559);
or U12631 (N_12631,N_12597,N_12423);
and U12632 (N_12632,N_12493,N_12410);
nand U12633 (N_12633,N_12581,N_12462);
or U12634 (N_12634,N_12446,N_12550);
and U12635 (N_12635,N_12522,N_12486);
xor U12636 (N_12636,N_12557,N_12586);
and U12637 (N_12637,N_12499,N_12469);
xor U12638 (N_12638,N_12440,N_12565);
xor U12639 (N_12639,N_12471,N_12503);
xnor U12640 (N_12640,N_12598,N_12426);
or U12641 (N_12641,N_12443,N_12536);
or U12642 (N_12642,N_12519,N_12401);
xor U12643 (N_12643,N_12409,N_12496);
and U12644 (N_12644,N_12589,N_12428);
or U12645 (N_12645,N_12590,N_12452);
nor U12646 (N_12646,N_12419,N_12583);
and U12647 (N_12647,N_12448,N_12580);
and U12648 (N_12648,N_12406,N_12456);
and U12649 (N_12649,N_12450,N_12595);
nor U12650 (N_12650,N_12525,N_12593);
and U12651 (N_12651,N_12566,N_12512);
or U12652 (N_12652,N_12494,N_12530);
and U12653 (N_12653,N_12442,N_12575);
and U12654 (N_12654,N_12479,N_12430);
or U12655 (N_12655,N_12543,N_12468);
or U12656 (N_12656,N_12535,N_12495);
xnor U12657 (N_12657,N_12416,N_12524);
or U12658 (N_12658,N_12488,N_12408);
or U12659 (N_12659,N_12511,N_12485);
and U12660 (N_12660,N_12458,N_12472);
xnor U12661 (N_12661,N_12577,N_12599);
nor U12662 (N_12662,N_12424,N_12421);
xnor U12663 (N_12663,N_12504,N_12556);
nand U12664 (N_12664,N_12515,N_12432);
and U12665 (N_12665,N_12546,N_12473);
or U12666 (N_12666,N_12478,N_12507);
nor U12667 (N_12667,N_12520,N_12514);
or U12668 (N_12668,N_12492,N_12537);
nand U12669 (N_12669,N_12518,N_12402);
nor U12670 (N_12670,N_12510,N_12434);
or U12671 (N_12671,N_12553,N_12579);
nor U12672 (N_12672,N_12445,N_12501);
xnor U12673 (N_12673,N_12562,N_12427);
or U12674 (N_12674,N_12483,N_12502);
nor U12675 (N_12675,N_12560,N_12544);
xor U12676 (N_12676,N_12509,N_12484);
and U12677 (N_12677,N_12549,N_12444);
nand U12678 (N_12678,N_12439,N_12429);
and U12679 (N_12679,N_12407,N_12404);
and U12680 (N_12680,N_12563,N_12545);
and U12681 (N_12681,N_12481,N_12508);
nor U12682 (N_12682,N_12505,N_12455);
or U12683 (N_12683,N_12564,N_12576);
or U12684 (N_12684,N_12464,N_12465);
nor U12685 (N_12685,N_12588,N_12584);
xor U12686 (N_12686,N_12453,N_12491);
nand U12687 (N_12687,N_12461,N_12534);
xnor U12688 (N_12688,N_12463,N_12415);
or U12689 (N_12689,N_12436,N_12460);
nand U12690 (N_12690,N_12490,N_12418);
nand U12691 (N_12691,N_12542,N_12454);
and U12692 (N_12692,N_12475,N_12558);
nand U12693 (N_12693,N_12480,N_12438);
and U12694 (N_12694,N_12528,N_12457);
and U12695 (N_12695,N_12533,N_12527);
nand U12696 (N_12696,N_12526,N_12578);
nand U12697 (N_12697,N_12517,N_12539);
and U12698 (N_12698,N_12487,N_12538);
or U12699 (N_12699,N_12573,N_12405);
and U12700 (N_12700,N_12400,N_12416);
nand U12701 (N_12701,N_12502,N_12498);
xnor U12702 (N_12702,N_12471,N_12594);
or U12703 (N_12703,N_12478,N_12541);
or U12704 (N_12704,N_12508,N_12479);
nand U12705 (N_12705,N_12441,N_12590);
nor U12706 (N_12706,N_12504,N_12524);
or U12707 (N_12707,N_12400,N_12410);
and U12708 (N_12708,N_12429,N_12555);
and U12709 (N_12709,N_12560,N_12435);
xnor U12710 (N_12710,N_12476,N_12475);
or U12711 (N_12711,N_12448,N_12561);
xnor U12712 (N_12712,N_12562,N_12576);
nand U12713 (N_12713,N_12465,N_12569);
xnor U12714 (N_12714,N_12496,N_12524);
or U12715 (N_12715,N_12597,N_12534);
xnor U12716 (N_12716,N_12554,N_12565);
xor U12717 (N_12717,N_12542,N_12430);
and U12718 (N_12718,N_12515,N_12557);
xnor U12719 (N_12719,N_12526,N_12450);
xor U12720 (N_12720,N_12507,N_12456);
xnor U12721 (N_12721,N_12440,N_12412);
and U12722 (N_12722,N_12590,N_12599);
nor U12723 (N_12723,N_12552,N_12585);
nor U12724 (N_12724,N_12455,N_12568);
or U12725 (N_12725,N_12491,N_12492);
or U12726 (N_12726,N_12425,N_12589);
or U12727 (N_12727,N_12503,N_12427);
xor U12728 (N_12728,N_12416,N_12423);
or U12729 (N_12729,N_12596,N_12591);
nand U12730 (N_12730,N_12428,N_12515);
nand U12731 (N_12731,N_12427,N_12525);
xnor U12732 (N_12732,N_12481,N_12491);
xor U12733 (N_12733,N_12498,N_12440);
xnor U12734 (N_12734,N_12584,N_12568);
xnor U12735 (N_12735,N_12573,N_12423);
nor U12736 (N_12736,N_12442,N_12566);
nand U12737 (N_12737,N_12530,N_12462);
nand U12738 (N_12738,N_12525,N_12476);
nand U12739 (N_12739,N_12458,N_12492);
and U12740 (N_12740,N_12517,N_12544);
nor U12741 (N_12741,N_12460,N_12416);
nand U12742 (N_12742,N_12577,N_12591);
or U12743 (N_12743,N_12522,N_12500);
or U12744 (N_12744,N_12534,N_12521);
and U12745 (N_12745,N_12441,N_12531);
xnor U12746 (N_12746,N_12480,N_12492);
or U12747 (N_12747,N_12581,N_12432);
nor U12748 (N_12748,N_12479,N_12560);
or U12749 (N_12749,N_12560,N_12561);
nand U12750 (N_12750,N_12542,N_12502);
and U12751 (N_12751,N_12435,N_12544);
nor U12752 (N_12752,N_12423,N_12558);
nor U12753 (N_12753,N_12534,N_12546);
nand U12754 (N_12754,N_12552,N_12406);
or U12755 (N_12755,N_12452,N_12558);
xnor U12756 (N_12756,N_12510,N_12517);
or U12757 (N_12757,N_12507,N_12521);
xor U12758 (N_12758,N_12532,N_12463);
and U12759 (N_12759,N_12417,N_12561);
and U12760 (N_12760,N_12554,N_12532);
nand U12761 (N_12761,N_12564,N_12580);
nor U12762 (N_12762,N_12436,N_12474);
nor U12763 (N_12763,N_12591,N_12535);
or U12764 (N_12764,N_12584,N_12493);
xor U12765 (N_12765,N_12567,N_12528);
nor U12766 (N_12766,N_12525,N_12405);
nor U12767 (N_12767,N_12526,N_12428);
nor U12768 (N_12768,N_12523,N_12466);
xnor U12769 (N_12769,N_12446,N_12570);
nor U12770 (N_12770,N_12532,N_12501);
nor U12771 (N_12771,N_12441,N_12403);
xor U12772 (N_12772,N_12549,N_12468);
nand U12773 (N_12773,N_12522,N_12489);
nand U12774 (N_12774,N_12427,N_12527);
and U12775 (N_12775,N_12583,N_12441);
nand U12776 (N_12776,N_12527,N_12542);
or U12777 (N_12777,N_12552,N_12570);
xor U12778 (N_12778,N_12509,N_12461);
or U12779 (N_12779,N_12536,N_12403);
and U12780 (N_12780,N_12435,N_12542);
and U12781 (N_12781,N_12493,N_12490);
nand U12782 (N_12782,N_12491,N_12532);
xor U12783 (N_12783,N_12435,N_12559);
or U12784 (N_12784,N_12504,N_12454);
or U12785 (N_12785,N_12433,N_12460);
xor U12786 (N_12786,N_12536,N_12572);
xor U12787 (N_12787,N_12536,N_12535);
xnor U12788 (N_12788,N_12494,N_12446);
and U12789 (N_12789,N_12592,N_12581);
nand U12790 (N_12790,N_12499,N_12569);
nand U12791 (N_12791,N_12585,N_12560);
and U12792 (N_12792,N_12525,N_12485);
xnor U12793 (N_12793,N_12430,N_12552);
and U12794 (N_12794,N_12416,N_12554);
xnor U12795 (N_12795,N_12486,N_12523);
nand U12796 (N_12796,N_12564,N_12536);
or U12797 (N_12797,N_12494,N_12513);
nand U12798 (N_12798,N_12561,N_12527);
and U12799 (N_12799,N_12589,N_12477);
or U12800 (N_12800,N_12748,N_12610);
nor U12801 (N_12801,N_12692,N_12649);
and U12802 (N_12802,N_12660,N_12686);
nor U12803 (N_12803,N_12755,N_12792);
or U12804 (N_12804,N_12664,N_12679);
nor U12805 (N_12805,N_12689,N_12645);
and U12806 (N_12806,N_12776,N_12684);
or U12807 (N_12807,N_12608,N_12713);
and U12808 (N_12808,N_12743,N_12670);
or U12809 (N_12809,N_12709,N_12668);
or U12810 (N_12810,N_12667,N_12678);
or U12811 (N_12811,N_12632,N_12751);
and U12812 (N_12812,N_12688,N_12785);
nand U12813 (N_12813,N_12798,N_12745);
nor U12814 (N_12814,N_12711,N_12677);
nand U12815 (N_12815,N_12734,N_12676);
or U12816 (N_12816,N_12714,N_12696);
and U12817 (N_12817,N_12768,N_12741);
nor U12818 (N_12818,N_12720,N_12631);
xor U12819 (N_12819,N_12702,N_12630);
or U12820 (N_12820,N_12726,N_12722);
nor U12821 (N_12821,N_12760,N_12795);
or U12822 (N_12822,N_12721,N_12646);
nand U12823 (N_12823,N_12700,N_12765);
nand U12824 (N_12824,N_12715,N_12797);
or U12825 (N_12825,N_12789,N_12611);
nand U12826 (N_12826,N_12782,N_12779);
xor U12827 (N_12827,N_12773,N_12603);
xor U12828 (N_12828,N_12612,N_12628);
or U12829 (N_12829,N_12730,N_12719);
or U12830 (N_12830,N_12793,N_12662);
or U12831 (N_12831,N_12787,N_12706);
xor U12832 (N_12832,N_12757,N_12669);
nand U12833 (N_12833,N_12724,N_12791);
nand U12834 (N_12834,N_12614,N_12665);
xor U12835 (N_12835,N_12694,N_12708);
or U12836 (N_12836,N_12749,N_12763);
xnor U12837 (N_12837,N_12635,N_12737);
and U12838 (N_12838,N_12777,N_12753);
or U12839 (N_12839,N_12717,N_12756);
nor U12840 (N_12840,N_12698,N_12659);
or U12841 (N_12841,N_12607,N_12761);
xor U12842 (N_12842,N_12727,N_12764);
and U12843 (N_12843,N_12732,N_12769);
nand U12844 (N_12844,N_12666,N_12639);
xor U12845 (N_12845,N_12775,N_12671);
nor U12846 (N_12846,N_12653,N_12729);
nand U12847 (N_12847,N_12752,N_12625);
nor U12848 (N_12848,N_12691,N_12739);
and U12849 (N_12849,N_12788,N_12786);
xor U12850 (N_12850,N_12673,N_12758);
or U12851 (N_12851,N_12606,N_12703);
nand U12852 (N_12852,N_12747,N_12643);
nor U12853 (N_12853,N_12601,N_12716);
and U12854 (N_12854,N_12731,N_12627);
and U12855 (N_12855,N_12622,N_12641);
nor U12856 (N_12856,N_12796,N_12783);
nand U12857 (N_12857,N_12693,N_12674);
or U12858 (N_12858,N_12634,N_12799);
and U12859 (N_12859,N_12762,N_12682);
nand U12860 (N_12860,N_12638,N_12617);
nand U12861 (N_12861,N_12784,N_12772);
or U12862 (N_12862,N_12636,N_12774);
and U12863 (N_12863,N_12633,N_12754);
or U12864 (N_12864,N_12781,N_12746);
and U12865 (N_12865,N_12623,N_12655);
nor U12866 (N_12866,N_12640,N_12613);
nor U12867 (N_12867,N_12705,N_12626);
xnor U12868 (N_12868,N_12750,N_12735);
xor U12869 (N_12869,N_12742,N_12728);
nand U12870 (N_12870,N_12766,N_12707);
xnor U12871 (N_12871,N_12605,N_12657);
nand U12872 (N_12872,N_12624,N_12699);
and U12873 (N_12873,N_12661,N_12740);
or U12874 (N_12874,N_12654,N_12770);
nor U12875 (N_12875,N_12680,N_12615);
or U12876 (N_12876,N_12650,N_12681);
nand U12877 (N_12877,N_12629,N_12663);
xnor U12878 (N_12878,N_12723,N_12790);
xor U12879 (N_12879,N_12652,N_12794);
or U12880 (N_12880,N_12736,N_12780);
xnor U12881 (N_12881,N_12609,N_12710);
nor U12882 (N_12882,N_12778,N_12771);
nor U12883 (N_12883,N_12733,N_12697);
and U12884 (N_12884,N_12738,N_12618);
xor U12885 (N_12885,N_12658,N_12725);
xnor U12886 (N_12886,N_12600,N_12685);
nand U12887 (N_12887,N_12687,N_12647);
or U12888 (N_12888,N_12704,N_12620);
or U12889 (N_12889,N_12619,N_12651);
and U12890 (N_12890,N_12616,N_12744);
and U12891 (N_12891,N_12672,N_12712);
xnor U12892 (N_12892,N_12690,N_12718);
xnor U12893 (N_12893,N_12637,N_12695);
and U12894 (N_12894,N_12701,N_12675);
nand U12895 (N_12895,N_12683,N_12648);
nand U12896 (N_12896,N_12602,N_12644);
nand U12897 (N_12897,N_12621,N_12656);
nand U12898 (N_12898,N_12767,N_12642);
or U12899 (N_12899,N_12759,N_12604);
xor U12900 (N_12900,N_12623,N_12752);
or U12901 (N_12901,N_12715,N_12716);
nor U12902 (N_12902,N_12602,N_12696);
nand U12903 (N_12903,N_12752,N_12697);
and U12904 (N_12904,N_12614,N_12729);
nand U12905 (N_12905,N_12789,N_12633);
nand U12906 (N_12906,N_12600,N_12703);
nor U12907 (N_12907,N_12788,N_12674);
xnor U12908 (N_12908,N_12712,N_12704);
nor U12909 (N_12909,N_12674,N_12727);
xnor U12910 (N_12910,N_12723,N_12611);
nand U12911 (N_12911,N_12685,N_12743);
xnor U12912 (N_12912,N_12668,N_12764);
and U12913 (N_12913,N_12652,N_12617);
and U12914 (N_12914,N_12717,N_12722);
and U12915 (N_12915,N_12662,N_12726);
nand U12916 (N_12916,N_12654,N_12629);
nand U12917 (N_12917,N_12641,N_12782);
nor U12918 (N_12918,N_12763,N_12670);
xnor U12919 (N_12919,N_12682,N_12713);
or U12920 (N_12920,N_12718,N_12739);
and U12921 (N_12921,N_12670,N_12681);
and U12922 (N_12922,N_12715,N_12792);
or U12923 (N_12923,N_12632,N_12778);
xor U12924 (N_12924,N_12745,N_12792);
nand U12925 (N_12925,N_12619,N_12766);
and U12926 (N_12926,N_12785,N_12609);
xor U12927 (N_12927,N_12780,N_12690);
nor U12928 (N_12928,N_12780,N_12685);
xor U12929 (N_12929,N_12693,N_12682);
nor U12930 (N_12930,N_12676,N_12723);
xnor U12931 (N_12931,N_12690,N_12737);
nor U12932 (N_12932,N_12627,N_12750);
nand U12933 (N_12933,N_12640,N_12793);
or U12934 (N_12934,N_12779,N_12768);
nor U12935 (N_12935,N_12741,N_12758);
nor U12936 (N_12936,N_12753,N_12756);
or U12937 (N_12937,N_12763,N_12618);
nor U12938 (N_12938,N_12713,N_12629);
or U12939 (N_12939,N_12769,N_12697);
nand U12940 (N_12940,N_12759,N_12735);
nand U12941 (N_12941,N_12784,N_12622);
nand U12942 (N_12942,N_12662,N_12686);
nor U12943 (N_12943,N_12675,N_12791);
or U12944 (N_12944,N_12748,N_12753);
nor U12945 (N_12945,N_12716,N_12704);
xor U12946 (N_12946,N_12601,N_12645);
or U12947 (N_12947,N_12751,N_12744);
nand U12948 (N_12948,N_12754,N_12720);
and U12949 (N_12949,N_12640,N_12641);
xnor U12950 (N_12950,N_12770,N_12636);
nor U12951 (N_12951,N_12613,N_12637);
nor U12952 (N_12952,N_12610,N_12617);
nand U12953 (N_12953,N_12667,N_12723);
or U12954 (N_12954,N_12641,N_12734);
nand U12955 (N_12955,N_12626,N_12716);
and U12956 (N_12956,N_12773,N_12745);
xor U12957 (N_12957,N_12627,N_12773);
or U12958 (N_12958,N_12654,N_12792);
nor U12959 (N_12959,N_12611,N_12691);
nor U12960 (N_12960,N_12648,N_12744);
nand U12961 (N_12961,N_12633,N_12768);
nand U12962 (N_12962,N_12764,N_12601);
and U12963 (N_12963,N_12611,N_12757);
xor U12964 (N_12964,N_12696,N_12604);
xor U12965 (N_12965,N_12678,N_12768);
nand U12966 (N_12966,N_12707,N_12638);
nor U12967 (N_12967,N_12697,N_12730);
nor U12968 (N_12968,N_12780,N_12768);
nand U12969 (N_12969,N_12754,N_12608);
nor U12970 (N_12970,N_12766,N_12765);
nor U12971 (N_12971,N_12725,N_12644);
xnor U12972 (N_12972,N_12697,N_12737);
xor U12973 (N_12973,N_12682,N_12615);
and U12974 (N_12974,N_12643,N_12665);
and U12975 (N_12975,N_12659,N_12749);
or U12976 (N_12976,N_12777,N_12637);
or U12977 (N_12977,N_12708,N_12652);
xnor U12978 (N_12978,N_12605,N_12621);
or U12979 (N_12979,N_12757,N_12733);
nor U12980 (N_12980,N_12621,N_12792);
xor U12981 (N_12981,N_12696,N_12742);
and U12982 (N_12982,N_12759,N_12731);
xnor U12983 (N_12983,N_12690,N_12714);
xnor U12984 (N_12984,N_12645,N_12646);
xnor U12985 (N_12985,N_12681,N_12608);
nand U12986 (N_12986,N_12651,N_12689);
xor U12987 (N_12987,N_12624,N_12720);
nor U12988 (N_12988,N_12604,N_12765);
and U12989 (N_12989,N_12753,N_12681);
or U12990 (N_12990,N_12782,N_12657);
nor U12991 (N_12991,N_12615,N_12608);
xnor U12992 (N_12992,N_12797,N_12703);
xor U12993 (N_12993,N_12758,N_12679);
and U12994 (N_12994,N_12775,N_12752);
and U12995 (N_12995,N_12622,N_12618);
and U12996 (N_12996,N_12728,N_12681);
nand U12997 (N_12997,N_12685,N_12675);
xnor U12998 (N_12998,N_12741,N_12619);
xor U12999 (N_12999,N_12696,N_12671);
and U13000 (N_13000,N_12854,N_12835);
nor U13001 (N_13001,N_12981,N_12831);
nand U13002 (N_13002,N_12915,N_12907);
nand U13003 (N_13003,N_12879,N_12962);
or U13004 (N_13004,N_12852,N_12996);
nor U13005 (N_13005,N_12971,N_12936);
nand U13006 (N_13006,N_12951,N_12955);
nand U13007 (N_13007,N_12860,N_12837);
or U13008 (N_13008,N_12894,N_12923);
or U13009 (N_13009,N_12901,N_12979);
nor U13010 (N_13010,N_12966,N_12851);
and U13011 (N_13011,N_12875,N_12819);
nand U13012 (N_13012,N_12980,N_12909);
or U13013 (N_13013,N_12813,N_12916);
and U13014 (N_13014,N_12914,N_12934);
nand U13015 (N_13015,N_12977,N_12919);
and U13016 (N_13016,N_12965,N_12821);
nor U13017 (N_13017,N_12843,N_12888);
nand U13018 (N_13018,N_12807,N_12994);
nand U13019 (N_13019,N_12815,N_12887);
or U13020 (N_13020,N_12844,N_12984);
and U13021 (N_13021,N_12929,N_12990);
and U13022 (N_13022,N_12858,N_12836);
nor U13023 (N_13023,N_12918,N_12871);
xor U13024 (N_13024,N_12989,N_12937);
nor U13025 (N_13025,N_12949,N_12926);
or U13026 (N_13026,N_12925,N_12892);
and U13027 (N_13027,N_12866,N_12886);
nor U13028 (N_13028,N_12822,N_12855);
xor U13029 (N_13029,N_12904,N_12896);
nor U13030 (N_13030,N_12933,N_12961);
xor U13031 (N_13031,N_12959,N_12868);
nand U13032 (N_13032,N_12898,N_12922);
nor U13033 (N_13033,N_12804,N_12972);
or U13034 (N_13034,N_12801,N_12912);
and U13035 (N_13035,N_12952,N_12803);
nand U13036 (N_13036,N_12833,N_12802);
nand U13037 (N_13037,N_12884,N_12825);
and U13038 (N_13038,N_12828,N_12842);
nor U13039 (N_13039,N_12985,N_12857);
nor U13040 (N_13040,N_12834,N_12908);
nand U13041 (N_13041,N_12905,N_12808);
nor U13042 (N_13042,N_12920,N_12900);
nand U13043 (N_13043,N_12805,N_12950);
xnor U13044 (N_13044,N_12917,N_12849);
or U13045 (N_13045,N_12800,N_12942);
nand U13046 (N_13046,N_12853,N_12811);
nand U13047 (N_13047,N_12978,N_12997);
xnor U13048 (N_13048,N_12903,N_12940);
and U13049 (N_13049,N_12998,N_12867);
xnor U13050 (N_13050,N_12812,N_12938);
nor U13051 (N_13051,N_12945,N_12986);
nand U13052 (N_13052,N_12932,N_12841);
or U13053 (N_13053,N_12885,N_12993);
xor U13054 (N_13054,N_12838,N_12935);
nand U13055 (N_13055,N_12873,N_12830);
or U13056 (N_13056,N_12969,N_12928);
nand U13057 (N_13057,N_12816,N_12818);
nor U13058 (N_13058,N_12839,N_12988);
or U13059 (N_13059,N_12899,N_12958);
or U13060 (N_13060,N_12939,N_12893);
xor U13061 (N_13061,N_12859,N_12829);
xor U13062 (N_13062,N_12881,N_12876);
nand U13063 (N_13063,N_12960,N_12814);
or U13064 (N_13064,N_12810,N_12957);
nand U13065 (N_13065,N_12954,N_12991);
nand U13066 (N_13066,N_12806,N_12877);
and U13067 (N_13067,N_12878,N_12906);
nand U13068 (N_13068,N_12883,N_12850);
nand U13069 (N_13069,N_12872,N_12891);
nor U13070 (N_13070,N_12832,N_12968);
nand U13071 (N_13071,N_12927,N_12889);
or U13072 (N_13072,N_12913,N_12987);
nor U13073 (N_13073,N_12953,N_12882);
or U13074 (N_13074,N_12847,N_12973);
nand U13075 (N_13075,N_12823,N_12826);
nand U13076 (N_13076,N_12943,N_12809);
and U13077 (N_13077,N_12967,N_12924);
nand U13078 (N_13078,N_12820,N_12911);
nor U13079 (N_13079,N_12846,N_12880);
xor U13080 (N_13080,N_12964,N_12948);
nand U13081 (N_13081,N_12863,N_12975);
nor U13082 (N_13082,N_12976,N_12970);
or U13083 (N_13083,N_12890,N_12992);
nand U13084 (N_13084,N_12946,N_12983);
and U13085 (N_13085,N_12874,N_12941);
and U13086 (N_13086,N_12944,N_12921);
nor U13087 (N_13087,N_12848,N_12817);
or U13088 (N_13088,N_12827,N_12963);
nand U13089 (N_13089,N_12895,N_12840);
nand U13090 (N_13090,N_12930,N_12869);
or U13091 (N_13091,N_12856,N_12870);
or U13092 (N_13092,N_12902,N_12931);
and U13093 (N_13093,N_12999,N_12824);
or U13094 (N_13094,N_12974,N_12995);
nand U13095 (N_13095,N_12910,N_12865);
and U13096 (N_13096,N_12864,N_12982);
nand U13097 (N_13097,N_12947,N_12861);
or U13098 (N_13098,N_12845,N_12956);
xnor U13099 (N_13099,N_12897,N_12862);
nor U13100 (N_13100,N_12990,N_12931);
nand U13101 (N_13101,N_12869,N_12815);
or U13102 (N_13102,N_12890,N_12900);
xnor U13103 (N_13103,N_12856,N_12995);
nand U13104 (N_13104,N_12871,N_12860);
and U13105 (N_13105,N_12891,N_12880);
xnor U13106 (N_13106,N_12892,N_12943);
and U13107 (N_13107,N_12807,N_12970);
xor U13108 (N_13108,N_12990,N_12840);
and U13109 (N_13109,N_12924,N_12841);
nor U13110 (N_13110,N_12874,N_12982);
or U13111 (N_13111,N_12814,N_12895);
nor U13112 (N_13112,N_12805,N_12840);
and U13113 (N_13113,N_12897,N_12985);
nand U13114 (N_13114,N_12822,N_12853);
and U13115 (N_13115,N_12944,N_12915);
or U13116 (N_13116,N_12832,N_12874);
xor U13117 (N_13117,N_12871,N_12898);
xnor U13118 (N_13118,N_12960,N_12987);
nor U13119 (N_13119,N_12913,N_12812);
or U13120 (N_13120,N_12823,N_12896);
or U13121 (N_13121,N_12988,N_12815);
xor U13122 (N_13122,N_12928,N_12945);
xnor U13123 (N_13123,N_12856,N_12822);
xnor U13124 (N_13124,N_12979,N_12976);
xor U13125 (N_13125,N_12832,N_12881);
and U13126 (N_13126,N_12925,N_12801);
nand U13127 (N_13127,N_12809,N_12845);
nand U13128 (N_13128,N_12925,N_12907);
xor U13129 (N_13129,N_12872,N_12967);
xnor U13130 (N_13130,N_12972,N_12949);
nor U13131 (N_13131,N_12875,N_12947);
nor U13132 (N_13132,N_12996,N_12907);
nand U13133 (N_13133,N_12904,N_12829);
and U13134 (N_13134,N_12900,N_12932);
nor U13135 (N_13135,N_12923,N_12880);
and U13136 (N_13136,N_12915,N_12912);
and U13137 (N_13137,N_12873,N_12855);
xnor U13138 (N_13138,N_12877,N_12900);
nand U13139 (N_13139,N_12806,N_12939);
nor U13140 (N_13140,N_12818,N_12825);
xnor U13141 (N_13141,N_12989,N_12837);
or U13142 (N_13142,N_12894,N_12931);
nand U13143 (N_13143,N_12989,N_12857);
and U13144 (N_13144,N_12897,N_12866);
and U13145 (N_13145,N_12929,N_12962);
or U13146 (N_13146,N_12943,N_12958);
xnor U13147 (N_13147,N_12807,N_12899);
nand U13148 (N_13148,N_12965,N_12982);
xor U13149 (N_13149,N_12956,N_12999);
nor U13150 (N_13150,N_12989,N_12870);
xnor U13151 (N_13151,N_12828,N_12989);
and U13152 (N_13152,N_12848,N_12829);
and U13153 (N_13153,N_12884,N_12957);
nor U13154 (N_13154,N_12992,N_12885);
nand U13155 (N_13155,N_12895,N_12986);
or U13156 (N_13156,N_12984,N_12941);
and U13157 (N_13157,N_12837,N_12905);
nand U13158 (N_13158,N_12845,N_12858);
or U13159 (N_13159,N_12923,N_12874);
and U13160 (N_13160,N_12862,N_12932);
nand U13161 (N_13161,N_12842,N_12973);
and U13162 (N_13162,N_12962,N_12865);
nand U13163 (N_13163,N_12849,N_12983);
nand U13164 (N_13164,N_12932,N_12918);
and U13165 (N_13165,N_12898,N_12901);
or U13166 (N_13166,N_12964,N_12930);
nand U13167 (N_13167,N_12979,N_12803);
nand U13168 (N_13168,N_12842,N_12998);
nor U13169 (N_13169,N_12855,N_12913);
nand U13170 (N_13170,N_12837,N_12906);
and U13171 (N_13171,N_12877,N_12807);
and U13172 (N_13172,N_12970,N_12834);
and U13173 (N_13173,N_12846,N_12848);
or U13174 (N_13174,N_12811,N_12992);
nor U13175 (N_13175,N_12824,N_12893);
nand U13176 (N_13176,N_12919,N_12984);
nand U13177 (N_13177,N_12968,N_12881);
xnor U13178 (N_13178,N_12990,N_12969);
or U13179 (N_13179,N_12886,N_12821);
nor U13180 (N_13180,N_12907,N_12979);
or U13181 (N_13181,N_12923,N_12994);
and U13182 (N_13182,N_12843,N_12990);
nand U13183 (N_13183,N_12841,N_12882);
nand U13184 (N_13184,N_12978,N_12921);
nor U13185 (N_13185,N_12885,N_12898);
xnor U13186 (N_13186,N_12912,N_12844);
and U13187 (N_13187,N_12999,N_12898);
and U13188 (N_13188,N_12947,N_12916);
nor U13189 (N_13189,N_12966,N_12913);
nand U13190 (N_13190,N_12886,N_12965);
nor U13191 (N_13191,N_12923,N_12876);
nor U13192 (N_13192,N_12898,N_12867);
xnor U13193 (N_13193,N_12943,N_12856);
or U13194 (N_13194,N_12996,N_12860);
xor U13195 (N_13195,N_12844,N_12914);
xnor U13196 (N_13196,N_12840,N_12802);
xor U13197 (N_13197,N_12900,N_12849);
and U13198 (N_13198,N_12954,N_12818);
and U13199 (N_13199,N_12942,N_12812);
nand U13200 (N_13200,N_13162,N_13115);
nor U13201 (N_13201,N_13000,N_13002);
or U13202 (N_13202,N_13193,N_13073);
or U13203 (N_13203,N_13160,N_13096);
nor U13204 (N_13204,N_13030,N_13171);
nor U13205 (N_13205,N_13014,N_13145);
or U13206 (N_13206,N_13147,N_13190);
and U13207 (N_13207,N_13048,N_13107);
or U13208 (N_13208,N_13062,N_13126);
nor U13209 (N_13209,N_13024,N_13165);
or U13210 (N_13210,N_13138,N_13117);
or U13211 (N_13211,N_13097,N_13125);
nand U13212 (N_13212,N_13188,N_13098);
nand U13213 (N_13213,N_13018,N_13122);
nor U13214 (N_13214,N_13156,N_13169);
and U13215 (N_13215,N_13144,N_13141);
and U13216 (N_13216,N_13075,N_13167);
nor U13217 (N_13217,N_13194,N_13198);
and U13218 (N_13218,N_13049,N_13146);
nor U13219 (N_13219,N_13152,N_13143);
and U13220 (N_13220,N_13140,N_13151);
xor U13221 (N_13221,N_13076,N_13134);
xor U13222 (N_13222,N_13094,N_13178);
xor U13223 (N_13223,N_13054,N_13072);
nand U13224 (N_13224,N_13181,N_13105);
nand U13225 (N_13225,N_13189,N_13050);
nand U13226 (N_13226,N_13116,N_13078);
nor U13227 (N_13227,N_13136,N_13088);
nor U13228 (N_13228,N_13191,N_13029);
xnor U13229 (N_13229,N_13103,N_13164);
xnor U13230 (N_13230,N_13043,N_13133);
nand U13231 (N_13231,N_13052,N_13187);
or U13232 (N_13232,N_13129,N_13020);
xor U13233 (N_13233,N_13081,N_13057);
or U13234 (N_13234,N_13006,N_13039);
and U13235 (N_13235,N_13074,N_13067);
or U13236 (N_13236,N_13085,N_13028);
nor U13237 (N_13237,N_13046,N_13058);
or U13238 (N_13238,N_13182,N_13055);
xor U13239 (N_13239,N_13118,N_13047);
xor U13240 (N_13240,N_13111,N_13172);
nand U13241 (N_13241,N_13149,N_13027);
nor U13242 (N_13242,N_13184,N_13110);
xor U13243 (N_13243,N_13173,N_13185);
nand U13244 (N_13244,N_13093,N_13180);
nand U13245 (N_13245,N_13089,N_13004);
or U13246 (N_13246,N_13044,N_13139);
or U13247 (N_13247,N_13168,N_13195);
nor U13248 (N_13248,N_13099,N_13021);
or U13249 (N_13249,N_13179,N_13092);
or U13250 (N_13250,N_13176,N_13061);
and U13251 (N_13251,N_13019,N_13183);
and U13252 (N_13252,N_13068,N_13148);
or U13253 (N_13253,N_13109,N_13102);
nor U13254 (N_13254,N_13013,N_13003);
or U13255 (N_13255,N_13154,N_13114);
nor U13256 (N_13256,N_13011,N_13128);
xor U13257 (N_13257,N_13192,N_13091);
nor U13258 (N_13258,N_13051,N_13012);
or U13259 (N_13259,N_13035,N_13010);
nor U13260 (N_13260,N_13009,N_13077);
nand U13261 (N_13261,N_13065,N_13060);
nand U13262 (N_13262,N_13095,N_13045);
and U13263 (N_13263,N_13036,N_13005);
or U13264 (N_13264,N_13042,N_13071);
xor U13265 (N_13265,N_13108,N_13124);
nor U13266 (N_13266,N_13080,N_13025);
or U13267 (N_13267,N_13120,N_13175);
and U13268 (N_13268,N_13022,N_13017);
or U13269 (N_13269,N_13007,N_13196);
nor U13270 (N_13270,N_13157,N_13023);
xor U13271 (N_13271,N_13158,N_13131);
xor U13272 (N_13272,N_13079,N_13100);
xnor U13273 (N_13273,N_13040,N_13070);
nand U13274 (N_13274,N_13163,N_13032);
xnor U13275 (N_13275,N_13159,N_13016);
nand U13276 (N_13276,N_13031,N_13166);
nand U13277 (N_13277,N_13170,N_13130);
and U13278 (N_13278,N_13177,N_13066);
nand U13279 (N_13279,N_13041,N_13059);
and U13280 (N_13280,N_13026,N_13199);
and U13281 (N_13281,N_13112,N_13104);
or U13282 (N_13282,N_13087,N_13053);
or U13283 (N_13283,N_13155,N_13132);
nand U13284 (N_13284,N_13084,N_13069);
nand U13285 (N_13285,N_13197,N_13142);
nor U13286 (N_13286,N_13150,N_13001);
and U13287 (N_13287,N_13101,N_13174);
nand U13288 (N_13288,N_13083,N_13015);
xor U13289 (N_13289,N_13153,N_13123);
nor U13290 (N_13290,N_13038,N_13113);
and U13291 (N_13291,N_13033,N_13121);
nor U13292 (N_13292,N_13127,N_13063);
or U13293 (N_13293,N_13161,N_13090);
and U13294 (N_13294,N_13064,N_13137);
or U13295 (N_13295,N_13082,N_13034);
and U13296 (N_13296,N_13056,N_13106);
or U13297 (N_13297,N_13119,N_13135);
nand U13298 (N_13298,N_13086,N_13037);
xor U13299 (N_13299,N_13008,N_13186);
or U13300 (N_13300,N_13092,N_13013);
xor U13301 (N_13301,N_13076,N_13177);
and U13302 (N_13302,N_13102,N_13140);
and U13303 (N_13303,N_13149,N_13018);
nand U13304 (N_13304,N_13070,N_13075);
and U13305 (N_13305,N_13074,N_13134);
and U13306 (N_13306,N_13124,N_13192);
nor U13307 (N_13307,N_13094,N_13197);
nand U13308 (N_13308,N_13088,N_13133);
or U13309 (N_13309,N_13156,N_13097);
and U13310 (N_13310,N_13011,N_13019);
xor U13311 (N_13311,N_13126,N_13128);
nor U13312 (N_13312,N_13143,N_13010);
xor U13313 (N_13313,N_13190,N_13160);
or U13314 (N_13314,N_13155,N_13030);
or U13315 (N_13315,N_13116,N_13051);
nor U13316 (N_13316,N_13009,N_13085);
or U13317 (N_13317,N_13049,N_13153);
xnor U13318 (N_13318,N_13143,N_13186);
nand U13319 (N_13319,N_13070,N_13000);
nor U13320 (N_13320,N_13007,N_13066);
and U13321 (N_13321,N_13119,N_13066);
nand U13322 (N_13322,N_13038,N_13089);
nand U13323 (N_13323,N_13079,N_13072);
nand U13324 (N_13324,N_13046,N_13028);
nand U13325 (N_13325,N_13054,N_13034);
or U13326 (N_13326,N_13032,N_13132);
nor U13327 (N_13327,N_13144,N_13192);
or U13328 (N_13328,N_13014,N_13115);
xnor U13329 (N_13329,N_13021,N_13130);
nor U13330 (N_13330,N_13007,N_13059);
or U13331 (N_13331,N_13166,N_13005);
nand U13332 (N_13332,N_13001,N_13025);
and U13333 (N_13333,N_13097,N_13040);
xor U13334 (N_13334,N_13190,N_13175);
nor U13335 (N_13335,N_13105,N_13151);
or U13336 (N_13336,N_13018,N_13074);
or U13337 (N_13337,N_13002,N_13066);
or U13338 (N_13338,N_13137,N_13154);
nor U13339 (N_13339,N_13124,N_13198);
or U13340 (N_13340,N_13163,N_13029);
and U13341 (N_13341,N_13153,N_13010);
xor U13342 (N_13342,N_13104,N_13128);
xnor U13343 (N_13343,N_13130,N_13177);
or U13344 (N_13344,N_13100,N_13092);
nor U13345 (N_13345,N_13154,N_13171);
and U13346 (N_13346,N_13118,N_13074);
and U13347 (N_13347,N_13193,N_13160);
nor U13348 (N_13348,N_13128,N_13194);
nand U13349 (N_13349,N_13175,N_13041);
xor U13350 (N_13350,N_13000,N_13120);
and U13351 (N_13351,N_13148,N_13043);
or U13352 (N_13352,N_13150,N_13153);
nor U13353 (N_13353,N_13036,N_13079);
or U13354 (N_13354,N_13173,N_13104);
nor U13355 (N_13355,N_13098,N_13035);
or U13356 (N_13356,N_13165,N_13152);
xor U13357 (N_13357,N_13092,N_13111);
and U13358 (N_13358,N_13132,N_13090);
nand U13359 (N_13359,N_13115,N_13187);
nand U13360 (N_13360,N_13079,N_13185);
nor U13361 (N_13361,N_13043,N_13076);
or U13362 (N_13362,N_13055,N_13060);
xor U13363 (N_13363,N_13066,N_13184);
or U13364 (N_13364,N_13175,N_13036);
nor U13365 (N_13365,N_13084,N_13096);
or U13366 (N_13366,N_13026,N_13153);
or U13367 (N_13367,N_13105,N_13046);
nor U13368 (N_13368,N_13144,N_13146);
nand U13369 (N_13369,N_13067,N_13091);
nor U13370 (N_13370,N_13114,N_13039);
xnor U13371 (N_13371,N_13059,N_13028);
or U13372 (N_13372,N_13062,N_13100);
or U13373 (N_13373,N_13069,N_13095);
xnor U13374 (N_13374,N_13056,N_13151);
nand U13375 (N_13375,N_13143,N_13084);
nor U13376 (N_13376,N_13000,N_13107);
nand U13377 (N_13377,N_13015,N_13071);
xor U13378 (N_13378,N_13037,N_13139);
nand U13379 (N_13379,N_13058,N_13050);
nand U13380 (N_13380,N_13134,N_13017);
nor U13381 (N_13381,N_13169,N_13191);
nand U13382 (N_13382,N_13011,N_13101);
xnor U13383 (N_13383,N_13181,N_13108);
or U13384 (N_13384,N_13023,N_13172);
nand U13385 (N_13385,N_13045,N_13054);
xor U13386 (N_13386,N_13066,N_13014);
xor U13387 (N_13387,N_13107,N_13080);
nor U13388 (N_13388,N_13135,N_13107);
nand U13389 (N_13389,N_13118,N_13116);
nor U13390 (N_13390,N_13109,N_13126);
nor U13391 (N_13391,N_13138,N_13160);
xor U13392 (N_13392,N_13154,N_13113);
nand U13393 (N_13393,N_13100,N_13195);
nand U13394 (N_13394,N_13066,N_13116);
or U13395 (N_13395,N_13161,N_13177);
xor U13396 (N_13396,N_13011,N_13198);
xnor U13397 (N_13397,N_13152,N_13040);
or U13398 (N_13398,N_13144,N_13062);
xnor U13399 (N_13399,N_13171,N_13100);
nor U13400 (N_13400,N_13282,N_13247);
or U13401 (N_13401,N_13263,N_13276);
nand U13402 (N_13402,N_13296,N_13298);
nor U13403 (N_13403,N_13229,N_13277);
nor U13404 (N_13404,N_13381,N_13346);
nand U13405 (N_13405,N_13215,N_13238);
or U13406 (N_13406,N_13332,N_13254);
nand U13407 (N_13407,N_13287,N_13274);
xor U13408 (N_13408,N_13278,N_13371);
or U13409 (N_13409,N_13375,N_13271);
and U13410 (N_13410,N_13377,N_13290);
nand U13411 (N_13411,N_13201,N_13295);
or U13412 (N_13412,N_13249,N_13213);
nand U13413 (N_13413,N_13361,N_13272);
and U13414 (N_13414,N_13344,N_13258);
or U13415 (N_13415,N_13235,N_13242);
nor U13416 (N_13416,N_13368,N_13341);
nand U13417 (N_13417,N_13246,N_13210);
and U13418 (N_13418,N_13357,N_13310);
nor U13419 (N_13419,N_13208,N_13364);
or U13420 (N_13420,N_13330,N_13230);
xor U13421 (N_13421,N_13345,N_13305);
or U13422 (N_13422,N_13264,N_13259);
nand U13423 (N_13423,N_13252,N_13214);
nor U13424 (N_13424,N_13311,N_13244);
nand U13425 (N_13425,N_13233,N_13237);
nand U13426 (N_13426,N_13321,N_13260);
and U13427 (N_13427,N_13343,N_13394);
nand U13428 (N_13428,N_13232,N_13391);
nand U13429 (N_13429,N_13337,N_13280);
or U13430 (N_13430,N_13307,N_13319);
nor U13431 (N_13431,N_13216,N_13382);
or U13432 (N_13432,N_13338,N_13253);
and U13433 (N_13433,N_13224,N_13358);
xnor U13434 (N_13434,N_13279,N_13331);
or U13435 (N_13435,N_13306,N_13302);
and U13436 (N_13436,N_13241,N_13348);
and U13437 (N_13437,N_13262,N_13309);
nand U13438 (N_13438,N_13202,N_13316);
nand U13439 (N_13439,N_13251,N_13362);
xnor U13440 (N_13440,N_13301,N_13267);
nor U13441 (N_13441,N_13236,N_13209);
xnor U13442 (N_13442,N_13312,N_13303);
and U13443 (N_13443,N_13227,N_13203);
nor U13444 (N_13444,N_13335,N_13231);
nand U13445 (N_13445,N_13388,N_13389);
or U13446 (N_13446,N_13286,N_13370);
or U13447 (N_13447,N_13320,N_13373);
or U13448 (N_13448,N_13217,N_13392);
nand U13449 (N_13449,N_13207,N_13220);
xnor U13450 (N_13450,N_13270,N_13355);
nor U13451 (N_13451,N_13376,N_13339);
and U13452 (N_13452,N_13265,N_13340);
and U13453 (N_13453,N_13349,N_13322);
or U13454 (N_13454,N_13275,N_13299);
and U13455 (N_13455,N_13378,N_13387);
nor U13456 (N_13456,N_13356,N_13256);
xnor U13457 (N_13457,N_13369,N_13334);
and U13458 (N_13458,N_13300,N_13329);
or U13459 (N_13459,N_13399,N_13308);
nor U13460 (N_13460,N_13313,N_13284);
xor U13461 (N_13461,N_13204,N_13297);
xnor U13462 (N_13462,N_13365,N_13360);
or U13463 (N_13463,N_13315,N_13380);
or U13464 (N_13464,N_13385,N_13283);
nor U13465 (N_13465,N_13292,N_13269);
or U13466 (N_13466,N_13323,N_13205);
xor U13467 (N_13467,N_13317,N_13383);
nor U13468 (N_13468,N_13354,N_13386);
nand U13469 (N_13469,N_13239,N_13390);
nand U13470 (N_13470,N_13366,N_13359);
and U13471 (N_13471,N_13342,N_13333);
xor U13472 (N_13472,N_13384,N_13225);
and U13473 (N_13473,N_13268,N_13218);
and U13474 (N_13474,N_13367,N_13223);
nor U13475 (N_13475,N_13248,N_13245);
nand U13476 (N_13476,N_13326,N_13293);
and U13477 (N_13477,N_13327,N_13395);
nor U13478 (N_13478,N_13200,N_13336);
nor U13479 (N_13479,N_13372,N_13324);
nand U13480 (N_13480,N_13211,N_13398);
nor U13481 (N_13481,N_13234,N_13240);
nor U13482 (N_13482,N_13288,N_13273);
and U13483 (N_13483,N_13351,N_13289);
and U13484 (N_13484,N_13257,N_13285);
or U13485 (N_13485,N_13226,N_13393);
and U13486 (N_13486,N_13347,N_13250);
nand U13487 (N_13487,N_13325,N_13379);
xnor U13488 (N_13488,N_13219,N_13291);
and U13489 (N_13489,N_13222,N_13397);
xor U13490 (N_13490,N_13228,N_13294);
and U13491 (N_13491,N_13374,N_13281);
nand U13492 (N_13492,N_13350,N_13255);
and U13493 (N_13493,N_13314,N_13221);
and U13494 (N_13494,N_13266,N_13353);
nor U13495 (N_13495,N_13206,N_13304);
xor U13496 (N_13496,N_13352,N_13212);
xor U13497 (N_13497,N_13243,N_13318);
nand U13498 (N_13498,N_13261,N_13328);
or U13499 (N_13499,N_13396,N_13363);
nand U13500 (N_13500,N_13251,N_13277);
or U13501 (N_13501,N_13303,N_13258);
nand U13502 (N_13502,N_13309,N_13279);
or U13503 (N_13503,N_13231,N_13338);
nor U13504 (N_13504,N_13237,N_13362);
or U13505 (N_13505,N_13286,N_13332);
nand U13506 (N_13506,N_13302,N_13303);
nand U13507 (N_13507,N_13211,N_13204);
nor U13508 (N_13508,N_13385,N_13252);
and U13509 (N_13509,N_13201,N_13371);
or U13510 (N_13510,N_13395,N_13247);
nand U13511 (N_13511,N_13304,N_13354);
and U13512 (N_13512,N_13226,N_13250);
and U13513 (N_13513,N_13288,N_13218);
and U13514 (N_13514,N_13286,N_13285);
or U13515 (N_13515,N_13317,N_13246);
xnor U13516 (N_13516,N_13314,N_13317);
nand U13517 (N_13517,N_13255,N_13261);
nor U13518 (N_13518,N_13293,N_13226);
nand U13519 (N_13519,N_13328,N_13215);
nand U13520 (N_13520,N_13269,N_13301);
or U13521 (N_13521,N_13241,N_13380);
nor U13522 (N_13522,N_13235,N_13219);
or U13523 (N_13523,N_13209,N_13343);
or U13524 (N_13524,N_13393,N_13256);
nor U13525 (N_13525,N_13237,N_13311);
or U13526 (N_13526,N_13225,N_13320);
nand U13527 (N_13527,N_13229,N_13294);
nand U13528 (N_13528,N_13364,N_13299);
or U13529 (N_13529,N_13262,N_13338);
or U13530 (N_13530,N_13353,N_13367);
xor U13531 (N_13531,N_13368,N_13330);
xor U13532 (N_13532,N_13257,N_13304);
and U13533 (N_13533,N_13361,N_13295);
nand U13534 (N_13534,N_13233,N_13334);
nor U13535 (N_13535,N_13317,N_13284);
or U13536 (N_13536,N_13310,N_13349);
and U13537 (N_13537,N_13291,N_13290);
and U13538 (N_13538,N_13214,N_13311);
xor U13539 (N_13539,N_13339,N_13258);
nand U13540 (N_13540,N_13330,N_13294);
and U13541 (N_13541,N_13335,N_13291);
and U13542 (N_13542,N_13273,N_13237);
and U13543 (N_13543,N_13319,N_13302);
nand U13544 (N_13544,N_13239,N_13370);
xor U13545 (N_13545,N_13219,N_13329);
nand U13546 (N_13546,N_13261,N_13322);
or U13547 (N_13547,N_13331,N_13266);
xnor U13548 (N_13548,N_13292,N_13264);
xnor U13549 (N_13549,N_13303,N_13361);
nand U13550 (N_13550,N_13210,N_13319);
nor U13551 (N_13551,N_13274,N_13253);
nand U13552 (N_13552,N_13378,N_13238);
or U13553 (N_13553,N_13336,N_13226);
and U13554 (N_13554,N_13399,N_13260);
or U13555 (N_13555,N_13355,N_13247);
nand U13556 (N_13556,N_13355,N_13388);
or U13557 (N_13557,N_13248,N_13265);
nand U13558 (N_13558,N_13296,N_13365);
nand U13559 (N_13559,N_13372,N_13266);
nand U13560 (N_13560,N_13385,N_13286);
and U13561 (N_13561,N_13300,N_13334);
xnor U13562 (N_13562,N_13235,N_13379);
nand U13563 (N_13563,N_13349,N_13365);
and U13564 (N_13564,N_13395,N_13289);
and U13565 (N_13565,N_13276,N_13211);
or U13566 (N_13566,N_13353,N_13361);
nor U13567 (N_13567,N_13282,N_13292);
nor U13568 (N_13568,N_13243,N_13219);
xor U13569 (N_13569,N_13267,N_13321);
xnor U13570 (N_13570,N_13207,N_13270);
and U13571 (N_13571,N_13237,N_13325);
nand U13572 (N_13572,N_13313,N_13380);
or U13573 (N_13573,N_13223,N_13272);
and U13574 (N_13574,N_13273,N_13255);
nor U13575 (N_13575,N_13344,N_13398);
nor U13576 (N_13576,N_13291,N_13390);
and U13577 (N_13577,N_13220,N_13350);
and U13578 (N_13578,N_13380,N_13266);
nand U13579 (N_13579,N_13337,N_13335);
and U13580 (N_13580,N_13391,N_13367);
nand U13581 (N_13581,N_13264,N_13301);
xor U13582 (N_13582,N_13201,N_13302);
nor U13583 (N_13583,N_13253,N_13233);
and U13584 (N_13584,N_13276,N_13384);
nor U13585 (N_13585,N_13304,N_13332);
xnor U13586 (N_13586,N_13329,N_13302);
and U13587 (N_13587,N_13387,N_13328);
xor U13588 (N_13588,N_13283,N_13265);
nand U13589 (N_13589,N_13242,N_13369);
xnor U13590 (N_13590,N_13268,N_13315);
nor U13591 (N_13591,N_13363,N_13232);
nor U13592 (N_13592,N_13229,N_13373);
or U13593 (N_13593,N_13335,N_13252);
and U13594 (N_13594,N_13235,N_13363);
or U13595 (N_13595,N_13205,N_13387);
or U13596 (N_13596,N_13388,N_13385);
xor U13597 (N_13597,N_13291,N_13387);
nand U13598 (N_13598,N_13283,N_13242);
and U13599 (N_13599,N_13218,N_13260);
xnor U13600 (N_13600,N_13569,N_13513);
and U13601 (N_13601,N_13438,N_13573);
or U13602 (N_13602,N_13499,N_13424);
and U13603 (N_13603,N_13530,N_13509);
and U13604 (N_13604,N_13577,N_13588);
xor U13605 (N_13605,N_13554,N_13437);
nand U13606 (N_13606,N_13562,N_13504);
or U13607 (N_13607,N_13474,N_13524);
xnor U13608 (N_13608,N_13548,N_13429);
nor U13609 (N_13609,N_13461,N_13512);
nand U13610 (N_13610,N_13511,N_13401);
nor U13611 (N_13611,N_13542,N_13468);
nand U13612 (N_13612,N_13455,N_13431);
or U13613 (N_13613,N_13518,N_13586);
and U13614 (N_13614,N_13458,N_13583);
xnor U13615 (N_13615,N_13430,N_13564);
and U13616 (N_13616,N_13568,N_13405);
or U13617 (N_13617,N_13408,N_13559);
nand U13618 (N_13618,N_13423,N_13479);
or U13619 (N_13619,N_13498,N_13400);
and U13620 (N_13620,N_13435,N_13407);
and U13621 (N_13621,N_13485,N_13445);
and U13622 (N_13622,N_13549,N_13507);
xor U13623 (N_13623,N_13517,N_13574);
and U13624 (N_13624,N_13403,N_13587);
xnor U13625 (N_13625,N_13506,N_13529);
and U13626 (N_13626,N_13589,N_13522);
or U13627 (N_13627,N_13567,N_13576);
or U13628 (N_13628,N_13497,N_13417);
or U13629 (N_13629,N_13406,N_13557);
or U13630 (N_13630,N_13457,N_13428);
nor U13631 (N_13631,N_13415,N_13436);
and U13632 (N_13632,N_13402,N_13503);
and U13633 (N_13633,N_13515,N_13508);
and U13634 (N_13634,N_13448,N_13416);
xor U13635 (N_13635,N_13502,N_13464);
xnor U13636 (N_13636,N_13533,N_13545);
xor U13637 (N_13637,N_13531,N_13505);
and U13638 (N_13638,N_13476,N_13496);
and U13639 (N_13639,N_13555,N_13527);
and U13640 (N_13640,N_13475,N_13447);
xnor U13641 (N_13641,N_13411,N_13450);
nand U13642 (N_13642,N_13422,N_13546);
nand U13643 (N_13643,N_13467,N_13595);
xor U13644 (N_13644,N_13456,N_13584);
xnor U13645 (N_13645,N_13570,N_13553);
nand U13646 (N_13646,N_13493,N_13451);
nor U13647 (N_13647,N_13528,N_13442);
xor U13648 (N_13648,N_13463,N_13578);
or U13649 (N_13649,N_13571,N_13520);
nor U13650 (N_13650,N_13414,N_13536);
or U13651 (N_13651,N_13452,N_13460);
and U13652 (N_13652,N_13566,N_13532);
and U13653 (N_13653,N_13472,N_13540);
nor U13654 (N_13654,N_13477,N_13488);
nor U13655 (N_13655,N_13537,N_13597);
nor U13656 (N_13656,N_13427,N_13575);
and U13657 (N_13657,N_13421,N_13500);
nand U13658 (N_13658,N_13501,N_13550);
nor U13659 (N_13659,N_13565,N_13534);
xnor U13660 (N_13660,N_13523,N_13409);
xnor U13661 (N_13661,N_13551,N_13579);
or U13662 (N_13662,N_13592,N_13572);
nor U13663 (N_13663,N_13494,N_13593);
nor U13664 (N_13664,N_13444,N_13454);
and U13665 (N_13665,N_13558,N_13591);
xor U13666 (N_13666,N_13469,N_13439);
nand U13667 (N_13667,N_13539,N_13466);
or U13668 (N_13668,N_13516,N_13543);
and U13669 (N_13669,N_13419,N_13561);
or U13670 (N_13670,N_13514,N_13560);
and U13671 (N_13671,N_13432,N_13487);
or U13672 (N_13672,N_13470,N_13510);
nand U13673 (N_13673,N_13473,N_13526);
nor U13674 (N_13674,N_13491,N_13420);
and U13675 (N_13675,N_13596,N_13547);
and U13676 (N_13676,N_13525,N_13480);
nor U13677 (N_13677,N_13433,N_13412);
nand U13678 (N_13678,N_13478,N_13598);
nor U13679 (N_13679,N_13599,N_13492);
and U13680 (N_13680,N_13544,N_13426);
and U13681 (N_13681,N_13410,N_13495);
xnor U13682 (N_13682,N_13541,N_13580);
nor U13683 (N_13683,N_13582,N_13489);
or U13684 (N_13684,N_13446,N_13585);
nor U13685 (N_13685,N_13471,N_13425);
or U13686 (N_13686,N_13404,N_13453);
and U13687 (N_13687,N_13443,N_13594);
xor U13688 (N_13688,N_13481,N_13434);
nand U13689 (N_13689,N_13590,N_13490);
nand U13690 (N_13690,N_13459,N_13552);
nor U13691 (N_13691,N_13418,N_13519);
xnor U13692 (N_13692,N_13449,N_13440);
nor U13693 (N_13693,N_13484,N_13538);
nor U13694 (N_13694,N_13563,N_13486);
or U13695 (N_13695,N_13556,N_13465);
xnor U13696 (N_13696,N_13535,N_13483);
and U13697 (N_13697,N_13521,N_13413);
xnor U13698 (N_13698,N_13441,N_13482);
or U13699 (N_13699,N_13581,N_13462);
and U13700 (N_13700,N_13402,N_13598);
and U13701 (N_13701,N_13576,N_13555);
xor U13702 (N_13702,N_13544,N_13587);
nor U13703 (N_13703,N_13404,N_13579);
xnor U13704 (N_13704,N_13422,N_13515);
nor U13705 (N_13705,N_13585,N_13518);
nand U13706 (N_13706,N_13572,N_13480);
nor U13707 (N_13707,N_13411,N_13408);
nor U13708 (N_13708,N_13562,N_13518);
and U13709 (N_13709,N_13588,N_13535);
xor U13710 (N_13710,N_13494,N_13419);
xnor U13711 (N_13711,N_13484,N_13471);
xnor U13712 (N_13712,N_13587,N_13415);
nor U13713 (N_13713,N_13475,N_13578);
or U13714 (N_13714,N_13416,N_13459);
or U13715 (N_13715,N_13461,N_13580);
or U13716 (N_13716,N_13599,N_13561);
nand U13717 (N_13717,N_13524,N_13466);
nor U13718 (N_13718,N_13466,N_13590);
nor U13719 (N_13719,N_13446,N_13475);
and U13720 (N_13720,N_13434,N_13535);
or U13721 (N_13721,N_13542,N_13445);
xor U13722 (N_13722,N_13469,N_13584);
or U13723 (N_13723,N_13592,N_13496);
nor U13724 (N_13724,N_13516,N_13496);
and U13725 (N_13725,N_13486,N_13550);
nor U13726 (N_13726,N_13508,N_13481);
nand U13727 (N_13727,N_13471,N_13566);
nor U13728 (N_13728,N_13520,N_13542);
nor U13729 (N_13729,N_13463,N_13574);
or U13730 (N_13730,N_13400,N_13448);
nand U13731 (N_13731,N_13576,N_13537);
or U13732 (N_13732,N_13504,N_13471);
and U13733 (N_13733,N_13524,N_13558);
or U13734 (N_13734,N_13447,N_13457);
xnor U13735 (N_13735,N_13500,N_13483);
nor U13736 (N_13736,N_13552,N_13443);
xnor U13737 (N_13737,N_13410,N_13484);
nor U13738 (N_13738,N_13485,N_13522);
and U13739 (N_13739,N_13546,N_13493);
nor U13740 (N_13740,N_13534,N_13442);
nand U13741 (N_13741,N_13470,N_13526);
nor U13742 (N_13742,N_13420,N_13543);
nor U13743 (N_13743,N_13555,N_13494);
nor U13744 (N_13744,N_13414,N_13438);
and U13745 (N_13745,N_13468,N_13532);
or U13746 (N_13746,N_13454,N_13417);
and U13747 (N_13747,N_13537,N_13440);
nand U13748 (N_13748,N_13544,N_13416);
and U13749 (N_13749,N_13536,N_13539);
xnor U13750 (N_13750,N_13427,N_13480);
nand U13751 (N_13751,N_13403,N_13554);
nor U13752 (N_13752,N_13583,N_13460);
or U13753 (N_13753,N_13592,N_13413);
and U13754 (N_13754,N_13579,N_13463);
nand U13755 (N_13755,N_13526,N_13481);
xnor U13756 (N_13756,N_13423,N_13520);
or U13757 (N_13757,N_13493,N_13599);
nor U13758 (N_13758,N_13429,N_13470);
nand U13759 (N_13759,N_13551,N_13467);
or U13760 (N_13760,N_13584,N_13428);
and U13761 (N_13761,N_13543,N_13511);
or U13762 (N_13762,N_13567,N_13514);
xor U13763 (N_13763,N_13521,N_13425);
or U13764 (N_13764,N_13450,N_13532);
or U13765 (N_13765,N_13550,N_13543);
or U13766 (N_13766,N_13599,N_13405);
xor U13767 (N_13767,N_13546,N_13427);
nor U13768 (N_13768,N_13511,N_13432);
nand U13769 (N_13769,N_13427,N_13596);
and U13770 (N_13770,N_13517,N_13538);
nor U13771 (N_13771,N_13552,N_13592);
or U13772 (N_13772,N_13474,N_13456);
and U13773 (N_13773,N_13500,N_13405);
nand U13774 (N_13774,N_13487,N_13453);
or U13775 (N_13775,N_13551,N_13428);
xnor U13776 (N_13776,N_13421,N_13527);
nand U13777 (N_13777,N_13510,N_13535);
nand U13778 (N_13778,N_13543,N_13483);
nand U13779 (N_13779,N_13444,N_13422);
nor U13780 (N_13780,N_13432,N_13549);
and U13781 (N_13781,N_13501,N_13542);
xnor U13782 (N_13782,N_13511,N_13501);
xnor U13783 (N_13783,N_13437,N_13571);
xor U13784 (N_13784,N_13578,N_13598);
xnor U13785 (N_13785,N_13564,N_13509);
and U13786 (N_13786,N_13408,N_13578);
nor U13787 (N_13787,N_13533,N_13591);
and U13788 (N_13788,N_13490,N_13517);
nor U13789 (N_13789,N_13493,N_13499);
nand U13790 (N_13790,N_13491,N_13572);
xor U13791 (N_13791,N_13592,N_13500);
nand U13792 (N_13792,N_13590,N_13586);
xor U13793 (N_13793,N_13496,N_13411);
nor U13794 (N_13794,N_13421,N_13455);
nand U13795 (N_13795,N_13576,N_13438);
or U13796 (N_13796,N_13581,N_13533);
nor U13797 (N_13797,N_13598,N_13584);
nand U13798 (N_13798,N_13545,N_13491);
nand U13799 (N_13799,N_13477,N_13472);
xnor U13800 (N_13800,N_13791,N_13604);
nand U13801 (N_13801,N_13730,N_13673);
and U13802 (N_13802,N_13734,N_13720);
xor U13803 (N_13803,N_13628,N_13721);
or U13804 (N_13804,N_13636,N_13697);
or U13805 (N_13805,N_13736,N_13646);
and U13806 (N_13806,N_13614,N_13744);
nand U13807 (N_13807,N_13603,N_13620);
or U13808 (N_13808,N_13626,N_13774);
nor U13809 (N_13809,N_13704,N_13715);
and U13810 (N_13810,N_13635,N_13638);
and U13811 (N_13811,N_13768,N_13747);
and U13812 (N_13812,N_13668,N_13687);
nor U13813 (N_13813,N_13759,N_13743);
and U13814 (N_13814,N_13776,N_13727);
xor U13815 (N_13815,N_13784,N_13731);
xnor U13816 (N_13816,N_13698,N_13672);
or U13817 (N_13817,N_13792,N_13773);
xnor U13818 (N_13818,N_13642,N_13685);
xnor U13819 (N_13819,N_13653,N_13767);
nand U13820 (N_13820,N_13650,N_13739);
or U13821 (N_13821,N_13610,N_13797);
or U13822 (N_13822,N_13782,N_13724);
and U13823 (N_13823,N_13651,N_13667);
or U13824 (N_13824,N_13600,N_13750);
or U13825 (N_13825,N_13758,N_13681);
and U13826 (N_13826,N_13694,N_13711);
xnor U13827 (N_13827,N_13796,N_13717);
or U13828 (N_13828,N_13772,N_13779);
xor U13829 (N_13829,N_13793,N_13798);
nand U13830 (N_13830,N_13702,N_13786);
nand U13831 (N_13831,N_13765,N_13611);
and U13832 (N_13832,N_13787,N_13749);
or U13833 (N_13833,N_13630,N_13669);
and U13834 (N_13834,N_13795,N_13617);
or U13835 (N_13835,N_13757,N_13643);
nand U13836 (N_13836,N_13741,N_13714);
nand U13837 (N_13837,N_13762,N_13686);
nor U13838 (N_13838,N_13608,N_13726);
xor U13839 (N_13839,N_13783,N_13718);
or U13840 (N_13840,N_13683,N_13612);
and U13841 (N_13841,N_13671,N_13602);
nand U13842 (N_13842,N_13699,N_13754);
xor U13843 (N_13843,N_13645,N_13661);
or U13844 (N_13844,N_13615,N_13679);
xor U13845 (N_13845,N_13627,N_13708);
xnor U13846 (N_13846,N_13794,N_13729);
and U13847 (N_13847,N_13735,N_13622);
and U13848 (N_13848,N_13664,N_13799);
and U13849 (N_13849,N_13690,N_13771);
and U13850 (N_13850,N_13705,N_13732);
nor U13851 (N_13851,N_13737,N_13745);
or U13852 (N_13852,N_13647,N_13780);
nand U13853 (N_13853,N_13701,N_13742);
or U13854 (N_13854,N_13616,N_13657);
nor U13855 (N_13855,N_13631,N_13781);
xor U13856 (N_13856,N_13706,N_13733);
nand U13857 (N_13857,N_13658,N_13777);
nor U13858 (N_13858,N_13625,N_13644);
xnor U13859 (N_13859,N_13695,N_13740);
nand U13860 (N_13860,N_13665,N_13723);
nor U13861 (N_13861,N_13623,N_13663);
nor U13862 (N_13862,N_13656,N_13738);
nand U13863 (N_13863,N_13713,N_13674);
and U13864 (N_13864,N_13649,N_13632);
nand U13865 (N_13865,N_13639,N_13682);
xnor U13866 (N_13866,N_13619,N_13692);
nand U13867 (N_13867,N_13637,N_13609);
and U13868 (N_13868,N_13752,N_13618);
and U13869 (N_13869,N_13677,N_13652);
nand U13870 (N_13870,N_13725,N_13689);
or U13871 (N_13871,N_13670,N_13696);
xor U13872 (N_13872,N_13753,N_13778);
and U13873 (N_13873,N_13760,N_13709);
xor U13874 (N_13874,N_13654,N_13751);
nand U13875 (N_13875,N_13691,N_13666);
and U13876 (N_13876,N_13660,N_13640);
xor U13877 (N_13877,N_13703,N_13641);
or U13878 (N_13878,N_13728,N_13716);
and U13879 (N_13879,N_13722,N_13710);
or U13880 (N_13880,N_13756,N_13748);
xor U13881 (N_13881,N_13684,N_13648);
nand U13882 (N_13882,N_13675,N_13688);
or U13883 (N_13883,N_13770,N_13790);
xor U13884 (N_13884,N_13761,N_13693);
and U13885 (N_13885,N_13769,N_13719);
nand U13886 (N_13886,N_13707,N_13788);
xor U13887 (N_13887,N_13789,N_13712);
nand U13888 (N_13888,N_13700,N_13755);
xnor U13889 (N_13889,N_13680,N_13775);
nor U13890 (N_13890,N_13766,N_13659);
or U13891 (N_13891,N_13634,N_13764);
xor U13892 (N_13892,N_13629,N_13607);
or U13893 (N_13893,N_13678,N_13601);
or U13894 (N_13894,N_13633,N_13605);
or U13895 (N_13895,N_13785,N_13655);
xnor U13896 (N_13896,N_13621,N_13676);
or U13897 (N_13897,N_13606,N_13763);
and U13898 (N_13898,N_13662,N_13613);
and U13899 (N_13899,N_13746,N_13624);
or U13900 (N_13900,N_13734,N_13778);
and U13901 (N_13901,N_13791,N_13698);
xnor U13902 (N_13902,N_13686,N_13638);
xnor U13903 (N_13903,N_13719,N_13775);
nor U13904 (N_13904,N_13774,N_13787);
and U13905 (N_13905,N_13633,N_13758);
and U13906 (N_13906,N_13711,N_13730);
nand U13907 (N_13907,N_13788,N_13710);
nor U13908 (N_13908,N_13704,N_13671);
nand U13909 (N_13909,N_13759,N_13638);
or U13910 (N_13910,N_13746,N_13702);
nor U13911 (N_13911,N_13662,N_13636);
xnor U13912 (N_13912,N_13751,N_13733);
or U13913 (N_13913,N_13701,N_13741);
nor U13914 (N_13914,N_13633,N_13704);
and U13915 (N_13915,N_13749,N_13799);
and U13916 (N_13916,N_13605,N_13781);
and U13917 (N_13917,N_13763,N_13732);
or U13918 (N_13918,N_13781,N_13613);
nand U13919 (N_13919,N_13616,N_13756);
and U13920 (N_13920,N_13791,N_13758);
and U13921 (N_13921,N_13709,N_13606);
xor U13922 (N_13922,N_13613,N_13752);
and U13923 (N_13923,N_13742,N_13653);
nor U13924 (N_13924,N_13653,N_13679);
and U13925 (N_13925,N_13688,N_13653);
and U13926 (N_13926,N_13779,N_13647);
or U13927 (N_13927,N_13679,N_13764);
and U13928 (N_13928,N_13605,N_13606);
or U13929 (N_13929,N_13645,N_13663);
or U13930 (N_13930,N_13631,N_13755);
or U13931 (N_13931,N_13736,N_13644);
xor U13932 (N_13932,N_13639,N_13631);
xnor U13933 (N_13933,N_13716,N_13765);
and U13934 (N_13934,N_13712,N_13772);
nand U13935 (N_13935,N_13645,N_13701);
or U13936 (N_13936,N_13735,N_13762);
and U13937 (N_13937,N_13602,N_13790);
nand U13938 (N_13938,N_13677,N_13635);
xor U13939 (N_13939,N_13684,N_13694);
xnor U13940 (N_13940,N_13628,N_13695);
nor U13941 (N_13941,N_13633,N_13780);
xnor U13942 (N_13942,N_13653,N_13745);
nand U13943 (N_13943,N_13605,N_13685);
nand U13944 (N_13944,N_13685,N_13798);
or U13945 (N_13945,N_13646,N_13677);
and U13946 (N_13946,N_13643,N_13707);
nor U13947 (N_13947,N_13680,N_13689);
or U13948 (N_13948,N_13727,N_13723);
xnor U13949 (N_13949,N_13710,N_13621);
and U13950 (N_13950,N_13749,N_13626);
or U13951 (N_13951,N_13621,N_13722);
and U13952 (N_13952,N_13735,N_13796);
nand U13953 (N_13953,N_13780,N_13602);
and U13954 (N_13954,N_13742,N_13678);
nor U13955 (N_13955,N_13659,N_13772);
xor U13956 (N_13956,N_13780,N_13661);
nand U13957 (N_13957,N_13677,N_13789);
and U13958 (N_13958,N_13778,N_13641);
or U13959 (N_13959,N_13615,N_13748);
xor U13960 (N_13960,N_13738,N_13652);
nand U13961 (N_13961,N_13775,N_13698);
xnor U13962 (N_13962,N_13612,N_13715);
or U13963 (N_13963,N_13798,N_13610);
xnor U13964 (N_13964,N_13693,N_13714);
and U13965 (N_13965,N_13774,N_13635);
nor U13966 (N_13966,N_13605,N_13696);
and U13967 (N_13967,N_13660,N_13688);
nand U13968 (N_13968,N_13614,N_13649);
or U13969 (N_13969,N_13734,N_13616);
or U13970 (N_13970,N_13689,N_13682);
and U13971 (N_13971,N_13625,N_13645);
or U13972 (N_13972,N_13697,N_13633);
nand U13973 (N_13973,N_13646,N_13639);
or U13974 (N_13974,N_13768,N_13664);
xnor U13975 (N_13975,N_13779,N_13734);
xor U13976 (N_13976,N_13768,N_13780);
or U13977 (N_13977,N_13622,N_13605);
xor U13978 (N_13978,N_13608,N_13668);
nand U13979 (N_13979,N_13787,N_13680);
nand U13980 (N_13980,N_13649,N_13765);
xor U13981 (N_13981,N_13653,N_13722);
nand U13982 (N_13982,N_13603,N_13735);
nand U13983 (N_13983,N_13656,N_13621);
and U13984 (N_13984,N_13656,N_13660);
and U13985 (N_13985,N_13702,N_13694);
or U13986 (N_13986,N_13631,N_13748);
nand U13987 (N_13987,N_13619,N_13702);
nor U13988 (N_13988,N_13672,N_13693);
xnor U13989 (N_13989,N_13734,N_13692);
nor U13990 (N_13990,N_13603,N_13623);
nand U13991 (N_13991,N_13665,N_13722);
xnor U13992 (N_13992,N_13622,N_13667);
nor U13993 (N_13993,N_13661,N_13791);
nand U13994 (N_13994,N_13628,N_13624);
xnor U13995 (N_13995,N_13603,N_13762);
and U13996 (N_13996,N_13695,N_13661);
nand U13997 (N_13997,N_13626,N_13715);
or U13998 (N_13998,N_13788,N_13678);
nor U13999 (N_13999,N_13619,N_13624);
xor U14000 (N_14000,N_13850,N_13887);
xnor U14001 (N_14001,N_13931,N_13870);
and U14002 (N_14002,N_13974,N_13920);
and U14003 (N_14003,N_13844,N_13873);
and U14004 (N_14004,N_13959,N_13990);
or U14005 (N_14005,N_13986,N_13951);
and U14006 (N_14006,N_13941,N_13992);
or U14007 (N_14007,N_13948,N_13968);
nor U14008 (N_14008,N_13852,N_13918);
or U14009 (N_14009,N_13814,N_13817);
and U14010 (N_14010,N_13864,N_13875);
and U14011 (N_14011,N_13988,N_13812);
nor U14012 (N_14012,N_13993,N_13881);
nor U14013 (N_14013,N_13947,N_13832);
or U14014 (N_14014,N_13804,N_13860);
nor U14015 (N_14015,N_13808,N_13859);
and U14016 (N_14016,N_13917,N_13954);
nor U14017 (N_14017,N_13910,N_13958);
and U14018 (N_14018,N_13802,N_13882);
or U14019 (N_14019,N_13806,N_13960);
nand U14020 (N_14020,N_13801,N_13924);
and U14021 (N_14021,N_13901,N_13907);
or U14022 (N_14022,N_13885,N_13983);
nand U14023 (N_14023,N_13807,N_13871);
nand U14024 (N_14024,N_13927,N_13841);
nor U14025 (N_14025,N_13865,N_13943);
xnor U14026 (N_14026,N_13888,N_13977);
xor U14027 (N_14027,N_13898,N_13833);
nor U14028 (N_14028,N_13953,N_13998);
xnor U14029 (N_14029,N_13851,N_13863);
and U14030 (N_14030,N_13830,N_13912);
xor U14031 (N_14031,N_13847,N_13827);
and U14032 (N_14032,N_13821,N_13899);
nor U14033 (N_14033,N_13890,N_13877);
or U14034 (N_14034,N_13957,N_13868);
xnor U14035 (N_14035,N_13837,N_13819);
or U14036 (N_14036,N_13962,N_13835);
nor U14037 (N_14037,N_13915,N_13858);
nor U14038 (N_14038,N_13862,N_13826);
nand U14039 (N_14039,N_13900,N_13816);
or U14040 (N_14040,N_13940,N_13911);
and U14041 (N_14041,N_13933,N_13896);
nor U14042 (N_14042,N_13934,N_13969);
and U14043 (N_14043,N_13999,N_13813);
nand U14044 (N_14044,N_13976,N_13800);
and U14045 (N_14045,N_13836,N_13903);
nor U14046 (N_14046,N_13884,N_13936);
and U14047 (N_14047,N_13922,N_13973);
and U14048 (N_14048,N_13838,N_13978);
or U14049 (N_14049,N_13989,N_13878);
nor U14050 (N_14050,N_13861,N_13942);
nor U14051 (N_14051,N_13815,N_13982);
nor U14052 (N_14052,N_13906,N_13995);
and U14053 (N_14053,N_13872,N_13949);
xnor U14054 (N_14054,N_13996,N_13856);
or U14055 (N_14055,N_13991,N_13913);
nand U14056 (N_14056,N_13939,N_13970);
or U14057 (N_14057,N_13874,N_13979);
nor U14058 (N_14058,N_13822,N_13975);
nand U14059 (N_14059,N_13803,N_13904);
xnor U14060 (N_14060,N_13916,N_13945);
nor U14061 (N_14061,N_13854,N_13955);
nand U14062 (N_14062,N_13902,N_13892);
or U14063 (N_14063,N_13805,N_13893);
xor U14064 (N_14064,N_13961,N_13842);
nand U14065 (N_14065,N_13925,N_13994);
and U14066 (N_14066,N_13937,N_13905);
or U14067 (N_14067,N_13981,N_13894);
and U14068 (N_14068,N_13883,N_13880);
or U14069 (N_14069,N_13853,N_13897);
nand U14070 (N_14070,N_13987,N_13971);
and U14071 (N_14071,N_13965,N_13810);
nand U14072 (N_14072,N_13818,N_13891);
xnor U14073 (N_14073,N_13908,N_13950);
xnor U14074 (N_14074,N_13849,N_13928);
nor U14075 (N_14075,N_13944,N_13825);
xnor U14076 (N_14076,N_13966,N_13895);
nand U14077 (N_14077,N_13930,N_13946);
xor U14078 (N_14078,N_13984,N_13811);
nor U14079 (N_14079,N_13926,N_13855);
or U14080 (N_14080,N_13840,N_13820);
and U14081 (N_14081,N_13831,N_13935);
xnor U14082 (N_14082,N_13829,N_13964);
or U14083 (N_14083,N_13980,N_13848);
and U14084 (N_14084,N_13839,N_13823);
nor U14085 (N_14085,N_13866,N_13889);
and U14086 (N_14086,N_13867,N_13809);
nand U14087 (N_14087,N_13919,N_13985);
nand U14088 (N_14088,N_13923,N_13843);
nor U14089 (N_14089,N_13909,N_13834);
nor U14090 (N_14090,N_13857,N_13929);
or U14091 (N_14091,N_13956,N_13886);
xor U14092 (N_14092,N_13952,N_13845);
or U14093 (N_14093,N_13869,N_13921);
nand U14094 (N_14094,N_13997,N_13846);
nand U14095 (N_14095,N_13828,N_13932);
or U14096 (N_14096,N_13824,N_13972);
or U14097 (N_14097,N_13967,N_13914);
and U14098 (N_14098,N_13876,N_13938);
or U14099 (N_14099,N_13879,N_13963);
nor U14100 (N_14100,N_13952,N_13842);
and U14101 (N_14101,N_13944,N_13855);
or U14102 (N_14102,N_13955,N_13917);
or U14103 (N_14103,N_13883,N_13865);
or U14104 (N_14104,N_13931,N_13932);
xor U14105 (N_14105,N_13924,N_13942);
xnor U14106 (N_14106,N_13949,N_13876);
and U14107 (N_14107,N_13858,N_13977);
or U14108 (N_14108,N_13898,N_13925);
or U14109 (N_14109,N_13942,N_13964);
nand U14110 (N_14110,N_13918,N_13988);
nand U14111 (N_14111,N_13976,N_13933);
nor U14112 (N_14112,N_13996,N_13898);
nand U14113 (N_14113,N_13808,N_13854);
or U14114 (N_14114,N_13832,N_13986);
and U14115 (N_14115,N_13868,N_13975);
or U14116 (N_14116,N_13954,N_13976);
or U14117 (N_14117,N_13930,N_13828);
or U14118 (N_14118,N_13942,N_13989);
xor U14119 (N_14119,N_13832,N_13985);
nor U14120 (N_14120,N_13938,N_13989);
or U14121 (N_14121,N_13838,N_13801);
nand U14122 (N_14122,N_13938,N_13909);
nand U14123 (N_14123,N_13908,N_13833);
nand U14124 (N_14124,N_13922,N_13804);
or U14125 (N_14125,N_13936,N_13899);
nand U14126 (N_14126,N_13831,N_13881);
nand U14127 (N_14127,N_13999,N_13986);
nand U14128 (N_14128,N_13805,N_13968);
or U14129 (N_14129,N_13969,N_13921);
and U14130 (N_14130,N_13916,N_13888);
or U14131 (N_14131,N_13806,N_13868);
or U14132 (N_14132,N_13936,N_13986);
or U14133 (N_14133,N_13928,N_13844);
xnor U14134 (N_14134,N_13838,N_13935);
xor U14135 (N_14135,N_13886,N_13917);
nor U14136 (N_14136,N_13809,N_13825);
nor U14137 (N_14137,N_13802,N_13804);
xor U14138 (N_14138,N_13833,N_13884);
or U14139 (N_14139,N_13952,N_13876);
xor U14140 (N_14140,N_13999,N_13994);
nand U14141 (N_14141,N_13978,N_13936);
nand U14142 (N_14142,N_13995,N_13877);
xnor U14143 (N_14143,N_13995,N_13896);
or U14144 (N_14144,N_13943,N_13983);
and U14145 (N_14145,N_13860,N_13808);
xor U14146 (N_14146,N_13878,N_13848);
and U14147 (N_14147,N_13842,N_13948);
and U14148 (N_14148,N_13800,N_13997);
or U14149 (N_14149,N_13882,N_13905);
xnor U14150 (N_14150,N_13883,N_13952);
nand U14151 (N_14151,N_13940,N_13839);
nand U14152 (N_14152,N_13975,N_13839);
nor U14153 (N_14153,N_13997,N_13907);
or U14154 (N_14154,N_13856,N_13971);
or U14155 (N_14155,N_13880,N_13955);
or U14156 (N_14156,N_13804,N_13876);
nor U14157 (N_14157,N_13853,N_13890);
nor U14158 (N_14158,N_13851,N_13922);
and U14159 (N_14159,N_13815,N_13996);
nor U14160 (N_14160,N_13822,N_13985);
nor U14161 (N_14161,N_13985,N_13895);
nor U14162 (N_14162,N_13987,N_13886);
xor U14163 (N_14163,N_13942,N_13911);
nor U14164 (N_14164,N_13973,N_13866);
nand U14165 (N_14165,N_13875,N_13959);
and U14166 (N_14166,N_13853,N_13841);
nand U14167 (N_14167,N_13856,N_13857);
and U14168 (N_14168,N_13840,N_13803);
and U14169 (N_14169,N_13953,N_13863);
nand U14170 (N_14170,N_13990,N_13938);
and U14171 (N_14171,N_13963,N_13973);
and U14172 (N_14172,N_13800,N_13856);
nor U14173 (N_14173,N_13897,N_13937);
nand U14174 (N_14174,N_13888,N_13852);
or U14175 (N_14175,N_13914,N_13996);
or U14176 (N_14176,N_13817,N_13952);
xnor U14177 (N_14177,N_13801,N_13951);
xor U14178 (N_14178,N_13921,N_13919);
and U14179 (N_14179,N_13993,N_13906);
nand U14180 (N_14180,N_13831,N_13839);
nor U14181 (N_14181,N_13906,N_13837);
or U14182 (N_14182,N_13855,N_13850);
nor U14183 (N_14183,N_13864,N_13812);
or U14184 (N_14184,N_13928,N_13813);
or U14185 (N_14185,N_13994,N_13969);
nor U14186 (N_14186,N_13828,N_13979);
nor U14187 (N_14187,N_13839,N_13993);
xor U14188 (N_14188,N_13997,N_13918);
and U14189 (N_14189,N_13990,N_13802);
xnor U14190 (N_14190,N_13923,N_13845);
nor U14191 (N_14191,N_13958,N_13887);
nand U14192 (N_14192,N_13960,N_13902);
nand U14193 (N_14193,N_13966,N_13891);
and U14194 (N_14194,N_13884,N_13886);
or U14195 (N_14195,N_13995,N_13850);
nor U14196 (N_14196,N_13954,N_13850);
nand U14197 (N_14197,N_13963,N_13827);
nor U14198 (N_14198,N_13915,N_13890);
nor U14199 (N_14199,N_13867,N_13886);
or U14200 (N_14200,N_14024,N_14195);
and U14201 (N_14201,N_14003,N_14156);
xnor U14202 (N_14202,N_14020,N_14180);
or U14203 (N_14203,N_14089,N_14187);
or U14204 (N_14204,N_14016,N_14033);
xnor U14205 (N_14205,N_14184,N_14196);
and U14206 (N_14206,N_14173,N_14080);
xor U14207 (N_14207,N_14158,N_14191);
nor U14208 (N_14208,N_14083,N_14039);
and U14209 (N_14209,N_14199,N_14120);
or U14210 (N_14210,N_14082,N_14185);
and U14211 (N_14211,N_14113,N_14155);
nand U14212 (N_14212,N_14028,N_14027);
xor U14213 (N_14213,N_14069,N_14143);
or U14214 (N_14214,N_14112,N_14059);
xnor U14215 (N_14215,N_14150,N_14002);
nor U14216 (N_14216,N_14161,N_14065);
nand U14217 (N_14217,N_14014,N_14122);
or U14218 (N_14218,N_14034,N_14148);
xor U14219 (N_14219,N_14124,N_14045);
xor U14220 (N_14220,N_14129,N_14179);
and U14221 (N_14221,N_14088,N_14031);
nor U14222 (N_14222,N_14183,N_14116);
or U14223 (N_14223,N_14070,N_14107);
or U14224 (N_14224,N_14073,N_14162);
and U14225 (N_14225,N_14035,N_14086);
and U14226 (N_14226,N_14093,N_14182);
nor U14227 (N_14227,N_14051,N_14167);
nand U14228 (N_14228,N_14101,N_14168);
nand U14229 (N_14229,N_14133,N_14140);
and U14230 (N_14230,N_14074,N_14063);
xnor U14231 (N_14231,N_14040,N_14165);
and U14232 (N_14232,N_14192,N_14068);
and U14233 (N_14233,N_14079,N_14160);
nor U14234 (N_14234,N_14021,N_14175);
or U14235 (N_14235,N_14006,N_14154);
xor U14236 (N_14236,N_14067,N_14009);
nand U14237 (N_14237,N_14139,N_14064);
and U14238 (N_14238,N_14055,N_14121);
or U14239 (N_14239,N_14011,N_14025);
xnor U14240 (N_14240,N_14110,N_14041);
or U14241 (N_14241,N_14166,N_14022);
or U14242 (N_14242,N_14001,N_14096);
nand U14243 (N_14243,N_14125,N_14057);
or U14244 (N_14244,N_14102,N_14012);
nand U14245 (N_14245,N_14193,N_14023);
nand U14246 (N_14246,N_14134,N_14157);
and U14247 (N_14247,N_14005,N_14037);
nor U14248 (N_14248,N_14013,N_14090);
nor U14249 (N_14249,N_14049,N_14015);
xnor U14250 (N_14250,N_14135,N_14106);
xnor U14251 (N_14251,N_14138,N_14131);
xnor U14252 (N_14252,N_14098,N_14109);
nor U14253 (N_14253,N_14117,N_14137);
nand U14254 (N_14254,N_14004,N_14078);
xnor U14255 (N_14255,N_14186,N_14111);
xor U14256 (N_14256,N_14099,N_14176);
and U14257 (N_14257,N_14050,N_14152);
or U14258 (N_14258,N_14164,N_14108);
and U14259 (N_14259,N_14052,N_14026);
nand U14260 (N_14260,N_14047,N_14123);
xor U14261 (N_14261,N_14159,N_14081);
and U14262 (N_14262,N_14172,N_14017);
nor U14263 (N_14263,N_14188,N_14128);
nand U14264 (N_14264,N_14092,N_14043);
xor U14265 (N_14265,N_14126,N_14007);
nor U14266 (N_14266,N_14147,N_14114);
or U14267 (N_14267,N_14077,N_14046);
or U14268 (N_14268,N_14054,N_14132);
xnor U14269 (N_14269,N_14136,N_14103);
nor U14270 (N_14270,N_14127,N_14105);
nor U14271 (N_14271,N_14032,N_14072);
xnor U14272 (N_14272,N_14169,N_14115);
xnor U14273 (N_14273,N_14042,N_14030);
xnor U14274 (N_14274,N_14000,N_14177);
nand U14275 (N_14275,N_14048,N_14095);
nor U14276 (N_14276,N_14170,N_14085);
xnor U14277 (N_14277,N_14174,N_14141);
nor U14278 (N_14278,N_14171,N_14142);
and U14279 (N_14279,N_14119,N_14178);
xnor U14280 (N_14280,N_14189,N_14190);
or U14281 (N_14281,N_14019,N_14076);
or U14282 (N_14282,N_14061,N_14008);
nor U14283 (N_14283,N_14053,N_14056);
or U14284 (N_14284,N_14097,N_14010);
xor U14285 (N_14285,N_14062,N_14194);
or U14286 (N_14286,N_14151,N_14198);
and U14287 (N_14287,N_14018,N_14104);
xor U14288 (N_14288,N_14100,N_14084);
and U14289 (N_14289,N_14181,N_14145);
xor U14290 (N_14290,N_14144,N_14044);
and U14291 (N_14291,N_14197,N_14075);
or U14292 (N_14292,N_14058,N_14163);
xor U14293 (N_14293,N_14066,N_14130);
and U14294 (N_14294,N_14071,N_14091);
xor U14295 (N_14295,N_14146,N_14087);
and U14296 (N_14296,N_14153,N_14118);
nand U14297 (N_14297,N_14060,N_14029);
nor U14298 (N_14298,N_14149,N_14094);
xnor U14299 (N_14299,N_14036,N_14038);
xnor U14300 (N_14300,N_14157,N_14193);
xnor U14301 (N_14301,N_14060,N_14065);
xnor U14302 (N_14302,N_14071,N_14161);
and U14303 (N_14303,N_14109,N_14056);
xnor U14304 (N_14304,N_14100,N_14167);
nor U14305 (N_14305,N_14052,N_14011);
nand U14306 (N_14306,N_14199,N_14046);
xnor U14307 (N_14307,N_14081,N_14130);
and U14308 (N_14308,N_14028,N_14048);
or U14309 (N_14309,N_14151,N_14178);
or U14310 (N_14310,N_14198,N_14059);
nor U14311 (N_14311,N_14007,N_14045);
nor U14312 (N_14312,N_14104,N_14197);
or U14313 (N_14313,N_14144,N_14101);
or U14314 (N_14314,N_14052,N_14162);
and U14315 (N_14315,N_14018,N_14132);
or U14316 (N_14316,N_14012,N_14060);
or U14317 (N_14317,N_14101,N_14183);
nor U14318 (N_14318,N_14120,N_14057);
nand U14319 (N_14319,N_14025,N_14045);
xnor U14320 (N_14320,N_14085,N_14098);
nor U14321 (N_14321,N_14160,N_14007);
xnor U14322 (N_14322,N_14162,N_14199);
and U14323 (N_14323,N_14177,N_14087);
xnor U14324 (N_14324,N_14103,N_14185);
and U14325 (N_14325,N_14177,N_14007);
xor U14326 (N_14326,N_14189,N_14061);
nor U14327 (N_14327,N_14165,N_14174);
nand U14328 (N_14328,N_14076,N_14080);
and U14329 (N_14329,N_14046,N_14083);
nor U14330 (N_14330,N_14069,N_14093);
and U14331 (N_14331,N_14111,N_14195);
and U14332 (N_14332,N_14095,N_14039);
or U14333 (N_14333,N_14107,N_14167);
nor U14334 (N_14334,N_14013,N_14065);
nor U14335 (N_14335,N_14156,N_14071);
and U14336 (N_14336,N_14051,N_14140);
and U14337 (N_14337,N_14006,N_14045);
or U14338 (N_14338,N_14165,N_14084);
and U14339 (N_14339,N_14180,N_14053);
nor U14340 (N_14340,N_14192,N_14152);
and U14341 (N_14341,N_14167,N_14115);
nand U14342 (N_14342,N_14190,N_14135);
or U14343 (N_14343,N_14101,N_14057);
and U14344 (N_14344,N_14145,N_14045);
xor U14345 (N_14345,N_14140,N_14040);
nor U14346 (N_14346,N_14044,N_14051);
and U14347 (N_14347,N_14045,N_14083);
and U14348 (N_14348,N_14061,N_14127);
xnor U14349 (N_14349,N_14199,N_14070);
and U14350 (N_14350,N_14177,N_14160);
xor U14351 (N_14351,N_14098,N_14080);
and U14352 (N_14352,N_14089,N_14070);
nand U14353 (N_14353,N_14023,N_14145);
and U14354 (N_14354,N_14096,N_14000);
nor U14355 (N_14355,N_14173,N_14163);
nand U14356 (N_14356,N_14145,N_14186);
and U14357 (N_14357,N_14159,N_14071);
or U14358 (N_14358,N_14170,N_14113);
nor U14359 (N_14359,N_14170,N_14114);
and U14360 (N_14360,N_14198,N_14055);
or U14361 (N_14361,N_14161,N_14020);
nand U14362 (N_14362,N_14159,N_14172);
nor U14363 (N_14363,N_14185,N_14147);
xnor U14364 (N_14364,N_14184,N_14006);
or U14365 (N_14365,N_14121,N_14151);
xnor U14366 (N_14366,N_14100,N_14116);
or U14367 (N_14367,N_14034,N_14075);
nor U14368 (N_14368,N_14036,N_14175);
and U14369 (N_14369,N_14133,N_14191);
nor U14370 (N_14370,N_14008,N_14094);
nor U14371 (N_14371,N_14072,N_14199);
or U14372 (N_14372,N_14161,N_14117);
xnor U14373 (N_14373,N_14061,N_14116);
nor U14374 (N_14374,N_14025,N_14048);
nand U14375 (N_14375,N_14009,N_14060);
xor U14376 (N_14376,N_14052,N_14184);
nor U14377 (N_14377,N_14173,N_14159);
and U14378 (N_14378,N_14036,N_14137);
and U14379 (N_14379,N_14002,N_14106);
and U14380 (N_14380,N_14146,N_14134);
xnor U14381 (N_14381,N_14044,N_14188);
nor U14382 (N_14382,N_14008,N_14099);
nand U14383 (N_14383,N_14188,N_14066);
nor U14384 (N_14384,N_14070,N_14073);
xnor U14385 (N_14385,N_14070,N_14014);
xnor U14386 (N_14386,N_14154,N_14073);
xnor U14387 (N_14387,N_14199,N_14035);
nor U14388 (N_14388,N_14092,N_14171);
nor U14389 (N_14389,N_14136,N_14124);
and U14390 (N_14390,N_14074,N_14092);
nand U14391 (N_14391,N_14021,N_14078);
nand U14392 (N_14392,N_14090,N_14052);
nor U14393 (N_14393,N_14177,N_14156);
and U14394 (N_14394,N_14008,N_14100);
nor U14395 (N_14395,N_14170,N_14165);
and U14396 (N_14396,N_14072,N_14166);
nor U14397 (N_14397,N_14199,N_14071);
nand U14398 (N_14398,N_14063,N_14101);
nor U14399 (N_14399,N_14180,N_14043);
and U14400 (N_14400,N_14315,N_14364);
nor U14401 (N_14401,N_14300,N_14309);
nand U14402 (N_14402,N_14322,N_14225);
and U14403 (N_14403,N_14356,N_14308);
nand U14404 (N_14404,N_14237,N_14351);
xnor U14405 (N_14405,N_14216,N_14330);
or U14406 (N_14406,N_14360,N_14213);
nor U14407 (N_14407,N_14376,N_14281);
or U14408 (N_14408,N_14236,N_14388);
nor U14409 (N_14409,N_14202,N_14374);
or U14410 (N_14410,N_14289,N_14269);
xor U14411 (N_14411,N_14250,N_14241);
nor U14412 (N_14412,N_14266,N_14215);
and U14413 (N_14413,N_14224,N_14354);
nor U14414 (N_14414,N_14341,N_14207);
and U14415 (N_14415,N_14307,N_14329);
nor U14416 (N_14416,N_14384,N_14353);
and U14417 (N_14417,N_14346,N_14321);
xor U14418 (N_14418,N_14357,N_14347);
xor U14419 (N_14419,N_14378,N_14242);
or U14420 (N_14420,N_14243,N_14331);
xnor U14421 (N_14421,N_14333,N_14375);
xnor U14422 (N_14422,N_14369,N_14277);
and U14423 (N_14423,N_14324,N_14220);
and U14424 (N_14424,N_14317,N_14370);
nand U14425 (N_14425,N_14340,N_14328);
nor U14426 (N_14426,N_14395,N_14203);
nor U14427 (N_14427,N_14211,N_14306);
or U14428 (N_14428,N_14390,N_14230);
and U14429 (N_14429,N_14342,N_14276);
or U14430 (N_14430,N_14280,N_14293);
or U14431 (N_14431,N_14337,N_14397);
nand U14432 (N_14432,N_14231,N_14362);
nand U14433 (N_14433,N_14234,N_14367);
nor U14434 (N_14434,N_14258,N_14286);
nand U14435 (N_14435,N_14217,N_14380);
xnor U14436 (N_14436,N_14348,N_14343);
and U14437 (N_14437,N_14361,N_14267);
nor U14438 (N_14438,N_14325,N_14392);
or U14439 (N_14439,N_14326,N_14232);
nor U14440 (N_14440,N_14229,N_14257);
nand U14441 (N_14441,N_14262,N_14264);
nand U14442 (N_14442,N_14246,N_14248);
nand U14443 (N_14443,N_14240,N_14278);
xnor U14444 (N_14444,N_14298,N_14201);
or U14445 (N_14445,N_14205,N_14373);
nor U14446 (N_14446,N_14285,N_14338);
nor U14447 (N_14447,N_14222,N_14239);
and U14448 (N_14448,N_14358,N_14323);
and U14449 (N_14449,N_14314,N_14394);
or U14450 (N_14450,N_14295,N_14252);
xnor U14451 (N_14451,N_14393,N_14382);
xor U14452 (N_14452,N_14320,N_14304);
nor U14453 (N_14453,N_14235,N_14312);
or U14454 (N_14454,N_14208,N_14218);
and U14455 (N_14455,N_14279,N_14303);
nand U14456 (N_14456,N_14270,N_14251);
or U14457 (N_14457,N_14292,N_14254);
and U14458 (N_14458,N_14399,N_14272);
or U14459 (N_14459,N_14214,N_14332);
xor U14460 (N_14460,N_14396,N_14352);
or U14461 (N_14461,N_14227,N_14386);
or U14462 (N_14462,N_14368,N_14260);
xor U14463 (N_14463,N_14311,N_14391);
nand U14464 (N_14464,N_14296,N_14389);
nand U14465 (N_14465,N_14398,N_14297);
xnor U14466 (N_14466,N_14290,N_14349);
xnor U14467 (N_14467,N_14233,N_14355);
or U14468 (N_14468,N_14263,N_14316);
and U14469 (N_14469,N_14228,N_14274);
nor U14470 (N_14470,N_14345,N_14282);
and U14471 (N_14471,N_14283,N_14249);
and U14472 (N_14472,N_14383,N_14245);
nand U14473 (N_14473,N_14359,N_14256);
and U14474 (N_14474,N_14291,N_14265);
and U14475 (N_14475,N_14336,N_14288);
nor U14476 (N_14476,N_14261,N_14363);
or U14477 (N_14477,N_14226,N_14223);
or U14478 (N_14478,N_14255,N_14287);
nor U14479 (N_14479,N_14302,N_14221);
or U14480 (N_14480,N_14271,N_14313);
or U14481 (N_14481,N_14381,N_14247);
xnor U14482 (N_14482,N_14305,N_14204);
nand U14483 (N_14483,N_14200,N_14385);
or U14484 (N_14484,N_14371,N_14327);
and U14485 (N_14485,N_14318,N_14377);
or U14486 (N_14486,N_14334,N_14379);
and U14487 (N_14487,N_14210,N_14350);
nand U14488 (N_14488,N_14335,N_14275);
xnor U14489 (N_14489,N_14339,N_14372);
nor U14490 (N_14490,N_14212,N_14284);
xor U14491 (N_14491,N_14299,N_14209);
or U14492 (N_14492,N_14301,N_14294);
xor U14493 (N_14493,N_14259,N_14319);
nor U14494 (N_14494,N_14310,N_14344);
xor U14495 (N_14495,N_14253,N_14206);
nand U14496 (N_14496,N_14273,N_14268);
and U14497 (N_14497,N_14366,N_14244);
and U14498 (N_14498,N_14238,N_14219);
and U14499 (N_14499,N_14387,N_14365);
xor U14500 (N_14500,N_14287,N_14278);
or U14501 (N_14501,N_14204,N_14317);
xnor U14502 (N_14502,N_14374,N_14346);
nor U14503 (N_14503,N_14307,N_14230);
or U14504 (N_14504,N_14379,N_14310);
xnor U14505 (N_14505,N_14222,N_14250);
or U14506 (N_14506,N_14218,N_14324);
or U14507 (N_14507,N_14240,N_14279);
or U14508 (N_14508,N_14336,N_14281);
nor U14509 (N_14509,N_14383,N_14343);
and U14510 (N_14510,N_14274,N_14250);
nor U14511 (N_14511,N_14386,N_14286);
xnor U14512 (N_14512,N_14366,N_14205);
nor U14513 (N_14513,N_14224,N_14212);
xor U14514 (N_14514,N_14245,N_14201);
or U14515 (N_14515,N_14369,N_14387);
and U14516 (N_14516,N_14386,N_14202);
nor U14517 (N_14517,N_14375,N_14210);
xnor U14518 (N_14518,N_14365,N_14361);
and U14519 (N_14519,N_14364,N_14211);
or U14520 (N_14520,N_14336,N_14267);
xor U14521 (N_14521,N_14283,N_14369);
nor U14522 (N_14522,N_14384,N_14206);
nor U14523 (N_14523,N_14343,N_14321);
or U14524 (N_14524,N_14382,N_14343);
or U14525 (N_14525,N_14215,N_14222);
or U14526 (N_14526,N_14326,N_14390);
nor U14527 (N_14527,N_14221,N_14365);
xnor U14528 (N_14528,N_14314,N_14218);
nand U14529 (N_14529,N_14239,N_14365);
xnor U14530 (N_14530,N_14384,N_14236);
nand U14531 (N_14531,N_14268,N_14349);
nor U14532 (N_14532,N_14270,N_14205);
nand U14533 (N_14533,N_14363,N_14263);
or U14534 (N_14534,N_14259,N_14348);
xor U14535 (N_14535,N_14339,N_14293);
nor U14536 (N_14536,N_14290,N_14253);
and U14537 (N_14537,N_14377,N_14211);
nand U14538 (N_14538,N_14349,N_14396);
nand U14539 (N_14539,N_14348,N_14335);
nand U14540 (N_14540,N_14297,N_14345);
xor U14541 (N_14541,N_14285,N_14357);
or U14542 (N_14542,N_14240,N_14397);
nor U14543 (N_14543,N_14298,N_14360);
xor U14544 (N_14544,N_14289,N_14367);
xnor U14545 (N_14545,N_14328,N_14370);
xor U14546 (N_14546,N_14214,N_14317);
and U14547 (N_14547,N_14388,N_14316);
nor U14548 (N_14548,N_14276,N_14374);
or U14549 (N_14549,N_14317,N_14367);
nand U14550 (N_14550,N_14247,N_14204);
nand U14551 (N_14551,N_14256,N_14244);
nand U14552 (N_14552,N_14351,N_14315);
xnor U14553 (N_14553,N_14230,N_14260);
or U14554 (N_14554,N_14240,N_14319);
nand U14555 (N_14555,N_14313,N_14230);
and U14556 (N_14556,N_14362,N_14359);
nor U14557 (N_14557,N_14352,N_14202);
nor U14558 (N_14558,N_14386,N_14347);
nand U14559 (N_14559,N_14393,N_14392);
nand U14560 (N_14560,N_14292,N_14303);
nor U14561 (N_14561,N_14345,N_14313);
and U14562 (N_14562,N_14242,N_14396);
or U14563 (N_14563,N_14325,N_14377);
xor U14564 (N_14564,N_14321,N_14212);
nand U14565 (N_14565,N_14300,N_14259);
or U14566 (N_14566,N_14382,N_14252);
xor U14567 (N_14567,N_14226,N_14222);
nand U14568 (N_14568,N_14374,N_14213);
xor U14569 (N_14569,N_14235,N_14333);
or U14570 (N_14570,N_14338,N_14351);
nand U14571 (N_14571,N_14312,N_14386);
and U14572 (N_14572,N_14329,N_14281);
or U14573 (N_14573,N_14323,N_14350);
nor U14574 (N_14574,N_14310,N_14285);
or U14575 (N_14575,N_14295,N_14325);
nand U14576 (N_14576,N_14376,N_14301);
xor U14577 (N_14577,N_14266,N_14397);
and U14578 (N_14578,N_14272,N_14225);
and U14579 (N_14579,N_14327,N_14302);
or U14580 (N_14580,N_14267,N_14375);
nor U14581 (N_14581,N_14333,N_14299);
xnor U14582 (N_14582,N_14247,N_14289);
xor U14583 (N_14583,N_14264,N_14232);
nor U14584 (N_14584,N_14264,N_14399);
nand U14585 (N_14585,N_14311,N_14229);
and U14586 (N_14586,N_14258,N_14206);
nand U14587 (N_14587,N_14302,N_14332);
and U14588 (N_14588,N_14385,N_14214);
or U14589 (N_14589,N_14215,N_14216);
and U14590 (N_14590,N_14223,N_14387);
nand U14591 (N_14591,N_14266,N_14279);
or U14592 (N_14592,N_14324,N_14211);
nand U14593 (N_14593,N_14368,N_14342);
or U14594 (N_14594,N_14244,N_14296);
xnor U14595 (N_14595,N_14375,N_14391);
or U14596 (N_14596,N_14258,N_14342);
and U14597 (N_14597,N_14255,N_14317);
nor U14598 (N_14598,N_14257,N_14264);
and U14599 (N_14599,N_14369,N_14219);
and U14600 (N_14600,N_14529,N_14456);
xor U14601 (N_14601,N_14564,N_14496);
or U14602 (N_14602,N_14462,N_14511);
nor U14603 (N_14603,N_14576,N_14474);
and U14604 (N_14604,N_14436,N_14485);
nand U14605 (N_14605,N_14441,N_14579);
or U14606 (N_14606,N_14446,N_14415);
nand U14607 (N_14607,N_14443,N_14578);
and U14608 (N_14608,N_14480,N_14521);
nor U14609 (N_14609,N_14453,N_14586);
xor U14610 (N_14610,N_14585,N_14504);
and U14611 (N_14611,N_14520,N_14533);
nand U14612 (N_14612,N_14598,N_14503);
nor U14613 (N_14613,N_14522,N_14413);
or U14614 (N_14614,N_14572,N_14492);
nand U14615 (N_14615,N_14464,N_14475);
nand U14616 (N_14616,N_14563,N_14527);
xor U14617 (N_14617,N_14556,N_14541);
or U14618 (N_14618,N_14425,N_14554);
or U14619 (N_14619,N_14483,N_14481);
nor U14620 (N_14620,N_14531,N_14455);
and U14621 (N_14621,N_14591,N_14429);
nand U14622 (N_14622,N_14407,N_14452);
nand U14623 (N_14623,N_14549,N_14538);
nand U14624 (N_14624,N_14400,N_14547);
nor U14625 (N_14625,N_14442,N_14479);
or U14626 (N_14626,N_14587,N_14500);
or U14627 (N_14627,N_14592,N_14508);
or U14628 (N_14628,N_14582,N_14553);
xor U14629 (N_14629,N_14583,N_14566);
xnor U14630 (N_14630,N_14548,N_14427);
and U14631 (N_14631,N_14417,N_14408);
nand U14632 (N_14632,N_14515,N_14433);
nor U14633 (N_14633,N_14416,N_14546);
and U14634 (N_14634,N_14575,N_14532);
nand U14635 (N_14635,N_14469,N_14580);
and U14636 (N_14636,N_14482,N_14505);
or U14637 (N_14637,N_14457,N_14570);
or U14638 (N_14638,N_14422,N_14523);
xnor U14639 (N_14639,N_14439,N_14435);
xnor U14640 (N_14640,N_14471,N_14526);
nor U14641 (N_14641,N_14489,N_14516);
and U14642 (N_14642,N_14589,N_14424);
nor U14643 (N_14643,N_14560,N_14594);
and U14644 (N_14644,N_14445,N_14565);
and U14645 (N_14645,N_14537,N_14423);
or U14646 (N_14646,N_14571,N_14402);
nor U14647 (N_14647,N_14599,N_14409);
or U14648 (N_14648,N_14498,N_14567);
nand U14649 (N_14649,N_14406,N_14448);
nor U14650 (N_14650,N_14460,N_14535);
nor U14651 (N_14651,N_14545,N_14596);
or U14652 (N_14652,N_14552,N_14488);
xnor U14653 (N_14653,N_14540,N_14414);
xor U14654 (N_14654,N_14447,N_14420);
or U14655 (N_14655,N_14590,N_14404);
nand U14656 (N_14656,N_14426,N_14536);
xnor U14657 (N_14657,N_14430,N_14454);
or U14658 (N_14658,N_14486,N_14517);
and U14659 (N_14659,N_14450,N_14559);
or U14660 (N_14660,N_14476,N_14419);
nor U14661 (N_14661,N_14530,N_14444);
xor U14662 (N_14662,N_14493,N_14451);
nand U14663 (N_14663,N_14544,N_14405);
xnor U14664 (N_14664,N_14461,N_14421);
nor U14665 (N_14665,N_14459,N_14495);
xor U14666 (N_14666,N_14558,N_14513);
xnor U14667 (N_14667,N_14525,N_14431);
or U14668 (N_14668,N_14524,N_14501);
and U14669 (N_14669,N_14449,N_14597);
nor U14670 (N_14670,N_14411,N_14550);
and U14671 (N_14671,N_14588,N_14438);
and U14672 (N_14672,N_14519,N_14502);
xor U14673 (N_14673,N_14418,N_14428);
nor U14674 (N_14674,N_14568,N_14403);
and U14675 (N_14675,N_14542,N_14487);
and U14676 (N_14676,N_14466,N_14410);
and U14677 (N_14677,N_14593,N_14539);
nor U14678 (N_14678,N_14412,N_14490);
nand U14679 (N_14679,N_14465,N_14509);
and U14680 (N_14680,N_14432,N_14584);
xnor U14681 (N_14681,N_14468,N_14561);
xor U14682 (N_14682,N_14595,N_14573);
nor U14683 (N_14683,N_14497,N_14534);
xnor U14684 (N_14684,N_14551,N_14514);
xor U14685 (N_14685,N_14477,N_14574);
xor U14686 (N_14686,N_14478,N_14499);
xnor U14687 (N_14687,N_14562,N_14555);
xor U14688 (N_14688,N_14557,N_14440);
nand U14689 (N_14689,N_14491,N_14458);
nor U14690 (N_14690,N_14512,N_14434);
nand U14691 (N_14691,N_14528,N_14473);
or U14692 (N_14692,N_14463,N_14543);
nor U14693 (N_14693,N_14401,N_14569);
xor U14694 (N_14694,N_14510,N_14507);
nor U14695 (N_14695,N_14577,N_14470);
nand U14696 (N_14696,N_14494,N_14518);
and U14697 (N_14697,N_14472,N_14437);
nor U14698 (N_14698,N_14467,N_14506);
or U14699 (N_14699,N_14581,N_14484);
and U14700 (N_14700,N_14490,N_14525);
nor U14701 (N_14701,N_14584,N_14492);
nand U14702 (N_14702,N_14522,N_14478);
xor U14703 (N_14703,N_14504,N_14502);
xnor U14704 (N_14704,N_14591,N_14499);
xor U14705 (N_14705,N_14407,N_14513);
or U14706 (N_14706,N_14543,N_14478);
and U14707 (N_14707,N_14543,N_14512);
or U14708 (N_14708,N_14517,N_14465);
nand U14709 (N_14709,N_14460,N_14580);
and U14710 (N_14710,N_14567,N_14587);
nor U14711 (N_14711,N_14411,N_14598);
and U14712 (N_14712,N_14499,N_14567);
xnor U14713 (N_14713,N_14554,N_14497);
nand U14714 (N_14714,N_14419,N_14552);
xnor U14715 (N_14715,N_14479,N_14539);
nand U14716 (N_14716,N_14502,N_14493);
xnor U14717 (N_14717,N_14502,N_14479);
and U14718 (N_14718,N_14581,N_14439);
and U14719 (N_14719,N_14586,N_14432);
nand U14720 (N_14720,N_14441,N_14596);
xor U14721 (N_14721,N_14484,N_14554);
xnor U14722 (N_14722,N_14504,N_14596);
or U14723 (N_14723,N_14546,N_14460);
nor U14724 (N_14724,N_14441,N_14515);
nand U14725 (N_14725,N_14414,N_14587);
and U14726 (N_14726,N_14459,N_14536);
and U14727 (N_14727,N_14471,N_14527);
or U14728 (N_14728,N_14483,N_14460);
or U14729 (N_14729,N_14416,N_14585);
and U14730 (N_14730,N_14540,N_14458);
nand U14731 (N_14731,N_14584,N_14547);
nand U14732 (N_14732,N_14503,N_14455);
xor U14733 (N_14733,N_14493,N_14403);
nand U14734 (N_14734,N_14430,N_14511);
and U14735 (N_14735,N_14427,N_14444);
and U14736 (N_14736,N_14571,N_14532);
and U14737 (N_14737,N_14509,N_14442);
xor U14738 (N_14738,N_14585,N_14580);
and U14739 (N_14739,N_14510,N_14458);
or U14740 (N_14740,N_14483,N_14417);
xnor U14741 (N_14741,N_14512,N_14410);
nand U14742 (N_14742,N_14495,N_14430);
xnor U14743 (N_14743,N_14527,N_14554);
nor U14744 (N_14744,N_14493,N_14439);
or U14745 (N_14745,N_14445,N_14532);
nor U14746 (N_14746,N_14571,N_14425);
nor U14747 (N_14747,N_14452,N_14403);
xor U14748 (N_14748,N_14480,N_14445);
and U14749 (N_14749,N_14486,N_14525);
and U14750 (N_14750,N_14578,N_14558);
and U14751 (N_14751,N_14588,N_14492);
nand U14752 (N_14752,N_14476,N_14576);
nor U14753 (N_14753,N_14590,N_14468);
and U14754 (N_14754,N_14425,N_14433);
nor U14755 (N_14755,N_14445,N_14568);
nor U14756 (N_14756,N_14571,N_14477);
nand U14757 (N_14757,N_14520,N_14446);
xor U14758 (N_14758,N_14506,N_14495);
nand U14759 (N_14759,N_14529,N_14448);
xor U14760 (N_14760,N_14464,N_14521);
nand U14761 (N_14761,N_14518,N_14501);
or U14762 (N_14762,N_14429,N_14521);
xnor U14763 (N_14763,N_14526,N_14496);
and U14764 (N_14764,N_14474,N_14561);
nor U14765 (N_14765,N_14504,N_14430);
or U14766 (N_14766,N_14570,N_14556);
and U14767 (N_14767,N_14432,N_14509);
xor U14768 (N_14768,N_14507,N_14531);
and U14769 (N_14769,N_14572,N_14557);
nor U14770 (N_14770,N_14479,N_14453);
xnor U14771 (N_14771,N_14564,N_14431);
nand U14772 (N_14772,N_14536,N_14462);
or U14773 (N_14773,N_14566,N_14559);
xor U14774 (N_14774,N_14581,N_14448);
or U14775 (N_14775,N_14502,N_14420);
and U14776 (N_14776,N_14436,N_14557);
nor U14777 (N_14777,N_14582,N_14530);
nand U14778 (N_14778,N_14435,N_14535);
or U14779 (N_14779,N_14502,N_14500);
and U14780 (N_14780,N_14438,N_14552);
or U14781 (N_14781,N_14582,N_14575);
nand U14782 (N_14782,N_14448,N_14468);
and U14783 (N_14783,N_14500,N_14526);
nor U14784 (N_14784,N_14563,N_14403);
nand U14785 (N_14785,N_14436,N_14498);
and U14786 (N_14786,N_14510,N_14433);
nor U14787 (N_14787,N_14487,N_14520);
xor U14788 (N_14788,N_14588,N_14400);
nand U14789 (N_14789,N_14504,N_14414);
nor U14790 (N_14790,N_14486,N_14573);
and U14791 (N_14791,N_14573,N_14574);
xnor U14792 (N_14792,N_14538,N_14544);
nand U14793 (N_14793,N_14536,N_14532);
nor U14794 (N_14794,N_14483,N_14594);
and U14795 (N_14795,N_14597,N_14470);
nand U14796 (N_14796,N_14553,N_14483);
and U14797 (N_14797,N_14528,N_14401);
xor U14798 (N_14798,N_14464,N_14476);
nand U14799 (N_14799,N_14531,N_14465);
or U14800 (N_14800,N_14799,N_14751);
nor U14801 (N_14801,N_14794,N_14640);
xor U14802 (N_14802,N_14612,N_14710);
xor U14803 (N_14803,N_14724,N_14634);
xor U14804 (N_14804,N_14742,N_14678);
nand U14805 (N_14805,N_14778,N_14711);
xor U14806 (N_14806,N_14667,N_14691);
nand U14807 (N_14807,N_14623,N_14665);
xnor U14808 (N_14808,N_14684,N_14779);
nand U14809 (N_14809,N_14690,N_14693);
nor U14810 (N_14810,N_14686,N_14628);
or U14811 (N_14811,N_14732,N_14659);
and U14812 (N_14812,N_14645,N_14703);
nor U14813 (N_14813,N_14635,N_14602);
nor U14814 (N_14814,N_14715,N_14739);
xor U14815 (N_14815,N_14696,N_14780);
nor U14816 (N_14816,N_14603,N_14611);
xnor U14817 (N_14817,N_14615,N_14601);
and U14818 (N_14818,N_14661,N_14781);
and U14819 (N_14819,N_14642,N_14728);
nor U14820 (N_14820,N_14735,N_14760);
and U14821 (N_14821,N_14750,N_14796);
and U14822 (N_14822,N_14713,N_14643);
nand U14823 (N_14823,N_14670,N_14788);
or U14824 (N_14824,N_14625,N_14725);
xnor U14825 (N_14825,N_14764,N_14669);
nand U14826 (N_14826,N_14707,N_14610);
or U14827 (N_14827,N_14649,N_14626);
or U14828 (N_14828,N_14644,N_14700);
xnor U14829 (N_14829,N_14738,N_14662);
nor U14830 (N_14830,N_14631,N_14740);
and U14831 (N_14831,N_14632,N_14789);
or U14832 (N_14832,N_14749,N_14687);
nand U14833 (N_14833,N_14666,N_14655);
nand U14834 (N_14834,N_14747,N_14638);
and U14835 (N_14835,N_14766,N_14716);
and U14836 (N_14836,N_14608,N_14718);
or U14837 (N_14837,N_14671,N_14775);
and U14838 (N_14838,N_14694,N_14726);
nand U14839 (N_14839,N_14748,N_14768);
and U14840 (N_14840,N_14736,N_14784);
nor U14841 (N_14841,N_14737,N_14629);
or U14842 (N_14842,N_14759,N_14656);
nor U14843 (N_14843,N_14787,N_14609);
nand U14844 (N_14844,N_14795,N_14639);
xnor U14845 (N_14845,N_14674,N_14754);
nor U14846 (N_14846,N_14654,N_14746);
nand U14847 (N_14847,N_14723,N_14791);
and U14848 (N_14848,N_14614,N_14769);
and U14849 (N_14849,N_14752,N_14774);
nor U14850 (N_14850,N_14708,N_14743);
and U14851 (N_14851,N_14681,N_14650);
and U14852 (N_14852,N_14660,N_14653);
and U14853 (N_14853,N_14731,N_14651);
nor U14854 (N_14854,N_14677,N_14619);
nor U14855 (N_14855,N_14744,N_14706);
xor U14856 (N_14856,N_14604,N_14721);
or U14857 (N_14857,N_14673,N_14636);
and U14858 (N_14858,N_14633,N_14792);
or U14859 (N_14859,N_14757,N_14782);
nor U14860 (N_14860,N_14600,N_14717);
xor U14861 (N_14861,N_14730,N_14705);
and U14862 (N_14862,N_14648,N_14652);
nor U14863 (N_14863,N_14712,N_14704);
nor U14864 (N_14864,N_14701,N_14770);
or U14865 (N_14865,N_14745,N_14605);
nor U14866 (N_14866,N_14679,N_14698);
nor U14867 (N_14867,N_14692,N_14699);
nor U14868 (N_14868,N_14767,N_14756);
nor U14869 (N_14869,N_14630,N_14772);
and U14870 (N_14870,N_14727,N_14785);
xnor U14871 (N_14871,N_14607,N_14761);
xor U14872 (N_14872,N_14624,N_14771);
and U14873 (N_14873,N_14627,N_14797);
xor U14874 (N_14874,N_14790,N_14672);
or U14875 (N_14875,N_14641,N_14657);
xnor U14876 (N_14876,N_14719,N_14663);
or U14877 (N_14877,N_14777,N_14668);
nor U14878 (N_14878,N_14755,N_14675);
nand U14879 (N_14879,N_14613,N_14664);
or U14880 (N_14880,N_14682,N_14773);
and U14881 (N_14881,N_14729,N_14617);
and U14882 (N_14882,N_14702,N_14753);
and U14883 (N_14883,N_14714,N_14763);
nor U14884 (N_14884,N_14637,N_14722);
nand U14885 (N_14885,N_14606,N_14733);
xor U14886 (N_14886,N_14646,N_14658);
nand U14887 (N_14887,N_14762,N_14783);
nor U14888 (N_14888,N_14616,N_14697);
nor U14889 (N_14889,N_14798,N_14621);
xnor U14890 (N_14890,N_14688,N_14741);
nor U14891 (N_14891,N_14720,N_14689);
xnor U14892 (N_14892,N_14765,N_14622);
nor U14893 (N_14893,N_14793,N_14695);
nand U14894 (N_14894,N_14776,N_14620);
xnor U14895 (N_14895,N_14676,N_14685);
xor U14896 (N_14896,N_14680,N_14786);
xor U14897 (N_14897,N_14647,N_14683);
nor U14898 (N_14898,N_14618,N_14758);
xnor U14899 (N_14899,N_14734,N_14709);
and U14900 (N_14900,N_14708,N_14790);
xor U14901 (N_14901,N_14658,N_14749);
and U14902 (N_14902,N_14753,N_14698);
and U14903 (N_14903,N_14640,N_14651);
nand U14904 (N_14904,N_14728,N_14617);
nor U14905 (N_14905,N_14686,N_14688);
and U14906 (N_14906,N_14682,N_14677);
and U14907 (N_14907,N_14779,N_14644);
nand U14908 (N_14908,N_14731,N_14728);
nor U14909 (N_14909,N_14680,N_14619);
xor U14910 (N_14910,N_14728,N_14768);
nor U14911 (N_14911,N_14667,N_14749);
and U14912 (N_14912,N_14797,N_14723);
xnor U14913 (N_14913,N_14610,N_14687);
nand U14914 (N_14914,N_14691,N_14793);
nor U14915 (N_14915,N_14600,N_14607);
and U14916 (N_14916,N_14768,N_14708);
or U14917 (N_14917,N_14684,N_14767);
xor U14918 (N_14918,N_14634,N_14717);
nand U14919 (N_14919,N_14697,N_14639);
nor U14920 (N_14920,N_14730,N_14759);
nor U14921 (N_14921,N_14687,N_14672);
nor U14922 (N_14922,N_14778,N_14663);
nand U14923 (N_14923,N_14675,N_14649);
xor U14924 (N_14924,N_14781,N_14611);
xor U14925 (N_14925,N_14681,N_14757);
or U14926 (N_14926,N_14603,N_14698);
xnor U14927 (N_14927,N_14717,N_14757);
and U14928 (N_14928,N_14764,N_14787);
nand U14929 (N_14929,N_14646,N_14767);
or U14930 (N_14930,N_14690,N_14725);
xnor U14931 (N_14931,N_14741,N_14740);
or U14932 (N_14932,N_14617,N_14726);
nor U14933 (N_14933,N_14644,N_14623);
or U14934 (N_14934,N_14626,N_14732);
and U14935 (N_14935,N_14782,N_14781);
and U14936 (N_14936,N_14765,N_14758);
nand U14937 (N_14937,N_14722,N_14796);
nand U14938 (N_14938,N_14602,N_14642);
nand U14939 (N_14939,N_14771,N_14710);
or U14940 (N_14940,N_14753,N_14697);
and U14941 (N_14941,N_14728,N_14761);
and U14942 (N_14942,N_14655,N_14609);
xnor U14943 (N_14943,N_14719,N_14743);
and U14944 (N_14944,N_14697,N_14739);
nand U14945 (N_14945,N_14670,N_14601);
or U14946 (N_14946,N_14756,N_14625);
nand U14947 (N_14947,N_14658,N_14694);
nor U14948 (N_14948,N_14782,N_14755);
nand U14949 (N_14949,N_14688,N_14606);
xnor U14950 (N_14950,N_14768,N_14658);
nand U14951 (N_14951,N_14729,N_14697);
nand U14952 (N_14952,N_14724,N_14651);
nor U14953 (N_14953,N_14725,N_14706);
xnor U14954 (N_14954,N_14692,N_14751);
nand U14955 (N_14955,N_14641,N_14782);
nor U14956 (N_14956,N_14712,N_14618);
and U14957 (N_14957,N_14769,N_14720);
or U14958 (N_14958,N_14625,N_14712);
nand U14959 (N_14959,N_14705,N_14653);
xnor U14960 (N_14960,N_14713,N_14667);
xor U14961 (N_14961,N_14602,N_14631);
and U14962 (N_14962,N_14776,N_14615);
nand U14963 (N_14963,N_14760,N_14747);
or U14964 (N_14964,N_14657,N_14764);
nand U14965 (N_14965,N_14639,N_14663);
nor U14966 (N_14966,N_14649,N_14769);
nor U14967 (N_14967,N_14623,N_14764);
or U14968 (N_14968,N_14785,N_14617);
xnor U14969 (N_14969,N_14628,N_14762);
nand U14970 (N_14970,N_14674,N_14775);
or U14971 (N_14971,N_14645,N_14602);
and U14972 (N_14972,N_14675,N_14703);
nor U14973 (N_14973,N_14650,N_14687);
xor U14974 (N_14974,N_14798,N_14724);
or U14975 (N_14975,N_14630,N_14680);
xnor U14976 (N_14976,N_14694,N_14627);
or U14977 (N_14977,N_14796,N_14719);
nor U14978 (N_14978,N_14675,N_14655);
or U14979 (N_14979,N_14743,N_14796);
nand U14980 (N_14980,N_14649,N_14640);
nand U14981 (N_14981,N_14705,N_14689);
nor U14982 (N_14982,N_14628,N_14665);
nor U14983 (N_14983,N_14787,N_14691);
xor U14984 (N_14984,N_14758,N_14728);
nand U14985 (N_14985,N_14663,N_14695);
nor U14986 (N_14986,N_14790,N_14783);
or U14987 (N_14987,N_14702,N_14761);
and U14988 (N_14988,N_14756,N_14673);
nand U14989 (N_14989,N_14787,N_14791);
or U14990 (N_14990,N_14776,N_14642);
or U14991 (N_14991,N_14783,N_14734);
nor U14992 (N_14992,N_14751,N_14601);
nand U14993 (N_14993,N_14686,N_14745);
or U14994 (N_14994,N_14667,N_14777);
or U14995 (N_14995,N_14738,N_14794);
nand U14996 (N_14996,N_14700,N_14721);
or U14997 (N_14997,N_14695,N_14612);
xor U14998 (N_14998,N_14659,N_14711);
nand U14999 (N_14999,N_14699,N_14610);
nor U15000 (N_15000,N_14816,N_14828);
xnor U15001 (N_15001,N_14862,N_14940);
nor U15002 (N_15002,N_14970,N_14952);
or U15003 (N_15003,N_14817,N_14997);
or U15004 (N_15004,N_14872,N_14993);
nand U15005 (N_15005,N_14875,N_14936);
and U15006 (N_15006,N_14827,N_14867);
nand U15007 (N_15007,N_14995,N_14841);
nand U15008 (N_15008,N_14966,N_14825);
nor U15009 (N_15009,N_14985,N_14939);
or U15010 (N_15010,N_14865,N_14990);
xnor U15011 (N_15011,N_14992,N_14961);
xnor U15012 (N_15012,N_14916,N_14886);
and U15013 (N_15013,N_14891,N_14978);
xnor U15014 (N_15014,N_14861,N_14920);
xor U15015 (N_15015,N_14975,N_14803);
xnor U15016 (N_15016,N_14996,N_14955);
nand U15017 (N_15017,N_14931,N_14963);
nor U15018 (N_15018,N_14819,N_14911);
xor U15019 (N_15019,N_14932,N_14994);
or U15020 (N_15020,N_14831,N_14974);
nor U15021 (N_15021,N_14950,N_14833);
xor U15022 (N_15022,N_14938,N_14956);
xor U15023 (N_15023,N_14856,N_14802);
nand U15024 (N_15024,N_14881,N_14925);
xnor U15025 (N_15025,N_14818,N_14953);
xor U15026 (N_15026,N_14937,N_14988);
xor U15027 (N_15027,N_14846,N_14915);
nand U15028 (N_15028,N_14839,N_14922);
xnor U15029 (N_15029,N_14933,N_14903);
xnor U15030 (N_15030,N_14951,N_14830);
nor U15031 (N_15031,N_14873,N_14926);
xnor U15032 (N_15032,N_14840,N_14980);
or U15033 (N_15033,N_14853,N_14929);
xor U15034 (N_15034,N_14912,N_14851);
nand U15035 (N_15035,N_14800,N_14834);
nor U15036 (N_15036,N_14899,N_14913);
and U15037 (N_15037,N_14812,N_14887);
nor U15038 (N_15038,N_14969,N_14957);
and U15039 (N_15039,N_14835,N_14808);
nor U15040 (N_15040,N_14981,N_14845);
and U15041 (N_15041,N_14900,N_14858);
xnor U15042 (N_15042,N_14890,N_14894);
nor U15043 (N_15043,N_14857,N_14815);
or U15044 (N_15044,N_14882,N_14810);
or U15045 (N_15045,N_14965,N_14917);
nand U15046 (N_15046,N_14863,N_14941);
xor U15047 (N_15047,N_14914,N_14968);
or U15048 (N_15048,N_14962,N_14804);
nand U15049 (N_15049,N_14944,N_14870);
nand U15050 (N_15050,N_14885,N_14811);
and U15051 (N_15051,N_14901,N_14945);
xnor U15052 (N_15052,N_14877,N_14964);
nand U15053 (N_15053,N_14924,N_14888);
nand U15054 (N_15054,N_14972,N_14847);
xnor U15055 (N_15055,N_14868,N_14906);
or U15056 (N_15056,N_14871,N_14838);
xnor U15057 (N_15057,N_14942,N_14849);
nand U15058 (N_15058,N_14948,N_14971);
nor U15059 (N_15059,N_14976,N_14860);
and U15060 (N_15060,N_14934,N_14908);
nand U15061 (N_15061,N_14984,N_14904);
or U15062 (N_15062,N_14927,N_14977);
nand U15063 (N_15063,N_14859,N_14866);
nor U15064 (N_15064,N_14943,N_14910);
or U15065 (N_15065,N_14928,N_14854);
nor U15066 (N_15066,N_14883,N_14880);
and U15067 (N_15067,N_14909,N_14844);
nand U15068 (N_15068,N_14892,N_14829);
xor U15069 (N_15069,N_14954,N_14842);
and U15070 (N_15070,N_14991,N_14878);
and U15071 (N_15071,N_14923,N_14823);
or U15072 (N_15072,N_14850,N_14983);
or U15073 (N_15073,N_14999,N_14869);
xor U15074 (N_15074,N_14998,N_14879);
xor U15075 (N_15075,N_14801,N_14832);
xnor U15076 (N_15076,N_14826,N_14813);
xnor U15077 (N_15077,N_14837,N_14960);
or U15078 (N_15078,N_14874,N_14876);
xnor U15079 (N_15079,N_14987,N_14864);
nand U15080 (N_15080,N_14958,N_14986);
or U15081 (N_15081,N_14895,N_14852);
and U15082 (N_15082,N_14949,N_14982);
xnor U15083 (N_15083,N_14855,N_14902);
and U15084 (N_15084,N_14824,N_14820);
or U15085 (N_15085,N_14809,N_14946);
or U15086 (N_15086,N_14989,N_14905);
or U15087 (N_15087,N_14947,N_14889);
or U15088 (N_15088,N_14930,N_14935);
and U15089 (N_15089,N_14843,N_14805);
nor U15090 (N_15090,N_14821,N_14907);
nor U15091 (N_15091,N_14979,N_14893);
or U15092 (N_15092,N_14806,N_14807);
nand U15093 (N_15093,N_14967,N_14814);
nor U15094 (N_15094,N_14973,N_14884);
nand U15095 (N_15095,N_14919,N_14822);
and U15096 (N_15096,N_14896,N_14898);
and U15097 (N_15097,N_14959,N_14836);
or U15098 (N_15098,N_14848,N_14921);
and U15099 (N_15099,N_14897,N_14918);
and U15100 (N_15100,N_14861,N_14843);
nor U15101 (N_15101,N_14888,N_14812);
nand U15102 (N_15102,N_14958,N_14947);
nor U15103 (N_15103,N_14887,N_14801);
and U15104 (N_15104,N_14833,N_14987);
and U15105 (N_15105,N_14887,N_14926);
or U15106 (N_15106,N_14975,N_14925);
nor U15107 (N_15107,N_14854,N_14898);
nand U15108 (N_15108,N_14943,N_14841);
nor U15109 (N_15109,N_14856,N_14939);
nand U15110 (N_15110,N_14904,N_14913);
nor U15111 (N_15111,N_14863,N_14969);
and U15112 (N_15112,N_14800,N_14946);
nand U15113 (N_15113,N_14864,N_14845);
xnor U15114 (N_15114,N_14916,N_14899);
or U15115 (N_15115,N_14825,N_14900);
nor U15116 (N_15116,N_14918,N_14811);
nand U15117 (N_15117,N_14993,N_14972);
and U15118 (N_15118,N_14941,N_14936);
nor U15119 (N_15119,N_14926,N_14964);
and U15120 (N_15120,N_14971,N_14915);
xnor U15121 (N_15121,N_14835,N_14999);
xnor U15122 (N_15122,N_14970,N_14865);
nand U15123 (N_15123,N_14909,N_14908);
and U15124 (N_15124,N_14972,N_14917);
xnor U15125 (N_15125,N_14830,N_14938);
and U15126 (N_15126,N_14890,N_14860);
and U15127 (N_15127,N_14873,N_14812);
or U15128 (N_15128,N_14819,N_14855);
or U15129 (N_15129,N_14893,N_14895);
and U15130 (N_15130,N_14934,N_14883);
nand U15131 (N_15131,N_14874,N_14975);
xnor U15132 (N_15132,N_14831,N_14817);
nor U15133 (N_15133,N_14875,N_14965);
nand U15134 (N_15134,N_14914,N_14850);
xor U15135 (N_15135,N_14960,N_14879);
or U15136 (N_15136,N_14941,N_14803);
nand U15137 (N_15137,N_14817,N_14905);
and U15138 (N_15138,N_14977,N_14831);
and U15139 (N_15139,N_14958,N_14981);
xnor U15140 (N_15140,N_14891,N_14803);
and U15141 (N_15141,N_14902,N_14926);
and U15142 (N_15142,N_14935,N_14806);
xor U15143 (N_15143,N_14974,N_14888);
nor U15144 (N_15144,N_14944,N_14980);
xnor U15145 (N_15145,N_14810,N_14892);
nor U15146 (N_15146,N_14921,N_14912);
nand U15147 (N_15147,N_14972,N_14965);
nand U15148 (N_15148,N_14991,N_14974);
xnor U15149 (N_15149,N_14863,N_14803);
xnor U15150 (N_15150,N_14923,N_14945);
nor U15151 (N_15151,N_14975,N_14905);
xnor U15152 (N_15152,N_14857,N_14943);
and U15153 (N_15153,N_14956,N_14884);
and U15154 (N_15154,N_14951,N_14870);
or U15155 (N_15155,N_14952,N_14901);
nand U15156 (N_15156,N_14899,N_14864);
or U15157 (N_15157,N_14859,N_14984);
nand U15158 (N_15158,N_14914,N_14980);
and U15159 (N_15159,N_14861,N_14973);
nand U15160 (N_15160,N_14979,N_14910);
nand U15161 (N_15161,N_14802,N_14990);
and U15162 (N_15162,N_14864,N_14906);
or U15163 (N_15163,N_14964,N_14958);
nor U15164 (N_15164,N_14860,N_14937);
nand U15165 (N_15165,N_14821,N_14964);
nand U15166 (N_15166,N_14816,N_14848);
nor U15167 (N_15167,N_14873,N_14859);
and U15168 (N_15168,N_14982,N_14846);
nand U15169 (N_15169,N_14805,N_14992);
xnor U15170 (N_15170,N_14858,N_14817);
and U15171 (N_15171,N_14800,N_14964);
nand U15172 (N_15172,N_14807,N_14842);
or U15173 (N_15173,N_14891,N_14845);
nand U15174 (N_15174,N_14802,N_14807);
nand U15175 (N_15175,N_14922,N_14968);
xnor U15176 (N_15176,N_14806,N_14886);
nand U15177 (N_15177,N_14971,N_14945);
or U15178 (N_15178,N_14806,N_14992);
and U15179 (N_15179,N_14813,N_14980);
xor U15180 (N_15180,N_14913,N_14942);
nor U15181 (N_15181,N_14885,N_14914);
nor U15182 (N_15182,N_14930,N_14829);
nor U15183 (N_15183,N_14990,N_14915);
nand U15184 (N_15184,N_14956,N_14992);
and U15185 (N_15185,N_14990,N_14848);
and U15186 (N_15186,N_14882,N_14977);
and U15187 (N_15187,N_14955,N_14879);
xnor U15188 (N_15188,N_14999,N_14849);
nand U15189 (N_15189,N_14966,N_14919);
and U15190 (N_15190,N_14975,N_14985);
xnor U15191 (N_15191,N_14942,N_14969);
nor U15192 (N_15192,N_14998,N_14995);
nand U15193 (N_15193,N_14980,N_14983);
nor U15194 (N_15194,N_14925,N_14852);
or U15195 (N_15195,N_14936,N_14831);
or U15196 (N_15196,N_14878,N_14822);
xor U15197 (N_15197,N_14915,N_14967);
and U15198 (N_15198,N_14833,N_14894);
or U15199 (N_15199,N_14831,N_14924);
xor U15200 (N_15200,N_15030,N_15045);
nor U15201 (N_15201,N_15049,N_15118);
and U15202 (N_15202,N_15007,N_15038);
xor U15203 (N_15203,N_15072,N_15074);
or U15204 (N_15204,N_15155,N_15044);
xnor U15205 (N_15205,N_15008,N_15025);
and U15206 (N_15206,N_15097,N_15145);
nor U15207 (N_15207,N_15116,N_15054);
xnor U15208 (N_15208,N_15157,N_15112);
and U15209 (N_15209,N_15115,N_15184);
and U15210 (N_15210,N_15031,N_15075);
xor U15211 (N_15211,N_15013,N_15056);
nand U15212 (N_15212,N_15053,N_15103);
nor U15213 (N_15213,N_15125,N_15175);
xnor U15214 (N_15214,N_15179,N_15099);
nor U15215 (N_15215,N_15083,N_15046);
or U15216 (N_15216,N_15197,N_15114);
xor U15217 (N_15217,N_15111,N_15003);
nor U15218 (N_15218,N_15084,N_15193);
nand U15219 (N_15219,N_15036,N_15019);
or U15220 (N_15220,N_15077,N_15015);
nand U15221 (N_15221,N_15109,N_15011);
nor U15222 (N_15222,N_15186,N_15004);
or U15223 (N_15223,N_15119,N_15037);
xnor U15224 (N_15224,N_15141,N_15024);
or U15225 (N_15225,N_15107,N_15171);
and U15226 (N_15226,N_15117,N_15068);
nand U15227 (N_15227,N_15100,N_15079);
xor U15228 (N_15228,N_15034,N_15195);
nand U15229 (N_15229,N_15090,N_15060);
nand U15230 (N_15230,N_15105,N_15156);
nand U15231 (N_15231,N_15122,N_15110);
xor U15232 (N_15232,N_15067,N_15163);
xnor U15233 (N_15233,N_15026,N_15069);
nand U15234 (N_15234,N_15050,N_15042);
nor U15235 (N_15235,N_15108,N_15148);
nand U15236 (N_15236,N_15087,N_15198);
xnor U15237 (N_15237,N_15023,N_15086);
nand U15238 (N_15238,N_15048,N_15135);
and U15239 (N_15239,N_15059,N_15160);
nand U15240 (N_15240,N_15181,N_15137);
xor U15241 (N_15241,N_15169,N_15094);
nand U15242 (N_15242,N_15180,N_15168);
and U15243 (N_15243,N_15158,N_15129);
nand U15244 (N_15244,N_15029,N_15088);
and U15245 (N_15245,N_15071,N_15021);
nand U15246 (N_15246,N_15058,N_15190);
or U15247 (N_15247,N_15096,N_15188);
nor U15248 (N_15248,N_15147,N_15126);
nor U15249 (N_15249,N_15081,N_15170);
nor U15250 (N_15250,N_15017,N_15027);
and U15251 (N_15251,N_15093,N_15095);
or U15252 (N_15252,N_15080,N_15066);
and U15253 (N_15253,N_15123,N_15043);
xnor U15254 (N_15254,N_15178,N_15020);
xor U15255 (N_15255,N_15154,N_15151);
xor U15256 (N_15256,N_15033,N_15166);
nor U15257 (N_15257,N_15173,N_15127);
nand U15258 (N_15258,N_15062,N_15032);
nor U15259 (N_15259,N_15085,N_15082);
nor U15260 (N_15260,N_15150,N_15018);
and U15261 (N_15261,N_15187,N_15101);
or U15262 (N_15262,N_15124,N_15136);
and U15263 (N_15263,N_15113,N_15022);
nor U15264 (N_15264,N_15040,N_15153);
nand U15265 (N_15265,N_15005,N_15041);
and U15266 (N_15266,N_15132,N_15051);
nand U15267 (N_15267,N_15006,N_15191);
or U15268 (N_15268,N_15014,N_15089);
nor U15269 (N_15269,N_15120,N_15194);
xor U15270 (N_15270,N_15012,N_15001);
or U15271 (N_15271,N_15138,N_15065);
nor U15272 (N_15272,N_15177,N_15078);
xor U15273 (N_15273,N_15098,N_15131);
nor U15274 (N_15274,N_15172,N_15159);
or U15275 (N_15275,N_15164,N_15121);
xor U15276 (N_15276,N_15162,N_15144);
and U15277 (N_15277,N_15189,N_15035);
nand U15278 (N_15278,N_15047,N_15061);
and U15279 (N_15279,N_15146,N_15152);
or U15280 (N_15280,N_15134,N_15106);
xnor U15281 (N_15281,N_15140,N_15057);
xor U15282 (N_15282,N_15143,N_15174);
nor U15283 (N_15283,N_15133,N_15161);
or U15284 (N_15284,N_15039,N_15064);
nand U15285 (N_15285,N_15076,N_15104);
nor U15286 (N_15286,N_15055,N_15000);
xor U15287 (N_15287,N_15192,N_15182);
nor U15288 (N_15288,N_15183,N_15010);
nand U15289 (N_15289,N_15028,N_15139);
and U15290 (N_15290,N_15070,N_15130);
or U15291 (N_15291,N_15091,N_15016);
and U15292 (N_15292,N_15073,N_15149);
nand U15293 (N_15293,N_15196,N_15052);
or U15294 (N_15294,N_15167,N_15092);
nor U15295 (N_15295,N_15142,N_15002);
xor U15296 (N_15296,N_15063,N_15009);
nor U15297 (N_15297,N_15128,N_15199);
and U15298 (N_15298,N_15102,N_15165);
nand U15299 (N_15299,N_15185,N_15176);
xor U15300 (N_15300,N_15170,N_15137);
nor U15301 (N_15301,N_15080,N_15008);
nor U15302 (N_15302,N_15021,N_15106);
and U15303 (N_15303,N_15116,N_15075);
xor U15304 (N_15304,N_15030,N_15134);
or U15305 (N_15305,N_15060,N_15000);
nand U15306 (N_15306,N_15102,N_15047);
nand U15307 (N_15307,N_15079,N_15171);
xnor U15308 (N_15308,N_15147,N_15015);
nor U15309 (N_15309,N_15139,N_15091);
or U15310 (N_15310,N_15098,N_15037);
or U15311 (N_15311,N_15010,N_15127);
or U15312 (N_15312,N_15126,N_15072);
nor U15313 (N_15313,N_15178,N_15042);
or U15314 (N_15314,N_15052,N_15167);
xnor U15315 (N_15315,N_15031,N_15155);
xnor U15316 (N_15316,N_15053,N_15098);
xnor U15317 (N_15317,N_15185,N_15149);
and U15318 (N_15318,N_15116,N_15108);
and U15319 (N_15319,N_15183,N_15008);
xor U15320 (N_15320,N_15130,N_15110);
nand U15321 (N_15321,N_15040,N_15157);
or U15322 (N_15322,N_15171,N_15162);
xnor U15323 (N_15323,N_15141,N_15121);
xor U15324 (N_15324,N_15177,N_15136);
nand U15325 (N_15325,N_15023,N_15003);
nand U15326 (N_15326,N_15106,N_15179);
nor U15327 (N_15327,N_15068,N_15195);
nand U15328 (N_15328,N_15130,N_15103);
nand U15329 (N_15329,N_15005,N_15092);
and U15330 (N_15330,N_15028,N_15154);
nor U15331 (N_15331,N_15159,N_15166);
or U15332 (N_15332,N_15073,N_15097);
xnor U15333 (N_15333,N_15145,N_15039);
or U15334 (N_15334,N_15158,N_15075);
xnor U15335 (N_15335,N_15028,N_15062);
or U15336 (N_15336,N_15050,N_15106);
and U15337 (N_15337,N_15065,N_15038);
or U15338 (N_15338,N_15079,N_15130);
or U15339 (N_15339,N_15036,N_15089);
and U15340 (N_15340,N_15020,N_15012);
xor U15341 (N_15341,N_15172,N_15094);
nand U15342 (N_15342,N_15097,N_15182);
and U15343 (N_15343,N_15012,N_15099);
xor U15344 (N_15344,N_15157,N_15138);
nand U15345 (N_15345,N_15191,N_15163);
or U15346 (N_15346,N_15019,N_15134);
or U15347 (N_15347,N_15037,N_15160);
and U15348 (N_15348,N_15067,N_15118);
and U15349 (N_15349,N_15121,N_15044);
xnor U15350 (N_15350,N_15075,N_15154);
nor U15351 (N_15351,N_15108,N_15139);
nand U15352 (N_15352,N_15127,N_15140);
xor U15353 (N_15353,N_15012,N_15121);
or U15354 (N_15354,N_15060,N_15003);
and U15355 (N_15355,N_15124,N_15057);
nand U15356 (N_15356,N_15075,N_15065);
nor U15357 (N_15357,N_15154,N_15184);
and U15358 (N_15358,N_15070,N_15081);
and U15359 (N_15359,N_15058,N_15083);
nand U15360 (N_15360,N_15189,N_15172);
or U15361 (N_15361,N_15121,N_15074);
or U15362 (N_15362,N_15079,N_15155);
xnor U15363 (N_15363,N_15130,N_15181);
and U15364 (N_15364,N_15191,N_15107);
and U15365 (N_15365,N_15046,N_15011);
and U15366 (N_15366,N_15030,N_15006);
or U15367 (N_15367,N_15058,N_15156);
or U15368 (N_15368,N_15067,N_15016);
nor U15369 (N_15369,N_15158,N_15079);
or U15370 (N_15370,N_15052,N_15099);
and U15371 (N_15371,N_15181,N_15092);
or U15372 (N_15372,N_15103,N_15005);
xor U15373 (N_15373,N_15175,N_15051);
nand U15374 (N_15374,N_15017,N_15112);
xnor U15375 (N_15375,N_15094,N_15144);
nor U15376 (N_15376,N_15048,N_15133);
xor U15377 (N_15377,N_15129,N_15099);
xnor U15378 (N_15378,N_15197,N_15167);
or U15379 (N_15379,N_15014,N_15069);
or U15380 (N_15380,N_15157,N_15059);
xor U15381 (N_15381,N_15168,N_15012);
nor U15382 (N_15382,N_15180,N_15112);
and U15383 (N_15383,N_15171,N_15010);
xor U15384 (N_15384,N_15139,N_15177);
nand U15385 (N_15385,N_15140,N_15101);
xor U15386 (N_15386,N_15027,N_15078);
nor U15387 (N_15387,N_15038,N_15064);
nand U15388 (N_15388,N_15084,N_15078);
and U15389 (N_15389,N_15110,N_15154);
xnor U15390 (N_15390,N_15025,N_15141);
and U15391 (N_15391,N_15194,N_15007);
nand U15392 (N_15392,N_15159,N_15180);
xor U15393 (N_15393,N_15073,N_15098);
xnor U15394 (N_15394,N_15055,N_15105);
nand U15395 (N_15395,N_15197,N_15140);
nor U15396 (N_15396,N_15018,N_15151);
xnor U15397 (N_15397,N_15003,N_15063);
nand U15398 (N_15398,N_15001,N_15043);
or U15399 (N_15399,N_15153,N_15066);
nand U15400 (N_15400,N_15236,N_15316);
xnor U15401 (N_15401,N_15234,N_15366);
nand U15402 (N_15402,N_15332,N_15306);
xnor U15403 (N_15403,N_15295,N_15380);
or U15404 (N_15404,N_15394,N_15344);
nor U15405 (N_15405,N_15274,N_15279);
and U15406 (N_15406,N_15389,N_15395);
or U15407 (N_15407,N_15314,N_15305);
nor U15408 (N_15408,N_15377,N_15354);
or U15409 (N_15409,N_15388,N_15367);
nor U15410 (N_15410,N_15379,N_15398);
nand U15411 (N_15411,N_15341,N_15286);
and U15412 (N_15412,N_15378,N_15269);
or U15413 (N_15413,N_15368,N_15291);
nor U15414 (N_15414,N_15239,N_15308);
or U15415 (N_15415,N_15261,N_15302);
nor U15416 (N_15416,N_15242,N_15347);
and U15417 (N_15417,N_15205,N_15243);
nor U15418 (N_15418,N_15249,N_15386);
or U15419 (N_15419,N_15376,N_15357);
xor U15420 (N_15420,N_15225,N_15244);
xnor U15421 (N_15421,N_15227,N_15211);
and U15422 (N_15422,N_15229,N_15233);
nor U15423 (N_15423,N_15319,N_15215);
nand U15424 (N_15424,N_15200,N_15251);
or U15425 (N_15425,N_15263,N_15396);
nor U15426 (N_15426,N_15385,N_15355);
and U15427 (N_15427,N_15217,N_15320);
or U15428 (N_15428,N_15277,N_15348);
or U15429 (N_15429,N_15276,N_15324);
nor U15430 (N_15430,N_15289,N_15315);
nor U15431 (N_15431,N_15255,N_15253);
xor U15432 (N_15432,N_15201,N_15349);
nor U15433 (N_15433,N_15299,N_15247);
and U15434 (N_15434,N_15293,N_15387);
xor U15435 (N_15435,N_15262,N_15397);
nor U15436 (N_15436,N_15343,N_15370);
xnor U15437 (N_15437,N_15248,N_15222);
xnor U15438 (N_15438,N_15301,N_15311);
nor U15439 (N_15439,N_15207,N_15384);
nand U15440 (N_15440,N_15338,N_15252);
and U15441 (N_15441,N_15219,N_15393);
nor U15442 (N_15442,N_15326,N_15330);
nand U15443 (N_15443,N_15290,N_15391);
xor U15444 (N_15444,N_15235,N_15221);
xnor U15445 (N_15445,N_15309,N_15283);
xnor U15446 (N_15446,N_15298,N_15220);
nand U15447 (N_15447,N_15230,N_15213);
nand U15448 (N_15448,N_15296,N_15327);
nand U15449 (N_15449,N_15267,N_15206);
nand U15450 (N_15450,N_15365,N_15231);
nor U15451 (N_15451,N_15304,N_15223);
nand U15452 (N_15452,N_15282,N_15258);
nor U15453 (N_15453,N_15224,N_15292);
xor U15454 (N_15454,N_15208,N_15323);
nand U15455 (N_15455,N_15226,N_15335);
nand U15456 (N_15456,N_15246,N_15212);
and U15457 (N_15457,N_15353,N_15294);
or U15458 (N_15458,N_15356,N_15214);
nand U15459 (N_15459,N_15218,N_15245);
nor U15460 (N_15460,N_15369,N_15361);
xor U15461 (N_15461,N_15241,N_15270);
or U15462 (N_15462,N_15297,N_15358);
xnor U15463 (N_15463,N_15390,N_15303);
nor U15464 (N_15464,N_15203,N_15254);
nand U15465 (N_15465,N_15381,N_15352);
nand U15466 (N_15466,N_15250,N_15285);
xnor U15467 (N_15467,N_15336,N_15266);
or U15468 (N_15468,N_15337,N_15374);
nand U15469 (N_15469,N_15373,N_15240);
and U15470 (N_15470,N_15322,N_15259);
xor U15471 (N_15471,N_15260,N_15371);
nor U15472 (N_15472,N_15272,N_15275);
or U15473 (N_15473,N_15273,N_15307);
and U15474 (N_15474,N_15325,N_15329);
xor U15475 (N_15475,N_15287,N_15202);
and U15476 (N_15476,N_15350,N_15232);
nor U15477 (N_15477,N_15238,N_15264);
nor U15478 (N_15478,N_15333,N_15257);
or U15479 (N_15479,N_15346,N_15383);
xnor U15480 (N_15480,N_15313,N_15328);
and U15481 (N_15481,N_15288,N_15362);
nand U15482 (N_15482,N_15204,N_15256);
and U15483 (N_15483,N_15392,N_15345);
xnor U15484 (N_15484,N_15331,N_15271);
and U15485 (N_15485,N_15216,N_15278);
nand U15486 (N_15486,N_15237,N_15312);
nand U15487 (N_15487,N_15318,N_15360);
and U15488 (N_15488,N_15359,N_15284);
nor U15489 (N_15489,N_15281,N_15372);
xor U15490 (N_15490,N_15399,N_15339);
xor U15491 (N_15491,N_15317,N_15351);
nand U15492 (N_15492,N_15300,N_15321);
xor U15493 (N_15493,N_15375,N_15228);
xnor U15494 (N_15494,N_15210,N_15280);
or U15495 (N_15495,N_15364,N_15265);
or U15496 (N_15496,N_15334,N_15342);
or U15497 (N_15497,N_15382,N_15363);
nand U15498 (N_15498,N_15310,N_15268);
or U15499 (N_15499,N_15340,N_15209);
nor U15500 (N_15500,N_15337,N_15358);
or U15501 (N_15501,N_15231,N_15352);
xnor U15502 (N_15502,N_15345,N_15201);
and U15503 (N_15503,N_15386,N_15281);
xnor U15504 (N_15504,N_15381,N_15205);
xor U15505 (N_15505,N_15336,N_15341);
or U15506 (N_15506,N_15232,N_15206);
nand U15507 (N_15507,N_15218,N_15360);
xor U15508 (N_15508,N_15327,N_15263);
or U15509 (N_15509,N_15245,N_15219);
or U15510 (N_15510,N_15340,N_15276);
and U15511 (N_15511,N_15394,N_15335);
and U15512 (N_15512,N_15265,N_15215);
nand U15513 (N_15513,N_15271,N_15370);
nand U15514 (N_15514,N_15249,N_15358);
or U15515 (N_15515,N_15285,N_15261);
nand U15516 (N_15516,N_15327,N_15275);
xor U15517 (N_15517,N_15368,N_15361);
nor U15518 (N_15518,N_15281,N_15221);
nor U15519 (N_15519,N_15327,N_15306);
xor U15520 (N_15520,N_15365,N_15375);
nand U15521 (N_15521,N_15326,N_15283);
nor U15522 (N_15522,N_15215,N_15229);
nand U15523 (N_15523,N_15322,N_15251);
nand U15524 (N_15524,N_15241,N_15299);
nor U15525 (N_15525,N_15345,N_15298);
nor U15526 (N_15526,N_15245,N_15223);
xnor U15527 (N_15527,N_15397,N_15301);
nand U15528 (N_15528,N_15321,N_15250);
and U15529 (N_15529,N_15229,N_15350);
nor U15530 (N_15530,N_15219,N_15249);
or U15531 (N_15531,N_15356,N_15343);
xnor U15532 (N_15532,N_15313,N_15254);
or U15533 (N_15533,N_15218,N_15396);
nand U15534 (N_15534,N_15328,N_15365);
xor U15535 (N_15535,N_15271,N_15378);
or U15536 (N_15536,N_15283,N_15288);
nor U15537 (N_15537,N_15221,N_15366);
and U15538 (N_15538,N_15392,N_15365);
and U15539 (N_15539,N_15331,N_15307);
xor U15540 (N_15540,N_15360,N_15300);
xor U15541 (N_15541,N_15285,N_15201);
xnor U15542 (N_15542,N_15273,N_15344);
and U15543 (N_15543,N_15363,N_15343);
and U15544 (N_15544,N_15319,N_15397);
nor U15545 (N_15545,N_15391,N_15341);
nand U15546 (N_15546,N_15377,N_15230);
xor U15547 (N_15547,N_15242,N_15216);
or U15548 (N_15548,N_15227,N_15277);
nor U15549 (N_15549,N_15241,N_15354);
nand U15550 (N_15550,N_15205,N_15213);
nand U15551 (N_15551,N_15333,N_15374);
xor U15552 (N_15552,N_15378,N_15393);
nor U15553 (N_15553,N_15247,N_15382);
xor U15554 (N_15554,N_15374,N_15282);
nor U15555 (N_15555,N_15356,N_15394);
nand U15556 (N_15556,N_15202,N_15381);
nor U15557 (N_15557,N_15397,N_15371);
and U15558 (N_15558,N_15209,N_15210);
nor U15559 (N_15559,N_15236,N_15376);
nor U15560 (N_15560,N_15360,N_15394);
xor U15561 (N_15561,N_15246,N_15269);
nand U15562 (N_15562,N_15375,N_15303);
xnor U15563 (N_15563,N_15306,N_15339);
nor U15564 (N_15564,N_15208,N_15275);
or U15565 (N_15565,N_15344,N_15217);
and U15566 (N_15566,N_15231,N_15339);
xnor U15567 (N_15567,N_15334,N_15330);
and U15568 (N_15568,N_15361,N_15273);
xnor U15569 (N_15569,N_15329,N_15359);
nor U15570 (N_15570,N_15335,N_15299);
or U15571 (N_15571,N_15227,N_15220);
nor U15572 (N_15572,N_15308,N_15397);
and U15573 (N_15573,N_15245,N_15222);
and U15574 (N_15574,N_15325,N_15320);
or U15575 (N_15575,N_15395,N_15251);
nor U15576 (N_15576,N_15204,N_15213);
and U15577 (N_15577,N_15202,N_15260);
xor U15578 (N_15578,N_15258,N_15225);
or U15579 (N_15579,N_15363,N_15205);
nand U15580 (N_15580,N_15212,N_15330);
or U15581 (N_15581,N_15236,N_15328);
nor U15582 (N_15582,N_15345,N_15223);
xor U15583 (N_15583,N_15266,N_15306);
nand U15584 (N_15584,N_15353,N_15225);
xor U15585 (N_15585,N_15348,N_15333);
and U15586 (N_15586,N_15355,N_15251);
nand U15587 (N_15587,N_15367,N_15377);
and U15588 (N_15588,N_15308,N_15234);
nor U15589 (N_15589,N_15324,N_15240);
and U15590 (N_15590,N_15374,N_15315);
nor U15591 (N_15591,N_15265,N_15325);
xor U15592 (N_15592,N_15271,N_15280);
nor U15593 (N_15593,N_15318,N_15385);
or U15594 (N_15594,N_15323,N_15226);
nor U15595 (N_15595,N_15347,N_15259);
or U15596 (N_15596,N_15390,N_15392);
or U15597 (N_15597,N_15295,N_15388);
xor U15598 (N_15598,N_15243,N_15388);
nor U15599 (N_15599,N_15280,N_15215);
and U15600 (N_15600,N_15569,N_15406);
xnor U15601 (N_15601,N_15445,N_15500);
nand U15602 (N_15602,N_15449,N_15555);
and U15603 (N_15603,N_15462,N_15537);
and U15604 (N_15604,N_15487,N_15505);
or U15605 (N_15605,N_15433,N_15479);
nand U15606 (N_15606,N_15531,N_15522);
or U15607 (N_15607,N_15426,N_15469);
or U15608 (N_15608,N_15442,N_15436);
or U15609 (N_15609,N_15557,N_15453);
and U15610 (N_15610,N_15539,N_15415);
and U15611 (N_15611,N_15508,N_15421);
nand U15612 (N_15612,N_15596,N_15597);
xnor U15613 (N_15613,N_15548,N_15488);
nor U15614 (N_15614,N_15571,N_15441);
or U15615 (N_15615,N_15452,N_15575);
and U15616 (N_15616,N_15425,N_15551);
and U15617 (N_15617,N_15470,N_15521);
or U15618 (N_15618,N_15475,N_15430);
and U15619 (N_15619,N_15409,N_15550);
nand U15620 (N_15620,N_15559,N_15413);
or U15621 (N_15621,N_15513,N_15437);
or U15622 (N_15622,N_15553,N_15585);
nand U15623 (N_15623,N_15402,N_15407);
nand U15624 (N_15624,N_15595,N_15463);
xnor U15625 (N_15625,N_15588,N_15440);
nand U15626 (N_15626,N_15471,N_15416);
and U15627 (N_15627,N_15501,N_15561);
and U15628 (N_15628,N_15486,N_15526);
nor U15629 (N_15629,N_15458,N_15444);
nand U15630 (N_15630,N_15474,N_15494);
and U15631 (N_15631,N_15564,N_15574);
xnor U15632 (N_15632,N_15515,N_15456);
xnor U15633 (N_15633,N_15464,N_15503);
and U15634 (N_15634,N_15577,N_15461);
and U15635 (N_15635,N_15514,N_15482);
xnor U15636 (N_15636,N_15447,N_15599);
or U15637 (N_15637,N_15438,N_15586);
nor U15638 (N_15638,N_15459,N_15593);
or U15639 (N_15639,N_15431,N_15560);
nor U15640 (N_15640,N_15582,N_15420);
and U15641 (N_15641,N_15480,N_15497);
and U15642 (N_15642,N_15566,N_15589);
nor U15643 (N_15643,N_15401,N_15506);
nand U15644 (N_15644,N_15478,N_15570);
xor U15645 (N_15645,N_15519,N_15490);
or U15646 (N_15646,N_15535,N_15423);
and U15647 (N_15647,N_15411,N_15554);
nand U15648 (N_15648,N_15547,N_15516);
or U15649 (N_15649,N_15563,N_15476);
or U15650 (N_15650,N_15422,N_15405);
and U15651 (N_15651,N_15427,N_15408);
and U15652 (N_15652,N_15491,N_15528);
nand U15653 (N_15653,N_15435,N_15573);
nor U15654 (N_15654,N_15450,N_15484);
or U15655 (N_15655,N_15466,N_15568);
and U15656 (N_15656,N_15446,N_15467);
and U15657 (N_15657,N_15556,N_15529);
and U15658 (N_15658,N_15419,N_15579);
or U15659 (N_15659,N_15443,N_15572);
xor U15660 (N_15660,N_15473,N_15424);
nand U15661 (N_15661,N_15552,N_15496);
and U15662 (N_15662,N_15455,N_15502);
nand U15663 (N_15663,N_15525,N_15495);
nor U15664 (N_15664,N_15404,N_15590);
nand U15665 (N_15665,N_15460,N_15592);
and U15666 (N_15666,N_15524,N_15439);
nand U15667 (N_15667,N_15536,N_15417);
and U15668 (N_15668,N_15454,N_15581);
xnor U15669 (N_15669,N_15523,N_15498);
or U15670 (N_15670,N_15538,N_15549);
or U15671 (N_15671,N_15511,N_15512);
nand U15672 (N_15672,N_15565,N_15448);
nand U15673 (N_15673,N_15434,N_15400);
or U15674 (N_15674,N_15493,N_15534);
or U15675 (N_15675,N_15451,N_15492);
xor U15676 (N_15676,N_15418,N_15562);
or U15677 (N_15677,N_15509,N_15510);
or U15678 (N_15678,N_15591,N_15533);
or U15679 (N_15679,N_15468,N_15598);
xnor U15680 (N_15680,N_15410,N_15481);
xor U15681 (N_15681,N_15432,N_15576);
xor U15682 (N_15682,N_15540,N_15542);
nor U15683 (N_15683,N_15580,N_15594);
or U15684 (N_15684,N_15472,N_15518);
xnor U15685 (N_15685,N_15527,N_15584);
xnor U15686 (N_15686,N_15532,N_15583);
or U15687 (N_15687,N_15587,N_15429);
and U15688 (N_15688,N_15541,N_15567);
and U15689 (N_15689,N_15414,N_15507);
nand U15690 (N_15690,N_15403,N_15485);
or U15691 (N_15691,N_15483,N_15530);
and U15692 (N_15692,N_15517,N_15499);
or U15693 (N_15693,N_15544,N_15457);
xnor U15694 (N_15694,N_15489,N_15545);
xor U15695 (N_15695,N_15504,N_15578);
or U15696 (N_15696,N_15520,N_15543);
or U15697 (N_15697,N_15428,N_15412);
and U15698 (N_15698,N_15465,N_15477);
xnor U15699 (N_15699,N_15558,N_15546);
nand U15700 (N_15700,N_15581,N_15435);
nor U15701 (N_15701,N_15517,N_15472);
or U15702 (N_15702,N_15504,N_15575);
xor U15703 (N_15703,N_15486,N_15510);
nand U15704 (N_15704,N_15505,N_15467);
and U15705 (N_15705,N_15597,N_15540);
and U15706 (N_15706,N_15538,N_15406);
nand U15707 (N_15707,N_15528,N_15464);
nand U15708 (N_15708,N_15401,N_15524);
or U15709 (N_15709,N_15578,N_15409);
or U15710 (N_15710,N_15548,N_15446);
nor U15711 (N_15711,N_15451,N_15453);
nand U15712 (N_15712,N_15539,N_15408);
and U15713 (N_15713,N_15444,N_15417);
xnor U15714 (N_15714,N_15532,N_15435);
nor U15715 (N_15715,N_15476,N_15426);
xor U15716 (N_15716,N_15400,N_15561);
nor U15717 (N_15717,N_15593,N_15415);
and U15718 (N_15718,N_15547,N_15477);
xor U15719 (N_15719,N_15518,N_15563);
and U15720 (N_15720,N_15599,N_15548);
nand U15721 (N_15721,N_15522,N_15539);
or U15722 (N_15722,N_15544,N_15499);
nor U15723 (N_15723,N_15517,N_15409);
and U15724 (N_15724,N_15443,N_15417);
or U15725 (N_15725,N_15475,N_15592);
nand U15726 (N_15726,N_15506,N_15413);
nand U15727 (N_15727,N_15547,N_15419);
xor U15728 (N_15728,N_15517,N_15544);
nand U15729 (N_15729,N_15437,N_15425);
and U15730 (N_15730,N_15453,N_15569);
and U15731 (N_15731,N_15565,N_15462);
and U15732 (N_15732,N_15474,N_15581);
xnor U15733 (N_15733,N_15466,N_15443);
or U15734 (N_15734,N_15537,N_15577);
nand U15735 (N_15735,N_15542,N_15481);
xnor U15736 (N_15736,N_15420,N_15502);
and U15737 (N_15737,N_15552,N_15422);
and U15738 (N_15738,N_15418,N_15467);
and U15739 (N_15739,N_15446,N_15524);
nor U15740 (N_15740,N_15510,N_15456);
xor U15741 (N_15741,N_15474,N_15443);
nor U15742 (N_15742,N_15507,N_15467);
or U15743 (N_15743,N_15461,N_15407);
nand U15744 (N_15744,N_15577,N_15584);
and U15745 (N_15745,N_15436,N_15506);
nand U15746 (N_15746,N_15460,N_15538);
or U15747 (N_15747,N_15470,N_15549);
or U15748 (N_15748,N_15518,N_15578);
xnor U15749 (N_15749,N_15510,N_15424);
or U15750 (N_15750,N_15487,N_15418);
nor U15751 (N_15751,N_15486,N_15406);
nand U15752 (N_15752,N_15548,N_15448);
nand U15753 (N_15753,N_15518,N_15531);
nor U15754 (N_15754,N_15486,N_15574);
nor U15755 (N_15755,N_15442,N_15513);
or U15756 (N_15756,N_15506,N_15447);
or U15757 (N_15757,N_15592,N_15532);
and U15758 (N_15758,N_15494,N_15460);
and U15759 (N_15759,N_15528,N_15516);
nand U15760 (N_15760,N_15523,N_15489);
or U15761 (N_15761,N_15415,N_15558);
or U15762 (N_15762,N_15476,N_15544);
nor U15763 (N_15763,N_15505,N_15441);
nor U15764 (N_15764,N_15465,N_15420);
and U15765 (N_15765,N_15493,N_15422);
or U15766 (N_15766,N_15467,N_15572);
and U15767 (N_15767,N_15545,N_15531);
nand U15768 (N_15768,N_15523,N_15516);
xnor U15769 (N_15769,N_15483,N_15525);
nand U15770 (N_15770,N_15439,N_15429);
nand U15771 (N_15771,N_15572,N_15582);
nor U15772 (N_15772,N_15405,N_15466);
nor U15773 (N_15773,N_15525,N_15486);
nand U15774 (N_15774,N_15500,N_15417);
and U15775 (N_15775,N_15475,N_15561);
xor U15776 (N_15776,N_15444,N_15586);
or U15777 (N_15777,N_15460,N_15471);
xor U15778 (N_15778,N_15569,N_15459);
or U15779 (N_15779,N_15496,N_15520);
nor U15780 (N_15780,N_15555,N_15538);
or U15781 (N_15781,N_15426,N_15545);
and U15782 (N_15782,N_15442,N_15474);
and U15783 (N_15783,N_15506,N_15408);
nand U15784 (N_15784,N_15417,N_15556);
and U15785 (N_15785,N_15496,N_15414);
xnor U15786 (N_15786,N_15470,N_15517);
nor U15787 (N_15787,N_15529,N_15507);
nand U15788 (N_15788,N_15479,N_15455);
nand U15789 (N_15789,N_15497,N_15525);
xnor U15790 (N_15790,N_15474,N_15560);
or U15791 (N_15791,N_15500,N_15563);
nor U15792 (N_15792,N_15576,N_15587);
xnor U15793 (N_15793,N_15515,N_15482);
nor U15794 (N_15794,N_15403,N_15562);
nor U15795 (N_15795,N_15405,N_15571);
xor U15796 (N_15796,N_15579,N_15556);
or U15797 (N_15797,N_15484,N_15546);
nand U15798 (N_15798,N_15414,N_15446);
nor U15799 (N_15799,N_15435,N_15520);
nand U15800 (N_15800,N_15700,N_15755);
nor U15801 (N_15801,N_15696,N_15757);
nand U15802 (N_15802,N_15678,N_15751);
and U15803 (N_15803,N_15600,N_15787);
and U15804 (N_15804,N_15632,N_15789);
xnor U15805 (N_15805,N_15779,N_15732);
and U15806 (N_15806,N_15691,N_15672);
nor U15807 (N_15807,N_15660,N_15796);
nand U15808 (N_15808,N_15610,N_15724);
or U15809 (N_15809,N_15701,N_15611);
nand U15810 (N_15810,N_15639,N_15669);
or U15811 (N_15811,N_15729,N_15640);
xor U15812 (N_15812,N_15622,N_15728);
xor U15813 (N_15813,N_15780,N_15615);
nor U15814 (N_15814,N_15767,N_15624);
or U15815 (N_15815,N_15720,N_15708);
nor U15816 (N_15816,N_15777,N_15671);
nand U15817 (N_15817,N_15730,N_15707);
nand U15818 (N_15818,N_15731,N_15604);
or U15819 (N_15819,N_15737,N_15713);
or U15820 (N_15820,N_15771,N_15790);
or U15821 (N_15821,N_15627,N_15741);
nand U15822 (N_15822,N_15699,N_15712);
or U15823 (N_15823,N_15617,N_15653);
nand U15824 (N_15824,N_15776,N_15618);
nand U15825 (N_15825,N_15683,N_15775);
and U15826 (N_15826,N_15794,N_15655);
or U15827 (N_15827,N_15753,N_15763);
and U15828 (N_15828,N_15676,N_15652);
nand U15829 (N_15829,N_15654,N_15650);
nor U15830 (N_15830,N_15603,N_15735);
xnor U15831 (N_15831,N_15759,N_15685);
xor U15832 (N_15832,N_15733,N_15630);
nand U15833 (N_15833,N_15714,N_15710);
and U15834 (N_15834,N_15770,N_15711);
nor U15835 (N_15835,N_15721,N_15665);
and U15836 (N_15836,N_15608,N_15666);
xnor U15837 (N_15837,N_15768,N_15749);
or U15838 (N_15838,N_15716,N_15791);
or U15839 (N_15839,N_15781,N_15705);
nand U15840 (N_15840,N_15677,N_15667);
or U15841 (N_15841,N_15687,N_15747);
nor U15842 (N_15842,N_15657,N_15693);
nand U15843 (N_15843,N_15785,N_15746);
and U15844 (N_15844,N_15761,N_15798);
xnor U15845 (N_15845,N_15692,N_15760);
and U15846 (N_15846,N_15682,N_15621);
xnor U15847 (N_15847,N_15668,N_15778);
or U15848 (N_15848,N_15756,N_15612);
xnor U15849 (N_15849,N_15726,N_15722);
or U15850 (N_15850,N_15647,N_15658);
and U15851 (N_15851,N_15725,N_15616);
and U15852 (N_15852,N_15744,N_15742);
nand U15853 (N_15853,N_15606,N_15631);
nor U15854 (N_15854,N_15626,N_15629);
or U15855 (N_15855,N_15782,N_15605);
nor U15856 (N_15856,N_15634,N_15642);
nand U15857 (N_15857,N_15795,N_15689);
nor U15858 (N_15858,N_15686,N_15734);
or U15859 (N_15859,N_15706,N_15602);
xnor U15860 (N_15860,N_15613,N_15675);
xor U15861 (N_15861,N_15614,N_15679);
and U15862 (N_15862,N_15688,N_15793);
xnor U15863 (N_15863,N_15740,N_15638);
nor U15864 (N_15864,N_15628,N_15718);
and U15865 (N_15865,N_15680,N_15703);
nand U15866 (N_15866,N_15772,N_15752);
or U15867 (N_15867,N_15766,N_15697);
nor U15868 (N_15868,N_15681,N_15643);
or U15869 (N_15869,N_15695,N_15649);
and U15870 (N_15870,N_15662,N_15635);
or U15871 (N_15871,N_15673,N_15698);
or U15872 (N_15872,N_15754,N_15661);
or U15873 (N_15873,N_15601,N_15764);
nand U15874 (N_15874,N_15799,N_15792);
and U15875 (N_15875,N_15644,N_15633);
nor U15876 (N_15876,N_15797,N_15619);
xor U15877 (N_15877,N_15736,N_15715);
nand U15878 (N_15878,N_15723,N_15762);
nand U15879 (N_15879,N_15625,N_15773);
or U15880 (N_15880,N_15784,N_15709);
xnor U15881 (N_15881,N_15620,N_15663);
nor U15882 (N_15882,N_15637,N_15783);
nor U15883 (N_15883,N_15623,N_15674);
nor U15884 (N_15884,N_15769,N_15743);
and U15885 (N_15885,N_15745,N_15646);
xor U15886 (N_15886,N_15609,N_15786);
xor U15887 (N_15887,N_15738,N_15788);
xor U15888 (N_15888,N_15684,N_15694);
nand U15889 (N_15889,N_15739,N_15750);
or U15890 (N_15890,N_15664,N_15765);
xor U15891 (N_15891,N_15717,N_15719);
nor U15892 (N_15892,N_15659,N_15702);
nand U15893 (N_15893,N_15670,N_15704);
xnor U15894 (N_15894,N_15641,N_15645);
xor U15895 (N_15895,N_15748,N_15648);
or U15896 (N_15896,N_15656,N_15636);
or U15897 (N_15897,N_15607,N_15758);
xor U15898 (N_15898,N_15690,N_15727);
or U15899 (N_15899,N_15651,N_15774);
or U15900 (N_15900,N_15753,N_15749);
and U15901 (N_15901,N_15644,N_15625);
xor U15902 (N_15902,N_15621,N_15722);
nand U15903 (N_15903,N_15635,N_15700);
and U15904 (N_15904,N_15785,N_15745);
and U15905 (N_15905,N_15707,N_15602);
or U15906 (N_15906,N_15771,N_15784);
and U15907 (N_15907,N_15730,N_15640);
and U15908 (N_15908,N_15643,N_15768);
or U15909 (N_15909,N_15677,N_15732);
and U15910 (N_15910,N_15656,N_15709);
nor U15911 (N_15911,N_15721,N_15642);
and U15912 (N_15912,N_15646,N_15765);
nor U15913 (N_15913,N_15714,N_15600);
and U15914 (N_15914,N_15709,N_15681);
and U15915 (N_15915,N_15671,N_15604);
xor U15916 (N_15916,N_15714,N_15607);
or U15917 (N_15917,N_15611,N_15767);
nor U15918 (N_15918,N_15637,N_15639);
or U15919 (N_15919,N_15698,N_15790);
xnor U15920 (N_15920,N_15785,N_15789);
nand U15921 (N_15921,N_15698,N_15721);
nand U15922 (N_15922,N_15744,N_15678);
and U15923 (N_15923,N_15650,N_15661);
nand U15924 (N_15924,N_15737,N_15785);
nand U15925 (N_15925,N_15672,N_15663);
or U15926 (N_15926,N_15620,N_15611);
or U15927 (N_15927,N_15685,N_15688);
or U15928 (N_15928,N_15769,N_15686);
nor U15929 (N_15929,N_15771,N_15648);
nand U15930 (N_15930,N_15777,N_15730);
xnor U15931 (N_15931,N_15610,N_15741);
xor U15932 (N_15932,N_15617,N_15619);
nand U15933 (N_15933,N_15727,N_15670);
nor U15934 (N_15934,N_15659,N_15626);
and U15935 (N_15935,N_15600,N_15680);
nand U15936 (N_15936,N_15633,N_15754);
nor U15937 (N_15937,N_15629,N_15681);
and U15938 (N_15938,N_15678,N_15659);
nand U15939 (N_15939,N_15644,N_15600);
nor U15940 (N_15940,N_15723,N_15796);
or U15941 (N_15941,N_15788,N_15649);
and U15942 (N_15942,N_15635,N_15726);
nor U15943 (N_15943,N_15743,N_15641);
and U15944 (N_15944,N_15757,N_15706);
xnor U15945 (N_15945,N_15693,N_15644);
nor U15946 (N_15946,N_15611,N_15741);
or U15947 (N_15947,N_15764,N_15733);
or U15948 (N_15948,N_15799,N_15787);
nor U15949 (N_15949,N_15632,N_15685);
nor U15950 (N_15950,N_15772,N_15609);
or U15951 (N_15951,N_15719,N_15704);
and U15952 (N_15952,N_15649,N_15787);
and U15953 (N_15953,N_15741,N_15629);
and U15954 (N_15954,N_15777,N_15638);
nor U15955 (N_15955,N_15744,N_15643);
xor U15956 (N_15956,N_15620,N_15621);
or U15957 (N_15957,N_15751,N_15796);
xnor U15958 (N_15958,N_15767,N_15790);
nor U15959 (N_15959,N_15742,N_15765);
xor U15960 (N_15960,N_15767,N_15635);
and U15961 (N_15961,N_15707,N_15663);
and U15962 (N_15962,N_15746,N_15603);
and U15963 (N_15963,N_15623,N_15798);
or U15964 (N_15964,N_15755,N_15686);
nor U15965 (N_15965,N_15616,N_15679);
xor U15966 (N_15966,N_15745,N_15685);
nor U15967 (N_15967,N_15765,N_15677);
nand U15968 (N_15968,N_15677,N_15613);
nand U15969 (N_15969,N_15637,N_15631);
nand U15970 (N_15970,N_15764,N_15709);
nand U15971 (N_15971,N_15768,N_15794);
or U15972 (N_15972,N_15678,N_15694);
xor U15973 (N_15973,N_15729,N_15757);
or U15974 (N_15974,N_15702,N_15754);
nand U15975 (N_15975,N_15713,N_15694);
nand U15976 (N_15976,N_15653,N_15772);
and U15977 (N_15977,N_15788,N_15796);
nor U15978 (N_15978,N_15685,N_15723);
nor U15979 (N_15979,N_15661,N_15748);
nor U15980 (N_15980,N_15664,N_15654);
and U15981 (N_15981,N_15759,N_15740);
xor U15982 (N_15982,N_15722,N_15680);
xor U15983 (N_15983,N_15602,N_15747);
xor U15984 (N_15984,N_15622,N_15763);
nand U15985 (N_15985,N_15750,N_15648);
or U15986 (N_15986,N_15706,N_15638);
nand U15987 (N_15987,N_15656,N_15640);
nand U15988 (N_15988,N_15726,N_15668);
and U15989 (N_15989,N_15794,N_15647);
nor U15990 (N_15990,N_15647,N_15782);
nand U15991 (N_15991,N_15750,N_15706);
or U15992 (N_15992,N_15733,N_15756);
xor U15993 (N_15993,N_15673,N_15791);
xnor U15994 (N_15994,N_15785,N_15621);
and U15995 (N_15995,N_15728,N_15696);
and U15996 (N_15996,N_15741,N_15711);
and U15997 (N_15997,N_15692,N_15796);
nand U15998 (N_15998,N_15661,N_15729);
or U15999 (N_15999,N_15740,N_15640);
nor U16000 (N_16000,N_15999,N_15985);
xnor U16001 (N_16001,N_15898,N_15945);
xnor U16002 (N_16002,N_15861,N_15805);
nor U16003 (N_16003,N_15828,N_15986);
and U16004 (N_16004,N_15883,N_15915);
and U16005 (N_16005,N_15908,N_15943);
and U16006 (N_16006,N_15866,N_15970);
and U16007 (N_16007,N_15889,N_15809);
or U16008 (N_16008,N_15899,N_15872);
xor U16009 (N_16009,N_15918,N_15919);
and U16010 (N_16010,N_15801,N_15982);
or U16011 (N_16011,N_15856,N_15987);
nand U16012 (N_16012,N_15959,N_15927);
nor U16013 (N_16013,N_15863,N_15910);
or U16014 (N_16014,N_15834,N_15956);
or U16015 (N_16015,N_15800,N_15854);
and U16016 (N_16016,N_15818,N_15830);
nand U16017 (N_16017,N_15835,N_15853);
nand U16018 (N_16018,N_15873,N_15803);
or U16019 (N_16019,N_15868,N_15802);
and U16020 (N_16020,N_15932,N_15810);
nor U16021 (N_16021,N_15973,N_15876);
nor U16022 (N_16022,N_15971,N_15991);
xnor U16023 (N_16023,N_15848,N_15875);
or U16024 (N_16024,N_15886,N_15814);
xnor U16025 (N_16025,N_15892,N_15912);
or U16026 (N_16026,N_15832,N_15994);
and U16027 (N_16027,N_15947,N_15896);
or U16028 (N_16028,N_15894,N_15965);
nor U16029 (N_16029,N_15840,N_15869);
nor U16030 (N_16030,N_15807,N_15820);
and U16031 (N_16031,N_15909,N_15953);
nand U16032 (N_16032,N_15907,N_15995);
or U16033 (N_16033,N_15860,N_15998);
xor U16034 (N_16034,N_15992,N_15904);
and U16035 (N_16035,N_15859,N_15833);
nor U16036 (N_16036,N_15900,N_15879);
and U16037 (N_16037,N_15881,N_15989);
nor U16038 (N_16038,N_15817,N_15938);
nor U16039 (N_16039,N_15857,N_15816);
or U16040 (N_16040,N_15895,N_15822);
nand U16041 (N_16041,N_15984,N_15922);
xor U16042 (N_16042,N_15901,N_15939);
or U16043 (N_16043,N_15944,N_15906);
nand U16044 (N_16044,N_15942,N_15969);
or U16045 (N_16045,N_15951,N_15829);
nor U16046 (N_16046,N_15940,N_15815);
xnor U16047 (N_16047,N_15988,N_15937);
xor U16048 (N_16048,N_15911,N_15865);
xnor U16049 (N_16049,N_15893,N_15831);
or U16050 (N_16050,N_15924,N_15930);
nor U16051 (N_16051,N_15955,N_15950);
nor U16052 (N_16052,N_15913,N_15882);
nand U16053 (N_16053,N_15888,N_15978);
nor U16054 (N_16054,N_15825,N_15862);
nand U16055 (N_16055,N_15847,N_15972);
xor U16056 (N_16056,N_15941,N_15975);
nor U16057 (N_16057,N_15926,N_15842);
nor U16058 (N_16058,N_15871,N_15851);
xnor U16059 (N_16059,N_15877,N_15958);
and U16060 (N_16060,N_15852,N_15819);
nand U16061 (N_16061,N_15976,N_15917);
nor U16062 (N_16062,N_15845,N_15931);
nor U16063 (N_16063,N_15843,N_15983);
nor U16064 (N_16064,N_15890,N_15827);
nand U16065 (N_16065,N_15821,N_15966);
nand U16066 (N_16066,N_15903,N_15849);
and U16067 (N_16067,N_15846,N_15838);
or U16068 (N_16068,N_15874,N_15960);
nand U16069 (N_16069,N_15977,N_15864);
nand U16070 (N_16070,N_15916,N_15997);
or U16071 (N_16071,N_15885,N_15936);
nand U16072 (N_16072,N_15981,N_15884);
or U16073 (N_16073,N_15914,N_15855);
xor U16074 (N_16074,N_15850,N_15806);
nor U16075 (N_16075,N_15957,N_15920);
nand U16076 (N_16076,N_15946,N_15826);
nand U16077 (N_16077,N_15804,N_15933);
or U16078 (N_16078,N_15812,N_15929);
xnor U16079 (N_16079,N_15878,N_15887);
and U16080 (N_16080,N_15921,N_15836);
nand U16081 (N_16081,N_15928,N_15844);
nand U16082 (N_16082,N_15841,N_15858);
nor U16083 (N_16083,N_15993,N_15935);
and U16084 (N_16084,N_15962,N_15974);
and U16085 (N_16085,N_15954,N_15925);
nor U16086 (N_16086,N_15963,N_15952);
nor U16087 (N_16087,N_15811,N_15870);
xnor U16088 (N_16088,N_15823,N_15967);
xor U16089 (N_16089,N_15961,N_15964);
and U16090 (N_16090,N_15934,N_15897);
or U16091 (N_16091,N_15891,N_15979);
and U16092 (N_16092,N_15837,N_15990);
or U16093 (N_16093,N_15948,N_15905);
nor U16094 (N_16094,N_15902,N_15880);
and U16095 (N_16095,N_15813,N_15980);
or U16096 (N_16096,N_15867,N_15968);
nor U16097 (N_16097,N_15949,N_15808);
and U16098 (N_16098,N_15923,N_15839);
nor U16099 (N_16099,N_15824,N_15996);
and U16100 (N_16100,N_15960,N_15945);
xor U16101 (N_16101,N_15946,N_15878);
nor U16102 (N_16102,N_15876,N_15909);
nand U16103 (N_16103,N_15926,N_15828);
and U16104 (N_16104,N_15880,N_15897);
nor U16105 (N_16105,N_15855,N_15867);
nor U16106 (N_16106,N_15848,N_15817);
and U16107 (N_16107,N_15986,N_15832);
nor U16108 (N_16108,N_15882,N_15838);
nor U16109 (N_16109,N_15986,N_15982);
nand U16110 (N_16110,N_15852,N_15953);
or U16111 (N_16111,N_15929,N_15938);
or U16112 (N_16112,N_15866,N_15833);
xor U16113 (N_16113,N_15834,N_15896);
and U16114 (N_16114,N_15962,N_15923);
nand U16115 (N_16115,N_15914,N_15830);
and U16116 (N_16116,N_15866,N_15879);
nand U16117 (N_16117,N_15808,N_15952);
and U16118 (N_16118,N_15920,N_15954);
xnor U16119 (N_16119,N_15865,N_15803);
xor U16120 (N_16120,N_15978,N_15816);
xor U16121 (N_16121,N_15928,N_15913);
nand U16122 (N_16122,N_15851,N_15966);
xnor U16123 (N_16123,N_15914,N_15875);
and U16124 (N_16124,N_15858,N_15803);
nand U16125 (N_16125,N_15812,N_15925);
and U16126 (N_16126,N_15889,N_15974);
xor U16127 (N_16127,N_15941,N_15834);
or U16128 (N_16128,N_15958,N_15808);
and U16129 (N_16129,N_15979,N_15987);
and U16130 (N_16130,N_15830,N_15982);
and U16131 (N_16131,N_15927,N_15901);
nand U16132 (N_16132,N_15823,N_15802);
nand U16133 (N_16133,N_15921,N_15868);
nand U16134 (N_16134,N_15826,N_15915);
nor U16135 (N_16135,N_15802,N_15875);
or U16136 (N_16136,N_15987,N_15981);
xor U16137 (N_16137,N_15811,N_15927);
nand U16138 (N_16138,N_15835,N_15915);
xnor U16139 (N_16139,N_15895,N_15926);
or U16140 (N_16140,N_15910,N_15979);
nand U16141 (N_16141,N_15842,N_15972);
or U16142 (N_16142,N_15892,N_15897);
nor U16143 (N_16143,N_15958,N_15866);
xor U16144 (N_16144,N_15921,N_15886);
xnor U16145 (N_16145,N_15885,N_15942);
xnor U16146 (N_16146,N_15834,N_15872);
and U16147 (N_16147,N_15860,N_15839);
and U16148 (N_16148,N_15948,N_15913);
or U16149 (N_16149,N_15805,N_15818);
xor U16150 (N_16150,N_15904,N_15975);
or U16151 (N_16151,N_15828,N_15881);
nand U16152 (N_16152,N_15993,N_15975);
nor U16153 (N_16153,N_15822,N_15928);
xnor U16154 (N_16154,N_15838,N_15868);
xor U16155 (N_16155,N_15888,N_15907);
nor U16156 (N_16156,N_15968,N_15881);
xnor U16157 (N_16157,N_15889,N_15943);
xor U16158 (N_16158,N_15975,N_15806);
nand U16159 (N_16159,N_15882,N_15860);
and U16160 (N_16160,N_15821,N_15938);
and U16161 (N_16161,N_15868,N_15903);
or U16162 (N_16162,N_15959,N_15864);
xnor U16163 (N_16163,N_15826,N_15855);
and U16164 (N_16164,N_15870,N_15857);
or U16165 (N_16165,N_15971,N_15883);
and U16166 (N_16166,N_15981,N_15875);
xnor U16167 (N_16167,N_15942,N_15992);
nor U16168 (N_16168,N_15808,N_15919);
or U16169 (N_16169,N_15880,N_15863);
nor U16170 (N_16170,N_15877,N_15928);
xor U16171 (N_16171,N_15856,N_15955);
and U16172 (N_16172,N_15999,N_15874);
and U16173 (N_16173,N_15884,N_15900);
or U16174 (N_16174,N_15942,N_15993);
nor U16175 (N_16175,N_15844,N_15825);
or U16176 (N_16176,N_15824,N_15937);
nor U16177 (N_16177,N_15823,N_15917);
xor U16178 (N_16178,N_15944,N_15892);
or U16179 (N_16179,N_15917,N_15897);
and U16180 (N_16180,N_15958,N_15961);
nand U16181 (N_16181,N_15819,N_15918);
nand U16182 (N_16182,N_15865,N_15995);
or U16183 (N_16183,N_15991,N_15944);
xor U16184 (N_16184,N_15851,N_15993);
and U16185 (N_16185,N_15949,N_15993);
and U16186 (N_16186,N_15952,N_15851);
nor U16187 (N_16187,N_15883,N_15888);
nand U16188 (N_16188,N_15949,N_15905);
and U16189 (N_16189,N_15951,N_15969);
and U16190 (N_16190,N_15943,N_15826);
xor U16191 (N_16191,N_15931,N_15857);
nor U16192 (N_16192,N_15982,N_15863);
and U16193 (N_16193,N_15987,N_15967);
nand U16194 (N_16194,N_15975,N_15945);
xnor U16195 (N_16195,N_15876,N_15847);
nand U16196 (N_16196,N_15819,N_15899);
and U16197 (N_16197,N_15801,N_15800);
or U16198 (N_16198,N_15980,N_15931);
or U16199 (N_16199,N_15956,N_15974);
nand U16200 (N_16200,N_16032,N_16062);
or U16201 (N_16201,N_16095,N_16077);
xor U16202 (N_16202,N_16158,N_16033);
nor U16203 (N_16203,N_16053,N_16137);
nor U16204 (N_16204,N_16189,N_16117);
nand U16205 (N_16205,N_16188,N_16193);
xnor U16206 (N_16206,N_16026,N_16004);
nand U16207 (N_16207,N_16112,N_16041);
nand U16208 (N_16208,N_16142,N_16124);
nor U16209 (N_16209,N_16145,N_16102);
and U16210 (N_16210,N_16114,N_16167);
xnor U16211 (N_16211,N_16049,N_16156);
and U16212 (N_16212,N_16161,N_16196);
or U16213 (N_16213,N_16022,N_16164);
nor U16214 (N_16214,N_16039,N_16088);
and U16215 (N_16215,N_16075,N_16104);
and U16216 (N_16216,N_16173,N_16105);
nor U16217 (N_16217,N_16072,N_16118);
nand U16218 (N_16218,N_16011,N_16038);
nand U16219 (N_16219,N_16058,N_16151);
nor U16220 (N_16220,N_16127,N_16150);
nor U16221 (N_16221,N_16012,N_16037);
and U16222 (N_16222,N_16110,N_16008);
or U16223 (N_16223,N_16101,N_16094);
nor U16224 (N_16224,N_16185,N_16071);
nor U16225 (N_16225,N_16122,N_16040);
xor U16226 (N_16226,N_16093,N_16177);
and U16227 (N_16227,N_16030,N_16163);
or U16228 (N_16228,N_16172,N_16059);
nor U16229 (N_16229,N_16152,N_16194);
nor U16230 (N_16230,N_16016,N_16149);
nand U16231 (N_16231,N_16089,N_16179);
xnor U16232 (N_16232,N_16159,N_16096);
and U16233 (N_16233,N_16092,N_16044);
or U16234 (N_16234,N_16045,N_16182);
nand U16235 (N_16235,N_16147,N_16010);
nor U16236 (N_16236,N_16090,N_16064);
xor U16237 (N_16237,N_16057,N_16065);
nor U16238 (N_16238,N_16115,N_16015);
xnor U16239 (N_16239,N_16157,N_16166);
nor U16240 (N_16240,N_16153,N_16107);
nor U16241 (N_16241,N_16160,N_16195);
or U16242 (N_16242,N_16046,N_16130);
xnor U16243 (N_16243,N_16029,N_16125);
nor U16244 (N_16244,N_16055,N_16025);
and U16245 (N_16245,N_16132,N_16097);
xnor U16246 (N_16246,N_16080,N_16054);
or U16247 (N_16247,N_16141,N_16067);
and U16248 (N_16248,N_16148,N_16126);
or U16249 (N_16249,N_16063,N_16139);
nand U16250 (N_16250,N_16129,N_16134);
nor U16251 (N_16251,N_16081,N_16003);
or U16252 (N_16252,N_16165,N_16131);
xor U16253 (N_16253,N_16001,N_16184);
or U16254 (N_16254,N_16191,N_16079);
xor U16255 (N_16255,N_16047,N_16070);
nand U16256 (N_16256,N_16060,N_16140);
nor U16257 (N_16257,N_16176,N_16128);
or U16258 (N_16258,N_16168,N_16024);
nand U16259 (N_16259,N_16048,N_16146);
nor U16260 (N_16260,N_16043,N_16017);
xor U16261 (N_16261,N_16109,N_16169);
xor U16262 (N_16262,N_16183,N_16187);
xor U16263 (N_16263,N_16068,N_16190);
and U16264 (N_16264,N_16056,N_16121);
nor U16265 (N_16265,N_16116,N_16018);
nand U16266 (N_16266,N_16181,N_16023);
and U16267 (N_16267,N_16174,N_16136);
and U16268 (N_16268,N_16050,N_16098);
or U16269 (N_16269,N_16027,N_16103);
or U16270 (N_16270,N_16019,N_16082);
nor U16271 (N_16271,N_16028,N_16086);
and U16272 (N_16272,N_16135,N_16155);
nand U16273 (N_16273,N_16006,N_16111);
xnor U16274 (N_16274,N_16061,N_16034);
nand U16275 (N_16275,N_16171,N_16078);
xnor U16276 (N_16276,N_16123,N_16178);
nand U16277 (N_16277,N_16162,N_16036);
nand U16278 (N_16278,N_16084,N_16180);
nand U16279 (N_16279,N_16000,N_16113);
nand U16280 (N_16280,N_16031,N_16020);
xnor U16281 (N_16281,N_16073,N_16052);
xor U16282 (N_16282,N_16143,N_16076);
nand U16283 (N_16283,N_16138,N_16144);
and U16284 (N_16284,N_16051,N_16192);
nand U16285 (N_16285,N_16100,N_16106);
or U16286 (N_16286,N_16085,N_16035);
or U16287 (N_16287,N_16013,N_16014);
xnor U16288 (N_16288,N_16021,N_16133);
nand U16289 (N_16289,N_16066,N_16099);
nand U16290 (N_16290,N_16087,N_16175);
nand U16291 (N_16291,N_16009,N_16198);
or U16292 (N_16292,N_16074,N_16083);
nand U16293 (N_16293,N_16007,N_16197);
xnor U16294 (N_16294,N_16108,N_16119);
and U16295 (N_16295,N_16120,N_16002);
or U16296 (N_16296,N_16091,N_16069);
xnor U16297 (N_16297,N_16186,N_16199);
xnor U16298 (N_16298,N_16170,N_16154);
nand U16299 (N_16299,N_16042,N_16005);
and U16300 (N_16300,N_16146,N_16160);
nor U16301 (N_16301,N_16093,N_16001);
nor U16302 (N_16302,N_16006,N_16029);
or U16303 (N_16303,N_16001,N_16029);
nor U16304 (N_16304,N_16052,N_16031);
or U16305 (N_16305,N_16110,N_16000);
nand U16306 (N_16306,N_16180,N_16155);
and U16307 (N_16307,N_16001,N_16128);
nand U16308 (N_16308,N_16128,N_16167);
or U16309 (N_16309,N_16161,N_16055);
xnor U16310 (N_16310,N_16188,N_16148);
or U16311 (N_16311,N_16063,N_16124);
and U16312 (N_16312,N_16087,N_16050);
nand U16313 (N_16313,N_16019,N_16034);
nand U16314 (N_16314,N_16008,N_16037);
nor U16315 (N_16315,N_16102,N_16056);
xor U16316 (N_16316,N_16045,N_16013);
xor U16317 (N_16317,N_16021,N_16079);
or U16318 (N_16318,N_16126,N_16140);
nand U16319 (N_16319,N_16021,N_16017);
nand U16320 (N_16320,N_16162,N_16008);
nand U16321 (N_16321,N_16149,N_16141);
or U16322 (N_16322,N_16090,N_16042);
nor U16323 (N_16323,N_16028,N_16122);
xnor U16324 (N_16324,N_16067,N_16041);
and U16325 (N_16325,N_16075,N_16177);
nor U16326 (N_16326,N_16046,N_16146);
and U16327 (N_16327,N_16118,N_16147);
nand U16328 (N_16328,N_16030,N_16156);
xnor U16329 (N_16329,N_16140,N_16170);
or U16330 (N_16330,N_16121,N_16170);
or U16331 (N_16331,N_16055,N_16167);
or U16332 (N_16332,N_16022,N_16037);
or U16333 (N_16333,N_16022,N_16020);
nor U16334 (N_16334,N_16017,N_16065);
xnor U16335 (N_16335,N_16195,N_16012);
and U16336 (N_16336,N_16193,N_16183);
and U16337 (N_16337,N_16067,N_16155);
nand U16338 (N_16338,N_16108,N_16165);
or U16339 (N_16339,N_16071,N_16075);
nand U16340 (N_16340,N_16162,N_16150);
nand U16341 (N_16341,N_16137,N_16154);
nor U16342 (N_16342,N_16102,N_16144);
and U16343 (N_16343,N_16159,N_16025);
nor U16344 (N_16344,N_16047,N_16190);
or U16345 (N_16345,N_16008,N_16035);
xor U16346 (N_16346,N_16080,N_16085);
nor U16347 (N_16347,N_16129,N_16062);
nor U16348 (N_16348,N_16033,N_16126);
nand U16349 (N_16349,N_16062,N_16141);
nand U16350 (N_16350,N_16118,N_16139);
nand U16351 (N_16351,N_16132,N_16008);
nand U16352 (N_16352,N_16161,N_16079);
and U16353 (N_16353,N_16151,N_16136);
nand U16354 (N_16354,N_16028,N_16033);
nand U16355 (N_16355,N_16089,N_16017);
and U16356 (N_16356,N_16198,N_16155);
nor U16357 (N_16357,N_16019,N_16137);
nand U16358 (N_16358,N_16047,N_16026);
or U16359 (N_16359,N_16101,N_16172);
nor U16360 (N_16360,N_16129,N_16100);
xnor U16361 (N_16361,N_16168,N_16151);
xnor U16362 (N_16362,N_16004,N_16120);
nor U16363 (N_16363,N_16120,N_16189);
and U16364 (N_16364,N_16117,N_16057);
nor U16365 (N_16365,N_16140,N_16091);
nand U16366 (N_16366,N_16018,N_16091);
or U16367 (N_16367,N_16022,N_16130);
or U16368 (N_16368,N_16164,N_16035);
nand U16369 (N_16369,N_16159,N_16111);
nand U16370 (N_16370,N_16089,N_16150);
nand U16371 (N_16371,N_16083,N_16075);
and U16372 (N_16372,N_16169,N_16011);
nand U16373 (N_16373,N_16126,N_16031);
nor U16374 (N_16374,N_16057,N_16196);
and U16375 (N_16375,N_16082,N_16178);
nand U16376 (N_16376,N_16115,N_16118);
nor U16377 (N_16377,N_16053,N_16021);
or U16378 (N_16378,N_16023,N_16018);
nand U16379 (N_16379,N_16170,N_16005);
xor U16380 (N_16380,N_16072,N_16009);
xor U16381 (N_16381,N_16109,N_16072);
nor U16382 (N_16382,N_16122,N_16185);
nor U16383 (N_16383,N_16064,N_16019);
nand U16384 (N_16384,N_16142,N_16054);
or U16385 (N_16385,N_16072,N_16114);
nor U16386 (N_16386,N_16160,N_16012);
nor U16387 (N_16387,N_16092,N_16165);
xor U16388 (N_16388,N_16134,N_16158);
or U16389 (N_16389,N_16000,N_16177);
nand U16390 (N_16390,N_16167,N_16025);
or U16391 (N_16391,N_16083,N_16079);
nand U16392 (N_16392,N_16198,N_16053);
nand U16393 (N_16393,N_16167,N_16092);
xor U16394 (N_16394,N_16119,N_16165);
nand U16395 (N_16395,N_16087,N_16071);
nor U16396 (N_16396,N_16085,N_16123);
or U16397 (N_16397,N_16108,N_16053);
nand U16398 (N_16398,N_16150,N_16059);
xnor U16399 (N_16399,N_16125,N_16122);
nand U16400 (N_16400,N_16258,N_16385);
and U16401 (N_16401,N_16346,N_16205);
nor U16402 (N_16402,N_16314,N_16269);
and U16403 (N_16403,N_16274,N_16340);
or U16404 (N_16404,N_16290,N_16344);
nand U16405 (N_16405,N_16337,N_16382);
and U16406 (N_16406,N_16345,N_16372);
nand U16407 (N_16407,N_16300,N_16243);
nand U16408 (N_16408,N_16284,N_16266);
and U16409 (N_16409,N_16376,N_16309);
or U16410 (N_16410,N_16220,N_16260);
and U16411 (N_16411,N_16254,N_16371);
xnor U16412 (N_16412,N_16328,N_16226);
xor U16413 (N_16413,N_16280,N_16292);
and U16414 (N_16414,N_16291,N_16281);
and U16415 (N_16415,N_16233,N_16366);
nor U16416 (N_16416,N_16253,N_16207);
and U16417 (N_16417,N_16246,N_16302);
nor U16418 (N_16418,N_16377,N_16388);
or U16419 (N_16419,N_16327,N_16383);
nor U16420 (N_16420,N_16390,N_16311);
and U16421 (N_16421,N_16235,N_16204);
xnor U16422 (N_16422,N_16331,N_16395);
nand U16423 (N_16423,N_16361,N_16293);
xor U16424 (N_16424,N_16347,N_16353);
nand U16425 (N_16425,N_16209,N_16273);
nor U16426 (N_16426,N_16219,N_16329);
nor U16427 (N_16427,N_16267,N_16387);
or U16428 (N_16428,N_16319,N_16248);
and U16429 (N_16429,N_16301,N_16368);
nand U16430 (N_16430,N_16306,N_16268);
xor U16431 (N_16431,N_16252,N_16239);
and U16432 (N_16432,N_16283,N_16285);
nor U16433 (N_16433,N_16223,N_16230);
nand U16434 (N_16434,N_16249,N_16251);
nor U16435 (N_16435,N_16365,N_16245);
and U16436 (N_16436,N_16375,N_16271);
nand U16437 (N_16437,N_16351,N_16210);
xnor U16438 (N_16438,N_16272,N_16338);
xor U16439 (N_16439,N_16391,N_16392);
xnor U16440 (N_16440,N_16255,N_16213);
nor U16441 (N_16441,N_16221,N_16229);
nor U16442 (N_16442,N_16201,N_16240);
nor U16443 (N_16443,N_16307,N_16325);
nor U16444 (N_16444,N_16367,N_16288);
nand U16445 (N_16445,N_16242,N_16360);
and U16446 (N_16446,N_16378,N_16282);
or U16447 (N_16447,N_16217,N_16208);
and U16448 (N_16448,N_16363,N_16312);
or U16449 (N_16449,N_16355,N_16370);
nand U16450 (N_16450,N_16305,N_16335);
nand U16451 (N_16451,N_16278,N_16234);
xnor U16452 (N_16452,N_16238,N_16336);
and U16453 (N_16453,N_16275,N_16295);
nand U16454 (N_16454,N_16334,N_16308);
and U16455 (N_16455,N_16237,N_16236);
or U16456 (N_16456,N_16304,N_16381);
nand U16457 (N_16457,N_16399,N_16202);
or U16458 (N_16458,N_16206,N_16393);
and U16459 (N_16459,N_16369,N_16222);
nor U16460 (N_16460,N_16384,N_16320);
nand U16461 (N_16461,N_16277,N_16398);
nor U16462 (N_16462,N_16287,N_16270);
nand U16463 (N_16463,N_16321,N_16261);
xnor U16464 (N_16464,N_16330,N_16265);
nand U16465 (N_16465,N_16386,N_16303);
or U16466 (N_16466,N_16232,N_16279);
nand U16467 (N_16467,N_16379,N_16244);
xor U16468 (N_16468,N_16215,N_16397);
xor U16469 (N_16469,N_16348,N_16374);
nor U16470 (N_16470,N_16396,N_16228);
xor U16471 (N_16471,N_16225,N_16324);
nand U16472 (N_16472,N_16256,N_16212);
or U16473 (N_16473,N_16394,N_16241);
nor U16474 (N_16474,N_16299,N_16264);
nand U16475 (N_16475,N_16263,N_16200);
nand U16476 (N_16476,N_16203,N_16296);
nand U16477 (N_16477,N_16316,N_16364);
or U16478 (N_16478,N_16373,N_16250);
and U16479 (N_16479,N_16313,N_16317);
nand U16480 (N_16480,N_16343,N_16333);
and U16481 (N_16481,N_16218,N_16259);
xor U16482 (N_16482,N_16354,N_16318);
and U16483 (N_16483,N_16276,N_16350);
and U16484 (N_16484,N_16341,N_16357);
or U16485 (N_16485,N_16289,N_16227);
or U16486 (N_16486,N_16332,N_16214);
nand U16487 (N_16487,N_16315,N_16322);
nand U16488 (N_16488,N_16297,N_16342);
or U16489 (N_16489,N_16298,N_16362);
nor U16490 (N_16490,N_16211,N_16358);
nor U16491 (N_16491,N_16359,N_16380);
and U16492 (N_16492,N_16294,N_16216);
and U16493 (N_16493,N_16323,N_16352);
or U16494 (N_16494,N_16286,N_16231);
nand U16495 (N_16495,N_16339,N_16247);
or U16496 (N_16496,N_16356,N_16262);
or U16497 (N_16497,N_16310,N_16389);
xor U16498 (N_16498,N_16224,N_16257);
nand U16499 (N_16499,N_16349,N_16326);
xnor U16500 (N_16500,N_16377,N_16244);
or U16501 (N_16501,N_16258,N_16222);
nor U16502 (N_16502,N_16351,N_16254);
xnor U16503 (N_16503,N_16272,N_16378);
and U16504 (N_16504,N_16339,N_16350);
nor U16505 (N_16505,N_16321,N_16228);
and U16506 (N_16506,N_16203,N_16341);
and U16507 (N_16507,N_16297,N_16320);
or U16508 (N_16508,N_16262,N_16357);
or U16509 (N_16509,N_16284,N_16336);
xor U16510 (N_16510,N_16285,N_16307);
or U16511 (N_16511,N_16273,N_16205);
nand U16512 (N_16512,N_16342,N_16205);
or U16513 (N_16513,N_16227,N_16235);
nor U16514 (N_16514,N_16321,N_16274);
xnor U16515 (N_16515,N_16298,N_16204);
or U16516 (N_16516,N_16285,N_16361);
or U16517 (N_16517,N_16277,N_16387);
and U16518 (N_16518,N_16314,N_16389);
nand U16519 (N_16519,N_16202,N_16318);
nand U16520 (N_16520,N_16273,N_16217);
or U16521 (N_16521,N_16208,N_16259);
nor U16522 (N_16522,N_16308,N_16317);
and U16523 (N_16523,N_16283,N_16321);
or U16524 (N_16524,N_16376,N_16276);
or U16525 (N_16525,N_16379,N_16229);
nor U16526 (N_16526,N_16265,N_16257);
nor U16527 (N_16527,N_16223,N_16370);
nand U16528 (N_16528,N_16276,N_16358);
nand U16529 (N_16529,N_16364,N_16214);
xnor U16530 (N_16530,N_16249,N_16354);
xnor U16531 (N_16531,N_16347,N_16218);
or U16532 (N_16532,N_16201,N_16262);
nor U16533 (N_16533,N_16348,N_16272);
or U16534 (N_16534,N_16299,N_16237);
xnor U16535 (N_16535,N_16352,N_16303);
or U16536 (N_16536,N_16373,N_16339);
nor U16537 (N_16537,N_16237,N_16305);
or U16538 (N_16538,N_16354,N_16369);
nor U16539 (N_16539,N_16281,N_16296);
nor U16540 (N_16540,N_16213,N_16246);
xnor U16541 (N_16541,N_16236,N_16228);
or U16542 (N_16542,N_16345,N_16251);
nand U16543 (N_16543,N_16315,N_16266);
or U16544 (N_16544,N_16282,N_16381);
or U16545 (N_16545,N_16355,N_16313);
or U16546 (N_16546,N_16254,N_16262);
and U16547 (N_16547,N_16230,N_16384);
nor U16548 (N_16548,N_16231,N_16269);
or U16549 (N_16549,N_16274,N_16271);
and U16550 (N_16550,N_16327,N_16216);
and U16551 (N_16551,N_16313,N_16376);
nand U16552 (N_16552,N_16247,N_16257);
and U16553 (N_16553,N_16296,N_16384);
nor U16554 (N_16554,N_16277,N_16351);
and U16555 (N_16555,N_16269,N_16258);
xor U16556 (N_16556,N_16332,N_16294);
nand U16557 (N_16557,N_16253,N_16212);
xnor U16558 (N_16558,N_16382,N_16274);
or U16559 (N_16559,N_16271,N_16229);
or U16560 (N_16560,N_16381,N_16316);
nand U16561 (N_16561,N_16306,N_16258);
and U16562 (N_16562,N_16288,N_16354);
and U16563 (N_16563,N_16221,N_16318);
and U16564 (N_16564,N_16310,N_16396);
nand U16565 (N_16565,N_16219,N_16209);
nor U16566 (N_16566,N_16283,N_16393);
nand U16567 (N_16567,N_16278,N_16217);
nand U16568 (N_16568,N_16228,N_16286);
nor U16569 (N_16569,N_16222,N_16356);
or U16570 (N_16570,N_16384,N_16377);
nor U16571 (N_16571,N_16251,N_16378);
xor U16572 (N_16572,N_16374,N_16333);
nor U16573 (N_16573,N_16370,N_16281);
and U16574 (N_16574,N_16278,N_16362);
nor U16575 (N_16575,N_16382,N_16297);
or U16576 (N_16576,N_16213,N_16248);
or U16577 (N_16577,N_16299,N_16284);
xnor U16578 (N_16578,N_16355,N_16270);
and U16579 (N_16579,N_16342,N_16262);
and U16580 (N_16580,N_16327,N_16315);
or U16581 (N_16581,N_16368,N_16366);
nand U16582 (N_16582,N_16381,N_16237);
or U16583 (N_16583,N_16235,N_16334);
or U16584 (N_16584,N_16382,N_16291);
and U16585 (N_16585,N_16270,N_16209);
xor U16586 (N_16586,N_16318,N_16300);
nand U16587 (N_16587,N_16215,N_16331);
xor U16588 (N_16588,N_16314,N_16377);
and U16589 (N_16589,N_16286,N_16323);
nand U16590 (N_16590,N_16341,N_16371);
or U16591 (N_16591,N_16382,N_16305);
nand U16592 (N_16592,N_16392,N_16397);
xor U16593 (N_16593,N_16393,N_16291);
nand U16594 (N_16594,N_16226,N_16314);
xor U16595 (N_16595,N_16321,N_16357);
nand U16596 (N_16596,N_16240,N_16354);
xor U16597 (N_16597,N_16329,N_16264);
or U16598 (N_16598,N_16239,N_16212);
and U16599 (N_16599,N_16246,N_16398);
or U16600 (N_16600,N_16583,N_16461);
nand U16601 (N_16601,N_16518,N_16510);
nor U16602 (N_16602,N_16590,N_16435);
nor U16603 (N_16603,N_16584,N_16530);
or U16604 (N_16604,N_16438,N_16483);
xor U16605 (N_16605,N_16443,N_16559);
or U16606 (N_16606,N_16488,N_16515);
xnor U16607 (N_16607,N_16407,N_16522);
or U16608 (N_16608,N_16529,N_16411);
nor U16609 (N_16609,N_16416,N_16497);
or U16610 (N_16610,N_16418,N_16534);
and U16611 (N_16611,N_16444,N_16553);
nor U16612 (N_16612,N_16431,N_16539);
nor U16613 (N_16613,N_16567,N_16524);
nand U16614 (N_16614,N_16410,N_16491);
nand U16615 (N_16615,N_16588,N_16420);
nand U16616 (N_16616,N_16423,N_16500);
nor U16617 (N_16617,N_16473,N_16544);
nor U16618 (N_16618,N_16472,N_16533);
nor U16619 (N_16619,N_16548,N_16597);
nor U16620 (N_16620,N_16437,N_16477);
nand U16621 (N_16621,N_16479,N_16469);
or U16622 (N_16622,N_16463,N_16555);
and U16623 (N_16623,N_16591,N_16512);
xor U16624 (N_16624,N_16465,N_16426);
or U16625 (N_16625,N_16458,N_16536);
nand U16626 (N_16626,N_16422,N_16504);
nand U16627 (N_16627,N_16576,N_16565);
xnor U16628 (N_16628,N_16511,N_16467);
nand U16629 (N_16629,N_16439,N_16414);
or U16630 (N_16630,N_16447,N_16545);
nor U16631 (N_16631,N_16503,N_16543);
nor U16632 (N_16632,N_16489,N_16546);
and U16633 (N_16633,N_16542,N_16450);
nor U16634 (N_16634,N_16428,N_16487);
nor U16635 (N_16635,N_16560,N_16550);
or U16636 (N_16636,N_16580,N_16474);
or U16637 (N_16637,N_16404,N_16434);
xnor U16638 (N_16638,N_16578,N_16554);
or U16639 (N_16639,N_16599,N_16471);
nor U16640 (N_16640,N_16528,N_16574);
nor U16641 (N_16641,N_16573,N_16502);
xor U16642 (N_16642,N_16486,N_16401);
nor U16643 (N_16643,N_16424,N_16509);
nor U16644 (N_16644,N_16594,N_16452);
nand U16645 (N_16645,N_16442,N_16476);
nand U16646 (N_16646,N_16531,N_16429);
and U16647 (N_16647,N_16457,N_16492);
nor U16648 (N_16648,N_16540,N_16455);
xnor U16649 (N_16649,N_16592,N_16495);
nand U16650 (N_16650,N_16541,N_16448);
nor U16651 (N_16651,N_16451,N_16508);
nand U16652 (N_16652,N_16566,N_16460);
xnor U16653 (N_16653,N_16482,N_16570);
nand U16654 (N_16654,N_16409,N_16552);
or U16655 (N_16655,N_16490,N_16568);
nand U16656 (N_16656,N_16513,N_16475);
or U16657 (N_16657,N_16517,N_16516);
nand U16658 (N_16658,N_16433,N_16572);
xnor U16659 (N_16659,N_16470,N_16499);
or U16660 (N_16660,N_16459,N_16532);
nand U16661 (N_16661,N_16419,N_16596);
or U16662 (N_16662,N_16595,N_16480);
nor U16663 (N_16663,N_16462,N_16408);
nand U16664 (N_16664,N_16558,N_16525);
or U16665 (N_16665,N_16430,N_16449);
xor U16666 (N_16666,N_16454,N_16582);
nor U16667 (N_16667,N_16400,N_16445);
or U16668 (N_16668,N_16405,N_16575);
nor U16669 (N_16669,N_16577,N_16535);
xnor U16670 (N_16670,N_16579,N_16406);
or U16671 (N_16671,N_16417,N_16468);
nand U16672 (N_16672,N_16441,N_16571);
and U16673 (N_16673,N_16464,N_16507);
and U16674 (N_16674,N_16557,N_16569);
and U16675 (N_16675,N_16563,N_16506);
xnor U16676 (N_16676,N_16466,N_16593);
nand U16677 (N_16677,N_16586,N_16425);
xnor U16678 (N_16678,N_16427,N_16456);
or U16679 (N_16679,N_16432,N_16523);
and U16680 (N_16680,N_16562,N_16478);
nand U16681 (N_16681,N_16527,N_16453);
and U16682 (N_16682,N_16440,N_16538);
nor U16683 (N_16683,N_16587,N_16520);
and U16684 (N_16684,N_16521,N_16537);
nor U16685 (N_16685,N_16484,N_16561);
and U16686 (N_16686,N_16412,N_16446);
and U16687 (N_16687,N_16549,N_16403);
xnor U16688 (N_16688,N_16581,N_16505);
nor U16689 (N_16689,N_16551,N_16421);
or U16690 (N_16690,N_16514,N_16498);
nand U16691 (N_16691,N_16519,N_16402);
nor U16692 (N_16692,N_16413,N_16494);
or U16693 (N_16693,N_16481,N_16496);
nor U16694 (N_16694,N_16493,N_16585);
or U16695 (N_16695,N_16436,N_16526);
nand U16696 (N_16696,N_16415,N_16598);
or U16697 (N_16697,N_16589,N_16556);
or U16698 (N_16698,N_16547,N_16485);
or U16699 (N_16699,N_16501,N_16564);
or U16700 (N_16700,N_16530,N_16454);
xnor U16701 (N_16701,N_16569,N_16462);
and U16702 (N_16702,N_16486,N_16589);
nand U16703 (N_16703,N_16542,N_16530);
xor U16704 (N_16704,N_16520,N_16476);
nor U16705 (N_16705,N_16522,N_16514);
nand U16706 (N_16706,N_16417,N_16501);
nor U16707 (N_16707,N_16425,N_16599);
nand U16708 (N_16708,N_16571,N_16409);
nor U16709 (N_16709,N_16536,N_16488);
nor U16710 (N_16710,N_16403,N_16529);
or U16711 (N_16711,N_16574,N_16577);
and U16712 (N_16712,N_16413,N_16481);
nand U16713 (N_16713,N_16533,N_16470);
and U16714 (N_16714,N_16510,N_16541);
and U16715 (N_16715,N_16452,N_16471);
and U16716 (N_16716,N_16412,N_16527);
or U16717 (N_16717,N_16401,N_16569);
nor U16718 (N_16718,N_16585,N_16548);
nor U16719 (N_16719,N_16495,N_16568);
nor U16720 (N_16720,N_16495,N_16598);
and U16721 (N_16721,N_16563,N_16531);
xor U16722 (N_16722,N_16553,N_16568);
and U16723 (N_16723,N_16457,N_16519);
xnor U16724 (N_16724,N_16544,N_16519);
xnor U16725 (N_16725,N_16535,N_16406);
or U16726 (N_16726,N_16470,N_16438);
xnor U16727 (N_16727,N_16451,N_16484);
nor U16728 (N_16728,N_16433,N_16592);
and U16729 (N_16729,N_16495,N_16522);
nand U16730 (N_16730,N_16578,N_16493);
xor U16731 (N_16731,N_16477,N_16566);
or U16732 (N_16732,N_16567,N_16433);
and U16733 (N_16733,N_16514,N_16546);
nand U16734 (N_16734,N_16474,N_16517);
xor U16735 (N_16735,N_16429,N_16505);
and U16736 (N_16736,N_16465,N_16444);
nor U16737 (N_16737,N_16515,N_16485);
nand U16738 (N_16738,N_16548,N_16420);
nor U16739 (N_16739,N_16509,N_16473);
nand U16740 (N_16740,N_16488,N_16489);
or U16741 (N_16741,N_16538,N_16542);
nor U16742 (N_16742,N_16547,N_16483);
xor U16743 (N_16743,N_16455,N_16481);
xor U16744 (N_16744,N_16449,N_16536);
and U16745 (N_16745,N_16403,N_16496);
and U16746 (N_16746,N_16556,N_16425);
or U16747 (N_16747,N_16565,N_16524);
nor U16748 (N_16748,N_16426,N_16515);
xor U16749 (N_16749,N_16532,N_16401);
or U16750 (N_16750,N_16530,N_16573);
and U16751 (N_16751,N_16478,N_16450);
nand U16752 (N_16752,N_16522,N_16556);
or U16753 (N_16753,N_16587,N_16482);
xnor U16754 (N_16754,N_16510,N_16585);
xnor U16755 (N_16755,N_16444,N_16449);
or U16756 (N_16756,N_16541,N_16497);
nor U16757 (N_16757,N_16415,N_16402);
and U16758 (N_16758,N_16473,N_16578);
or U16759 (N_16759,N_16404,N_16406);
nor U16760 (N_16760,N_16409,N_16481);
nand U16761 (N_16761,N_16411,N_16450);
nand U16762 (N_16762,N_16493,N_16599);
or U16763 (N_16763,N_16421,N_16509);
or U16764 (N_16764,N_16522,N_16442);
and U16765 (N_16765,N_16465,N_16524);
xor U16766 (N_16766,N_16414,N_16461);
xor U16767 (N_16767,N_16594,N_16481);
xnor U16768 (N_16768,N_16539,N_16461);
nor U16769 (N_16769,N_16400,N_16453);
xnor U16770 (N_16770,N_16467,N_16589);
nand U16771 (N_16771,N_16474,N_16520);
and U16772 (N_16772,N_16593,N_16504);
or U16773 (N_16773,N_16526,N_16403);
xnor U16774 (N_16774,N_16507,N_16535);
nand U16775 (N_16775,N_16518,N_16421);
or U16776 (N_16776,N_16474,N_16591);
nor U16777 (N_16777,N_16427,N_16447);
or U16778 (N_16778,N_16570,N_16430);
or U16779 (N_16779,N_16566,N_16406);
or U16780 (N_16780,N_16488,N_16571);
and U16781 (N_16781,N_16560,N_16526);
xnor U16782 (N_16782,N_16481,N_16422);
nor U16783 (N_16783,N_16518,N_16549);
and U16784 (N_16784,N_16536,N_16437);
nor U16785 (N_16785,N_16455,N_16572);
nor U16786 (N_16786,N_16498,N_16527);
nor U16787 (N_16787,N_16434,N_16403);
and U16788 (N_16788,N_16496,N_16433);
nor U16789 (N_16789,N_16443,N_16460);
xor U16790 (N_16790,N_16550,N_16418);
xor U16791 (N_16791,N_16591,N_16500);
xnor U16792 (N_16792,N_16411,N_16536);
or U16793 (N_16793,N_16436,N_16449);
and U16794 (N_16794,N_16511,N_16464);
or U16795 (N_16795,N_16516,N_16486);
xor U16796 (N_16796,N_16457,N_16445);
nand U16797 (N_16797,N_16525,N_16430);
nor U16798 (N_16798,N_16445,N_16474);
nor U16799 (N_16799,N_16519,N_16495);
nand U16800 (N_16800,N_16798,N_16727);
nor U16801 (N_16801,N_16690,N_16643);
or U16802 (N_16802,N_16601,N_16788);
xnor U16803 (N_16803,N_16617,N_16696);
nor U16804 (N_16804,N_16740,N_16768);
and U16805 (N_16805,N_16650,N_16634);
nand U16806 (N_16806,N_16778,N_16691);
xor U16807 (N_16807,N_16780,N_16717);
xor U16808 (N_16808,N_16793,N_16746);
nand U16809 (N_16809,N_16797,N_16687);
or U16810 (N_16810,N_16639,N_16608);
or U16811 (N_16811,N_16708,N_16674);
nor U16812 (N_16812,N_16737,N_16695);
nand U16813 (N_16813,N_16733,N_16613);
or U16814 (N_16814,N_16722,N_16711);
nand U16815 (N_16815,N_16720,N_16747);
nor U16816 (N_16816,N_16671,N_16624);
nand U16817 (N_16817,N_16610,N_16673);
nor U16818 (N_16818,N_16661,N_16680);
or U16819 (N_16819,N_16623,N_16799);
nor U16820 (N_16820,N_16700,N_16646);
xor U16821 (N_16821,N_16606,N_16714);
or U16822 (N_16822,N_16692,N_16609);
or U16823 (N_16823,N_16640,N_16642);
and U16824 (N_16824,N_16775,N_16723);
xor U16825 (N_16825,N_16618,N_16677);
xor U16826 (N_16826,N_16704,N_16686);
nand U16827 (N_16827,N_16731,N_16754);
and U16828 (N_16828,N_16653,N_16765);
nand U16829 (N_16829,N_16785,N_16626);
nor U16830 (N_16830,N_16666,N_16726);
nand U16831 (N_16831,N_16651,N_16647);
xnor U16832 (N_16832,N_16749,N_16752);
and U16833 (N_16833,N_16628,N_16763);
and U16834 (N_16834,N_16667,N_16648);
or U16835 (N_16835,N_16706,N_16622);
xor U16836 (N_16836,N_16777,N_16629);
nor U16837 (N_16837,N_16762,N_16728);
nor U16838 (N_16838,N_16770,N_16794);
nand U16839 (N_16839,N_16619,N_16683);
or U16840 (N_16840,N_16758,N_16791);
and U16841 (N_16841,N_16774,N_16644);
xor U16842 (N_16842,N_16718,N_16753);
nor U16843 (N_16843,N_16668,N_16678);
nand U16844 (N_16844,N_16605,N_16709);
and U16845 (N_16845,N_16724,N_16741);
nand U16846 (N_16846,N_16730,N_16681);
nor U16847 (N_16847,N_16755,N_16764);
nor U16848 (N_16848,N_16672,N_16664);
nor U16849 (N_16849,N_16790,N_16638);
nor U16850 (N_16850,N_16734,N_16698);
nor U16851 (N_16851,N_16669,N_16693);
xnor U16852 (N_16852,N_16748,N_16710);
or U16853 (N_16853,N_16766,N_16782);
nor U16854 (N_16854,N_16614,N_16676);
xor U16855 (N_16855,N_16738,N_16776);
and U16856 (N_16856,N_16659,N_16627);
xnor U16857 (N_16857,N_16652,N_16633);
or U16858 (N_16858,N_16771,N_16649);
or U16859 (N_16859,N_16773,N_16611);
or U16860 (N_16860,N_16707,N_16732);
nor U16861 (N_16861,N_16725,N_16744);
nand U16862 (N_16862,N_16645,N_16607);
xnor U16863 (N_16863,N_16625,N_16615);
or U16864 (N_16864,N_16654,N_16689);
nand U16865 (N_16865,N_16713,N_16787);
or U16866 (N_16866,N_16760,N_16739);
or U16867 (N_16867,N_16742,N_16719);
nand U16868 (N_16868,N_16701,N_16796);
nor U16869 (N_16869,N_16602,N_16757);
nor U16870 (N_16870,N_16702,N_16662);
or U16871 (N_16871,N_16703,N_16759);
nor U16872 (N_16872,N_16715,N_16616);
or U16873 (N_16873,N_16637,N_16721);
xnor U16874 (N_16874,N_16743,N_16631);
nor U16875 (N_16875,N_16621,N_16665);
xnor U16876 (N_16876,N_16761,N_16751);
and U16877 (N_16877,N_16736,N_16660);
and U16878 (N_16878,N_16767,N_16769);
xor U16879 (N_16879,N_16656,N_16735);
nor U16880 (N_16880,N_16783,N_16675);
and U16881 (N_16881,N_16685,N_16779);
xor U16882 (N_16882,N_16657,N_16786);
and U16883 (N_16883,N_16620,N_16635);
nor U16884 (N_16884,N_16603,N_16772);
nor U16885 (N_16885,N_16682,N_16694);
or U16886 (N_16886,N_16636,N_16756);
or U16887 (N_16887,N_16699,N_16655);
nor U16888 (N_16888,N_16705,N_16641);
nor U16889 (N_16889,N_16745,N_16604);
xnor U16890 (N_16890,N_16729,N_16658);
nand U16891 (N_16891,N_16663,N_16600);
xnor U16892 (N_16892,N_16716,N_16792);
xor U16893 (N_16893,N_16795,N_16630);
nor U16894 (N_16894,N_16784,N_16750);
xor U16895 (N_16895,N_16789,N_16612);
nor U16896 (N_16896,N_16670,N_16781);
nor U16897 (N_16897,N_16697,N_16688);
xnor U16898 (N_16898,N_16679,N_16632);
xor U16899 (N_16899,N_16684,N_16712);
and U16900 (N_16900,N_16661,N_16759);
nand U16901 (N_16901,N_16702,N_16744);
and U16902 (N_16902,N_16776,N_16614);
nand U16903 (N_16903,N_16614,N_16662);
nor U16904 (N_16904,N_16774,N_16790);
xnor U16905 (N_16905,N_16722,N_16611);
xnor U16906 (N_16906,N_16708,N_16626);
or U16907 (N_16907,N_16687,N_16741);
and U16908 (N_16908,N_16657,N_16676);
nor U16909 (N_16909,N_16705,N_16730);
xnor U16910 (N_16910,N_16662,N_16732);
xnor U16911 (N_16911,N_16726,N_16651);
nand U16912 (N_16912,N_16637,N_16681);
nand U16913 (N_16913,N_16753,N_16686);
xor U16914 (N_16914,N_16716,N_16730);
and U16915 (N_16915,N_16716,N_16751);
or U16916 (N_16916,N_16627,N_16680);
nor U16917 (N_16917,N_16781,N_16692);
xor U16918 (N_16918,N_16716,N_16609);
nor U16919 (N_16919,N_16655,N_16697);
and U16920 (N_16920,N_16732,N_16631);
nor U16921 (N_16921,N_16653,N_16641);
xnor U16922 (N_16922,N_16619,N_16687);
nand U16923 (N_16923,N_16663,N_16623);
nand U16924 (N_16924,N_16646,N_16620);
or U16925 (N_16925,N_16670,N_16677);
xnor U16926 (N_16926,N_16692,N_16770);
nand U16927 (N_16927,N_16699,N_16640);
nand U16928 (N_16928,N_16686,N_16609);
and U16929 (N_16929,N_16757,N_16758);
nor U16930 (N_16930,N_16601,N_16656);
or U16931 (N_16931,N_16780,N_16673);
nand U16932 (N_16932,N_16656,N_16774);
nor U16933 (N_16933,N_16647,N_16637);
nor U16934 (N_16934,N_16759,N_16708);
xnor U16935 (N_16935,N_16613,N_16791);
nand U16936 (N_16936,N_16725,N_16740);
and U16937 (N_16937,N_16719,N_16630);
xnor U16938 (N_16938,N_16746,N_16731);
and U16939 (N_16939,N_16650,N_16733);
or U16940 (N_16940,N_16756,N_16644);
nor U16941 (N_16941,N_16620,N_16789);
xor U16942 (N_16942,N_16614,N_16642);
nand U16943 (N_16943,N_16791,N_16636);
nand U16944 (N_16944,N_16657,N_16604);
or U16945 (N_16945,N_16701,N_16712);
nor U16946 (N_16946,N_16614,N_16611);
xnor U16947 (N_16947,N_16721,N_16758);
and U16948 (N_16948,N_16685,N_16787);
nand U16949 (N_16949,N_16721,N_16791);
or U16950 (N_16950,N_16762,N_16793);
nand U16951 (N_16951,N_16765,N_16718);
nand U16952 (N_16952,N_16605,N_16783);
and U16953 (N_16953,N_16742,N_16695);
xor U16954 (N_16954,N_16715,N_16669);
xor U16955 (N_16955,N_16605,N_16774);
xnor U16956 (N_16956,N_16736,N_16664);
nor U16957 (N_16957,N_16642,N_16776);
or U16958 (N_16958,N_16768,N_16775);
or U16959 (N_16959,N_16732,N_16773);
nand U16960 (N_16960,N_16744,N_16692);
nor U16961 (N_16961,N_16621,N_16611);
and U16962 (N_16962,N_16655,N_16772);
nor U16963 (N_16963,N_16756,N_16624);
nand U16964 (N_16964,N_16784,N_16740);
or U16965 (N_16965,N_16723,N_16707);
nand U16966 (N_16966,N_16701,N_16771);
nand U16967 (N_16967,N_16787,N_16640);
nand U16968 (N_16968,N_16694,N_16662);
xnor U16969 (N_16969,N_16709,N_16750);
or U16970 (N_16970,N_16735,N_16628);
and U16971 (N_16971,N_16709,N_16639);
or U16972 (N_16972,N_16724,N_16768);
xor U16973 (N_16973,N_16668,N_16777);
or U16974 (N_16974,N_16737,N_16633);
nand U16975 (N_16975,N_16633,N_16654);
or U16976 (N_16976,N_16643,N_16713);
nor U16977 (N_16977,N_16649,N_16720);
xnor U16978 (N_16978,N_16670,N_16775);
nand U16979 (N_16979,N_16634,N_16645);
nor U16980 (N_16980,N_16672,N_16700);
xor U16981 (N_16981,N_16767,N_16711);
nor U16982 (N_16982,N_16618,N_16626);
and U16983 (N_16983,N_16746,N_16718);
xor U16984 (N_16984,N_16705,N_16648);
and U16985 (N_16985,N_16751,N_16726);
or U16986 (N_16986,N_16759,N_16717);
nor U16987 (N_16987,N_16641,N_16750);
and U16988 (N_16988,N_16722,N_16736);
and U16989 (N_16989,N_16680,N_16667);
nand U16990 (N_16990,N_16641,N_16637);
xnor U16991 (N_16991,N_16719,N_16694);
nand U16992 (N_16992,N_16663,N_16607);
or U16993 (N_16993,N_16758,N_16764);
or U16994 (N_16994,N_16791,N_16733);
or U16995 (N_16995,N_16748,N_16758);
and U16996 (N_16996,N_16749,N_16610);
nand U16997 (N_16997,N_16778,N_16792);
and U16998 (N_16998,N_16728,N_16662);
or U16999 (N_16999,N_16620,N_16679);
or U17000 (N_17000,N_16817,N_16806);
or U17001 (N_17001,N_16950,N_16876);
and U17002 (N_17002,N_16991,N_16915);
or U17003 (N_17003,N_16814,N_16914);
xor U17004 (N_17004,N_16923,N_16829);
xor U17005 (N_17005,N_16909,N_16944);
and U17006 (N_17006,N_16938,N_16962);
nor U17007 (N_17007,N_16896,N_16833);
and U17008 (N_17008,N_16828,N_16847);
nand U17009 (N_17009,N_16903,N_16910);
and U17010 (N_17010,N_16984,N_16993);
or U17011 (N_17011,N_16958,N_16924);
or U17012 (N_17012,N_16873,N_16827);
xor U17013 (N_17013,N_16875,N_16839);
nand U17014 (N_17014,N_16865,N_16819);
or U17015 (N_17015,N_16888,N_16826);
or U17016 (N_17016,N_16967,N_16853);
or U17017 (N_17017,N_16862,N_16840);
xnor U17018 (N_17018,N_16927,N_16882);
xor U17019 (N_17019,N_16985,N_16831);
and U17020 (N_17020,N_16990,N_16821);
nand U17021 (N_17021,N_16845,N_16884);
and U17022 (N_17022,N_16911,N_16897);
nor U17023 (N_17023,N_16982,N_16926);
or U17024 (N_17024,N_16930,N_16918);
xor U17025 (N_17025,N_16912,N_16932);
or U17026 (N_17026,N_16994,N_16964);
nor U17027 (N_17027,N_16823,N_16913);
and U17028 (N_17028,N_16928,N_16816);
or U17029 (N_17029,N_16992,N_16843);
and U17030 (N_17030,N_16906,N_16988);
and U17031 (N_17031,N_16802,N_16830);
nor U17032 (N_17032,N_16810,N_16883);
nand U17033 (N_17033,N_16997,N_16933);
xor U17034 (N_17034,N_16860,N_16822);
nand U17035 (N_17035,N_16968,N_16981);
nor U17036 (N_17036,N_16919,N_16902);
and U17037 (N_17037,N_16866,N_16809);
and U17038 (N_17038,N_16979,N_16801);
or U17039 (N_17039,N_16940,N_16942);
xor U17040 (N_17040,N_16920,N_16959);
and U17041 (N_17041,N_16807,N_16929);
and U17042 (N_17042,N_16879,N_16935);
nand U17043 (N_17043,N_16948,N_16945);
nor U17044 (N_17044,N_16877,N_16846);
or U17045 (N_17045,N_16832,N_16811);
or U17046 (N_17046,N_16841,N_16898);
nor U17047 (N_17047,N_16998,N_16859);
and U17048 (N_17048,N_16978,N_16961);
nand U17049 (N_17049,N_16863,N_16867);
and U17050 (N_17050,N_16868,N_16854);
xnor U17051 (N_17051,N_16901,N_16999);
nand U17052 (N_17052,N_16818,N_16971);
or U17053 (N_17053,N_16989,N_16842);
xor U17054 (N_17054,N_16825,N_16889);
and U17055 (N_17055,N_16983,N_16916);
nand U17056 (N_17056,N_16857,N_16917);
or U17057 (N_17057,N_16960,N_16872);
or U17058 (N_17058,N_16874,N_16943);
or U17059 (N_17059,N_16800,N_16925);
xor U17060 (N_17060,N_16815,N_16931);
xor U17061 (N_17061,N_16895,N_16974);
nor U17062 (N_17062,N_16855,N_16891);
or U17063 (N_17063,N_16837,N_16892);
nor U17064 (N_17064,N_16952,N_16951);
or U17065 (N_17065,N_16856,N_16835);
or U17066 (N_17066,N_16805,N_16957);
nand U17067 (N_17067,N_16954,N_16880);
and U17068 (N_17068,N_16849,N_16834);
or U17069 (N_17069,N_16864,N_16858);
xnor U17070 (N_17070,N_16976,N_16852);
nand U17071 (N_17071,N_16899,N_16808);
nand U17072 (N_17072,N_16969,N_16995);
xnor U17073 (N_17073,N_16836,N_16956);
and U17074 (N_17074,N_16812,N_16813);
or U17075 (N_17075,N_16986,N_16949);
nand U17076 (N_17076,N_16922,N_16886);
xnor U17077 (N_17077,N_16838,N_16861);
and U17078 (N_17078,N_16881,N_16975);
xor U17079 (N_17079,N_16851,N_16885);
or U17080 (N_17080,N_16871,N_16820);
nand U17081 (N_17081,N_16996,N_16947);
or U17082 (N_17082,N_16887,N_16904);
and U17083 (N_17083,N_16905,N_16804);
xor U17084 (N_17084,N_16946,N_16921);
nand U17085 (N_17085,N_16850,N_16900);
nand U17086 (N_17086,N_16894,N_16907);
nor U17087 (N_17087,N_16980,N_16941);
xnor U17088 (N_17088,N_16934,N_16977);
xor U17089 (N_17089,N_16878,N_16803);
xnor U17090 (N_17090,N_16955,N_16953);
or U17091 (N_17091,N_16893,N_16970);
nor U17092 (N_17092,N_16848,N_16939);
nand U17093 (N_17093,N_16963,N_16973);
or U17094 (N_17094,N_16890,N_16869);
nand U17095 (N_17095,N_16972,N_16824);
nor U17096 (N_17096,N_16844,N_16987);
xor U17097 (N_17097,N_16870,N_16965);
nor U17098 (N_17098,N_16908,N_16937);
xor U17099 (N_17099,N_16966,N_16936);
or U17100 (N_17100,N_16814,N_16932);
nor U17101 (N_17101,N_16950,N_16895);
and U17102 (N_17102,N_16853,N_16986);
nand U17103 (N_17103,N_16809,N_16916);
or U17104 (N_17104,N_16964,N_16835);
xnor U17105 (N_17105,N_16879,N_16896);
and U17106 (N_17106,N_16972,N_16874);
xor U17107 (N_17107,N_16833,N_16883);
and U17108 (N_17108,N_16971,N_16906);
nand U17109 (N_17109,N_16874,N_16928);
or U17110 (N_17110,N_16850,N_16819);
nor U17111 (N_17111,N_16874,N_16933);
nand U17112 (N_17112,N_16965,N_16921);
or U17113 (N_17113,N_16816,N_16877);
nor U17114 (N_17114,N_16895,N_16880);
xor U17115 (N_17115,N_16867,N_16928);
xor U17116 (N_17116,N_16827,N_16960);
nor U17117 (N_17117,N_16904,N_16924);
or U17118 (N_17118,N_16930,N_16826);
nor U17119 (N_17119,N_16820,N_16850);
or U17120 (N_17120,N_16891,N_16979);
nand U17121 (N_17121,N_16861,N_16898);
or U17122 (N_17122,N_16941,N_16854);
and U17123 (N_17123,N_16805,N_16929);
xor U17124 (N_17124,N_16961,N_16875);
nand U17125 (N_17125,N_16817,N_16966);
nand U17126 (N_17126,N_16810,N_16897);
or U17127 (N_17127,N_16958,N_16997);
xor U17128 (N_17128,N_16805,N_16944);
or U17129 (N_17129,N_16810,N_16949);
nor U17130 (N_17130,N_16906,N_16969);
nor U17131 (N_17131,N_16924,N_16944);
nor U17132 (N_17132,N_16870,N_16923);
or U17133 (N_17133,N_16968,N_16894);
nor U17134 (N_17134,N_16923,N_16876);
nand U17135 (N_17135,N_16824,N_16881);
nand U17136 (N_17136,N_16931,N_16849);
or U17137 (N_17137,N_16898,N_16813);
nor U17138 (N_17138,N_16909,N_16999);
or U17139 (N_17139,N_16977,N_16886);
xor U17140 (N_17140,N_16888,N_16818);
and U17141 (N_17141,N_16907,N_16948);
xnor U17142 (N_17142,N_16837,N_16820);
nor U17143 (N_17143,N_16890,N_16910);
nor U17144 (N_17144,N_16806,N_16893);
and U17145 (N_17145,N_16993,N_16975);
xnor U17146 (N_17146,N_16830,N_16978);
nor U17147 (N_17147,N_16986,N_16822);
xnor U17148 (N_17148,N_16887,N_16818);
and U17149 (N_17149,N_16934,N_16874);
nand U17150 (N_17150,N_16934,N_16844);
or U17151 (N_17151,N_16851,N_16881);
and U17152 (N_17152,N_16806,N_16975);
and U17153 (N_17153,N_16975,N_16898);
nand U17154 (N_17154,N_16975,N_16836);
nor U17155 (N_17155,N_16999,N_16852);
xnor U17156 (N_17156,N_16974,N_16921);
nor U17157 (N_17157,N_16827,N_16938);
and U17158 (N_17158,N_16927,N_16895);
nor U17159 (N_17159,N_16823,N_16849);
xnor U17160 (N_17160,N_16833,N_16902);
nand U17161 (N_17161,N_16903,N_16940);
or U17162 (N_17162,N_16990,N_16862);
or U17163 (N_17163,N_16961,N_16889);
xnor U17164 (N_17164,N_16977,N_16935);
and U17165 (N_17165,N_16957,N_16934);
xor U17166 (N_17166,N_16938,N_16845);
nor U17167 (N_17167,N_16995,N_16939);
xor U17168 (N_17168,N_16891,N_16936);
nand U17169 (N_17169,N_16996,N_16870);
and U17170 (N_17170,N_16833,N_16948);
or U17171 (N_17171,N_16873,N_16863);
nor U17172 (N_17172,N_16900,N_16916);
or U17173 (N_17173,N_16920,N_16834);
or U17174 (N_17174,N_16902,N_16907);
or U17175 (N_17175,N_16859,N_16962);
and U17176 (N_17176,N_16824,N_16982);
nor U17177 (N_17177,N_16871,N_16934);
nand U17178 (N_17178,N_16958,N_16886);
xnor U17179 (N_17179,N_16867,N_16890);
or U17180 (N_17180,N_16865,N_16915);
nor U17181 (N_17181,N_16802,N_16800);
xor U17182 (N_17182,N_16885,N_16915);
or U17183 (N_17183,N_16856,N_16875);
nor U17184 (N_17184,N_16893,N_16867);
or U17185 (N_17185,N_16933,N_16876);
and U17186 (N_17186,N_16912,N_16937);
and U17187 (N_17187,N_16854,N_16802);
nand U17188 (N_17188,N_16865,N_16855);
or U17189 (N_17189,N_16966,N_16941);
or U17190 (N_17190,N_16954,N_16998);
and U17191 (N_17191,N_16896,N_16843);
xor U17192 (N_17192,N_16977,N_16975);
or U17193 (N_17193,N_16826,N_16849);
or U17194 (N_17194,N_16973,N_16939);
or U17195 (N_17195,N_16996,N_16953);
and U17196 (N_17196,N_16897,N_16872);
and U17197 (N_17197,N_16916,N_16852);
and U17198 (N_17198,N_16843,N_16832);
xnor U17199 (N_17199,N_16981,N_16876);
and U17200 (N_17200,N_17040,N_17058);
xnor U17201 (N_17201,N_17027,N_17000);
and U17202 (N_17202,N_17089,N_17032);
nor U17203 (N_17203,N_17025,N_17116);
nand U17204 (N_17204,N_17043,N_17097);
xor U17205 (N_17205,N_17086,N_17037);
or U17206 (N_17206,N_17149,N_17185);
xor U17207 (N_17207,N_17019,N_17077);
and U17208 (N_17208,N_17134,N_17189);
or U17209 (N_17209,N_17157,N_17059);
xnor U17210 (N_17210,N_17009,N_17052);
xnor U17211 (N_17211,N_17156,N_17187);
nor U17212 (N_17212,N_17140,N_17135);
or U17213 (N_17213,N_17041,N_17030);
or U17214 (N_17214,N_17055,N_17186);
nand U17215 (N_17215,N_17083,N_17144);
xnor U17216 (N_17216,N_17068,N_17105);
nand U17217 (N_17217,N_17170,N_17125);
xor U17218 (N_17218,N_17153,N_17173);
and U17219 (N_17219,N_17106,N_17117);
xnor U17220 (N_17220,N_17123,N_17179);
and U17221 (N_17221,N_17092,N_17014);
or U17222 (N_17222,N_17182,N_17151);
or U17223 (N_17223,N_17063,N_17064);
and U17224 (N_17224,N_17061,N_17191);
or U17225 (N_17225,N_17109,N_17008);
nor U17226 (N_17226,N_17172,N_17017);
nand U17227 (N_17227,N_17071,N_17120);
nand U17228 (N_17228,N_17127,N_17056);
or U17229 (N_17229,N_17142,N_17108);
xor U17230 (N_17230,N_17107,N_17021);
nor U17231 (N_17231,N_17033,N_17079);
or U17232 (N_17232,N_17137,N_17065);
and U17233 (N_17233,N_17168,N_17048);
and U17234 (N_17234,N_17088,N_17198);
and U17235 (N_17235,N_17013,N_17139);
nor U17236 (N_17236,N_17152,N_17023);
nor U17237 (N_17237,N_17118,N_17146);
xor U17238 (N_17238,N_17007,N_17085);
xor U17239 (N_17239,N_17073,N_17148);
nor U17240 (N_17240,N_17110,N_17184);
nand U17241 (N_17241,N_17130,N_17102);
nor U17242 (N_17242,N_17093,N_17199);
nand U17243 (N_17243,N_17035,N_17003);
xnor U17244 (N_17244,N_17101,N_17046);
nor U17245 (N_17245,N_17129,N_17180);
nor U17246 (N_17246,N_17006,N_17181);
nand U17247 (N_17247,N_17169,N_17070);
xnor U17248 (N_17248,N_17190,N_17047);
nand U17249 (N_17249,N_17174,N_17154);
or U17250 (N_17250,N_17002,N_17038);
nor U17251 (N_17251,N_17018,N_17178);
nor U17252 (N_17252,N_17094,N_17166);
nor U17253 (N_17253,N_17004,N_17145);
nor U17254 (N_17254,N_17016,N_17143);
or U17255 (N_17255,N_17119,N_17076);
nand U17256 (N_17256,N_17060,N_17162);
nand U17257 (N_17257,N_17044,N_17112);
nor U17258 (N_17258,N_17126,N_17104);
nor U17259 (N_17259,N_17141,N_17010);
and U17260 (N_17260,N_17133,N_17028);
nor U17261 (N_17261,N_17005,N_17163);
and U17262 (N_17262,N_17087,N_17057);
nor U17263 (N_17263,N_17171,N_17165);
nor U17264 (N_17264,N_17113,N_17012);
nand U17265 (N_17265,N_17159,N_17195);
xor U17266 (N_17266,N_17011,N_17082);
nand U17267 (N_17267,N_17015,N_17081);
nand U17268 (N_17268,N_17196,N_17136);
nor U17269 (N_17269,N_17069,N_17177);
nor U17270 (N_17270,N_17124,N_17050);
or U17271 (N_17271,N_17193,N_17051);
and U17272 (N_17272,N_17099,N_17020);
or U17273 (N_17273,N_17078,N_17036);
or U17274 (N_17274,N_17183,N_17026);
nor U17275 (N_17275,N_17155,N_17049);
nor U17276 (N_17276,N_17175,N_17034);
nand U17277 (N_17277,N_17098,N_17084);
and U17278 (N_17278,N_17128,N_17054);
and U17279 (N_17279,N_17100,N_17031);
or U17280 (N_17280,N_17121,N_17192);
or U17281 (N_17281,N_17045,N_17067);
nor U17282 (N_17282,N_17080,N_17167);
nor U17283 (N_17283,N_17158,N_17160);
nand U17284 (N_17284,N_17066,N_17095);
and U17285 (N_17285,N_17062,N_17114);
xor U17286 (N_17286,N_17022,N_17150);
xor U17287 (N_17287,N_17024,N_17194);
nor U17288 (N_17288,N_17138,N_17115);
and U17289 (N_17289,N_17053,N_17132);
xnor U17290 (N_17290,N_17096,N_17197);
xor U17291 (N_17291,N_17039,N_17042);
nor U17292 (N_17292,N_17147,N_17074);
and U17293 (N_17293,N_17001,N_17176);
xor U17294 (N_17294,N_17090,N_17075);
xnor U17295 (N_17295,N_17131,N_17091);
or U17296 (N_17296,N_17161,N_17122);
nor U17297 (N_17297,N_17164,N_17103);
or U17298 (N_17298,N_17029,N_17072);
nand U17299 (N_17299,N_17111,N_17188);
and U17300 (N_17300,N_17139,N_17048);
nor U17301 (N_17301,N_17009,N_17059);
or U17302 (N_17302,N_17174,N_17008);
nor U17303 (N_17303,N_17041,N_17039);
and U17304 (N_17304,N_17096,N_17091);
or U17305 (N_17305,N_17010,N_17069);
nand U17306 (N_17306,N_17127,N_17152);
nor U17307 (N_17307,N_17071,N_17059);
or U17308 (N_17308,N_17103,N_17020);
and U17309 (N_17309,N_17169,N_17135);
and U17310 (N_17310,N_17178,N_17122);
nor U17311 (N_17311,N_17150,N_17161);
xor U17312 (N_17312,N_17122,N_17163);
nor U17313 (N_17313,N_17150,N_17038);
xor U17314 (N_17314,N_17098,N_17021);
nand U17315 (N_17315,N_17013,N_17044);
and U17316 (N_17316,N_17128,N_17051);
nor U17317 (N_17317,N_17115,N_17087);
nor U17318 (N_17318,N_17162,N_17194);
or U17319 (N_17319,N_17105,N_17169);
nand U17320 (N_17320,N_17031,N_17051);
or U17321 (N_17321,N_17158,N_17037);
nor U17322 (N_17322,N_17068,N_17131);
xnor U17323 (N_17323,N_17045,N_17069);
xor U17324 (N_17324,N_17075,N_17077);
and U17325 (N_17325,N_17087,N_17093);
or U17326 (N_17326,N_17084,N_17022);
nand U17327 (N_17327,N_17009,N_17122);
nand U17328 (N_17328,N_17097,N_17098);
nand U17329 (N_17329,N_17130,N_17192);
or U17330 (N_17330,N_17060,N_17044);
xnor U17331 (N_17331,N_17022,N_17042);
or U17332 (N_17332,N_17191,N_17129);
nor U17333 (N_17333,N_17179,N_17178);
xor U17334 (N_17334,N_17038,N_17069);
nand U17335 (N_17335,N_17054,N_17040);
and U17336 (N_17336,N_17022,N_17128);
nand U17337 (N_17337,N_17099,N_17159);
nand U17338 (N_17338,N_17014,N_17164);
xnor U17339 (N_17339,N_17126,N_17131);
xor U17340 (N_17340,N_17095,N_17155);
nor U17341 (N_17341,N_17009,N_17145);
and U17342 (N_17342,N_17021,N_17195);
nand U17343 (N_17343,N_17035,N_17053);
xor U17344 (N_17344,N_17088,N_17146);
nand U17345 (N_17345,N_17129,N_17045);
or U17346 (N_17346,N_17125,N_17104);
and U17347 (N_17347,N_17164,N_17128);
xor U17348 (N_17348,N_17090,N_17179);
and U17349 (N_17349,N_17151,N_17030);
xor U17350 (N_17350,N_17177,N_17168);
or U17351 (N_17351,N_17160,N_17009);
or U17352 (N_17352,N_17153,N_17023);
nor U17353 (N_17353,N_17040,N_17174);
xnor U17354 (N_17354,N_17169,N_17177);
nor U17355 (N_17355,N_17057,N_17133);
nor U17356 (N_17356,N_17080,N_17000);
xnor U17357 (N_17357,N_17165,N_17173);
or U17358 (N_17358,N_17161,N_17073);
nand U17359 (N_17359,N_17022,N_17155);
xor U17360 (N_17360,N_17082,N_17166);
or U17361 (N_17361,N_17100,N_17138);
xor U17362 (N_17362,N_17181,N_17007);
nand U17363 (N_17363,N_17015,N_17089);
nor U17364 (N_17364,N_17168,N_17146);
xnor U17365 (N_17365,N_17106,N_17083);
and U17366 (N_17366,N_17125,N_17070);
or U17367 (N_17367,N_17010,N_17133);
nor U17368 (N_17368,N_17161,N_17025);
or U17369 (N_17369,N_17016,N_17115);
xor U17370 (N_17370,N_17165,N_17019);
nor U17371 (N_17371,N_17097,N_17085);
or U17372 (N_17372,N_17027,N_17186);
xnor U17373 (N_17373,N_17053,N_17011);
or U17374 (N_17374,N_17186,N_17103);
nand U17375 (N_17375,N_17173,N_17111);
nor U17376 (N_17376,N_17059,N_17077);
nand U17377 (N_17377,N_17165,N_17031);
and U17378 (N_17378,N_17120,N_17082);
xnor U17379 (N_17379,N_17188,N_17079);
or U17380 (N_17380,N_17055,N_17022);
or U17381 (N_17381,N_17027,N_17189);
and U17382 (N_17382,N_17003,N_17026);
nor U17383 (N_17383,N_17070,N_17177);
nor U17384 (N_17384,N_17013,N_17116);
or U17385 (N_17385,N_17072,N_17160);
nand U17386 (N_17386,N_17084,N_17081);
and U17387 (N_17387,N_17040,N_17132);
nand U17388 (N_17388,N_17165,N_17085);
nor U17389 (N_17389,N_17147,N_17116);
and U17390 (N_17390,N_17091,N_17153);
or U17391 (N_17391,N_17025,N_17194);
nand U17392 (N_17392,N_17147,N_17056);
xor U17393 (N_17393,N_17140,N_17074);
nand U17394 (N_17394,N_17034,N_17179);
or U17395 (N_17395,N_17072,N_17182);
xnor U17396 (N_17396,N_17082,N_17096);
xnor U17397 (N_17397,N_17067,N_17061);
and U17398 (N_17398,N_17072,N_17104);
xnor U17399 (N_17399,N_17032,N_17144);
nor U17400 (N_17400,N_17212,N_17391);
nand U17401 (N_17401,N_17382,N_17265);
nor U17402 (N_17402,N_17210,N_17291);
nand U17403 (N_17403,N_17348,N_17344);
nand U17404 (N_17404,N_17211,N_17328);
or U17405 (N_17405,N_17274,N_17288);
and U17406 (N_17406,N_17377,N_17280);
nand U17407 (N_17407,N_17335,N_17392);
nand U17408 (N_17408,N_17366,N_17379);
or U17409 (N_17409,N_17236,N_17368);
and U17410 (N_17410,N_17287,N_17258);
xnor U17411 (N_17411,N_17246,N_17385);
nor U17412 (N_17412,N_17389,N_17352);
xor U17413 (N_17413,N_17360,N_17203);
xnor U17414 (N_17414,N_17397,N_17256);
and U17415 (N_17415,N_17329,N_17311);
or U17416 (N_17416,N_17342,N_17350);
nand U17417 (N_17417,N_17234,N_17270);
and U17418 (N_17418,N_17355,N_17218);
nand U17419 (N_17419,N_17354,N_17373);
or U17420 (N_17420,N_17371,N_17240);
and U17421 (N_17421,N_17244,N_17302);
nand U17422 (N_17422,N_17387,N_17297);
nor U17423 (N_17423,N_17241,N_17305);
nor U17424 (N_17424,N_17278,N_17320);
xnor U17425 (N_17425,N_17266,N_17245);
nor U17426 (N_17426,N_17393,N_17358);
and U17427 (N_17427,N_17248,N_17318);
xnor U17428 (N_17428,N_17359,N_17390);
nand U17429 (N_17429,N_17296,N_17381);
or U17430 (N_17430,N_17252,N_17281);
xor U17431 (N_17431,N_17238,N_17298);
xor U17432 (N_17432,N_17243,N_17294);
and U17433 (N_17433,N_17289,N_17314);
and U17434 (N_17434,N_17331,N_17208);
nor U17435 (N_17435,N_17399,N_17227);
nor U17436 (N_17436,N_17233,N_17217);
nand U17437 (N_17437,N_17398,N_17362);
or U17438 (N_17438,N_17306,N_17250);
nand U17439 (N_17439,N_17273,N_17339);
nand U17440 (N_17440,N_17378,N_17285);
xnor U17441 (N_17441,N_17284,N_17215);
xor U17442 (N_17442,N_17300,N_17223);
and U17443 (N_17443,N_17376,N_17200);
and U17444 (N_17444,N_17259,N_17263);
or U17445 (N_17445,N_17361,N_17315);
nor U17446 (N_17446,N_17386,N_17347);
and U17447 (N_17447,N_17365,N_17260);
nand U17448 (N_17448,N_17257,N_17202);
or U17449 (N_17449,N_17269,N_17303);
nand U17450 (N_17450,N_17367,N_17224);
and U17451 (N_17451,N_17345,N_17374);
xnor U17452 (N_17452,N_17220,N_17316);
and U17453 (N_17453,N_17254,N_17231);
or U17454 (N_17454,N_17372,N_17356);
and U17455 (N_17455,N_17299,N_17321);
xor U17456 (N_17456,N_17225,N_17222);
nand U17457 (N_17457,N_17255,N_17226);
nor U17458 (N_17458,N_17330,N_17332);
or U17459 (N_17459,N_17308,N_17313);
nand U17460 (N_17460,N_17346,N_17395);
and U17461 (N_17461,N_17207,N_17249);
and U17462 (N_17462,N_17276,N_17295);
nor U17463 (N_17463,N_17232,N_17323);
nor U17464 (N_17464,N_17214,N_17349);
or U17465 (N_17465,N_17307,N_17264);
xnor U17466 (N_17466,N_17267,N_17219);
nor U17467 (N_17467,N_17262,N_17221);
nor U17468 (N_17468,N_17235,N_17340);
and U17469 (N_17469,N_17351,N_17279);
and U17470 (N_17470,N_17353,N_17333);
xnor U17471 (N_17471,N_17237,N_17357);
or U17472 (N_17472,N_17216,N_17268);
xor U17473 (N_17473,N_17292,N_17201);
and U17474 (N_17474,N_17326,N_17228);
nor U17475 (N_17475,N_17204,N_17230);
nand U17476 (N_17476,N_17325,N_17336);
nand U17477 (N_17477,N_17290,N_17363);
xnor U17478 (N_17478,N_17205,N_17277);
and U17479 (N_17479,N_17209,N_17301);
and U17480 (N_17480,N_17338,N_17370);
nand U17481 (N_17481,N_17239,N_17380);
nand U17482 (N_17482,N_17213,N_17327);
and U17483 (N_17483,N_17322,N_17261);
nand U17484 (N_17484,N_17242,N_17251);
xor U17485 (N_17485,N_17304,N_17229);
or U17486 (N_17486,N_17319,N_17369);
or U17487 (N_17487,N_17247,N_17293);
nor U17488 (N_17488,N_17312,N_17283);
or U17489 (N_17489,N_17309,N_17343);
or U17490 (N_17490,N_17388,N_17206);
nand U17491 (N_17491,N_17324,N_17337);
xor U17492 (N_17492,N_17364,N_17341);
xor U17493 (N_17493,N_17271,N_17396);
nand U17494 (N_17494,N_17334,N_17384);
nor U17495 (N_17495,N_17275,N_17272);
or U17496 (N_17496,N_17383,N_17394);
nor U17497 (N_17497,N_17375,N_17310);
and U17498 (N_17498,N_17317,N_17253);
or U17499 (N_17499,N_17286,N_17282);
nor U17500 (N_17500,N_17214,N_17201);
or U17501 (N_17501,N_17286,N_17398);
xor U17502 (N_17502,N_17343,N_17217);
nor U17503 (N_17503,N_17355,N_17310);
or U17504 (N_17504,N_17338,N_17238);
xor U17505 (N_17505,N_17394,N_17399);
and U17506 (N_17506,N_17245,N_17236);
nand U17507 (N_17507,N_17327,N_17364);
nor U17508 (N_17508,N_17336,N_17382);
nor U17509 (N_17509,N_17243,N_17364);
nand U17510 (N_17510,N_17280,N_17345);
and U17511 (N_17511,N_17222,N_17208);
nor U17512 (N_17512,N_17245,N_17237);
xor U17513 (N_17513,N_17265,N_17218);
and U17514 (N_17514,N_17356,N_17299);
nand U17515 (N_17515,N_17238,N_17356);
nor U17516 (N_17516,N_17337,N_17384);
or U17517 (N_17517,N_17271,N_17234);
nand U17518 (N_17518,N_17326,N_17323);
and U17519 (N_17519,N_17354,N_17324);
nor U17520 (N_17520,N_17359,N_17376);
or U17521 (N_17521,N_17215,N_17226);
nor U17522 (N_17522,N_17361,N_17352);
or U17523 (N_17523,N_17387,N_17247);
xor U17524 (N_17524,N_17296,N_17339);
xnor U17525 (N_17525,N_17216,N_17343);
or U17526 (N_17526,N_17351,N_17360);
and U17527 (N_17527,N_17299,N_17385);
xnor U17528 (N_17528,N_17385,N_17329);
xor U17529 (N_17529,N_17257,N_17329);
and U17530 (N_17530,N_17264,N_17206);
xnor U17531 (N_17531,N_17217,N_17206);
xor U17532 (N_17532,N_17382,N_17345);
nor U17533 (N_17533,N_17365,N_17318);
or U17534 (N_17534,N_17345,N_17275);
nor U17535 (N_17535,N_17224,N_17298);
or U17536 (N_17536,N_17249,N_17385);
or U17537 (N_17537,N_17391,N_17284);
xor U17538 (N_17538,N_17355,N_17350);
xor U17539 (N_17539,N_17308,N_17386);
nor U17540 (N_17540,N_17344,N_17305);
and U17541 (N_17541,N_17322,N_17331);
nor U17542 (N_17542,N_17322,N_17233);
or U17543 (N_17543,N_17352,N_17242);
nand U17544 (N_17544,N_17323,N_17239);
nand U17545 (N_17545,N_17360,N_17309);
nor U17546 (N_17546,N_17338,N_17274);
xor U17547 (N_17547,N_17251,N_17361);
or U17548 (N_17548,N_17229,N_17220);
or U17549 (N_17549,N_17328,N_17368);
and U17550 (N_17550,N_17276,N_17237);
and U17551 (N_17551,N_17360,N_17206);
nor U17552 (N_17552,N_17260,N_17380);
xor U17553 (N_17553,N_17349,N_17208);
xor U17554 (N_17554,N_17288,N_17266);
and U17555 (N_17555,N_17309,N_17247);
nor U17556 (N_17556,N_17307,N_17223);
nand U17557 (N_17557,N_17347,N_17287);
xor U17558 (N_17558,N_17246,N_17247);
xor U17559 (N_17559,N_17284,N_17241);
and U17560 (N_17560,N_17284,N_17205);
or U17561 (N_17561,N_17207,N_17322);
and U17562 (N_17562,N_17286,N_17378);
nand U17563 (N_17563,N_17321,N_17359);
nor U17564 (N_17564,N_17339,N_17226);
or U17565 (N_17565,N_17310,N_17259);
nand U17566 (N_17566,N_17382,N_17251);
xnor U17567 (N_17567,N_17327,N_17302);
and U17568 (N_17568,N_17276,N_17380);
xnor U17569 (N_17569,N_17200,N_17214);
nand U17570 (N_17570,N_17201,N_17350);
xor U17571 (N_17571,N_17298,N_17373);
xnor U17572 (N_17572,N_17222,N_17356);
nand U17573 (N_17573,N_17361,N_17205);
and U17574 (N_17574,N_17233,N_17346);
nor U17575 (N_17575,N_17247,N_17235);
nand U17576 (N_17576,N_17340,N_17387);
or U17577 (N_17577,N_17232,N_17263);
or U17578 (N_17578,N_17368,N_17243);
xnor U17579 (N_17579,N_17382,N_17376);
and U17580 (N_17580,N_17381,N_17240);
xor U17581 (N_17581,N_17266,N_17374);
nor U17582 (N_17582,N_17394,N_17256);
nor U17583 (N_17583,N_17328,N_17294);
and U17584 (N_17584,N_17343,N_17368);
nand U17585 (N_17585,N_17313,N_17298);
and U17586 (N_17586,N_17253,N_17244);
xnor U17587 (N_17587,N_17269,N_17271);
and U17588 (N_17588,N_17342,N_17353);
nor U17589 (N_17589,N_17232,N_17341);
nor U17590 (N_17590,N_17297,N_17285);
nand U17591 (N_17591,N_17279,N_17299);
xor U17592 (N_17592,N_17244,N_17336);
nand U17593 (N_17593,N_17293,N_17383);
and U17594 (N_17594,N_17214,N_17398);
nand U17595 (N_17595,N_17367,N_17336);
xnor U17596 (N_17596,N_17203,N_17357);
xor U17597 (N_17597,N_17261,N_17391);
and U17598 (N_17598,N_17274,N_17231);
nor U17599 (N_17599,N_17389,N_17259);
nor U17600 (N_17600,N_17544,N_17551);
or U17601 (N_17601,N_17558,N_17414);
or U17602 (N_17602,N_17443,N_17451);
nand U17603 (N_17603,N_17432,N_17404);
or U17604 (N_17604,N_17530,N_17526);
and U17605 (N_17605,N_17520,N_17472);
nor U17606 (N_17606,N_17476,N_17435);
nand U17607 (N_17607,N_17517,N_17511);
nor U17608 (N_17608,N_17518,N_17545);
xor U17609 (N_17609,N_17462,N_17563);
xnor U17610 (N_17610,N_17429,N_17521);
xor U17611 (N_17611,N_17473,N_17492);
or U17612 (N_17612,N_17466,N_17585);
nor U17613 (N_17613,N_17495,N_17539);
xnor U17614 (N_17614,N_17457,N_17580);
nand U17615 (N_17615,N_17405,N_17549);
or U17616 (N_17616,N_17550,N_17489);
nand U17617 (N_17617,N_17506,N_17468);
and U17618 (N_17618,N_17562,N_17553);
xnor U17619 (N_17619,N_17433,N_17500);
nor U17620 (N_17620,N_17465,N_17401);
nand U17621 (N_17621,N_17407,N_17477);
nor U17622 (N_17622,N_17437,N_17515);
nand U17623 (N_17623,N_17421,N_17471);
nand U17624 (N_17624,N_17486,N_17430);
nand U17625 (N_17625,N_17535,N_17494);
nand U17626 (N_17626,N_17543,N_17527);
or U17627 (N_17627,N_17469,N_17504);
nand U17628 (N_17628,N_17528,N_17560);
nor U17629 (N_17629,N_17496,N_17408);
or U17630 (N_17630,N_17582,N_17566);
nor U17631 (N_17631,N_17581,N_17485);
nor U17632 (N_17632,N_17482,N_17509);
xnor U17633 (N_17633,N_17596,N_17510);
xor U17634 (N_17634,N_17565,N_17428);
nor U17635 (N_17635,N_17552,N_17592);
and U17636 (N_17636,N_17400,N_17569);
xnor U17637 (N_17637,N_17455,N_17416);
xnor U17638 (N_17638,N_17478,N_17426);
nand U17639 (N_17639,N_17480,N_17519);
xor U17640 (N_17640,N_17556,N_17578);
nand U17641 (N_17641,N_17450,N_17501);
xnor U17642 (N_17642,N_17431,N_17567);
nand U17643 (N_17643,N_17547,N_17570);
nor U17644 (N_17644,N_17591,N_17534);
nor U17645 (N_17645,N_17442,N_17564);
or U17646 (N_17646,N_17475,N_17412);
or U17647 (N_17647,N_17590,N_17419);
nor U17648 (N_17648,N_17554,N_17522);
and U17649 (N_17649,N_17499,N_17409);
nand U17650 (N_17650,N_17542,N_17446);
or U17651 (N_17651,N_17513,N_17548);
and U17652 (N_17652,N_17445,N_17481);
and U17653 (N_17653,N_17597,N_17541);
nor U17654 (N_17654,N_17503,N_17434);
or U17655 (N_17655,N_17454,N_17479);
and U17656 (N_17656,N_17423,N_17448);
nor U17657 (N_17657,N_17557,N_17525);
nand U17658 (N_17658,N_17470,N_17461);
nand U17659 (N_17659,N_17508,N_17577);
nor U17660 (N_17660,N_17595,N_17540);
nand U17661 (N_17661,N_17484,N_17410);
xor U17662 (N_17662,N_17452,N_17536);
or U17663 (N_17663,N_17533,N_17463);
xor U17664 (N_17664,N_17436,N_17574);
nand U17665 (N_17665,N_17420,N_17579);
nand U17666 (N_17666,N_17524,N_17425);
xnor U17667 (N_17667,N_17415,N_17411);
and U17668 (N_17668,N_17444,N_17458);
and U17669 (N_17669,N_17586,N_17439);
xnor U17670 (N_17670,N_17537,N_17474);
nor U17671 (N_17671,N_17529,N_17531);
xnor U17672 (N_17672,N_17402,N_17447);
and U17673 (N_17673,N_17523,N_17424);
and U17674 (N_17674,N_17491,N_17587);
nor U17675 (N_17675,N_17588,N_17546);
nand U17676 (N_17676,N_17573,N_17417);
and U17677 (N_17677,N_17427,N_17413);
or U17678 (N_17678,N_17512,N_17441);
nor U17679 (N_17679,N_17576,N_17490);
nand U17680 (N_17680,N_17505,N_17594);
nor U17681 (N_17681,N_17599,N_17493);
or U17682 (N_17682,N_17575,N_17438);
nand U17683 (N_17683,N_17418,N_17488);
and U17684 (N_17684,N_17403,N_17406);
nand U17685 (N_17685,N_17559,N_17561);
nor U17686 (N_17686,N_17498,N_17514);
or U17687 (N_17687,N_17571,N_17464);
nand U17688 (N_17688,N_17584,N_17568);
nor U17689 (N_17689,N_17456,N_17467);
nor U17690 (N_17690,N_17583,N_17483);
nand U17691 (N_17691,N_17422,N_17459);
or U17692 (N_17692,N_17538,N_17460);
nand U17693 (N_17693,N_17598,N_17487);
nor U17694 (N_17694,N_17449,N_17502);
nor U17695 (N_17695,N_17507,N_17532);
xor U17696 (N_17696,N_17497,N_17453);
xor U17697 (N_17697,N_17589,N_17555);
and U17698 (N_17698,N_17572,N_17593);
nor U17699 (N_17699,N_17440,N_17516);
and U17700 (N_17700,N_17423,N_17463);
xor U17701 (N_17701,N_17574,N_17555);
nand U17702 (N_17702,N_17422,N_17466);
or U17703 (N_17703,N_17519,N_17465);
xnor U17704 (N_17704,N_17431,N_17459);
xnor U17705 (N_17705,N_17564,N_17559);
xor U17706 (N_17706,N_17441,N_17471);
nand U17707 (N_17707,N_17558,N_17453);
xnor U17708 (N_17708,N_17556,N_17440);
and U17709 (N_17709,N_17594,N_17482);
nand U17710 (N_17710,N_17572,N_17418);
nor U17711 (N_17711,N_17589,N_17404);
and U17712 (N_17712,N_17442,N_17538);
xnor U17713 (N_17713,N_17553,N_17490);
or U17714 (N_17714,N_17491,N_17403);
and U17715 (N_17715,N_17532,N_17450);
xor U17716 (N_17716,N_17410,N_17530);
xor U17717 (N_17717,N_17570,N_17540);
and U17718 (N_17718,N_17505,N_17423);
nor U17719 (N_17719,N_17531,N_17598);
nor U17720 (N_17720,N_17441,N_17555);
nor U17721 (N_17721,N_17544,N_17538);
and U17722 (N_17722,N_17500,N_17462);
and U17723 (N_17723,N_17575,N_17452);
xnor U17724 (N_17724,N_17402,N_17587);
or U17725 (N_17725,N_17561,N_17450);
nand U17726 (N_17726,N_17567,N_17503);
nand U17727 (N_17727,N_17487,N_17588);
nor U17728 (N_17728,N_17494,N_17595);
nand U17729 (N_17729,N_17583,N_17554);
nand U17730 (N_17730,N_17511,N_17541);
or U17731 (N_17731,N_17516,N_17537);
nand U17732 (N_17732,N_17552,N_17593);
nand U17733 (N_17733,N_17450,N_17568);
nand U17734 (N_17734,N_17454,N_17583);
or U17735 (N_17735,N_17530,N_17565);
or U17736 (N_17736,N_17481,N_17531);
or U17737 (N_17737,N_17543,N_17560);
and U17738 (N_17738,N_17592,N_17459);
nand U17739 (N_17739,N_17596,N_17452);
xnor U17740 (N_17740,N_17563,N_17419);
and U17741 (N_17741,N_17596,N_17400);
and U17742 (N_17742,N_17424,N_17427);
nor U17743 (N_17743,N_17572,N_17491);
xnor U17744 (N_17744,N_17500,N_17591);
xnor U17745 (N_17745,N_17442,N_17573);
xor U17746 (N_17746,N_17487,N_17501);
nand U17747 (N_17747,N_17527,N_17470);
or U17748 (N_17748,N_17498,N_17591);
and U17749 (N_17749,N_17503,N_17546);
xor U17750 (N_17750,N_17559,N_17409);
nand U17751 (N_17751,N_17435,N_17463);
nor U17752 (N_17752,N_17406,N_17567);
or U17753 (N_17753,N_17410,N_17499);
or U17754 (N_17754,N_17462,N_17567);
nor U17755 (N_17755,N_17444,N_17586);
or U17756 (N_17756,N_17598,N_17441);
nand U17757 (N_17757,N_17557,N_17470);
xnor U17758 (N_17758,N_17408,N_17503);
nor U17759 (N_17759,N_17442,N_17549);
nand U17760 (N_17760,N_17572,N_17460);
nor U17761 (N_17761,N_17437,N_17439);
and U17762 (N_17762,N_17444,N_17410);
xnor U17763 (N_17763,N_17486,N_17474);
and U17764 (N_17764,N_17479,N_17418);
xor U17765 (N_17765,N_17405,N_17566);
or U17766 (N_17766,N_17439,N_17458);
nand U17767 (N_17767,N_17438,N_17471);
nand U17768 (N_17768,N_17573,N_17527);
and U17769 (N_17769,N_17426,N_17459);
or U17770 (N_17770,N_17567,N_17477);
xor U17771 (N_17771,N_17415,N_17581);
xor U17772 (N_17772,N_17481,N_17558);
xor U17773 (N_17773,N_17469,N_17540);
nor U17774 (N_17774,N_17595,N_17575);
nand U17775 (N_17775,N_17501,N_17546);
nand U17776 (N_17776,N_17530,N_17513);
and U17777 (N_17777,N_17483,N_17410);
nand U17778 (N_17778,N_17540,N_17529);
nand U17779 (N_17779,N_17465,N_17505);
or U17780 (N_17780,N_17583,N_17542);
xor U17781 (N_17781,N_17560,N_17440);
and U17782 (N_17782,N_17489,N_17573);
nor U17783 (N_17783,N_17486,N_17456);
and U17784 (N_17784,N_17473,N_17554);
xor U17785 (N_17785,N_17502,N_17592);
or U17786 (N_17786,N_17569,N_17490);
nor U17787 (N_17787,N_17459,N_17531);
nand U17788 (N_17788,N_17576,N_17554);
or U17789 (N_17789,N_17480,N_17401);
nor U17790 (N_17790,N_17428,N_17442);
and U17791 (N_17791,N_17479,N_17569);
nand U17792 (N_17792,N_17528,N_17547);
nand U17793 (N_17793,N_17526,N_17490);
or U17794 (N_17794,N_17558,N_17400);
xor U17795 (N_17795,N_17405,N_17479);
nand U17796 (N_17796,N_17487,N_17421);
nand U17797 (N_17797,N_17419,N_17476);
nand U17798 (N_17798,N_17468,N_17411);
nor U17799 (N_17799,N_17528,N_17430);
nor U17800 (N_17800,N_17715,N_17782);
nand U17801 (N_17801,N_17629,N_17620);
and U17802 (N_17802,N_17703,N_17655);
nor U17803 (N_17803,N_17750,N_17705);
and U17804 (N_17804,N_17669,N_17709);
nand U17805 (N_17805,N_17607,N_17712);
nand U17806 (N_17806,N_17685,N_17732);
nand U17807 (N_17807,N_17762,N_17713);
and U17808 (N_17808,N_17768,N_17640);
nor U17809 (N_17809,N_17614,N_17769);
xor U17810 (N_17810,N_17630,N_17797);
xnor U17811 (N_17811,N_17752,N_17626);
nor U17812 (N_17812,N_17741,N_17653);
nor U17813 (N_17813,N_17722,N_17689);
and U17814 (N_17814,N_17603,N_17729);
xor U17815 (N_17815,N_17618,N_17758);
and U17816 (N_17816,N_17794,N_17785);
nand U17817 (N_17817,N_17706,N_17771);
xnor U17818 (N_17818,N_17682,N_17748);
nand U17819 (N_17819,N_17641,N_17661);
xor U17820 (N_17820,N_17651,N_17781);
nor U17821 (N_17821,N_17680,N_17720);
and U17822 (N_17822,N_17738,N_17683);
and U17823 (N_17823,N_17749,N_17613);
and U17824 (N_17824,N_17791,N_17757);
xor U17825 (N_17825,N_17666,N_17663);
and U17826 (N_17826,N_17612,N_17635);
nor U17827 (N_17827,N_17723,N_17650);
xor U17828 (N_17828,N_17649,N_17701);
nor U17829 (N_17829,N_17658,N_17615);
and U17830 (N_17830,N_17727,N_17724);
and U17831 (N_17831,N_17660,N_17644);
nor U17832 (N_17832,N_17743,N_17792);
nor U17833 (N_17833,N_17774,N_17617);
or U17834 (N_17834,N_17604,N_17754);
xor U17835 (N_17835,N_17605,N_17725);
or U17836 (N_17836,N_17687,N_17796);
or U17837 (N_17837,N_17765,N_17790);
nor U17838 (N_17838,N_17675,N_17773);
xor U17839 (N_17839,N_17733,N_17601);
xor U17840 (N_17840,N_17672,N_17780);
and U17841 (N_17841,N_17783,N_17737);
nand U17842 (N_17842,N_17728,N_17795);
or U17843 (N_17843,N_17721,N_17759);
nor U17844 (N_17844,N_17788,N_17695);
or U17845 (N_17845,N_17735,N_17642);
or U17846 (N_17846,N_17704,N_17657);
and U17847 (N_17847,N_17787,N_17659);
and U17848 (N_17848,N_17770,N_17710);
or U17849 (N_17849,N_17625,N_17609);
or U17850 (N_17850,N_17686,N_17702);
and U17851 (N_17851,N_17673,N_17691);
and U17852 (N_17852,N_17767,N_17714);
or U17853 (N_17853,N_17678,N_17652);
or U17854 (N_17854,N_17654,N_17627);
nor U17855 (N_17855,N_17624,N_17693);
xnor U17856 (N_17856,N_17608,N_17646);
and U17857 (N_17857,N_17690,N_17700);
xor U17858 (N_17858,N_17667,N_17632);
nor U17859 (N_17859,N_17799,N_17622);
or U17860 (N_17860,N_17677,N_17662);
or U17861 (N_17861,N_17637,N_17668);
xnor U17862 (N_17862,N_17656,N_17761);
or U17863 (N_17863,N_17764,N_17692);
and U17864 (N_17864,N_17665,N_17776);
nor U17865 (N_17865,N_17602,N_17756);
xor U17866 (N_17866,N_17789,N_17708);
or U17867 (N_17867,N_17763,N_17694);
and U17868 (N_17868,N_17621,N_17736);
nand U17869 (N_17869,N_17634,N_17628);
and U17870 (N_17870,N_17619,N_17639);
nand U17871 (N_17871,N_17740,N_17718);
nand U17872 (N_17872,N_17631,N_17623);
nor U17873 (N_17873,N_17747,N_17647);
nand U17874 (N_17874,N_17734,N_17670);
xor U17875 (N_17875,N_17664,N_17676);
nand U17876 (N_17876,N_17636,N_17679);
xor U17877 (N_17877,N_17742,N_17755);
nor U17878 (N_17878,N_17674,N_17645);
and U17879 (N_17879,N_17648,N_17600);
nand U17880 (N_17880,N_17730,N_17699);
or U17881 (N_17881,N_17611,N_17616);
nor U17882 (N_17882,N_17638,N_17779);
nor U17883 (N_17883,N_17746,N_17731);
or U17884 (N_17884,N_17711,N_17726);
nor U17885 (N_17885,N_17610,N_17745);
xor U17886 (N_17886,N_17798,N_17793);
nor U17887 (N_17887,N_17778,N_17744);
xor U17888 (N_17888,N_17753,N_17698);
and U17889 (N_17889,N_17633,N_17772);
nor U17890 (N_17890,N_17707,N_17684);
and U17891 (N_17891,N_17681,N_17751);
or U17892 (N_17892,N_17688,N_17643);
and U17893 (N_17893,N_17696,N_17775);
and U17894 (N_17894,N_17760,N_17717);
or U17895 (N_17895,N_17766,N_17719);
or U17896 (N_17896,N_17784,N_17697);
nand U17897 (N_17897,N_17777,N_17606);
xnor U17898 (N_17898,N_17716,N_17786);
xnor U17899 (N_17899,N_17739,N_17671);
xor U17900 (N_17900,N_17782,N_17689);
and U17901 (N_17901,N_17652,N_17743);
nor U17902 (N_17902,N_17792,N_17706);
xnor U17903 (N_17903,N_17624,N_17676);
or U17904 (N_17904,N_17671,N_17630);
xnor U17905 (N_17905,N_17632,N_17729);
and U17906 (N_17906,N_17754,N_17762);
nor U17907 (N_17907,N_17792,N_17709);
and U17908 (N_17908,N_17670,N_17744);
nand U17909 (N_17909,N_17660,N_17694);
or U17910 (N_17910,N_17604,N_17665);
and U17911 (N_17911,N_17703,N_17626);
or U17912 (N_17912,N_17724,N_17634);
nand U17913 (N_17913,N_17627,N_17721);
or U17914 (N_17914,N_17791,N_17721);
nor U17915 (N_17915,N_17619,N_17745);
xor U17916 (N_17916,N_17729,N_17680);
nor U17917 (N_17917,N_17793,N_17660);
nand U17918 (N_17918,N_17724,N_17694);
nor U17919 (N_17919,N_17713,N_17613);
xnor U17920 (N_17920,N_17660,N_17705);
nand U17921 (N_17921,N_17787,N_17611);
xnor U17922 (N_17922,N_17696,N_17614);
xnor U17923 (N_17923,N_17747,N_17699);
or U17924 (N_17924,N_17768,N_17692);
nand U17925 (N_17925,N_17694,N_17606);
and U17926 (N_17926,N_17676,N_17797);
nand U17927 (N_17927,N_17670,N_17622);
nand U17928 (N_17928,N_17741,N_17647);
nand U17929 (N_17929,N_17762,N_17751);
or U17930 (N_17930,N_17736,N_17797);
nor U17931 (N_17931,N_17601,N_17640);
and U17932 (N_17932,N_17638,N_17616);
and U17933 (N_17933,N_17658,N_17611);
nand U17934 (N_17934,N_17678,N_17797);
nand U17935 (N_17935,N_17664,N_17633);
nor U17936 (N_17936,N_17604,N_17631);
xnor U17937 (N_17937,N_17774,N_17698);
nor U17938 (N_17938,N_17798,N_17749);
or U17939 (N_17939,N_17695,N_17653);
nor U17940 (N_17940,N_17625,N_17631);
or U17941 (N_17941,N_17703,N_17686);
or U17942 (N_17942,N_17744,N_17715);
nor U17943 (N_17943,N_17734,N_17620);
xor U17944 (N_17944,N_17728,N_17796);
and U17945 (N_17945,N_17634,N_17774);
xor U17946 (N_17946,N_17622,N_17721);
nor U17947 (N_17947,N_17762,N_17698);
xnor U17948 (N_17948,N_17781,N_17618);
nand U17949 (N_17949,N_17772,N_17750);
and U17950 (N_17950,N_17721,N_17712);
or U17951 (N_17951,N_17642,N_17660);
and U17952 (N_17952,N_17785,N_17648);
and U17953 (N_17953,N_17797,N_17776);
nor U17954 (N_17954,N_17658,N_17746);
and U17955 (N_17955,N_17682,N_17733);
nor U17956 (N_17956,N_17655,N_17736);
or U17957 (N_17957,N_17773,N_17693);
or U17958 (N_17958,N_17636,N_17613);
nor U17959 (N_17959,N_17706,N_17635);
nand U17960 (N_17960,N_17684,N_17733);
and U17961 (N_17961,N_17738,N_17703);
xnor U17962 (N_17962,N_17759,N_17718);
or U17963 (N_17963,N_17776,N_17640);
xnor U17964 (N_17964,N_17646,N_17684);
and U17965 (N_17965,N_17729,N_17740);
and U17966 (N_17966,N_17686,N_17679);
nand U17967 (N_17967,N_17704,N_17613);
and U17968 (N_17968,N_17792,N_17641);
xor U17969 (N_17969,N_17784,N_17642);
or U17970 (N_17970,N_17656,N_17631);
and U17971 (N_17971,N_17629,N_17645);
and U17972 (N_17972,N_17618,N_17755);
nand U17973 (N_17973,N_17701,N_17792);
xnor U17974 (N_17974,N_17755,N_17605);
nand U17975 (N_17975,N_17630,N_17602);
and U17976 (N_17976,N_17749,N_17746);
xnor U17977 (N_17977,N_17723,N_17632);
and U17978 (N_17978,N_17751,N_17618);
or U17979 (N_17979,N_17682,N_17609);
or U17980 (N_17980,N_17757,N_17701);
nor U17981 (N_17981,N_17661,N_17724);
or U17982 (N_17982,N_17735,N_17797);
nor U17983 (N_17983,N_17624,N_17787);
nor U17984 (N_17984,N_17662,N_17718);
or U17985 (N_17985,N_17650,N_17734);
xor U17986 (N_17986,N_17724,N_17745);
or U17987 (N_17987,N_17644,N_17707);
xor U17988 (N_17988,N_17674,N_17627);
and U17989 (N_17989,N_17619,N_17731);
nor U17990 (N_17990,N_17714,N_17660);
nor U17991 (N_17991,N_17661,N_17779);
or U17992 (N_17992,N_17712,N_17625);
xor U17993 (N_17993,N_17783,N_17656);
nand U17994 (N_17994,N_17776,N_17771);
and U17995 (N_17995,N_17777,N_17734);
or U17996 (N_17996,N_17687,N_17619);
nor U17997 (N_17997,N_17736,N_17713);
nor U17998 (N_17998,N_17702,N_17661);
nand U17999 (N_17999,N_17676,N_17693);
or U18000 (N_18000,N_17825,N_17849);
nor U18001 (N_18001,N_17941,N_17930);
nand U18002 (N_18002,N_17815,N_17926);
or U18003 (N_18003,N_17963,N_17996);
nor U18004 (N_18004,N_17982,N_17861);
nand U18005 (N_18005,N_17838,N_17855);
and U18006 (N_18006,N_17836,N_17826);
or U18007 (N_18007,N_17893,N_17839);
nand U18008 (N_18008,N_17809,N_17810);
nand U18009 (N_18009,N_17949,N_17890);
and U18010 (N_18010,N_17846,N_17806);
nand U18011 (N_18011,N_17980,N_17901);
or U18012 (N_18012,N_17962,N_17969);
xor U18013 (N_18013,N_17921,N_17805);
and U18014 (N_18014,N_17957,N_17852);
and U18015 (N_18015,N_17970,N_17801);
and U18016 (N_18016,N_17959,N_17932);
xor U18017 (N_18017,N_17985,N_17802);
nand U18018 (N_18018,N_17975,N_17814);
and U18019 (N_18019,N_17920,N_17891);
or U18020 (N_18020,N_17915,N_17879);
or U18021 (N_18021,N_17813,N_17874);
and U18022 (N_18022,N_17875,N_17888);
nor U18023 (N_18023,N_17840,N_17865);
nor U18024 (N_18024,N_17859,N_17967);
xor U18025 (N_18025,N_17881,N_17880);
nor U18026 (N_18026,N_17974,N_17908);
nor U18027 (N_18027,N_17884,N_17848);
xnor U18028 (N_18028,N_17837,N_17856);
or U18029 (N_18029,N_17863,N_17913);
xnor U18030 (N_18030,N_17943,N_17945);
xor U18031 (N_18031,N_17953,N_17803);
or U18032 (N_18032,N_17937,N_17811);
and U18033 (N_18033,N_17955,N_17981);
or U18034 (N_18034,N_17800,N_17958);
and U18035 (N_18035,N_17829,N_17894);
or U18036 (N_18036,N_17822,N_17964);
nor U18037 (N_18037,N_17978,N_17971);
nor U18038 (N_18038,N_17951,N_17897);
and U18039 (N_18039,N_17946,N_17999);
nor U18040 (N_18040,N_17912,N_17834);
nand U18041 (N_18041,N_17895,N_17997);
xnor U18042 (N_18042,N_17979,N_17988);
xor U18043 (N_18043,N_17927,N_17887);
nor U18044 (N_18044,N_17995,N_17992);
nand U18045 (N_18045,N_17910,N_17807);
nor U18046 (N_18046,N_17972,N_17867);
xnor U18047 (N_18047,N_17832,N_17854);
xnor U18048 (N_18048,N_17804,N_17876);
nand U18049 (N_18049,N_17853,N_17914);
and U18050 (N_18050,N_17886,N_17917);
nor U18051 (N_18051,N_17878,N_17847);
or U18052 (N_18052,N_17872,N_17828);
nor U18053 (N_18053,N_17823,N_17862);
and U18054 (N_18054,N_17821,N_17960);
xor U18055 (N_18055,N_17950,N_17973);
nor U18056 (N_18056,N_17991,N_17843);
or U18057 (N_18057,N_17983,N_17864);
nand U18058 (N_18058,N_17952,N_17860);
nor U18059 (N_18059,N_17904,N_17889);
nand U18060 (N_18060,N_17909,N_17812);
or U18061 (N_18061,N_17850,N_17934);
xor U18062 (N_18062,N_17907,N_17986);
xnor U18063 (N_18063,N_17936,N_17905);
or U18064 (N_18064,N_17948,N_17844);
nand U18065 (N_18065,N_17987,N_17883);
or U18066 (N_18066,N_17977,N_17922);
nand U18067 (N_18067,N_17870,N_17871);
nand U18068 (N_18068,N_17944,N_17831);
nand U18069 (N_18069,N_17947,N_17841);
xnor U18070 (N_18070,N_17956,N_17898);
nor U18071 (N_18071,N_17998,N_17994);
nor U18072 (N_18072,N_17954,N_17976);
nand U18073 (N_18073,N_17938,N_17919);
or U18074 (N_18074,N_17818,N_17918);
or U18075 (N_18075,N_17924,N_17935);
xor U18076 (N_18076,N_17906,N_17896);
xnor U18077 (N_18077,N_17830,N_17989);
nor U18078 (N_18078,N_17965,N_17961);
or U18079 (N_18079,N_17868,N_17869);
or U18080 (N_18080,N_17928,N_17824);
and U18081 (N_18081,N_17816,N_17851);
or U18082 (N_18082,N_17968,N_17903);
nor U18083 (N_18083,N_17808,N_17873);
and U18084 (N_18084,N_17916,N_17990);
xor U18085 (N_18085,N_17827,N_17931);
xnor U18086 (N_18086,N_17925,N_17842);
or U18087 (N_18087,N_17845,N_17833);
or U18088 (N_18088,N_17885,N_17933);
xor U18089 (N_18089,N_17858,N_17899);
or U18090 (N_18090,N_17929,N_17866);
or U18091 (N_18091,N_17984,N_17900);
nor U18092 (N_18092,N_17942,N_17940);
and U18093 (N_18093,N_17923,N_17877);
xor U18094 (N_18094,N_17902,N_17819);
and U18095 (N_18095,N_17835,N_17966);
nand U18096 (N_18096,N_17817,N_17993);
or U18097 (N_18097,N_17857,N_17892);
nor U18098 (N_18098,N_17911,N_17820);
xor U18099 (N_18099,N_17882,N_17939);
nand U18100 (N_18100,N_17945,N_17933);
or U18101 (N_18101,N_17959,N_17871);
xor U18102 (N_18102,N_17856,N_17816);
and U18103 (N_18103,N_17829,N_17832);
nand U18104 (N_18104,N_17874,N_17938);
nor U18105 (N_18105,N_17910,N_17876);
or U18106 (N_18106,N_17823,N_17802);
xor U18107 (N_18107,N_17872,N_17847);
and U18108 (N_18108,N_17957,N_17977);
nor U18109 (N_18109,N_17998,N_17995);
nor U18110 (N_18110,N_17801,N_17943);
nand U18111 (N_18111,N_17965,N_17981);
nor U18112 (N_18112,N_17850,N_17959);
nand U18113 (N_18113,N_17985,N_17839);
nand U18114 (N_18114,N_17814,N_17884);
nand U18115 (N_18115,N_17915,N_17858);
nor U18116 (N_18116,N_17893,N_17829);
nand U18117 (N_18117,N_17908,N_17977);
xor U18118 (N_18118,N_17853,N_17957);
nand U18119 (N_18119,N_17967,N_17808);
xnor U18120 (N_18120,N_17822,N_17938);
nand U18121 (N_18121,N_17807,N_17934);
nand U18122 (N_18122,N_17970,N_17941);
nor U18123 (N_18123,N_17806,N_17927);
nand U18124 (N_18124,N_17828,N_17875);
xor U18125 (N_18125,N_17943,N_17930);
nand U18126 (N_18126,N_17993,N_17917);
nor U18127 (N_18127,N_17995,N_17990);
nand U18128 (N_18128,N_17854,N_17839);
or U18129 (N_18129,N_17863,N_17930);
nor U18130 (N_18130,N_17957,N_17940);
nor U18131 (N_18131,N_17916,N_17889);
xor U18132 (N_18132,N_17858,N_17830);
or U18133 (N_18133,N_17842,N_17837);
nor U18134 (N_18134,N_17990,N_17828);
and U18135 (N_18135,N_17863,N_17961);
nand U18136 (N_18136,N_17802,N_17942);
xor U18137 (N_18137,N_17978,N_17997);
and U18138 (N_18138,N_17887,N_17991);
nor U18139 (N_18139,N_17904,N_17935);
xor U18140 (N_18140,N_17988,N_17829);
or U18141 (N_18141,N_17876,N_17987);
xor U18142 (N_18142,N_17882,N_17904);
and U18143 (N_18143,N_17944,N_17836);
nand U18144 (N_18144,N_17880,N_17885);
nor U18145 (N_18145,N_17942,N_17923);
nand U18146 (N_18146,N_17878,N_17920);
nor U18147 (N_18147,N_17814,N_17862);
nand U18148 (N_18148,N_17943,N_17968);
nor U18149 (N_18149,N_17917,N_17921);
nand U18150 (N_18150,N_17990,N_17895);
and U18151 (N_18151,N_17877,N_17800);
xor U18152 (N_18152,N_17849,N_17905);
xnor U18153 (N_18153,N_17807,N_17913);
xor U18154 (N_18154,N_17948,N_17926);
xnor U18155 (N_18155,N_17969,N_17942);
xor U18156 (N_18156,N_17921,N_17959);
xor U18157 (N_18157,N_17905,N_17809);
nand U18158 (N_18158,N_17879,N_17887);
nand U18159 (N_18159,N_17966,N_17971);
nand U18160 (N_18160,N_17887,N_17847);
xnor U18161 (N_18161,N_17952,N_17964);
nand U18162 (N_18162,N_17814,N_17930);
nor U18163 (N_18163,N_17979,N_17969);
xor U18164 (N_18164,N_17945,N_17897);
or U18165 (N_18165,N_17890,N_17909);
or U18166 (N_18166,N_17845,N_17893);
nand U18167 (N_18167,N_17844,N_17821);
nand U18168 (N_18168,N_17829,N_17905);
nor U18169 (N_18169,N_17961,N_17825);
xnor U18170 (N_18170,N_17910,N_17863);
or U18171 (N_18171,N_17961,N_17851);
or U18172 (N_18172,N_17908,N_17897);
nand U18173 (N_18173,N_17903,N_17805);
or U18174 (N_18174,N_17905,N_17804);
or U18175 (N_18175,N_17823,N_17806);
nand U18176 (N_18176,N_17970,N_17830);
nor U18177 (N_18177,N_17888,N_17857);
xor U18178 (N_18178,N_17912,N_17824);
nand U18179 (N_18179,N_17928,N_17985);
and U18180 (N_18180,N_17889,N_17857);
or U18181 (N_18181,N_17812,N_17824);
and U18182 (N_18182,N_17893,N_17997);
nor U18183 (N_18183,N_17958,N_17889);
or U18184 (N_18184,N_17978,N_17814);
xor U18185 (N_18185,N_17886,N_17951);
nor U18186 (N_18186,N_17943,N_17999);
or U18187 (N_18187,N_17826,N_17874);
and U18188 (N_18188,N_17998,N_17990);
or U18189 (N_18189,N_17871,N_17844);
and U18190 (N_18190,N_17944,N_17876);
nor U18191 (N_18191,N_17964,N_17911);
and U18192 (N_18192,N_17899,N_17945);
and U18193 (N_18193,N_17991,N_17840);
xor U18194 (N_18194,N_17983,N_17914);
or U18195 (N_18195,N_17963,N_17843);
and U18196 (N_18196,N_17911,N_17876);
or U18197 (N_18197,N_17833,N_17842);
nor U18198 (N_18198,N_17950,N_17822);
or U18199 (N_18199,N_17900,N_17963);
nor U18200 (N_18200,N_18051,N_18143);
nand U18201 (N_18201,N_18106,N_18163);
nand U18202 (N_18202,N_18138,N_18112);
xnor U18203 (N_18203,N_18150,N_18126);
nand U18204 (N_18204,N_18152,N_18041);
nor U18205 (N_18205,N_18077,N_18118);
and U18206 (N_18206,N_18119,N_18030);
nor U18207 (N_18207,N_18181,N_18107);
xnor U18208 (N_18208,N_18039,N_18148);
and U18209 (N_18209,N_18100,N_18146);
and U18210 (N_18210,N_18042,N_18014);
or U18211 (N_18211,N_18010,N_18123);
nand U18212 (N_18212,N_18061,N_18131);
or U18213 (N_18213,N_18125,N_18103);
nor U18214 (N_18214,N_18018,N_18104);
and U18215 (N_18215,N_18044,N_18004);
nor U18216 (N_18216,N_18006,N_18159);
xor U18217 (N_18217,N_18192,N_18080);
or U18218 (N_18218,N_18083,N_18048);
xor U18219 (N_18219,N_18066,N_18183);
and U18220 (N_18220,N_18057,N_18108);
or U18221 (N_18221,N_18185,N_18087);
xnor U18222 (N_18222,N_18137,N_18120);
nand U18223 (N_18223,N_18016,N_18176);
xnor U18224 (N_18224,N_18151,N_18145);
or U18225 (N_18225,N_18160,N_18015);
nand U18226 (N_18226,N_18035,N_18179);
and U18227 (N_18227,N_18020,N_18177);
nand U18228 (N_18228,N_18095,N_18170);
nor U18229 (N_18229,N_18058,N_18194);
and U18230 (N_18230,N_18188,N_18136);
nor U18231 (N_18231,N_18054,N_18189);
nor U18232 (N_18232,N_18111,N_18141);
and U18233 (N_18233,N_18115,N_18047);
and U18234 (N_18234,N_18193,N_18049);
or U18235 (N_18235,N_18062,N_18088);
or U18236 (N_18236,N_18195,N_18199);
nand U18237 (N_18237,N_18075,N_18026);
and U18238 (N_18238,N_18040,N_18074);
nand U18239 (N_18239,N_18086,N_18182);
nor U18240 (N_18240,N_18069,N_18122);
and U18241 (N_18241,N_18024,N_18096);
and U18242 (N_18242,N_18158,N_18187);
nand U18243 (N_18243,N_18029,N_18157);
xnor U18244 (N_18244,N_18171,N_18084);
nand U18245 (N_18245,N_18129,N_18021);
and U18246 (N_18246,N_18027,N_18005);
nor U18247 (N_18247,N_18043,N_18133);
xnor U18248 (N_18248,N_18135,N_18144);
and U18249 (N_18249,N_18071,N_18003);
xnor U18250 (N_18250,N_18037,N_18156);
nor U18251 (N_18251,N_18079,N_18031);
nor U18252 (N_18252,N_18046,N_18117);
and U18253 (N_18253,N_18198,N_18009);
xnor U18254 (N_18254,N_18007,N_18025);
nor U18255 (N_18255,N_18164,N_18134);
nand U18256 (N_18256,N_18022,N_18165);
nand U18257 (N_18257,N_18000,N_18184);
nor U18258 (N_18258,N_18169,N_18056);
or U18259 (N_18259,N_18168,N_18196);
xnor U18260 (N_18260,N_18110,N_18081);
nand U18261 (N_18261,N_18068,N_18052);
or U18262 (N_18262,N_18094,N_18162);
and U18263 (N_18263,N_18154,N_18050);
and U18264 (N_18264,N_18023,N_18078);
and U18265 (N_18265,N_18028,N_18127);
nor U18266 (N_18266,N_18032,N_18002);
nor U18267 (N_18267,N_18105,N_18017);
xor U18268 (N_18268,N_18113,N_18167);
or U18269 (N_18269,N_18091,N_18019);
nor U18270 (N_18270,N_18067,N_18098);
nand U18271 (N_18271,N_18053,N_18197);
and U18272 (N_18272,N_18063,N_18101);
xnor U18273 (N_18273,N_18139,N_18099);
xor U18274 (N_18274,N_18011,N_18178);
nor U18275 (N_18275,N_18155,N_18092);
nor U18276 (N_18276,N_18102,N_18116);
nand U18277 (N_18277,N_18036,N_18038);
nor U18278 (N_18278,N_18045,N_18161);
nand U18279 (N_18279,N_18173,N_18034);
nand U18280 (N_18280,N_18191,N_18085);
xor U18281 (N_18281,N_18093,N_18072);
and U18282 (N_18282,N_18142,N_18012);
or U18283 (N_18283,N_18090,N_18166);
and U18284 (N_18284,N_18008,N_18064);
nor U18285 (N_18285,N_18121,N_18060);
and U18286 (N_18286,N_18132,N_18082);
xor U18287 (N_18287,N_18186,N_18055);
xor U18288 (N_18288,N_18073,N_18109);
or U18289 (N_18289,N_18114,N_18070);
and U18290 (N_18290,N_18190,N_18001);
xor U18291 (N_18291,N_18097,N_18147);
nand U18292 (N_18292,N_18149,N_18130);
nor U18293 (N_18293,N_18174,N_18089);
or U18294 (N_18294,N_18128,N_18153);
nor U18295 (N_18295,N_18140,N_18124);
nand U18296 (N_18296,N_18059,N_18076);
xor U18297 (N_18297,N_18013,N_18065);
nor U18298 (N_18298,N_18180,N_18175);
or U18299 (N_18299,N_18172,N_18033);
or U18300 (N_18300,N_18120,N_18096);
or U18301 (N_18301,N_18191,N_18047);
and U18302 (N_18302,N_18173,N_18078);
nand U18303 (N_18303,N_18178,N_18027);
and U18304 (N_18304,N_18196,N_18017);
and U18305 (N_18305,N_18116,N_18160);
and U18306 (N_18306,N_18154,N_18003);
nand U18307 (N_18307,N_18123,N_18120);
or U18308 (N_18308,N_18055,N_18026);
nand U18309 (N_18309,N_18032,N_18125);
and U18310 (N_18310,N_18115,N_18174);
xor U18311 (N_18311,N_18043,N_18187);
and U18312 (N_18312,N_18172,N_18159);
and U18313 (N_18313,N_18066,N_18005);
xor U18314 (N_18314,N_18135,N_18072);
and U18315 (N_18315,N_18035,N_18037);
and U18316 (N_18316,N_18030,N_18135);
nand U18317 (N_18317,N_18193,N_18097);
nand U18318 (N_18318,N_18133,N_18178);
and U18319 (N_18319,N_18120,N_18185);
nor U18320 (N_18320,N_18097,N_18014);
xnor U18321 (N_18321,N_18052,N_18193);
or U18322 (N_18322,N_18147,N_18051);
nor U18323 (N_18323,N_18139,N_18164);
and U18324 (N_18324,N_18135,N_18164);
xor U18325 (N_18325,N_18000,N_18089);
nor U18326 (N_18326,N_18166,N_18106);
nand U18327 (N_18327,N_18086,N_18161);
and U18328 (N_18328,N_18031,N_18045);
nor U18329 (N_18329,N_18094,N_18135);
nand U18330 (N_18330,N_18001,N_18182);
and U18331 (N_18331,N_18134,N_18109);
xor U18332 (N_18332,N_18044,N_18023);
xor U18333 (N_18333,N_18151,N_18199);
nor U18334 (N_18334,N_18122,N_18189);
nor U18335 (N_18335,N_18045,N_18177);
nand U18336 (N_18336,N_18111,N_18191);
nor U18337 (N_18337,N_18043,N_18188);
or U18338 (N_18338,N_18062,N_18020);
and U18339 (N_18339,N_18024,N_18004);
nor U18340 (N_18340,N_18192,N_18155);
xnor U18341 (N_18341,N_18131,N_18013);
and U18342 (N_18342,N_18126,N_18180);
or U18343 (N_18343,N_18168,N_18072);
xnor U18344 (N_18344,N_18003,N_18048);
nor U18345 (N_18345,N_18098,N_18013);
and U18346 (N_18346,N_18092,N_18175);
nor U18347 (N_18347,N_18011,N_18047);
xor U18348 (N_18348,N_18116,N_18001);
nand U18349 (N_18349,N_18053,N_18100);
nor U18350 (N_18350,N_18061,N_18179);
nand U18351 (N_18351,N_18020,N_18023);
xor U18352 (N_18352,N_18157,N_18036);
nor U18353 (N_18353,N_18047,N_18104);
nand U18354 (N_18354,N_18180,N_18107);
nand U18355 (N_18355,N_18190,N_18193);
nor U18356 (N_18356,N_18172,N_18088);
and U18357 (N_18357,N_18096,N_18094);
or U18358 (N_18358,N_18071,N_18125);
or U18359 (N_18359,N_18114,N_18173);
or U18360 (N_18360,N_18167,N_18052);
or U18361 (N_18361,N_18045,N_18043);
nand U18362 (N_18362,N_18171,N_18142);
nand U18363 (N_18363,N_18127,N_18085);
nand U18364 (N_18364,N_18130,N_18122);
or U18365 (N_18365,N_18071,N_18154);
xor U18366 (N_18366,N_18051,N_18013);
xor U18367 (N_18367,N_18055,N_18166);
and U18368 (N_18368,N_18047,N_18125);
and U18369 (N_18369,N_18177,N_18046);
and U18370 (N_18370,N_18019,N_18030);
nor U18371 (N_18371,N_18068,N_18039);
and U18372 (N_18372,N_18155,N_18046);
nor U18373 (N_18373,N_18040,N_18008);
xor U18374 (N_18374,N_18067,N_18157);
nand U18375 (N_18375,N_18133,N_18080);
and U18376 (N_18376,N_18071,N_18149);
or U18377 (N_18377,N_18131,N_18184);
nor U18378 (N_18378,N_18105,N_18179);
nor U18379 (N_18379,N_18155,N_18089);
nand U18380 (N_18380,N_18055,N_18156);
xor U18381 (N_18381,N_18055,N_18125);
nand U18382 (N_18382,N_18112,N_18007);
and U18383 (N_18383,N_18197,N_18064);
xnor U18384 (N_18384,N_18166,N_18069);
or U18385 (N_18385,N_18189,N_18143);
and U18386 (N_18386,N_18133,N_18007);
nand U18387 (N_18387,N_18154,N_18198);
nor U18388 (N_18388,N_18050,N_18021);
or U18389 (N_18389,N_18146,N_18020);
nand U18390 (N_18390,N_18097,N_18107);
or U18391 (N_18391,N_18060,N_18017);
or U18392 (N_18392,N_18066,N_18046);
and U18393 (N_18393,N_18004,N_18131);
or U18394 (N_18394,N_18177,N_18010);
or U18395 (N_18395,N_18072,N_18080);
or U18396 (N_18396,N_18135,N_18126);
and U18397 (N_18397,N_18138,N_18050);
nand U18398 (N_18398,N_18102,N_18105);
nand U18399 (N_18399,N_18196,N_18003);
xnor U18400 (N_18400,N_18231,N_18359);
nor U18401 (N_18401,N_18273,N_18242);
nor U18402 (N_18402,N_18220,N_18236);
nand U18403 (N_18403,N_18375,N_18331);
and U18404 (N_18404,N_18216,N_18207);
nor U18405 (N_18405,N_18298,N_18230);
or U18406 (N_18406,N_18218,N_18263);
nor U18407 (N_18407,N_18338,N_18381);
xnor U18408 (N_18408,N_18264,N_18366);
nor U18409 (N_18409,N_18357,N_18363);
or U18410 (N_18410,N_18252,N_18208);
and U18411 (N_18411,N_18307,N_18310);
or U18412 (N_18412,N_18294,N_18389);
and U18413 (N_18413,N_18232,N_18267);
nand U18414 (N_18414,N_18392,N_18314);
nand U18415 (N_18415,N_18300,N_18317);
xor U18416 (N_18416,N_18391,N_18385);
or U18417 (N_18417,N_18274,N_18271);
nor U18418 (N_18418,N_18316,N_18374);
nor U18419 (N_18419,N_18334,N_18202);
and U18420 (N_18420,N_18382,N_18203);
nor U18421 (N_18421,N_18255,N_18305);
nand U18422 (N_18422,N_18272,N_18283);
xor U18423 (N_18423,N_18353,N_18379);
nor U18424 (N_18424,N_18284,N_18365);
or U18425 (N_18425,N_18348,N_18269);
nand U18426 (N_18426,N_18393,N_18318);
nand U18427 (N_18427,N_18280,N_18336);
xor U18428 (N_18428,N_18278,N_18251);
and U18429 (N_18429,N_18350,N_18211);
nand U18430 (N_18430,N_18356,N_18341);
xor U18431 (N_18431,N_18398,N_18384);
or U18432 (N_18432,N_18219,N_18226);
nor U18433 (N_18433,N_18282,N_18248);
xnor U18434 (N_18434,N_18210,N_18227);
or U18435 (N_18435,N_18320,N_18339);
nand U18436 (N_18436,N_18308,N_18299);
nand U18437 (N_18437,N_18249,N_18370);
or U18438 (N_18438,N_18289,N_18337);
nand U18439 (N_18439,N_18261,N_18325);
and U18440 (N_18440,N_18380,N_18228);
nand U18441 (N_18441,N_18394,N_18346);
nor U18442 (N_18442,N_18286,N_18266);
xnor U18443 (N_18443,N_18367,N_18340);
or U18444 (N_18444,N_18277,N_18215);
nand U18445 (N_18445,N_18200,N_18313);
or U18446 (N_18446,N_18291,N_18332);
nor U18447 (N_18447,N_18268,N_18324);
nor U18448 (N_18448,N_18352,N_18262);
or U18449 (N_18449,N_18281,N_18302);
and U18450 (N_18450,N_18354,N_18233);
xnor U18451 (N_18451,N_18209,N_18238);
nor U18452 (N_18452,N_18279,N_18388);
and U18453 (N_18453,N_18396,N_18201);
nand U18454 (N_18454,N_18378,N_18344);
nor U18455 (N_18455,N_18383,N_18377);
and U18456 (N_18456,N_18223,N_18214);
nand U18457 (N_18457,N_18270,N_18371);
or U18458 (N_18458,N_18257,N_18205);
and U18459 (N_18459,N_18247,N_18326);
xnor U18460 (N_18460,N_18243,N_18303);
xor U18461 (N_18461,N_18204,N_18306);
or U18462 (N_18462,N_18234,N_18329);
or U18463 (N_18463,N_18321,N_18225);
and U18464 (N_18464,N_18342,N_18237);
or U18465 (N_18465,N_18309,N_18369);
xor U18466 (N_18466,N_18387,N_18241);
or U18467 (N_18467,N_18295,N_18217);
nand U18468 (N_18468,N_18358,N_18376);
or U18469 (N_18469,N_18304,N_18287);
nor U18470 (N_18470,N_18292,N_18256);
nor U18471 (N_18471,N_18285,N_18355);
and U18472 (N_18472,N_18347,N_18296);
nand U18473 (N_18473,N_18399,N_18301);
and U18474 (N_18474,N_18319,N_18293);
nand U18475 (N_18475,N_18290,N_18361);
xnor U18476 (N_18476,N_18327,N_18253);
nor U18477 (N_18477,N_18235,N_18351);
xor U18478 (N_18478,N_18259,N_18275);
or U18479 (N_18479,N_18260,N_18240);
nor U18480 (N_18480,N_18335,N_18222);
nor U18481 (N_18481,N_18213,N_18312);
and U18482 (N_18482,N_18245,N_18368);
nand U18483 (N_18483,N_18328,N_18323);
nor U18484 (N_18484,N_18349,N_18244);
nor U18485 (N_18485,N_18360,N_18288);
and U18486 (N_18486,N_18362,N_18212);
xor U18487 (N_18487,N_18311,N_18390);
or U18488 (N_18488,N_18386,N_18246);
nand U18489 (N_18489,N_18250,N_18221);
or U18490 (N_18490,N_18297,N_18315);
or U18491 (N_18491,N_18254,N_18372);
and U18492 (N_18492,N_18239,N_18343);
or U18493 (N_18493,N_18322,N_18206);
xor U18494 (N_18494,N_18373,N_18276);
xnor U18495 (N_18495,N_18265,N_18224);
xor U18496 (N_18496,N_18333,N_18258);
nand U18497 (N_18497,N_18345,N_18395);
nand U18498 (N_18498,N_18397,N_18229);
nand U18499 (N_18499,N_18364,N_18330);
nor U18500 (N_18500,N_18230,N_18297);
xor U18501 (N_18501,N_18326,N_18371);
nor U18502 (N_18502,N_18380,N_18260);
nand U18503 (N_18503,N_18253,N_18284);
nand U18504 (N_18504,N_18338,N_18218);
nor U18505 (N_18505,N_18247,N_18292);
and U18506 (N_18506,N_18234,N_18328);
nor U18507 (N_18507,N_18385,N_18216);
or U18508 (N_18508,N_18349,N_18201);
and U18509 (N_18509,N_18292,N_18344);
xnor U18510 (N_18510,N_18348,N_18355);
xnor U18511 (N_18511,N_18367,N_18398);
nand U18512 (N_18512,N_18353,N_18242);
xnor U18513 (N_18513,N_18301,N_18277);
nor U18514 (N_18514,N_18399,N_18356);
and U18515 (N_18515,N_18258,N_18292);
and U18516 (N_18516,N_18330,N_18219);
nand U18517 (N_18517,N_18306,N_18220);
nand U18518 (N_18518,N_18366,N_18356);
nand U18519 (N_18519,N_18206,N_18202);
or U18520 (N_18520,N_18220,N_18276);
nor U18521 (N_18521,N_18239,N_18318);
nand U18522 (N_18522,N_18263,N_18357);
and U18523 (N_18523,N_18357,N_18318);
or U18524 (N_18524,N_18389,N_18342);
and U18525 (N_18525,N_18339,N_18282);
and U18526 (N_18526,N_18298,N_18287);
and U18527 (N_18527,N_18374,N_18335);
or U18528 (N_18528,N_18275,N_18391);
or U18529 (N_18529,N_18291,N_18339);
xnor U18530 (N_18530,N_18352,N_18322);
nand U18531 (N_18531,N_18358,N_18353);
and U18532 (N_18532,N_18244,N_18237);
xnor U18533 (N_18533,N_18342,N_18378);
nor U18534 (N_18534,N_18325,N_18210);
nor U18535 (N_18535,N_18248,N_18207);
nor U18536 (N_18536,N_18214,N_18213);
xnor U18537 (N_18537,N_18211,N_18393);
nand U18538 (N_18538,N_18211,N_18294);
nor U18539 (N_18539,N_18300,N_18256);
xnor U18540 (N_18540,N_18308,N_18318);
xor U18541 (N_18541,N_18219,N_18207);
and U18542 (N_18542,N_18320,N_18274);
xor U18543 (N_18543,N_18215,N_18261);
nor U18544 (N_18544,N_18254,N_18398);
or U18545 (N_18545,N_18257,N_18250);
nor U18546 (N_18546,N_18231,N_18303);
nand U18547 (N_18547,N_18388,N_18226);
nor U18548 (N_18548,N_18336,N_18293);
xnor U18549 (N_18549,N_18227,N_18350);
xor U18550 (N_18550,N_18301,N_18272);
or U18551 (N_18551,N_18359,N_18308);
nor U18552 (N_18552,N_18218,N_18330);
or U18553 (N_18553,N_18384,N_18365);
nor U18554 (N_18554,N_18232,N_18224);
and U18555 (N_18555,N_18303,N_18366);
xnor U18556 (N_18556,N_18390,N_18382);
and U18557 (N_18557,N_18233,N_18257);
nand U18558 (N_18558,N_18288,N_18286);
and U18559 (N_18559,N_18252,N_18342);
and U18560 (N_18560,N_18271,N_18210);
nand U18561 (N_18561,N_18354,N_18257);
or U18562 (N_18562,N_18282,N_18369);
or U18563 (N_18563,N_18227,N_18379);
and U18564 (N_18564,N_18268,N_18313);
xnor U18565 (N_18565,N_18363,N_18372);
and U18566 (N_18566,N_18294,N_18276);
nand U18567 (N_18567,N_18260,N_18379);
xor U18568 (N_18568,N_18366,N_18240);
nor U18569 (N_18569,N_18241,N_18252);
xnor U18570 (N_18570,N_18262,N_18277);
and U18571 (N_18571,N_18305,N_18385);
nor U18572 (N_18572,N_18210,N_18207);
xnor U18573 (N_18573,N_18224,N_18345);
nand U18574 (N_18574,N_18278,N_18315);
xor U18575 (N_18575,N_18338,N_18251);
and U18576 (N_18576,N_18263,N_18377);
nand U18577 (N_18577,N_18215,N_18229);
nand U18578 (N_18578,N_18256,N_18330);
or U18579 (N_18579,N_18344,N_18348);
or U18580 (N_18580,N_18299,N_18372);
nor U18581 (N_18581,N_18332,N_18388);
nand U18582 (N_18582,N_18285,N_18385);
nor U18583 (N_18583,N_18229,N_18331);
and U18584 (N_18584,N_18393,N_18346);
and U18585 (N_18585,N_18271,N_18212);
or U18586 (N_18586,N_18208,N_18356);
nand U18587 (N_18587,N_18232,N_18373);
xnor U18588 (N_18588,N_18267,N_18295);
xor U18589 (N_18589,N_18392,N_18273);
and U18590 (N_18590,N_18201,N_18218);
or U18591 (N_18591,N_18227,N_18214);
and U18592 (N_18592,N_18315,N_18263);
nand U18593 (N_18593,N_18278,N_18255);
or U18594 (N_18594,N_18329,N_18213);
and U18595 (N_18595,N_18303,N_18235);
xnor U18596 (N_18596,N_18280,N_18350);
xor U18597 (N_18597,N_18293,N_18215);
xnor U18598 (N_18598,N_18264,N_18327);
and U18599 (N_18599,N_18380,N_18232);
or U18600 (N_18600,N_18532,N_18483);
nand U18601 (N_18601,N_18589,N_18482);
and U18602 (N_18602,N_18590,N_18449);
and U18603 (N_18603,N_18547,N_18453);
and U18604 (N_18604,N_18518,N_18406);
xnor U18605 (N_18605,N_18447,N_18462);
or U18606 (N_18606,N_18527,N_18591);
nand U18607 (N_18607,N_18520,N_18558);
nand U18608 (N_18608,N_18515,N_18461);
nand U18609 (N_18609,N_18409,N_18481);
or U18610 (N_18610,N_18470,N_18567);
nor U18611 (N_18611,N_18427,N_18487);
or U18612 (N_18612,N_18469,N_18566);
nor U18613 (N_18613,N_18542,N_18458);
nor U18614 (N_18614,N_18457,N_18504);
and U18615 (N_18615,N_18599,N_18555);
xnor U18616 (N_18616,N_18577,N_18440);
xor U18617 (N_18617,N_18403,N_18534);
nor U18618 (N_18618,N_18522,N_18404);
and U18619 (N_18619,N_18552,N_18425);
xnor U18620 (N_18620,N_18432,N_18421);
nand U18621 (N_18621,N_18438,N_18492);
xnor U18622 (N_18622,N_18490,N_18581);
xor U18623 (N_18623,N_18560,N_18557);
nor U18624 (N_18624,N_18586,N_18410);
or U18625 (N_18625,N_18496,N_18569);
or U18626 (N_18626,N_18538,N_18422);
nor U18627 (N_18627,N_18519,N_18476);
and U18628 (N_18628,N_18594,N_18511);
or U18629 (N_18629,N_18510,N_18420);
nor U18630 (N_18630,N_18582,N_18587);
or U18631 (N_18631,N_18568,N_18465);
xor U18632 (N_18632,N_18554,N_18486);
or U18633 (N_18633,N_18544,N_18494);
or U18634 (N_18634,N_18405,N_18443);
xor U18635 (N_18635,N_18561,N_18417);
or U18636 (N_18636,N_18489,N_18573);
nor U18637 (N_18637,N_18502,N_18508);
nand U18638 (N_18638,N_18549,N_18578);
or U18639 (N_18639,N_18446,N_18546);
xnor U18640 (N_18640,N_18479,N_18433);
and U18641 (N_18641,N_18407,N_18435);
nor U18642 (N_18642,N_18436,N_18588);
nand U18643 (N_18643,N_18414,N_18450);
and U18644 (N_18644,N_18467,N_18595);
and U18645 (N_18645,N_18418,N_18439);
nor U18646 (N_18646,N_18579,N_18500);
nand U18647 (N_18647,N_18553,N_18529);
nand U18648 (N_18648,N_18548,N_18495);
nor U18649 (N_18649,N_18451,N_18575);
or U18650 (N_18650,N_18545,N_18408);
nand U18651 (N_18651,N_18464,N_18456);
nor U18652 (N_18652,N_18572,N_18583);
nand U18653 (N_18653,N_18434,N_18537);
nor U18654 (N_18654,N_18517,N_18499);
or U18655 (N_18655,N_18525,N_18412);
or U18656 (N_18656,N_18400,N_18463);
or U18657 (N_18657,N_18533,N_18541);
nand U18658 (N_18658,N_18513,N_18441);
xor U18659 (N_18659,N_18478,N_18426);
or U18660 (N_18660,N_18585,N_18563);
nor U18661 (N_18661,N_18430,N_18593);
nor U18662 (N_18662,N_18562,N_18550);
nand U18663 (N_18663,N_18480,N_18459);
nand U18664 (N_18664,N_18523,N_18471);
and U18665 (N_18665,N_18466,N_18570);
nor U18666 (N_18666,N_18592,N_18484);
nand U18667 (N_18667,N_18423,N_18431);
nor U18668 (N_18668,N_18503,N_18596);
nand U18669 (N_18669,N_18419,N_18536);
nand U18670 (N_18670,N_18597,N_18501);
xnor U18671 (N_18671,N_18401,N_18576);
xnor U18672 (N_18672,N_18428,N_18516);
xnor U18673 (N_18673,N_18580,N_18477);
nand U18674 (N_18674,N_18551,N_18565);
xnor U18675 (N_18675,N_18488,N_18455);
and U18676 (N_18676,N_18413,N_18507);
nor U18677 (N_18677,N_18564,N_18584);
nor U18678 (N_18678,N_18506,N_18543);
and U18679 (N_18679,N_18528,N_18474);
nor U18680 (N_18680,N_18472,N_18445);
nand U18681 (N_18681,N_18402,N_18497);
nand U18682 (N_18682,N_18574,N_18505);
or U18683 (N_18683,N_18416,N_18512);
nand U18684 (N_18684,N_18415,N_18468);
nor U18685 (N_18685,N_18526,N_18571);
and U18686 (N_18686,N_18460,N_18521);
nand U18687 (N_18687,N_18559,N_18429);
xnor U18688 (N_18688,N_18444,N_18454);
nand U18689 (N_18689,N_18539,N_18473);
nand U18690 (N_18690,N_18491,N_18485);
or U18691 (N_18691,N_18411,N_18540);
and U18692 (N_18692,N_18509,N_18448);
xor U18693 (N_18693,N_18475,N_18598);
nor U18694 (N_18694,N_18493,N_18531);
nand U18695 (N_18695,N_18437,N_18524);
or U18696 (N_18696,N_18424,N_18442);
nand U18697 (N_18697,N_18556,N_18530);
and U18698 (N_18698,N_18514,N_18535);
or U18699 (N_18699,N_18498,N_18452);
or U18700 (N_18700,N_18449,N_18473);
xor U18701 (N_18701,N_18465,N_18446);
nor U18702 (N_18702,N_18446,N_18484);
nor U18703 (N_18703,N_18481,N_18525);
nand U18704 (N_18704,N_18545,N_18527);
nand U18705 (N_18705,N_18556,N_18580);
and U18706 (N_18706,N_18492,N_18594);
xnor U18707 (N_18707,N_18549,N_18453);
nor U18708 (N_18708,N_18423,N_18500);
or U18709 (N_18709,N_18407,N_18419);
xnor U18710 (N_18710,N_18566,N_18461);
nor U18711 (N_18711,N_18564,N_18524);
xor U18712 (N_18712,N_18553,N_18592);
or U18713 (N_18713,N_18470,N_18585);
nand U18714 (N_18714,N_18581,N_18574);
nor U18715 (N_18715,N_18553,N_18593);
and U18716 (N_18716,N_18481,N_18569);
nand U18717 (N_18717,N_18499,N_18405);
nor U18718 (N_18718,N_18561,N_18477);
nand U18719 (N_18719,N_18494,N_18516);
nor U18720 (N_18720,N_18514,N_18599);
and U18721 (N_18721,N_18544,N_18430);
nand U18722 (N_18722,N_18506,N_18420);
and U18723 (N_18723,N_18495,N_18550);
or U18724 (N_18724,N_18528,N_18502);
nor U18725 (N_18725,N_18415,N_18524);
or U18726 (N_18726,N_18505,N_18441);
nor U18727 (N_18727,N_18562,N_18422);
and U18728 (N_18728,N_18423,N_18568);
or U18729 (N_18729,N_18494,N_18413);
and U18730 (N_18730,N_18500,N_18433);
xor U18731 (N_18731,N_18498,N_18460);
or U18732 (N_18732,N_18591,N_18590);
or U18733 (N_18733,N_18494,N_18545);
and U18734 (N_18734,N_18505,N_18474);
nor U18735 (N_18735,N_18462,N_18544);
nor U18736 (N_18736,N_18419,N_18498);
and U18737 (N_18737,N_18520,N_18559);
or U18738 (N_18738,N_18558,N_18567);
and U18739 (N_18739,N_18410,N_18429);
or U18740 (N_18740,N_18483,N_18543);
xor U18741 (N_18741,N_18498,N_18437);
nand U18742 (N_18742,N_18530,N_18554);
or U18743 (N_18743,N_18512,N_18460);
nand U18744 (N_18744,N_18432,N_18437);
and U18745 (N_18745,N_18519,N_18412);
xor U18746 (N_18746,N_18450,N_18515);
and U18747 (N_18747,N_18462,N_18507);
xnor U18748 (N_18748,N_18463,N_18451);
nand U18749 (N_18749,N_18438,N_18555);
and U18750 (N_18750,N_18442,N_18553);
xor U18751 (N_18751,N_18402,N_18417);
or U18752 (N_18752,N_18506,N_18462);
or U18753 (N_18753,N_18516,N_18507);
or U18754 (N_18754,N_18421,N_18427);
and U18755 (N_18755,N_18582,N_18471);
nand U18756 (N_18756,N_18477,N_18542);
and U18757 (N_18757,N_18599,N_18407);
nor U18758 (N_18758,N_18408,N_18419);
nor U18759 (N_18759,N_18504,N_18403);
or U18760 (N_18760,N_18456,N_18457);
nand U18761 (N_18761,N_18573,N_18524);
and U18762 (N_18762,N_18564,N_18550);
nor U18763 (N_18763,N_18584,N_18523);
nand U18764 (N_18764,N_18596,N_18492);
and U18765 (N_18765,N_18515,N_18498);
nor U18766 (N_18766,N_18584,N_18583);
and U18767 (N_18767,N_18592,N_18545);
and U18768 (N_18768,N_18568,N_18410);
nor U18769 (N_18769,N_18551,N_18574);
and U18770 (N_18770,N_18461,N_18428);
xor U18771 (N_18771,N_18404,N_18421);
nor U18772 (N_18772,N_18574,N_18404);
and U18773 (N_18773,N_18570,N_18531);
nor U18774 (N_18774,N_18441,N_18457);
xnor U18775 (N_18775,N_18505,N_18466);
nand U18776 (N_18776,N_18474,N_18539);
xor U18777 (N_18777,N_18441,N_18596);
nor U18778 (N_18778,N_18579,N_18596);
nand U18779 (N_18779,N_18522,N_18447);
and U18780 (N_18780,N_18455,N_18542);
nand U18781 (N_18781,N_18481,N_18484);
and U18782 (N_18782,N_18452,N_18427);
nand U18783 (N_18783,N_18530,N_18492);
and U18784 (N_18784,N_18462,N_18527);
and U18785 (N_18785,N_18473,N_18466);
or U18786 (N_18786,N_18521,N_18426);
and U18787 (N_18787,N_18503,N_18499);
and U18788 (N_18788,N_18442,N_18432);
xnor U18789 (N_18789,N_18405,N_18541);
nor U18790 (N_18790,N_18521,N_18583);
xnor U18791 (N_18791,N_18541,N_18583);
nand U18792 (N_18792,N_18593,N_18427);
or U18793 (N_18793,N_18417,N_18504);
or U18794 (N_18794,N_18461,N_18431);
nor U18795 (N_18795,N_18438,N_18436);
nand U18796 (N_18796,N_18571,N_18542);
and U18797 (N_18797,N_18492,N_18475);
xor U18798 (N_18798,N_18400,N_18518);
nor U18799 (N_18799,N_18417,N_18472);
nor U18800 (N_18800,N_18617,N_18784);
nor U18801 (N_18801,N_18774,N_18745);
nand U18802 (N_18802,N_18685,N_18664);
nand U18803 (N_18803,N_18792,N_18741);
nand U18804 (N_18804,N_18688,N_18608);
and U18805 (N_18805,N_18750,N_18666);
nor U18806 (N_18806,N_18739,N_18692);
or U18807 (N_18807,N_18781,N_18706);
and U18808 (N_18808,N_18621,N_18683);
nand U18809 (N_18809,N_18655,N_18768);
nand U18810 (N_18810,N_18734,N_18767);
nor U18811 (N_18811,N_18737,N_18749);
and U18812 (N_18812,N_18636,N_18733);
xor U18813 (N_18813,N_18738,N_18678);
nand U18814 (N_18814,N_18607,N_18791);
xnor U18815 (N_18815,N_18799,N_18662);
nand U18816 (N_18816,N_18728,N_18712);
nor U18817 (N_18817,N_18777,N_18732);
nand U18818 (N_18818,N_18795,N_18744);
and U18819 (N_18819,N_18703,N_18796);
nand U18820 (N_18820,N_18619,N_18691);
or U18821 (N_18821,N_18758,N_18632);
and U18822 (N_18822,N_18742,N_18793);
and U18823 (N_18823,N_18725,N_18652);
or U18824 (N_18824,N_18630,N_18711);
nand U18825 (N_18825,N_18633,N_18762);
or U18826 (N_18826,N_18714,N_18629);
or U18827 (N_18827,N_18623,N_18708);
nor U18828 (N_18828,N_18650,N_18618);
nand U18829 (N_18829,N_18794,N_18746);
nor U18830 (N_18830,N_18600,N_18788);
xor U18831 (N_18831,N_18686,N_18769);
nand U18832 (N_18832,N_18626,N_18753);
xnor U18833 (N_18833,N_18687,N_18727);
or U18834 (N_18834,N_18716,N_18743);
nor U18835 (N_18835,N_18614,N_18783);
nand U18836 (N_18836,N_18681,N_18748);
xor U18837 (N_18837,N_18730,N_18698);
xnor U18838 (N_18838,N_18635,N_18710);
or U18839 (N_18839,N_18722,N_18751);
or U18840 (N_18840,N_18644,N_18773);
xnor U18841 (N_18841,N_18663,N_18640);
xnor U18842 (N_18842,N_18606,N_18676);
xor U18843 (N_18843,N_18785,N_18638);
and U18844 (N_18844,N_18603,N_18671);
and U18845 (N_18845,N_18694,N_18651);
and U18846 (N_18846,N_18770,N_18693);
nor U18847 (N_18847,N_18735,N_18756);
nor U18848 (N_18848,N_18709,N_18639);
and U18849 (N_18849,N_18720,N_18726);
nor U18850 (N_18850,N_18721,N_18778);
nor U18851 (N_18851,N_18604,N_18715);
or U18852 (N_18852,N_18675,N_18602);
or U18853 (N_18853,N_18622,N_18661);
xor U18854 (N_18854,N_18699,N_18659);
xor U18855 (N_18855,N_18754,N_18631);
nor U18856 (N_18856,N_18667,N_18747);
or U18857 (N_18857,N_18647,N_18787);
xnor U18858 (N_18858,N_18625,N_18776);
or U18859 (N_18859,N_18701,N_18723);
or U18860 (N_18860,N_18665,N_18763);
nor U18861 (N_18861,N_18757,N_18643);
and U18862 (N_18862,N_18615,N_18702);
xor U18863 (N_18863,N_18717,N_18668);
nand U18864 (N_18864,N_18772,N_18680);
and U18865 (N_18865,N_18616,N_18609);
nand U18866 (N_18866,N_18660,N_18782);
and U18867 (N_18867,N_18786,N_18764);
nor U18868 (N_18868,N_18775,N_18677);
xor U18869 (N_18869,N_18620,N_18766);
or U18870 (N_18870,N_18779,N_18612);
nand U18871 (N_18871,N_18718,N_18637);
nor U18872 (N_18872,N_18642,N_18752);
nor U18873 (N_18873,N_18755,N_18765);
and U18874 (N_18874,N_18627,N_18669);
xnor U18875 (N_18875,N_18780,N_18670);
nand U18876 (N_18876,N_18611,N_18713);
nand U18877 (N_18877,N_18628,N_18649);
nor U18878 (N_18878,N_18634,N_18695);
and U18879 (N_18879,N_18696,N_18736);
nand U18880 (N_18880,N_18624,N_18648);
or U18881 (N_18881,N_18673,N_18760);
or U18882 (N_18882,N_18790,N_18724);
or U18883 (N_18883,N_18672,N_18689);
xnor U18884 (N_18884,N_18731,N_18697);
or U18885 (N_18885,N_18729,N_18700);
or U18886 (N_18886,N_18719,N_18707);
nor U18887 (N_18887,N_18674,N_18771);
or U18888 (N_18888,N_18605,N_18601);
or U18889 (N_18889,N_18789,N_18658);
and U18890 (N_18890,N_18656,N_18797);
xnor U18891 (N_18891,N_18645,N_18653);
or U18892 (N_18892,N_18682,N_18798);
or U18893 (N_18893,N_18613,N_18704);
xor U18894 (N_18894,N_18610,N_18740);
or U18895 (N_18895,N_18690,N_18641);
or U18896 (N_18896,N_18759,N_18646);
or U18897 (N_18897,N_18679,N_18761);
or U18898 (N_18898,N_18684,N_18654);
and U18899 (N_18899,N_18705,N_18657);
and U18900 (N_18900,N_18775,N_18641);
or U18901 (N_18901,N_18652,N_18608);
and U18902 (N_18902,N_18725,N_18624);
or U18903 (N_18903,N_18791,N_18634);
xnor U18904 (N_18904,N_18671,N_18679);
nor U18905 (N_18905,N_18714,N_18666);
nand U18906 (N_18906,N_18659,N_18786);
and U18907 (N_18907,N_18712,N_18788);
and U18908 (N_18908,N_18665,N_18768);
nor U18909 (N_18909,N_18604,N_18703);
nand U18910 (N_18910,N_18794,N_18766);
nand U18911 (N_18911,N_18678,N_18797);
nor U18912 (N_18912,N_18664,N_18677);
or U18913 (N_18913,N_18646,N_18674);
nand U18914 (N_18914,N_18673,N_18654);
and U18915 (N_18915,N_18625,N_18757);
nand U18916 (N_18916,N_18703,N_18631);
and U18917 (N_18917,N_18690,N_18627);
xor U18918 (N_18918,N_18629,N_18762);
xnor U18919 (N_18919,N_18735,N_18777);
xor U18920 (N_18920,N_18694,N_18797);
xnor U18921 (N_18921,N_18676,N_18603);
and U18922 (N_18922,N_18707,N_18755);
and U18923 (N_18923,N_18771,N_18621);
or U18924 (N_18924,N_18675,N_18716);
and U18925 (N_18925,N_18786,N_18629);
nand U18926 (N_18926,N_18632,N_18785);
and U18927 (N_18927,N_18631,N_18740);
nand U18928 (N_18928,N_18758,N_18714);
nand U18929 (N_18929,N_18760,N_18645);
or U18930 (N_18930,N_18795,N_18774);
nor U18931 (N_18931,N_18636,N_18713);
and U18932 (N_18932,N_18713,N_18666);
or U18933 (N_18933,N_18685,N_18757);
or U18934 (N_18934,N_18750,N_18608);
xnor U18935 (N_18935,N_18794,N_18792);
and U18936 (N_18936,N_18615,N_18745);
nand U18937 (N_18937,N_18618,N_18633);
nor U18938 (N_18938,N_18653,N_18796);
or U18939 (N_18939,N_18731,N_18632);
or U18940 (N_18940,N_18718,N_18795);
or U18941 (N_18941,N_18734,N_18777);
xor U18942 (N_18942,N_18688,N_18772);
nand U18943 (N_18943,N_18709,N_18757);
xnor U18944 (N_18944,N_18788,N_18617);
nand U18945 (N_18945,N_18711,N_18769);
nor U18946 (N_18946,N_18637,N_18639);
or U18947 (N_18947,N_18617,N_18746);
nand U18948 (N_18948,N_18706,N_18613);
xnor U18949 (N_18949,N_18766,N_18626);
xor U18950 (N_18950,N_18600,N_18755);
nor U18951 (N_18951,N_18726,N_18762);
nor U18952 (N_18952,N_18684,N_18677);
and U18953 (N_18953,N_18739,N_18630);
or U18954 (N_18954,N_18679,N_18663);
nor U18955 (N_18955,N_18633,N_18613);
nor U18956 (N_18956,N_18748,N_18790);
xor U18957 (N_18957,N_18740,N_18767);
nand U18958 (N_18958,N_18687,N_18611);
nor U18959 (N_18959,N_18743,N_18677);
or U18960 (N_18960,N_18704,N_18731);
nand U18961 (N_18961,N_18679,N_18745);
nand U18962 (N_18962,N_18667,N_18690);
xnor U18963 (N_18963,N_18642,N_18679);
or U18964 (N_18964,N_18646,N_18673);
nand U18965 (N_18965,N_18680,N_18603);
nand U18966 (N_18966,N_18784,N_18640);
xnor U18967 (N_18967,N_18705,N_18656);
or U18968 (N_18968,N_18600,N_18724);
nor U18969 (N_18969,N_18767,N_18656);
nor U18970 (N_18970,N_18750,N_18681);
and U18971 (N_18971,N_18734,N_18794);
nand U18972 (N_18972,N_18733,N_18642);
or U18973 (N_18973,N_18669,N_18601);
nand U18974 (N_18974,N_18649,N_18717);
nor U18975 (N_18975,N_18786,N_18756);
nor U18976 (N_18976,N_18739,N_18656);
nor U18977 (N_18977,N_18611,N_18607);
and U18978 (N_18978,N_18696,N_18751);
nor U18979 (N_18979,N_18671,N_18698);
nor U18980 (N_18980,N_18683,N_18676);
or U18981 (N_18981,N_18604,N_18682);
nor U18982 (N_18982,N_18682,N_18786);
xnor U18983 (N_18983,N_18609,N_18783);
or U18984 (N_18984,N_18780,N_18621);
and U18985 (N_18985,N_18674,N_18742);
nand U18986 (N_18986,N_18674,N_18774);
or U18987 (N_18987,N_18606,N_18636);
nor U18988 (N_18988,N_18789,N_18666);
or U18989 (N_18989,N_18636,N_18660);
and U18990 (N_18990,N_18679,N_18694);
or U18991 (N_18991,N_18667,N_18792);
nor U18992 (N_18992,N_18635,N_18645);
nand U18993 (N_18993,N_18724,N_18631);
or U18994 (N_18994,N_18663,N_18779);
xnor U18995 (N_18995,N_18621,N_18654);
nand U18996 (N_18996,N_18726,N_18772);
and U18997 (N_18997,N_18739,N_18661);
and U18998 (N_18998,N_18797,N_18767);
nor U18999 (N_18999,N_18696,N_18622);
xor U19000 (N_19000,N_18870,N_18992);
nor U19001 (N_19001,N_18809,N_18942);
and U19002 (N_19002,N_18977,N_18833);
nand U19003 (N_19003,N_18903,N_18879);
nor U19004 (N_19004,N_18963,N_18839);
nor U19005 (N_19005,N_18905,N_18914);
and U19006 (N_19006,N_18834,N_18867);
or U19007 (N_19007,N_18873,N_18869);
and U19008 (N_19008,N_18924,N_18910);
nor U19009 (N_19009,N_18849,N_18952);
or U19010 (N_19010,N_18934,N_18904);
nand U19011 (N_19011,N_18965,N_18956);
nor U19012 (N_19012,N_18872,N_18909);
or U19013 (N_19013,N_18936,N_18827);
or U19014 (N_19014,N_18915,N_18962);
xnor U19015 (N_19015,N_18807,N_18967);
nand U19016 (N_19016,N_18832,N_18989);
xor U19017 (N_19017,N_18923,N_18955);
and U19018 (N_19018,N_18864,N_18803);
nand U19019 (N_19019,N_18902,N_18928);
xnor U19020 (N_19020,N_18874,N_18985);
or U19021 (N_19021,N_18953,N_18950);
and U19022 (N_19022,N_18811,N_18815);
and U19023 (N_19023,N_18971,N_18932);
xnor U19024 (N_19024,N_18845,N_18906);
and U19025 (N_19025,N_18972,N_18897);
and U19026 (N_19026,N_18899,N_18895);
xor U19027 (N_19027,N_18861,N_18947);
nor U19028 (N_19028,N_18812,N_18964);
nand U19029 (N_19029,N_18958,N_18853);
or U19030 (N_19030,N_18800,N_18920);
nand U19031 (N_19031,N_18898,N_18841);
xor U19032 (N_19032,N_18860,N_18970);
xnor U19033 (N_19033,N_18913,N_18959);
xnor U19034 (N_19034,N_18865,N_18939);
or U19035 (N_19035,N_18856,N_18945);
and U19036 (N_19036,N_18886,N_18810);
nand U19037 (N_19037,N_18937,N_18922);
and U19038 (N_19038,N_18966,N_18896);
xnor U19039 (N_19039,N_18804,N_18995);
and U19040 (N_19040,N_18911,N_18976);
nor U19041 (N_19041,N_18818,N_18877);
xor U19042 (N_19042,N_18883,N_18900);
and U19043 (N_19043,N_18929,N_18893);
xor U19044 (N_19044,N_18984,N_18931);
and U19045 (N_19045,N_18851,N_18823);
nand U19046 (N_19046,N_18938,N_18921);
and U19047 (N_19047,N_18979,N_18829);
xor U19048 (N_19048,N_18933,N_18871);
or U19049 (N_19049,N_18948,N_18862);
nor U19050 (N_19050,N_18978,N_18935);
xnor U19051 (N_19051,N_18944,N_18997);
nor U19052 (N_19052,N_18987,N_18875);
nor U19053 (N_19053,N_18954,N_18941);
nor U19054 (N_19054,N_18943,N_18863);
and U19055 (N_19055,N_18822,N_18973);
and U19056 (N_19056,N_18847,N_18859);
nor U19057 (N_19057,N_18991,N_18806);
and U19058 (N_19058,N_18828,N_18908);
xor U19059 (N_19059,N_18994,N_18982);
nor U19060 (N_19060,N_18890,N_18835);
nand U19061 (N_19061,N_18918,N_18986);
or U19062 (N_19062,N_18820,N_18830);
nand U19063 (N_19063,N_18961,N_18843);
and U19064 (N_19064,N_18996,N_18848);
and U19065 (N_19065,N_18892,N_18831);
xor U19066 (N_19066,N_18891,N_18983);
xor U19067 (N_19067,N_18808,N_18825);
nand U19068 (N_19068,N_18840,N_18975);
and U19069 (N_19069,N_18889,N_18949);
nand U19070 (N_19070,N_18878,N_18926);
or U19071 (N_19071,N_18824,N_18907);
nand U19072 (N_19072,N_18998,N_18802);
and U19073 (N_19073,N_18855,N_18940);
and U19074 (N_19074,N_18946,N_18917);
xor U19075 (N_19075,N_18858,N_18816);
nand U19076 (N_19076,N_18842,N_18990);
nor U19077 (N_19077,N_18969,N_18957);
nand U19078 (N_19078,N_18857,N_18838);
nand U19079 (N_19079,N_18801,N_18854);
nor U19080 (N_19080,N_18876,N_18805);
xor U19081 (N_19081,N_18852,N_18814);
nand U19082 (N_19082,N_18999,N_18884);
or U19083 (N_19083,N_18960,N_18826);
nand U19084 (N_19084,N_18881,N_18837);
nor U19085 (N_19085,N_18819,N_18988);
nor U19086 (N_19086,N_18916,N_18912);
and U19087 (N_19087,N_18919,N_18821);
or U19088 (N_19088,N_18813,N_18974);
nor U19089 (N_19089,N_18885,N_18846);
xnor U19090 (N_19090,N_18981,N_18887);
and U19091 (N_19091,N_18980,N_18868);
nand U19092 (N_19092,N_18880,N_18968);
xor U19093 (N_19093,N_18866,N_18993);
nand U19094 (N_19094,N_18850,N_18894);
xnor U19095 (N_19095,N_18927,N_18888);
nand U19096 (N_19096,N_18836,N_18951);
or U19097 (N_19097,N_18817,N_18901);
and U19098 (N_19098,N_18882,N_18925);
nand U19099 (N_19099,N_18844,N_18930);
nor U19100 (N_19100,N_18947,N_18877);
xnor U19101 (N_19101,N_18994,N_18902);
nand U19102 (N_19102,N_18878,N_18991);
nand U19103 (N_19103,N_18925,N_18885);
xnor U19104 (N_19104,N_18811,N_18802);
nand U19105 (N_19105,N_18945,N_18847);
and U19106 (N_19106,N_18990,N_18848);
or U19107 (N_19107,N_18818,N_18934);
or U19108 (N_19108,N_18951,N_18967);
nor U19109 (N_19109,N_18801,N_18950);
or U19110 (N_19110,N_18940,N_18995);
nand U19111 (N_19111,N_18966,N_18986);
or U19112 (N_19112,N_18843,N_18865);
xnor U19113 (N_19113,N_18821,N_18881);
and U19114 (N_19114,N_18973,N_18885);
nand U19115 (N_19115,N_18919,N_18837);
or U19116 (N_19116,N_18976,N_18929);
xnor U19117 (N_19117,N_18801,N_18803);
and U19118 (N_19118,N_18968,N_18916);
xnor U19119 (N_19119,N_18997,N_18815);
nand U19120 (N_19120,N_18814,N_18937);
or U19121 (N_19121,N_18817,N_18902);
and U19122 (N_19122,N_18859,N_18866);
or U19123 (N_19123,N_18916,N_18951);
xor U19124 (N_19124,N_18934,N_18876);
or U19125 (N_19125,N_18865,N_18946);
nand U19126 (N_19126,N_18974,N_18821);
nor U19127 (N_19127,N_18841,N_18862);
or U19128 (N_19128,N_18810,N_18955);
nor U19129 (N_19129,N_18879,N_18957);
or U19130 (N_19130,N_18925,N_18836);
xnor U19131 (N_19131,N_18976,N_18952);
and U19132 (N_19132,N_18975,N_18842);
nand U19133 (N_19133,N_18985,N_18826);
nand U19134 (N_19134,N_18963,N_18908);
and U19135 (N_19135,N_18829,N_18846);
or U19136 (N_19136,N_18939,N_18932);
and U19137 (N_19137,N_18804,N_18828);
and U19138 (N_19138,N_18834,N_18981);
xnor U19139 (N_19139,N_18837,N_18930);
nor U19140 (N_19140,N_18873,N_18941);
nand U19141 (N_19141,N_18989,N_18852);
xor U19142 (N_19142,N_18839,N_18970);
or U19143 (N_19143,N_18815,N_18976);
and U19144 (N_19144,N_18885,N_18826);
nor U19145 (N_19145,N_18888,N_18938);
xor U19146 (N_19146,N_18908,N_18877);
nor U19147 (N_19147,N_18898,N_18980);
or U19148 (N_19148,N_18942,N_18832);
nor U19149 (N_19149,N_18954,N_18835);
or U19150 (N_19150,N_18966,N_18848);
nor U19151 (N_19151,N_18915,N_18936);
and U19152 (N_19152,N_18974,N_18842);
and U19153 (N_19153,N_18859,N_18846);
or U19154 (N_19154,N_18983,N_18995);
or U19155 (N_19155,N_18847,N_18811);
nand U19156 (N_19156,N_18866,N_18896);
xor U19157 (N_19157,N_18901,N_18822);
nand U19158 (N_19158,N_18953,N_18934);
xnor U19159 (N_19159,N_18856,N_18988);
nor U19160 (N_19160,N_18917,N_18809);
and U19161 (N_19161,N_18886,N_18824);
xnor U19162 (N_19162,N_18971,N_18909);
xor U19163 (N_19163,N_18966,N_18835);
nor U19164 (N_19164,N_18805,N_18961);
xor U19165 (N_19165,N_18803,N_18971);
and U19166 (N_19166,N_18899,N_18967);
xnor U19167 (N_19167,N_18882,N_18802);
nor U19168 (N_19168,N_18948,N_18898);
or U19169 (N_19169,N_18944,N_18821);
nand U19170 (N_19170,N_18829,N_18921);
nand U19171 (N_19171,N_18852,N_18913);
and U19172 (N_19172,N_18898,N_18833);
nand U19173 (N_19173,N_18948,N_18927);
xor U19174 (N_19174,N_18921,N_18903);
or U19175 (N_19175,N_18988,N_18899);
xnor U19176 (N_19176,N_18865,N_18901);
nor U19177 (N_19177,N_18945,N_18992);
nor U19178 (N_19178,N_18984,N_18899);
or U19179 (N_19179,N_18826,N_18814);
or U19180 (N_19180,N_18898,N_18803);
nor U19181 (N_19181,N_18903,N_18984);
xor U19182 (N_19182,N_18849,N_18902);
nor U19183 (N_19183,N_18802,N_18833);
and U19184 (N_19184,N_18801,N_18973);
xnor U19185 (N_19185,N_18997,N_18859);
xnor U19186 (N_19186,N_18909,N_18862);
xor U19187 (N_19187,N_18923,N_18925);
or U19188 (N_19188,N_18938,N_18908);
or U19189 (N_19189,N_18962,N_18929);
and U19190 (N_19190,N_18988,N_18801);
xnor U19191 (N_19191,N_18924,N_18884);
nor U19192 (N_19192,N_18996,N_18905);
and U19193 (N_19193,N_18865,N_18917);
nand U19194 (N_19194,N_18904,N_18834);
nand U19195 (N_19195,N_18962,N_18996);
and U19196 (N_19196,N_18931,N_18954);
xnor U19197 (N_19197,N_18993,N_18951);
and U19198 (N_19198,N_18918,N_18942);
or U19199 (N_19199,N_18824,N_18919);
nand U19200 (N_19200,N_19121,N_19011);
or U19201 (N_19201,N_19094,N_19108);
nor U19202 (N_19202,N_19080,N_19020);
nand U19203 (N_19203,N_19050,N_19199);
and U19204 (N_19204,N_19099,N_19107);
and U19205 (N_19205,N_19089,N_19082);
or U19206 (N_19206,N_19017,N_19132);
nand U19207 (N_19207,N_19163,N_19119);
xnor U19208 (N_19208,N_19019,N_19183);
or U19209 (N_19209,N_19178,N_19090);
or U19210 (N_19210,N_19148,N_19113);
nand U19211 (N_19211,N_19028,N_19127);
or U19212 (N_19212,N_19155,N_19047);
nor U19213 (N_19213,N_19006,N_19154);
and U19214 (N_19214,N_19166,N_19065);
or U19215 (N_19215,N_19165,N_19152);
nor U19216 (N_19216,N_19110,N_19038);
or U19217 (N_19217,N_19195,N_19035);
or U19218 (N_19218,N_19077,N_19109);
and U19219 (N_19219,N_19069,N_19133);
nand U19220 (N_19220,N_19198,N_19051);
or U19221 (N_19221,N_19029,N_19180);
xor U19222 (N_19222,N_19040,N_19004);
or U19223 (N_19223,N_19140,N_19061);
or U19224 (N_19224,N_19088,N_19106);
and U19225 (N_19225,N_19102,N_19086);
xnor U19226 (N_19226,N_19056,N_19101);
xnor U19227 (N_19227,N_19042,N_19012);
nor U19228 (N_19228,N_19066,N_19062);
nand U19229 (N_19229,N_19150,N_19024);
xor U19230 (N_19230,N_19187,N_19045);
nor U19231 (N_19231,N_19126,N_19072);
xor U19232 (N_19232,N_19001,N_19125);
nand U19233 (N_19233,N_19085,N_19075);
or U19234 (N_19234,N_19139,N_19067);
nor U19235 (N_19235,N_19158,N_19053);
or U19236 (N_19236,N_19087,N_19117);
or U19237 (N_19237,N_19189,N_19096);
xnor U19238 (N_19238,N_19197,N_19058);
xor U19239 (N_19239,N_19172,N_19073);
nand U19240 (N_19240,N_19013,N_19091);
nor U19241 (N_19241,N_19185,N_19000);
nor U19242 (N_19242,N_19100,N_19010);
or U19243 (N_19243,N_19151,N_19179);
and U19244 (N_19244,N_19092,N_19167);
nor U19245 (N_19245,N_19002,N_19046);
or U19246 (N_19246,N_19134,N_19018);
xor U19247 (N_19247,N_19142,N_19093);
and U19248 (N_19248,N_19146,N_19039);
xnor U19249 (N_19249,N_19049,N_19016);
xnor U19250 (N_19250,N_19015,N_19120);
xor U19251 (N_19251,N_19114,N_19115);
xor U19252 (N_19252,N_19057,N_19111);
nand U19253 (N_19253,N_19025,N_19141);
and U19254 (N_19254,N_19164,N_19123);
or U19255 (N_19255,N_19138,N_19174);
and U19256 (N_19256,N_19009,N_19043);
and U19257 (N_19257,N_19005,N_19149);
xor U19258 (N_19258,N_19177,N_19124);
nor U19259 (N_19259,N_19137,N_19135);
and U19260 (N_19260,N_19034,N_19031);
nand U19261 (N_19261,N_19162,N_19054);
nor U19262 (N_19262,N_19129,N_19190);
nor U19263 (N_19263,N_19191,N_19157);
nand U19264 (N_19264,N_19169,N_19003);
nor U19265 (N_19265,N_19014,N_19036);
nor U19266 (N_19266,N_19026,N_19098);
or U19267 (N_19267,N_19032,N_19084);
nor U19268 (N_19268,N_19074,N_19192);
and U19269 (N_19269,N_19181,N_19131);
nor U19270 (N_19270,N_19112,N_19143);
nor U19271 (N_19271,N_19173,N_19027);
or U19272 (N_19272,N_19136,N_19064);
nand U19273 (N_19273,N_19048,N_19168);
and U19274 (N_19274,N_19188,N_19156);
nor U19275 (N_19275,N_19153,N_19081);
xor U19276 (N_19276,N_19170,N_19122);
nor U19277 (N_19277,N_19193,N_19184);
nor U19278 (N_19278,N_19159,N_19083);
nor U19279 (N_19279,N_19097,N_19052);
xnor U19280 (N_19280,N_19104,N_19145);
or U19281 (N_19281,N_19030,N_19182);
nor U19282 (N_19282,N_19186,N_19079);
nand U19283 (N_19283,N_19007,N_19130);
and U19284 (N_19284,N_19055,N_19196);
nor U19285 (N_19285,N_19095,N_19071);
nand U19286 (N_19286,N_19068,N_19171);
nand U19287 (N_19287,N_19144,N_19037);
xnor U19288 (N_19288,N_19175,N_19022);
xor U19289 (N_19289,N_19076,N_19103);
nand U19290 (N_19290,N_19060,N_19023);
nor U19291 (N_19291,N_19070,N_19078);
nand U19292 (N_19292,N_19128,N_19059);
nand U19293 (N_19293,N_19118,N_19063);
nand U19294 (N_19294,N_19041,N_19021);
and U19295 (N_19295,N_19160,N_19161);
xor U19296 (N_19296,N_19194,N_19147);
xor U19297 (N_19297,N_19033,N_19176);
nand U19298 (N_19298,N_19008,N_19105);
and U19299 (N_19299,N_19116,N_19044);
and U19300 (N_19300,N_19035,N_19011);
nor U19301 (N_19301,N_19162,N_19158);
nand U19302 (N_19302,N_19047,N_19014);
nand U19303 (N_19303,N_19135,N_19151);
nor U19304 (N_19304,N_19121,N_19095);
nor U19305 (N_19305,N_19159,N_19041);
nor U19306 (N_19306,N_19164,N_19126);
xor U19307 (N_19307,N_19195,N_19052);
xnor U19308 (N_19308,N_19157,N_19051);
and U19309 (N_19309,N_19102,N_19026);
xnor U19310 (N_19310,N_19159,N_19169);
or U19311 (N_19311,N_19105,N_19178);
or U19312 (N_19312,N_19101,N_19052);
nor U19313 (N_19313,N_19140,N_19000);
or U19314 (N_19314,N_19184,N_19009);
xor U19315 (N_19315,N_19041,N_19191);
xnor U19316 (N_19316,N_19179,N_19113);
nor U19317 (N_19317,N_19044,N_19022);
nor U19318 (N_19318,N_19093,N_19105);
nor U19319 (N_19319,N_19088,N_19001);
and U19320 (N_19320,N_19006,N_19014);
xor U19321 (N_19321,N_19139,N_19158);
or U19322 (N_19322,N_19089,N_19171);
nand U19323 (N_19323,N_19153,N_19092);
xnor U19324 (N_19324,N_19027,N_19071);
or U19325 (N_19325,N_19074,N_19091);
nor U19326 (N_19326,N_19057,N_19191);
and U19327 (N_19327,N_19131,N_19092);
and U19328 (N_19328,N_19110,N_19190);
or U19329 (N_19329,N_19104,N_19191);
and U19330 (N_19330,N_19068,N_19128);
nor U19331 (N_19331,N_19091,N_19114);
or U19332 (N_19332,N_19086,N_19167);
and U19333 (N_19333,N_19059,N_19083);
xnor U19334 (N_19334,N_19136,N_19162);
and U19335 (N_19335,N_19050,N_19131);
or U19336 (N_19336,N_19044,N_19185);
nand U19337 (N_19337,N_19157,N_19131);
or U19338 (N_19338,N_19191,N_19096);
nor U19339 (N_19339,N_19184,N_19145);
or U19340 (N_19340,N_19120,N_19148);
nor U19341 (N_19341,N_19147,N_19076);
nand U19342 (N_19342,N_19033,N_19180);
xnor U19343 (N_19343,N_19080,N_19196);
and U19344 (N_19344,N_19029,N_19068);
or U19345 (N_19345,N_19110,N_19162);
nand U19346 (N_19346,N_19179,N_19152);
nand U19347 (N_19347,N_19136,N_19134);
or U19348 (N_19348,N_19137,N_19166);
nand U19349 (N_19349,N_19123,N_19011);
nand U19350 (N_19350,N_19138,N_19188);
nor U19351 (N_19351,N_19172,N_19001);
or U19352 (N_19352,N_19033,N_19061);
xor U19353 (N_19353,N_19048,N_19023);
nor U19354 (N_19354,N_19181,N_19157);
and U19355 (N_19355,N_19159,N_19121);
nor U19356 (N_19356,N_19081,N_19172);
nor U19357 (N_19357,N_19111,N_19054);
and U19358 (N_19358,N_19134,N_19185);
xnor U19359 (N_19359,N_19114,N_19056);
xnor U19360 (N_19360,N_19027,N_19157);
nand U19361 (N_19361,N_19018,N_19006);
nor U19362 (N_19362,N_19067,N_19085);
or U19363 (N_19363,N_19085,N_19171);
xor U19364 (N_19364,N_19132,N_19150);
nor U19365 (N_19365,N_19067,N_19025);
and U19366 (N_19366,N_19055,N_19054);
nand U19367 (N_19367,N_19071,N_19113);
nand U19368 (N_19368,N_19030,N_19148);
and U19369 (N_19369,N_19061,N_19043);
nor U19370 (N_19370,N_19084,N_19186);
nor U19371 (N_19371,N_19136,N_19127);
nor U19372 (N_19372,N_19188,N_19185);
nor U19373 (N_19373,N_19107,N_19071);
xor U19374 (N_19374,N_19033,N_19079);
xor U19375 (N_19375,N_19197,N_19087);
nand U19376 (N_19376,N_19015,N_19081);
xor U19377 (N_19377,N_19022,N_19080);
or U19378 (N_19378,N_19183,N_19099);
or U19379 (N_19379,N_19088,N_19135);
nand U19380 (N_19380,N_19102,N_19177);
nor U19381 (N_19381,N_19177,N_19072);
or U19382 (N_19382,N_19047,N_19173);
nor U19383 (N_19383,N_19021,N_19113);
nor U19384 (N_19384,N_19196,N_19026);
nor U19385 (N_19385,N_19120,N_19051);
nor U19386 (N_19386,N_19174,N_19197);
nor U19387 (N_19387,N_19100,N_19058);
xor U19388 (N_19388,N_19112,N_19187);
xor U19389 (N_19389,N_19067,N_19140);
nand U19390 (N_19390,N_19016,N_19161);
xor U19391 (N_19391,N_19088,N_19095);
nand U19392 (N_19392,N_19084,N_19063);
and U19393 (N_19393,N_19027,N_19174);
and U19394 (N_19394,N_19109,N_19062);
or U19395 (N_19395,N_19192,N_19148);
nor U19396 (N_19396,N_19038,N_19098);
and U19397 (N_19397,N_19155,N_19073);
xor U19398 (N_19398,N_19053,N_19127);
xnor U19399 (N_19399,N_19042,N_19056);
xnor U19400 (N_19400,N_19287,N_19312);
nand U19401 (N_19401,N_19371,N_19222);
xnor U19402 (N_19402,N_19214,N_19364);
nand U19403 (N_19403,N_19323,N_19201);
xor U19404 (N_19404,N_19205,N_19279);
nand U19405 (N_19405,N_19254,N_19224);
and U19406 (N_19406,N_19383,N_19392);
nand U19407 (N_19407,N_19345,N_19285);
xor U19408 (N_19408,N_19225,N_19235);
xor U19409 (N_19409,N_19342,N_19290);
nor U19410 (N_19410,N_19284,N_19256);
or U19411 (N_19411,N_19202,N_19221);
and U19412 (N_19412,N_19395,N_19275);
and U19413 (N_19413,N_19307,N_19367);
nand U19414 (N_19414,N_19289,N_19300);
and U19415 (N_19415,N_19396,N_19208);
and U19416 (N_19416,N_19231,N_19210);
nand U19417 (N_19417,N_19283,N_19369);
or U19418 (N_19418,N_19291,N_19313);
xor U19419 (N_19419,N_19380,N_19309);
nor U19420 (N_19420,N_19314,N_19232);
nand U19421 (N_19421,N_19237,N_19343);
or U19422 (N_19422,N_19244,N_19393);
nor U19423 (N_19423,N_19228,N_19213);
or U19424 (N_19424,N_19203,N_19271);
xnor U19425 (N_19425,N_19379,N_19250);
xnor U19426 (N_19426,N_19229,N_19247);
nor U19427 (N_19427,N_19305,N_19399);
or U19428 (N_19428,N_19292,N_19370);
nor U19429 (N_19429,N_19268,N_19324);
nor U19430 (N_19430,N_19373,N_19209);
or U19431 (N_19431,N_19260,N_19277);
xor U19432 (N_19432,N_19257,N_19385);
and U19433 (N_19433,N_19372,N_19328);
xor U19434 (N_19434,N_19263,N_19219);
and U19435 (N_19435,N_19234,N_19280);
or U19436 (N_19436,N_19262,N_19375);
or U19437 (N_19437,N_19365,N_19223);
and U19438 (N_19438,N_19286,N_19267);
nor U19439 (N_19439,N_19226,N_19363);
nand U19440 (N_19440,N_19391,N_19346);
nor U19441 (N_19441,N_19357,N_19252);
and U19442 (N_19442,N_19274,N_19243);
nor U19443 (N_19443,N_19282,N_19317);
nand U19444 (N_19444,N_19200,N_19242);
xnor U19445 (N_19445,N_19241,N_19227);
xor U19446 (N_19446,N_19264,N_19358);
xnor U19447 (N_19447,N_19337,N_19315);
and U19448 (N_19448,N_19297,N_19253);
xnor U19449 (N_19449,N_19356,N_19335);
nor U19450 (N_19450,N_19384,N_19390);
or U19451 (N_19451,N_19261,N_19397);
xor U19452 (N_19452,N_19293,N_19269);
nand U19453 (N_19453,N_19368,N_19398);
or U19454 (N_19454,N_19251,N_19249);
nor U19455 (N_19455,N_19296,N_19276);
nor U19456 (N_19456,N_19281,N_19361);
nand U19457 (N_19457,N_19360,N_19386);
or U19458 (N_19458,N_19327,N_19359);
and U19459 (N_19459,N_19374,N_19294);
nand U19460 (N_19460,N_19378,N_19388);
nand U19461 (N_19461,N_19216,N_19320);
xnor U19462 (N_19462,N_19303,N_19347);
and U19463 (N_19463,N_19206,N_19270);
nand U19464 (N_19464,N_19204,N_19349);
nand U19465 (N_19465,N_19353,N_19310);
or U19466 (N_19466,N_19322,N_19255);
xnor U19467 (N_19467,N_19248,N_19265);
and U19468 (N_19468,N_19332,N_19236);
xor U19469 (N_19469,N_19341,N_19319);
xnor U19470 (N_19470,N_19301,N_19304);
and U19471 (N_19471,N_19302,N_19215);
and U19472 (N_19472,N_19266,N_19207);
xor U19473 (N_19473,N_19258,N_19344);
nor U19474 (N_19474,N_19339,N_19218);
and U19475 (N_19475,N_19288,N_19212);
xor U19476 (N_19476,N_19362,N_19298);
or U19477 (N_19477,N_19352,N_19336);
nor U19478 (N_19478,N_19311,N_19299);
nor U19479 (N_19479,N_19382,N_19351);
nor U19480 (N_19480,N_19217,N_19338);
or U19481 (N_19481,N_19245,N_19389);
and U19482 (N_19482,N_19321,N_19238);
and U19483 (N_19483,N_19278,N_19259);
xor U19484 (N_19484,N_19220,N_19381);
and U19485 (N_19485,N_19334,N_19239);
or U19486 (N_19486,N_19330,N_19350);
nor U19487 (N_19487,N_19355,N_19333);
nor U19488 (N_19488,N_19211,N_19377);
or U19489 (N_19489,N_19295,N_19326);
and U19490 (N_19490,N_19348,N_19233);
nand U19491 (N_19491,N_19394,N_19246);
xor U19492 (N_19492,N_19272,N_19354);
xnor U19493 (N_19493,N_19308,N_19306);
xnor U19494 (N_19494,N_19230,N_19387);
nand U19495 (N_19495,N_19240,N_19318);
xnor U19496 (N_19496,N_19316,N_19329);
nand U19497 (N_19497,N_19273,N_19376);
nor U19498 (N_19498,N_19340,N_19331);
nand U19499 (N_19499,N_19366,N_19325);
or U19500 (N_19500,N_19340,N_19218);
xnor U19501 (N_19501,N_19288,N_19363);
and U19502 (N_19502,N_19351,N_19364);
and U19503 (N_19503,N_19399,N_19280);
nor U19504 (N_19504,N_19208,N_19369);
nor U19505 (N_19505,N_19306,N_19222);
and U19506 (N_19506,N_19268,N_19261);
and U19507 (N_19507,N_19350,N_19383);
xnor U19508 (N_19508,N_19341,N_19240);
xor U19509 (N_19509,N_19304,N_19261);
or U19510 (N_19510,N_19204,N_19338);
or U19511 (N_19511,N_19390,N_19338);
nand U19512 (N_19512,N_19250,N_19350);
and U19513 (N_19513,N_19355,N_19229);
nor U19514 (N_19514,N_19252,N_19335);
and U19515 (N_19515,N_19336,N_19230);
nor U19516 (N_19516,N_19245,N_19375);
xor U19517 (N_19517,N_19388,N_19368);
nand U19518 (N_19518,N_19280,N_19227);
xor U19519 (N_19519,N_19330,N_19288);
nor U19520 (N_19520,N_19209,N_19249);
nor U19521 (N_19521,N_19374,N_19236);
or U19522 (N_19522,N_19364,N_19251);
or U19523 (N_19523,N_19328,N_19359);
nand U19524 (N_19524,N_19344,N_19224);
or U19525 (N_19525,N_19359,N_19246);
nand U19526 (N_19526,N_19355,N_19349);
or U19527 (N_19527,N_19338,N_19328);
and U19528 (N_19528,N_19357,N_19308);
xnor U19529 (N_19529,N_19245,N_19235);
and U19530 (N_19530,N_19215,N_19337);
or U19531 (N_19531,N_19334,N_19217);
nand U19532 (N_19532,N_19358,N_19288);
and U19533 (N_19533,N_19299,N_19252);
nor U19534 (N_19534,N_19200,N_19260);
and U19535 (N_19535,N_19328,N_19203);
nand U19536 (N_19536,N_19278,N_19327);
or U19537 (N_19537,N_19345,N_19281);
nor U19538 (N_19538,N_19397,N_19211);
nand U19539 (N_19539,N_19270,N_19346);
or U19540 (N_19540,N_19338,N_19391);
xor U19541 (N_19541,N_19232,N_19219);
xnor U19542 (N_19542,N_19240,N_19268);
nand U19543 (N_19543,N_19259,N_19284);
and U19544 (N_19544,N_19255,N_19216);
xor U19545 (N_19545,N_19266,N_19344);
and U19546 (N_19546,N_19276,N_19218);
and U19547 (N_19547,N_19295,N_19373);
nor U19548 (N_19548,N_19248,N_19252);
or U19549 (N_19549,N_19237,N_19335);
or U19550 (N_19550,N_19392,N_19349);
nand U19551 (N_19551,N_19321,N_19265);
xnor U19552 (N_19552,N_19350,N_19355);
nand U19553 (N_19553,N_19342,N_19387);
and U19554 (N_19554,N_19255,N_19214);
and U19555 (N_19555,N_19217,N_19396);
and U19556 (N_19556,N_19362,N_19300);
nor U19557 (N_19557,N_19345,N_19377);
or U19558 (N_19558,N_19344,N_19306);
nor U19559 (N_19559,N_19269,N_19288);
xor U19560 (N_19560,N_19215,N_19351);
nor U19561 (N_19561,N_19380,N_19376);
nor U19562 (N_19562,N_19210,N_19225);
nand U19563 (N_19563,N_19259,N_19369);
nor U19564 (N_19564,N_19304,N_19298);
nor U19565 (N_19565,N_19397,N_19254);
or U19566 (N_19566,N_19209,N_19277);
and U19567 (N_19567,N_19324,N_19248);
xnor U19568 (N_19568,N_19382,N_19250);
or U19569 (N_19569,N_19230,N_19326);
nor U19570 (N_19570,N_19258,N_19225);
and U19571 (N_19571,N_19309,N_19298);
xor U19572 (N_19572,N_19268,N_19239);
nor U19573 (N_19573,N_19363,N_19371);
xnor U19574 (N_19574,N_19214,N_19305);
nand U19575 (N_19575,N_19217,N_19261);
nand U19576 (N_19576,N_19252,N_19238);
nor U19577 (N_19577,N_19265,N_19256);
or U19578 (N_19578,N_19341,N_19386);
or U19579 (N_19579,N_19235,N_19340);
nand U19580 (N_19580,N_19372,N_19252);
nor U19581 (N_19581,N_19301,N_19314);
or U19582 (N_19582,N_19348,N_19271);
and U19583 (N_19583,N_19311,N_19266);
or U19584 (N_19584,N_19306,N_19237);
xnor U19585 (N_19585,N_19270,N_19220);
and U19586 (N_19586,N_19269,N_19393);
and U19587 (N_19587,N_19264,N_19230);
nor U19588 (N_19588,N_19201,N_19384);
nor U19589 (N_19589,N_19339,N_19330);
nor U19590 (N_19590,N_19200,N_19287);
nor U19591 (N_19591,N_19342,N_19209);
and U19592 (N_19592,N_19315,N_19357);
nor U19593 (N_19593,N_19375,N_19331);
xor U19594 (N_19594,N_19314,N_19210);
or U19595 (N_19595,N_19388,N_19331);
nand U19596 (N_19596,N_19396,N_19210);
xor U19597 (N_19597,N_19375,N_19272);
and U19598 (N_19598,N_19382,N_19252);
nand U19599 (N_19599,N_19398,N_19268);
or U19600 (N_19600,N_19520,N_19470);
or U19601 (N_19601,N_19583,N_19566);
nand U19602 (N_19602,N_19533,N_19547);
or U19603 (N_19603,N_19413,N_19549);
or U19604 (N_19604,N_19429,N_19440);
and U19605 (N_19605,N_19585,N_19589);
or U19606 (N_19606,N_19419,N_19528);
xor U19607 (N_19607,N_19442,N_19456);
xor U19608 (N_19608,N_19510,N_19477);
nor U19609 (N_19609,N_19525,N_19410);
xor U19610 (N_19610,N_19581,N_19472);
nor U19611 (N_19611,N_19457,N_19481);
nand U19612 (N_19612,N_19513,N_19522);
or U19613 (N_19613,N_19479,N_19400);
xor U19614 (N_19614,N_19438,N_19582);
and U19615 (N_19615,N_19548,N_19455);
and U19616 (N_19616,N_19478,N_19441);
or U19617 (N_19617,N_19484,N_19565);
or U19618 (N_19618,N_19515,N_19524);
or U19619 (N_19619,N_19507,N_19437);
and U19620 (N_19620,N_19551,N_19532);
or U19621 (N_19621,N_19518,N_19444);
xor U19622 (N_19622,N_19468,N_19415);
and U19623 (N_19623,N_19490,N_19402);
nand U19624 (N_19624,N_19534,N_19414);
or U19625 (N_19625,N_19473,N_19476);
nand U19626 (N_19626,N_19516,N_19506);
nand U19627 (N_19627,N_19588,N_19469);
and U19628 (N_19628,N_19491,N_19480);
and U19629 (N_19629,N_19598,N_19521);
or U19630 (N_19630,N_19563,N_19475);
or U19631 (N_19631,N_19591,N_19462);
and U19632 (N_19632,N_19536,N_19535);
nand U19633 (N_19633,N_19540,N_19417);
nand U19634 (N_19634,N_19531,N_19500);
nor U19635 (N_19635,N_19492,N_19517);
or U19636 (N_19636,N_19488,N_19450);
xnor U19637 (N_19637,N_19504,N_19508);
and U19638 (N_19638,N_19554,N_19493);
nand U19639 (N_19639,N_19422,N_19505);
nand U19640 (N_19640,N_19543,N_19542);
nand U19641 (N_19641,N_19497,N_19486);
and U19642 (N_19642,N_19599,N_19575);
nand U19643 (N_19643,N_19502,N_19466);
nand U19644 (N_19644,N_19496,N_19436);
nand U19645 (N_19645,N_19460,N_19573);
xnor U19646 (N_19646,N_19593,N_19541);
or U19647 (N_19647,N_19538,N_19559);
nor U19648 (N_19648,N_19596,N_19576);
or U19649 (N_19649,N_19499,N_19537);
xnor U19650 (N_19650,N_19577,N_19403);
nand U19651 (N_19651,N_19430,N_19560);
nor U19652 (N_19652,N_19443,N_19580);
and U19653 (N_19653,N_19587,N_19544);
nand U19654 (N_19654,N_19571,N_19514);
and U19655 (N_19655,N_19574,N_19511);
or U19656 (N_19656,N_19449,N_19404);
and U19657 (N_19657,N_19446,N_19420);
or U19658 (N_19658,N_19451,N_19545);
nand U19659 (N_19659,N_19459,N_19586);
xor U19660 (N_19660,N_19495,N_19458);
and U19661 (N_19661,N_19552,N_19401);
nor U19662 (N_19662,N_19439,N_19423);
nor U19663 (N_19663,N_19546,N_19562);
nand U19664 (N_19664,N_19454,N_19595);
xor U19665 (N_19665,N_19426,N_19594);
xnor U19666 (N_19666,N_19526,N_19447);
or U19667 (N_19667,N_19408,N_19445);
or U19668 (N_19668,N_19570,N_19428);
nor U19669 (N_19669,N_19503,N_19501);
xnor U19670 (N_19670,N_19579,N_19561);
nand U19671 (N_19671,N_19523,N_19452);
xnor U19672 (N_19672,N_19569,N_19416);
nand U19673 (N_19673,N_19421,N_19409);
xnor U19674 (N_19674,N_19578,N_19572);
nand U19675 (N_19675,N_19530,N_19418);
or U19676 (N_19676,N_19461,N_19432);
and U19677 (N_19677,N_19467,N_19558);
nor U19678 (N_19678,N_19427,N_19550);
xor U19679 (N_19679,N_19555,N_19568);
and U19680 (N_19680,N_19498,N_19494);
xnor U19681 (N_19681,N_19471,N_19509);
or U19682 (N_19682,N_19406,N_19519);
nor U19683 (N_19683,N_19405,N_19590);
nor U19684 (N_19684,N_19407,N_19485);
nor U19685 (N_19685,N_19556,N_19527);
nor U19686 (N_19686,N_19539,N_19564);
or U19687 (N_19687,N_19425,N_19584);
or U19688 (N_19688,N_19448,N_19483);
or U19689 (N_19689,N_19592,N_19431);
nor U19690 (N_19690,N_19435,N_19465);
and U19691 (N_19691,N_19434,N_19412);
and U19692 (N_19692,N_19487,N_19557);
nand U19693 (N_19693,N_19512,N_19567);
nor U19694 (N_19694,N_19433,N_19529);
and U19695 (N_19695,N_19463,N_19482);
and U19696 (N_19696,N_19424,N_19411);
and U19697 (N_19697,N_19597,N_19489);
nor U19698 (N_19698,N_19453,N_19474);
or U19699 (N_19699,N_19553,N_19464);
or U19700 (N_19700,N_19426,N_19556);
nor U19701 (N_19701,N_19403,N_19592);
nand U19702 (N_19702,N_19431,N_19453);
xnor U19703 (N_19703,N_19596,N_19520);
nand U19704 (N_19704,N_19500,N_19476);
nand U19705 (N_19705,N_19452,N_19426);
xor U19706 (N_19706,N_19546,N_19466);
and U19707 (N_19707,N_19569,N_19581);
and U19708 (N_19708,N_19517,N_19580);
xnor U19709 (N_19709,N_19444,N_19595);
nor U19710 (N_19710,N_19516,N_19450);
and U19711 (N_19711,N_19596,N_19571);
xnor U19712 (N_19712,N_19446,N_19449);
nand U19713 (N_19713,N_19544,N_19425);
and U19714 (N_19714,N_19579,N_19482);
nor U19715 (N_19715,N_19527,N_19594);
xor U19716 (N_19716,N_19500,N_19432);
nand U19717 (N_19717,N_19523,N_19513);
xor U19718 (N_19718,N_19462,N_19470);
nor U19719 (N_19719,N_19534,N_19404);
and U19720 (N_19720,N_19476,N_19467);
nor U19721 (N_19721,N_19537,N_19425);
nor U19722 (N_19722,N_19583,N_19537);
nand U19723 (N_19723,N_19554,N_19423);
nor U19724 (N_19724,N_19489,N_19450);
or U19725 (N_19725,N_19430,N_19459);
xor U19726 (N_19726,N_19589,N_19488);
and U19727 (N_19727,N_19436,N_19520);
and U19728 (N_19728,N_19515,N_19453);
xor U19729 (N_19729,N_19585,N_19465);
nor U19730 (N_19730,N_19550,N_19480);
nor U19731 (N_19731,N_19568,N_19407);
nor U19732 (N_19732,N_19429,N_19567);
or U19733 (N_19733,N_19510,N_19503);
nor U19734 (N_19734,N_19534,N_19562);
nand U19735 (N_19735,N_19538,N_19418);
nand U19736 (N_19736,N_19460,N_19411);
nor U19737 (N_19737,N_19578,N_19559);
nand U19738 (N_19738,N_19454,N_19438);
nor U19739 (N_19739,N_19568,N_19530);
xnor U19740 (N_19740,N_19537,N_19475);
nand U19741 (N_19741,N_19490,N_19515);
and U19742 (N_19742,N_19418,N_19445);
nand U19743 (N_19743,N_19523,N_19586);
nor U19744 (N_19744,N_19458,N_19567);
nand U19745 (N_19745,N_19584,N_19509);
nor U19746 (N_19746,N_19496,N_19501);
and U19747 (N_19747,N_19505,N_19502);
or U19748 (N_19748,N_19546,N_19523);
and U19749 (N_19749,N_19511,N_19599);
nor U19750 (N_19750,N_19499,N_19415);
and U19751 (N_19751,N_19528,N_19476);
and U19752 (N_19752,N_19542,N_19569);
and U19753 (N_19753,N_19599,N_19547);
nand U19754 (N_19754,N_19537,N_19547);
and U19755 (N_19755,N_19527,N_19427);
nor U19756 (N_19756,N_19419,N_19420);
nor U19757 (N_19757,N_19502,N_19511);
nor U19758 (N_19758,N_19439,N_19502);
xor U19759 (N_19759,N_19549,N_19449);
nor U19760 (N_19760,N_19469,N_19459);
nor U19761 (N_19761,N_19590,N_19472);
xnor U19762 (N_19762,N_19567,N_19409);
or U19763 (N_19763,N_19564,N_19506);
and U19764 (N_19764,N_19573,N_19474);
and U19765 (N_19765,N_19481,N_19402);
nor U19766 (N_19766,N_19443,N_19474);
and U19767 (N_19767,N_19400,N_19511);
xor U19768 (N_19768,N_19427,N_19424);
xnor U19769 (N_19769,N_19460,N_19544);
nand U19770 (N_19770,N_19479,N_19528);
nor U19771 (N_19771,N_19577,N_19408);
nor U19772 (N_19772,N_19457,N_19419);
and U19773 (N_19773,N_19418,N_19484);
nor U19774 (N_19774,N_19425,N_19559);
nor U19775 (N_19775,N_19463,N_19574);
xor U19776 (N_19776,N_19547,N_19485);
and U19777 (N_19777,N_19472,N_19597);
or U19778 (N_19778,N_19407,N_19582);
and U19779 (N_19779,N_19414,N_19419);
nor U19780 (N_19780,N_19542,N_19433);
or U19781 (N_19781,N_19584,N_19545);
nor U19782 (N_19782,N_19570,N_19496);
xor U19783 (N_19783,N_19596,N_19588);
nor U19784 (N_19784,N_19529,N_19545);
nand U19785 (N_19785,N_19452,N_19532);
and U19786 (N_19786,N_19484,N_19496);
and U19787 (N_19787,N_19532,N_19478);
nand U19788 (N_19788,N_19440,N_19586);
and U19789 (N_19789,N_19489,N_19471);
or U19790 (N_19790,N_19570,N_19525);
nand U19791 (N_19791,N_19543,N_19423);
nand U19792 (N_19792,N_19566,N_19530);
or U19793 (N_19793,N_19494,N_19499);
nor U19794 (N_19794,N_19510,N_19401);
nand U19795 (N_19795,N_19418,N_19453);
and U19796 (N_19796,N_19438,N_19526);
or U19797 (N_19797,N_19408,N_19549);
and U19798 (N_19798,N_19536,N_19509);
and U19799 (N_19799,N_19422,N_19423);
and U19800 (N_19800,N_19696,N_19681);
nor U19801 (N_19801,N_19632,N_19634);
or U19802 (N_19802,N_19617,N_19780);
nor U19803 (N_19803,N_19788,N_19714);
xnor U19804 (N_19804,N_19642,N_19736);
nand U19805 (N_19805,N_19633,N_19742);
or U19806 (N_19806,N_19740,N_19691);
and U19807 (N_19807,N_19627,N_19741);
or U19808 (N_19808,N_19684,N_19675);
and U19809 (N_19809,N_19783,N_19699);
or U19810 (N_19810,N_19784,N_19777);
or U19811 (N_19811,N_19618,N_19694);
xnor U19812 (N_19812,N_19720,N_19762);
nand U19813 (N_19813,N_19707,N_19797);
xor U19814 (N_19814,N_19705,N_19790);
nor U19815 (N_19815,N_19725,N_19671);
nand U19816 (N_19816,N_19676,N_19735);
nor U19817 (N_19817,N_19654,N_19674);
and U19818 (N_19818,N_19731,N_19653);
and U19819 (N_19819,N_19704,N_19739);
nor U19820 (N_19820,N_19737,N_19635);
nand U19821 (N_19821,N_19779,N_19668);
nor U19822 (N_19822,N_19649,N_19610);
xor U19823 (N_19823,N_19764,N_19672);
or U19824 (N_19824,N_19716,N_19601);
nor U19825 (N_19825,N_19785,N_19636);
xnor U19826 (N_19826,N_19662,N_19756);
xor U19827 (N_19827,N_19670,N_19752);
nand U19828 (N_19828,N_19757,N_19614);
nand U19829 (N_19829,N_19769,N_19693);
and U19830 (N_19830,N_19746,N_19792);
nor U19831 (N_19831,N_19755,N_19713);
xnor U19832 (N_19832,N_19639,N_19602);
and U19833 (N_19833,N_19648,N_19774);
xor U19834 (N_19834,N_19603,N_19655);
nand U19835 (N_19835,N_19629,N_19787);
nor U19836 (N_19836,N_19759,N_19724);
and U19837 (N_19837,N_19747,N_19703);
nor U19838 (N_19838,N_19753,N_19718);
xnor U19839 (N_19839,N_19700,N_19600);
xor U19840 (N_19840,N_19721,N_19715);
nand U19841 (N_19841,N_19607,N_19640);
xor U19842 (N_19842,N_19750,N_19651);
or U19843 (N_19843,N_19701,N_19658);
or U19844 (N_19844,N_19767,N_19604);
nand U19845 (N_19845,N_19786,N_19766);
and U19846 (N_19846,N_19719,N_19773);
or U19847 (N_19847,N_19761,N_19734);
nand U19848 (N_19848,N_19758,N_19744);
nor U19849 (N_19849,N_19677,N_19789);
xor U19850 (N_19850,N_19717,N_19637);
or U19851 (N_19851,N_19765,N_19667);
nand U19852 (N_19852,N_19751,N_19605);
xor U19853 (N_19853,N_19771,N_19791);
nand U19854 (N_19854,N_19729,N_19619);
and U19855 (N_19855,N_19659,N_19775);
nor U19856 (N_19856,N_19664,N_19624);
xnor U19857 (N_19857,N_19623,N_19683);
nor U19858 (N_19858,N_19690,N_19692);
or U19859 (N_19859,N_19781,N_19772);
and U19860 (N_19860,N_19641,N_19666);
nor U19861 (N_19861,N_19776,N_19680);
xor U19862 (N_19862,N_19687,N_19673);
nor U19863 (N_19863,N_19743,N_19749);
nor U19864 (N_19864,N_19625,N_19616);
or U19865 (N_19865,N_19768,N_19613);
nor U19866 (N_19866,N_19795,N_19685);
nand U19867 (N_19867,N_19622,N_19621);
nand U19868 (N_19868,N_19709,N_19799);
and U19869 (N_19869,N_19615,N_19794);
nor U19870 (N_19870,N_19712,N_19708);
nor U19871 (N_19871,N_19727,N_19643);
nand U19872 (N_19872,N_19723,N_19732);
or U19873 (N_19873,N_19660,N_19650);
nor U19874 (N_19874,N_19611,N_19688);
and U19875 (N_19875,N_19733,N_19682);
nor U19876 (N_19876,N_19652,N_19665);
nor U19877 (N_19877,N_19745,N_19695);
nand U19878 (N_19878,N_19728,N_19798);
xor U19879 (N_19879,N_19628,N_19738);
nor U19880 (N_19880,N_19644,N_19697);
nor U19881 (N_19881,N_19706,N_19631);
or U19882 (N_19882,N_19645,N_19661);
nand U19883 (N_19883,N_19698,N_19770);
or U19884 (N_19884,N_19657,N_19748);
xnor U19885 (N_19885,N_19612,N_19702);
or U19886 (N_19886,N_19710,N_19793);
nand U19887 (N_19887,N_19726,N_19646);
nor U19888 (N_19888,N_19778,N_19730);
xnor U19889 (N_19889,N_19796,N_19647);
nor U19890 (N_19890,N_19669,N_19760);
nor U19891 (N_19891,N_19626,N_19663);
or U19892 (N_19892,N_19722,N_19620);
xor U19893 (N_19893,N_19608,N_19606);
nor U19894 (N_19894,N_19686,N_19630);
nor U19895 (N_19895,N_19763,N_19679);
and U19896 (N_19896,N_19711,N_19754);
or U19897 (N_19897,N_19638,N_19678);
nand U19898 (N_19898,N_19689,N_19656);
and U19899 (N_19899,N_19782,N_19609);
or U19900 (N_19900,N_19794,N_19700);
nor U19901 (N_19901,N_19631,N_19774);
nand U19902 (N_19902,N_19777,N_19620);
or U19903 (N_19903,N_19678,N_19641);
xnor U19904 (N_19904,N_19675,N_19657);
xnor U19905 (N_19905,N_19652,N_19606);
and U19906 (N_19906,N_19659,N_19611);
and U19907 (N_19907,N_19615,N_19629);
nor U19908 (N_19908,N_19625,N_19760);
xor U19909 (N_19909,N_19682,N_19779);
nand U19910 (N_19910,N_19671,N_19653);
xor U19911 (N_19911,N_19671,N_19656);
xor U19912 (N_19912,N_19650,N_19719);
or U19913 (N_19913,N_19795,N_19646);
or U19914 (N_19914,N_19699,N_19628);
nor U19915 (N_19915,N_19701,N_19783);
nand U19916 (N_19916,N_19676,N_19689);
and U19917 (N_19917,N_19624,N_19646);
xor U19918 (N_19918,N_19608,N_19761);
nor U19919 (N_19919,N_19625,N_19709);
xnor U19920 (N_19920,N_19697,N_19604);
nand U19921 (N_19921,N_19747,N_19700);
and U19922 (N_19922,N_19712,N_19633);
and U19923 (N_19923,N_19616,N_19663);
nor U19924 (N_19924,N_19633,N_19607);
nor U19925 (N_19925,N_19722,N_19717);
or U19926 (N_19926,N_19660,N_19651);
nand U19927 (N_19927,N_19671,N_19651);
nand U19928 (N_19928,N_19670,N_19720);
xnor U19929 (N_19929,N_19645,N_19660);
xnor U19930 (N_19930,N_19711,N_19792);
and U19931 (N_19931,N_19622,N_19736);
nand U19932 (N_19932,N_19706,N_19607);
nor U19933 (N_19933,N_19737,N_19601);
or U19934 (N_19934,N_19760,N_19667);
and U19935 (N_19935,N_19732,N_19683);
or U19936 (N_19936,N_19635,N_19665);
nand U19937 (N_19937,N_19782,N_19716);
or U19938 (N_19938,N_19690,N_19651);
or U19939 (N_19939,N_19744,N_19701);
and U19940 (N_19940,N_19714,N_19733);
nand U19941 (N_19941,N_19601,N_19741);
xnor U19942 (N_19942,N_19778,N_19741);
or U19943 (N_19943,N_19755,N_19693);
and U19944 (N_19944,N_19700,N_19758);
or U19945 (N_19945,N_19629,N_19642);
and U19946 (N_19946,N_19685,N_19701);
nor U19947 (N_19947,N_19662,N_19761);
or U19948 (N_19948,N_19799,N_19789);
or U19949 (N_19949,N_19608,N_19700);
xnor U19950 (N_19950,N_19666,N_19631);
xnor U19951 (N_19951,N_19779,N_19746);
or U19952 (N_19952,N_19753,N_19765);
xnor U19953 (N_19953,N_19693,N_19732);
or U19954 (N_19954,N_19709,N_19635);
or U19955 (N_19955,N_19603,N_19606);
nor U19956 (N_19956,N_19608,N_19738);
or U19957 (N_19957,N_19698,N_19694);
nor U19958 (N_19958,N_19736,N_19603);
or U19959 (N_19959,N_19799,N_19663);
nor U19960 (N_19960,N_19680,N_19686);
nor U19961 (N_19961,N_19632,N_19611);
and U19962 (N_19962,N_19726,N_19752);
and U19963 (N_19963,N_19746,N_19754);
xnor U19964 (N_19964,N_19731,N_19606);
nand U19965 (N_19965,N_19746,N_19695);
nor U19966 (N_19966,N_19715,N_19682);
and U19967 (N_19967,N_19658,N_19763);
xnor U19968 (N_19968,N_19741,N_19725);
xor U19969 (N_19969,N_19791,N_19657);
nand U19970 (N_19970,N_19788,N_19626);
or U19971 (N_19971,N_19711,N_19702);
and U19972 (N_19972,N_19615,N_19770);
or U19973 (N_19973,N_19700,N_19739);
nor U19974 (N_19974,N_19725,N_19780);
nand U19975 (N_19975,N_19651,N_19723);
or U19976 (N_19976,N_19637,N_19636);
nor U19977 (N_19977,N_19634,N_19722);
nor U19978 (N_19978,N_19774,N_19640);
nand U19979 (N_19979,N_19749,N_19745);
and U19980 (N_19980,N_19678,N_19751);
and U19981 (N_19981,N_19746,N_19644);
nor U19982 (N_19982,N_19634,N_19693);
nand U19983 (N_19983,N_19667,N_19731);
nand U19984 (N_19984,N_19660,N_19642);
nand U19985 (N_19985,N_19721,N_19669);
xnor U19986 (N_19986,N_19679,N_19782);
or U19987 (N_19987,N_19734,N_19639);
and U19988 (N_19988,N_19661,N_19742);
and U19989 (N_19989,N_19683,N_19676);
or U19990 (N_19990,N_19603,N_19775);
nand U19991 (N_19991,N_19614,N_19720);
nand U19992 (N_19992,N_19737,N_19651);
xnor U19993 (N_19993,N_19626,N_19667);
and U19994 (N_19994,N_19637,N_19778);
xor U19995 (N_19995,N_19692,N_19792);
or U19996 (N_19996,N_19681,N_19758);
or U19997 (N_19997,N_19647,N_19723);
and U19998 (N_19998,N_19650,N_19708);
nor U19999 (N_19999,N_19707,N_19769);
and UO_0 (O_0,N_19956,N_19979);
nor UO_1 (O_1,N_19854,N_19968);
nor UO_2 (O_2,N_19865,N_19939);
or UO_3 (O_3,N_19924,N_19872);
and UO_4 (O_4,N_19955,N_19947);
nor UO_5 (O_5,N_19990,N_19839);
nor UO_6 (O_6,N_19893,N_19934);
or UO_7 (O_7,N_19940,N_19927);
or UO_8 (O_8,N_19988,N_19842);
xor UO_9 (O_9,N_19853,N_19830);
xnor UO_10 (O_10,N_19961,N_19954);
and UO_11 (O_11,N_19910,N_19944);
nor UO_12 (O_12,N_19963,N_19846);
or UO_13 (O_13,N_19884,N_19804);
or UO_14 (O_14,N_19829,N_19819);
or UO_15 (O_15,N_19802,N_19848);
xnor UO_16 (O_16,N_19908,N_19953);
or UO_17 (O_17,N_19827,N_19887);
or UO_18 (O_18,N_19816,N_19815);
and UO_19 (O_19,N_19952,N_19950);
and UO_20 (O_20,N_19964,N_19957);
nor UO_21 (O_21,N_19824,N_19917);
or UO_22 (O_22,N_19946,N_19851);
or UO_23 (O_23,N_19981,N_19805);
or UO_24 (O_24,N_19862,N_19828);
nand UO_25 (O_25,N_19921,N_19926);
nand UO_26 (O_26,N_19883,N_19810);
or UO_27 (O_27,N_19850,N_19896);
nor UO_28 (O_28,N_19903,N_19969);
or UO_29 (O_29,N_19911,N_19881);
nand UO_30 (O_30,N_19831,N_19876);
and UO_31 (O_31,N_19864,N_19959);
nand UO_32 (O_32,N_19966,N_19977);
and UO_33 (O_33,N_19832,N_19936);
xor UO_34 (O_34,N_19965,N_19880);
and UO_35 (O_35,N_19877,N_19840);
and UO_36 (O_36,N_19995,N_19945);
nor UO_37 (O_37,N_19942,N_19837);
nand UO_38 (O_38,N_19986,N_19971);
nor UO_39 (O_39,N_19897,N_19807);
and UO_40 (O_40,N_19879,N_19998);
or UO_41 (O_41,N_19809,N_19992);
nor UO_42 (O_42,N_19937,N_19803);
or UO_43 (O_43,N_19889,N_19976);
or UO_44 (O_44,N_19991,N_19980);
or UO_45 (O_45,N_19800,N_19983);
xnor UO_46 (O_46,N_19873,N_19808);
nand UO_47 (O_47,N_19820,N_19861);
nand UO_48 (O_48,N_19962,N_19907);
or UO_49 (O_49,N_19943,N_19974);
xnor UO_50 (O_50,N_19929,N_19886);
and UO_51 (O_51,N_19882,N_19823);
and UO_52 (O_52,N_19948,N_19875);
and UO_53 (O_53,N_19960,N_19817);
and UO_54 (O_54,N_19989,N_19899);
xor UO_55 (O_55,N_19930,N_19871);
nor UO_56 (O_56,N_19825,N_19931);
or UO_57 (O_57,N_19890,N_19868);
nor UO_58 (O_58,N_19985,N_19993);
xnor UO_59 (O_59,N_19812,N_19860);
nor UO_60 (O_60,N_19863,N_19814);
or UO_61 (O_61,N_19847,N_19938);
nand UO_62 (O_62,N_19925,N_19919);
nor UO_63 (O_63,N_19958,N_19826);
or UO_64 (O_64,N_19999,N_19904);
xor UO_65 (O_65,N_19866,N_19973);
or UO_66 (O_66,N_19836,N_19898);
or UO_67 (O_67,N_19894,N_19935);
nor UO_68 (O_68,N_19891,N_19902);
nand UO_69 (O_69,N_19801,N_19916);
and UO_70 (O_70,N_19834,N_19909);
xnor UO_71 (O_71,N_19841,N_19813);
nand UO_72 (O_72,N_19970,N_19845);
nand UO_73 (O_73,N_19835,N_19994);
xnor UO_74 (O_74,N_19849,N_19913);
and UO_75 (O_75,N_19912,N_19982);
or UO_76 (O_76,N_19878,N_19895);
nand UO_77 (O_77,N_19905,N_19967);
and UO_78 (O_78,N_19806,N_19858);
xnor UO_79 (O_79,N_19838,N_19918);
nand UO_80 (O_80,N_19811,N_19885);
xnor UO_81 (O_81,N_19933,N_19843);
and UO_82 (O_82,N_19888,N_19874);
and UO_83 (O_83,N_19941,N_19928);
nand UO_84 (O_84,N_19857,N_19869);
xnor UO_85 (O_85,N_19920,N_19900);
nor UO_86 (O_86,N_19923,N_19972);
nor UO_87 (O_87,N_19996,N_19922);
nor UO_88 (O_88,N_19867,N_19987);
nor UO_89 (O_89,N_19901,N_19852);
and UO_90 (O_90,N_19951,N_19833);
xor UO_91 (O_91,N_19949,N_19844);
nand UO_92 (O_92,N_19915,N_19821);
xnor UO_93 (O_93,N_19822,N_19818);
and UO_94 (O_94,N_19856,N_19914);
nor UO_95 (O_95,N_19975,N_19978);
nor UO_96 (O_96,N_19892,N_19997);
nand UO_97 (O_97,N_19932,N_19906);
and UO_98 (O_98,N_19859,N_19870);
nand UO_99 (O_99,N_19855,N_19984);
nand UO_100 (O_100,N_19945,N_19895);
or UO_101 (O_101,N_19845,N_19928);
or UO_102 (O_102,N_19859,N_19898);
nor UO_103 (O_103,N_19821,N_19831);
xnor UO_104 (O_104,N_19809,N_19843);
or UO_105 (O_105,N_19836,N_19925);
xnor UO_106 (O_106,N_19999,N_19984);
nor UO_107 (O_107,N_19953,N_19880);
xor UO_108 (O_108,N_19866,N_19913);
xor UO_109 (O_109,N_19867,N_19805);
or UO_110 (O_110,N_19906,N_19918);
nand UO_111 (O_111,N_19816,N_19827);
nor UO_112 (O_112,N_19931,N_19972);
and UO_113 (O_113,N_19880,N_19958);
xnor UO_114 (O_114,N_19826,N_19857);
xnor UO_115 (O_115,N_19906,N_19804);
and UO_116 (O_116,N_19853,N_19998);
nor UO_117 (O_117,N_19993,N_19921);
or UO_118 (O_118,N_19981,N_19837);
xnor UO_119 (O_119,N_19868,N_19983);
and UO_120 (O_120,N_19806,N_19866);
or UO_121 (O_121,N_19814,N_19852);
nand UO_122 (O_122,N_19933,N_19847);
nor UO_123 (O_123,N_19960,N_19875);
or UO_124 (O_124,N_19900,N_19908);
or UO_125 (O_125,N_19819,N_19901);
nand UO_126 (O_126,N_19805,N_19952);
or UO_127 (O_127,N_19841,N_19890);
or UO_128 (O_128,N_19839,N_19918);
xor UO_129 (O_129,N_19845,N_19889);
xnor UO_130 (O_130,N_19980,N_19815);
nor UO_131 (O_131,N_19856,N_19930);
or UO_132 (O_132,N_19931,N_19927);
and UO_133 (O_133,N_19862,N_19845);
nor UO_134 (O_134,N_19957,N_19914);
nor UO_135 (O_135,N_19960,N_19958);
nand UO_136 (O_136,N_19820,N_19868);
and UO_137 (O_137,N_19866,N_19938);
nand UO_138 (O_138,N_19894,N_19866);
or UO_139 (O_139,N_19817,N_19830);
and UO_140 (O_140,N_19955,N_19814);
xnor UO_141 (O_141,N_19906,N_19902);
and UO_142 (O_142,N_19814,N_19827);
and UO_143 (O_143,N_19951,N_19873);
nor UO_144 (O_144,N_19928,N_19919);
xnor UO_145 (O_145,N_19946,N_19856);
or UO_146 (O_146,N_19925,N_19962);
and UO_147 (O_147,N_19992,N_19861);
xnor UO_148 (O_148,N_19985,N_19829);
nor UO_149 (O_149,N_19877,N_19938);
nor UO_150 (O_150,N_19845,N_19909);
nand UO_151 (O_151,N_19974,N_19930);
and UO_152 (O_152,N_19983,N_19919);
nor UO_153 (O_153,N_19892,N_19889);
or UO_154 (O_154,N_19968,N_19847);
xor UO_155 (O_155,N_19893,N_19864);
or UO_156 (O_156,N_19874,N_19934);
nand UO_157 (O_157,N_19844,N_19993);
nand UO_158 (O_158,N_19959,N_19983);
and UO_159 (O_159,N_19993,N_19949);
nor UO_160 (O_160,N_19882,N_19843);
or UO_161 (O_161,N_19948,N_19842);
nor UO_162 (O_162,N_19820,N_19803);
nor UO_163 (O_163,N_19845,N_19999);
xnor UO_164 (O_164,N_19825,N_19834);
nand UO_165 (O_165,N_19864,N_19912);
and UO_166 (O_166,N_19853,N_19903);
xor UO_167 (O_167,N_19918,N_19972);
nor UO_168 (O_168,N_19828,N_19925);
xnor UO_169 (O_169,N_19812,N_19853);
and UO_170 (O_170,N_19996,N_19883);
nor UO_171 (O_171,N_19961,N_19957);
nor UO_172 (O_172,N_19831,N_19906);
or UO_173 (O_173,N_19966,N_19859);
xnor UO_174 (O_174,N_19901,N_19982);
nand UO_175 (O_175,N_19929,N_19835);
or UO_176 (O_176,N_19904,N_19822);
xnor UO_177 (O_177,N_19856,N_19876);
or UO_178 (O_178,N_19930,N_19903);
xnor UO_179 (O_179,N_19987,N_19980);
xnor UO_180 (O_180,N_19969,N_19834);
nand UO_181 (O_181,N_19899,N_19863);
xnor UO_182 (O_182,N_19973,N_19888);
and UO_183 (O_183,N_19939,N_19977);
nor UO_184 (O_184,N_19849,N_19914);
nor UO_185 (O_185,N_19854,N_19904);
nor UO_186 (O_186,N_19827,N_19931);
and UO_187 (O_187,N_19974,N_19917);
xor UO_188 (O_188,N_19860,N_19938);
and UO_189 (O_189,N_19991,N_19998);
nand UO_190 (O_190,N_19973,N_19850);
or UO_191 (O_191,N_19835,N_19951);
nand UO_192 (O_192,N_19903,N_19914);
or UO_193 (O_193,N_19989,N_19851);
xnor UO_194 (O_194,N_19939,N_19829);
xnor UO_195 (O_195,N_19870,N_19924);
and UO_196 (O_196,N_19828,N_19839);
xor UO_197 (O_197,N_19982,N_19880);
nor UO_198 (O_198,N_19872,N_19987);
and UO_199 (O_199,N_19862,N_19995);
or UO_200 (O_200,N_19905,N_19856);
xor UO_201 (O_201,N_19931,N_19943);
and UO_202 (O_202,N_19872,N_19920);
nor UO_203 (O_203,N_19847,N_19854);
or UO_204 (O_204,N_19881,N_19833);
xnor UO_205 (O_205,N_19855,N_19922);
and UO_206 (O_206,N_19891,N_19941);
and UO_207 (O_207,N_19814,N_19824);
and UO_208 (O_208,N_19807,N_19842);
nand UO_209 (O_209,N_19980,N_19994);
and UO_210 (O_210,N_19905,N_19808);
nor UO_211 (O_211,N_19988,N_19992);
xnor UO_212 (O_212,N_19984,N_19983);
xnor UO_213 (O_213,N_19920,N_19851);
and UO_214 (O_214,N_19817,N_19959);
or UO_215 (O_215,N_19907,N_19867);
xor UO_216 (O_216,N_19826,N_19999);
or UO_217 (O_217,N_19900,N_19845);
xor UO_218 (O_218,N_19870,N_19821);
or UO_219 (O_219,N_19918,N_19934);
or UO_220 (O_220,N_19944,N_19879);
xor UO_221 (O_221,N_19936,N_19943);
nor UO_222 (O_222,N_19925,N_19939);
nor UO_223 (O_223,N_19811,N_19940);
or UO_224 (O_224,N_19908,N_19804);
or UO_225 (O_225,N_19985,N_19947);
nor UO_226 (O_226,N_19878,N_19820);
and UO_227 (O_227,N_19868,N_19949);
xnor UO_228 (O_228,N_19870,N_19998);
nor UO_229 (O_229,N_19983,N_19944);
nor UO_230 (O_230,N_19980,N_19849);
nor UO_231 (O_231,N_19832,N_19969);
nand UO_232 (O_232,N_19909,N_19981);
and UO_233 (O_233,N_19894,N_19837);
and UO_234 (O_234,N_19988,N_19821);
and UO_235 (O_235,N_19911,N_19809);
nor UO_236 (O_236,N_19939,N_19839);
and UO_237 (O_237,N_19803,N_19947);
nor UO_238 (O_238,N_19981,N_19999);
and UO_239 (O_239,N_19947,N_19861);
or UO_240 (O_240,N_19927,N_19989);
xnor UO_241 (O_241,N_19952,N_19973);
xor UO_242 (O_242,N_19906,N_19861);
xor UO_243 (O_243,N_19931,N_19966);
or UO_244 (O_244,N_19873,N_19890);
and UO_245 (O_245,N_19877,N_19904);
xor UO_246 (O_246,N_19813,N_19858);
xor UO_247 (O_247,N_19964,N_19916);
nor UO_248 (O_248,N_19836,N_19860);
and UO_249 (O_249,N_19821,N_19839);
nor UO_250 (O_250,N_19856,N_19916);
xor UO_251 (O_251,N_19898,N_19967);
xnor UO_252 (O_252,N_19837,N_19877);
nand UO_253 (O_253,N_19834,N_19963);
nor UO_254 (O_254,N_19897,N_19969);
or UO_255 (O_255,N_19826,N_19802);
or UO_256 (O_256,N_19886,N_19969);
xnor UO_257 (O_257,N_19857,N_19911);
nor UO_258 (O_258,N_19845,N_19947);
nor UO_259 (O_259,N_19885,N_19809);
nand UO_260 (O_260,N_19927,N_19819);
and UO_261 (O_261,N_19904,N_19865);
or UO_262 (O_262,N_19974,N_19978);
xor UO_263 (O_263,N_19935,N_19940);
and UO_264 (O_264,N_19911,N_19878);
and UO_265 (O_265,N_19826,N_19913);
xor UO_266 (O_266,N_19881,N_19850);
nand UO_267 (O_267,N_19926,N_19876);
nand UO_268 (O_268,N_19985,N_19977);
nand UO_269 (O_269,N_19998,N_19946);
and UO_270 (O_270,N_19891,N_19844);
xnor UO_271 (O_271,N_19806,N_19860);
and UO_272 (O_272,N_19942,N_19823);
or UO_273 (O_273,N_19898,N_19869);
xor UO_274 (O_274,N_19846,N_19900);
xor UO_275 (O_275,N_19965,N_19991);
nor UO_276 (O_276,N_19854,N_19810);
and UO_277 (O_277,N_19803,N_19905);
xnor UO_278 (O_278,N_19822,N_19938);
nand UO_279 (O_279,N_19998,N_19932);
xnor UO_280 (O_280,N_19917,N_19994);
and UO_281 (O_281,N_19815,N_19996);
or UO_282 (O_282,N_19905,N_19879);
and UO_283 (O_283,N_19896,N_19839);
nor UO_284 (O_284,N_19818,N_19976);
xor UO_285 (O_285,N_19838,N_19926);
nor UO_286 (O_286,N_19964,N_19917);
and UO_287 (O_287,N_19999,N_19895);
or UO_288 (O_288,N_19907,N_19862);
nor UO_289 (O_289,N_19825,N_19999);
xor UO_290 (O_290,N_19884,N_19963);
and UO_291 (O_291,N_19859,N_19809);
nand UO_292 (O_292,N_19902,N_19848);
nand UO_293 (O_293,N_19803,N_19977);
or UO_294 (O_294,N_19827,N_19940);
xnor UO_295 (O_295,N_19988,N_19935);
nor UO_296 (O_296,N_19927,N_19920);
nor UO_297 (O_297,N_19866,N_19979);
nand UO_298 (O_298,N_19956,N_19952);
nor UO_299 (O_299,N_19982,N_19807);
nor UO_300 (O_300,N_19846,N_19940);
nand UO_301 (O_301,N_19977,N_19940);
or UO_302 (O_302,N_19999,N_19839);
xnor UO_303 (O_303,N_19972,N_19810);
nand UO_304 (O_304,N_19847,N_19921);
or UO_305 (O_305,N_19952,N_19967);
and UO_306 (O_306,N_19847,N_19899);
nand UO_307 (O_307,N_19901,N_19958);
and UO_308 (O_308,N_19925,N_19931);
and UO_309 (O_309,N_19855,N_19977);
nand UO_310 (O_310,N_19826,N_19902);
and UO_311 (O_311,N_19965,N_19886);
and UO_312 (O_312,N_19939,N_19927);
or UO_313 (O_313,N_19809,N_19916);
xor UO_314 (O_314,N_19948,N_19965);
and UO_315 (O_315,N_19801,N_19878);
or UO_316 (O_316,N_19903,N_19887);
xor UO_317 (O_317,N_19870,N_19908);
or UO_318 (O_318,N_19907,N_19932);
xnor UO_319 (O_319,N_19824,N_19909);
xnor UO_320 (O_320,N_19845,N_19878);
or UO_321 (O_321,N_19941,N_19816);
nor UO_322 (O_322,N_19954,N_19977);
nor UO_323 (O_323,N_19945,N_19803);
nand UO_324 (O_324,N_19901,N_19836);
and UO_325 (O_325,N_19865,N_19954);
and UO_326 (O_326,N_19912,N_19961);
or UO_327 (O_327,N_19874,N_19940);
and UO_328 (O_328,N_19861,N_19994);
nor UO_329 (O_329,N_19928,N_19896);
and UO_330 (O_330,N_19941,N_19914);
xnor UO_331 (O_331,N_19900,N_19916);
nor UO_332 (O_332,N_19921,N_19872);
xor UO_333 (O_333,N_19955,N_19839);
nor UO_334 (O_334,N_19982,N_19852);
nor UO_335 (O_335,N_19993,N_19956);
nor UO_336 (O_336,N_19870,N_19888);
or UO_337 (O_337,N_19977,N_19830);
nor UO_338 (O_338,N_19975,N_19879);
or UO_339 (O_339,N_19949,N_19845);
and UO_340 (O_340,N_19989,N_19850);
or UO_341 (O_341,N_19977,N_19868);
and UO_342 (O_342,N_19915,N_19989);
and UO_343 (O_343,N_19960,N_19967);
nor UO_344 (O_344,N_19863,N_19862);
or UO_345 (O_345,N_19979,N_19828);
nor UO_346 (O_346,N_19945,N_19831);
nor UO_347 (O_347,N_19962,N_19850);
xor UO_348 (O_348,N_19853,N_19939);
nand UO_349 (O_349,N_19804,N_19934);
nor UO_350 (O_350,N_19916,N_19968);
or UO_351 (O_351,N_19958,N_19903);
xor UO_352 (O_352,N_19824,N_19880);
or UO_353 (O_353,N_19895,N_19817);
or UO_354 (O_354,N_19919,N_19878);
and UO_355 (O_355,N_19835,N_19808);
and UO_356 (O_356,N_19928,N_19902);
or UO_357 (O_357,N_19889,N_19970);
and UO_358 (O_358,N_19918,N_19925);
nand UO_359 (O_359,N_19870,N_19914);
and UO_360 (O_360,N_19880,N_19983);
and UO_361 (O_361,N_19921,N_19959);
nand UO_362 (O_362,N_19830,N_19857);
or UO_363 (O_363,N_19938,N_19970);
nand UO_364 (O_364,N_19961,N_19905);
nor UO_365 (O_365,N_19985,N_19921);
or UO_366 (O_366,N_19952,N_19804);
xnor UO_367 (O_367,N_19973,N_19915);
or UO_368 (O_368,N_19890,N_19821);
nor UO_369 (O_369,N_19847,N_19924);
or UO_370 (O_370,N_19957,N_19991);
nor UO_371 (O_371,N_19817,N_19999);
or UO_372 (O_372,N_19859,N_19894);
nand UO_373 (O_373,N_19855,N_19976);
or UO_374 (O_374,N_19953,N_19943);
and UO_375 (O_375,N_19898,N_19977);
nor UO_376 (O_376,N_19836,N_19965);
and UO_377 (O_377,N_19945,N_19941);
nand UO_378 (O_378,N_19954,N_19875);
or UO_379 (O_379,N_19910,N_19952);
nand UO_380 (O_380,N_19849,N_19838);
nor UO_381 (O_381,N_19828,N_19969);
and UO_382 (O_382,N_19994,N_19991);
nor UO_383 (O_383,N_19814,N_19823);
xnor UO_384 (O_384,N_19876,N_19940);
xor UO_385 (O_385,N_19962,N_19848);
and UO_386 (O_386,N_19808,N_19892);
nor UO_387 (O_387,N_19960,N_19870);
nor UO_388 (O_388,N_19852,N_19934);
nand UO_389 (O_389,N_19935,N_19969);
xnor UO_390 (O_390,N_19810,N_19969);
nor UO_391 (O_391,N_19842,N_19803);
nor UO_392 (O_392,N_19821,N_19974);
nor UO_393 (O_393,N_19903,N_19989);
or UO_394 (O_394,N_19985,N_19967);
xnor UO_395 (O_395,N_19891,N_19975);
nand UO_396 (O_396,N_19863,N_19833);
xnor UO_397 (O_397,N_19971,N_19891);
and UO_398 (O_398,N_19914,N_19894);
or UO_399 (O_399,N_19806,N_19890);
or UO_400 (O_400,N_19807,N_19989);
nor UO_401 (O_401,N_19802,N_19996);
xnor UO_402 (O_402,N_19852,N_19909);
nand UO_403 (O_403,N_19865,N_19804);
xnor UO_404 (O_404,N_19884,N_19952);
nor UO_405 (O_405,N_19868,N_19960);
and UO_406 (O_406,N_19934,N_19947);
xnor UO_407 (O_407,N_19879,N_19899);
xor UO_408 (O_408,N_19981,N_19861);
nand UO_409 (O_409,N_19818,N_19912);
xnor UO_410 (O_410,N_19909,N_19881);
nor UO_411 (O_411,N_19957,N_19947);
or UO_412 (O_412,N_19929,N_19820);
nand UO_413 (O_413,N_19851,N_19858);
and UO_414 (O_414,N_19829,N_19984);
nor UO_415 (O_415,N_19946,N_19835);
xnor UO_416 (O_416,N_19974,N_19896);
and UO_417 (O_417,N_19856,N_19826);
nor UO_418 (O_418,N_19962,N_19844);
nor UO_419 (O_419,N_19820,N_19937);
xor UO_420 (O_420,N_19989,N_19907);
xor UO_421 (O_421,N_19886,N_19872);
or UO_422 (O_422,N_19882,N_19983);
and UO_423 (O_423,N_19832,N_19917);
xor UO_424 (O_424,N_19953,N_19925);
nor UO_425 (O_425,N_19967,N_19989);
xor UO_426 (O_426,N_19992,N_19915);
nor UO_427 (O_427,N_19845,N_19912);
and UO_428 (O_428,N_19849,N_19955);
or UO_429 (O_429,N_19888,N_19805);
or UO_430 (O_430,N_19977,N_19936);
nand UO_431 (O_431,N_19895,N_19826);
and UO_432 (O_432,N_19840,N_19872);
xor UO_433 (O_433,N_19926,N_19958);
nor UO_434 (O_434,N_19966,N_19981);
nor UO_435 (O_435,N_19922,N_19859);
xor UO_436 (O_436,N_19828,N_19883);
nand UO_437 (O_437,N_19966,N_19876);
nor UO_438 (O_438,N_19804,N_19979);
xnor UO_439 (O_439,N_19976,N_19904);
xnor UO_440 (O_440,N_19802,N_19982);
xor UO_441 (O_441,N_19802,N_19872);
nor UO_442 (O_442,N_19992,N_19848);
or UO_443 (O_443,N_19863,N_19933);
nor UO_444 (O_444,N_19871,N_19831);
xnor UO_445 (O_445,N_19808,N_19828);
xor UO_446 (O_446,N_19969,N_19916);
nor UO_447 (O_447,N_19888,N_19934);
nand UO_448 (O_448,N_19901,N_19804);
and UO_449 (O_449,N_19843,N_19940);
nand UO_450 (O_450,N_19889,N_19927);
or UO_451 (O_451,N_19845,N_19828);
and UO_452 (O_452,N_19881,N_19817);
xnor UO_453 (O_453,N_19931,N_19935);
nor UO_454 (O_454,N_19810,N_19908);
and UO_455 (O_455,N_19910,N_19897);
xor UO_456 (O_456,N_19988,N_19852);
xor UO_457 (O_457,N_19985,N_19870);
or UO_458 (O_458,N_19936,N_19955);
and UO_459 (O_459,N_19880,N_19898);
nand UO_460 (O_460,N_19904,N_19860);
nor UO_461 (O_461,N_19894,N_19990);
xnor UO_462 (O_462,N_19843,N_19975);
nor UO_463 (O_463,N_19959,N_19951);
and UO_464 (O_464,N_19914,N_19988);
nor UO_465 (O_465,N_19802,N_19863);
nor UO_466 (O_466,N_19921,N_19918);
and UO_467 (O_467,N_19851,N_19845);
and UO_468 (O_468,N_19934,N_19863);
xnor UO_469 (O_469,N_19889,N_19935);
and UO_470 (O_470,N_19922,N_19957);
xnor UO_471 (O_471,N_19845,N_19925);
xor UO_472 (O_472,N_19980,N_19867);
xnor UO_473 (O_473,N_19913,N_19976);
or UO_474 (O_474,N_19990,N_19868);
and UO_475 (O_475,N_19842,N_19909);
and UO_476 (O_476,N_19838,N_19803);
nand UO_477 (O_477,N_19818,N_19890);
xor UO_478 (O_478,N_19868,N_19814);
or UO_479 (O_479,N_19904,N_19951);
or UO_480 (O_480,N_19891,N_19958);
xor UO_481 (O_481,N_19937,N_19953);
nand UO_482 (O_482,N_19812,N_19849);
or UO_483 (O_483,N_19966,N_19813);
xnor UO_484 (O_484,N_19800,N_19904);
or UO_485 (O_485,N_19869,N_19801);
nand UO_486 (O_486,N_19916,N_19976);
nor UO_487 (O_487,N_19980,N_19888);
or UO_488 (O_488,N_19997,N_19809);
nand UO_489 (O_489,N_19939,N_19800);
xor UO_490 (O_490,N_19969,N_19911);
or UO_491 (O_491,N_19830,N_19874);
and UO_492 (O_492,N_19961,N_19953);
or UO_493 (O_493,N_19987,N_19998);
nor UO_494 (O_494,N_19810,N_19851);
or UO_495 (O_495,N_19927,N_19986);
or UO_496 (O_496,N_19822,N_19844);
or UO_497 (O_497,N_19829,N_19976);
or UO_498 (O_498,N_19855,N_19859);
or UO_499 (O_499,N_19982,N_19834);
or UO_500 (O_500,N_19965,N_19831);
and UO_501 (O_501,N_19907,N_19971);
or UO_502 (O_502,N_19807,N_19965);
or UO_503 (O_503,N_19930,N_19936);
and UO_504 (O_504,N_19921,N_19871);
and UO_505 (O_505,N_19984,N_19843);
or UO_506 (O_506,N_19844,N_19861);
and UO_507 (O_507,N_19813,N_19911);
nor UO_508 (O_508,N_19880,N_19948);
or UO_509 (O_509,N_19878,N_19839);
nor UO_510 (O_510,N_19834,N_19813);
nand UO_511 (O_511,N_19878,N_19891);
nor UO_512 (O_512,N_19829,N_19843);
xor UO_513 (O_513,N_19805,N_19930);
nor UO_514 (O_514,N_19950,N_19886);
or UO_515 (O_515,N_19921,N_19978);
and UO_516 (O_516,N_19933,N_19934);
or UO_517 (O_517,N_19909,N_19958);
or UO_518 (O_518,N_19937,N_19861);
and UO_519 (O_519,N_19833,N_19992);
nand UO_520 (O_520,N_19877,N_19918);
and UO_521 (O_521,N_19993,N_19890);
nand UO_522 (O_522,N_19906,N_19949);
or UO_523 (O_523,N_19890,N_19832);
xor UO_524 (O_524,N_19898,N_19986);
nor UO_525 (O_525,N_19854,N_19930);
xor UO_526 (O_526,N_19934,N_19999);
xnor UO_527 (O_527,N_19873,N_19848);
xnor UO_528 (O_528,N_19977,N_19958);
or UO_529 (O_529,N_19994,N_19876);
nor UO_530 (O_530,N_19815,N_19884);
and UO_531 (O_531,N_19938,N_19928);
and UO_532 (O_532,N_19850,N_19935);
xor UO_533 (O_533,N_19991,N_19920);
nand UO_534 (O_534,N_19886,N_19840);
nand UO_535 (O_535,N_19957,N_19913);
xor UO_536 (O_536,N_19809,N_19855);
or UO_537 (O_537,N_19988,N_19811);
or UO_538 (O_538,N_19883,N_19811);
nor UO_539 (O_539,N_19947,N_19828);
xnor UO_540 (O_540,N_19961,N_19801);
xor UO_541 (O_541,N_19940,N_19873);
nand UO_542 (O_542,N_19932,N_19888);
and UO_543 (O_543,N_19802,N_19887);
nor UO_544 (O_544,N_19988,N_19939);
and UO_545 (O_545,N_19866,N_19909);
or UO_546 (O_546,N_19936,N_19863);
xor UO_547 (O_547,N_19949,N_19862);
and UO_548 (O_548,N_19920,N_19887);
and UO_549 (O_549,N_19860,N_19803);
nor UO_550 (O_550,N_19974,N_19808);
nand UO_551 (O_551,N_19817,N_19824);
xor UO_552 (O_552,N_19824,N_19842);
nand UO_553 (O_553,N_19875,N_19835);
or UO_554 (O_554,N_19934,N_19891);
xor UO_555 (O_555,N_19800,N_19855);
nor UO_556 (O_556,N_19961,N_19844);
or UO_557 (O_557,N_19965,N_19951);
and UO_558 (O_558,N_19924,N_19819);
nor UO_559 (O_559,N_19837,N_19804);
or UO_560 (O_560,N_19982,N_19915);
and UO_561 (O_561,N_19972,N_19838);
nand UO_562 (O_562,N_19929,N_19934);
nand UO_563 (O_563,N_19973,N_19846);
nand UO_564 (O_564,N_19951,N_19812);
and UO_565 (O_565,N_19996,N_19914);
nand UO_566 (O_566,N_19805,N_19959);
or UO_567 (O_567,N_19853,N_19865);
and UO_568 (O_568,N_19843,N_19857);
nand UO_569 (O_569,N_19947,N_19938);
or UO_570 (O_570,N_19873,N_19846);
and UO_571 (O_571,N_19896,N_19854);
and UO_572 (O_572,N_19987,N_19883);
or UO_573 (O_573,N_19951,N_19997);
nor UO_574 (O_574,N_19978,N_19871);
or UO_575 (O_575,N_19829,N_19857);
nand UO_576 (O_576,N_19904,N_19992);
and UO_577 (O_577,N_19881,N_19843);
and UO_578 (O_578,N_19842,N_19809);
nand UO_579 (O_579,N_19855,N_19872);
or UO_580 (O_580,N_19859,N_19924);
and UO_581 (O_581,N_19990,N_19889);
and UO_582 (O_582,N_19953,N_19996);
nand UO_583 (O_583,N_19941,N_19919);
and UO_584 (O_584,N_19811,N_19834);
nor UO_585 (O_585,N_19809,N_19816);
or UO_586 (O_586,N_19936,N_19973);
or UO_587 (O_587,N_19959,N_19891);
and UO_588 (O_588,N_19858,N_19824);
nor UO_589 (O_589,N_19876,N_19863);
xor UO_590 (O_590,N_19995,N_19982);
and UO_591 (O_591,N_19887,N_19912);
nor UO_592 (O_592,N_19896,N_19936);
and UO_593 (O_593,N_19906,N_19942);
xnor UO_594 (O_594,N_19800,N_19962);
xor UO_595 (O_595,N_19966,N_19885);
nand UO_596 (O_596,N_19822,N_19912);
and UO_597 (O_597,N_19880,N_19804);
xor UO_598 (O_598,N_19857,N_19929);
nand UO_599 (O_599,N_19982,N_19858);
or UO_600 (O_600,N_19845,N_19945);
or UO_601 (O_601,N_19871,N_19867);
nand UO_602 (O_602,N_19915,N_19809);
nor UO_603 (O_603,N_19805,N_19954);
and UO_604 (O_604,N_19858,N_19895);
nand UO_605 (O_605,N_19817,N_19967);
xnor UO_606 (O_606,N_19953,N_19831);
nor UO_607 (O_607,N_19815,N_19943);
or UO_608 (O_608,N_19849,N_19817);
nand UO_609 (O_609,N_19893,N_19868);
and UO_610 (O_610,N_19972,N_19953);
and UO_611 (O_611,N_19873,N_19932);
nand UO_612 (O_612,N_19936,N_19921);
and UO_613 (O_613,N_19865,N_19827);
nand UO_614 (O_614,N_19809,N_19965);
or UO_615 (O_615,N_19841,N_19879);
xor UO_616 (O_616,N_19935,N_19992);
xnor UO_617 (O_617,N_19961,N_19979);
or UO_618 (O_618,N_19920,N_19822);
and UO_619 (O_619,N_19920,N_19996);
nand UO_620 (O_620,N_19990,N_19996);
nand UO_621 (O_621,N_19871,N_19932);
and UO_622 (O_622,N_19838,N_19806);
nand UO_623 (O_623,N_19867,N_19925);
xnor UO_624 (O_624,N_19937,N_19900);
and UO_625 (O_625,N_19918,N_19939);
and UO_626 (O_626,N_19958,N_19873);
nand UO_627 (O_627,N_19802,N_19937);
or UO_628 (O_628,N_19874,N_19948);
and UO_629 (O_629,N_19989,N_19808);
and UO_630 (O_630,N_19970,N_19895);
or UO_631 (O_631,N_19959,N_19907);
xnor UO_632 (O_632,N_19946,N_19926);
nand UO_633 (O_633,N_19827,N_19920);
xor UO_634 (O_634,N_19893,N_19902);
and UO_635 (O_635,N_19897,N_19928);
nand UO_636 (O_636,N_19815,N_19840);
nor UO_637 (O_637,N_19979,N_19879);
xor UO_638 (O_638,N_19804,N_19964);
or UO_639 (O_639,N_19831,N_19957);
and UO_640 (O_640,N_19939,N_19862);
or UO_641 (O_641,N_19921,N_19983);
and UO_642 (O_642,N_19916,N_19860);
nand UO_643 (O_643,N_19841,N_19850);
or UO_644 (O_644,N_19838,N_19902);
xnor UO_645 (O_645,N_19800,N_19899);
or UO_646 (O_646,N_19864,N_19890);
and UO_647 (O_647,N_19928,N_19994);
or UO_648 (O_648,N_19893,N_19944);
nand UO_649 (O_649,N_19979,N_19859);
and UO_650 (O_650,N_19998,N_19887);
nand UO_651 (O_651,N_19878,N_19852);
nor UO_652 (O_652,N_19857,N_19920);
xnor UO_653 (O_653,N_19810,N_19871);
xnor UO_654 (O_654,N_19818,N_19847);
nand UO_655 (O_655,N_19980,N_19827);
nand UO_656 (O_656,N_19889,N_19983);
or UO_657 (O_657,N_19816,N_19968);
nor UO_658 (O_658,N_19957,N_19936);
and UO_659 (O_659,N_19838,N_19981);
nand UO_660 (O_660,N_19953,N_19951);
or UO_661 (O_661,N_19913,N_19948);
nand UO_662 (O_662,N_19915,N_19987);
nand UO_663 (O_663,N_19817,N_19856);
and UO_664 (O_664,N_19973,N_19985);
and UO_665 (O_665,N_19966,N_19802);
nor UO_666 (O_666,N_19915,N_19868);
nand UO_667 (O_667,N_19946,N_19897);
xnor UO_668 (O_668,N_19955,N_19820);
or UO_669 (O_669,N_19834,N_19915);
and UO_670 (O_670,N_19872,N_19957);
nand UO_671 (O_671,N_19912,N_19820);
nor UO_672 (O_672,N_19819,N_19835);
nand UO_673 (O_673,N_19823,N_19897);
nand UO_674 (O_674,N_19860,N_19981);
nand UO_675 (O_675,N_19807,N_19846);
and UO_676 (O_676,N_19991,N_19815);
and UO_677 (O_677,N_19929,N_19804);
or UO_678 (O_678,N_19803,N_19844);
or UO_679 (O_679,N_19952,N_19968);
nor UO_680 (O_680,N_19817,N_19885);
xnor UO_681 (O_681,N_19985,N_19911);
nand UO_682 (O_682,N_19814,N_19907);
and UO_683 (O_683,N_19927,N_19817);
nor UO_684 (O_684,N_19916,N_19957);
and UO_685 (O_685,N_19851,N_19900);
nor UO_686 (O_686,N_19959,N_19847);
xnor UO_687 (O_687,N_19986,N_19800);
and UO_688 (O_688,N_19856,N_19945);
and UO_689 (O_689,N_19967,N_19857);
xor UO_690 (O_690,N_19875,N_19903);
nor UO_691 (O_691,N_19977,N_19970);
nor UO_692 (O_692,N_19809,N_19928);
xor UO_693 (O_693,N_19873,N_19899);
nor UO_694 (O_694,N_19986,N_19946);
nor UO_695 (O_695,N_19914,N_19800);
and UO_696 (O_696,N_19842,N_19904);
xor UO_697 (O_697,N_19990,N_19908);
nor UO_698 (O_698,N_19912,N_19941);
and UO_699 (O_699,N_19874,N_19943);
nand UO_700 (O_700,N_19845,N_19895);
or UO_701 (O_701,N_19927,N_19981);
or UO_702 (O_702,N_19860,N_19857);
nor UO_703 (O_703,N_19813,N_19868);
nor UO_704 (O_704,N_19850,N_19875);
nand UO_705 (O_705,N_19961,N_19813);
and UO_706 (O_706,N_19936,N_19953);
or UO_707 (O_707,N_19995,N_19970);
and UO_708 (O_708,N_19802,N_19986);
or UO_709 (O_709,N_19877,N_19946);
nand UO_710 (O_710,N_19976,N_19885);
and UO_711 (O_711,N_19863,N_19935);
and UO_712 (O_712,N_19800,N_19888);
nor UO_713 (O_713,N_19805,N_19925);
or UO_714 (O_714,N_19859,N_19851);
xnor UO_715 (O_715,N_19899,N_19906);
xor UO_716 (O_716,N_19822,N_19848);
nand UO_717 (O_717,N_19917,N_19888);
nor UO_718 (O_718,N_19845,N_19820);
nor UO_719 (O_719,N_19903,N_19970);
xnor UO_720 (O_720,N_19916,N_19862);
xnor UO_721 (O_721,N_19800,N_19875);
nand UO_722 (O_722,N_19988,N_19889);
and UO_723 (O_723,N_19931,N_19823);
or UO_724 (O_724,N_19807,N_19905);
and UO_725 (O_725,N_19932,N_19846);
xnor UO_726 (O_726,N_19839,N_19905);
xnor UO_727 (O_727,N_19802,N_19867);
nor UO_728 (O_728,N_19827,N_19941);
nor UO_729 (O_729,N_19811,N_19807);
nor UO_730 (O_730,N_19857,N_19988);
nand UO_731 (O_731,N_19825,N_19944);
and UO_732 (O_732,N_19817,N_19980);
xor UO_733 (O_733,N_19889,N_19993);
nor UO_734 (O_734,N_19815,N_19960);
nor UO_735 (O_735,N_19898,N_19846);
xnor UO_736 (O_736,N_19906,N_19894);
nor UO_737 (O_737,N_19932,N_19852);
nor UO_738 (O_738,N_19916,N_19889);
nand UO_739 (O_739,N_19861,N_19944);
xnor UO_740 (O_740,N_19962,N_19816);
xnor UO_741 (O_741,N_19856,N_19878);
xnor UO_742 (O_742,N_19961,N_19972);
or UO_743 (O_743,N_19919,N_19999);
nor UO_744 (O_744,N_19827,N_19967);
nand UO_745 (O_745,N_19808,N_19921);
xor UO_746 (O_746,N_19868,N_19979);
nor UO_747 (O_747,N_19924,N_19857);
xor UO_748 (O_748,N_19884,N_19857);
nand UO_749 (O_749,N_19927,N_19961);
nand UO_750 (O_750,N_19897,N_19896);
xor UO_751 (O_751,N_19953,N_19939);
xor UO_752 (O_752,N_19818,N_19983);
and UO_753 (O_753,N_19874,N_19901);
or UO_754 (O_754,N_19840,N_19989);
nand UO_755 (O_755,N_19876,N_19869);
and UO_756 (O_756,N_19862,N_19885);
nand UO_757 (O_757,N_19895,N_19949);
nand UO_758 (O_758,N_19877,N_19868);
and UO_759 (O_759,N_19919,N_19890);
nand UO_760 (O_760,N_19918,N_19932);
nor UO_761 (O_761,N_19952,N_19890);
or UO_762 (O_762,N_19886,N_19930);
nor UO_763 (O_763,N_19801,N_19937);
and UO_764 (O_764,N_19893,N_19838);
and UO_765 (O_765,N_19984,N_19867);
or UO_766 (O_766,N_19995,N_19988);
xor UO_767 (O_767,N_19947,N_19882);
or UO_768 (O_768,N_19821,N_19902);
nor UO_769 (O_769,N_19824,N_19984);
xor UO_770 (O_770,N_19833,N_19957);
or UO_771 (O_771,N_19826,N_19971);
or UO_772 (O_772,N_19865,N_19974);
nor UO_773 (O_773,N_19936,N_19923);
xnor UO_774 (O_774,N_19945,N_19927);
nand UO_775 (O_775,N_19863,N_19906);
nor UO_776 (O_776,N_19949,N_19903);
nand UO_777 (O_777,N_19949,N_19893);
xor UO_778 (O_778,N_19859,N_19896);
nand UO_779 (O_779,N_19981,N_19867);
xnor UO_780 (O_780,N_19832,N_19868);
or UO_781 (O_781,N_19882,N_19996);
nand UO_782 (O_782,N_19872,N_19832);
and UO_783 (O_783,N_19826,N_19835);
and UO_784 (O_784,N_19808,N_19983);
nor UO_785 (O_785,N_19862,N_19905);
nor UO_786 (O_786,N_19909,N_19829);
nand UO_787 (O_787,N_19800,N_19849);
nor UO_788 (O_788,N_19998,N_19905);
nand UO_789 (O_789,N_19828,N_19953);
and UO_790 (O_790,N_19847,N_19922);
and UO_791 (O_791,N_19993,N_19947);
or UO_792 (O_792,N_19849,N_19854);
nor UO_793 (O_793,N_19978,N_19857);
and UO_794 (O_794,N_19944,N_19981);
or UO_795 (O_795,N_19880,N_19916);
nand UO_796 (O_796,N_19876,N_19841);
nand UO_797 (O_797,N_19827,N_19932);
xor UO_798 (O_798,N_19930,N_19812);
xnor UO_799 (O_799,N_19954,N_19986);
nand UO_800 (O_800,N_19928,N_19856);
xnor UO_801 (O_801,N_19995,N_19973);
nor UO_802 (O_802,N_19888,N_19884);
nand UO_803 (O_803,N_19896,N_19914);
and UO_804 (O_804,N_19991,N_19915);
nor UO_805 (O_805,N_19874,N_19989);
nor UO_806 (O_806,N_19853,N_19944);
or UO_807 (O_807,N_19993,N_19959);
xor UO_808 (O_808,N_19808,N_19836);
nor UO_809 (O_809,N_19929,N_19863);
or UO_810 (O_810,N_19942,N_19889);
nand UO_811 (O_811,N_19970,N_19953);
or UO_812 (O_812,N_19942,N_19893);
and UO_813 (O_813,N_19991,N_19983);
xnor UO_814 (O_814,N_19945,N_19889);
or UO_815 (O_815,N_19816,N_19889);
nor UO_816 (O_816,N_19889,N_19936);
nand UO_817 (O_817,N_19903,N_19900);
nor UO_818 (O_818,N_19984,N_19813);
and UO_819 (O_819,N_19872,N_19926);
nor UO_820 (O_820,N_19933,N_19980);
or UO_821 (O_821,N_19991,N_19832);
xor UO_822 (O_822,N_19897,N_19906);
nand UO_823 (O_823,N_19867,N_19846);
nor UO_824 (O_824,N_19925,N_19929);
or UO_825 (O_825,N_19956,N_19837);
or UO_826 (O_826,N_19866,N_19837);
nor UO_827 (O_827,N_19858,N_19976);
nand UO_828 (O_828,N_19920,N_19839);
nand UO_829 (O_829,N_19812,N_19962);
and UO_830 (O_830,N_19808,N_19926);
nand UO_831 (O_831,N_19881,N_19852);
or UO_832 (O_832,N_19954,N_19836);
or UO_833 (O_833,N_19998,N_19880);
xor UO_834 (O_834,N_19804,N_19826);
and UO_835 (O_835,N_19803,N_19996);
or UO_836 (O_836,N_19823,N_19826);
nand UO_837 (O_837,N_19856,N_19988);
xor UO_838 (O_838,N_19823,N_19821);
nor UO_839 (O_839,N_19876,N_19937);
or UO_840 (O_840,N_19801,N_19988);
and UO_841 (O_841,N_19853,N_19809);
nor UO_842 (O_842,N_19813,N_19963);
or UO_843 (O_843,N_19930,N_19975);
nor UO_844 (O_844,N_19956,N_19891);
xor UO_845 (O_845,N_19844,N_19965);
nor UO_846 (O_846,N_19840,N_19828);
and UO_847 (O_847,N_19817,N_19971);
and UO_848 (O_848,N_19898,N_19802);
nor UO_849 (O_849,N_19916,N_19911);
nand UO_850 (O_850,N_19860,N_19832);
and UO_851 (O_851,N_19943,N_19924);
or UO_852 (O_852,N_19955,N_19995);
nor UO_853 (O_853,N_19929,N_19948);
nand UO_854 (O_854,N_19870,N_19977);
xnor UO_855 (O_855,N_19949,N_19873);
or UO_856 (O_856,N_19947,N_19881);
or UO_857 (O_857,N_19817,N_19816);
nor UO_858 (O_858,N_19919,N_19961);
and UO_859 (O_859,N_19952,N_19875);
nand UO_860 (O_860,N_19938,N_19918);
and UO_861 (O_861,N_19837,N_19963);
xor UO_862 (O_862,N_19990,N_19800);
nand UO_863 (O_863,N_19894,N_19950);
xor UO_864 (O_864,N_19811,N_19962);
or UO_865 (O_865,N_19998,N_19802);
and UO_866 (O_866,N_19966,N_19892);
nor UO_867 (O_867,N_19881,N_19831);
nand UO_868 (O_868,N_19894,N_19981);
nor UO_869 (O_869,N_19866,N_19838);
and UO_870 (O_870,N_19953,N_19817);
nor UO_871 (O_871,N_19850,N_19807);
nand UO_872 (O_872,N_19837,N_19835);
or UO_873 (O_873,N_19842,N_19810);
nand UO_874 (O_874,N_19954,N_19911);
nor UO_875 (O_875,N_19918,N_19887);
nand UO_876 (O_876,N_19857,N_19899);
and UO_877 (O_877,N_19932,N_19968);
nor UO_878 (O_878,N_19872,N_19873);
nor UO_879 (O_879,N_19924,N_19986);
nor UO_880 (O_880,N_19874,N_19996);
xor UO_881 (O_881,N_19940,N_19885);
nand UO_882 (O_882,N_19820,N_19971);
xor UO_883 (O_883,N_19805,N_19934);
or UO_884 (O_884,N_19901,N_19985);
xor UO_885 (O_885,N_19883,N_19801);
xnor UO_886 (O_886,N_19865,N_19977);
xnor UO_887 (O_887,N_19979,N_19924);
nand UO_888 (O_888,N_19857,N_19864);
or UO_889 (O_889,N_19918,N_19982);
nand UO_890 (O_890,N_19838,N_19983);
xor UO_891 (O_891,N_19997,N_19915);
and UO_892 (O_892,N_19960,N_19830);
nand UO_893 (O_893,N_19873,N_19983);
nand UO_894 (O_894,N_19908,N_19864);
xnor UO_895 (O_895,N_19841,N_19917);
nand UO_896 (O_896,N_19861,N_19978);
or UO_897 (O_897,N_19875,N_19984);
and UO_898 (O_898,N_19993,N_19835);
and UO_899 (O_899,N_19984,N_19947);
and UO_900 (O_900,N_19978,N_19836);
nor UO_901 (O_901,N_19904,N_19845);
or UO_902 (O_902,N_19859,N_19828);
nor UO_903 (O_903,N_19879,N_19837);
nand UO_904 (O_904,N_19824,N_19860);
and UO_905 (O_905,N_19941,N_19826);
nand UO_906 (O_906,N_19985,N_19958);
or UO_907 (O_907,N_19915,N_19938);
and UO_908 (O_908,N_19841,N_19989);
or UO_909 (O_909,N_19802,N_19995);
xnor UO_910 (O_910,N_19855,N_19960);
nor UO_911 (O_911,N_19867,N_19848);
nor UO_912 (O_912,N_19965,N_19878);
or UO_913 (O_913,N_19978,N_19864);
and UO_914 (O_914,N_19975,N_19921);
nor UO_915 (O_915,N_19892,N_19944);
and UO_916 (O_916,N_19986,N_19903);
nand UO_917 (O_917,N_19951,N_19822);
nor UO_918 (O_918,N_19892,N_19941);
nor UO_919 (O_919,N_19915,N_19843);
xor UO_920 (O_920,N_19970,N_19971);
xnor UO_921 (O_921,N_19808,N_19993);
nor UO_922 (O_922,N_19842,N_19975);
and UO_923 (O_923,N_19872,N_19876);
nor UO_924 (O_924,N_19920,N_19952);
nand UO_925 (O_925,N_19821,N_19953);
nand UO_926 (O_926,N_19824,N_19848);
and UO_927 (O_927,N_19826,N_19806);
nand UO_928 (O_928,N_19918,N_19884);
or UO_929 (O_929,N_19839,N_19825);
or UO_930 (O_930,N_19997,N_19811);
and UO_931 (O_931,N_19958,N_19801);
nand UO_932 (O_932,N_19849,N_19893);
or UO_933 (O_933,N_19989,N_19938);
xor UO_934 (O_934,N_19911,N_19804);
nor UO_935 (O_935,N_19867,N_19955);
nand UO_936 (O_936,N_19878,N_19962);
or UO_937 (O_937,N_19872,N_19841);
xor UO_938 (O_938,N_19836,N_19815);
xor UO_939 (O_939,N_19821,N_19910);
nor UO_940 (O_940,N_19951,N_19849);
nor UO_941 (O_941,N_19965,N_19980);
or UO_942 (O_942,N_19917,N_19861);
or UO_943 (O_943,N_19907,N_19824);
xor UO_944 (O_944,N_19881,N_19860);
or UO_945 (O_945,N_19867,N_19850);
nand UO_946 (O_946,N_19900,N_19850);
and UO_947 (O_947,N_19844,N_19969);
nor UO_948 (O_948,N_19859,N_19860);
xor UO_949 (O_949,N_19909,N_19801);
nor UO_950 (O_950,N_19876,N_19849);
or UO_951 (O_951,N_19957,N_19996);
or UO_952 (O_952,N_19892,N_19872);
xor UO_953 (O_953,N_19952,N_19913);
nand UO_954 (O_954,N_19830,N_19988);
xnor UO_955 (O_955,N_19892,N_19809);
nand UO_956 (O_956,N_19911,N_19997);
nor UO_957 (O_957,N_19942,N_19892);
and UO_958 (O_958,N_19859,N_19868);
or UO_959 (O_959,N_19816,N_19843);
nor UO_960 (O_960,N_19847,N_19802);
and UO_961 (O_961,N_19942,N_19867);
xor UO_962 (O_962,N_19917,N_19987);
nor UO_963 (O_963,N_19938,N_19829);
and UO_964 (O_964,N_19941,N_19802);
or UO_965 (O_965,N_19991,N_19812);
or UO_966 (O_966,N_19869,N_19973);
or UO_967 (O_967,N_19824,N_19826);
nor UO_968 (O_968,N_19883,N_19911);
nor UO_969 (O_969,N_19980,N_19998);
nor UO_970 (O_970,N_19935,N_19813);
and UO_971 (O_971,N_19884,N_19808);
nand UO_972 (O_972,N_19881,N_19826);
or UO_973 (O_973,N_19850,N_19844);
xor UO_974 (O_974,N_19866,N_19883);
and UO_975 (O_975,N_19895,N_19996);
or UO_976 (O_976,N_19960,N_19833);
xor UO_977 (O_977,N_19801,N_19802);
nor UO_978 (O_978,N_19800,N_19822);
xor UO_979 (O_979,N_19855,N_19908);
or UO_980 (O_980,N_19900,N_19855);
or UO_981 (O_981,N_19910,N_19819);
or UO_982 (O_982,N_19895,N_19926);
nor UO_983 (O_983,N_19855,N_19823);
nand UO_984 (O_984,N_19987,N_19898);
nand UO_985 (O_985,N_19894,N_19908);
xor UO_986 (O_986,N_19949,N_19902);
nor UO_987 (O_987,N_19927,N_19993);
nand UO_988 (O_988,N_19828,N_19975);
or UO_989 (O_989,N_19907,N_19927);
or UO_990 (O_990,N_19840,N_19972);
or UO_991 (O_991,N_19900,N_19830);
nor UO_992 (O_992,N_19832,N_19912);
or UO_993 (O_993,N_19802,N_19906);
and UO_994 (O_994,N_19980,N_19826);
or UO_995 (O_995,N_19948,N_19860);
nand UO_996 (O_996,N_19988,N_19878);
xnor UO_997 (O_997,N_19987,N_19916);
nor UO_998 (O_998,N_19970,N_19881);
nand UO_999 (O_999,N_19948,N_19873);
and UO_1000 (O_1000,N_19979,N_19845);
and UO_1001 (O_1001,N_19833,N_19868);
or UO_1002 (O_1002,N_19960,N_19819);
nor UO_1003 (O_1003,N_19842,N_19991);
or UO_1004 (O_1004,N_19875,N_19889);
nor UO_1005 (O_1005,N_19856,N_19969);
and UO_1006 (O_1006,N_19933,N_19801);
nor UO_1007 (O_1007,N_19970,N_19824);
xnor UO_1008 (O_1008,N_19958,N_19839);
xor UO_1009 (O_1009,N_19980,N_19851);
or UO_1010 (O_1010,N_19882,N_19908);
nand UO_1011 (O_1011,N_19981,N_19880);
nand UO_1012 (O_1012,N_19996,N_19926);
or UO_1013 (O_1013,N_19861,N_19965);
and UO_1014 (O_1014,N_19954,N_19987);
and UO_1015 (O_1015,N_19901,N_19837);
nand UO_1016 (O_1016,N_19985,N_19806);
xor UO_1017 (O_1017,N_19946,N_19951);
xor UO_1018 (O_1018,N_19842,N_19929);
nand UO_1019 (O_1019,N_19879,N_19824);
and UO_1020 (O_1020,N_19934,N_19969);
xnor UO_1021 (O_1021,N_19893,N_19966);
nand UO_1022 (O_1022,N_19980,N_19836);
xnor UO_1023 (O_1023,N_19930,N_19881);
xnor UO_1024 (O_1024,N_19923,N_19909);
and UO_1025 (O_1025,N_19887,N_19987);
nor UO_1026 (O_1026,N_19942,N_19827);
nand UO_1027 (O_1027,N_19874,N_19889);
nor UO_1028 (O_1028,N_19830,N_19980);
and UO_1029 (O_1029,N_19916,N_19807);
and UO_1030 (O_1030,N_19861,N_19990);
nor UO_1031 (O_1031,N_19924,N_19917);
and UO_1032 (O_1032,N_19970,N_19874);
nor UO_1033 (O_1033,N_19941,N_19937);
nor UO_1034 (O_1034,N_19967,N_19982);
nor UO_1035 (O_1035,N_19824,N_19800);
nand UO_1036 (O_1036,N_19896,N_19972);
xor UO_1037 (O_1037,N_19989,N_19969);
nand UO_1038 (O_1038,N_19862,N_19997);
nor UO_1039 (O_1039,N_19915,N_19965);
nor UO_1040 (O_1040,N_19918,N_19910);
nand UO_1041 (O_1041,N_19966,N_19805);
nor UO_1042 (O_1042,N_19806,N_19977);
xor UO_1043 (O_1043,N_19894,N_19857);
or UO_1044 (O_1044,N_19820,N_19808);
nand UO_1045 (O_1045,N_19913,N_19839);
nor UO_1046 (O_1046,N_19964,N_19990);
nand UO_1047 (O_1047,N_19985,N_19915);
nand UO_1048 (O_1048,N_19894,N_19909);
and UO_1049 (O_1049,N_19975,N_19816);
xnor UO_1050 (O_1050,N_19962,N_19959);
xor UO_1051 (O_1051,N_19856,N_19875);
or UO_1052 (O_1052,N_19819,N_19988);
nor UO_1053 (O_1053,N_19813,N_19948);
or UO_1054 (O_1054,N_19927,N_19955);
or UO_1055 (O_1055,N_19800,N_19853);
nor UO_1056 (O_1056,N_19909,N_19844);
or UO_1057 (O_1057,N_19855,N_19885);
nor UO_1058 (O_1058,N_19963,N_19962);
xnor UO_1059 (O_1059,N_19938,N_19981);
nand UO_1060 (O_1060,N_19895,N_19821);
xor UO_1061 (O_1061,N_19879,N_19909);
nor UO_1062 (O_1062,N_19945,N_19866);
or UO_1063 (O_1063,N_19882,N_19925);
xor UO_1064 (O_1064,N_19849,N_19874);
nor UO_1065 (O_1065,N_19940,N_19907);
nor UO_1066 (O_1066,N_19938,N_19913);
or UO_1067 (O_1067,N_19851,N_19993);
nand UO_1068 (O_1068,N_19861,N_19957);
xnor UO_1069 (O_1069,N_19890,N_19947);
or UO_1070 (O_1070,N_19985,N_19807);
xnor UO_1071 (O_1071,N_19921,N_19817);
xnor UO_1072 (O_1072,N_19882,N_19857);
and UO_1073 (O_1073,N_19864,N_19807);
nand UO_1074 (O_1074,N_19880,N_19864);
nor UO_1075 (O_1075,N_19992,N_19865);
and UO_1076 (O_1076,N_19972,N_19836);
or UO_1077 (O_1077,N_19927,N_19862);
nand UO_1078 (O_1078,N_19999,N_19966);
or UO_1079 (O_1079,N_19911,N_19905);
and UO_1080 (O_1080,N_19913,N_19845);
or UO_1081 (O_1081,N_19957,N_19909);
or UO_1082 (O_1082,N_19808,N_19906);
xor UO_1083 (O_1083,N_19899,N_19900);
xnor UO_1084 (O_1084,N_19951,N_19810);
and UO_1085 (O_1085,N_19981,N_19973);
nor UO_1086 (O_1086,N_19857,N_19879);
and UO_1087 (O_1087,N_19858,N_19969);
nor UO_1088 (O_1088,N_19894,N_19998);
or UO_1089 (O_1089,N_19836,N_19873);
and UO_1090 (O_1090,N_19968,N_19899);
or UO_1091 (O_1091,N_19820,N_19828);
nand UO_1092 (O_1092,N_19800,N_19992);
and UO_1093 (O_1093,N_19936,N_19944);
nor UO_1094 (O_1094,N_19997,N_19921);
nand UO_1095 (O_1095,N_19994,N_19984);
nand UO_1096 (O_1096,N_19923,N_19965);
nor UO_1097 (O_1097,N_19940,N_19881);
or UO_1098 (O_1098,N_19921,N_19803);
nand UO_1099 (O_1099,N_19869,N_19823);
and UO_1100 (O_1100,N_19875,N_19986);
xnor UO_1101 (O_1101,N_19926,N_19842);
or UO_1102 (O_1102,N_19950,N_19866);
nor UO_1103 (O_1103,N_19843,N_19885);
nand UO_1104 (O_1104,N_19841,N_19921);
or UO_1105 (O_1105,N_19815,N_19850);
or UO_1106 (O_1106,N_19870,N_19811);
nand UO_1107 (O_1107,N_19844,N_19805);
xor UO_1108 (O_1108,N_19945,N_19959);
and UO_1109 (O_1109,N_19835,N_19863);
nand UO_1110 (O_1110,N_19924,N_19901);
nor UO_1111 (O_1111,N_19940,N_19963);
nand UO_1112 (O_1112,N_19893,N_19895);
xnor UO_1113 (O_1113,N_19953,N_19998);
and UO_1114 (O_1114,N_19800,N_19928);
nor UO_1115 (O_1115,N_19828,N_19987);
nor UO_1116 (O_1116,N_19889,N_19896);
or UO_1117 (O_1117,N_19996,N_19861);
nor UO_1118 (O_1118,N_19807,N_19839);
or UO_1119 (O_1119,N_19921,N_19966);
xor UO_1120 (O_1120,N_19989,N_19936);
nand UO_1121 (O_1121,N_19948,N_19832);
xnor UO_1122 (O_1122,N_19801,N_19920);
and UO_1123 (O_1123,N_19995,N_19999);
or UO_1124 (O_1124,N_19828,N_19830);
or UO_1125 (O_1125,N_19892,N_19839);
or UO_1126 (O_1126,N_19975,N_19867);
xnor UO_1127 (O_1127,N_19962,N_19926);
nand UO_1128 (O_1128,N_19957,N_19945);
nor UO_1129 (O_1129,N_19958,N_19971);
or UO_1130 (O_1130,N_19949,N_19877);
xor UO_1131 (O_1131,N_19887,N_19845);
and UO_1132 (O_1132,N_19943,N_19970);
nor UO_1133 (O_1133,N_19819,N_19978);
xor UO_1134 (O_1134,N_19949,N_19840);
nand UO_1135 (O_1135,N_19918,N_19948);
and UO_1136 (O_1136,N_19907,N_19833);
nor UO_1137 (O_1137,N_19907,N_19957);
nor UO_1138 (O_1138,N_19836,N_19927);
xnor UO_1139 (O_1139,N_19910,N_19946);
nand UO_1140 (O_1140,N_19905,N_19861);
and UO_1141 (O_1141,N_19878,N_19951);
nand UO_1142 (O_1142,N_19864,N_19850);
nand UO_1143 (O_1143,N_19961,N_19938);
and UO_1144 (O_1144,N_19897,N_19987);
and UO_1145 (O_1145,N_19825,N_19948);
or UO_1146 (O_1146,N_19813,N_19827);
nor UO_1147 (O_1147,N_19879,N_19910);
nand UO_1148 (O_1148,N_19828,N_19871);
nor UO_1149 (O_1149,N_19912,N_19824);
nor UO_1150 (O_1150,N_19898,N_19912);
and UO_1151 (O_1151,N_19887,N_19929);
xor UO_1152 (O_1152,N_19892,N_19902);
and UO_1153 (O_1153,N_19835,N_19877);
or UO_1154 (O_1154,N_19801,N_19900);
or UO_1155 (O_1155,N_19991,N_19850);
nor UO_1156 (O_1156,N_19870,N_19832);
nand UO_1157 (O_1157,N_19883,N_19837);
and UO_1158 (O_1158,N_19973,N_19942);
and UO_1159 (O_1159,N_19849,N_19832);
xnor UO_1160 (O_1160,N_19898,N_19980);
nand UO_1161 (O_1161,N_19827,N_19860);
or UO_1162 (O_1162,N_19867,N_19890);
or UO_1163 (O_1163,N_19848,N_19919);
or UO_1164 (O_1164,N_19867,N_19986);
nor UO_1165 (O_1165,N_19851,N_19977);
nand UO_1166 (O_1166,N_19989,N_19892);
nor UO_1167 (O_1167,N_19832,N_19846);
nor UO_1168 (O_1168,N_19900,N_19949);
nand UO_1169 (O_1169,N_19899,N_19883);
xnor UO_1170 (O_1170,N_19819,N_19931);
nand UO_1171 (O_1171,N_19985,N_19878);
nor UO_1172 (O_1172,N_19907,N_19832);
or UO_1173 (O_1173,N_19812,N_19967);
and UO_1174 (O_1174,N_19970,N_19827);
nand UO_1175 (O_1175,N_19930,N_19987);
and UO_1176 (O_1176,N_19807,N_19972);
or UO_1177 (O_1177,N_19854,N_19940);
or UO_1178 (O_1178,N_19997,N_19840);
nor UO_1179 (O_1179,N_19906,N_19810);
nand UO_1180 (O_1180,N_19966,N_19930);
nor UO_1181 (O_1181,N_19948,N_19849);
xor UO_1182 (O_1182,N_19880,N_19906);
or UO_1183 (O_1183,N_19937,N_19980);
and UO_1184 (O_1184,N_19993,N_19885);
nand UO_1185 (O_1185,N_19938,N_19982);
nand UO_1186 (O_1186,N_19943,N_19865);
and UO_1187 (O_1187,N_19996,N_19821);
xnor UO_1188 (O_1188,N_19961,N_19976);
and UO_1189 (O_1189,N_19836,N_19941);
nor UO_1190 (O_1190,N_19807,N_19995);
or UO_1191 (O_1191,N_19907,N_19924);
xnor UO_1192 (O_1192,N_19832,N_19853);
xnor UO_1193 (O_1193,N_19851,N_19967);
nand UO_1194 (O_1194,N_19837,N_19842);
nand UO_1195 (O_1195,N_19881,N_19823);
nand UO_1196 (O_1196,N_19944,N_19840);
xor UO_1197 (O_1197,N_19970,N_19954);
nand UO_1198 (O_1198,N_19981,N_19891);
or UO_1199 (O_1199,N_19890,N_19881);
nand UO_1200 (O_1200,N_19935,N_19927);
or UO_1201 (O_1201,N_19901,N_19859);
and UO_1202 (O_1202,N_19802,N_19921);
nor UO_1203 (O_1203,N_19890,N_19964);
or UO_1204 (O_1204,N_19988,N_19919);
nor UO_1205 (O_1205,N_19992,N_19978);
and UO_1206 (O_1206,N_19979,N_19898);
or UO_1207 (O_1207,N_19983,N_19950);
and UO_1208 (O_1208,N_19870,N_19929);
and UO_1209 (O_1209,N_19839,N_19951);
nor UO_1210 (O_1210,N_19814,N_19993);
xnor UO_1211 (O_1211,N_19952,N_19863);
nand UO_1212 (O_1212,N_19951,N_19974);
nor UO_1213 (O_1213,N_19987,N_19895);
or UO_1214 (O_1214,N_19915,N_19984);
and UO_1215 (O_1215,N_19892,N_19830);
or UO_1216 (O_1216,N_19880,N_19900);
xnor UO_1217 (O_1217,N_19990,N_19923);
or UO_1218 (O_1218,N_19878,N_19877);
or UO_1219 (O_1219,N_19959,N_19841);
nand UO_1220 (O_1220,N_19849,N_19915);
and UO_1221 (O_1221,N_19883,N_19867);
nor UO_1222 (O_1222,N_19957,N_19980);
nand UO_1223 (O_1223,N_19935,N_19842);
nor UO_1224 (O_1224,N_19941,N_19841);
nand UO_1225 (O_1225,N_19997,N_19917);
nand UO_1226 (O_1226,N_19978,N_19980);
nor UO_1227 (O_1227,N_19836,N_19912);
nor UO_1228 (O_1228,N_19972,N_19855);
nor UO_1229 (O_1229,N_19859,N_19842);
nand UO_1230 (O_1230,N_19905,N_19999);
nand UO_1231 (O_1231,N_19940,N_19814);
nor UO_1232 (O_1232,N_19827,N_19917);
nor UO_1233 (O_1233,N_19938,N_19922);
nor UO_1234 (O_1234,N_19835,N_19860);
nor UO_1235 (O_1235,N_19978,N_19940);
or UO_1236 (O_1236,N_19904,N_19997);
xnor UO_1237 (O_1237,N_19815,N_19879);
or UO_1238 (O_1238,N_19800,N_19917);
nand UO_1239 (O_1239,N_19949,N_19802);
or UO_1240 (O_1240,N_19851,N_19833);
nor UO_1241 (O_1241,N_19873,N_19802);
nor UO_1242 (O_1242,N_19826,N_19841);
nand UO_1243 (O_1243,N_19907,N_19967);
nand UO_1244 (O_1244,N_19957,N_19827);
or UO_1245 (O_1245,N_19961,N_19888);
nand UO_1246 (O_1246,N_19824,N_19897);
nor UO_1247 (O_1247,N_19808,N_19859);
nand UO_1248 (O_1248,N_19846,N_19965);
nand UO_1249 (O_1249,N_19923,N_19837);
nand UO_1250 (O_1250,N_19828,N_19849);
or UO_1251 (O_1251,N_19908,N_19913);
nand UO_1252 (O_1252,N_19965,N_19979);
xnor UO_1253 (O_1253,N_19971,N_19840);
and UO_1254 (O_1254,N_19852,N_19955);
or UO_1255 (O_1255,N_19911,N_19959);
nor UO_1256 (O_1256,N_19989,N_19988);
nand UO_1257 (O_1257,N_19833,N_19925);
and UO_1258 (O_1258,N_19821,N_19881);
nand UO_1259 (O_1259,N_19810,N_19838);
nor UO_1260 (O_1260,N_19931,N_19859);
nand UO_1261 (O_1261,N_19838,N_19835);
xor UO_1262 (O_1262,N_19804,N_19997);
and UO_1263 (O_1263,N_19911,N_19906);
or UO_1264 (O_1264,N_19975,N_19815);
nor UO_1265 (O_1265,N_19949,N_19919);
xor UO_1266 (O_1266,N_19935,N_19991);
nor UO_1267 (O_1267,N_19980,N_19845);
nor UO_1268 (O_1268,N_19834,N_19877);
or UO_1269 (O_1269,N_19815,N_19858);
or UO_1270 (O_1270,N_19810,N_19934);
nor UO_1271 (O_1271,N_19825,N_19883);
nor UO_1272 (O_1272,N_19859,N_19970);
and UO_1273 (O_1273,N_19910,N_19990);
xnor UO_1274 (O_1274,N_19916,N_19980);
nor UO_1275 (O_1275,N_19975,N_19979);
nand UO_1276 (O_1276,N_19848,N_19862);
or UO_1277 (O_1277,N_19926,N_19959);
or UO_1278 (O_1278,N_19994,N_19822);
or UO_1279 (O_1279,N_19877,N_19974);
or UO_1280 (O_1280,N_19887,N_19953);
nand UO_1281 (O_1281,N_19975,N_19833);
xor UO_1282 (O_1282,N_19871,N_19826);
nand UO_1283 (O_1283,N_19854,N_19953);
nand UO_1284 (O_1284,N_19815,N_19898);
or UO_1285 (O_1285,N_19934,N_19958);
nand UO_1286 (O_1286,N_19946,N_19915);
nor UO_1287 (O_1287,N_19907,N_19870);
nor UO_1288 (O_1288,N_19830,N_19832);
and UO_1289 (O_1289,N_19831,N_19979);
xnor UO_1290 (O_1290,N_19955,N_19912);
xor UO_1291 (O_1291,N_19832,N_19982);
or UO_1292 (O_1292,N_19974,N_19806);
and UO_1293 (O_1293,N_19899,N_19850);
and UO_1294 (O_1294,N_19976,N_19967);
and UO_1295 (O_1295,N_19947,N_19969);
and UO_1296 (O_1296,N_19841,N_19939);
or UO_1297 (O_1297,N_19975,N_19980);
nor UO_1298 (O_1298,N_19865,N_19998);
nand UO_1299 (O_1299,N_19990,N_19860);
nor UO_1300 (O_1300,N_19996,N_19973);
and UO_1301 (O_1301,N_19830,N_19885);
nand UO_1302 (O_1302,N_19981,N_19872);
xor UO_1303 (O_1303,N_19845,N_19834);
nand UO_1304 (O_1304,N_19844,N_19977);
or UO_1305 (O_1305,N_19836,N_19961);
xor UO_1306 (O_1306,N_19844,N_19997);
and UO_1307 (O_1307,N_19970,N_19872);
nand UO_1308 (O_1308,N_19963,N_19953);
and UO_1309 (O_1309,N_19923,N_19893);
and UO_1310 (O_1310,N_19898,N_19857);
and UO_1311 (O_1311,N_19850,N_19849);
and UO_1312 (O_1312,N_19882,N_19910);
nand UO_1313 (O_1313,N_19993,N_19816);
and UO_1314 (O_1314,N_19840,N_19832);
or UO_1315 (O_1315,N_19803,N_19885);
nor UO_1316 (O_1316,N_19809,N_19889);
nand UO_1317 (O_1317,N_19892,N_19806);
nor UO_1318 (O_1318,N_19910,N_19926);
nand UO_1319 (O_1319,N_19896,N_19982);
and UO_1320 (O_1320,N_19907,N_19908);
or UO_1321 (O_1321,N_19863,N_19843);
or UO_1322 (O_1322,N_19947,N_19837);
or UO_1323 (O_1323,N_19949,N_19956);
and UO_1324 (O_1324,N_19829,N_19848);
nand UO_1325 (O_1325,N_19899,N_19936);
and UO_1326 (O_1326,N_19980,N_19812);
nand UO_1327 (O_1327,N_19866,N_19911);
and UO_1328 (O_1328,N_19933,N_19945);
nand UO_1329 (O_1329,N_19936,N_19998);
nand UO_1330 (O_1330,N_19940,N_19897);
nand UO_1331 (O_1331,N_19974,N_19958);
nand UO_1332 (O_1332,N_19992,N_19965);
nand UO_1333 (O_1333,N_19838,N_19999);
nand UO_1334 (O_1334,N_19823,N_19852);
xor UO_1335 (O_1335,N_19990,N_19801);
nor UO_1336 (O_1336,N_19987,N_19907);
and UO_1337 (O_1337,N_19855,N_19961);
and UO_1338 (O_1338,N_19898,N_19842);
nor UO_1339 (O_1339,N_19847,N_19863);
nor UO_1340 (O_1340,N_19831,N_19968);
or UO_1341 (O_1341,N_19834,N_19991);
and UO_1342 (O_1342,N_19897,N_19872);
and UO_1343 (O_1343,N_19999,N_19994);
and UO_1344 (O_1344,N_19819,N_19998);
and UO_1345 (O_1345,N_19899,N_19814);
xnor UO_1346 (O_1346,N_19907,N_19834);
or UO_1347 (O_1347,N_19868,N_19931);
or UO_1348 (O_1348,N_19819,N_19890);
xor UO_1349 (O_1349,N_19924,N_19997);
or UO_1350 (O_1350,N_19836,N_19946);
nor UO_1351 (O_1351,N_19870,N_19910);
and UO_1352 (O_1352,N_19875,N_19976);
xor UO_1353 (O_1353,N_19872,N_19953);
nor UO_1354 (O_1354,N_19927,N_19991);
or UO_1355 (O_1355,N_19997,N_19995);
nor UO_1356 (O_1356,N_19920,N_19870);
or UO_1357 (O_1357,N_19962,N_19842);
xnor UO_1358 (O_1358,N_19852,N_19851);
or UO_1359 (O_1359,N_19823,N_19911);
or UO_1360 (O_1360,N_19933,N_19800);
or UO_1361 (O_1361,N_19965,N_19832);
xor UO_1362 (O_1362,N_19817,N_19928);
nor UO_1363 (O_1363,N_19846,N_19962);
nand UO_1364 (O_1364,N_19882,N_19976);
nand UO_1365 (O_1365,N_19941,N_19865);
nor UO_1366 (O_1366,N_19900,N_19909);
xnor UO_1367 (O_1367,N_19969,N_19809);
or UO_1368 (O_1368,N_19923,N_19998);
nand UO_1369 (O_1369,N_19904,N_19903);
nand UO_1370 (O_1370,N_19923,N_19878);
xnor UO_1371 (O_1371,N_19924,N_19838);
and UO_1372 (O_1372,N_19879,N_19934);
and UO_1373 (O_1373,N_19814,N_19973);
or UO_1374 (O_1374,N_19993,N_19907);
nor UO_1375 (O_1375,N_19968,N_19956);
nor UO_1376 (O_1376,N_19864,N_19866);
and UO_1377 (O_1377,N_19837,N_19878);
and UO_1378 (O_1378,N_19915,N_19815);
nand UO_1379 (O_1379,N_19913,N_19931);
nand UO_1380 (O_1380,N_19979,N_19901);
nor UO_1381 (O_1381,N_19981,N_19816);
nand UO_1382 (O_1382,N_19972,N_19945);
and UO_1383 (O_1383,N_19988,N_19879);
xor UO_1384 (O_1384,N_19820,N_19831);
xnor UO_1385 (O_1385,N_19976,N_19869);
nand UO_1386 (O_1386,N_19823,N_19961);
nand UO_1387 (O_1387,N_19890,N_19956);
nor UO_1388 (O_1388,N_19838,N_19874);
and UO_1389 (O_1389,N_19940,N_19957);
nand UO_1390 (O_1390,N_19825,N_19990);
or UO_1391 (O_1391,N_19986,N_19846);
xor UO_1392 (O_1392,N_19958,N_19968);
nand UO_1393 (O_1393,N_19816,N_19895);
xnor UO_1394 (O_1394,N_19806,N_19904);
nor UO_1395 (O_1395,N_19901,N_19999);
nand UO_1396 (O_1396,N_19941,N_19932);
or UO_1397 (O_1397,N_19966,N_19838);
and UO_1398 (O_1398,N_19885,N_19821);
or UO_1399 (O_1399,N_19880,N_19921);
or UO_1400 (O_1400,N_19815,N_19801);
nand UO_1401 (O_1401,N_19951,N_19998);
xor UO_1402 (O_1402,N_19950,N_19937);
nor UO_1403 (O_1403,N_19853,N_19849);
nand UO_1404 (O_1404,N_19800,N_19984);
nor UO_1405 (O_1405,N_19859,N_19974);
or UO_1406 (O_1406,N_19839,N_19919);
nand UO_1407 (O_1407,N_19999,N_19932);
nand UO_1408 (O_1408,N_19878,N_19955);
and UO_1409 (O_1409,N_19923,N_19829);
or UO_1410 (O_1410,N_19846,N_19968);
xor UO_1411 (O_1411,N_19907,N_19846);
or UO_1412 (O_1412,N_19839,N_19984);
or UO_1413 (O_1413,N_19991,N_19851);
xnor UO_1414 (O_1414,N_19960,N_19974);
and UO_1415 (O_1415,N_19969,N_19971);
nor UO_1416 (O_1416,N_19808,N_19981);
and UO_1417 (O_1417,N_19820,N_19834);
and UO_1418 (O_1418,N_19924,N_19821);
and UO_1419 (O_1419,N_19951,N_19906);
or UO_1420 (O_1420,N_19932,N_19804);
xnor UO_1421 (O_1421,N_19942,N_19976);
nor UO_1422 (O_1422,N_19899,N_19891);
and UO_1423 (O_1423,N_19860,N_19884);
or UO_1424 (O_1424,N_19836,N_19959);
nand UO_1425 (O_1425,N_19883,N_19935);
xor UO_1426 (O_1426,N_19972,N_19874);
nand UO_1427 (O_1427,N_19867,N_19923);
nor UO_1428 (O_1428,N_19906,N_19909);
nor UO_1429 (O_1429,N_19963,N_19807);
nor UO_1430 (O_1430,N_19996,N_19968);
nor UO_1431 (O_1431,N_19986,N_19999);
and UO_1432 (O_1432,N_19858,N_19907);
or UO_1433 (O_1433,N_19918,N_19964);
nor UO_1434 (O_1434,N_19888,N_19856);
nor UO_1435 (O_1435,N_19974,N_19929);
nor UO_1436 (O_1436,N_19841,N_19979);
and UO_1437 (O_1437,N_19880,N_19889);
nand UO_1438 (O_1438,N_19839,N_19994);
nand UO_1439 (O_1439,N_19917,N_19811);
xor UO_1440 (O_1440,N_19919,N_19963);
xnor UO_1441 (O_1441,N_19863,N_19967);
or UO_1442 (O_1442,N_19966,N_19908);
and UO_1443 (O_1443,N_19870,N_19847);
nor UO_1444 (O_1444,N_19976,N_19886);
and UO_1445 (O_1445,N_19803,N_19825);
nand UO_1446 (O_1446,N_19860,N_19842);
nand UO_1447 (O_1447,N_19937,N_19867);
or UO_1448 (O_1448,N_19943,N_19990);
and UO_1449 (O_1449,N_19951,N_19834);
nor UO_1450 (O_1450,N_19853,N_19874);
or UO_1451 (O_1451,N_19872,N_19808);
and UO_1452 (O_1452,N_19993,N_19988);
or UO_1453 (O_1453,N_19972,N_19868);
or UO_1454 (O_1454,N_19804,N_19971);
nand UO_1455 (O_1455,N_19957,N_19810);
nand UO_1456 (O_1456,N_19909,N_19851);
or UO_1457 (O_1457,N_19876,N_19996);
and UO_1458 (O_1458,N_19931,N_19961);
nor UO_1459 (O_1459,N_19912,N_19986);
nor UO_1460 (O_1460,N_19804,N_19898);
and UO_1461 (O_1461,N_19842,N_19857);
nor UO_1462 (O_1462,N_19856,N_19921);
nor UO_1463 (O_1463,N_19951,N_19841);
nor UO_1464 (O_1464,N_19873,N_19938);
nand UO_1465 (O_1465,N_19933,N_19858);
nand UO_1466 (O_1466,N_19849,N_19805);
nor UO_1467 (O_1467,N_19851,N_19971);
xnor UO_1468 (O_1468,N_19988,N_19942);
nand UO_1469 (O_1469,N_19997,N_19800);
and UO_1470 (O_1470,N_19867,N_19865);
nand UO_1471 (O_1471,N_19965,N_19989);
or UO_1472 (O_1472,N_19844,N_19839);
nand UO_1473 (O_1473,N_19953,N_19994);
xnor UO_1474 (O_1474,N_19996,N_19872);
nand UO_1475 (O_1475,N_19878,N_19912);
nor UO_1476 (O_1476,N_19816,N_19835);
xor UO_1477 (O_1477,N_19855,N_19861);
xor UO_1478 (O_1478,N_19956,N_19973);
nor UO_1479 (O_1479,N_19899,N_19866);
and UO_1480 (O_1480,N_19884,N_19946);
or UO_1481 (O_1481,N_19967,N_19986);
nor UO_1482 (O_1482,N_19802,N_19943);
nand UO_1483 (O_1483,N_19957,N_19836);
xor UO_1484 (O_1484,N_19896,N_19866);
and UO_1485 (O_1485,N_19953,N_19894);
and UO_1486 (O_1486,N_19808,N_19995);
and UO_1487 (O_1487,N_19841,N_19895);
and UO_1488 (O_1488,N_19925,N_19928);
or UO_1489 (O_1489,N_19893,N_19890);
nor UO_1490 (O_1490,N_19801,N_19865);
nand UO_1491 (O_1491,N_19908,N_19827);
and UO_1492 (O_1492,N_19856,N_19972);
nor UO_1493 (O_1493,N_19862,N_19913);
nand UO_1494 (O_1494,N_19944,N_19883);
or UO_1495 (O_1495,N_19900,N_19951);
nand UO_1496 (O_1496,N_19927,N_19978);
nor UO_1497 (O_1497,N_19973,N_19899);
or UO_1498 (O_1498,N_19957,N_19988);
nand UO_1499 (O_1499,N_19976,N_19905);
nor UO_1500 (O_1500,N_19991,N_19938);
nand UO_1501 (O_1501,N_19896,N_19819);
and UO_1502 (O_1502,N_19994,N_19960);
or UO_1503 (O_1503,N_19994,N_19901);
nand UO_1504 (O_1504,N_19855,N_19989);
xor UO_1505 (O_1505,N_19887,N_19900);
or UO_1506 (O_1506,N_19915,N_19909);
or UO_1507 (O_1507,N_19945,N_19916);
or UO_1508 (O_1508,N_19821,N_19937);
and UO_1509 (O_1509,N_19848,N_19956);
xnor UO_1510 (O_1510,N_19811,N_19830);
xor UO_1511 (O_1511,N_19861,N_19874);
and UO_1512 (O_1512,N_19924,N_19972);
xnor UO_1513 (O_1513,N_19988,N_19958);
nor UO_1514 (O_1514,N_19936,N_19925);
and UO_1515 (O_1515,N_19851,N_19825);
and UO_1516 (O_1516,N_19811,N_19847);
nor UO_1517 (O_1517,N_19933,N_19872);
nand UO_1518 (O_1518,N_19928,N_19940);
and UO_1519 (O_1519,N_19890,N_19897);
nand UO_1520 (O_1520,N_19855,N_19920);
and UO_1521 (O_1521,N_19932,N_19936);
and UO_1522 (O_1522,N_19831,N_19864);
nor UO_1523 (O_1523,N_19881,N_19989);
and UO_1524 (O_1524,N_19897,N_19881);
xnor UO_1525 (O_1525,N_19914,N_19985);
nand UO_1526 (O_1526,N_19875,N_19863);
nor UO_1527 (O_1527,N_19915,N_19974);
nand UO_1528 (O_1528,N_19833,N_19813);
nor UO_1529 (O_1529,N_19937,N_19933);
nor UO_1530 (O_1530,N_19977,N_19841);
nor UO_1531 (O_1531,N_19895,N_19968);
xnor UO_1532 (O_1532,N_19814,N_19919);
nor UO_1533 (O_1533,N_19811,N_19829);
xnor UO_1534 (O_1534,N_19822,N_19972);
or UO_1535 (O_1535,N_19955,N_19812);
and UO_1536 (O_1536,N_19948,N_19953);
or UO_1537 (O_1537,N_19880,N_19971);
nor UO_1538 (O_1538,N_19971,N_19872);
nand UO_1539 (O_1539,N_19997,N_19996);
nand UO_1540 (O_1540,N_19862,N_19882);
or UO_1541 (O_1541,N_19912,N_19870);
nor UO_1542 (O_1542,N_19909,N_19868);
and UO_1543 (O_1543,N_19915,N_19913);
nor UO_1544 (O_1544,N_19879,N_19997);
nand UO_1545 (O_1545,N_19989,N_19837);
or UO_1546 (O_1546,N_19916,N_19825);
xor UO_1547 (O_1547,N_19904,N_19898);
nand UO_1548 (O_1548,N_19844,N_19811);
or UO_1549 (O_1549,N_19835,N_19969);
nor UO_1550 (O_1550,N_19939,N_19990);
nand UO_1551 (O_1551,N_19805,N_19942);
nand UO_1552 (O_1552,N_19970,N_19861);
or UO_1553 (O_1553,N_19967,N_19926);
nor UO_1554 (O_1554,N_19966,N_19957);
and UO_1555 (O_1555,N_19852,N_19864);
xnor UO_1556 (O_1556,N_19824,N_19945);
xor UO_1557 (O_1557,N_19999,N_19945);
xor UO_1558 (O_1558,N_19846,N_19945);
or UO_1559 (O_1559,N_19900,N_19852);
nand UO_1560 (O_1560,N_19951,N_19821);
nor UO_1561 (O_1561,N_19854,N_19913);
or UO_1562 (O_1562,N_19860,N_19985);
xnor UO_1563 (O_1563,N_19822,N_19893);
nand UO_1564 (O_1564,N_19892,N_19802);
nand UO_1565 (O_1565,N_19971,N_19903);
nor UO_1566 (O_1566,N_19856,N_19967);
and UO_1567 (O_1567,N_19949,N_19922);
or UO_1568 (O_1568,N_19844,N_19847);
nand UO_1569 (O_1569,N_19938,N_19846);
or UO_1570 (O_1570,N_19995,N_19829);
nand UO_1571 (O_1571,N_19865,N_19966);
nand UO_1572 (O_1572,N_19841,N_19812);
nand UO_1573 (O_1573,N_19975,N_19871);
nand UO_1574 (O_1574,N_19824,N_19892);
nor UO_1575 (O_1575,N_19960,N_19961);
nand UO_1576 (O_1576,N_19957,N_19902);
or UO_1577 (O_1577,N_19959,N_19963);
and UO_1578 (O_1578,N_19814,N_19800);
and UO_1579 (O_1579,N_19876,N_19890);
or UO_1580 (O_1580,N_19952,N_19990);
nor UO_1581 (O_1581,N_19999,N_19833);
and UO_1582 (O_1582,N_19869,N_19907);
nand UO_1583 (O_1583,N_19841,N_19844);
xor UO_1584 (O_1584,N_19898,N_19850);
or UO_1585 (O_1585,N_19944,N_19954);
nor UO_1586 (O_1586,N_19947,N_19897);
nor UO_1587 (O_1587,N_19869,N_19956);
nor UO_1588 (O_1588,N_19800,N_19810);
nand UO_1589 (O_1589,N_19993,N_19925);
and UO_1590 (O_1590,N_19866,N_19948);
nor UO_1591 (O_1591,N_19910,N_19943);
nand UO_1592 (O_1592,N_19846,N_19916);
xor UO_1593 (O_1593,N_19942,N_19834);
or UO_1594 (O_1594,N_19920,N_19939);
or UO_1595 (O_1595,N_19965,N_19908);
nand UO_1596 (O_1596,N_19944,N_19926);
or UO_1597 (O_1597,N_19950,N_19925);
xor UO_1598 (O_1598,N_19889,N_19864);
xnor UO_1599 (O_1599,N_19856,N_19982);
and UO_1600 (O_1600,N_19949,N_19977);
and UO_1601 (O_1601,N_19921,N_19829);
nor UO_1602 (O_1602,N_19949,N_19871);
or UO_1603 (O_1603,N_19826,N_19893);
or UO_1604 (O_1604,N_19958,N_19981);
and UO_1605 (O_1605,N_19883,N_19809);
and UO_1606 (O_1606,N_19908,N_19820);
nand UO_1607 (O_1607,N_19915,N_19871);
xnor UO_1608 (O_1608,N_19828,N_19824);
and UO_1609 (O_1609,N_19973,N_19965);
nand UO_1610 (O_1610,N_19871,N_19935);
nor UO_1611 (O_1611,N_19892,N_19879);
and UO_1612 (O_1612,N_19859,N_19830);
or UO_1613 (O_1613,N_19864,N_19971);
nand UO_1614 (O_1614,N_19978,N_19906);
xnor UO_1615 (O_1615,N_19849,N_19958);
xnor UO_1616 (O_1616,N_19837,N_19824);
or UO_1617 (O_1617,N_19802,N_19846);
nor UO_1618 (O_1618,N_19920,N_19966);
nor UO_1619 (O_1619,N_19949,N_19874);
xor UO_1620 (O_1620,N_19971,N_19972);
nand UO_1621 (O_1621,N_19830,N_19933);
nor UO_1622 (O_1622,N_19987,N_19940);
xnor UO_1623 (O_1623,N_19880,N_19847);
nand UO_1624 (O_1624,N_19836,N_19879);
and UO_1625 (O_1625,N_19913,N_19844);
nand UO_1626 (O_1626,N_19983,N_19968);
nand UO_1627 (O_1627,N_19959,N_19970);
xnor UO_1628 (O_1628,N_19863,N_19853);
and UO_1629 (O_1629,N_19902,N_19954);
and UO_1630 (O_1630,N_19867,N_19845);
nand UO_1631 (O_1631,N_19945,N_19975);
nand UO_1632 (O_1632,N_19983,N_19975);
nor UO_1633 (O_1633,N_19906,N_19856);
nand UO_1634 (O_1634,N_19953,N_19971);
nand UO_1635 (O_1635,N_19914,N_19979);
nor UO_1636 (O_1636,N_19815,N_19828);
and UO_1637 (O_1637,N_19837,N_19821);
nor UO_1638 (O_1638,N_19886,N_19987);
nor UO_1639 (O_1639,N_19967,N_19945);
and UO_1640 (O_1640,N_19870,N_19963);
xor UO_1641 (O_1641,N_19852,N_19905);
xor UO_1642 (O_1642,N_19886,N_19978);
nor UO_1643 (O_1643,N_19975,N_19996);
nand UO_1644 (O_1644,N_19910,N_19989);
or UO_1645 (O_1645,N_19883,N_19890);
nand UO_1646 (O_1646,N_19888,N_19920);
or UO_1647 (O_1647,N_19899,N_19938);
or UO_1648 (O_1648,N_19804,N_19813);
nand UO_1649 (O_1649,N_19931,N_19988);
xnor UO_1650 (O_1650,N_19818,N_19940);
xnor UO_1651 (O_1651,N_19864,N_19942);
and UO_1652 (O_1652,N_19866,N_19901);
xnor UO_1653 (O_1653,N_19887,N_19995);
xnor UO_1654 (O_1654,N_19806,N_19907);
nand UO_1655 (O_1655,N_19994,N_19855);
or UO_1656 (O_1656,N_19912,N_19895);
and UO_1657 (O_1657,N_19872,N_19972);
nor UO_1658 (O_1658,N_19819,N_19834);
xor UO_1659 (O_1659,N_19885,N_19901);
nor UO_1660 (O_1660,N_19939,N_19915);
or UO_1661 (O_1661,N_19978,N_19809);
and UO_1662 (O_1662,N_19983,N_19877);
or UO_1663 (O_1663,N_19989,N_19822);
nand UO_1664 (O_1664,N_19968,N_19995);
or UO_1665 (O_1665,N_19878,N_19957);
nand UO_1666 (O_1666,N_19935,N_19981);
or UO_1667 (O_1667,N_19831,N_19921);
or UO_1668 (O_1668,N_19847,N_19829);
xor UO_1669 (O_1669,N_19977,N_19839);
and UO_1670 (O_1670,N_19801,N_19959);
xor UO_1671 (O_1671,N_19867,N_19926);
and UO_1672 (O_1672,N_19814,N_19883);
xor UO_1673 (O_1673,N_19932,N_19912);
nand UO_1674 (O_1674,N_19850,N_19985);
or UO_1675 (O_1675,N_19998,N_19964);
and UO_1676 (O_1676,N_19885,N_19831);
nand UO_1677 (O_1677,N_19908,N_19991);
and UO_1678 (O_1678,N_19884,N_19875);
nand UO_1679 (O_1679,N_19982,N_19921);
and UO_1680 (O_1680,N_19969,N_19813);
and UO_1681 (O_1681,N_19819,N_19899);
xnor UO_1682 (O_1682,N_19959,N_19804);
xor UO_1683 (O_1683,N_19958,N_19868);
xnor UO_1684 (O_1684,N_19962,N_19999);
nor UO_1685 (O_1685,N_19857,N_19856);
nor UO_1686 (O_1686,N_19812,N_19922);
or UO_1687 (O_1687,N_19932,N_19886);
xnor UO_1688 (O_1688,N_19807,N_19918);
or UO_1689 (O_1689,N_19947,N_19999);
or UO_1690 (O_1690,N_19981,N_19895);
nor UO_1691 (O_1691,N_19872,N_19838);
nor UO_1692 (O_1692,N_19876,N_19810);
or UO_1693 (O_1693,N_19987,N_19839);
and UO_1694 (O_1694,N_19917,N_19869);
nor UO_1695 (O_1695,N_19962,N_19919);
xor UO_1696 (O_1696,N_19967,N_19801);
and UO_1697 (O_1697,N_19882,N_19812);
xor UO_1698 (O_1698,N_19867,N_19970);
nor UO_1699 (O_1699,N_19929,N_19855);
nand UO_1700 (O_1700,N_19895,N_19861);
nand UO_1701 (O_1701,N_19959,N_19885);
xor UO_1702 (O_1702,N_19940,N_19951);
and UO_1703 (O_1703,N_19849,N_19830);
or UO_1704 (O_1704,N_19899,N_19804);
xnor UO_1705 (O_1705,N_19828,N_19831);
and UO_1706 (O_1706,N_19960,N_19983);
and UO_1707 (O_1707,N_19966,N_19847);
nand UO_1708 (O_1708,N_19907,N_19807);
nor UO_1709 (O_1709,N_19902,N_19938);
nand UO_1710 (O_1710,N_19921,N_19901);
and UO_1711 (O_1711,N_19911,N_19830);
nand UO_1712 (O_1712,N_19988,N_19941);
nand UO_1713 (O_1713,N_19888,N_19882);
xor UO_1714 (O_1714,N_19987,N_19949);
xnor UO_1715 (O_1715,N_19866,N_19919);
nor UO_1716 (O_1716,N_19913,N_19892);
nor UO_1717 (O_1717,N_19870,N_19990);
xor UO_1718 (O_1718,N_19845,N_19968);
and UO_1719 (O_1719,N_19864,N_19854);
xnor UO_1720 (O_1720,N_19905,N_19977);
or UO_1721 (O_1721,N_19957,N_19846);
or UO_1722 (O_1722,N_19856,N_19835);
or UO_1723 (O_1723,N_19888,N_19851);
and UO_1724 (O_1724,N_19847,N_19833);
xor UO_1725 (O_1725,N_19898,N_19868);
or UO_1726 (O_1726,N_19887,N_19806);
nor UO_1727 (O_1727,N_19893,N_19801);
nor UO_1728 (O_1728,N_19874,N_19964);
nor UO_1729 (O_1729,N_19883,N_19868);
xor UO_1730 (O_1730,N_19910,N_19820);
or UO_1731 (O_1731,N_19821,N_19936);
xor UO_1732 (O_1732,N_19879,N_19877);
xnor UO_1733 (O_1733,N_19809,N_19891);
xor UO_1734 (O_1734,N_19850,N_19995);
nand UO_1735 (O_1735,N_19929,N_19944);
nand UO_1736 (O_1736,N_19891,N_19876);
and UO_1737 (O_1737,N_19858,N_19943);
xor UO_1738 (O_1738,N_19856,N_19959);
nand UO_1739 (O_1739,N_19895,N_19887);
or UO_1740 (O_1740,N_19960,N_19884);
nand UO_1741 (O_1741,N_19929,N_19861);
and UO_1742 (O_1742,N_19858,N_19861);
and UO_1743 (O_1743,N_19915,N_19953);
and UO_1744 (O_1744,N_19916,N_19827);
and UO_1745 (O_1745,N_19932,N_19842);
or UO_1746 (O_1746,N_19830,N_19877);
xnor UO_1747 (O_1747,N_19858,N_19986);
or UO_1748 (O_1748,N_19834,N_19955);
and UO_1749 (O_1749,N_19818,N_19906);
nand UO_1750 (O_1750,N_19962,N_19968);
nand UO_1751 (O_1751,N_19957,N_19958);
nor UO_1752 (O_1752,N_19805,N_19961);
xnor UO_1753 (O_1753,N_19984,N_19935);
xnor UO_1754 (O_1754,N_19802,N_19874);
and UO_1755 (O_1755,N_19870,N_19994);
and UO_1756 (O_1756,N_19956,N_19814);
xnor UO_1757 (O_1757,N_19843,N_19835);
nand UO_1758 (O_1758,N_19964,N_19961);
or UO_1759 (O_1759,N_19816,N_19883);
nand UO_1760 (O_1760,N_19954,N_19914);
nand UO_1761 (O_1761,N_19965,N_19993);
and UO_1762 (O_1762,N_19918,N_19996);
or UO_1763 (O_1763,N_19837,N_19933);
and UO_1764 (O_1764,N_19818,N_19871);
nand UO_1765 (O_1765,N_19909,N_19896);
nor UO_1766 (O_1766,N_19933,N_19845);
nand UO_1767 (O_1767,N_19841,N_19839);
nor UO_1768 (O_1768,N_19903,N_19946);
nor UO_1769 (O_1769,N_19895,N_19953);
xnor UO_1770 (O_1770,N_19801,N_19880);
nand UO_1771 (O_1771,N_19989,N_19982);
xnor UO_1772 (O_1772,N_19996,N_19885);
nand UO_1773 (O_1773,N_19884,N_19955);
nor UO_1774 (O_1774,N_19839,N_19818);
and UO_1775 (O_1775,N_19905,N_19810);
or UO_1776 (O_1776,N_19811,N_19845);
nand UO_1777 (O_1777,N_19984,N_19882);
or UO_1778 (O_1778,N_19989,N_19919);
and UO_1779 (O_1779,N_19823,N_19984);
xor UO_1780 (O_1780,N_19863,N_19900);
nand UO_1781 (O_1781,N_19889,N_19869);
nor UO_1782 (O_1782,N_19919,N_19847);
or UO_1783 (O_1783,N_19913,N_19943);
xnor UO_1784 (O_1784,N_19929,N_19950);
nand UO_1785 (O_1785,N_19855,N_19924);
nor UO_1786 (O_1786,N_19944,N_19872);
and UO_1787 (O_1787,N_19845,N_19944);
xnor UO_1788 (O_1788,N_19987,N_19819);
nand UO_1789 (O_1789,N_19881,N_19836);
nand UO_1790 (O_1790,N_19970,N_19807);
or UO_1791 (O_1791,N_19854,N_19803);
xor UO_1792 (O_1792,N_19826,N_19878);
and UO_1793 (O_1793,N_19867,N_19869);
xor UO_1794 (O_1794,N_19997,N_19810);
and UO_1795 (O_1795,N_19835,N_19900);
nor UO_1796 (O_1796,N_19901,N_19856);
nand UO_1797 (O_1797,N_19822,N_19849);
nand UO_1798 (O_1798,N_19857,N_19964);
or UO_1799 (O_1799,N_19870,N_19850);
xor UO_1800 (O_1800,N_19994,N_19942);
or UO_1801 (O_1801,N_19933,N_19947);
and UO_1802 (O_1802,N_19828,N_19885);
or UO_1803 (O_1803,N_19880,N_19812);
nor UO_1804 (O_1804,N_19915,N_19962);
nand UO_1805 (O_1805,N_19968,N_19910);
or UO_1806 (O_1806,N_19959,N_19890);
xor UO_1807 (O_1807,N_19805,N_19809);
xor UO_1808 (O_1808,N_19846,N_19953);
or UO_1809 (O_1809,N_19858,N_19950);
nor UO_1810 (O_1810,N_19848,N_19984);
xor UO_1811 (O_1811,N_19918,N_19800);
xnor UO_1812 (O_1812,N_19997,N_19847);
nand UO_1813 (O_1813,N_19836,N_19821);
nand UO_1814 (O_1814,N_19979,N_19834);
or UO_1815 (O_1815,N_19843,N_19886);
or UO_1816 (O_1816,N_19828,N_19944);
and UO_1817 (O_1817,N_19828,N_19878);
xor UO_1818 (O_1818,N_19828,N_19971);
or UO_1819 (O_1819,N_19900,N_19931);
xnor UO_1820 (O_1820,N_19955,N_19830);
nor UO_1821 (O_1821,N_19968,N_19973);
and UO_1822 (O_1822,N_19833,N_19839);
xnor UO_1823 (O_1823,N_19808,N_19986);
and UO_1824 (O_1824,N_19908,N_19932);
nor UO_1825 (O_1825,N_19930,N_19880);
nand UO_1826 (O_1826,N_19993,N_19887);
or UO_1827 (O_1827,N_19826,N_19861);
xor UO_1828 (O_1828,N_19942,N_19961);
nor UO_1829 (O_1829,N_19905,N_19970);
and UO_1830 (O_1830,N_19803,N_19928);
and UO_1831 (O_1831,N_19841,N_19842);
nor UO_1832 (O_1832,N_19906,N_19988);
nor UO_1833 (O_1833,N_19877,N_19803);
nand UO_1834 (O_1834,N_19994,N_19854);
or UO_1835 (O_1835,N_19935,N_19899);
or UO_1836 (O_1836,N_19874,N_19813);
and UO_1837 (O_1837,N_19863,N_19998);
and UO_1838 (O_1838,N_19940,N_19906);
and UO_1839 (O_1839,N_19804,N_19866);
and UO_1840 (O_1840,N_19878,N_19952);
xor UO_1841 (O_1841,N_19977,N_19876);
nand UO_1842 (O_1842,N_19995,N_19914);
or UO_1843 (O_1843,N_19919,N_19832);
nand UO_1844 (O_1844,N_19943,N_19844);
nor UO_1845 (O_1845,N_19829,N_19908);
or UO_1846 (O_1846,N_19910,N_19863);
or UO_1847 (O_1847,N_19825,N_19852);
xor UO_1848 (O_1848,N_19880,N_19881);
and UO_1849 (O_1849,N_19815,N_19869);
nor UO_1850 (O_1850,N_19847,N_19888);
nor UO_1851 (O_1851,N_19917,N_19807);
nor UO_1852 (O_1852,N_19911,N_19886);
nand UO_1853 (O_1853,N_19850,N_19958);
or UO_1854 (O_1854,N_19998,N_19960);
nor UO_1855 (O_1855,N_19939,N_19989);
and UO_1856 (O_1856,N_19820,N_19835);
xor UO_1857 (O_1857,N_19852,N_19887);
or UO_1858 (O_1858,N_19965,N_19914);
and UO_1859 (O_1859,N_19998,N_19826);
and UO_1860 (O_1860,N_19931,N_19923);
nand UO_1861 (O_1861,N_19883,N_19919);
or UO_1862 (O_1862,N_19929,N_19860);
nand UO_1863 (O_1863,N_19912,N_19897);
nand UO_1864 (O_1864,N_19963,N_19929);
xor UO_1865 (O_1865,N_19913,N_19991);
or UO_1866 (O_1866,N_19926,N_19950);
and UO_1867 (O_1867,N_19856,N_19850);
nor UO_1868 (O_1868,N_19981,N_19918);
and UO_1869 (O_1869,N_19908,N_19878);
nor UO_1870 (O_1870,N_19814,N_19905);
xor UO_1871 (O_1871,N_19908,N_19914);
and UO_1872 (O_1872,N_19917,N_19818);
and UO_1873 (O_1873,N_19840,N_19873);
xor UO_1874 (O_1874,N_19982,N_19903);
nor UO_1875 (O_1875,N_19945,N_19850);
nor UO_1876 (O_1876,N_19805,N_19971);
nand UO_1877 (O_1877,N_19906,N_19985);
xnor UO_1878 (O_1878,N_19930,N_19905);
and UO_1879 (O_1879,N_19841,N_19994);
nor UO_1880 (O_1880,N_19804,N_19948);
nand UO_1881 (O_1881,N_19971,N_19869);
nor UO_1882 (O_1882,N_19875,N_19919);
xnor UO_1883 (O_1883,N_19897,N_19886);
nor UO_1884 (O_1884,N_19871,N_19804);
nor UO_1885 (O_1885,N_19880,N_19887);
nand UO_1886 (O_1886,N_19991,N_19902);
nand UO_1887 (O_1887,N_19875,N_19997);
nand UO_1888 (O_1888,N_19836,N_19884);
nand UO_1889 (O_1889,N_19897,N_19863);
nand UO_1890 (O_1890,N_19953,N_19847);
or UO_1891 (O_1891,N_19971,N_19848);
nand UO_1892 (O_1892,N_19988,N_19880);
or UO_1893 (O_1893,N_19803,N_19880);
or UO_1894 (O_1894,N_19854,N_19906);
xor UO_1895 (O_1895,N_19815,N_19844);
and UO_1896 (O_1896,N_19809,N_19959);
or UO_1897 (O_1897,N_19915,N_19817);
nor UO_1898 (O_1898,N_19971,N_19928);
xor UO_1899 (O_1899,N_19829,N_19942);
nand UO_1900 (O_1900,N_19848,N_19814);
nor UO_1901 (O_1901,N_19877,N_19836);
and UO_1902 (O_1902,N_19985,N_19904);
and UO_1903 (O_1903,N_19861,N_19869);
nor UO_1904 (O_1904,N_19971,N_19879);
or UO_1905 (O_1905,N_19958,N_19845);
nor UO_1906 (O_1906,N_19919,N_19912);
nand UO_1907 (O_1907,N_19907,N_19836);
nand UO_1908 (O_1908,N_19839,N_19875);
and UO_1909 (O_1909,N_19818,N_19978);
xor UO_1910 (O_1910,N_19843,N_19997);
nand UO_1911 (O_1911,N_19978,N_19937);
xor UO_1912 (O_1912,N_19884,N_19931);
xor UO_1913 (O_1913,N_19803,N_19805);
xnor UO_1914 (O_1914,N_19857,N_19881);
or UO_1915 (O_1915,N_19992,N_19909);
or UO_1916 (O_1916,N_19811,N_19859);
nor UO_1917 (O_1917,N_19808,N_19991);
and UO_1918 (O_1918,N_19866,N_19955);
or UO_1919 (O_1919,N_19869,N_19944);
or UO_1920 (O_1920,N_19864,N_19897);
and UO_1921 (O_1921,N_19831,N_19997);
nand UO_1922 (O_1922,N_19892,N_19926);
and UO_1923 (O_1923,N_19948,N_19933);
and UO_1924 (O_1924,N_19958,N_19972);
nor UO_1925 (O_1925,N_19954,N_19871);
xor UO_1926 (O_1926,N_19814,N_19934);
and UO_1927 (O_1927,N_19845,N_19880);
xor UO_1928 (O_1928,N_19875,N_19836);
nor UO_1929 (O_1929,N_19871,N_19999);
nand UO_1930 (O_1930,N_19981,N_19946);
nand UO_1931 (O_1931,N_19841,N_19883);
or UO_1932 (O_1932,N_19949,N_19967);
and UO_1933 (O_1933,N_19832,N_19813);
xnor UO_1934 (O_1934,N_19858,N_19944);
nor UO_1935 (O_1935,N_19940,N_19877);
xnor UO_1936 (O_1936,N_19899,N_19886);
nand UO_1937 (O_1937,N_19835,N_19928);
or UO_1938 (O_1938,N_19963,N_19954);
or UO_1939 (O_1939,N_19832,N_19992);
or UO_1940 (O_1940,N_19910,N_19980);
nor UO_1941 (O_1941,N_19988,N_19940);
xnor UO_1942 (O_1942,N_19907,N_19902);
or UO_1943 (O_1943,N_19952,N_19817);
nand UO_1944 (O_1944,N_19830,N_19864);
and UO_1945 (O_1945,N_19982,N_19867);
xor UO_1946 (O_1946,N_19925,N_19959);
xnor UO_1947 (O_1947,N_19904,N_19802);
and UO_1948 (O_1948,N_19966,N_19963);
nor UO_1949 (O_1949,N_19896,N_19834);
nand UO_1950 (O_1950,N_19842,N_19835);
nor UO_1951 (O_1951,N_19873,N_19883);
nand UO_1952 (O_1952,N_19813,N_19826);
nand UO_1953 (O_1953,N_19979,N_19890);
xnor UO_1954 (O_1954,N_19963,N_19801);
and UO_1955 (O_1955,N_19905,N_19996);
or UO_1956 (O_1956,N_19930,N_19874);
xor UO_1957 (O_1957,N_19980,N_19808);
nand UO_1958 (O_1958,N_19960,N_19859);
nor UO_1959 (O_1959,N_19949,N_19820);
nor UO_1960 (O_1960,N_19835,N_19855);
nand UO_1961 (O_1961,N_19852,N_19883);
or UO_1962 (O_1962,N_19995,N_19964);
and UO_1963 (O_1963,N_19850,N_19888);
and UO_1964 (O_1964,N_19950,N_19957);
or UO_1965 (O_1965,N_19850,N_19851);
and UO_1966 (O_1966,N_19807,N_19969);
xnor UO_1967 (O_1967,N_19932,N_19858);
nor UO_1968 (O_1968,N_19990,N_19942);
and UO_1969 (O_1969,N_19934,N_19815);
nand UO_1970 (O_1970,N_19835,N_19942);
nand UO_1971 (O_1971,N_19856,N_19827);
nor UO_1972 (O_1972,N_19978,N_19973);
and UO_1973 (O_1973,N_19903,N_19915);
xnor UO_1974 (O_1974,N_19826,N_19808);
nand UO_1975 (O_1975,N_19826,N_19968);
and UO_1976 (O_1976,N_19903,N_19801);
nand UO_1977 (O_1977,N_19924,N_19969);
nand UO_1978 (O_1978,N_19993,N_19954);
or UO_1979 (O_1979,N_19874,N_19867);
nand UO_1980 (O_1980,N_19944,N_19911);
nand UO_1981 (O_1981,N_19979,N_19872);
nand UO_1982 (O_1982,N_19956,N_19864);
nand UO_1983 (O_1983,N_19854,N_19898);
nand UO_1984 (O_1984,N_19832,N_19950);
nand UO_1985 (O_1985,N_19998,N_19917);
nor UO_1986 (O_1986,N_19980,N_19803);
or UO_1987 (O_1987,N_19903,N_19892);
nand UO_1988 (O_1988,N_19945,N_19930);
xor UO_1989 (O_1989,N_19802,N_19926);
and UO_1990 (O_1990,N_19893,N_19919);
nand UO_1991 (O_1991,N_19999,N_19964);
nand UO_1992 (O_1992,N_19942,N_19939);
nand UO_1993 (O_1993,N_19959,N_19927);
xnor UO_1994 (O_1994,N_19838,N_19953);
nor UO_1995 (O_1995,N_19988,N_19837);
nand UO_1996 (O_1996,N_19881,N_19954);
nor UO_1997 (O_1997,N_19928,N_19950);
or UO_1998 (O_1998,N_19854,N_19944);
nand UO_1999 (O_1999,N_19814,N_19859);
and UO_2000 (O_2000,N_19925,N_19984);
nand UO_2001 (O_2001,N_19884,N_19850);
xor UO_2002 (O_2002,N_19963,N_19817);
or UO_2003 (O_2003,N_19983,N_19874);
nand UO_2004 (O_2004,N_19851,N_19860);
nor UO_2005 (O_2005,N_19967,N_19900);
or UO_2006 (O_2006,N_19940,N_19917);
xor UO_2007 (O_2007,N_19808,N_19887);
xnor UO_2008 (O_2008,N_19877,N_19890);
nor UO_2009 (O_2009,N_19969,N_19902);
nor UO_2010 (O_2010,N_19854,N_19808);
xor UO_2011 (O_2011,N_19847,N_19998);
nand UO_2012 (O_2012,N_19954,N_19855);
and UO_2013 (O_2013,N_19833,N_19966);
nor UO_2014 (O_2014,N_19903,N_19846);
xnor UO_2015 (O_2015,N_19828,N_19910);
and UO_2016 (O_2016,N_19928,N_19972);
and UO_2017 (O_2017,N_19825,N_19804);
xor UO_2018 (O_2018,N_19854,N_19974);
and UO_2019 (O_2019,N_19901,N_19967);
nor UO_2020 (O_2020,N_19809,N_19874);
xnor UO_2021 (O_2021,N_19816,N_19864);
nor UO_2022 (O_2022,N_19884,N_19882);
or UO_2023 (O_2023,N_19808,N_19952);
nand UO_2024 (O_2024,N_19901,N_19987);
xnor UO_2025 (O_2025,N_19859,N_19875);
nand UO_2026 (O_2026,N_19959,N_19824);
nor UO_2027 (O_2027,N_19849,N_19840);
and UO_2028 (O_2028,N_19921,N_19899);
xnor UO_2029 (O_2029,N_19835,N_19881);
nand UO_2030 (O_2030,N_19825,N_19847);
nand UO_2031 (O_2031,N_19851,N_19821);
and UO_2032 (O_2032,N_19934,N_19853);
nand UO_2033 (O_2033,N_19897,N_19908);
xor UO_2034 (O_2034,N_19897,N_19992);
nor UO_2035 (O_2035,N_19812,N_19976);
or UO_2036 (O_2036,N_19933,N_19875);
nor UO_2037 (O_2037,N_19895,N_19854);
nor UO_2038 (O_2038,N_19866,N_19944);
or UO_2039 (O_2039,N_19925,N_19869);
nand UO_2040 (O_2040,N_19969,N_19845);
nor UO_2041 (O_2041,N_19912,N_19858);
nor UO_2042 (O_2042,N_19875,N_19927);
xnor UO_2043 (O_2043,N_19881,N_19873);
nand UO_2044 (O_2044,N_19885,N_19801);
nand UO_2045 (O_2045,N_19978,N_19949);
and UO_2046 (O_2046,N_19805,N_19897);
xnor UO_2047 (O_2047,N_19817,N_19993);
or UO_2048 (O_2048,N_19800,N_19836);
and UO_2049 (O_2049,N_19975,N_19911);
nor UO_2050 (O_2050,N_19851,N_19873);
nor UO_2051 (O_2051,N_19941,N_19921);
nand UO_2052 (O_2052,N_19912,N_19871);
nand UO_2053 (O_2053,N_19831,N_19925);
and UO_2054 (O_2054,N_19825,N_19871);
or UO_2055 (O_2055,N_19898,N_19991);
xor UO_2056 (O_2056,N_19898,N_19915);
xor UO_2057 (O_2057,N_19951,N_19949);
nor UO_2058 (O_2058,N_19838,N_19965);
and UO_2059 (O_2059,N_19966,N_19806);
nand UO_2060 (O_2060,N_19821,N_19989);
and UO_2061 (O_2061,N_19903,N_19856);
xnor UO_2062 (O_2062,N_19811,N_19938);
nand UO_2063 (O_2063,N_19861,N_19862);
and UO_2064 (O_2064,N_19850,N_19996);
xor UO_2065 (O_2065,N_19882,N_19836);
nand UO_2066 (O_2066,N_19810,N_19938);
and UO_2067 (O_2067,N_19935,N_19827);
and UO_2068 (O_2068,N_19866,N_19954);
nor UO_2069 (O_2069,N_19887,N_19946);
xnor UO_2070 (O_2070,N_19806,N_19871);
nand UO_2071 (O_2071,N_19879,N_19947);
nor UO_2072 (O_2072,N_19970,N_19883);
or UO_2073 (O_2073,N_19849,N_19892);
or UO_2074 (O_2074,N_19909,N_19800);
nand UO_2075 (O_2075,N_19983,N_19883);
or UO_2076 (O_2076,N_19825,N_19837);
or UO_2077 (O_2077,N_19929,N_19971);
or UO_2078 (O_2078,N_19837,N_19888);
and UO_2079 (O_2079,N_19842,N_19949);
and UO_2080 (O_2080,N_19929,N_19847);
nand UO_2081 (O_2081,N_19881,N_19986);
or UO_2082 (O_2082,N_19994,N_19865);
or UO_2083 (O_2083,N_19849,N_19868);
xor UO_2084 (O_2084,N_19860,N_19994);
and UO_2085 (O_2085,N_19847,N_19931);
nand UO_2086 (O_2086,N_19924,N_19841);
or UO_2087 (O_2087,N_19802,N_19854);
nand UO_2088 (O_2088,N_19810,N_19809);
xnor UO_2089 (O_2089,N_19953,N_19962);
or UO_2090 (O_2090,N_19896,N_19864);
nor UO_2091 (O_2091,N_19912,N_19957);
nand UO_2092 (O_2092,N_19955,N_19841);
and UO_2093 (O_2093,N_19984,N_19836);
nand UO_2094 (O_2094,N_19833,N_19876);
xnor UO_2095 (O_2095,N_19988,N_19861);
xor UO_2096 (O_2096,N_19876,N_19824);
or UO_2097 (O_2097,N_19933,N_19876);
nor UO_2098 (O_2098,N_19961,N_19808);
and UO_2099 (O_2099,N_19954,N_19903);
xor UO_2100 (O_2100,N_19838,N_19841);
nand UO_2101 (O_2101,N_19941,N_19978);
or UO_2102 (O_2102,N_19863,N_19856);
nand UO_2103 (O_2103,N_19870,N_19863);
nor UO_2104 (O_2104,N_19970,N_19863);
xnor UO_2105 (O_2105,N_19909,N_19883);
nor UO_2106 (O_2106,N_19833,N_19871);
nor UO_2107 (O_2107,N_19978,N_19942);
and UO_2108 (O_2108,N_19925,N_19880);
nand UO_2109 (O_2109,N_19831,N_19890);
nand UO_2110 (O_2110,N_19945,N_19827);
or UO_2111 (O_2111,N_19995,N_19953);
xor UO_2112 (O_2112,N_19987,N_19962);
and UO_2113 (O_2113,N_19836,N_19938);
and UO_2114 (O_2114,N_19996,N_19966);
and UO_2115 (O_2115,N_19961,N_19907);
nor UO_2116 (O_2116,N_19978,N_19913);
nand UO_2117 (O_2117,N_19836,N_19864);
xnor UO_2118 (O_2118,N_19950,N_19980);
nor UO_2119 (O_2119,N_19925,N_19864);
or UO_2120 (O_2120,N_19968,N_19834);
xnor UO_2121 (O_2121,N_19974,N_19962);
xor UO_2122 (O_2122,N_19900,N_19866);
nor UO_2123 (O_2123,N_19873,N_19859);
xor UO_2124 (O_2124,N_19834,N_19853);
xnor UO_2125 (O_2125,N_19993,N_19847);
nand UO_2126 (O_2126,N_19993,N_19829);
nand UO_2127 (O_2127,N_19961,N_19994);
nand UO_2128 (O_2128,N_19818,N_19927);
xor UO_2129 (O_2129,N_19919,N_19969);
or UO_2130 (O_2130,N_19875,N_19858);
xor UO_2131 (O_2131,N_19932,N_19863);
and UO_2132 (O_2132,N_19924,N_19865);
and UO_2133 (O_2133,N_19857,N_19956);
or UO_2134 (O_2134,N_19896,N_19883);
xnor UO_2135 (O_2135,N_19844,N_19878);
xnor UO_2136 (O_2136,N_19953,N_19938);
nand UO_2137 (O_2137,N_19940,N_19983);
or UO_2138 (O_2138,N_19897,N_19959);
nor UO_2139 (O_2139,N_19961,N_19874);
nand UO_2140 (O_2140,N_19887,N_19938);
nor UO_2141 (O_2141,N_19986,N_19820);
or UO_2142 (O_2142,N_19816,N_19857);
xor UO_2143 (O_2143,N_19838,N_19847);
nand UO_2144 (O_2144,N_19911,N_19914);
nor UO_2145 (O_2145,N_19874,N_19941);
nor UO_2146 (O_2146,N_19941,N_19824);
or UO_2147 (O_2147,N_19968,N_19936);
or UO_2148 (O_2148,N_19937,N_19814);
xnor UO_2149 (O_2149,N_19838,N_19962);
nand UO_2150 (O_2150,N_19949,N_19829);
xnor UO_2151 (O_2151,N_19843,N_19937);
nor UO_2152 (O_2152,N_19851,N_19872);
nand UO_2153 (O_2153,N_19898,N_19936);
nor UO_2154 (O_2154,N_19805,N_19960);
and UO_2155 (O_2155,N_19919,N_19882);
and UO_2156 (O_2156,N_19943,N_19960);
xor UO_2157 (O_2157,N_19805,N_19827);
nor UO_2158 (O_2158,N_19973,N_19959);
nor UO_2159 (O_2159,N_19922,N_19984);
or UO_2160 (O_2160,N_19828,N_19861);
or UO_2161 (O_2161,N_19901,N_19847);
and UO_2162 (O_2162,N_19890,N_19900);
nand UO_2163 (O_2163,N_19920,N_19935);
and UO_2164 (O_2164,N_19995,N_19881);
xor UO_2165 (O_2165,N_19818,N_19926);
or UO_2166 (O_2166,N_19968,N_19925);
or UO_2167 (O_2167,N_19808,N_19946);
and UO_2168 (O_2168,N_19897,N_19853);
or UO_2169 (O_2169,N_19825,N_19882);
or UO_2170 (O_2170,N_19922,N_19883);
xor UO_2171 (O_2171,N_19975,N_19884);
or UO_2172 (O_2172,N_19847,N_19957);
nand UO_2173 (O_2173,N_19833,N_19968);
or UO_2174 (O_2174,N_19813,N_19979);
or UO_2175 (O_2175,N_19875,N_19876);
nor UO_2176 (O_2176,N_19983,N_19852);
nand UO_2177 (O_2177,N_19867,N_19832);
and UO_2178 (O_2178,N_19876,N_19857);
or UO_2179 (O_2179,N_19944,N_19924);
nor UO_2180 (O_2180,N_19875,N_19965);
xor UO_2181 (O_2181,N_19820,N_19843);
nor UO_2182 (O_2182,N_19974,N_19949);
nor UO_2183 (O_2183,N_19914,N_19980);
or UO_2184 (O_2184,N_19943,N_19917);
nand UO_2185 (O_2185,N_19905,N_19918);
or UO_2186 (O_2186,N_19954,N_19928);
xor UO_2187 (O_2187,N_19951,N_19930);
nor UO_2188 (O_2188,N_19955,N_19877);
xnor UO_2189 (O_2189,N_19972,N_19823);
nand UO_2190 (O_2190,N_19863,N_19943);
and UO_2191 (O_2191,N_19857,N_19902);
or UO_2192 (O_2192,N_19984,N_19933);
nor UO_2193 (O_2193,N_19912,N_19917);
nand UO_2194 (O_2194,N_19876,N_19864);
and UO_2195 (O_2195,N_19908,N_19886);
nor UO_2196 (O_2196,N_19874,N_19993);
xor UO_2197 (O_2197,N_19959,N_19823);
nor UO_2198 (O_2198,N_19894,N_19800);
or UO_2199 (O_2199,N_19933,N_19988);
or UO_2200 (O_2200,N_19908,N_19833);
xor UO_2201 (O_2201,N_19929,N_19919);
and UO_2202 (O_2202,N_19913,N_19887);
and UO_2203 (O_2203,N_19944,N_19942);
xnor UO_2204 (O_2204,N_19914,N_19852);
nor UO_2205 (O_2205,N_19802,N_19994);
and UO_2206 (O_2206,N_19821,N_19981);
or UO_2207 (O_2207,N_19867,N_19991);
xnor UO_2208 (O_2208,N_19885,N_19884);
or UO_2209 (O_2209,N_19804,N_19922);
xor UO_2210 (O_2210,N_19838,N_19840);
nor UO_2211 (O_2211,N_19965,N_19902);
xnor UO_2212 (O_2212,N_19874,N_19986);
xor UO_2213 (O_2213,N_19887,N_19899);
or UO_2214 (O_2214,N_19884,N_19986);
or UO_2215 (O_2215,N_19941,N_19905);
xnor UO_2216 (O_2216,N_19868,N_19801);
and UO_2217 (O_2217,N_19922,N_19997);
nor UO_2218 (O_2218,N_19943,N_19905);
nand UO_2219 (O_2219,N_19848,N_19922);
or UO_2220 (O_2220,N_19957,N_19823);
or UO_2221 (O_2221,N_19977,N_19964);
xnor UO_2222 (O_2222,N_19921,N_19940);
or UO_2223 (O_2223,N_19852,N_19906);
and UO_2224 (O_2224,N_19988,N_19904);
nor UO_2225 (O_2225,N_19824,N_19972);
or UO_2226 (O_2226,N_19884,N_19976);
nand UO_2227 (O_2227,N_19896,N_19835);
xor UO_2228 (O_2228,N_19971,N_19941);
or UO_2229 (O_2229,N_19888,N_19988);
and UO_2230 (O_2230,N_19863,N_19810);
nor UO_2231 (O_2231,N_19968,N_19904);
and UO_2232 (O_2232,N_19990,N_19966);
or UO_2233 (O_2233,N_19973,N_19961);
nor UO_2234 (O_2234,N_19975,N_19822);
nor UO_2235 (O_2235,N_19978,N_19812);
or UO_2236 (O_2236,N_19868,N_19808);
xnor UO_2237 (O_2237,N_19994,N_19959);
nor UO_2238 (O_2238,N_19909,N_19999);
xor UO_2239 (O_2239,N_19999,N_19941);
nor UO_2240 (O_2240,N_19806,N_19938);
nor UO_2241 (O_2241,N_19819,N_19972);
xnor UO_2242 (O_2242,N_19834,N_19995);
or UO_2243 (O_2243,N_19867,N_19905);
xor UO_2244 (O_2244,N_19906,N_19901);
or UO_2245 (O_2245,N_19946,N_19975);
xnor UO_2246 (O_2246,N_19945,N_19899);
xor UO_2247 (O_2247,N_19988,N_19859);
or UO_2248 (O_2248,N_19920,N_19950);
nand UO_2249 (O_2249,N_19954,N_19951);
and UO_2250 (O_2250,N_19810,N_19853);
or UO_2251 (O_2251,N_19987,N_19854);
nand UO_2252 (O_2252,N_19837,N_19830);
or UO_2253 (O_2253,N_19883,N_19853);
and UO_2254 (O_2254,N_19820,N_19976);
and UO_2255 (O_2255,N_19888,N_19945);
xor UO_2256 (O_2256,N_19938,N_19879);
nand UO_2257 (O_2257,N_19972,N_19899);
and UO_2258 (O_2258,N_19979,N_19986);
or UO_2259 (O_2259,N_19869,N_19924);
xor UO_2260 (O_2260,N_19851,N_19939);
xor UO_2261 (O_2261,N_19956,N_19803);
xor UO_2262 (O_2262,N_19871,N_19995);
xor UO_2263 (O_2263,N_19864,N_19845);
nor UO_2264 (O_2264,N_19867,N_19915);
or UO_2265 (O_2265,N_19844,N_19959);
xnor UO_2266 (O_2266,N_19876,N_19999);
nor UO_2267 (O_2267,N_19859,N_19930);
and UO_2268 (O_2268,N_19808,N_19978);
nor UO_2269 (O_2269,N_19819,N_19869);
or UO_2270 (O_2270,N_19958,N_19863);
or UO_2271 (O_2271,N_19922,N_19929);
or UO_2272 (O_2272,N_19892,N_19891);
or UO_2273 (O_2273,N_19980,N_19833);
xor UO_2274 (O_2274,N_19887,N_19925);
or UO_2275 (O_2275,N_19891,N_19835);
and UO_2276 (O_2276,N_19930,N_19963);
nand UO_2277 (O_2277,N_19899,N_19912);
nand UO_2278 (O_2278,N_19989,N_19884);
nand UO_2279 (O_2279,N_19892,N_19952);
nand UO_2280 (O_2280,N_19905,N_19972);
or UO_2281 (O_2281,N_19885,N_19832);
xnor UO_2282 (O_2282,N_19962,N_19930);
and UO_2283 (O_2283,N_19955,N_19949);
nor UO_2284 (O_2284,N_19805,N_19884);
xor UO_2285 (O_2285,N_19925,N_19979);
nand UO_2286 (O_2286,N_19809,N_19818);
xor UO_2287 (O_2287,N_19989,N_19834);
nand UO_2288 (O_2288,N_19814,N_19980);
nand UO_2289 (O_2289,N_19886,N_19906);
or UO_2290 (O_2290,N_19965,N_19887);
xnor UO_2291 (O_2291,N_19829,N_19872);
xnor UO_2292 (O_2292,N_19973,N_19812);
xnor UO_2293 (O_2293,N_19884,N_19824);
nor UO_2294 (O_2294,N_19966,N_19826);
and UO_2295 (O_2295,N_19863,N_19836);
or UO_2296 (O_2296,N_19882,N_19814);
and UO_2297 (O_2297,N_19823,N_19889);
or UO_2298 (O_2298,N_19840,N_19874);
and UO_2299 (O_2299,N_19896,N_19824);
nand UO_2300 (O_2300,N_19876,N_19895);
nand UO_2301 (O_2301,N_19902,N_19924);
nor UO_2302 (O_2302,N_19862,N_19851);
or UO_2303 (O_2303,N_19928,N_19996);
nor UO_2304 (O_2304,N_19879,N_19983);
xor UO_2305 (O_2305,N_19961,N_19848);
xnor UO_2306 (O_2306,N_19954,N_19882);
nor UO_2307 (O_2307,N_19965,N_19976);
xor UO_2308 (O_2308,N_19986,N_19857);
nor UO_2309 (O_2309,N_19906,N_19931);
xnor UO_2310 (O_2310,N_19882,N_19904);
and UO_2311 (O_2311,N_19975,N_19986);
and UO_2312 (O_2312,N_19807,N_19978);
or UO_2313 (O_2313,N_19963,N_19828);
or UO_2314 (O_2314,N_19832,N_19914);
nor UO_2315 (O_2315,N_19824,N_19977);
xnor UO_2316 (O_2316,N_19873,N_19995);
and UO_2317 (O_2317,N_19862,N_19842);
and UO_2318 (O_2318,N_19997,N_19919);
and UO_2319 (O_2319,N_19957,N_19970);
or UO_2320 (O_2320,N_19978,N_19806);
nand UO_2321 (O_2321,N_19872,N_19952);
or UO_2322 (O_2322,N_19827,N_19900);
and UO_2323 (O_2323,N_19923,N_19846);
and UO_2324 (O_2324,N_19988,N_19972);
or UO_2325 (O_2325,N_19824,N_19881);
and UO_2326 (O_2326,N_19947,N_19964);
or UO_2327 (O_2327,N_19976,N_19823);
or UO_2328 (O_2328,N_19956,N_19962);
nor UO_2329 (O_2329,N_19883,N_19994);
or UO_2330 (O_2330,N_19885,N_19973);
xor UO_2331 (O_2331,N_19815,N_19857);
nor UO_2332 (O_2332,N_19963,N_19869);
or UO_2333 (O_2333,N_19831,N_19886);
or UO_2334 (O_2334,N_19878,N_19901);
nor UO_2335 (O_2335,N_19968,N_19950);
nand UO_2336 (O_2336,N_19804,N_19895);
nor UO_2337 (O_2337,N_19807,N_19816);
nor UO_2338 (O_2338,N_19891,N_19966);
xor UO_2339 (O_2339,N_19811,N_19956);
or UO_2340 (O_2340,N_19852,N_19940);
nor UO_2341 (O_2341,N_19941,N_19861);
nor UO_2342 (O_2342,N_19899,N_19807);
xor UO_2343 (O_2343,N_19831,N_19844);
and UO_2344 (O_2344,N_19843,N_19841);
xnor UO_2345 (O_2345,N_19812,N_19832);
nor UO_2346 (O_2346,N_19817,N_19851);
nand UO_2347 (O_2347,N_19935,N_19954);
nand UO_2348 (O_2348,N_19963,N_19970);
nand UO_2349 (O_2349,N_19952,N_19947);
and UO_2350 (O_2350,N_19982,N_19846);
nor UO_2351 (O_2351,N_19898,N_19805);
nor UO_2352 (O_2352,N_19844,N_19908);
xor UO_2353 (O_2353,N_19806,N_19869);
nor UO_2354 (O_2354,N_19896,N_19991);
nor UO_2355 (O_2355,N_19924,N_19953);
nand UO_2356 (O_2356,N_19929,N_19992);
and UO_2357 (O_2357,N_19884,N_19959);
nand UO_2358 (O_2358,N_19895,N_19932);
nor UO_2359 (O_2359,N_19858,N_19963);
or UO_2360 (O_2360,N_19959,N_19946);
nand UO_2361 (O_2361,N_19819,N_19971);
and UO_2362 (O_2362,N_19867,N_19884);
nor UO_2363 (O_2363,N_19936,N_19934);
or UO_2364 (O_2364,N_19856,N_19872);
nand UO_2365 (O_2365,N_19860,N_19949);
nand UO_2366 (O_2366,N_19859,N_19848);
nor UO_2367 (O_2367,N_19855,N_19959);
or UO_2368 (O_2368,N_19973,N_19901);
xor UO_2369 (O_2369,N_19920,N_19803);
nor UO_2370 (O_2370,N_19974,N_19912);
xnor UO_2371 (O_2371,N_19981,N_19840);
xnor UO_2372 (O_2372,N_19835,N_19811);
or UO_2373 (O_2373,N_19801,N_19989);
and UO_2374 (O_2374,N_19903,N_19828);
nor UO_2375 (O_2375,N_19944,N_19947);
and UO_2376 (O_2376,N_19990,N_19836);
nand UO_2377 (O_2377,N_19935,N_19928);
nand UO_2378 (O_2378,N_19862,N_19918);
nand UO_2379 (O_2379,N_19901,N_19867);
nand UO_2380 (O_2380,N_19893,N_19876);
or UO_2381 (O_2381,N_19823,N_19993);
nor UO_2382 (O_2382,N_19825,N_19913);
and UO_2383 (O_2383,N_19841,N_19942);
or UO_2384 (O_2384,N_19894,N_19920);
xor UO_2385 (O_2385,N_19906,N_19844);
nand UO_2386 (O_2386,N_19845,N_19810);
or UO_2387 (O_2387,N_19914,N_19999);
or UO_2388 (O_2388,N_19852,N_19855);
and UO_2389 (O_2389,N_19996,N_19962);
nand UO_2390 (O_2390,N_19904,N_19873);
nand UO_2391 (O_2391,N_19820,N_19901);
nor UO_2392 (O_2392,N_19986,N_19955);
nor UO_2393 (O_2393,N_19841,N_19950);
xnor UO_2394 (O_2394,N_19969,N_19926);
or UO_2395 (O_2395,N_19867,N_19854);
nor UO_2396 (O_2396,N_19889,N_19995);
nor UO_2397 (O_2397,N_19981,N_19818);
xor UO_2398 (O_2398,N_19806,N_19849);
nand UO_2399 (O_2399,N_19958,N_19944);
and UO_2400 (O_2400,N_19900,N_19915);
nor UO_2401 (O_2401,N_19945,N_19996);
xnor UO_2402 (O_2402,N_19971,N_19935);
xor UO_2403 (O_2403,N_19980,N_19897);
xor UO_2404 (O_2404,N_19951,N_19801);
and UO_2405 (O_2405,N_19946,N_19904);
nand UO_2406 (O_2406,N_19979,N_19909);
xor UO_2407 (O_2407,N_19844,N_19897);
xor UO_2408 (O_2408,N_19822,N_19863);
and UO_2409 (O_2409,N_19818,N_19932);
xor UO_2410 (O_2410,N_19913,N_19848);
and UO_2411 (O_2411,N_19807,N_19855);
and UO_2412 (O_2412,N_19909,N_19991);
or UO_2413 (O_2413,N_19869,N_19899);
nand UO_2414 (O_2414,N_19852,N_19816);
and UO_2415 (O_2415,N_19981,N_19971);
xnor UO_2416 (O_2416,N_19872,N_19881);
or UO_2417 (O_2417,N_19859,N_19963);
or UO_2418 (O_2418,N_19982,N_19925);
or UO_2419 (O_2419,N_19848,N_19864);
or UO_2420 (O_2420,N_19811,N_19889);
xnor UO_2421 (O_2421,N_19935,N_19972);
nand UO_2422 (O_2422,N_19879,N_19867);
or UO_2423 (O_2423,N_19956,N_19842);
or UO_2424 (O_2424,N_19917,N_19985);
nand UO_2425 (O_2425,N_19916,N_19892);
nor UO_2426 (O_2426,N_19842,N_19897);
xor UO_2427 (O_2427,N_19884,N_19889);
xnor UO_2428 (O_2428,N_19978,N_19804);
nor UO_2429 (O_2429,N_19860,N_19888);
nor UO_2430 (O_2430,N_19983,N_19946);
nor UO_2431 (O_2431,N_19889,N_19901);
nor UO_2432 (O_2432,N_19819,N_19959);
and UO_2433 (O_2433,N_19825,N_19827);
and UO_2434 (O_2434,N_19910,N_19887);
xnor UO_2435 (O_2435,N_19995,N_19815);
nand UO_2436 (O_2436,N_19939,N_19936);
or UO_2437 (O_2437,N_19898,N_19937);
nor UO_2438 (O_2438,N_19826,N_19851);
xnor UO_2439 (O_2439,N_19826,N_19926);
xor UO_2440 (O_2440,N_19823,N_19983);
or UO_2441 (O_2441,N_19963,N_19998);
and UO_2442 (O_2442,N_19903,N_19945);
nor UO_2443 (O_2443,N_19864,N_19847);
xnor UO_2444 (O_2444,N_19942,N_19812);
nor UO_2445 (O_2445,N_19981,N_19851);
nand UO_2446 (O_2446,N_19971,N_19844);
xnor UO_2447 (O_2447,N_19812,N_19953);
nand UO_2448 (O_2448,N_19944,N_19875);
or UO_2449 (O_2449,N_19809,N_19962);
nand UO_2450 (O_2450,N_19968,N_19947);
or UO_2451 (O_2451,N_19990,N_19956);
xnor UO_2452 (O_2452,N_19974,N_19899);
and UO_2453 (O_2453,N_19880,N_19857);
nand UO_2454 (O_2454,N_19927,N_19966);
nand UO_2455 (O_2455,N_19969,N_19818);
nor UO_2456 (O_2456,N_19828,N_19897);
or UO_2457 (O_2457,N_19874,N_19880);
and UO_2458 (O_2458,N_19957,N_19999);
or UO_2459 (O_2459,N_19907,N_19881);
nor UO_2460 (O_2460,N_19844,N_19800);
xnor UO_2461 (O_2461,N_19917,N_19979);
and UO_2462 (O_2462,N_19818,N_19995);
and UO_2463 (O_2463,N_19960,N_19970);
nand UO_2464 (O_2464,N_19993,N_19916);
nor UO_2465 (O_2465,N_19923,N_19920);
nand UO_2466 (O_2466,N_19922,N_19851);
or UO_2467 (O_2467,N_19903,N_19826);
nor UO_2468 (O_2468,N_19981,N_19800);
and UO_2469 (O_2469,N_19961,N_19899);
or UO_2470 (O_2470,N_19926,N_19976);
xnor UO_2471 (O_2471,N_19969,N_19853);
nand UO_2472 (O_2472,N_19851,N_19942);
and UO_2473 (O_2473,N_19956,N_19980);
xnor UO_2474 (O_2474,N_19876,N_19948);
xnor UO_2475 (O_2475,N_19888,N_19807);
or UO_2476 (O_2476,N_19919,N_19932);
and UO_2477 (O_2477,N_19991,N_19863);
and UO_2478 (O_2478,N_19805,N_19926);
or UO_2479 (O_2479,N_19882,N_19803);
nor UO_2480 (O_2480,N_19803,N_19915);
nand UO_2481 (O_2481,N_19810,N_19850);
xnor UO_2482 (O_2482,N_19918,N_19866);
xor UO_2483 (O_2483,N_19827,N_19884);
and UO_2484 (O_2484,N_19912,N_19876);
nor UO_2485 (O_2485,N_19815,N_19901);
xor UO_2486 (O_2486,N_19999,N_19873);
nor UO_2487 (O_2487,N_19919,N_19881);
or UO_2488 (O_2488,N_19984,N_19801);
xor UO_2489 (O_2489,N_19954,N_19991);
and UO_2490 (O_2490,N_19866,N_19881);
nand UO_2491 (O_2491,N_19928,N_19931);
nand UO_2492 (O_2492,N_19891,N_19814);
xnor UO_2493 (O_2493,N_19810,N_19890);
nand UO_2494 (O_2494,N_19940,N_19896);
or UO_2495 (O_2495,N_19932,N_19994);
and UO_2496 (O_2496,N_19929,N_19850);
nand UO_2497 (O_2497,N_19877,N_19854);
xnor UO_2498 (O_2498,N_19892,N_19960);
nor UO_2499 (O_2499,N_19944,N_19802);
endmodule