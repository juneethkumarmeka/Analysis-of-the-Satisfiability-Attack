module basic_500_3000_500_40_levels_2xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nor U0 (N_0,In_480,In_446);
or U1 (N_1,In_200,In_283);
or U2 (N_2,In_67,In_358);
nor U3 (N_3,In_222,In_389);
nor U4 (N_4,In_455,In_101);
and U5 (N_5,In_125,In_103);
and U6 (N_6,In_193,In_47);
or U7 (N_7,In_132,In_366);
or U8 (N_8,In_292,In_403);
nor U9 (N_9,In_196,In_182);
nor U10 (N_10,In_391,In_40);
nor U11 (N_11,In_102,In_170);
and U12 (N_12,In_290,In_225);
and U13 (N_13,In_160,In_422);
xor U14 (N_14,In_487,In_38);
or U15 (N_15,In_398,In_131);
nand U16 (N_16,In_489,In_134);
and U17 (N_17,In_232,In_151);
nand U18 (N_18,In_167,In_371);
xor U19 (N_19,In_337,In_89);
or U20 (N_20,In_43,In_338);
nor U21 (N_21,In_297,In_479);
and U22 (N_22,In_7,In_359);
or U23 (N_23,In_64,In_344);
or U24 (N_24,In_1,In_330);
or U25 (N_25,In_60,In_17);
or U26 (N_26,In_152,In_115);
nor U27 (N_27,In_255,In_381);
nor U28 (N_28,In_8,In_208);
nor U29 (N_29,In_28,In_133);
and U30 (N_30,In_155,In_448);
or U31 (N_31,In_173,In_25);
nor U32 (N_32,In_267,In_294);
and U33 (N_33,In_457,In_444);
nand U34 (N_34,In_246,In_124);
and U35 (N_35,In_185,In_368);
and U36 (N_36,In_62,In_150);
nand U37 (N_37,In_51,In_107);
and U38 (N_38,In_194,In_270);
nand U39 (N_39,In_135,In_295);
nand U40 (N_40,In_498,In_276);
nand U41 (N_41,In_471,In_78);
nand U42 (N_42,In_311,In_187);
nor U43 (N_43,In_254,In_15);
or U44 (N_44,In_401,In_443);
and U45 (N_45,In_179,In_220);
nand U46 (N_46,In_218,In_321);
nand U47 (N_47,In_251,In_5);
nor U48 (N_48,In_24,In_203);
and U49 (N_49,In_215,In_53);
nor U50 (N_50,In_13,In_345);
nor U51 (N_51,In_360,In_104);
nand U52 (N_52,In_109,In_221);
nor U53 (N_53,In_364,In_326);
nor U54 (N_54,In_416,In_273);
nand U55 (N_55,In_198,In_259);
or U56 (N_56,In_219,In_165);
and U57 (N_57,In_91,In_210);
nand U58 (N_58,In_212,In_450);
and U59 (N_59,In_404,In_305);
and U60 (N_60,In_98,In_23);
or U61 (N_61,In_442,In_306);
nor U62 (N_62,In_61,In_117);
and U63 (N_63,In_320,In_148);
and U64 (N_64,In_417,In_88);
nand U65 (N_65,In_296,In_138);
and U66 (N_66,In_315,In_157);
nand U67 (N_67,In_57,In_411);
nor U68 (N_68,In_237,In_226);
or U69 (N_69,In_0,In_18);
or U70 (N_70,In_146,In_482);
nor U71 (N_71,In_129,In_153);
nor U72 (N_72,In_385,In_94);
or U73 (N_73,In_235,In_491);
and U74 (N_74,In_264,In_477);
and U75 (N_75,In_463,In_488);
or U76 (N_76,N_0,In_351);
xor U77 (N_77,N_70,In_348);
nor U78 (N_78,In_189,In_4);
nor U79 (N_79,N_45,In_263);
nor U80 (N_80,In_402,In_336);
nor U81 (N_81,In_32,In_37);
or U82 (N_82,In_497,N_46);
nor U83 (N_83,In_393,In_406);
or U84 (N_84,In_353,In_298);
and U85 (N_85,In_286,In_407);
and U86 (N_86,In_373,In_340);
nand U87 (N_87,In_245,In_44);
nor U88 (N_88,In_478,In_303);
nand U89 (N_89,In_121,In_58);
and U90 (N_90,In_192,In_413);
xnor U91 (N_91,N_52,N_34);
nand U92 (N_92,In_425,In_269);
or U93 (N_93,In_204,In_207);
or U94 (N_94,In_361,N_19);
and U95 (N_95,In_171,In_45);
nand U96 (N_96,In_438,N_68);
and U97 (N_97,In_378,In_106);
and U98 (N_98,In_395,In_241);
nand U99 (N_99,In_445,N_14);
and U100 (N_100,In_352,N_2);
or U101 (N_101,In_56,In_357);
and U102 (N_102,N_39,In_486);
nand U103 (N_103,In_289,N_67);
or U104 (N_104,In_470,In_92);
nor U105 (N_105,In_496,In_467);
and U106 (N_106,In_48,In_33);
nand U107 (N_107,N_30,In_343);
or U108 (N_108,In_327,In_166);
and U109 (N_109,In_396,In_287);
nor U110 (N_110,In_257,In_128);
nor U111 (N_111,In_399,In_316);
nand U112 (N_112,In_113,In_213);
nand U113 (N_113,In_265,N_51);
or U114 (N_114,In_71,In_2);
and U115 (N_115,In_30,N_5);
nor U116 (N_116,In_97,In_461);
nor U117 (N_117,N_47,In_432);
nor U118 (N_118,In_145,In_464);
nor U119 (N_119,In_469,N_65);
nor U120 (N_120,In_239,In_142);
or U121 (N_121,In_325,In_21);
and U122 (N_122,N_12,In_177);
and U123 (N_123,N_27,In_79);
and U124 (N_124,In_85,In_191);
and U125 (N_125,In_184,In_392);
and U126 (N_126,N_37,In_231);
or U127 (N_127,In_211,In_383);
nor U128 (N_128,In_492,In_230);
nor U129 (N_129,In_427,N_24);
or U130 (N_130,In_346,In_449);
and U131 (N_131,In_453,N_32);
nor U132 (N_132,In_332,In_388);
nand U133 (N_133,In_280,In_119);
or U134 (N_134,N_28,In_268);
nor U135 (N_135,In_339,N_21);
and U136 (N_136,In_175,In_68);
and U137 (N_137,In_136,In_77);
nand U138 (N_138,N_8,In_195);
or U139 (N_139,In_462,In_281);
nor U140 (N_140,In_460,N_3);
nor U141 (N_141,In_39,N_16);
nand U142 (N_142,N_74,In_390);
or U143 (N_143,In_247,In_279);
nor U144 (N_144,In_374,In_55);
or U145 (N_145,N_40,In_139);
or U146 (N_146,In_242,N_48);
and U147 (N_147,In_307,In_329);
nand U148 (N_148,In_258,In_437);
and U149 (N_149,N_17,In_334);
nor U150 (N_150,N_86,In_410);
nor U151 (N_151,In_190,In_441);
and U152 (N_152,N_106,In_349);
nor U153 (N_153,In_253,In_228);
and U154 (N_154,In_217,N_101);
or U155 (N_155,N_77,In_156);
nor U156 (N_156,In_6,N_136);
nand U157 (N_157,N_132,In_436);
and U158 (N_158,In_154,In_485);
or U159 (N_159,In_110,N_29);
nand U160 (N_160,N_149,N_130);
nor U161 (N_161,N_129,In_111);
xnor U162 (N_162,N_99,In_319);
nand U163 (N_163,In_476,In_172);
nand U164 (N_164,In_481,N_102);
or U165 (N_165,N_127,In_274);
and U166 (N_166,N_71,In_66);
or U167 (N_167,In_468,In_69);
xnor U168 (N_168,N_58,In_178);
nand U169 (N_169,In_299,In_309);
nand U170 (N_170,In_452,In_169);
and U171 (N_171,In_31,In_342);
nor U172 (N_172,In_168,In_466);
or U173 (N_173,In_494,In_261);
nor U174 (N_174,In_293,In_424);
nand U175 (N_175,In_302,In_84);
or U176 (N_176,In_243,In_147);
nand U177 (N_177,In_414,N_128);
or U178 (N_178,N_1,In_14);
nor U179 (N_179,N_54,In_300);
or U180 (N_180,N_89,In_206);
nand U181 (N_181,In_74,N_80);
or U182 (N_182,N_35,N_22);
nor U183 (N_183,In_236,In_421);
and U184 (N_184,In_250,In_161);
and U185 (N_185,N_85,N_138);
nand U186 (N_186,N_126,N_118);
or U187 (N_187,In_186,In_408);
nor U188 (N_188,In_380,In_419);
nor U189 (N_189,In_181,N_81);
or U190 (N_190,In_188,N_83);
nor U191 (N_191,In_341,N_100);
or U192 (N_192,In_35,N_142);
or U193 (N_193,In_63,In_318);
nor U194 (N_194,In_127,N_49);
nand U195 (N_195,In_42,In_256);
and U196 (N_196,In_46,In_116);
nor U197 (N_197,In_301,N_18);
nand U198 (N_198,In_130,N_144);
nor U199 (N_199,In_123,In_99);
and U200 (N_200,In_75,N_145);
and U201 (N_201,In_426,In_429);
and U202 (N_202,In_205,In_209);
nand U203 (N_203,In_122,In_499);
nor U204 (N_204,In_52,N_15);
and U205 (N_205,In_288,In_176);
and U206 (N_206,In_137,N_4);
nand U207 (N_207,In_400,N_66);
or U208 (N_208,In_65,In_365);
nand U209 (N_209,In_54,N_38);
nor U210 (N_210,In_224,In_22);
or U211 (N_211,In_120,In_379);
nor U212 (N_212,N_146,In_376);
and U213 (N_213,N_69,In_83);
nand U214 (N_214,In_11,In_314);
or U215 (N_215,In_362,In_227);
or U216 (N_216,In_394,In_451);
or U217 (N_217,N_61,In_459);
or U218 (N_218,N_112,In_95);
nand U219 (N_219,In_397,N_137);
nor U220 (N_220,In_335,N_96);
and U221 (N_221,In_143,In_483);
or U222 (N_222,In_439,In_275);
or U223 (N_223,N_91,In_412);
nor U224 (N_224,N_50,N_64);
nand U225 (N_225,N_171,In_323);
nand U226 (N_226,In_199,N_107);
nand U227 (N_227,In_3,N_151);
or U228 (N_228,In_308,N_214);
and U229 (N_229,In_282,N_199);
nor U230 (N_230,In_105,N_147);
or U231 (N_231,In_9,N_11);
nand U232 (N_232,In_72,N_150);
nand U233 (N_233,In_159,N_53);
or U234 (N_234,N_43,N_159);
or U235 (N_235,In_214,N_203);
and U236 (N_236,N_93,N_103);
nor U237 (N_237,In_440,In_141);
and U238 (N_238,N_75,In_456);
xnor U239 (N_239,N_211,N_41);
nor U240 (N_240,In_114,In_272);
and U241 (N_241,In_447,N_161);
and U242 (N_242,In_409,In_473);
nand U243 (N_243,N_206,N_44);
nor U244 (N_244,In_80,In_29);
or U245 (N_245,N_208,In_370);
and U246 (N_246,N_182,N_201);
and U247 (N_247,In_108,N_215);
nand U248 (N_248,N_25,N_36);
nor U249 (N_249,N_176,N_148);
and U250 (N_250,In_118,In_197);
and U251 (N_251,In_73,N_72);
nand U252 (N_252,N_42,N_82);
and U253 (N_253,N_196,N_57);
nand U254 (N_254,In_495,N_59);
nand U255 (N_255,N_23,N_180);
nor U256 (N_256,In_87,N_205);
or U257 (N_257,N_200,N_60);
xnor U258 (N_258,In_331,In_34);
nand U259 (N_259,In_201,In_284);
or U260 (N_260,N_153,N_220);
and U261 (N_261,N_90,In_50);
or U262 (N_262,In_100,N_116);
and U263 (N_263,N_97,In_82);
nand U264 (N_264,In_183,In_70);
and U265 (N_265,N_179,In_36);
nand U266 (N_266,In_180,N_6);
and U267 (N_267,N_192,N_56);
nor U268 (N_268,N_139,In_355);
and U269 (N_269,In_86,In_10);
nor U270 (N_270,N_221,N_155);
or U271 (N_271,N_10,N_131);
and U272 (N_272,In_140,In_271);
and U273 (N_273,In_262,N_135);
or U274 (N_274,N_123,N_168);
nor U275 (N_275,N_113,In_405);
nor U276 (N_276,N_198,N_186);
and U277 (N_277,N_117,In_252);
nand U278 (N_278,N_163,N_207);
or U279 (N_279,In_285,N_219);
and U280 (N_280,N_189,N_187);
nand U281 (N_281,In_20,In_313);
nand U282 (N_282,N_78,In_423);
nand U283 (N_283,In_350,N_156);
or U284 (N_284,N_178,N_63);
and U285 (N_285,N_183,N_95);
or U286 (N_286,In_12,N_193);
or U287 (N_287,In_266,In_312);
nor U288 (N_288,In_433,In_163);
nand U289 (N_289,In_244,N_216);
and U290 (N_290,In_328,N_224);
nand U291 (N_291,In_26,N_191);
or U292 (N_292,In_278,N_158);
xor U293 (N_293,In_216,In_310);
or U294 (N_294,N_114,In_490);
nor U295 (N_295,N_104,N_194);
xnor U296 (N_296,In_484,In_304);
or U297 (N_297,In_356,In_164);
xor U298 (N_298,In_49,In_415);
nand U299 (N_299,In_126,In_435);
or U300 (N_300,N_141,N_164);
and U301 (N_301,N_284,N_202);
or U302 (N_302,N_247,In_27);
nor U303 (N_303,N_209,N_291);
nand U304 (N_304,N_280,N_249);
xnor U305 (N_305,In_317,N_231);
nor U306 (N_306,N_288,N_293);
nand U307 (N_307,N_223,N_267);
or U308 (N_308,N_84,N_258);
xnor U309 (N_309,N_275,N_253);
nor U310 (N_310,N_261,In_249);
nand U311 (N_311,In_322,In_458);
xor U312 (N_312,N_55,In_41);
nand U313 (N_313,N_110,N_279);
and U314 (N_314,N_268,In_367);
nor U315 (N_315,N_264,N_184);
or U316 (N_316,N_259,N_143);
and U317 (N_317,N_277,In_93);
nor U318 (N_318,In_384,N_98);
and U319 (N_319,In_162,N_140);
nor U320 (N_320,In_96,N_181);
and U321 (N_321,N_166,N_266);
and U322 (N_322,N_230,N_297);
nand U323 (N_323,In_363,N_238);
nor U324 (N_324,N_262,In_431);
or U325 (N_325,N_119,In_333);
or U326 (N_326,In_158,In_375);
nor U327 (N_327,N_190,N_177);
nor U328 (N_328,N_122,N_105);
xor U329 (N_329,N_239,N_73);
or U330 (N_330,N_235,N_20);
nand U331 (N_331,In_76,N_295);
or U332 (N_332,In_229,N_269);
nand U333 (N_333,N_294,N_229);
or U334 (N_334,In_260,N_263);
or U335 (N_335,N_165,N_62);
nand U336 (N_336,In_387,In_382);
nand U337 (N_337,N_170,N_188);
and U338 (N_338,N_125,N_271);
nand U339 (N_339,N_250,N_133);
or U340 (N_340,N_197,N_232);
and U341 (N_341,In_354,In_144);
and U342 (N_342,In_372,In_234);
nor U343 (N_343,N_257,N_157);
and U344 (N_344,N_174,N_276);
xor U345 (N_345,In_420,N_120);
nor U346 (N_346,N_270,N_242);
or U347 (N_347,In_19,N_172);
nor U348 (N_348,N_226,In_90);
xor U349 (N_349,N_195,In_112);
and U350 (N_350,N_88,N_237);
nand U351 (N_351,In_377,N_236);
or U352 (N_352,In_174,N_76);
and U353 (N_353,N_299,N_245);
and U354 (N_354,In_324,N_278);
nor U355 (N_355,N_260,In_248);
and U356 (N_356,In_386,N_283);
nand U357 (N_357,N_108,In_238);
nor U358 (N_358,In_202,N_218);
nand U359 (N_359,N_134,N_296);
nor U360 (N_360,In_434,N_274);
nor U361 (N_361,In_277,In_465);
or U362 (N_362,N_227,N_152);
or U363 (N_363,N_87,In_81);
xor U364 (N_364,In_240,N_212);
nor U365 (N_365,N_241,N_167);
or U366 (N_366,N_109,N_162);
nor U367 (N_367,N_298,N_79);
nor U368 (N_368,N_154,N_160);
or U369 (N_369,N_173,N_234);
and U370 (N_370,N_265,In_149);
nand U371 (N_371,N_185,N_273);
nand U372 (N_372,In_418,N_124);
nor U373 (N_373,In_472,In_475);
nor U374 (N_374,In_233,N_255);
nand U375 (N_375,N_353,N_341);
and U376 (N_376,N_307,N_335);
nand U377 (N_377,N_309,In_291);
or U378 (N_378,N_210,N_287);
and U379 (N_379,In_59,N_301);
nand U380 (N_380,N_94,N_370);
or U381 (N_381,N_312,N_334);
nor U382 (N_382,N_286,N_281);
or U383 (N_383,N_333,N_347);
nand U384 (N_384,N_360,N_240);
or U385 (N_385,N_372,N_361);
nor U386 (N_386,N_304,N_339);
nand U387 (N_387,N_308,N_355);
or U388 (N_388,N_323,In_369);
nor U389 (N_389,N_349,N_332);
or U390 (N_390,N_244,N_337);
or U391 (N_391,N_31,N_302);
or U392 (N_392,N_292,N_317);
nor U393 (N_393,N_305,N_311);
nor U394 (N_394,N_314,N_356);
and U395 (N_395,N_285,N_364);
nor U396 (N_396,N_121,In_223);
and U397 (N_397,N_225,In_454);
and U398 (N_398,N_315,N_7);
or U399 (N_399,N_316,N_325);
and U400 (N_400,N_217,N_330);
nand U401 (N_401,N_228,In_493);
xnor U402 (N_402,N_9,N_357);
or U403 (N_403,N_324,N_254);
nand U404 (N_404,N_352,N_246);
or U405 (N_405,N_367,In_428);
and U406 (N_406,N_222,N_175);
nand U407 (N_407,N_233,N_213);
nor U408 (N_408,In_430,N_362);
and U409 (N_409,N_248,N_33);
and U410 (N_410,N_338,N_13);
nand U411 (N_411,N_169,In_347);
or U412 (N_412,N_318,N_346);
nor U413 (N_413,N_26,N_303);
or U414 (N_414,N_272,N_328);
nand U415 (N_415,N_331,N_340);
and U416 (N_416,N_365,N_369);
nand U417 (N_417,N_343,N_336);
or U418 (N_418,N_322,In_474);
and U419 (N_419,N_348,N_319);
and U420 (N_420,N_251,N_368);
or U421 (N_421,N_350,N_342);
and U422 (N_422,N_290,N_351);
nor U423 (N_423,N_111,N_320);
nor U424 (N_424,N_374,N_204);
nor U425 (N_425,N_282,N_363);
nand U426 (N_426,N_354,N_358);
and U427 (N_427,N_256,N_313);
nand U428 (N_428,N_289,N_300);
or U429 (N_429,N_373,N_345);
nand U430 (N_430,N_371,N_92);
nor U431 (N_431,N_310,In_16);
or U432 (N_432,N_321,N_326);
nor U433 (N_433,N_243,N_344);
nand U434 (N_434,N_306,N_327);
nor U435 (N_435,N_329,N_359);
nor U436 (N_436,N_115,N_366);
or U437 (N_437,N_252,N_370);
nor U438 (N_438,N_290,N_240);
and U439 (N_439,N_310,N_369);
or U440 (N_440,N_329,N_305);
nand U441 (N_441,N_121,N_213);
or U442 (N_442,N_345,In_347);
nor U443 (N_443,N_204,N_314);
and U444 (N_444,In_430,In_493);
nand U445 (N_445,N_330,N_319);
and U446 (N_446,N_315,N_313);
nand U447 (N_447,N_233,N_370);
or U448 (N_448,N_358,In_369);
and U449 (N_449,N_358,N_334);
xor U450 (N_450,N_412,N_438);
nor U451 (N_451,N_400,N_388);
nand U452 (N_452,N_445,N_380);
and U453 (N_453,N_396,N_430);
nor U454 (N_454,N_383,N_416);
or U455 (N_455,N_397,N_446);
nand U456 (N_456,N_387,N_434);
nand U457 (N_457,N_391,N_385);
or U458 (N_458,N_377,N_414);
nor U459 (N_459,N_398,N_449);
nor U460 (N_460,N_403,N_427);
nor U461 (N_461,N_384,N_417);
nand U462 (N_462,N_435,N_401);
and U463 (N_463,N_404,N_386);
nor U464 (N_464,N_443,N_410);
nor U465 (N_465,N_395,N_418);
and U466 (N_466,N_407,N_411);
nor U467 (N_467,N_389,N_433);
or U468 (N_468,N_413,N_440);
and U469 (N_469,N_381,N_425);
or U470 (N_470,N_415,N_393);
or U471 (N_471,N_390,N_422);
nor U472 (N_472,N_376,N_432);
nand U473 (N_473,N_406,N_409);
and U474 (N_474,N_408,N_424);
nand U475 (N_475,N_419,N_436);
nor U476 (N_476,N_448,N_378);
and U477 (N_477,N_439,N_405);
and U478 (N_478,N_447,N_399);
nand U479 (N_479,N_402,N_444);
or U480 (N_480,N_420,N_426);
and U481 (N_481,N_429,N_431);
or U482 (N_482,N_421,N_382);
nand U483 (N_483,N_423,N_441);
nor U484 (N_484,N_428,N_442);
nand U485 (N_485,N_379,N_375);
nand U486 (N_486,N_394,N_392);
nand U487 (N_487,N_437,N_436);
nand U488 (N_488,N_376,N_436);
or U489 (N_489,N_402,N_394);
nor U490 (N_490,N_396,N_421);
nand U491 (N_491,N_380,N_426);
nor U492 (N_492,N_449,N_414);
or U493 (N_493,N_427,N_413);
nor U494 (N_494,N_440,N_433);
or U495 (N_495,N_375,N_382);
nand U496 (N_496,N_390,N_414);
nand U497 (N_497,N_402,N_379);
or U498 (N_498,N_430,N_433);
and U499 (N_499,N_385,N_419);
and U500 (N_500,N_379,N_449);
nor U501 (N_501,N_423,N_445);
or U502 (N_502,N_397,N_398);
nand U503 (N_503,N_416,N_440);
and U504 (N_504,N_404,N_435);
nand U505 (N_505,N_395,N_415);
or U506 (N_506,N_396,N_380);
or U507 (N_507,N_391,N_383);
nand U508 (N_508,N_396,N_443);
or U509 (N_509,N_443,N_439);
nor U510 (N_510,N_423,N_394);
or U511 (N_511,N_437,N_394);
nand U512 (N_512,N_437,N_418);
or U513 (N_513,N_422,N_425);
nand U514 (N_514,N_425,N_420);
nor U515 (N_515,N_390,N_441);
xor U516 (N_516,N_431,N_408);
or U517 (N_517,N_410,N_440);
nand U518 (N_518,N_406,N_426);
nand U519 (N_519,N_405,N_417);
or U520 (N_520,N_399,N_386);
nor U521 (N_521,N_392,N_437);
or U522 (N_522,N_392,N_382);
xnor U523 (N_523,N_436,N_406);
nor U524 (N_524,N_417,N_387);
and U525 (N_525,N_513,N_491);
nor U526 (N_526,N_475,N_518);
and U527 (N_527,N_472,N_521);
nor U528 (N_528,N_457,N_495);
nor U529 (N_529,N_512,N_450);
or U530 (N_530,N_468,N_464);
nand U531 (N_531,N_501,N_458);
xor U532 (N_532,N_510,N_520);
and U533 (N_533,N_470,N_524);
nand U534 (N_534,N_484,N_481);
and U535 (N_535,N_455,N_471);
nor U536 (N_536,N_483,N_489);
or U537 (N_537,N_463,N_469);
or U538 (N_538,N_508,N_485);
and U539 (N_539,N_493,N_462);
or U540 (N_540,N_522,N_503);
nand U541 (N_541,N_500,N_502);
or U542 (N_542,N_473,N_476);
and U543 (N_543,N_461,N_466);
or U544 (N_544,N_514,N_515);
nand U545 (N_545,N_519,N_453);
and U546 (N_546,N_516,N_465);
and U547 (N_547,N_479,N_486);
and U548 (N_548,N_456,N_490);
nand U549 (N_549,N_523,N_459);
and U550 (N_550,N_487,N_451);
or U551 (N_551,N_454,N_507);
nand U552 (N_552,N_478,N_460);
nor U553 (N_553,N_511,N_494);
nand U554 (N_554,N_499,N_488);
nand U555 (N_555,N_509,N_480);
or U556 (N_556,N_505,N_467);
and U557 (N_557,N_492,N_496);
or U558 (N_558,N_452,N_498);
nor U559 (N_559,N_482,N_474);
nand U560 (N_560,N_477,N_517);
and U561 (N_561,N_504,N_497);
nor U562 (N_562,N_506,N_450);
nand U563 (N_563,N_493,N_497);
and U564 (N_564,N_483,N_479);
and U565 (N_565,N_465,N_489);
nor U566 (N_566,N_501,N_467);
nand U567 (N_567,N_511,N_499);
nor U568 (N_568,N_463,N_503);
or U569 (N_569,N_463,N_501);
or U570 (N_570,N_460,N_509);
and U571 (N_571,N_512,N_483);
and U572 (N_572,N_493,N_507);
xor U573 (N_573,N_494,N_471);
nand U574 (N_574,N_518,N_469);
and U575 (N_575,N_521,N_515);
or U576 (N_576,N_495,N_458);
nand U577 (N_577,N_506,N_471);
and U578 (N_578,N_496,N_457);
xnor U579 (N_579,N_498,N_491);
and U580 (N_580,N_475,N_473);
nand U581 (N_581,N_467,N_455);
and U582 (N_582,N_503,N_452);
and U583 (N_583,N_454,N_520);
and U584 (N_584,N_472,N_478);
and U585 (N_585,N_472,N_518);
nor U586 (N_586,N_522,N_458);
and U587 (N_587,N_457,N_503);
nor U588 (N_588,N_489,N_488);
nor U589 (N_589,N_464,N_509);
and U590 (N_590,N_494,N_476);
nand U591 (N_591,N_511,N_451);
nor U592 (N_592,N_455,N_484);
or U593 (N_593,N_473,N_451);
and U594 (N_594,N_507,N_522);
nor U595 (N_595,N_455,N_511);
nor U596 (N_596,N_483,N_460);
nor U597 (N_597,N_463,N_497);
and U598 (N_598,N_518,N_522);
or U599 (N_599,N_453,N_494);
or U600 (N_600,N_569,N_595);
nor U601 (N_601,N_561,N_568);
nor U602 (N_602,N_543,N_548);
or U603 (N_603,N_582,N_578);
nand U604 (N_604,N_598,N_587);
and U605 (N_605,N_563,N_533);
and U606 (N_606,N_579,N_546);
nand U607 (N_607,N_529,N_538);
nor U608 (N_608,N_570,N_550);
nor U609 (N_609,N_585,N_581);
xnor U610 (N_610,N_527,N_542);
xor U611 (N_611,N_534,N_531);
and U612 (N_612,N_562,N_584);
nand U613 (N_613,N_592,N_556);
nor U614 (N_614,N_594,N_567);
nor U615 (N_615,N_544,N_557);
or U616 (N_616,N_560,N_573);
or U617 (N_617,N_597,N_580);
nor U618 (N_618,N_565,N_590);
or U619 (N_619,N_547,N_599);
nand U620 (N_620,N_589,N_535);
and U621 (N_621,N_576,N_558);
nor U622 (N_622,N_549,N_575);
or U623 (N_623,N_588,N_572);
nor U624 (N_624,N_539,N_545);
or U625 (N_625,N_526,N_586);
nor U626 (N_626,N_541,N_537);
or U627 (N_627,N_530,N_555);
nor U628 (N_628,N_574,N_591);
nand U629 (N_629,N_566,N_551);
nor U630 (N_630,N_593,N_559);
nand U631 (N_631,N_525,N_564);
or U632 (N_632,N_532,N_583);
nand U633 (N_633,N_554,N_596);
and U634 (N_634,N_528,N_552);
nor U635 (N_635,N_536,N_577);
and U636 (N_636,N_571,N_553);
nor U637 (N_637,N_540,N_526);
nand U638 (N_638,N_588,N_546);
or U639 (N_639,N_525,N_581);
or U640 (N_640,N_599,N_572);
and U641 (N_641,N_555,N_570);
or U642 (N_642,N_526,N_547);
and U643 (N_643,N_578,N_525);
xnor U644 (N_644,N_578,N_595);
nor U645 (N_645,N_557,N_548);
or U646 (N_646,N_596,N_581);
and U647 (N_647,N_542,N_540);
nor U648 (N_648,N_585,N_565);
nand U649 (N_649,N_550,N_589);
nand U650 (N_650,N_588,N_530);
nand U651 (N_651,N_560,N_531);
nor U652 (N_652,N_537,N_566);
or U653 (N_653,N_537,N_526);
or U654 (N_654,N_542,N_574);
xor U655 (N_655,N_581,N_563);
or U656 (N_656,N_568,N_536);
or U657 (N_657,N_591,N_599);
nand U658 (N_658,N_574,N_593);
and U659 (N_659,N_571,N_550);
nor U660 (N_660,N_589,N_536);
and U661 (N_661,N_562,N_594);
or U662 (N_662,N_589,N_575);
nor U663 (N_663,N_562,N_557);
or U664 (N_664,N_576,N_557);
nand U665 (N_665,N_589,N_541);
and U666 (N_666,N_594,N_568);
and U667 (N_667,N_597,N_546);
nor U668 (N_668,N_575,N_538);
nand U669 (N_669,N_585,N_538);
nand U670 (N_670,N_550,N_566);
nor U671 (N_671,N_562,N_529);
nand U672 (N_672,N_525,N_554);
or U673 (N_673,N_572,N_526);
nand U674 (N_674,N_571,N_547);
nor U675 (N_675,N_611,N_605);
and U676 (N_676,N_622,N_641);
nor U677 (N_677,N_646,N_644);
and U678 (N_678,N_639,N_658);
and U679 (N_679,N_632,N_607);
nor U680 (N_680,N_652,N_637);
nand U681 (N_681,N_660,N_617);
nor U682 (N_682,N_618,N_620);
nand U683 (N_683,N_661,N_645);
nor U684 (N_684,N_649,N_648);
and U685 (N_685,N_643,N_606);
and U686 (N_686,N_621,N_608);
nand U687 (N_687,N_631,N_610);
or U688 (N_688,N_633,N_613);
or U689 (N_689,N_600,N_668);
and U690 (N_690,N_651,N_656);
or U691 (N_691,N_669,N_657);
or U692 (N_692,N_638,N_604);
and U693 (N_693,N_653,N_629);
nor U694 (N_694,N_619,N_665);
or U695 (N_695,N_674,N_628);
or U696 (N_696,N_626,N_635);
or U697 (N_697,N_663,N_601);
nand U698 (N_698,N_666,N_655);
nor U699 (N_699,N_624,N_615);
or U700 (N_700,N_642,N_636);
nand U701 (N_701,N_603,N_640);
or U702 (N_702,N_673,N_614);
nor U703 (N_703,N_664,N_654);
or U704 (N_704,N_672,N_667);
nor U705 (N_705,N_623,N_612);
nor U706 (N_706,N_650,N_616);
nor U707 (N_707,N_659,N_625);
nand U708 (N_708,N_662,N_671);
nor U709 (N_709,N_609,N_630);
and U710 (N_710,N_627,N_670);
nor U711 (N_711,N_634,N_647);
nand U712 (N_712,N_602,N_615);
nor U713 (N_713,N_636,N_667);
nand U714 (N_714,N_611,N_616);
nand U715 (N_715,N_651,N_629);
or U716 (N_716,N_631,N_644);
nor U717 (N_717,N_672,N_616);
or U718 (N_718,N_606,N_625);
and U719 (N_719,N_643,N_629);
nor U720 (N_720,N_665,N_611);
nor U721 (N_721,N_672,N_646);
nand U722 (N_722,N_609,N_672);
nor U723 (N_723,N_658,N_640);
xnor U724 (N_724,N_672,N_612);
and U725 (N_725,N_644,N_668);
nor U726 (N_726,N_620,N_630);
nor U727 (N_727,N_672,N_674);
nand U728 (N_728,N_610,N_647);
or U729 (N_729,N_621,N_629);
and U730 (N_730,N_655,N_641);
nand U731 (N_731,N_618,N_645);
and U732 (N_732,N_605,N_661);
or U733 (N_733,N_627,N_616);
and U734 (N_734,N_605,N_609);
nor U735 (N_735,N_642,N_644);
nand U736 (N_736,N_606,N_667);
nor U737 (N_737,N_649,N_625);
nor U738 (N_738,N_626,N_605);
nand U739 (N_739,N_613,N_601);
nor U740 (N_740,N_644,N_602);
and U741 (N_741,N_609,N_652);
nand U742 (N_742,N_634,N_654);
and U743 (N_743,N_607,N_641);
nor U744 (N_744,N_633,N_615);
nor U745 (N_745,N_605,N_624);
or U746 (N_746,N_608,N_652);
nor U747 (N_747,N_628,N_616);
nor U748 (N_748,N_663,N_649);
nor U749 (N_749,N_620,N_604);
and U750 (N_750,N_699,N_727);
or U751 (N_751,N_748,N_726);
nor U752 (N_752,N_728,N_679);
nand U753 (N_753,N_698,N_685);
nand U754 (N_754,N_683,N_720);
nand U755 (N_755,N_745,N_737);
nor U756 (N_756,N_702,N_693);
or U757 (N_757,N_690,N_684);
nand U758 (N_758,N_716,N_749);
or U759 (N_759,N_678,N_707);
nand U760 (N_760,N_715,N_709);
nor U761 (N_761,N_740,N_736);
nand U762 (N_762,N_700,N_746);
nand U763 (N_763,N_724,N_688);
nor U764 (N_764,N_689,N_739);
nand U765 (N_765,N_695,N_729);
or U766 (N_766,N_676,N_718);
nand U767 (N_767,N_744,N_742);
nand U768 (N_768,N_686,N_704);
nor U769 (N_769,N_697,N_701);
xor U770 (N_770,N_721,N_692);
nor U771 (N_771,N_733,N_741);
nor U772 (N_772,N_732,N_722);
or U773 (N_773,N_734,N_711);
nor U774 (N_774,N_691,N_710);
xnor U775 (N_775,N_705,N_696);
and U776 (N_776,N_680,N_694);
nor U777 (N_777,N_706,N_687);
or U778 (N_778,N_713,N_730);
nand U779 (N_779,N_747,N_708);
nand U780 (N_780,N_731,N_743);
nand U781 (N_781,N_717,N_714);
nand U782 (N_782,N_681,N_738);
nor U783 (N_783,N_723,N_719);
and U784 (N_784,N_703,N_682);
or U785 (N_785,N_675,N_677);
nand U786 (N_786,N_725,N_735);
nor U787 (N_787,N_712,N_705);
nand U788 (N_788,N_703,N_737);
nand U789 (N_789,N_720,N_706);
or U790 (N_790,N_728,N_733);
and U791 (N_791,N_737,N_741);
or U792 (N_792,N_694,N_717);
nand U793 (N_793,N_677,N_692);
nand U794 (N_794,N_707,N_718);
and U795 (N_795,N_744,N_731);
nand U796 (N_796,N_690,N_743);
nor U797 (N_797,N_731,N_723);
nor U798 (N_798,N_703,N_711);
nor U799 (N_799,N_744,N_708);
or U800 (N_800,N_690,N_739);
or U801 (N_801,N_716,N_734);
and U802 (N_802,N_676,N_732);
or U803 (N_803,N_734,N_681);
and U804 (N_804,N_714,N_681);
nor U805 (N_805,N_732,N_718);
nand U806 (N_806,N_726,N_725);
nor U807 (N_807,N_710,N_746);
nor U808 (N_808,N_701,N_749);
and U809 (N_809,N_705,N_719);
and U810 (N_810,N_732,N_720);
and U811 (N_811,N_708,N_690);
or U812 (N_812,N_719,N_704);
nand U813 (N_813,N_703,N_720);
and U814 (N_814,N_721,N_741);
nand U815 (N_815,N_697,N_684);
nor U816 (N_816,N_705,N_706);
and U817 (N_817,N_683,N_675);
and U818 (N_818,N_735,N_731);
and U819 (N_819,N_691,N_738);
and U820 (N_820,N_696,N_734);
or U821 (N_821,N_734,N_686);
nand U822 (N_822,N_689,N_696);
nor U823 (N_823,N_731,N_675);
nand U824 (N_824,N_729,N_720);
and U825 (N_825,N_785,N_799);
nand U826 (N_826,N_761,N_765);
or U827 (N_827,N_812,N_791);
nand U828 (N_828,N_777,N_783);
and U829 (N_829,N_795,N_750);
nand U830 (N_830,N_816,N_753);
and U831 (N_831,N_770,N_803);
nor U832 (N_832,N_817,N_782);
and U833 (N_833,N_787,N_822);
or U834 (N_834,N_772,N_773);
nor U835 (N_835,N_823,N_819);
or U836 (N_836,N_781,N_784);
nor U837 (N_837,N_759,N_775);
nor U838 (N_838,N_762,N_810);
nand U839 (N_839,N_807,N_767);
or U840 (N_840,N_756,N_808);
nor U841 (N_841,N_786,N_776);
nor U842 (N_842,N_804,N_755);
and U843 (N_843,N_780,N_815);
nor U844 (N_844,N_818,N_824);
nand U845 (N_845,N_800,N_774);
or U846 (N_846,N_814,N_796);
and U847 (N_847,N_764,N_792);
nor U848 (N_848,N_752,N_758);
nor U849 (N_849,N_754,N_768);
nor U850 (N_850,N_779,N_769);
or U851 (N_851,N_813,N_794);
or U852 (N_852,N_788,N_778);
or U853 (N_853,N_821,N_771);
nor U854 (N_854,N_797,N_789);
and U855 (N_855,N_760,N_811);
or U856 (N_856,N_820,N_801);
and U857 (N_857,N_757,N_763);
nor U858 (N_858,N_793,N_798);
or U859 (N_859,N_806,N_805);
nor U860 (N_860,N_809,N_751);
nor U861 (N_861,N_766,N_802);
or U862 (N_862,N_790,N_816);
and U863 (N_863,N_785,N_808);
and U864 (N_864,N_784,N_785);
and U865 (N_865,N_809,N_767);
nor U866 (N_866,N_799,N_772);
and U867 (N_867,N_818,N_786);
nand U868 (N_868,N_803,N_812);
nand U869 (N_869,N_765,N_776);
nor U870 (N_870,N_771,N_795);
nor U871 (N_871,N_750,N_764);
nor U872 (N_872,N_779,N_763);
and U873 (N_873,N_783,N_813);
and U874 (N_874,N_779,N_804);
and U875 (N_875,N_800,N_759);
nand U876 (N_876,N_757,N_779);
or U877 (N_877,N_756,N_817);
nor U878 (N_878,N_760,N_822);
nor U879 (N_879,N_750,N_776);
nor U880 (N_880,N_758,N_796);
or U881 (N_881,N_798,N_761);
nand U882 (N_882,N_811,N_810);
nor U883 (N_883,N_753,N_776);
nor U884 (N_884,N_803,N_763);
and U885 (N_885,N_774,N_798);
and U886 (N_886,N_788,N_824);
and U887 (N_887,N_752,N_783);
nand U888 (N_888,N_815,N_817);
and U889 (N_889,N_776,N_815);
or U890 (N_890,N_811,N_771);
and U891 (N_891,N_791,N_779);
and U892 (N_892,N_759,N_786);
or U893 (N_893,N_805,N_803);
nor U894 (N_894,N_814,N_806);
or U895 (N_895,N_810,N_803);
nand U896 (N_896,N_788,N_800);
xor U897 (N_897,N_755,N_779);
and U898 (N_898,N_814,N_756);
and U899 (N_899,N_773,N_810);
or U900 (N_900,N_895,N_862);
xor U901 (N_901,N_890,N_886);
and U902 (N_902,N_857,N_850);
nand U903 (N_903,N_896,N_847);
nand U904 (N_904,N_830,N_884);
or U905 (N_905,N_838,N_826);
nand U906 (N_906,N_869,N_832);
nor U907 (N_907,N_825,N_897);
nor U908 (N_908,N_834,N_898);
nand U909 (N_909,N_892,N_833);
or U910 (N_910,N_882,N_881);
nand U911 (N_911,N_863,N_864);
and U912 (N_912,N_854,N_837);
or U913 (N_913,N_880,N_894);
nor U914 (N_914,N_879,N_871);
nor U915 (N_915,N_887,N_843);
nand U916 (N_916,N_885,N_870);
and U917 (N_917,N_899,N_867);
nand U918 (N_918,N_878,N_852);
nor U919 (N_919,N_872,N_855);
nor U920 (N_920,N_859,N_875);
nor U921 (N_921,N_874,N_865);
or U922 (N_922,N_831,N_845);
nand U923 (N_923,N_868,N_893);
nor U924 (N_924,N_848,N_849);
and U925 (N_925,N_853,N_840);
nand U926 (N_926,N_883,N_888);
nor U927 (N_927,N_866,N_829);
and U928 (N_928,N_842,N_877);
nor U929 (N_929,N_827,N_861);
or U930 (N_930,N_839,N_889);
nor U931 (N_931,N_851,N_841);
nor U932 (N_932,N_846,N_835);
nor U933 (N_933,N_873,N_836);
nor U934 (N_934,N_844,N_860);
or U935 (N_935,N_828,N_858);
nor U936 (N_936,N_891,N_876);
nor U937 (N_937,N_856,N_843);
or U938 (N_938,N_829,N_864);
or U939 (N_939,N_866,N_826);
and U940 (N_940,N_840,N_834);
and U941 (N_941,N_847,N_872);
nor U942 (N_942,N_877,N_839);
nor U943 (N_943,N_826,N_825);
or U944 (N_944,N_842,N_884);
and U945 (N_945,N_883,N_847);
nor U946 (N_946,N_831,N_840);
nand U947 (N_947,N_836,N_871);
and U948 (N_948,N_896,N_866);
and U949 (N_949,N_833,N_895);
nand U950 (N_950,N_844,N_850);
and U951 (N_951,N_885,N_834);
nor U952 (N_952,N_871,N_830);
or U953 (N_953,N_862,N_841);
xor U954 (N_954,N_838,N_843);
and U955 (N_955,N_878,N_847);
nor U956 (N_956,N_876,N_873);
or U957 (N_957,N_868,N_864);
or U958 (N_958,N_851,N_848);
nand U959 (N_959,N_834,N_892);
and U960 (N_960,N_871,N_894);
nand U961 (N_961,N_868,N_847);
nor U962 (N_962,N_854,N_882);
nor U963 (N_963,N_862,N_890);
nand U964 (N_964,N_879,N_883);
nand U965 (N_965,N_855,N_895);
and U966 (N_966,N_841,N_889);
nand U967 (N_967,N_835,N_839);
and U968 (N_968,N_856,N_825);
nand U969 (N_969,N_888,N_870);
xor U970 (N_970,N_891,N_879);
and U971 (N_971,N_870,N_829);
nand U972 (N_972,N_858,N_897);
nor U973 (N_973,N_881,N_892);
and U974 (N_974,N_860,N_897);
and U975 (N_975,N_944,N_913);
nand U976 (N_976,N_964,N_966);
or U977 (N_977,N_926,N_946);
nor U978 (N_978,N_922,N_952);
nor U979 (N_979,N_901,N_931);
nand U980 (N_980,N_941,N_961);
or U981 (N_981,N_935,N_930);
or U982 (N_982,N_917,N_920);
nor U983 (N_983,N_965,N_967);
nand U984 (N_984,N_924,N_905);
nor U985 (N_985,N_974,N_951);
or U986 (N_986,N_968,N_919);
nand U987 (N_987,N_923,N_939);
nor U988 (N_988,N_908,N_972);
nor U989 (N_989,N_918,N_929);
or U990 (N_990,N_936,N_949);
nand U991 (N_991,N_963,N_903);
or U992 (N_992,N_938,N_959);
and U993 (N_993,N_927,N_958);
and U994 (N_994,N_945,N_942);
and U995 (N_995,N_969,N_960);
nor U996 (N_996,N_954,N_947);
xnor U997 (N_997,N_955,N_940);
or U998 (N_998,N_911,N_933);
nand U999 (N_999,N_925,N_906);
nand U1000 (N_1000,N_962,N_956);
or U1001 (N_1001,N_900,N_943);
nor U1002 (N_1002,N_950,N_910);
nand U1003 (N_1003,N_912,N_971);
or U1004 (N_1004,N_934,N_914);
nand U1005 (N_1005,N_948,N_937);
nor U1006 (N_1006,N_904,N_932);
nor U1007 (N_1007,N_953,N_957);
nand U1008 (N_1008,N_907,N_916);
or U1009 (N_1009,N_909,N_928);
and U1010 (N_1010,N_921,N_973);
nor U1011 (N_1011,N_970,N_915);
nand U1012 (N_1012,N_902,N_959);
or U1013 (N_1013,N_939,N_924);
and U1014 (N_1014,N_956,N_903);
nand U1015 (N_1015,N_958,N_955);
xnor U1016 (N_1016,N_949,N_905);
and U1017 (N_1017,N_961,N_921);
and U1018 (N_1018,N_954,N_923);
nor U1019 (N_1019,N_901,N_948);
nor U1020 (N_1020,N_943,N_970);
and U1021 (N_1021,N_913,N_926);
and U1022 (N_1022,N_929,N_956);
and U1023 (N_1023,N_903,N_929);
nor U1024 (N_1024,N_974,N_947);
or U1025 (N_1025,N_968,N_936);
nand U1026 (N_1026,N_961,N_936);
nor U1027 (N_1027,N_962,N_915);
and U1028 (N_1028,N_956,N_911);
or U1029 (N_1029,N_968,N_924);
and U1030 (N_1030,N_957,N_903);
and U1031 (N_1031,N_968,N_928);
or U1032 (N_1032,N_937,N_945);
nand U1033 (N_1033,N_927,N_942);
or U1034 (N_1034,N_915,N_910);
nor U1035 (N_1035,N_936,N_971);
nor U1036 (N_1036,N_933,N_938);
nand U1037 (N_1037,N_943,N_951);
nor U1038 (N_1038,N_909,N_903);
and U1039 (N_1039,N_917,N_939);
nand U1040 (N_1040,N_938,N_963);
and U1041 (N_1041,N_955,N_965);
and U1042 (N_1042,N_958,N_940);
and U1043 (N_1043,N_911,N_922);
or U1044 (N_1044,N_942,N_937);
nor U1045 (N_1045,N_906,N_965);
nand U1046 (N_1046,N_966,N_926);
nor U1047 (N_1047,N_945,N_918);
nor U1048 (N_1048,N_904,N_946);
or U1049 (N_1049,N_909,N_945);
nor U1050 (N_1050,N_1012,N_1040);
or U1051 (N_1051,N_987,N_1004);
nor U1052 (N_1052,N_993,N_981);
nor U1053 (N_1053,N_1047,N_995);
or U1054 (N_1054,N_1010,N_982);
nand U1055 (N_1055,N_991,N_1023);
nand U1056 (N_1056,N_1024,N_1046);
nand U1057 (N_1057,N_1019,N_1020);
nor U1058 (N_1058,N_1021,N_976);
or U1059 (N_1059,N_1031,N_1026);
or U1060 (N_1060,N_998,N_1025);
or U1061 (N_1061,N_1014,N_1038);
nor U1062 (N_1062,N_1016,N_980);
and U1063 (N_1063,N_975,N_977);
or U1064 (N_1064,N_989,N_990);
and U1065 (N_1065,N_1030,N_979);
and U1066 (N_1066,N_1036,N_1042);
or U1067 (N_1067,N_1033,N_1035);
nand U1068 (N_1068,N_978,N_996);
xnor U1069 (N_1069,N_1018,N_1006);
xnor U1070 (N_1070,N_1044,N_984);
or U1071 (N_1071,N_1043,N_1002);
nor U1072 (N_1072,N_1022,N_1032);
nor U1073 (N_1073,N_986,N_999);
and U1074 (N_1074,N_1045,N_1048);
and U1075 (N_1075,N_1015,N_1001);
nand U1076 (N_1076,N_1007,N_1034);
nor U1077 (N_1077,N_1028,N_983);
or U1078 (N_1078,N_1011,N_1008);
xor U1079 (N_1079,N_1037,N_1039);
nand U1080 (N_1080,N_1041,N_1005);
or U1081 (N_1081,N_1017,N_1009);
or U1082 (N_1082,N_997,N_1000);
or U1083 (N_1083,N_1049,N_994);
or U1084 (N_1084,N_1027,N_992);
nand U1085 (N_1085,N_985,N_1013);
nor U1086 (N_1086,N_1003,N_1029);
and U1087 (N_1087,N_988,N_1044);
nand U1088 (N_1088,N_1006,N_987);
and U1089 (N_1089,N_1016,N_977);
nor U1090 (N_1090,N_1037,N_1025);
or U1091 (N_1091,N_1005,N_977);
nor U1092 (N_1092,N_975,N_992);
nor U1093 (N_1093,N_1006,N_1003);
nand U1094 (N_1094,N_1020,N_1035);
and U1095 (N_1095,N_1040,N_1018);
nand U1096 (N_1096,N_1026,N_1001);
nor U1097 (N_1097,N_1049,N_1024);
and U1098 (N_1098,N_1019,N_1035);
nor U1099 (N_1099,N_1030,N_1023);
nor U1100 (N_1100,N_1002,N_1041);
and U1101 (N_1101,N_983,N_1030);
nor U1102 (N_1102,N_977,N_1041);
nand U1103 (N_1103,N_1007,N_1030);
nand U1104 (N_1104,N_1038,N_996);
nor U1105 (N_1105,N_1001,N_1039);
nor U1106 (N_1106,N_983,N_1032);
and U1107 (N_1107,N_1035,N_1023);
nand U1108 (N_1108,N_1030,N_1027);
or U1109 (N_1109,N_1002,N_1048);
or U1110 (N_1110,N_1018,N_1020);
nand U1111 (N_1111,N_1004,N_1036);
nor U1112 (N_1112,N_1027,N_1003);
nand U1113 (N_1113,N_1018,N_990);
nor U1114 (N_1114,N_1019,N_1047);
nand U1115 (N_1115,N_986,N_1047);
xnor U1116 (N_1116,N_997,N_993);
nand U1117 (N_1117,N_1011,N_1003);
and U1118 (N_1118,N_1010,N_1021);
or U1119 (N_1119,N_995,N_1021);
nor U1120 (N_1120,N_1026,N_1046);
nor U1121 (N_1121,N_1040,N_977);
xor U1122 (N_1122,N_994,N_1031);
and U1123 (N_1123,N_1004,N_1018);
or U1124 (N_1124,N_975,N_1010);
or U1125 (N_1125,N_1096,N_1060);
and U1126 (N_1126,N_1056,N_1057);
nor U1127 (N_1127,N_1055,N_1065);
or U1128 (N_1128,N_1087,N_1119);
nand U1129 (N_1129,N_1068,N_1117);
or U1130 (N_1130,N_1110,N_1118);
nor U1131 (N_1131,N_1072,N_1050);
nor U1132 (N_1132,N_1075,N_1073);
or U1133 (N_1133,N_1114,N_1107);
nor U1134 (N_1134,N_1090,N_1082);
nor U1135 (N_1135,N_1102,N_1054);
and U1136 (N_1136,N_1121,N_1097);
or U1137 (N_1137,N_1120,N_1078);
or U1138 (N_1138,N_1115,N_1083);
nand U1139 (N_1139,N_1098,N_1099);
nor U1140 (N_1140,N_1081,N_1124);
or U1141 (N_1141,N_1061,N_1052);
nand U1142 (N_1142,N_1109,N_1085);
nand U1143 (N_1143,N_1086,N_1091);
or U1144 (N_1144,N_1064,N_1104);
or U1145 (N_1145,N_1058,N_1108);
nor U1146 (N_1146,N_1100,N_1070);
and U1147 (N_1147,N_1062,N_1051);
or U1148 (N_1148,N_1053,N_1077);
nor U1149 (N_1149,N_1059,N_1094);
xor U1150 (N_1150,N_1103,N_1122);
and U1151 (N_1151,N_1079,N_1093);
nor U1152 (N_1152,N_1123,N_1101);
xor U1153 (N_1153,N_1089,N_1080);
nand U1154 (N_1154,N_1088,N_1074);
nand U1155 (N_1155,N_1116,N_1105);
nor U1156 (N_1156,N_1112,N_1106);
or U1157 (N_1157,N_1113,N_1066);
or U1158 (N_1158,N_1069,N_1076);
nor U1159 (N_1159,N_1092,N_1095);
and U1160 (N_1160,N_1111,N_1084);
nor U1161 (N_1161,N_1067,N_1063);
nand U1162 (N_1162,N_1071,N_1110);
nand U1163 (N_1163,N_1067,N_1111);
or U1164 (N_1164,N_1114,N_1062);
nand U1165 (N_1165,N_1061,N_1091);
nor U1166 (N_1166,N_1069,N_1056);
nor U1167 (N_1167,N_1088,N_1109);
nor U1168 (N_1168,N_1102,N_1124);
and U1169 (N_1169,N_1070,N_1120);
or U1170 (N_1170,N_1109,N_1099);
nand U1171 (N_1171,N_1104,N_1107);
or U1172 (N_1172,N_1116,N_1118);
or U1173 (N_1173,N_1089,N_1083);
or U1174 (N_1174,N_1109,N_1100);
and U1175 (N_1175,N_1051,N_1116);
and U1176 (N_1176,N_1088,N_1087);
nor U1177 (N_1177,N_1101,N_1066);
and U1178 (N_1178,N_1084,N_1069);
or U1179 (N_1179,N_1094,N_1082);
nor U1180 (N_1180,N_1050,N_1103);
and U1181 (N_1181,N_1122,N_1076);
nor U1182 (N_1182,N_1089,N_1070);
or U1183 (N_1183,N_1064,N_1070);
and U1184 (N_1184,N_1058,N_1098);
nor U1185 (N_1185,N_1124,N_1111);
and U1186 (N_1186,N_1052,N_1109);
nand U1187 (N_1187,N_1065,N_1087);
nand U1188 (N_1188,N_1119,N_1072);
and U1189 (N_1189,N_1119,N_1106);
nand U1190 (N_1190,N_1119,N_1050);
nand U1191 (N_1191,N_1072,N_1116);
nand U1192 (N_1192,N_1052,N_1076);
nor U1193 (N_1193,N_1101,N_1107);
and U1194 (N_1194,N_1111,N_1079);
nand U1195 (N_1195,N_1051,N_1112);
nand U1196 (N_1196,N_1097,N_1051);
nor U1197 (N_1197,N_1116,N_1065);
and U1198 (N_1198,N_1071,N_1086);
and U1199 (N_1199,N_1076,N_1119);
nor U1200 (N_1200,N_1143,N_1141);
nand U1201 (N_1201,N_1137,N_1128);
nor U1202 (N_1202,N_1135,N_1176);
nor U1203 (N_1203,N_1142,N_1184);
and U1204 (N_1204,N_1185,N_1190);
nor U1205 (N_1205,N_1181,N_1127);
or U1206 (N_1206,N_1178,N_1154);
nor U1207 (N_1207,N_1188,N_1150);
or U1208 (N_1208,N_1187,N_1167);
nor U1209 (N_1209,N_1172,N_1194);
nor U1210 (N_1210,N_1131,N_1168);
or U1211 (N_1211,N_1169,N_1139);
or U1212 (N_1212,N_1155,N_1191);
nand U1213 (N_1213,N_1159,N_1189);
and U1214 (N_1214,N_1152,N_1138);
and U1215 (N_1215,N_1149,N_1173);
nor U1216 (N_1216,N_1158,N_1179);
or U1217 (N_1217,N_1145,N_1199);
nor U1218 (N_1218,N_1193,N_1146);
nor U1219 (N_1219,N_1133,N_1136);
or U1220 (N_1220,N_1197,N_1162);
nor U1221 (N_1221,N_1177,N_1175);
and U1222 (N_1222,N_1151,N_1171);
and U1223 (N_1223,N_1153,N_1164);
nand U1224 (N_1224,N_1130,N_1170);
nor U1225 (N_1225,N_1125,N_1163);
or U1226 (N_1226,N_1166,N_1134);
nand U1227 (N_1227,N_1160,N_1148);
and U1228 (N_1228,N_1180,N_1129);
xor U1229 (N_1229,N_1165,N_1126);
nor U1230 (N_1230,N_1140,N_1198);
nor U1231 (N_1231,N_1186,N_1157);
and U1232 (N_1232,N_1196,N_1147);
or U1233 (N_1233,N_1144,N_1161);
and U1234 (N_1234,N_1183,N_1174);
and U1235 (N_1235,N_1195,N_1192);
nor U1236 (N_1236,N_1156,N_1182);
xnor U1237 (N_1237,N_1132,N_1153);
nor U1238 (N_1238,N_1179,N_1162);
nor U1239 (N_1239,N_1150,N_1184);
and U1240 (N_1240,N_1198,N_1155);
xnor U1241 (N_1241,N_1168,N_1135);
nor U1242 (N_1242,N_1157,N_1159);
and U1243 (N_1243,N_1125,N_1134);
or U1244 (N_1244,N_1171,N_1176);
nand U1245 (N_1245,N_1128,N_1179);
and U1246 (N_1246,N_1170,N_1169);
and U1247 (N_1247,N_1199,N_1171);
nand U1248 (N_1248,N_1182,N_1129);
nand U1249 (N_1249,N_1144,N_1168);
or U1250 (N_1250,N_1149,N_1192);
and U1251 (N_1251,N_1182,N_1186);
and U1252 (N_1252,N_1182,N_1171);
nor U1253 (N_1253,N_1197,N_1184);
nor U1254 (N_1254,N_1143,N_1172);
and U1255 (N_1255,N_1183,N_1152);
nor U1256 (N_1256,N_1193,N_1148);
nor U1257 (N_1257,N_1142,N_1190);
nand U1258 (N_1258,N_1129,N_1161);
nand U1259 (N_1259,N_1172,N_1179);
or U1260 (N_1260,N_1161,N_1127);
and U1261 (N_1261,N_1171,N_1166);
nor U1262 (N_1262,N_1191,N_1172);
nor U1263 (N_1263,N_1144,N_1166);
nor U1264 (N_1264,N_1170,N_1199);
nor U1265 (N_1265,N_1148,N_1186);
nor U1266 (N_1266,N_1178,N_1180);
nor U1267 (N_1267,N_1150,N_1171);
or U1268 (N_1268,N_1132,N_1161);
nor U1269 (N_1269,N_1151,N_1190);
and U1270 (N_1270,N_1159,N_1155);
or U1271 (N_1271,N_1147,N_1185);
nor U1272 (N_1272,N_1156,N_1150);
and U1273 (N_1273,N_1142,N_1139);
or U1274 (N_1274,N_1189,N_1157);
or U1275 (N_1275,N_1258,N_1256);
and U1276 (N_1276,N_1210,N_1266);
nand U1277 (N_1277,N_1216,N_1233);
nand U1278 (N_1278,N_1209,N_1203);
nand U1279 (N_1279,N_1260,N_1219);
xor U1280 (N_1280,N_1265,N_1224);
nor U1281 (N_1281,N_1230,N_1274);
or U1282 (N_1282,N_1226,N_1238);
nor U1283 (N_1283,N_1268,N_1247);
and U1284 (N_1284,N_1225,N_1255);
nor U1285 (N_1285,N_1237,N_1259);
and U1286 (N_1286,N_1261,N_1232);
and U1287 (N_1287,N_1202,N_1215);
or U1288 (N_1288,N_1234,N_1221);
or U1289 (N_1289,N_1217,N_1227);
nand U1290 (N_1290,N_1240,N_1248);
and U1291 (N_1291,N_1207,N_1264);
nand U1292 (N_1292,N_1231,N_1213);
or U1293 (N_1293,N_1241,N_1249);
or U1294 (N_1294,N_1271,N_1242);
xnor U1295 (N_1295,N_1252,N_1223);
nor U1296 (N_1296,N_1244,N_1204);
nor U1297 (N_1297,N_1269,N_1262);
nor U1298 (N_1298,N_1250,N_1245);
and U1299 (N_1299,N_1243,N_1257);
nand U1300 (N_1300,N_1206,N_1251);
nor U1301 (N_1301,N_1246,N_1201);
nand U1302 (N_1302,N_1200,N_1211);
and U1303 (N_1303,N_1235,N_1208);
nand U1304 (N_1304,N_1228,N_1220);
nor U1305 (N_1305,N_1218,N_1212);
xor U1306 (N_1306,N_1254,N_1205);
xnor U1307 (N_1307,N_1272,N_1267);
nor U1308 (N_1308,N_1239,N_1273);
nor U1309 (N_1309,N_1229,N_1236);
xor U1310 (N_1310,N_1270,N_1222);
nor U1311 (N_1311,N_1253,N_1214);
xnor U1312 (N_1312,N_1263,N_1236);
nand U1313 (N_1313,N_1207,N_1248);
and U1314 (N_1314,N_1212,N_1241);
nor U1315 (N_1315,N_1202,N_1241);
and U1316 (N_1316,N_1204,N_1271);
and U1317 (N_1317,N_1249,N_1274);
and U1318 (N_1318,N_1220,N_1202);
nor U1319 (N_1319,N_1245,N_1267);
and U1320 (N_1320,N_1212,N_1253);
or U1321 (N_1321,N_1247,N_1200);
nor U1322 (N_1322,N_1251,N_1218);
and U1323 (N_1323,N_1200,N_1259);
and U1324 (N_1324,N_1265,N_1227);
and U1325 (N_1325,N_1270,N_1252);
and U1326 (N_1326,N_1257,N_1206);
and U1327 (N_1327,N_1259,N_1273);
or U1328 (N_1328,N_1248,N_1243);
nor U1329 (N_1329,N_1202,N_1255);
nand U1330 (N_1330,N_1265,N_1270);
nor U1331 (N_1331,N_1232,N_1269);
or U1332 (N_1332,N_1274,N_1273);
nand U1333 (N_1333,N_1247,N_1263);
or U1334 (N_1334,N_1205,N_1255);
or U1335 (N_1335,N_1248,N_1266);
or U1336 (N_1336,N_1239,N_1240);
nor U1337 (N_1337,N_1206,N_1250);
and U1338 (N_1338,N_1273,N_1217);
and U1339 (N_1339,N_1249,N_1273);
and U1340 (N_1340,N_1204,N_1221);
or U1341 (N_1341,N_1208,N_1262);
nand U1342 (N_1342,N_1263,N_1246);
nand U1343 (N_1343,N_1219,N_1202);
nor U1344 (N_1344,N_1227,N_1262);
and U1345 (N_1345,N_1246,N_1251);
nand U1346 (N_1346,N_1207,N_1221);
nor U1347 (N_1347,N_1209,N_1249);
nor U1348 (N_1348,N_1253,N_1257);
or U1349 (N_1349,N_1239,N_1243);
nor U1350 (N_1350,N_1316,N_1331);
or U1351 (N_1351,N_1317,N_1297);
and U1352 (N_1352,N_1280,N_1285);
nor U1353 (N_1353,N_1307,N_1311);
nand U1354 (N_1354,N_1278,N_1279);
nor U1355 (N_1355,N_1320,N_1332);
nor U1356 (N_1356,N_1283,N_1294);
or U1357 (N_1357,N_1341,N_1328);
nand U1358 (N_1358,N_1309,N_1275);
and U1359 (N_1359,N_1304,N_1288);
or U1360 (N_1360,N_1345,N_1286);
and U1361 (N_1361,N_1338,N_1292);
nor U1362 (N_1362,N_1287,N_1324);
nor U1363 (N_1363,N_1302,N_1339);
or U1364 (N_1364,N_1323,N_1310);
and U1365 (N_1365,N_1299,N_1333);
xnor U1366 (N_1366,N_1290,N_1291);
and U1367 (N_1367,N_1346,N_1347);
nand U1368 (N_1368,N_1296,N_1276);
nand U1369 (N_1369,N_1301,N_1334);
or U1370 (N_1370,N_1293,N_1330);
and U1371 (N_1371,N_1313,N_1336);
nand U1372 (N_1372,N_1342,N_1348);
nor U1373 (N_1373,N_1343,N_1306);
and U1374 (N_1374,N_1337,N_1295);
nor U1375 (N_1375,N_1308,N_1315);
nor U1376 (N_1376,N_1335,N_1300);
and U1377 (N_1377,N_1318,N_1327);
nor U1378 (N_1378,N_1349,N_1314);
and U1379 (N_1379,N_1281,N_1298);
or U1380 (N_1380,N_1289,N_1284);
nand U1381 (N_1381,N_1282,N_1322);
xor U1382 (N_1382,N_1303,N_1344);
or U1383 (N_1383,N_1340,N_1312);
nand U1384 (N_1384,N_1321,N_1305);
nor U1385 (N_1385,N_1277,N_1326);
nand U1386 (N_1386,N_1319,N_1329);
nor U1387 (N_1387,N_1325,N_1313);
or U1388 (N_1388,N_1335,N_1316);
or U1389 (N_1389,N_1292,N_1334);
nor U1390 (N_1390,N_1292,N_1308);
nand U1391 (N_1391,N_1319,N_1282);
or U1392 (N_1392,N_1304,N_1330);
nand U1393 (N_1393,N_1297,N_1347);
or U1394 (N_1394,N_1332,N_1314);
or U1395 (N_1395,N_1320,N_1345);
nand U1396 (N_1396,N_1304,N_1338);
and U1397 (N_1397,N_1292,N_1295);
xor U1398 (N_1398,N_1288,N_1277);
and U1399 (N_1399,N_1322,N_1302);
or U1400 (N_1400,N_1333,N_1297);
nor U1401 (N_1401,N_1320,N_1276);
nor U1402 (N_1402,N_1347,N_1277);
xor U1403 (N_1403,N_1348,N_1328);
and U1404 (N_1404,N_1345,N_1277);
nor U1405 (N_1405,N_1283,N_1275);
or U1406 (N_1406,N_1288,N_1287);
nor U1407 (N_1407,N_1324,N_1280);
or U1408 (N_1408,N_1341,N_1312);
or U1409 (N_1409,N_1287,N_1286);
nand U1410 (N_1410,N_1295,N_1304);
nor U1411 (N_1411,N_1325,N_1279);
nor U1412 (N_1412,N_1300,N_1306);
or U1413 (N_1413,N_1329,N_1332);
and U1414 (N_1414,N_1310,N_1299);
or U1415 (N_1415,N_1276,N_1279);
and U1416 (N_1416,N_1284,N_1277);
nor U1417 (N_1417,N_1301,N_1277);
or U1418 (N_1418,N_1336,N_1346);
nand U1419 (N_1419,N_1288,N_1326);
nor U1420 (N_1420,N_1303,N_1292);
or U1421 (N_1421,N_1278,N_1334);
nand U1422 (N_1422,N_1286,N_1326);
or U1423 (N_1423,N_1304,N_1325);
nor U1424 (N_1424,N_1275,N_1343);
xor U1425 (N_1425,N_1418,N_1424);
or U1426 (N_1426,N_1398,N_1382);
nand U1427 (N_1427,N_1369,N_1413);
or U1428 (N_1428,N_1386,N_1399);
and U1429 (N_1429,N_1391,N_1360);
or U1430 (N_1430,N_1420,N_1367);
and U1431 (N_1431,N_1394,N_1415);
nand U1432 (N_1432,N_1392,N_1387);
nand U1433 (N_1433,N_1361,N_1354);
nor U1434 (N_1434,N_1384,N_1381);
nand U1435 (N_1435,N_1390,N_1419);
nand U1436 (N_1436,N_1396,N_1417);
nor U1437 (N_1437,N_1356,N_1383);
nor U1438 (N_1438,N_1421,N_1378);
and U1439 (N_1439,N_1351,N_1423);
nor U1440 (N_1440,N_1397,N_1357);
xnor U1441 (N_1441,N_1379,N_1364);
and U1442 (N_1442,N_1389,N_1414);
and U1443 (N_1443,N_1403,N_1411);
nor U1444 (N_1444,N_1393,N_1366);
nand U1445 (N_1445,N_1373,N_1358);
or U1446 (N_1446,N_1375,N_1365);
nor U1447 (N_1447,N_1409,N_1402);
nor U1448 (N_1448,N_1395,N_1376);
or U1449 (N_1449,N_1401,N_1353);
or U1450 (N_1450,N_1355,N_1412);
and U1451 (N_1451,N_1374,N_1422);
nand U1452 (N_1452,N_1368,N_1388);
and U1453 (N_1453,N_1406,N_1416);
and U1454 (N_1454,N_1352,N_1380);
nor U1455 (N_1455,N_1410,N_1377);
and U1456 (N_1456,N_1363,N_1362);
nand U1457 (N_1457,N_1370,N_1407);
and U1458 (N_1458,N_1372,N_1359);
nor U1459 (N_1459,N_1408,N_1371);
and U1460 (N_1460,N_1404,N_1405);
nor U1461 (N_1461,N_1400,N_1385);
nor U1462 (N_1462,N_1350,N_1390);
or U1463 (N_1463,N_1422,N_1350);
and U1464 (N_1464,N_1409,N_1405);
or U1465 (N_1465,N_1418,N_1355);
nand U1466 (N_1466,N_1421,N_1367);
or U1467 (N_1467,N_1351,N_1357);
nor U1468 (N_1468,N_1366,N_1409);
and U1469 (N_1469,N_1417,N_1378);
nor U1470 (N_1470,N_1385,N_1388);
nor U1471 (N_1471,N_1359,N_1351);
and U1472 (N_1472,N_1368,N_1384);
nand U1473 (N_1473,N_1352,N_1408);
nor U1474 (N_1474,N_1387,N_1395);
or U1475 (N_1475,N_1377,N_1380);
nand U1476 (N_1476,N_1417,N_1367);
and U1477 (N_1477,N_1373,N_1385);
or U1478 (N_1478,N_1378,N_1380);
nand U1479 (N_1479,N_1367,N_1406);
or U1480 (N_1480,N_1364,N_1371);
and U1481 (N_1481,N_1411,N_1368);
and U1482 (N_1482,N_1417,N_1368);
nor U1483 (N_1483,N_1377,N_1373);
nand U1484 (N_1484,N_1368,N_1383);
nand U1485 (N_1485,N_1422,N_1406);
nand U1486 (N_1486,N_1377,N_1351);
or U1487 (N_1487,N_1398,N_1368);
nor U1488 (N_1488,N_1420,N_1364);
or U1489 (N_1489,N_1368,N_1400);
and U1490 (N_1490,N_1387,N_1391);
nor U1491 (N_1491,N_1351,N_1410);
nand U1492 (N_1492,N_1380,N_1390);
or U1493 (N_1493,N_1392,N_1388);
nand U1494 (N_1494,N_1408,N_1400);
nand U1495 (N_1495,N_1369,N_1401);
nor U1496 (N_1496,N_1391,N_1355);
or U1497 (N_1497,N_1420,N_1358);
and U1498 (N_1498,N_1414,N_1388);
and U1499 (N_1499,N_1387,N_1401);
nand U1500 (N_1500,N_1462,N_1483);
nor U1501 (N_1501,N_1463,N_1452);
nand U1502 (N_1502,N_1427,N_1484);
nand U1503 (N_1503,N_1443,N_1458);
nand U1504 (N_1504,N_1490,N_1441);
or U1505 (N_1505,N_1476,N_1453);
and U1506 (N_1506,N_1466,N_1464);
xor U1507 (N_1507,N_1498,N_1440);
nor U1508 (N_1508,N_1426,N_1485);
nor U1509 (N_1509,N_1432,N_1425);
or U1510 (N_1510,N_1497,N_1492);
or U1511 (N_1511,N_1455,N_1437);
nor U1512 (N_1512,N_1428,N_1496);
nor U1513 (N_1513,N_1436,N_1480);
nor U1514 (N_1514,N_1435,N_1487);
nor U1515 (N_1515,N_1470,N_1486);
nand U1516 (N_1516,N_1446,N_1489);
nand U1517 (N_1517,N_1454,N_1444);
nand U1518 (N_1518,N_1451,N_1450);
nand U1519 (N_1519,N_1445,N_1442);
nand U1520 (N_1520,N_1429,N_1469);
or U1521 (N_1521,N_1491,N_1456);
xor U1522 (N_1522,N_1431,N_1449);
nand U1523 (N_1523,N_1474,N_1459);
or U1524 (N_1524,N_1499,N_1467);
or U1525 (N_1525,N_1461,N_1448);
nor U1526 (N_1526,N_1473,N_1439);
nand U1527 (N_1527,N_1472,N_1471);
nor U1528 (N_1528,N_1468,N_1488);
nand U1529 (N_1529,N_1475,N_1465);
nand U1530 (N_1530,N_1493,N_1457);
nor U1531 (N_1531,N_1434,N_1460);
nand U1532 (N_1532,N_1482,N_1447);
or U1533 (N_1533,N_1478,N_1479);
nor U1534 (N_1534,N_1481,N_1495);
nor U1535 (N_1535,N_1430,N_1438);
and U1536 (N_1536,N_1433,N_1494);
or U1537 (N_1537,N_1477,N_1467);
nand U1538 (N_1538,N_1485,N_1484);
or U1539 (N_1539,N_1466,N_1481);
or U1540 (N_1540,N_1487,N_1459);
or U1541 (N_1541,N_1469,N_1477);
xnor U1542 (N_1542,N_1447,N_1498);
nor U1543 (N_1543,N_1479,N_1491);
nor U1544 (N_1544,N_1451,N_1473);
nor U1545 (N_1545,N_1448,N_1455);
nor U1546 (N_1546,N_1461,N_1440);
or U1547 (N_1547,N_1441,N_1480);
nand U1548 (N_1548,N_1492,N_1426);
nor U1549 (N_1549,N_1464,N_1453);
and U1550 (N_1550,N_1428,N_1429);
or U1551 (N_1551,N_1493,N_1450);
nand U1552 (N_1552,N_1431,N_1479);
and U1553 (N_1553,N_1499,N_1482);
nand U1554 (N_1554,N_1475,N_1441);
nand U1555 (N_1555,N_1466,N_1433);
and U1556 (N_1556,N_1499,N_1439);
nor U1557 (N_1557,N_1475,N_1438);
nand U1558 (N_1558,N_1437,N_1487);
or U1559 (N_1559,N_1464,N_1437);
and U1560 (N_1560,N_1471,N_1485);
nor U1561 (N_1561,N_1467,N_1452);
nand U1562 (N_1562,N_1453,N_1443);
and U1563 (N_1563,N_1468,N_1452);
nor U1564 (N_1564,N_1426,N_1482);
and U1565 (N_1565,N_1439,N_1442);
nand U1566 (N_1566,N_1437,N_1483);
nor U1567 (N_1567,N_1459,N_1428);
nor U1568 (N_1568,N_1480,N_1499);
nor U1569 (N_1569,N_1429,N_1491);
nor U1570 (N_1570,N_1459,N_1497);
and U1571 (N_1571,N_1478,N_1460);
nor U1572 (N_1572,N_1488,N_1453);
or U1573 (N_1573,N_1480,N_1481);
xor U1574 (N_1574,N_1426,N_1455);
nand U1575 (N_1575,N_1540,N_1538);
or U1576 (N_1576,N_1521,N_1519);
and U1577 (N_1577,N_1502,N_1568);
or U1578 (N_1578,N_1541,N_1550);
nand U1579 (N_1579,N_1534,N_1552);
nor U1580 (N_1580,N_1559,N_1536);
or U1581 (N_1581,N_1517,N_1562);
or U1582 (N_1582,N_1542,N_1547);
nand U1583 (N_1583,N_1535,N_1513);
and U1584 (N_1584,N_1564,N_1523);
or U1585 (N_1585,N_1510,N_1555);
xor U1586 (N_1586,N_1505,N_1558);
nand U1587 (N_1587,N_1512,N_1549);
nor U1588 (N_1588,N_1574,N_1573);
or U1589 (N_1589,N_1561,N_1514);
and U1590 (N_1590,N_1501,N_1557);
nand U1591 (N_1591,N_1506,N_1503);
nand U1592 (N_1592,N_1504,N_1544);
and U1593 (N_1593,N_1530,N_1511);
xor U1594 (N_1594,N_1524,N_1527);
nand U1595 (N_1595,N_1529,N_1525);
nor U1596 (N_1596,N_1516,N_1570);
nor U1597 (N_1597,N_1554,N_1548);
nand U1598 (N_1598,N_1526,N_1539);
or U1599 (N_1599,N_1567,N_1546);
nor U1600 (N_1600,N_1522,N_1572);
nor U1601 (N_1601,N_1532,N_1507);
and U1602 (N_1602,N_1556,N_1571);
nand U1603 (N_1603,N_1508,N_1500);
nand U1604 (N_1604,N_1551,N_1553);
nor U1605 (N_1605,N_1528,N_1509);
and U1606 (N_1606,N_1545,N_1569);
nor U1607 (N_1607,N_1560,N_1520);
or U1608 (N_1608,N_1531,N_1515);
nand U1609 (N_1609,N_1533,N_1543);
nor U1610 (N_1610,N_1537,N_1565);
or U1611 (N_1611,N_1566,N_1518);
or U1612 (N_1612,N_1563,N_1525);
nand U1613 (N_1613,N_1504,N_1528);
and U1614 (N_1614,N_1566,N_1556);
or U1615 (N_1615,N_1549,N_1538);
nand U1616 (N_1616,N_1500,N_1558);
nand U1617 (N_1617,N_1563,N_1560);
or U1618 (N_1618,N_1542,N_1564);
and U1619 (N_1619,N_1537,N_1528);
or U1620 (N_1620,N_1538,N_1528);
and U1621 (N_1621,N_1573,N_1519);
and U1622 (N_1622,N_1546,N_1513);
or U1623 (N_1623,N_1568,N_1540);
nand U1624 (N_1624,N_1556,N_1501);
or U1625 (N_1625,N_1519,N_1556);
nor U1626 (N_1626,N_1574,N_1532);
nor U1627 (N_1627,N_1525,N_1538);
or U1628 (N_1628,N_1502,N_1524);
and U1629 (N_1629,N_1542,N_1543);
and U1630 (N_1630,N_1531,N_1500);
or U1631 (N_1631,N_1551,N_1528);
or U1632 (N_1632,N_1502,N_1519);
or U1633 (N_1633,N_1573,N_1516);
or U1634 (N_1634,N_1546,N_1526);
xnor U1635 (N_1635,N_1530,N_1508);
or U1636 (N_1636,N_1563,N_1565);
nand U1637 (N_1637,N_1524,N_1500);
and U1638 (N_1638,N_1552,N_1540);
nor U1639 (N_1639,N_1558,N_1562);
nor U1640 (N_1640,N_1554,N_1557);
nand U1641 (N_1641,N_1523,N_1514);
xor U1642 (N_1642,N_1562,N_1504);
and U1643 (N_1643,N_1537,N_1530);
nor U1644 (N_1644,N_1514,N_1571);
and U1645 (N_1645,N_1542,N_1502);
nand U1646 (N_1646,N_1573,N_1561);
nand U1647 (N_1647,N_1532,N_1524);
xor U1648 (N_1648,N_1531,N_1558);
nor U1649 (N_1649,N_1547,N_1574);
nor U1650 (N_1650,N_1583,N_1577);
nor U1651 (N_1651,N_1579,N_1614);
and U1652 (N_1652,N_1602,N_1581);
xor U1653 (N_1653,N_1609,N_1601);
or U1654 (N_1654,N_1628,N_1632);
nand U1655 (N_1655,N_1630,N_1623);
nand U1656 (N_1656,N_1580,N_1624);
nor U1657 (N_1657,N_1610,N_1640);
and U1658 (N_1658,N_1578,N_1582);
nor U1659 (N_1659,N_1604,N_1600);
and U1660 (N_1660,N_1648,N_1576);
or U1661 (N_1661,N_1584,N_1616);
nor U1662 (N_1662,N_1622,N_1594);
and U1663 (N_1663,N_1606,N_1592);
nand U1664 (N_1664,N_1588,N_1618);
or U1665 (N_1665,N_1643,N_1617);
nor U1666 (N_1666,N_1631,N_1575);
nor U1667 (N_1667,N_1593,N_1615);
nand U1668 (N_1668,N_1597,N_1599);
nand U1669 (N_1669,N_1603,N_1627);
nand U1670 (N_1670,N_1598,N_1612);
xnor U1671 (N_1671,N_1626,N_1587);
nor U1672 (N_1672,N_1585,N_1636);
or U1673 (N_1673,N_1642,N_1586);
nand U1674 (N_1674,N_1621,N_1607);
nor U1675 (N_1675,N_1645,N_1619);
xor U1676 (N_1676,N_1620,N_1641);
and U1677 (N_1677,N_1629,N_1635);
and U1678 (N_1678,N_1596,N_1608);
nand U1679 (N_1679,N_1638,N_1591);
or U1680 (N_1680,N_1595,N_1589);
and U1681 (N_1681,N_1649,N_1590);
nand U1682 (N_1682,N_1644,N_1647);
or U1683 (N_1683,N_1646,N_1611);
nor U1684 (N_1684,N_1639,N_1633);
nand U1685 (N_1685,N_1637,N_1634);
nor U1686 (N_1686,N_1605,N_1625);
nand U1687 (N_1687,N_1613,N_1623);
nand U1688 (N_1688,N_1605,N_1576);
nor U1689 (N_1689,N_1639,N_1592);
nand U1690 (N_1690,N_1584,N_1644);
nor U1691 (N_1691,N_1600,N_1576);
nand U1692 (N_1692,N_1640,N_1635);
and U1693 (N_1693,N_1639,N_1638);
nor U1694 (N_1694,N_1596,N_1628);
or U1695 (N_1695,N_1632,N_1619);
nor U1696 (N_1696,N_1609,N_1600);
nor U1697 (N_1697,N_1620,N_1644);
and U1698 (N_1698,N_1629,N_1604);
nor U1699 (N_1699,N_1637,N_1644);
and U1700 (N_1700,N_1612,N_1603);
nor U1701 (N_1701,N_1638,N_1631);
or U1702 (N_1702,N_1587,N_1603);
nand U1703 (N_1703,N_1624,N_1600);
nand U1704 (N_1704,N_1607,N_1613);
and U1705 (N_1705,N_1613,N_1608);
or U1706 (N_1706,N_1588,N_1589);
nor U1707 (N_1707,N_1644,N_1633);
and U1708 (N_1708,N_1641,N_1630);
nor U1709 (N_1709,N_1636,N_1602);
nor U1710 (N_1710,N_1578,N_1610);
nand U1711 (N_1711,N_1610,N_1592);
nand U1712 (N_1712,N_1643,N_1622);
nor U1713 (N_1713,N_1628,N_1619);
nor U1714 (N_1714,N_1606,N_1629);
nand U1715 (N_1715,N_1587,N_1595);
nand U1716 (N_1716,N_1579,N_1612);
nor U1717 (N_1717,N_1583,N_1582);
and U1718 (N_1718,N_1579,N_1619);
and U1719 (N_1719,N_1617,N_1632);
or U1720 (N_1720,N_1603,N_1649);
or U1721 (N_1721,N_1595,N_1636);
nor U1722 (N_1722,N_1635,N_1644);
or U1723 (N_1723,N_1605,N_1612);
or U1724 (N_1724,N_1645,N_1589);
nand U1725 (N_1725,N_1650,N_1713);
nand U1726 (N_1726,N_1689,N_1683);
nor U1727 (N_1727,N_1692,N_1668);
and U1728 (N_1728,N_1672,N_1704);
and U1729 (N_1729,N_1708,N_1676);
nor U1730 (N_1730,N_1690,N_1662);
or U1731 (N_1731,N_1685,N_1652);
or U1732 (N_1732,N_1681,N_1712);
or U1733 (N_1733,N_1691,N_1719);
xnor U1734 (N_1734,N_1673,N_1653);
and U1735 (N_1735,N_1658,N_1663);
and U1736 (N_1736,N_1657,N_1682);
and U1737 (N_1737,N_1695,N_1655);
or U1738 (N_1738,N_1666,N_1667);
or U1739 (N_1739,N_1696,N_1687);
nor U1740 (N_1740,N_1665,N_1693);
nand U1741 (N_1741,N_1705,N_1697);
nand U1742 (N_1742,N_1675,N_1659);
nand U1743 (N_1743,N_1723,N_1709);
xor U1744 (N_1744,N_1686,N_1699);
and U1745 (N_1745,N_1660,N_1671);
and U1746 (N_1746,N_1707,N_1678);
nor U1747 (N_1747,N_1724,N_1670);
xor U1748 (N_1748,N_1706,N_1688);
nand U1749 (N_1749,N_1674,N_1722);
or U1750 (N_1750,N_1656,N_1698);
or U1751 (N_1751,N_1715,N_1718);
nand U1752 (N_1752,N_1694,N_1710);
nor U1753 (N_1753,N_1701,N_1679);
xor U1754 (N_1754,N_1700,N_1720);
nor U1755 (N_1755,N_1654,N_1661);
or U1756 (N_1756,N_1711,N_1669);
nor U1757 (N_1757,N_1703,N_1721);
or U1758 (N_1758,N_1664,N_1717);
nand U1759 (N_1759,N_1677,N_1680);
nand U1760 (N_1760,N_1684,N_1714);
nand U1761 (N_1761,N_1651,N_1716);
nand U1762 (N_1762,N_1702,N_1665);
nand U1763 (N_1763,N_1690,N_1650);
or U1764 (N_1764,N_1695,N_1707);
nor U1765 (N_1765,N_1681,N_1652);
and U1766 (N_1766,N_1719,N_1697);
nand U1767 (N_1767,N_1667,N_1703);
and U1768 (N_1768,N_1710,N_1701);
and U1769 (N_1769,N_1693,N_1677);
nand U1770 (N_1770,N_1703,N_1672);
or U1771 (N_1771,N_1679,N_1673);
nor U1772 (N_1772,N_1724,N_1715);
or U1773 (N_1773,N_1719,N_1656);
and U1774 (N_1774,N_1661,N_1695);
and U1775 (N_1775,N_1724,N_1669);
nor U1776 (N_1776,N_1667,N_1691);
or U1777 (N_1777,N_1699,N_1659);
nand U1778 (N_1778,N_1663,N_1656);
nand U1779 (N_1779,N_1660,N_1650);
or U1780 (N_1780,N_1710,N_1662);
nand U1781 (N_1781,N_1689,N_1687);
nor U1782 (N_1782,N_1714,N_1685);
nand U1783 (N_1783,N_1706,N_1692);
or U1784 (N_1784,N_1719,N_1690);
nand U1785 (N_1785,N_1657,N_1711);
nor U1786 (N_1786,N_1661,N_1709);
xnor U1787 (N_1787,N_1677,N_1650);
nand U1788 (N_1788,N_1690,N_1660);
or U1789 (N_1789,N_1658,N_1664);
nor U1790 (N_1790,N_1679,N_1709);
and U1791 (N_1791,N_1667,N_1660);
nor U1792 (N_1792,N_1706,N_1658);
and U1793 (N_1793,N_1691,N_1721);
nand U1794 (N_1794,N_1663,N_1711);
and U1795 (N_1795,N_1699,N_1715);
nand U1796 (N_1796,N_1717,N_1702);
nand U1797 (N_1797,N_1661,N_1706);
and U1798 (N_1798,N_1657,N_1680);
nor U1799 (N_1799,N_1672,N_1713);
or U1800 (N_1800,N_1740,N_1738);
nand U1801 (N_1801,N_1759,N_1741);
nor U1802 (N_1802,N_1776,N_1788);
nor U1803 (N_1803,N_1784,N_1747);
and U1804 (N_1804,N_1764,N_1780);
nor U1805 (N_1805,N_1760,N_1730);
nor U1806 (N_1806,N_1775,N_1797);
or U1807 (N_1807,N_1728,N_1729);
nor U1808 (N_1808,N_1725,N_1782);
nor U1809 (N_1809,N_1739,N_1766);
and U1810 (N_1810,N_1743,N_1787);
xnor U1811 (N_1811,N_1785,N_1726);
nor U1812 (N_1812,N_1774,N_1768);
nor U1813 (N_1813,N_1735,N_1734);
nand U1814 (N_1814,N_1794,N_1761);
nor U1815 (N_1815,N_1752,N_1736);
and U1816 (N_1816,N_1781,N_1790);
or U1817 (N_1817,N_1771,N_1744);
and U1818 (N_1818,N_1742,N_1750);
nand U1819 (N_1819,N_1762,N_1758);
nor U1820 (N_1820,N_1767,N_1748);
nand U1821 (N_1821,N_1798,N_1751);
nand U1822 (N_1822,N_1763,N_1753);
nor U1823 (N_1823,N_1754,N_1746);
or U1824 (N_1824,N_1731,N_1778);
or U1825 (N_1825,N_1791,N_1786);
nand U1826 (N_1826,N_1727,N_1757);
or U1827 (N_1827,N_1770,N_1732);
and U1828 (N_1828,N_1772,N_1796);
or U1829 (N_1829,N_1783,N_1779);
and U1830 (N_1830,N_1765,N_1749);
xnor U1831 (N_1831,N_1792,N_1789);
and U1832 (N_1832,N_1737,N_1793);
xor U1833 (N_1833,N_1756,N_1773);
and U1834 (N_1834,N_1745,N_1799);
and U1835 (N_1835,N_1769,N_1755);
nand U1836 (N_1836,N_1777,N_1733);
and U1837 (N_1837,N_1795,N_1755);
or U1838 (N_1838,N_1729,N_1748);
nand U1839 (N_1839,N_1727,N_1749);
and U1840 (N_1840,N_1792,N_1751);
nand U1841 (N_1841,N_1753,N_1745);
nand U1842 (N_1842,N_1795,N_1745);
and U1843 (N_1843,N_1792,N_1757);
nand U1844 (N_1844,N_1725,N_1751);
nor U1845 (N_1845,N_1759,N_1758);
or U1846 (N_1846,N_1785,N_1781);
and U1847 (N_1847,N_1747,N_1782);
nand U1848 (N_1848,N_1751,N_1749);
and U1849 (N_1849,N_1799,N_1748);
nand U1850 (N_1850,N_1771,N_1765);
and U1851 (N_1851,N_1739,N_1728);
nor U1852 (N_1852,N_1737,N_1751);
or U1853 (N_1853,N_1783,N_1757);
nor U1854 (N_1854,N_1764,N_1771);
nor U1855 (N_1855,N_1752,N_1774);
nor U1856 (N_1856,N_1798,N_1744);
nor U1857 (N_1857,N_1743,N_1799);
nand U1858 (N_1858,N_1731,N_1753);
xnor U1859 (N_1859,N_1785,N_1750);
xnor U1860 (N_1860,N_1752,N_1726);
xor U1861 (N_1861,N_1788,N_1779);
and U1862 (N_1862,N_1766,N_1733);
and U1863 (N_1863,N_1731,N_1769);
nor U1864 (N_1864,N_1741,N_1728);
nand U1865 (N_1865,N_1764,N_1743);
nor U1866 (N_1866,N_1767,N_1759);
and U1867 (N_1867,N_1773,N_1797);
nand U1868 (N_1868,N_1789,N_1737);
nand U1869 (N_1869,N_1744,N_1791);
and U1870 (N_1870,N_1792,N_1746);
or U1871 (N_1871,N_1788,N_1749);
and U1872 (N_1872,N_1729,N_1774);
nor U1873 (N_1873,N_1765,N_1728);
and U1874 (N_1874,N_1737,N_1755);
and U1875 (N_1875,N_1852,N_1856);
nor U1876 (N_1876,N_1853,N_1860);
or U1877 (N_1877,N_1813,N_1804);
nand U1878 (N_1878,N_1857,N_1859);
or U1879 (N_1879,N_1855,N_1843);
or U1880 (N_1880,N_1863,N_1874);
nor U1881 (N_1881,N_1817,N_1805);
and U1882 (N_1882,N_1824,N_1810);
or U1883 (N_1883,N_1827,N_1866);
nand U1884 (N_1884,N_1825,N_1838);
and U1885 (N_1885,N_1842,N_1867);
or U1886 (N_1886,N_1848,N_1829);
nor U1887 (N_1887,N_1832,N_1820);
and U1888 (N_1888,N_1873,N_1816);
or U1889 (N_1889,N_1801,N_1869);
nor U1890 (N_1890,N_1850,N_1809);
and U1891 (N_1891,N_1858,N_1822);
nand U1892 (N_1892,N_1851,N_1814);
nand U1893 (N_1893,N_1831,N_1839);
and U1894 (N_1894,N_1849,N_1830);
and U1895 (N_1895,N_1841,N_1802);
nand U1896 (N_1896,N_1870,N_1861);
nand U1897 (N_1897,N_1812,N_1840);
or U1898 (N_1898,N_1819,N_1847);
nor U1899 (N_1899,N_1845,N_1808);
xnor U1900 (N_1900,N_1854,N_1835);
and U1901 (N_1901,N_1868,N_1844);
and U1902 (N_1902,N_1871,N_1833);
nor U1903 (N_1903,N_1800,N_1872);
nand U1904 (N_1904,N_1807,N_1862);
and U1905 (N_1905,N_1803,N_1834);
or U1906 (N_1906,N_1836,N_1828);
nor U1907 (N_1907,N_1806,N_1815);
and U1908 (N_1908,N_1864,N_1826);
and U1909 (N_1909,N_1865,N_1818);
nor U1910 (N_1910,N_1837,N_1846);
or U1911 (N_1911,N_1811,N_1821);
nand U1912 (N_1912,N_1823,N_1858);
nand U1913 (N_1913,N_1847,N_1863);
and U1914 (N_1914,N_1861,N_1810);
and U1915 (N_1915,N_1848,N_1850);
or U1916 (N_1916,N_1840,N_1874);
or U1917 (N_1917,N_1808,N_1856);
nor U1918 (N_1918,N_1864,N_1818);
nor U1919 (N_1919,N_1832,N_1813);
nand U1920 (N_1920,N_1866,N_1834);
or U1921 (N_1921,N_1800,N_1870);
nor U1922 (N_1922,N_1872,N_1815);
nor U1923 (N_1923,N_1871,N_1870);
or U1924 (N_1924,N_1850,N_1839);
or U1925 (N_1925,N_1845,N_1838);
and U1926 (N_1926,N_1800,N_1812);
nand U1927 (N_1927,N_1836,N_1845);
or U1928 (N_1928,N_1865,N_1821);
or U1929 (N_1929,N_1809,N_1854);
or U1930 (N_1930,N_1812,N_1807);
or U1931 (N_1931,N_1861,N_1851);
or U1932 (N_1932,N_1852,N_1861);
or U1933 (N_1933,N_1850,N_1859);
and U1934 (N_1934,N_1863,N_1857);
and U1935 (N_1935,N_1863,N_1850);
and U1936 (N_1936,N_1854,N_1836);
nor U1937 (N_1937,N_1830,N_1815);
nor U1938 (N_1938,N_1849,N_1859);
nand U1939 (N_1939,N_1849,N_1851);
and U1940 (N_1940,N_1864,N_1851);
and U1941 (N_1941,N_1869,N_1855);
and U1942 (N_1942,N_1847,N_1859);
xor U1943 (N_1943,N_1806,N_1851);
nand U1944 (N_1944,N_1800,N_1818);
and U1945 (N_1945,N_1828,N_1851);
or U1946 (N_1946,N_1842,N_1808);
or U1947 (N_1947,N_1809,N_1871);
nand U1948 (N_1948,N_1806,N_1813);
nand U1949 (N_1949,N_1822,N_1845);
nand U1950 (N_1950,N_1902,N_1934);
nand U1951 (N_1951,N_1925,N_1946);
nand U1952 (N_1952,N_1918,N_1882);
and U1953 (N_1953,N_1877,N_1938);
nand U1954 (N_1954,N_1906,N_1891);
xnor U1955 (N_1955,N_1904,N_1905);
xnor U1956 (N_1956,N_1899,N_1915);
or U1957 (N_1957,N_1917,N_1909);
nand U1958 (N_1958,N_1920,N_1897);
nand U1959 (N_1959,N_1923,N_1942);
nor U1960 (N_1960,N_1895,N_1875);
or U1961 (N_1961,N_1886,N_1949);
nor U1962 (N_1962,N_1878,N_1935);
nor U1963 (N_1963,N_1928,N_1940);
and U1964 (N_1964,N_1910,N_1885);
nor U1965 (N_1965,N_1911,N_1884);
and U1966 (N_1966,N_1919,N_1936);
and U1967 (N_1967,N_1892,N_1908);
nor U1968 (N_1968,N_1901,N_1890);
nor U1969 (N_1969,N_1929,N_1883);
and U1970 (N_1970,N_1879,N_1894);
nor U1971 (N_1971,N_1893,N_1948);
nor U1972 (N_1972,N_1926,N_1907);
or U1973 (N_1973,N_1900,N_1903);
nand U1974 (N_1974,N_1933,N_1927);
nor U1975 (N_1975,N_1913,N_1932);
and U1976 (N_1976,N_1945,N_1881);
nor U1977 (N_1977,N_1924,N_1896);
or U1978 (N_1978,N_1944,N_1939);
nand U1979 (N_1979,N_1947,N_1912);
nand U1980 (N_1980,N_1931,N_1898);
and U1981 (N_1981,N_1930,N_1880);
or U1982 (N_1982,N_1941,N_1887);
and U1983 (N_1983,N_1916,N_1922);
or U1984 (N_1984,N_1914,N_1888);
and U1985 (N_1985,N_1943,N_1889);
nor U1986 (N_1986,N_1921,N_1876);
or U1987 (N_1987,N_1937,N_1888);
nor U1988 (N_1988,N_1933,N_1883);
nand U1989 (N_1989,N_1934,N_1935);
nor U1990 (N_1990,N_1893,N_1910);
nor U1991 (N_1991,N_1946,N_1877);
and U1992 (N_1992,N_1936,N_1916);
or U1993 (N_1993,N_1945,N_1933);
nor U1994 (N_1994,N_1922,N_1907);
nand U1995 (N_1995,N_1919,N_1938);
or U1996 (N_1996,N_1901,N_1933);
nor U1997 (N_1997,N_1883,N_1889);
or U1998 (N_1998,N_1892,N_1891);
and U1999 (N_1999,N_1881,N_1936);
and U2000 (N_2000,N_1934,N_1895);
or U2001 (N_2001,N_1931,N_1928);
nor U2002 (N_2002,N_1902,N_1940);
or U2003 (N_2003,N_1892,N_1921);
and U2004 (N_2004,N_1945,N_1929);
nor U2005 (N_2005,N_1928,N_1889);
nor U2006 (N_2006,N_1892,N_1896);
and U2007 (N_2007,N_1930,N_1934);
or U2008 (N_2008,N_1904,N_1927);
nand U2009 (N_2009,N_1906,N_1926);
nand U2010 (N_2010,N_1890,N_1905);
or U2011 (N_2011,N_1927,N_1883);
or U2012 (N_2012,N_1930,N_1928);
nand U2013 (N_2013,N_1935,N_1884);
nand U2014 (N_2014,N_1925,N_1889);
and U2015 (N_2015,N_1934,N_1892);
nand U2016 (N_2016,N_1905,N_1884);
nor U2017 (N_2017,N_1929,N_1880);
or U2018 (N_2018,N_1898,N_1893);
xnor U2019 (N_2019,N_1901,N_1888);
and U2020 (N_2020,N_1876,N_1905);
and U2021 (N_2021,N_1897,N_1909);
nor U2022 (N_2022,N_1885,N_1879);
or U2023 (N_2023,N_1911,N_1921);
or U2024 (N_2024,N_1922,N_1941);
nand U2025 (N_2025,N_2024,N_2023);
nor U2026 (N_2026,N_1978,N_1961);
and U2027 (N_2027,N_2003,N_1966);
nor U2028 (N_2028,N_1996,N_1998);
nor U2029 (N_2029,N_2011,N_1985);
and U2030 (N_2030,N_1991,N_1979);
nand U2031 (N_2031,N_1972,N_2010);
or U2032 (N_2032,N_1983,N_1981);
and U2033 (N_2033,N_2012,N_1951);
and U2034 (N_2034,N_2006,N_2015);
and U2035 (N_2035,N_1989,N_1960);
xnor U2036 (N_2036,N_1992,N_2002);
nor U2037 (N_2037,N_2016,N_1955);
nand U2038 (N_2038,N_1965,N_1963);
xnor U2039 (N_2039,N_2022,N_2009);
or U2040 (N_2040,N_1988,N_2001);
and U2041 (N_2041,N_2017,N_1997);
or U2042 (N_2042,N_1953,N_1982);
nor U2043 (N_2043,N_1962,N_2004);
and U2044 (N_2044,N_1990,N_2020);
xnor U2045 (N_2045,N_2021,N_2019);
nor U2046 (N_2046,N_1980,N_1994);
nor U2047 (N_2047,N_1958,N_1959);
nor U2048 (N_2048,N_1986,N_1957);
xor U2049 (N_2049,N_1954,N_1952);
or U2050 (N_2050,N_1995,N_1976);
nor U2051 (N_2051,N_2018,N_2013);
nand U2052 (N_2052,N_1974,N_1987);
and U2053 (N_2053,N_1977,N_1993);
and U2054 (N_2054,N_1970,N_1967);
nor U2055 (N_2055,N_2005,N_1973);
nand U2056 (N_2056,N_1956,N_1969);
or U2057 (N_2057,N_1984,N_2007);
and U2058 (N_2058,N_1950,N_1971);
nor U2059 (N_2059,N_1999,N_1968);
nor U2060 (N_2060,N_1964,N_2014);
nand U2061 (N_2061,N_2008,N_2000);
xnor U2062 (N_2062,N_1975,N_2004);
or U2063 (N_2063,N_2001,N_1981);
and U2064 (N_2064,N_1984,N_1972);
nor U2065 (N_2065,N_1983,N_1958);
nand U2066 (N_2066,N_1977,N_1951);
nor U2067 (N_2067,N_1957,N_1962);
nor U2068 (N_2068,N_2021,N_1973);
nor U2069 (N_2069,N_1957,N_1952);
or U2070 (N_2070,N_2014,N_2001);
nor U2071 (N_2071,N_1953,N_2008);
nor U2072 (N_2072,N_2023,N_2006);
xnor U2073 (N_2073,N_1962,N_1993);
or U2074 (N_2074,N_1952,N_2008);
and U2075 (N_2075,N_1998,N_2014);
and U2076 (N_2076,N_1993,N_1963);
nand U2077 (N_2077,N_2013,N_1978);
or U2078 (N_2078,N_1958,N_1961);
and U2079 (N_2079,N_1959,N_1951);
and U2080 (N_2080,N_1998,N_1995);
nand U2081 (N_2081,N_2002,N_1995);
nand U2082 (N_2082,N_1970,N_1977);
nor U2083 (N_2083,N_1955,N_2021);
or U2084 (N_2084,N_1996,N_1968);
nor U2085 (N_2085,N_1974,N_2013);
nand U2086 (N_2086,N_2024,N_2010);
and U2087 (N_2087,N_2019,N_2011);
nor U2088 (N_2088,N_1978,N_1951);
or U2089 (N_2089,N_1951,N_1965);
or U2090 (N_2090,N_1981,N_2006);
or U2091 (N_2091,N_1976,N_2001);
or U2092 (N_2092,N_1976,N_2005);
nor U2093 (N_2093,N_2022,N_1968);
and U2094 (N_2094,N_2021,N_2001);
nor U2095 (N_2095,N_2019,N_2007);
or U2096 (N_2096,N_1999,N_1990);
nor U2097 (N_2097,N_1996,N_1960);
and U2098 (N_2098,N_1986,N_1961);
nor U2099 (N_2099,N_1978,N_1974);
nor U2100 (N_2100,N_2048,N_2046);
or U2101 (N_2101,N_2044,N_2086);
nand U2102 (N_2102,N_2073,N_2074);
or U2103 (N_2103,N_2037,N_2090);
and U2104 (N_2104,N_2076,N_2084);
or U2105 (N_2105,N_2030,N_2039);
nand U2106 (N_2106,N_2087,N_2035);
nor U2107 (N_2107,N_2032,N_2094);
nor U2108 (N_2108,N_2027,N_2072);
or U2109 (N_2109,N_2066,N_2045);
or U2110 (N_2110,N_2042,N_2050);
nand U2111 (N_2111,N_2091,N_2069);
nor U2112 (N_2112,N_2096,N_2053);
and U2113 (N_2113,N_2059,N_2075);
or U2114 (N_2114,N_2036,N_2067);
and U2115 (N_2115,N_2047,N_2031);
nor U2116 (N_2116,N_2028,N_2026);
and U2117 (N_2117,N_2097,N_2071);
nor U2118 (N_2118,N_2040,N_2034);
nor U2119 (N_2119,N_2064,N_2041);
or U2120 (N_2120,N_2082,N_2070);
nand U2121 (N_2121,N_2052,N_2080);
xor U2122 (N_2122,N_2079,N_2055);
nor U2123 (N_2123,N_2077,N_2025);
nor U2124 (N_2124,N_2078,N_2049);
and U2125 (N_2125,N_2029,N_2098);
nor U2126 (N_2126,N_2038,N_2093);
nand U2127 (N_2127,N_2061,N_2065);
nor U2128 (N_2128,N_2083,N_2058);
nor U2129 (N_2129,N_2056,N_2088);
or U2130 (N_2130,N_2060,N_2057);
and U2131 (N_2131,N_2081,N_2062);
nor U2132 (N_2132,N_2085,N_2054);
nand U2133 (N_2133,N_2095,N_2099);
nand U2134 (N_2134,N_2043,N_2063);
nand U2135 (N_2135,N_2092,N_2089);
and U2136 (N_2136,N_2051,N_2068);
nor U2137 (N_2137,N_2033,N_2058);
and U2138 (N_2138,N_2047,N_2077);
nand U2139 (N_2139,N_2064,N_2051);
and U2140 (N_2140,N_2071,N_2058);
and U2141 (N_2141,N_2074,N_2072);
nand U2142 (N_2142,N_2051,N_2060);
or U2143 (N_2143,N_2042,N_2072);
nor U2144 (N_2144,N_2093,N_2086);
nor U2145 (N_2145,N_2058,N_2060);
and U2146 (N_2146,N_2061,N_2028);
nor U2147 (N_2147,N_2079,N_2035);
or U2148 (N_2148,N_2097,N_2049);
xor U2149 (N_2149,N_2072,N_2053);
or U2150 (N_2150,N_2036,N_2042);
or U2151 (N_2151,N_2044,N_2071);
and U2152 (N_2152,N_2084,N_2061);
or U2153 (N_2153,N_2033,N_2065);
nor U2154 (N_2154,N_2035,N_2065);
nor U2155 (N_2155,N_2070,N_2049);
or U2156 (N_2156,N_2058,N_2048);
nand U2157 (N_2157,N_2025,N_2026);
or U2158 (N_2158,N_2080,N_2068);
or U2159 (N_2159,N_2058,N_2034);
nor U2160 (N_2160,N_2036,N_2048);
nor U2161 (N_2161,N_2086,N_2076);
nor U2162 (N_2162,N_2082,N_2089);
nand U2163 (N_2163,N_2076,N_2087);
nor U2164 (N_2164,N_2096,N_2060);
xnor U2165 (N_2165,N_2028,N_2064);
or U2166 (N_2166,N_2079,N_2078);
or U2167 (N_2167,N_2081,N_2027);
xnor U2168 (N_2168,N_2062,N_2070);
or U2169 (N_2169,N_2048,N_2037);
or U2170 (N_2170,N_2033,N_2098);
and U2171 (N_2171,N_2092,N_2098);
nand U2172 (N_2172,N_2027,N_2099);
nor U2173 (N_2173,N_2048,N_2080);
nor U2174 (N_2174,N_2040,N_2045);
nor U2175 (N_2175,N_2138,N_2160);
and U2176 (N_2176,N_2115,N_2150);
xnor U2177 (N_2177,N_2161,N_2112);
or U2178 (N_2178,N_2171,N_2147);
nand U2179 (N_2179,N_2157,N_2141);
or U2180 (N_2180,N_2108,N_2142);
nor U2181 (N_2181,N_2123,N_2114);
or U2182 (N_2182,N_2168,N_2173);
and U2183 (N_2183,N_2103,N_2104);
nor U2184 (N_2184,N_2156,N_2120);
and U2185 (N_2185,N_2102,N_2131);
nand U2186 (N_2186,N_2170,N_2174);
nand U2187 (N_2187,N_2132,N_2149);
xnor U2188 (N_2188,N_2158,N_2127);
or U2189 (N_2189,N_2121,N_2151);
nand U2190 (N_2190,N_2105,N_2137);
nand U2191 (N_2191,N_2113,N_2136);
nor U2192 (N_2192,N_2152,N_2169);
and U2193 (N_2193,N_2110,N_2118);
nand U2194 (N_2194,N_2163,N_2143);
and U2195 (N_2195,N_2135,N_2144);
and U2196 (N_2196,N_2126,N_2140);
nand U2197 (N_2197,N_2125,N_2139);
or U2198 (N_2198,N_2134,N_2111);
and U2199 (N_2199,N_2129,N_2162);
or U2200 (N_2200,N_2124,N_2109);
and U2201 (N_2201,N_2128,N_2106);
or U2202 (N_2202,N_2107,N_2153);
nand U2203 (N_2203,N_2166,N_2165);
nand U2204 (N_2204,N_2167,N_2101);
or U2205 (N_2205,N_2133,N_2155);
or U2206 (N_2206,N_2154,N_2119);
or U2207 (N_2207,N_2100,N_2148);
nor U2208 (N_2208,N_2122,N_2117);
or U2209 (N_2209,N_2116,N_2172);
nand U2210 (N_2210,N_2159,N_2130);
and U2211 (N_2211,N_2164,N_2145);
nor U2212 (N_2212,N_2146,N_2117);
and U2213 (N_2213,N_2111,N_2170);
or U2214 (N_2214,N_2130,N_2102);
nor U2215 (N_2215,N_2116,N_2140);
and U2216 (N_2216,N_2104,N_2144);
nand U2217 (N_2217,N_2122,N_2158);
and U2218 (N_2218,N_2106,N_2112);
nor U2219 (N_2219,N_2166,N_2151);
or U2220 (N_2220,N_2165,N_2103);
nand U2221 (N_2221,N_2136,N_2110);
or U2222 (N_2222,N_2121,N_2122);
or U2223 (N_2223,N_2152,N_2135);
and U2224 (N_2224,N_2119,N_2152);
nand U2225 (N_2225,N_2116,N_2168);
or U2226 (N_2226,N_2115,N_2147);
nand U2227 (N_2227,N_2126,N_2152);
nand U2228 (N_2228,N_2133,N_2149);
or U2229 (N_2229,N_2104,N_2122);
or U2230 (N_2230,N_2167,N_2174);
or U2231 (N_2231,N_2138,N_2125);
or U2232 (N_2232,N_2121,N_2160);
nand U2233 (N_2233,N_2167,N_2120);
and U2234 (N_2234,N_2121,N_2170);
or U2235 (N_2235,N_2163,N_2156);
or U2236 (N_2236,N_2165,N_2144);
nor U2237 (N_2237,N_2109,N_2153);
xnor U2238 (N_2238,N_2113,N_2165);
nand U2239 (N_2239,N_2119,N_2146);
nor U2240 (N_2240,N_2129,N_2134);
nor U2241 (N_2241,N_2132,N_2169);
nor U2242 (N_2242,N_2128,N_2165);
and U2243 (N_2243,N_2155,N_2139);
or U2244 (N_2244,N_2168,N_2151);
nand U2245 (N_2245,N_2167,N_2141);
and U2246 (N_2246,N_2146,N_2104);
and U2247 (N_2247,N_2125,N_2148);
or U2248 (N_2248,N_2126,N_2135);
or U2249 (N_2249,N_2145,N_2151);
nor U2250 (N_2250,N_2245,N_2198);
xor U2251 (N_2251,N_2232,N_2199);
nor U2252 (N_2252,N_2185,N_2188);
or U2253 (N_2253,N_2244,N_2191);
or U2254 (N_2254,N_2216,N_2249);
nor U2255 (N_2255,N_2226,N_2192);
and U2256 (N_2256,N_2242,N_2222);
and U2257 (N_2257,N_2177,N_2219);
nand U2258 (N_2258,N_2205,N_2248);
nor U2259 (N_2259,N_2190,N_2221);
nor U2260 (N_2260,N_2233,N_2230);
nand U2261 (N_2261,N_2217,N_2215);
and U2262 (N_2262,N_2224,N_2189);
nor U2263 (N_2263,N_2218,N_2208);
and U2264 (N_2264,N_2212,N_2234);
and U2265 (N_2265,N_2179,N_2195);
nand U2266 (N_2266,N_2200,N_2202);
nand U2267 (N_2267,N_2238,N_2183);
and U2268 (N_2268,N_2180,N_2211);
or U2269 (N_2269,N_2209,N_2196);
nand U2270 (N_2270,N_2178,N_2236);
nor U2271 (N_2271,N_2237,N_2214);
nand U2272 (N_2272,N_2186,N_2220);
nand U2273 (N_2273,N_2213,N_2207);
nand U2274 (N_2274,N_2201,N_2193);
or U2275 (N_2275,N_2181,N_2204);
or U2276 (N_2276,N_2176,N_2210);
nand U2277 (N_2277,N_2197,N_2225);
nor U2278 (N_2278,N_2227,N_2247);
or U2279 (N_2279,N_2223,N_2184);
nand U2280 (N_2280,N_2187,N_2203);
or U2281 (N_2281,N_2235,N_2246);
and U2282 (N_2282,N_2231,N_2239);
or U2283 (N_2283,N_2194,N_2243);
nor U2284 (N_2284,N_2175,N_2241);
nor U2285 (N_2285,N_2182,N_2228);
nand U2286 (N_2286,N_2240,N_2229);
and U2287 (N_2287,N_2206,N_2196);
nand U2288 (N_2288,N_2178,N_2247);
and U2289 (N_2289,N_2236,N_2249);
and U2290 (N_2290,N_2221,N_2184);
and U2291 (N_2291,N_2200,N_2237);
or U2292 (N_2292,N_2229,N_2227);
nand U2293 (N_2293,N_2213,N_2242);
nor U2294 (N_2294,N_2236,N_2207);
nor U2295 (N_2295,N_2212,N_2201);
or U2296 (N_2296,N_2249,N_2199);
or U2297 (N_2297,N_2218,N_2188);
nor U2298 (N_2298,N_2202,N_2192);
nand U2299 (N_2299,N_2185,N_2216);
nor U2300 (N_2300,N_2192,N_2240);
xnor U2301 (N_2301,N_2191,N_2210);
or U2302 (N_2302,N_2224,N_2190);
nor U2303 (N_2303,N_2187,N_2211);
or U2304 (N_2304,N_2232,N_2198);
and U2305 (N_2305,N_2231,N_2182);
nor U2306 (N_2306,N_2229,N_2195);
or U2307 (N_2307,N_2213,N_2186);
nand U2308 (N_2308,N_2180,N_2223);
or U2309 (N_2309,N_2176,N_2226);
or U2310 (N_2310,N_2209,N_2187);
or U2311 (N_2311,N_2227,N_2244);
and U2312 (N_2312,N_2241,N_2240);
nand U2313 (N_2313,N_2201,N_2223);
nand U2314 (N_2314,N_2229,N_2234);
or U2315 (N_2315,N_2233,N_2235);
and U2316 (N_2316,N_2228,N_2221);
xor U2317 (N_2317,N_2181,N_2192);
or U2318 (N_2318,N_2200,N_2240);
or U2319 (N_2319,N_2226,N_2235);
nand U2320 (N_2320,N_2240,N_2191);
and U2321 (N_2321,N_2198,N_2201);
nand U2322 (N_2322,N_2246,N_2202);
or U2323 (N_2323,N_2245,N_2177);
or U2324 (N_2324,N_2239,N_2230);
and U2325 (N_2325,N_2310,N_2292);
nand U2326 (N_2326,N_2311,N_2306);
nand U2327 (N_2327,N_2258,N_2313);
nor U2328 (N_2328,N_2256,N_2262);
or U2329 (N_2329,N_2252,N_2300);
nor U2330 (N_2330,N_2280,N_2287);
or U2331 (N_2331,N_2291,N_2281);
and U2332 (N_2332,N_2303,N_2255);
or U2333 (N_2333,N_2295,N_2301);
nor U2334 (N_2334,N_2277,N_2305);
nand U2335 (N_2335,N_2251,N_2308);
xor U2336 (N_2336,N_2317,N_2273);
nand U2337 (N_2337,N_2307,N_2289);
nor U2338 (N_2338,N_2314,N_2284);
and U2339 (N_2339,N_2266,N_2318);
and U2340 (N_2340,N_2309,N_2322);
and U2341 (N_2341,N_2288,N_2267);
xnor U2342 (N_2342,N_2319,N_2250);
or U2343 (N_2343,N_2320,N_2294);
or U2344 (N_2344,N_2269,N_2264);
and U2345 (N_2345,N_2276,N_2272);
and U2346 (N_2346,N_2323,N_2283);
and U2347 (N_2347,N_2279,N_2253);
or U2348 (N_2348,N_2293,N_2286);
and U2349 (N_2349,N_2282,N_2285);
and U2350 (N_2350,N_2290,N_2275);
and U2351 (N_2351,N_2304,N_2312);
and U2352 (N_2352,N_2324,N_2297);
and U2353 (N_2353,N_2257,N_2260);
or U2354 (N_2354,N_2259,N_2302);
nand U2355 (N_2355,N_2270,N_2321);
nor U2356 (N_2356,N_2278,N_2254);
nor U2357 (N_2357,N_2298,N_2296);
nand U2358 (N_2358,N_2261,N_2265);
xor U2359 (N_2359,N_2315,N_2271);
nor U2360 (N_2360,N_2316,N_2268);
nor U2361 (N_2361,N_2274,N_2299);
and U2362 (N_2362,N_2263,N_2314);
or U2363 (N_2363,N_2323,N_2319);
and U2364 (N_2364,N_2319,N_2324);
or U2365 (N_2365,N_2268,N_2287);
or U2366 (N_2366,N_2290,N_2286);
and U2367 (N_2367,N_2313,N_2294);
nor U2368 (N_2368,N_2282,N_2259);
or U2369 (N_2369,N_2279,N_2311);
nor U2370 (N_2370,N_2267,N_2308);
nor U2371 (N_2371,N_2294,N_2262);
and U2372 (N_2372,N_2320,N_2306);
or U2373 (N_2373,N_2273,N_2287);
and U2374 (N_2374,N_2275,N_2309);
or U2375 (N_2375,N_2279,N_2292);
or U2376 (N_2376,N_2314,N_2318);
or U2377 (N_2377,N_2260,N_2270);
nand U2378 (N_2378,N_2291,N_2318);
and U2379 (N_2379,N_2321,N_2274);
and U2380 (N_2380,N_2266,N_2281);
nand U2381 (N_2381,N_2289,N_2259);
and U2382 (N_2382,N_2275,N_2272);
and U2383 (N_2383,N_2302,N_2305);
and U2384 (N_2384,N_2294,N_2301);
nor U2385 (N_2385,N_2287,N_2309);
nand U2386 (N_2386,N_2271,N_2282);
nor U2387 (N_2387,N_2311,N_2264);
nor U2388 (N_2388,N_2306,N_2300);
nor U2389 (N_2389,N_2286,N_2277);
nor U2390 (N_2390,N_2300,N_2299);
nand U2391 (N_2391,N_2311,N_2275);
nand U2392 (N_2392,N_2288,N_2308);
or U2393 (N_2393,N_2311,N_2257);
or U2394 (N_2394,N_2324,N_2317);
nor U2395 (N_2395,N_2283,N_2282);
nor U2396 (N_2396,N_2262,N_2299);
nor U2397 (N_2397,N_2311,N_2263);
and U2398 (N_2398,N_2290,N_2252);
and U2399 (N_2399,N_2265,N_2311);
nand U2400 (N_2400,N_2388,N_2335);
and U2401 (N_2401,N_2391,N_2348);
nand U2402 (N_2402,N_2379,N_2346);
and U2403 (N_2403,N_2373,N_2332);
and U2404 (N_2404,N_2381,N_2399);
or U2405 (N_2405,N_2331,N_2340);
and U2406 (N_2406,N_2366,N_2338);
or U2407 (N_2407,N_2330,N_2396);
or U2408 (N_2408,N_2394,N_2384);
nand U2409 (N_2409,N_2361,N_2343);
or U2410 (N_2410,N_2363,N_2352);
nand U2411 (N_2411,N_2393,N_2326);
or U2412 (N_2412,N_2350,N_2353);
nand U2413 (N_2413,N_2336,N_2337);
or U2414 (N_2414,N_2351,N_2378);
or U2415 (N_2415,N_2333,N_2385);
nand U2416 (N_2416,N_2344,N_2397);
and U2417 (N_2417,N_2367,N_2345);
and U2418 (N_2418,N_2398,N_2356);
or U2419 (N_2419,N_2325,N_2375);
nor U2420 (N_2420,N_2395,N_2328);
or U2421 (N_2421,N_2368,N_2386);
nand U2422 (N_2422,N_2372,N_2364);
nor U2423 (N_2423,N_2334,N_2342);
nor U2424 (N_2424,N_2389,N_2365);
or U2425 (N_2425,N_2392,N_2374);
and U2426 (N_2426,N_2371,N_2387);
nand U2427 (N_2427,N_2383,N_2329);
and U2428 (N_2428,N_2347,N_2380);
nor U2429 (N_2429,N_2377,N_2357);
nand U2430 (N_2430,N_2358,N_2355);
nor U2431 (N_2431,N_2360,N_2359);
or U2432 (N_2432,N_2382,N_2327);
and U2433 (N_2433,N_2370,N_2349);
nor U2434 (N_2434,N_2339,N_2341);
or U2435 (N_2435,N_2376,N_2369);
xor U2436 (N_2436,N_2390,N_2354);
or U2437 (N_2437,N_2362,N_2361);
and U2438 (N_2438,N_2336,N_2391);
and U2439 (N_2439,N_2381,N_2365);
nand U2440 (N_2440,N_2378,N_2376);
and U2441 (N_2441,N_2328,N_2385);
nor U2442 (N_2442,N_2364,N_2356);
or U2443 (N_2443,N_2394,N_2387);
and U2444 (N_2444,N_2366,N_2358);
or U2445 (N_2445,N_2373,N_2349);
nand U2446 (N_2446,N_2342,N_2328);
or U2447 (N_2447,N_2380,N_2378);
and U2448 (N_2448,N_2342,N_2395);
nor U2449 (N_2449,N_2395,N_2359);
or U2450 (N_2450,N_2374,N_2342);
and U2451 (N_2451,N_2366,N_2326);
and U2452 (N_2452,N_2380,N_2343);
and U2453 (N_2453,N_2357,N_2379);
nand U2454 (N_2454,N_2387,N_2390);
xor U2455 (N_2455,N_2346,N_2325);
and U2456 (N_2456,N_2390,N_2381);
nand U2457 (N_2457,N_2327,N_2375);
nor U2458 (N_2458,N_2329,N_2340);
and U2459 (N_2459,N_2357,N_2335);
and U2460 (N_2460,N_2340,N_2381);
and U2461 (N_2461,N_2351,N_2353);
nor U2462 (N_2462,N_2339,N_2357);
and U2463 (N_2463,N_2353,N_2365);
nand U2464 (N_2464,N_2326,N_2378);
nor U2465 (N_2465,N_2327,N_2337);
nor U2466 (N_2466,N_2331,N_2344);
nor U2467 (N_2467,N_2376,N_2386);
or U2468 (N_2468,N_2394,N_2377);
and U2469 (N_2469,N_2337,N_2339);
and U2470 (N_2470,N_2382,N_2369);
or U2471 (N_2471,N_2343,N_2397);
nand U2472 (N_2472,N_2348,N_2364);
nand U2473 (N_2473,N_2395,N_2369);
nand U2474 (N_2474,N_2343,N_2393);
nand U2475 (N_2475,N_2417,N_2461);
or U2476 (N_2476,N_2441,N_2448);
and U2477 (N_2477,N_2432,N_2426);
nand U2478 (N_2478,N_2460,N_2434);
nand U2479 (N_2479,N_2428,N_2452);
nand U2480 (N_2480,N_2474,N_2401);
nor U2481 (N_2481,N_2457,N_2408);
nand U2482 (N_2482,N_2421,N_2450);
nor U2483 (N_2483,N_2453,N_2471);
nor U2484 (N_2484,N_2456,N_2447);
nand U2485 (N_2485,N_2455,N_2416);
and U2486 (N_2486,N_2451,N_2402);
nand U2487 (N_2487,N_2438,N_2407);
or U2488 (N_2488,N_2435,N_2462);
nand U2489 (N_2489,N_2403,N_2444);
nand U2490 (N_2490,N_2466,N_2430);
nor U2491 (N_2491,N_2446,N_2463);
nand U2492 (N_2492,N_2419,N_2415);
and U2493 (N_2493,N_2413,N_2449);
nor U2494 (N_2494,N_2427,N_2445);
nor U2495 (N_2495,N_2439,N_2400);
and U2496 (N_2496,N_2422,N_2409);
nand U2497 (N_2497,N_2429,N_2442);
nand U2498 (N_2498,N_2414,N_2458);
or U2499 (N_2499,N_2406,N_2470);
and U2500 (N_2500,N_2431,N_2437);
nor U2501 (N_2501,N_2433,N_2418);
nand U2502 (N_2502,N_2454,N_2473);
and U2503 (N_2503,N_2468,N_2404);
or U2504 (N_2504,N_2440,N_2412);
nand U2505 (N_2505,N_2443,N_2425);
nand U2506 (N_2506,N_2423,N_2420);
nand U2507 (N_2507,N_2459,N_2424);
nor U2508 (N_2508,N_2436,N_2467);
and U2509 (N_2509,N_2464,N_2469);
nand U2510 (N_2510,N_2472,N_2411);
nand U2511 (N_2511,N_2465,N_2405);
or U2512 (N_2512,N_2410,N_2402);
or U2513 (N_2513,N_2423,N_2432);
or U2514 (N_2514,N_2414,N_2419);
and U2515 (N_2515,N_2423,N_2446);
and U2516 (N_2516,N_2402,N_2441);
or U2517 (N_2517,N_2458,N_2407);
nand U2518 (N_2518,N_2433,N_2447);
nor U2519 (N_2519,N_2466,N_2459);
nor U2520 (N_2520,N_2453,N_2400);
and U2521 (N_2521,N_2463,N_2415);
and U2522 (N_2522,N_2414,N_2436);
or U2523 (N_2523,N_2414,N_2417);
nor U2524 (N_2524,N_2422,N_2464);
nor U2525 (N_2525,N_2442,N_2428);
or U2526 (N_2526,N_2451,N_2409);
nor U2527 (N_2527,N_2455,N_2433);
nor U2528 (N_2528,N_2473,N_2449);
and U2529 (N_2529,N_2457,N_2411);
nand U2530 (N_2530,N_2453,N_2469);
or U2531 (N_2531,N_2439,N_2456);
and U2532 (N_2532,N_2422,N_2454);
or U2533 (N_2533,N_2449,N_2471);
nor U2534 (N_2534,N_2458,N_2400);
or U2535 (N_2535,N_2416,N_2444);
or U2536 (N_2536,N_2418,N_2437);
or U2537 (N_2537,N_2461,N_2400);
nor U2538 (N_2538,N_2404,N_2441);
or U2539 (N_2539,N_2429,N_2450);
and U2540 (N_2540,N_2424,N_2444);
nand U2541 (N_2541,N_2408,N_2415);
or U2542 (N_2542,N_2432,N_2452);
and U2543 (N_2543,N_2423,N_2471);
nor U2544 (N_2544,N_2426,N_2409);
nand U2545 (N_2545,N_2428,N_2423);
or U2546 (N_2546,N_2402,N_2449);
nand U2547 (N_2547,N_2444,N_2461);
nor U2548 (N_2548,N_2438,N_2410);
nand U2549 (N_2549,N_2438,N_2428);
and U2550 (N_2550,N_2506,N_2517);
and U2551 (N_2551,N_2486,N_2509);
or U2552 (N_2552,N_2503,N_2526);
and U2553 (N_2553,N_2540,N_2501);
or U2554 (N_2554,N_2488,N_2476);
nor U2555 (N_2555,N_2521,N_2481);
nor U2556 (N_2556,N_2527,N_2542);
or U2557 (N_2557,N_2516,N_2484);
xor U2558 (N_2558,N_2492,N_2479);
nand U2559 (N_2559,N_2538,N_2544);
nor U2560 (N_2560,N_2525,N_2500);
or U2561 (N_2561,N_2528,N_2537);
or U2562 (N_2562,N_2512,N_2498);
and U2563 (N_2563,N_2475,N_2531);
nor U2564 (N_2564,N_2532,N_2518);
nor U2565 (N_2565,N_2545,N_2504);
xnor U2566 (N_2566,N_2543,N_2522);
nor U2567 (N_2567,N_2497,N_2491);
nand U2568 (N_2568,N_2523,N_2487);
nor U2569 (N_2569,N_2477,N_2519);
or U2570 (N_2570,N_2502,N_2511);
or U2571 (N_2571,N_2546,N_2489);
or U2572 (N_2572,N_2496,N_2548);
nor U2573 (N_2573,N_2539,N_2541);
and U2574 (N_2574,N_2495,N_2478);
and U2575 (N_2575,N_2505,N_2535);
nand U2576 (N_2576,N_2530,N_2508);
nand U2577 (N_2577,N_2524,N_2515);
nand U2578 (N_2578,N_2507,N_2482);
or U2579 (N_2579,N_2533,N_2510);
nand U2580 (N_2580,N_2529,N_2547);
nand U2581 (N_2581,N_2494,N_2513);
nand U2582 (N_2582,N_2490,N_2536);
nand U2583 (N_2583,N_2493,N_2514);
nor U2584 (N_2584,N_2520,N_2549);
or U2585 (N_2585,N_2499,N_2483);
or U2586 (N_2586,N_2480,N_2485);
nand U2587 (N_2587,N_2534,N_2542);
nor U2588 (N_2588,N_2504,N_2517);
nand U2589 (N_2589,N_2489,N_2495);
and U2590 (N_2590,N_2496,N_2490);
nand U2591 (N_2591,N_2530,N_2493);
nor U2592 (N_2592,N_2525,N_2496);
and U2593 (N_2593,N_2477,N_2475);
and U2594 (N_2594,N_2527,N_2481);
and U2595 (N_2595,N_2527,N_2511);
and U2596 (N_2596,N_2533,N_2531);
and U2597 (N_2597,N_2541,N_2477);
nor U2598 (N_2598,N_2482,N_2478);
nand U2599 (N_2599,N_2482,N_2513);
nand U2600 (N_2600,N_2497,N_2489);
and U2601 (N_2601,N_2512,N_2526);
and U2602 (N_2602,N_2511,N_2530);
nand U2603 (N_2603,N_2501,N_2500);
nor U2604 (N_2604,N_2524,N_2478);
nor U2605 (N_2605,N_2543,N_2491);
nor U2606 (N_2606,N_2496,N_2513);
nor U2607 (N_2607,N_2530,N_2539);
nand U2608 (N_2608,N_2494,N_2512);
nand U2609 (N_2609,N_2496,N_2482);
xnor U2610 (N_2610,N_2520,N_2505);
and U2611 (N_2611,N_2536,N_2540);
xor U2612 (N_2612,N_2548,N_2484);
and U2613 (N_2613,N_2544,N_2485);
nand U2614 (N_2614,N_2520,N_2537);
nor U2615 (N_2615,N_2523,N_2530);
and U2616 (N_2616,N_2516,N_2537);
nand U2617 (N_2617,N_2487,N_2479);
and U2618 (N_2618,N_2523,N_2478);
or U2619 (N_2619,N_2498,N_2506);
and U2620 (N_2620,N_2523,N_2526);
and U2621 (N_2621,N_2517,N_2490);
nand U2622 (N_2622,N_2485,N_2499);
nor U2623 (N_2623,N_2507,N_2549);
nor U2624 (N_2624,N_2535,N_2483);
nand U2625 (N_2625,N_2578,N_2592);
nor U2626 (N_2626,N_2590,N_2586);
nor U2627 (N_2627,N_2572,N_2576);
nor U2628 (N_2628,N_2554,N_2589);
and U2629 (N_2629,N_2620,N_2574);
nor U2630 (N_2630,N_2597,N_2612);
nor U2631 (N_2631,N_2565,N_2596);
xor U2632 (N_2632,N_2558,N_2577);
xor U2633 (N_2633,N_2619,N_2568);
nand U2634 (N_2634,N_2608,N_2622);
nand U2635 (N_2635,N_2580,N_2553);
and U2636 (N_2636,N_2569,N_2606);
or U2637 (N_2637,N_2605,N_2551);
nor U2638 (N_2638,N_2595,N_2613);
nand U2639 (N_2639,N_2611,N_2579);
and U2640 (N_2640,N_2601,N_2618);
nand U2641 (N_2641,N_2567,N_2594);
nand U2642 (N_2642,N_2600,N_2584);
or U2643 (N_2643,N_2591,N_2621);
and U2644 (N_2644,N_2614,N_2583);
nand U2645 (N_2645,N_2552,N_2598);
or U2646 (N_2646,N_2602,N_2561);
nor U2647 (N_2647,N_2624,N_2563);
or U2648 (N_2648,N_2617,N_2571);
nor U2649 (N_2649,N_2610,N_2616);
nor U2650 (N_2650,N_2582,N_2559);
nand U2651 (N_2651,N_2585,N_2550);
nor U2652 (N_2652,N_2587,N_2599);
nand U2653 (N_2653,N_2615,N_2603);
nor U2654 (N_2654,N_2607,N_2555);
nor U2655 (N_2655,N_2573,N_2570);
and U2656 (N_2656,N_2556,N_2604);
nand U2657 (N_2657,N_2588,N_2609);
nor U2658 (N_2658,N_2566,N_2564);
nor U2659 (N_2659,N_2575,N_2623);
or U2660 (N_2660,N_2581,N_2557);
and U2661 (N_2661,N_2593,N_2560);
nor U2662 (N_2662,N_2562,N_2590);
or U2663 (N_2663,N_2551,N_2620);
nand U2664 (N_2664,N_2558,N_2619);
nand U2665 (N_2665,N_2604,N_2598);
and U2666 (N_2666,N_2565,N_2598);
nor U2667 (N_2667,N_2561,N_2586);
nand U2668 (N_2668,N_2585,N_2566);
nor U2669 (N_2669,N_2601,N_2593);
or U2670 (N_2670,N_2552,N_2578);
and U2671 (N_2671,N_2583,N_2586);
nand U2672 (N_2672,N_2575,N_2578);
xnor U2673 (N_2673,N_2569,N_2557);
nand U2674 (N_2674,N_2605,N_2622);
and U2675 (N_2675,N_2606,N_2609);
or U2676 (N_2676,N_2585,N_2590);
xnor U2677 (N_2677,N_2591,N_2610);
and U2678 (N_2678,N_2578,N_2572);
nor U2679 (N_2679,N_2618,N_2622);
or U2680 (N_2680,N_2551,N_2600);
nor U2681 (N_2681,N_2586,N_2572);
nand U2682 (N_2682,N_2601,N_2597);
nand U2683 (N_2683,N_2587,N_2552);
and U2684 (N_2684,N_2585,N_2573);
nor U2685 (N_2685,N_2604,N_2607);
or U2686 (N_2686,N_2623,N_2601);
or U2687 (N_2687,N_2551,N_2593);
and U2688 (N_2688,N_2572,N_2557);
or U2689 (N_2689,N_2592,N_2598);
nand U2690 (N_2690,N_2558,N_2620);
nand U2691 (N_2691,N_2575,N_2601);
nand U2692 (N_2692,N_2597,N_2575);
or U2693 (N_2693,N_2586,N_2551);
nor U2694 (N_2694,N_2614,N_2576);
nor U2695 (N_2695,N_2564,N_2604);
nor U2696 (N_2696,N_2607,N_2594);
nor U2697 (N_2697,N_2609,N_2599);
or U2698 (N_2698,N_2623,N_2591);
nand U2699 (N_2699,N_2602,N_2596);
or U2700 (N_2700,N_2630,N_2695);
or U2701 (N_2701,N_2625,N_2635);
and U2702 (N_2702,N_2669,N_2673);
or U2703 (N_2703,N_2670,N_2686);
nand U2704 (N_2704,N_2664,N_2639);
nand U2705 (N_2705,N_2658,N_2674);
nand U2706 (N_2706,N_2683,N_2638);
nor U2707 (N_2707,N_2634,N_2663);
or U2708 (N_2708,N_2648,N_2667);
nand U2709 (N_2709,N_2665,N_2641);
nor U2710 (N_2710,N_2629,N_2697);
nand U2711 (N_2711,N_2680,N_2644);
or U2712 (N_2712,N_2672,N_2685);
nand U2713 (N_2713,N_2666,N_2632);
nor U2714 (N_2714,N_2676,N_2653);
nand U2715 (N_2715,N_2668,N_2637);
nand U2716 (N_2716,N_2647,N_2691);
nand U2717 (N_2717,N_2699,N_2682);
or U2718 (N_2718,N_2677,N_2656);
or U2719 (N_2719,N_2687,N_2655);
and U2720 (N_2720,N_2675,N_2690);
nand U2721 (N_2721,N_2679,N_2633);
and U2722 (N_2722,N_2636,N_2631);
nand U2723 (N_2723,N_2696,N_2642);
and U2724 (N_2724,N_2694,N_2654);
nand U2725 (N_2725,N_2640,N_2643);
and U2726 (N_2726,N_2693,N_2627);
or U2727 (N_2727,N_2659,N_2698);
nor U2728 (N_2728,N_2657,N_2628);
or U2729 (N_2729,N_2651,N_2688);
nor U2730 (N_2730,N_2689,N_2662);
nor U2731 (N_2731,N_2661,N_2660);
nor U2732 (N_2732,N_2649,N_2646);
and U2733 (N_2733,N_2692,N_2671);
nor U2734 (N_2734,N_2681,N_2678);
nand U2735 (N_2735,N_2626,N_2684);
and U2736 (N_2736,N_2652,N_2645);
and U2737 (N_2737,N_2650,N_2638);
or U2738 (N_2738,N_2662,N_2677);
or U2739 (N_2739,N_2659,N_2642);
nor U2740 (N_2740,N_2650,N_2666);
nor U2741 (N_2741,N_2655,N_2691);
and U2742 (N_2742,N_2664,N_2688);
nand U2743 (N_2743,N_2647,N_2665);
nand U2744 (N_2744,N_2652,N_2625);
nand U2745 (N_2745,N_2687,N_2651);
nand U2746 (N_2746,N_2664,N_2647);
nor U2747 (N_2747,N_2670,N_2643);
and U2748 (N_2748,N_2656,N_2636);
and U2749 (N_2749,N_2643,N_2649);
and U2750 (N_2750,N_2662,N_2679);
nor U2751 (N_2751,N_2633,N_2698);
nand U2752 (N_2752,N_2693,N_2659);
nand U2753 (N_2753,N_2675,N_2669);
and U2754 (N_2754,N_2672,N_2662);
and U2755 (N_2755,N_2638,N_2676);
and U2756 (N_2756,N_2652,N_2634);
or U2757 (N_2757,N_2636,N_2671);
or U2758 (N_2758,N_2632,N_2643);
and U2759 (N_2759,N_2664,N_2634);
or U2760 (N_2760,N_2675,N_2695);
and U2761 (N_2761,N_2651,N_2670);
or U2762 (N_2762,N_2698,N_2649);
and U2763 (N_2763,N_2679,N_2625);
nor U2764 (N_2764,N_2690,N_2657);
xnor U2765 (N_2765,N_2683,N_2642);
and U2766 (N_2766,N_2691,N_2643);
nand U2767 (N_2767,N_2692,N_2665);
xnor U2768 (N_2768,N_2635,N_2685);
or U2769 (N_2769,N_2685,N_2642);
and U2770 (N_2770,N_2681,N_2652);
nor U2771 (N_2771,N_2674,N_2691);
nor U2772 (N_2772,N_2641,N_2675);
and U2773 (N_2773,N_2646,N_2633);
nor U2774 (N_2774,N_2642,N_2634);
or U2775 (N_2775,N_2719,N_2755);
and U2776 (N_2776,N_2760,N_2753);
or U2777 (N_2777,N_2750,N_2703);
or U2778 (N_2778,N_2739,N_2770);
or U2779 (N_2779,N_2705,N_2742);
or U2780 (N_2780,N_2730,N_2736);
nand U2781 (N_2781,N_2746,N_2731);
nor U2782 (N_2782,N_2749,N_2732);
nand U2783 (N_2783,N_2740,N_2704);
and U2784 (N_2784,N_2772,N_2737);
or U2785 (N_2785,N_2717,N_2774);
nand U2786 (N_2786,N_2728,N_2727);
xnor U2787 (N_2787,N_2744,N_2735);
and U2788 (N_2788,N_2706,N_2763);
nor U2789 (N_2789,N_2708,N_2764);
nor U2790 (N_2790,N_2715,N_2747);
and U2791 (N_2791,N_2700,N_2762);
and U2792 (N_2792,N_2748,N_2713);
and U2793 (N_2793,N_2765,N_2714);
or U2794 (N_2794,N_2771,N_2710);
nand U2795 (N_2795,N_2712,N_2720);
and U2796 (N_2796,N_2724,N_2722);
nand U2797 (N_2797,N_2701,N_2767);
nand U2798 (N_2798,N_2766,N_2752);
nand U2799 (N_2799,N_2745,N_2707);
xor U2800 (N_2800,N_2759,N_2768);
or U2801 (N_2801,N_2758,N_2729);
nand U2802 (N_2802,N_2723,N_2716);
and U2803 (N_2803,N_2733,N_2769);
nor U2804 (N_2804,N_2757,N_2711);
and U2805 (N_2805,N_2743,N_2751);
and U2806 (N_2806,N_2754,N_2726);
and U2807 (N_2807,N_2773,N_2709);
xnor U2808 (N_2808,N_2761,N_2718);
nand U2809 (N_2809,N_2738,N_2702);
and U2810 (N_2810,N_2741,N_2725);
and U2811 (N_2811,N_2721,N_2734);
or U2812 (N_2812,N_2756,N_2733);
nand U2813 (N_2813,N_2708,N_2721);
or U2814 (N_2814,N_2738,N_2720);
and U2815 (N_2815,N_2740,N_2724);
and U2816 (N_2816,N_2730,N_2747);
nand U2817 (N_2817,N_2716,N_2717);
nor U2818 (N_2818,N_2726,N_2700);
and U2819 (N_2819,N_2714,N_2752);
or U2820 (N_2820,N_2747,N_2772);
nor U2821 (N_2821,N_2762,N_2770);
nor U2822 (N_2822,N_2734,N_2770);
and U2823 (N_2823,N_2740,N_2703);
nor U2824 (N_2824,N_2765,N_2749);
or U2825 (N_2825,N_2742,N_2732);
nand U2826 (N_2826,N_2736,N_2709);
nand U2827 (N_2827,N_2709,N_2715);
or U2828 (N_2828,N_2770,N_2710);
nor U2829 (N_2829,N_2721,N_2771);
and U2830 (N_2830,N_2767,N_2765);
and U2831 (N_2831,N_2700,N_2737);
nand U2832 (N_2832,N_2767,N_2700);
nor U2833 (N_2833,N_2748,N_2762);
nor U2834 (N_2834,N_2757,N_2746);
nor U2835 (N_2835,N_2700,N_2707);
and U2836 (N_2836,N_2712,N_2736);
nor U2837 (N_2837,N_2768,N_2748);
and U2838 (N_2838,N_2725,N_2754);
xnor U2839 (N_2839,N_2745,N_2763);
and U2840 (N_2840,N_2741,N_2723);
nand U2841 (N_2841,N_2747,N_2755);
or U2842 (N_2842,N_2764,N_2710);
nand U2843 (N_2843,N_2730,N_2764);
and U2844 (N_2844,N_2708,N_2729);
and U2845 (N_2845,N_2735,N_2724);
or U2846 (N_2846,N_2720,N_2727);
nor U2847 (N_2847,N_2728,N_2719);
and U2848 (N_2848,N_2760,N_2740);
and U2849 (N_2849,N_2738,N_2743);
and U2850 (N_2850,N_2815,N_2810);
and U2851 (N_2851,N_2814,N_2777);
or U2852 (N_2852,N_2825,N_2835);
nor U2853 (N_2853,N_2782,N_2786);
nor U2854 (N_2854,N_2793,N_2802);
nor U2855 (N_2855,N_2827,N_2845);
nand U2856 (N_2856,N_2797,N_2840);
and U2857 (N_2857,N_2842,N_2824);
nand U2858 (N_2858,N_2809,N_2801);
and U2859 (N_2859,N_2785,N_2832);
and U2860 (N_2860,N_2843,N_2790);
nand U2861 (N_2861,N_2775,N_2778);
nand U2862 (N_2862,N_2780,N_2826);
xor U2863 (N_2863,N_2795,N_2818);
nand U2864 (N_2864,N_2804,N_2817);
nand U2865 (N_2865,N_2834,N_2830);
nor U2866 (N_2866,N_2807,N_2823);
nor U2867 (N_2867,N_2806,N_2787);
and U2868 (N_2868,N_2836,N_2816);
nor U2869 (N_2869,N_2811,N_2847);
nand U2870 (N_2870,N_2805,N_2789);
and U2871 (N_2871,N_2798,N_2821);
or U2872 (N_2872,N_2794,N_2819);
nor U2873 (N_2873,N_2800,N_2791);
or U2874 (N_2874,N_2783,N_2796);
or U2875 (N_2875,N_2779,N_2828);
nor U2876 (N_2876,N_2784,N_2838);
or U2877 (N_2877,N_2792,N_2788);
nand U2878 (N_2878,N_2822,N_2846);
and U2879 (N_2879,N_2820,N_2844);
nand U2880 (N_2880,N_2841,N_2839);
nor U2881 (N_2881,N_2808,N_2837);
nor U2882 (N_2882,N_2776,N_2849);
nand U2883 (N_2883,N_2813,N_2803);
and U2884 (N_2884,N_2812,N_2831);
or U2885 (N_2885,N_2833,N_2848);
and U2886 (N_2886,N_2829,N_2799);
nand U2887 (N_2887,N_2781,N_2826);
nand U2888 (N_2888,N_2833,N_2794);
xnor U2889 (N_2889,N_2835,N_2775);
nor U2890 (N_2890,N_2794,N_2811);
nor U2891 (N_2891,N_2791,N_2790);
or U2892 (N_2892,N_2784,N_2816);
nand U2893 (N_2893,N_2782,N_2796);
nor U2894 (N_2894,N_2836,N_2828);
and U2895 (N_2895,N_2840,N_2815);
nand U2896 (N_2896,N_2791,N_2844);
or U2897 (N_2897,N_2840,N_2847);
or U2898 (N_2898,N_2792,N_2797);
and U2899 (N_2899,N_2834,N_2811);
nand U2900 (N_2900,N_2847,N_2836);
nor U2901 (N_2901,N_2837,N_2795);
or U2902 (N_2902,N_2801,N_2844);
and U2903 (N_2903,N_2813,N_2806);
or U2904 (N_2904,N_2779,N_2838);
or U2905 (N_2905,N_2809,N_2806);
and U2906 (N_2906,N_2824,N_2783);
nand U2907 (N_2907,N_2781,N_2789);
nand U2908 (N_2908,N_2827,N_2800);
or U2909 (N_2909,N_2796,N_2787);
and U2910 (N_2910,N_2830,N_2841);
nor U2911 (N_2911,N_2787,N_2843);
or U2912 (N_2912,N_2823,N_2833);
nand U2913 (N_2913,N_2789,N_2808);
and U2914 (N_2914,N_2821,N_2834);
nor U2915 (N_2915,N_2849,N_2836);
nor U2916 (N_2916,N_2793,N_2848);
nor U2917 (N_2917,N_2781,N_2783);
nand U2918 (N_2918,N_2792,N_2841);
or U2919 (N_2919,N_2813,N_2825);
nor U2920 (N_2920,N_2779,N_2845);
and U2921 (N_2921,N_2817,N_2848);
xor U2922 (N_2922,N_2782,N_2803);
or U2923 (N_2923,N_2777,N_2783);
nand U2924 (N_2924,N_2782,N_2838);
nand U2925 (N_2925,N_2878,N_2885);
nor U2926 (N_2926,N_2888,N_2882);
nor U2927 (N_2927,N_2898,N_2879);
and U2928 (N_2928,N_2922,N_2902);
or U2929 (N_2929,N_2851,N_2856);
or U2930 (N_2930,N_2904,N_2874);
or U2931 (N_2931,N_2860,N_2894);
nand U2932 (N_2932,N_2899,N_2912);
nor U2933 (N_2933,N_2864,N_2896);
and U2934 (N_2934,N_2873,N_2900);
xor U2935 (N_2935,N_2881,N_2870);
nor U2936 (N_2936,N_2886,N_2923);
and U2937 (N_2937,N_2858,N_2869);
or U2938 (N_2938,N_2906,N_2872);
nor U2939 (N_2939,N_2855,N_2893);
and U2940 (N_2940,N_2891,N_2883);
nor U2941 (N_2941,N_2859,N_2853);
nand U2942 (N_2942,N_2863,N_2918);
or U2943 (N_2943,N_2911,N_2868);
nor U2944 (N_2944,N_2910,N_2915);
and U2945 (N_2945,N_2862,N_2887);
nor U2946 (N_2946,N_2895,N_2861);
nor U2947 (N_2947,N_2921,N_2850);
nand U2948 (N_2948,N_2852,N_2924);
and U2949 (N_2949,N_2857,N_2867);
or U2950 (N_2950,N_2909,N_2854);
or U2951 (N_2951,N_2917,N_2890);
or U2952 (N_2952,N_2884,N_2914);
nand U2953 (N_2953,N_2877,N_2875);
nor U2954 (N_2954,N_2871,N_2907);
and U2955 (N_2955,N_2901,N_2876);
nor U2956 (N_2956,N_2880,N_2903);
and U2957 (N_2957,N_2905,N_2892);
nand U2958 (N_2958,N_2908,N_2897);
and U2959 (N_2959,N_2866,N_2865);
nor U2960 (N_2960,N_2913,N_2919);
nand U2961 (N_2961,N_2920,N_2916);
nand U2962 (N_2962,N_2889,N_2856);
and U2963 (N_2963,N_2889,N_2920);
or U2964 (N_2964,N_2897,N_2864);
nand U2965 (N_2965,N_2890,N_2853);
and U2966 (N_2966,N_2872,N_2905);
nand U2967 (N_2967,N_2886,N_2858);
nand U2968 (N_2968,N_2909,N_2860);
nor U2969 (N_2969,N_2861,N_2875);
nor U2970 (N_2970,N_2867,N_2884);
or U2971 (N_2971,N_2912,N_2866);
nand U2972 (N_2972,N_2911,N_2881);
xnor U2973 (N_2973,N_2881,N_2918);
nand U2974 (N_2974,N_2898,N_2856);
nand U2975 (N_2975,N_2856,N_2899);
nor U2976 (N_2976,N_2869,N_2901);
nand U2977 (N_2977,N_2867,N_2862);
nor U2978 (N_2978,N_2881,N_2863);
or U2979 (N_2979,N_2905,N_2887);
or U2980 (N_2980,N_2878,N_2897);
nand U2981 (N_2981,N_2893,N_2882);
nand U2982 (N_2982,N_2878,N_2913);
and U2983 (N_2983,N_2922,N_2893);
nor U2984 (N_2984,N_2870,N_2890);
nand U2985 (N_2985,N_2919,N_2883);
or U2986 (N_2986,N_2854,N_2877);
nand U2987 (N_2987,N_2897,N_2895);
xor U2988 (N_2988,N_2886,N_2857);
and U2989 (N_2989,N_2919,N_2877);
and U2990 (N_2990,N_2920,N_2865);
nor U2991 (N_2991,N_2850,N_2867);
or U2992 (N_2992,N_2892,N_2924);
nor U2993 (N_2993,N_2910,N_2857);
nand U2994 (N_2994,N_2921,N_2851);
or U2995 (N_2995,N_2912,N_2852);
nand U2996 (N_2996,N_2850,N_2896);
nor U2997 (N_2997,N_2903,N_2874);
nor U2998 (N_2998,N_2924,N_2858);
and U2999 (N_2999,N_2897,N_2910);
nor UO_0 (O_0,N_2973,N_2986);
nor UO_1 (O_1,N_2985,N_2960);
nand UO_2 (O_2,N_2941,N_2980);
nor UO_3 (O_3,N_2938,N_2975);
nand UO_4 (O_4,N_2997,N_2961);
nand UO_5 (O_5,N_2929,N_2995);
nor UO_6 (O_6,N_2996,N_2981);
nor UO_7 (O_7,N_2943,N_2952);
or UO_8 (O_8,N_2939,N_2984);
or UO_9 (O_9,N_2954,N_2987);
or UO_10 (O_10,N_2971,N_2951);
nor UO_11 (O_11,N_2927,N_2982);
nand UO_12 (O_12,N_2963,N_2949);
nand UO_13 (O_13,N_2959,N_2940);
nor UO_14 (O_14,N_2978,N_2999);
or UO_15 (O_15,N_2931,N_2957);
nor UO_16 (O_16,N_2947,N_2958);
and UO_17 (O_17,N_2993,N_2983);
nor UO_18 (O_18,N_2990,N_2962);
and UO_19 (O_19,N_2968,N_2956);
nor UO_20 (O_20,N_2944,N_2969);
nor UO_21 (O_21,N_2942,N_2972);
nor UO_22 (O_22,N_2928,N_2964);
nor UO_23 (O_23,N_2953,N_2967);
nor UO_24 (O_24,N_2955,N_2970);
or UO_25 (O_25,N_2934,N_2988);
and UO_26 (O_26,N_2976,N_2925);
or UO_27 (O_27,N_2979,N_2992);
and UO_28 (O_28,N_2977,N_2965);
nor UO_29 (O_29,N_2932,N_2930);
or UO_30 (O_30,N_2948,N_2966);
nor UO_31 (O_31,N_2998,N_2974);
and UO_32 (O_32,N_2936,N_2933);
or UO_33 (O_33,N_2994,N_2991);
and UO_34 (O_34,N_2946,N_2935);
and UO_35 (O_35,N_2937,N_2950);
or UO_36 (O_36,N_2945,N_2989);
nand UO_37 (O_37,N_2926,N_2945);
nand UO_38 (O_38,N_2969,N_2997);
and UO_39 (O_39,N_2997,N_2973);
and UO_40 (O_40,N_2996,N_2980);
nand UO_41 (O_41,N_2992,N_2989);
nor UO_42 (O_42,N_2955,N_2969);
nor UO_43 (O_43,N_2958,N_2991);
and UO_44 (O_44,N_2945,N_2960);
or UO_45 (O_45,N_2950,N_2972);
or UO_46 (O_46,N_2930,N_2985);
nand UO_47 (O_47,N_2949,N_2929);
or UO_48 (O_48,N_2993,N_2928);
and UO_49 (O_49,N_2929,N_2933);
nand UO_50 (O_50,N_2980,N_2973);
or UO_51 (O_51,N_2974,N_2958);
and UO_52 (O_52,N_2982,N_2947);
or UO_53 (O_53,N_2976,N_2966);
nor UO_54 (O_54,N_2927,N_2964);
and UO_55 (O_55,N_2925,N_2994);
or UO_56 (O_56,N_2980,N_2969);
nor UO_57 (O_57,N_2994,N_2993);
or UO_58 (O_58,N_2933,N_2996);
nand UO_59 (O_59,N_2977,N_2979);
nor UO_60 (O_60,N_2983,N_2955);
nor UO_61 (O_61,N_2933,N_2950);
and UO_62 (O_62,N_2952,N_2973);
nor UO_63 (O_63,N_2970,N_2977);
nor UO_64 (O_64,N_2937,N_2945);
xor UO_65 (O_65,N_2970,N_2950);
or UO_66 (O_66,N_2926,N_2955);
nor UO_67 (O_67,N_2942,N_2943);
nor UO_68 (O_68,N_2933,N_2935);
or UO_69 (O_69,N_2951,N_2972);
and UO_70 (O_70,N_2953,N_2988);
nor UO_71 (O_71,N_2950,N_2941);
nand UO_72 (O_72,N_2961,N_2982);
nor UO_73 (O_73,N_2956,N_2941);
nor UO_74 (O_74,N_2954,N_2970);
or UO_75 (O_75,N_2997,N_2947);
and UO_76 (O_76,N_2959,N_2989);
nor UO_77 (O_77,N_2936,N_2938);
and UO_78 (O_78,N_2936,N_2989);
nand UO_79 (O_79,N_2941,N_2932);
or UO_80 (O_80,N_2975,N_2981);
nand UO_81 (O_81,N_2949,N_2948);
nor UO_82 (O_82,N_2992,N_2986);
nand UO_83 (O_83,N_2992,N_2972);
or UO_84 (O_84,N_2997,N_2938);
or UO_85 (O_85,N_2941,N_2975);
and UO_86 (O_86,N_2927,N_2933);
nor UO_87 (O_87,N_2934,N_2998);
xor UO_88 (O_88,N_2973,N_2994);
or UO_89 (O_89,N_2957,N_2999);
nor UO_90 (O_90,N_2963,N_2946);
nand UO_91 (O_91,N_2982,N_2925);
nand UO_92 (O_92,N_2979,N_2952);
nor UO_93 (O_93,N_2929,N_2957);
nor UO_94 (O_94,N_2973,N_2970);
or UO_95 (O_95,N_2937,N_2953);
and UO_96 (O_96,N_2987,N_2931);
nor UO_97 (O_97,N_2960,N_2993);
nor UO_98 (O_98,N_2952,N_2991);
xor UO_99 (O_99,N_2957,N_2958);
and UO_100 (O_100,N_2991,N_2941);
nand UO_101 (O_101,N_2957,N_2941);
nand UO_102 (O_102,N_2987,N_2934);
or UO_103 (O_103,N_2968,N_2970);
nand UO_104 (O_104,N_2925,N_2943);
or UO_105 (O_105,N_2974,N_2955);
nand UO_106 (O_106,N_2994,N_2946);
and UO_107 (O_107,N_2985,N_2978);
or UO_108 (O_108,N_2939,N_2998);
nor UO_109 (O_109,N_2955,N_2989);
and UO_110 (O_110,N_2953,N_2929);
nor UO_111 (O_111,N_2948,N_2994);
nand UO_112 (O_112,N_2988,N_2940);
and UO_113 (O_113,N_2929,N_2966);
or UO_114 (O_114,N_2998,N_2930);
or UO_115 (O_115,N_2955,N_2931);
nand UO_116 (O_116,N_2962,N_2963);
and UO_117 (O_117,N_2998,N_2989);
nor UO_118 (O_118,N_2951,N_2926);
nor UO_119 (O_119,N_2979,N_2968);
or UO_120 (O_120,N_2931,N_2990);
and UO_121 (O_121,N_2988,N_2941);
nand UO_122 (O_122,N_2959,N_2946);
nor UO_123 (O_123,N_2993,N_2967);
or UO_124 (O_124,N_2933,N_2969);
nand UO_125 (O_125,N_2947,N_2936);
or UO_126 (O_126,N_2984,N_2963);
and UO_127 (O_127,N_2996,N_2998);
nand UO_128 (O_128,N_2963,N_2985);
nand UO_129 (O_129,N_2992,N_2928);
nor UO_130 (O_130,N_2975,N_2930);
nor UO_131 (O_131,N_2935,N_2972);
and UO_132 (O_132,N_2929,N_2990);
or UO_133 (O_133,N_2996,N_2968);
nand UO_134 (O_134,N_2966,N_2928);
nor UO_135 (O_135,N_2945,N_2938);
nor UO_136 (O_136,N_2953,N_2948);
nor UO_137 (O_137,N_2958,N_2970);
nor UO_138 (O_138,N_2990,N_2954);
and UO_139 (O_139,N_2969,N_2952);
nor UO_140 (O_140,N_2987,N_2974);
nand UO_141 (O_141,N_2961,N_2929);
nor UO_142 (O_142,N_2960,N_2975);
nand UO_143 (O_143,N_2935,N_2950);
and UO_144 (O_144,N_2975,N_2979);
nor UO_145 (O_145,N_2996,N_2970);
and UO_146 (O_146,N_2945,N_2942);
and UO_147 (O_147,N_2999,N_2933);
or UO_148 (O_148,N_2980,N_2926);
and UO_149 (O_149,N_2946,N_2948);
nand UO_150 (O_150,N_2945,N_2946);
nor UO_151 (O_151,N_2973,N_2935);
nand UO_152 (O_152,N_2928,N_2937);
or UO_153 (O_153,N_2973,N_2927);
nor UO_154 (O_154,N_2947,N_2978);
nand UO_155 (O_155,N_2950,N_2994);
nor UO_156 (O_156,N_2969,N_2943);
nand UO_157 (O_157,N_2981,N_2943);
or UO_158 (O_158,N_2999,N_2965);
or UO_159 (O_159,N_2973,N_2962);
nor UO_160 (O_160,N_2945,N_2982);
nand UO_161 (O_161,N_2994,N_2971);
or UO_162 (O_162,N_2975,N_2937);
nand UO_163 (O_163,N_2940,N_2946);
nand UO_164 (O_164,N_2941,N_2928);
nor UO_165 (O_165,N_2962,N_2975);
nand UO_166 (O_166,N_2985,N_2936);
and UO_167 (O_167,N_2970,N_2964);
and UO_168 (O_168,N_2973,N_2940);
or UO_169 (O_169,N_2987,N_2978);
and UO_170 (O_170,N_2979,N_2934);
nor UO_171 (O_171,N_2949,N_2961);
nor UO_172 (O_172,N_2992,N_2935);
nand UO_173 (O_173,N_2958,N_2960);
and UO_174 (O_174,N_2998,N_2957);
and UO_175 (O_175,N_2985,N_2927);
nand UO_176 (O_176,N_2967,N_2958);
nand UO_177 (O_177,N_2955,N_2957);
or UO_178 (O_178,N_2975,N_2968);
and UO_179 (O_179,N_2980,N_2938);
nor UO_180 (O_180,N_2949,N_2930);
nor UO_181 (O_181,N_2926,N_2993);
or UO_182 (O_182,N_2974,N_2954);
nor UO_183 (O_183,N_2989,N_2928);
and UO_184 (O_184,N_2934,N_2931);
nor UO_185 (O_185,N_2993,N_2966);
nor UO_186 (O_186,N_2965,N_2968);
or UO_187 (O_187,N_2970,N_2928);
and UO_188 (O_188,N_2989,N_2991);
and UO_189 (O_189,N_2948,N_2969);
or UO_190 (O_190,N_2943,N_2982);
or UO_191 (O_191,N_2970,N_2961);
and UO_192 (O_192,N_2961,N_2995);
or UO_193 (O_193,N_2929,N_2940);
nor UO_194 (O_194,N_2958,N_2989);
nand UO_195 (O_195,N_2967,N_2980);
xor UO_196 (O_196,N_2966,N_2957);
xor UO_197 (O_197,N_2967,N_2974);
and UO_198 (O_198,N_2989,N_2954);
and UO_199 (O_199,N_2995,N_2936);
nor UO_200 (O_200,N_2943,N_2976);
nand UO_201 (O_201,N_2930,N_2957);
nor UO_202 (O_202,N_2936,N_2939);
nor UO_203 (O_203,N_2928,N_2945);
or UO_204 (O_204,N_2931,N_2977);
xor UO_205 (O_205,N_2945,N_2994);
nand UO_206 (O_206,N_2950,N_2969);
and UO_207 (O_207,N_2992,N_2991);
or UO_208 (O_208,N_2948,N_2957);
nor UO_209 (O_209,N_2940,N_2960);
nor UO_210 (O_210,N_2944,N_2947);
nand UO_211 (O_211,N_2958,N_2944);
or UO_212 (O_212,N_2928,N_2962);
nor UO_213 (O_213,N_2928,N_2996);
nor UO_214 (O_214,N_2982,N_2972);
nor UO_215 (O_215,N_2950,N_2962);
nand UO_216 (O_216,N_2950,N_2957);
nand UO_217 (O_217,N_2950,N_2985);
nor UO_218 (O_218,N_2989,N_2988);
or UO_219 (O_219,N_2938,N_2951);
or UO_220 (O_220,N_2983,N_2959);
nand UO_221 (O_221,N_2991,N_2956);
nor UO_222 (O_222,N_2957,N_2937);
or UO_223 (O_223,N_2976,N_2948);
nand UO_224 (O_224,N_2976,N_2947);
or UO_225 (O_225,N_2972,N_2934);
nor UO_226 (O_226,N_2952,N_2996);
and UO_227 (O_227,N_2981,N_2955);
and UO_228 (O_228,N_2977,N_2937);
and UO_229 (O_229,N_2961,N_2973);
nor UO_230 (O_230,N_2943,N_2961);
nand UO_231 (O_231,N_2963,N_2978);
or UO_232 (O_232,N_2937,N_2996);
and UO_233 (O_233,N_2935,N_2947);
or UO_234 (O_234,N_2979,N_2996);
and UO_235 (O_235,N_2969,N_2960);
or UO_236 (O_236,N_2947,N_2991);
nand UO_237 (O_237,N_2959,N_2969);
nand UO_238 (O_238,N_2945,N_2949);
nor UO_239 (O_239,N_2962,N_2992);
nand UO_240 (O_240,N_2971,N_2925);
nor UO_241 (O_241,N_2975,N_2949);
and UO_242 (O_242,N_2943,N_2958);
or UO_243 (O_243,N_2973,N_2950);
and UO_244 (O_244,N_2977,N_2957);
or UO_245 (O_245,N_2980,N_2940);
nor UO_246 (O_246,N_2939,N_2972);
nor UO_247 (O_247,N_2933,N_2932);
or UO_248 (O_248,N_2931,N_2952);
and UO_249 (O_249,N_2952,N_2939);
nor UO_250 (O_250,N_2932,N_2991);
and UO_251 (O_251,N_2930,N_2971);
and UO_252 (O_252,N_2973,N_2933);
and UO_253 (O_253,N_2989,N_2993);
or UO_254 (O_254,N_2977,N_2978);
nor UO_255 (O_255,N_2934,N_2996);
or UO_256 (O_256,N_2951,N_2963);
nor UO_257 (O_257,N_2927,N_2974);
or UO_258 (O_258,N_2992,N_2950);
nand UO_259 (O_259,N_2963,N_2993);
nor UO_260 (O_260,N_2977,N_2938);
or UO_261 (O_261,N_2927,N_2984);
nor UO_262 (O_262,N_2953,N_2993);
nand UO_263 (O_263,N_2958,N_2955);
or UO_264 (O_264,N_2995,N_2964);
or UO_265 (O_265,N_2979,N_2963);
or UO_266 (O_266,N_2951,N_2989);
and UO_267 (O_267,N_2992,N_2954);
nand UO_268 (O_268,N_2982,N_2967);
and UO_269 (O_269,N_2945,N_2985);
nand UO_270 (O_270,N_2994,N_2979);
nor UO_271 (O_271,N_2982,N_2987);
and UO_272 (O_272,N_2925,N_2929);
nor UO_273 (O_273,N_2929,N_2944);
nand UO_274 (O_274,N_2927,N_2966);
nand UO_275 (O_275,N_2991,N_2987);
nand UO_276 (O_276,N_2926,N_2943);
or UO_277 (O_277,N_2990,N_2935);
nor UO_278 (O_278,N_2989,N_2948);
and UO_279 (O_279,N_2998,N_2973);
nor UO_280 (O_280,N_2967,N_2946);
nor UO_281 (O_281,N_2979,N_2997);
or UO_282 (O_282,N_2992,N_2949);
or UO_283 (O_283,N_2955,N_2954);
or UO_284 (O_284,N_2942,N_2926);
nand UO_285 (O_285,N_2990,N_2956);
nand UO_286 (O_286,N_2964,N_2960);
nand UO_287 (O_287,N_2926,N_2944);
nand UO_288 (O_288,N_2979,N_2954);
nand UO_289 (O_289,N_2987,N_2933);
nand UO_290 (O_290,N_2981,N_2946);
or UO_291 (O_291,N_2980,N_2971);
nand UO_292 (O_292,N_2992,N_2975);
nand UO_293 (O_293,N_2928,N_2934);
and UO_294 (O_294,N_2955,N_2998);
and UO_295 (O_295,N_2991,N_2930);
nor UO_296 (O_296,N_2985,N_2977);
or UO_297 (O_297,N_2982,N_2979);
and UO_298 (O_298,N_2965,N_2930);
and UO_299 (O_299,N_2925,N_2964);
and UO_300 (O_300,N_2974,N_2945);
or UO_301 (O_301,N_2996,N_2950);
and UO_302 (O_302,N_2988,N_2927);
and UO_303 (O_303,N_2969,N_2928);
or UO_304 (O_304,N_2975,N_2931);
and UO_305 (O_305,N_2999,N_2937);
nor UO_306 (O_306,N_2997,N_2928);
nand UO_307 (O_307,N_2966,N_2988);
or UO_308 (O_308,N_2990,N_2998);
or UO_309 (O_309,N_2986,N_2929);
nand UO_310 (O_310,N_2993,N_2988);
and UO_311 (O_311,N_2953,N_2961);
nor UO_312 (O_312,N_2972,N_2929);
xor UO_313 (O_313,N_2999,N_2993);
and UO_314 (O_314,N_2956,N_2982);
nor UO_315 (O_315,N_2947,N_2948);
nand UO_316 (O_316,N_2940,N_2991);
or UO_317 (O_317,N_2946,N_2987);
or UO_318 (O_318,N_2938,N_2932);
nor UO_319 (O_319,N_2960,N_2989);
or UO_320 (O_320,N_2961,N_2989);
nor UO_321 (O_321,N_2969,N_2988);
or UO_322 (O_322,N_2968,N_2949);
xor UO_323 (O_323,N_2984,N_2962);
nand UO_324 (O_324,N_2942,N_2932);
nor UO_325 (O_325,N_2925,N_2992);
and UO_326 (O_326,N_2980,N_2939);
nand UO_327 (O_327,N_2937,N_2954);
or UO_328 (O_328,N_2990,N_2993);
nand UO_329 (O_329,N_2953,N_2925);
nor UO_330 (O_330,N_2974,N_2971);
nand UO_331 (O_331,N_2939,N_2944);
xor UO_332 (O_332,N_2932,N_2925);
or UO_333 (O_333,N_2944,N_2953);
nor UO_334 (O_334,N_2938,N_2978);
or UO_335 (O_335,N_2933,N_2960);
nor UO_336 (O_336,N_2986,N_2963);
and UO_337 (O_337,N_2942,N_2989);
nand UO_338 (O_338,N_2928,N_2952);
and UO_339 (O_339,N_2980,N_2952);
nand UO_340 (O_340,N_2951,N_2925);
or UO_341 (O_341,N_2985,N_2991);
nand UO_342 (O_342,N_2981,N_2971);
and UO_343 (O_343,N_2956,N_2997);
and UO_344 (O_344,N_2950,N_2965);
and UO_345 (O_345,N_2997,N_2945);
or UO_346 (O_346,N_2972,N_2966);
or UO_347 (O_347,N_2974,N_2943);
or UO_348 (O_348,N_2960,N_2943);
or UO_349 (O_349,N_2993,N_2951);
nand UO_350 (O_350,N_2983,N_2989);
nand UO_351 (O_351,N_2978,N_2956);
nand UO_352 (O_352,N_2981,N_2968);
nor UO_353 (O_353,N_2966,N_2973);
and UO_354 (O_354,N_2965,N_2945);
or UO_355 (O_355,N_2986,N_2939);
and UO_356 (O_356,N_2952,N_2998);
and UO_357 (O_357,N_2968,N_2953);
and UO_358 (O_358,N_2939,N_2958);
nor UO_359 (O_359,N_2983,N_2940);
nand UO_360 (O_360,N_2926,N_2970);
nand UO_361 (O_361,N_2971,N_2967);
nand UO_362 (O_362,N_2988,N_2929);
and UO_363 (O_363,N_2963,N_2954);
or UO_364 (O_364,N_2994,N_2953);
nor UO_365 (O_365,N_2994,N_2944);
or UO_366 (O_366,N_2978,N_2986);
nand UO_367 (O_367,N_2960,N_2944);
or UO_368 (O_368,N_2989,N_2934);
or UO_369 (O_369,N_2932,N_2974);
nor UO_370 (O_370,N_2944,N_2981);
nand UO_371 (O_371,N_2964,N_2965);
nand UO_372 (O_372,N_2976,N_2959);
and UO_373 (O_373,N_2963,N_2967);
nor UO_374 (O_374,N_2960,N_2996);
nand UO_375 (O_375,N_2962,N_2927);
nand UO_376 (O_376,N_2929,N_2962);
and UO_377 (O_377,N_2981,N_2939);
nor UO_378 (O_378,N_2968,N_2987);
xor UO_379 (O_379,N_2951,N_2964);
nand UO_380 (O_380,N_2994,N_2977);
nand UO_381 (O_381,N_2961,N_2993);
or UO_382 (O_382,N_2998,N_2967);
nand UO_383 (O_383,N_2989,N_2963);
and UO_384 (O_384,N_2957,N_2933);
nand UO_385 (O_385,N_2965,N_2959);
nor UO_386 (O_386,N_2969,N_2936);
and UO_387 (O_387,N_2990,N_2983);
or UO_388 (O_388,N_2934,N_2927);
nand UO_389 (O_389,N_2969,N_2949);
and UO_390 (O_390,N_2930,N_2942);
or UO_391 (O_391,N_2986,N_2935);
or UO_392 (O_392,N_2996,N_2965);
nand UO_393 (O_393,N_2972,N_2990);
or UO_394 (O_394,N_2954,N_2936);
or UO_395 (O_395,N_2988,N_2962);
nand UO_396 (O_396,N_2993,N_2935);
nand UO_397 (O_397,N_2984,N_2969);
nand UO_398 (O_398,N_2936,N_2940);
nand UO_399 (O_399,N_2974,N_2976);
or UO_400 (O_400,N_2952,N_2963);
nor UO_401 (O_401,N_2925,N_2997);
nand UO_402 (O_402,N_2934,N_2948);
xor UO_403 (O_403,N_2977,N_2999);
nand UO_404 (O_404,N_2962,N_2949);
and UO_405 (O_405,N_2983,N_2999);
nor UO_406 (O_406,N_2941,N_2951);
nor UO_407 (O_407,N_2981,N_2945);
nor UO_408 (O_408,N_2963,N_2928);
nand UO_409 (O_409,N_2952,N_2961);
nand UO_410 (O_410,N_2973,N_2981);
nor UO_411 (O_411,N_2993,N_2945);
nor UO_412 (O_412,N_2948,N_2962);
nor UO_413 (O_413,N_2944,N_2990);
or UO_414 (O_414,N_2994,N_2930);
or UO_415 (O_415,N_2957,N_2938);
nand UO_416 (O_416,N_2964,N_2963);
or UO_417 (O_417,N_2941,N_2949);
nor UO_418 (O_418,N_2983,N_2977);
or UO_419 (O_419,N_2947,N_2995);
and UO_420 (O_420,N_2951,N_2956);
and UO_421 (O_421,N_2964,N_2987);
nor UO_422 (O_422,N_2943,N_2956);
or UO_423 (O_423,N_2930,N_2952);
nand UO_424 (O_424,N_2972,N_2936);
or UO_425 (O_425,N_2957,N_2952);
nand UO_426 (O_426,N_2948,N_2932);
and UO_427 (O_427,N_2930,N_2943);
and UO_428 (O_428,N_2984,N_2973);
or UO_429 (O_429,N_2949,N_2967);
nor UO_430 (O_430,N_2928,N_2979);
xnor UO_431 (O_431,N_2950,N_2999);
nor UO_432 (O_432,N_2946,N_2936);
or UO_433 (O_433,N_2981,N_2947);
nand UO_434 (O_434,N_2934,N_2926);
and UO_435 (O_435,N_2990,N_2964);
nand UO_436 (O_436,N_2983,N_2986);
nor UO_437 (O_437,N_2997,N_2958);
xnor UO_438 (O_438,N_2995,N_2993);
and UO_439 (O_439,N_2994,N_2939);
nand UO_440 (O_440,N_2954,N_2981);
nor UO_441 (O_441,N_2962,N_2981);
or UO_442 (O_442,N_2974,N_2936);
or UO_443 (O_443,N_2981,N_2929);
or UO_444 (O_444,N_2996,N_2987);
or UO_445 (O_445,N_2989,N_2935);
or UO_446 (O_446,N_2951,N_2987);
nand UO_447 (O_447,N_2972,N_2969);
or UO_448 (O_448,N_2947,N_2951);
or UO_449 (O_449,N_2977,N_2929);
or UO_450 (O_450,N_2970,N_2972);
nor UO_451 (O_451,N_2986,N_2988);
nand UO_452 (O_452,N_2980,N_2990);
and UO_453 (O_453,N_2979,N_2981);
or UO_454 (O_454,N_2944,N_2982);
or UO_455 (O_455,N_2929,N_2950);
or UO_456 (O_456,N_2951,N_2952);
and UO_457 (O_457,N_2960,N_2931);
and UO_458 (O_458,N_2997,N_2986);
nand UO_459 (O_459,N_2958,N_2979);
nand UO_460 (O_460,N_2998,N_2977);
or UO_461 (O_461,N_2985,N_2962);
or UO_462 (O_462,N_2954,N_2929);
and UO_463 (O_463,N_2985,N_2972);
or UO_464 (O_464,N_2953,N_2992);
and UO_465 (O_465,N_2938,N_2965);
nor UO_466 (O_466,N_2971,N_2988);
and UO_467 (O_467,N_2952,N_2999);
or UO_468 (O_468,N_2943,N_2955);
nor UO_469 (O_469,N_2941,N_2994);
nand UO_470 (O_470,N_2975,N_2945);
and UO_471 (O_471,N_2974,N_2934);
nor UO_472 (O_472,N_2943,N_2991);
or UO_473 (O_473,N_2928,N_2951);
nor UO_474 (O_474,N_2987,N_2989);
nand UO_475 (O_475,N_2979,N_2998);
nand UO_476 (O_476,N_2962,N_2968);
or UO_477 (O_477,N_2974,N_2986);
nand UO_478 (O_478,N_2939,N_2991);
and UO_479 (O_479,N_2987,N_2949);
nor UO_480 (O_480,N_2994,N_2996);
nand UO_481 (O_481,N_2940,N_2927);
or UO_482 (O_482,N_2971,N_2950);
and UO_483 (O_483,N_2981,N_2966);
nand UO_484 (O_484,N_2947,N_2937);
and UO_485 (O_485,N_2989,N_2997);
and UO_486 (O_486,N_2945,N_2958);
nor UO_487 (O_487,N_2933,N_2939);
and UO_488 (O_488,N_2926,N_2995);
and UO_489 (O_489,N_2976,N_2993);
or UO_490 (O_490,N_2959,N_2927);
and UO_491 (O_491,N_2931,N_2966);
and UO_492 (O_492,N_2943,N_2940);
and UO_493 (O_493,N_2934,N_2933);
and UO_494 (O_494,N_2968,N_2995);
and UO_495 (O_495,N_2941,N_2938);
nand UO_496 (O_496,N_2977,N_2988);
nand UO_497 (O_497,N_2944,N_2936);
or UO_498 (O_498,N_2952,N_2949);
nor UO_499 (O_499,N_2929,N_2942);
endmodule