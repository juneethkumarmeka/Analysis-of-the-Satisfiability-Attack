module basic_1000_10000_1500_100_levels_10xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
nor U0 (N_0,In_655,In_437);
or U1 (N_1,In_218,In_408);
xor U2 (N_2,In_866,In_485);
nand U3 (N_3,In_449,In_644);
and U4 (N_4,In_529,In_468);
xnor U5 (N_5,In_349,In_877);
nor U6 (N_6,In_616,In_682);
or U7 (N_7,In_500,In_808);
xor U8 (N_8,In_994,In_499);
and U9 (N_9,In_951,In_634);
or U10 (N_10,In_27,In_62);
or U11 (N_11,In_947,In_691);
nor U12 (N_12,In_671,In_872);
xnor U13 (N_13,In_942,In_127);
nor U14 (N_14,In_102,In_716);
and U15 (N_15,In_64,In_521);
xor U16 (N_16,In_900,In_628);
and U17 (N_17,In_657,In_514);
nor U18 (N_18,In_411,In_4);
and U19 (N_19,In_472,In_201);
or U20 (N_20,In_256,In_15);
or U21 (N_21,In_280,In_344);
nand U22 (N_22,In_572,In_950);
or U23 (N_23,In_934,In_342);
nand U24 (N_24,In_215,In_152);
nand U25 (N_25,In_121,In_314);
nor U26 (N_26,In_621,In_43);
nand U27 (N_27,In_549,In_176);
and U28 (N_28,In_86,In_452);
nor U29 (N_29,In_260,In_10);
nand U30 (N_30,In_662,In_337);
and U31 (N_31,In_690,In_137);
and U32 (N_32,In_696,In_922);
and U33 (N_33,In_123,In_713);
nor U34 (N_34,In_269,In_124);
nand U35 (N_35,In_298,In_835);
nor U36 (N_36,In_493,In_492);
nor U37 (N_37,In_421,In_371);
and U38 (N_38,In_573,In_462);
nand U39 (N_39,In_415,In_223);
xnor U40 (N_40,In_322,In_802);
and U41 (N_41,In_561,In_976);
and U42 (N_42,In_860,In_667);
and U43 (N_43,In_839,In_692);
or U44 (N_44,In_724,In_455);
nor U45 (N_45,In_685,In_520);
xor U46 (N_46,In_425,In_585);
or U47 (N_47,In_620,In_166);
or U48 (N_48,In_974,In_413);
and U49 (N_49,In_547,In_801);
and U50 (N_50,In_525,In_285);
nor U51 (N_51,In_35,In_991);
nand U52 (N_52,In_210,In_790);
nor U53 (N_53,In_300,In_388);
and U54 (N_54,In_639,In_770);
nor U55 (N_55,In_793,In_862);
xnor U56 (N_56,In_595,In_477);
nor U57 (N_57,In_279,In_928);
nor U58 (N_58,In_737,In_308);
nor U59 (N_59,In_868,In_524);
and U60 (N_60,In_283,In_32);
xnor U61 (N_61,In_855,In_842);
xor U62 (N_62,In_214,In_483);
nand U63 (N_63,In_732,In_909);
nand U64 (N_64,In_471,In_753);
nand U65 (N_65,In_28,In_535);
nor U66 (N_66,In_112,In_828);
or U67 (N_67,In_486,In_744);
xor U68 (N_68,In_377,In_146);
and U69 (N_69,In_970,In_643);
or U70 (N_70,In_614,In_38);
nand U71 (N_71,In_911,In_319);
nor U72 (N_72,In_65,In_591);
xor U73 (N_73,In_673,In_943);
xor U74 (N_74,In_650,In_233);
and U75 (N_75,In_712,In_676);
nand U76 (N_76,In_542,In_764);
nand U77 (N_77,In_848,In_886);
and U78 (N_78,In_786,In_881);
xnor U79 (N_79,In_606,In_695);
or U80 (N_80,In_699,In_961);
nand U81 (N_81,In_783,In_661);
and U82 (N_82,In_597,In_553);
and U83 (N_83,In_904,In_754);
nor U84 (N_84,In_735,In_668);
or U85 (N_85,In_328,In_345);
nand U86 (N_86,In_659,In_321);
nand U87 (N_87,In_119,In_939);
or U88 (N_88,In_463,In_420);
and U89 (N_89,In_409,In_960);
or U90 (N_90,In_887,In_675);
or U91 (N_91,In_562,In_746);
nand U92 (N_92,In_927,In_816);
nand U93 (N_93,In_914,In_108);
nor U94 (N_94,In_265,In_326);
nand U95 (N_95,In_548,In_944);
xnor U96 (N_96,In_403,In_254);
nor U97 (N_97,In_310,In_327);
and U98 (N_98,In_434,In_892);
xnor U99 (N_99,In_987,In_821);
or U100 (N_100,In_282,In_711);
xnor U101 (N_101,In_384,In_787);
and U102 (N_102,In_966,N_71);
nand U103 (N_103,N_93,In_825);
and U104 (N_104,N_85,N_94);
and U105 (N_105,In_351,In_995);
and U106 (N_106,In_309,In_653);
nor U107 (N_107,In_580,In_334);
or U108 (N_108,In_229,In_759);
nor U109 (N_109,N_70,In_255);
or U110 (N_110,In_461,N_74);
nand U111 (N_111,In_583,In_853);
or U112 (N_112,In_350,In_154);
and U113 (N_113,In_332,N_43);
and U114 (N_114,In_743,In_507);
nand U115 (N_115,In_648,In_436);
nand U116 (N_116,In_165,In_680);
and U117 (N_117,In_83,In_728);
or U118 (N_118,In_14,In_438);
or U119 (N_119,In_479,In_523);
xor U120 (N_120,In_417,In_575);
xnor U121 (N_121,In_481,In_382);
and U122 (N_122,In_60,In_510);
or U123 (N_123,N_69,In_530);
nor U124 (N_124,In_141,In_456);
nor U125 (N_125,In_128,N_33);
xnor U126 (N_126,In_50,In_570);
nand U127 (N_127,In_103,In_160);
or U128 (N_128,In_593,In_80);
nor U129 (N_129,In_563,In_195);
and U130 (N_130,In_44,N_7);
xnor U131 (N_131,In_281,In_450);
nand U132 (N_132,In_404,In_66);
or U133 (N_133,In_819,In_244);
nand U134 (N_134,In_817,In_6);
and U135 (N_135,In_604,In_977);
and U136 (N_136,In_504,In_48);
nand U137 (N_137,In_249,N_22);
nand U138 (N_138,In_586,In_397);
or U139 (N_139,In_264,In_626);
nor U140 (N_140,In_767,N_28);
or U141 (N_141,In_227,In_320);
nand U142 (N_142,In_694,In_460);
nor U143 (N_143,In_174,In_473);
nor U144 (N_144,N_88,In_286);
and U145 (N_145,In_157,In_183);
nor U146 (N_146,In_115,N_58);
nand U147 (N_147,In_433,In_912);
and U148 (N_148,N_1,N_38);
xor U149 (N_149,In_221,In_708);
or U150 (N_150,In_815,N_8);
nand U151 (N_151,In_224,In_531);
nor U152 (N_152,In_181,In_372);
nand U153 (N_153,In_689,In_581);
nor U154 (N_154,In_278,In_142);
nor U155 (N_155,In_869,In_876);
or U156 (N_156,In_159,In_923);
and U157 (N_157,In_163,In_246);
nor U158 (N_158,In_515,In_637);
nor U159 (N_159,In_899,In_67);
xor U160 (N_160,In_739,In_932);
nor U161 (N_161,In_56,In_803);
and U162 (N_162,In_804,In_874);
xor U163 (N_163,In_807,In_954);
or U164 (N_164,In_406,In_967);
nand U165 (N_165,In_330,In_566);
or U166 (N_166,In_369,In_8);
and U167 (N_167,In_749,In_295);
and U168 (N_168,In_707,In_973);
or U169 (N_169,In_212,In_316);
nand U170 (N_170,In_182,In_550);
or U171 (N_171,N_76,In_258);
and U172 (N_172,In_543,In_715);
nor U173 (N_173,In_82,In_261);
or U174 (N_174,In_373,In_885);
and U175 (N_175,N_62,In_54);
xnor U176 (N_176,In_702,In_138);
and U177 (N_177,In_941,In_526);
nor U178 (N_178,In_164,In_870);
and U179 (N_179,In_444,In_396);
and U180 (N_180,In_379,In_688);
xor U181 (N_181,In_697,In_714);
or U182 (N_182,In_775,In_305);
or U183 (N_183,In_429,In_405);
and U184 (N_184,In_366,In_101);
xnor U185 (N_185,In_474,In_92);
nor U186 (N_186,In_601,In_883);
and U187 (N_187,In_225,In_672);
xor U188 (N_188,In_664,In_917);
nand U189 (N_189,In_70,In_552);
xor U190 (N_190,In_752,In_177);
nand U191 (N_191,In_796,In_774);
or U192 (N_192,N_2,In_447);
or U193 (N_193,In_636,In_660);
nor U194 (N_194,In_110,In_162);
xor U195 (N_195,In_454,In_567);
nor U196 (N_196,In_81,In_893);
nor U197 (N_197,In_367,In_556);
nor U198 (N_198,In_453,In_891);
nand U199 (N_199,N_29,In_841);
and U200 (N_200,In_791,In_632);
xnor U201 (N_201,In_414,In_299);
xor U202 (N_202,N_173,In_478);
xnor U203 (N_203,In_389,In_965);
and U204 (N_204,In_642,In_386);
or U205 (N_205,In_341,In_629);
nor U206 (N_206,N_80,In_107);
nand U207 (N_207,In_761,In_871);
or U208 (N_208,In_719,In_996);
or U209 (N_209,In_220,In_723);
and U210 (N_210,In_69,In_851);
nor U211 (N_211,N_198,In_41);
nand U212 (N_212,In_490,In_125);
and U213 (N_213,In_7,N_77);
nand U214 (N_214,In_998,In_703);
and U215 (N_215,N_106,In_983);
and U216 (N_216,N_79,In_969);
nand U217 (N_217,In_145,In_918);
nand U218 (N_218,In_935,N_151);
nand U219 (N_219,In_169,In_9);
nand U220 (N_220,In_925,In_262);
xnor U221 (N_221,N_9,In_494);
and U222 (N_222,In_538,N_23);
and U223 (N_223,In_779,In_230);
or U224 (N_224,In_442,N_159);
and U225 (N_225,In_859,In_518);
nor U226 (N_226,In_186,In_239);
nor U227 (N_227,In_47,In_968);
or U228 (N_228,In_370,In_380);
nand U229 (N_229,In_430,In_203);
xnor U230 (N_230,In_197,In_569);
and U231 (N_231,N_192,N_158);
nand U232 (N_232,N_135,In_226);
xnor U233 (N_233,In_68,In_532);
xnor U234 (N_234,N_175,In_778);
nor U235 (N_235,In_336,N_169);
xor U236 (N_236,In_938,In_503);
and U237 (N_237,In_199,In_780);
nor U238 (N_238,N_128,In_313);
or U239 (N_239,In_333,In_58);
nor U240 (N_240,In_762,N_30);
and U241 (N_241,In_533,In_20);
or U242 (N_242,N_5,N_60);
nor U243 (N_243,In_718,In_823);
nand U244 (N_244,In_589,N_105);
or U245 (N_245,In_559,N_87);
xnor U246 (N_246,In_989,In_958);
or U247 (N_247,In_856,In_191);
nor U248 (N_248,In_242,In_390);
nor U249 (N_249,In_439,In_211);
nand U250 (N_250,N_55,In_539);
xnor U251 (N_251,In_484,In_26);
or U252 (N_252,N_26,In_849);
nand U253 (N_253,In_505,In_475);
xnor U254 (N_254,N_82,N_162);
nor U255 (N_255,In_184,In_139);
and U256 (N_256,In_118,In_700);
nor U257 (N_257,N_152,In_179);
or U258 (N_258,N_16,In_432);
or U259 (N_259,N_91,In_480);
xnor U260 (N_260,In_957,In_832);
xnor U261 (N_261,N_103,In_104);
or U262 (N_262,In_301,In_150);
xor U263 (N_263,In_701,In_97);
or U264 (N_264,In_190,In_824);
and U265 (N_265,N_186,N_44);
nand U266 (N_266,N_10,N_63);
nor U267 (N_267,In_863,In_789);
nand U268 (N_268,N_72,In_122);
xnor U269 (N_269,In_198,N_78);
nor U270 (N_270,In_236,In_926);
nor U271 (N_271,In_564,N_117);
xor U272 (N_272,In_897,In_624);
nor U273 (N_273,N_126,N_189);
nand U274 (N_274,N_140,N_68);
or U275 (N_275,In_73,In_693);
xnor U276 (N_276,In_161,In_511);
xnor U277 (N_277,In_189,In_980);
nor U278 (N_278,In_888,In_906);
and U279 (N_279,In_440,In_206);
or U280 (N_280,In_272,In_394);
nor U281 (N_281,N_154,In_71);
nand U282 (N_282,N_65,N_143);
and U283 (N_283,In_311,In_428);
nor U284 (N_284,In_536,In_840);
or U285 (N_285,In_129,In_167);
and U286 (N_286,In_577,In_846);
and U287 (N_287,In_222,In_574);
or U288 (N_288,In_489,N_168);
or U289 (N_289,In_993,In_745);
nor U290 (N_290,In_674,In_130);
nand U291 (N_291,In_55,In_800);
xor U292 (N_292,In_259,In_677);
or U293 (N_293,N_111,In_395);
nor U294 (N_294,In_171,N_185);
or U295 (N_295,In_945,In_622);
xnor U296 (N_296,In_116,In_952);
nand U297 (N_297,In_738,In_276);
and U298 (N_298,In_908,In_940);
and U299 (N_299,In_847,In_348);
nor U300 (N_300,In_143,In_763);
nor U301 (N_301,N_209,N_132);
nor U302 (N_302,N_177,N_147);
nand U303 (N_303,N_206,In_740);
or U304 (N_304,In_376,In_464);
nor U305 (N_305,N_116,In_126);
or U306 (N_306,In_592,In_537);
xor U307 (N_307,N_59,N_190);
or U308 (N_308,In_134,N_96);
xor U309 (N_309,N_17,N_297);
nor U310 (N_310,In_173,In_470);
nor U311 (N_311,N_174,In_704);
nor U312 (N_312,In_57,N_246);
and U313 (N_313,In_458,In_865);
and U314 (N_314,In_878,In_905);
xor U315 (N_315,N_285,In_303);
nand U316 (N_316,N_12,In_245);
nand U317 (N_317,In_972,In_898);
or U318 (N_318,In_466,N_280);
or U319 (N_319,In_364,N_167);
xnor U320 (N_320,In_445,N_112);
nor U321 (N_321,In_85,In_997);
nand U322 (N_322,N_39,In_683);
and U323 (N_323,In_540,N_14);
and U324 (N_324,N_194,In_879);
xnor U325 (N_325,N_216,N_121);
and U326 (N_326,In_975,In_410);
xnor U327 (N_327,In_641,N_187);
xnor U328 (N_328,In_558,In_795);
and U329 (N_329,In_827,In_238);
nor U330 (N_330,N_281,In_231);
nand U331 (N_331,In_194,In_457);
xor U332 (N_332,In_111,N_11);
nand U333 (N_333,In_541,In_600);
and U334 (N_334,In_582,N_231);
and U335 (N_335,In_920,In_733);
or U336 (N_336,In_175,N_150);
or U337 (N_337,In_323,In_598);
nor U338 (N_338,In_826,In_810);
nor U339 (N_339,N_284,In_78);
and U340 (N_340,N_199,In_23);
nand U341 (N_341,N_250,N_272);
xnor U342 (N_342,N_273,In_751);
nor U343 (N_343,In_640,In_654);
or U344 (N_344,N_53,In_424);
and U345 (N_345,In_649,In_273);
and U346 (N_346,N_241,In_959);
or U347 (N_347,N_4,In_756);
xor U348 (N_348,In_106,In_773);
or U349 (N_349,In_284,N_97);
xor U350 (N_350,N_170,In_76);
xnor U351 (N_351,In_794,N_108);
or U352 (N_352,N_164,N_133);
xnor U353 (N_353,In_647,N_223);
and U354 (N_354,N_153,In_232);
and U355 (N_355,In_578,In_867);
or U356 (N_356,In_684,In_747);
xnor U357 (N_357,In_398,In_94);
nor U358 (N_358,In_750,In_843);
xor U359 (N_359,In_235,In_99);
or U360 (N_360,In_30,In_522);
nor U361 (N_361,N_15,In_882);
and U362 (N_362,In_978,In_208);
and U363 (N_363,N_86,In_555);
xnor U364 (N_364,In_240,In_519);
xor U365 (N_365,In_748,In_805);
or U366 (N_366,N_263,In_502);
nor U367 (N_367,In_427,In_347);
or U368 (N_368,In_39,In_512);
nor U369 (N_369,N_127,In_315);
xor U370 (N_370,In_721,N_269);
xor U371 (N_371,N_149,N_253);
nor U372 (N_372,In_401,In_557);
and U373 (N_373,N_19,In_374);
and U374 (N_374,In_187,In_607);
nor U375 (N_375,N_36,In_289);
or U376 (N_376,N_276,In_18);
nand U377 (N_377,In_33,In_652);
nor U378 (N_378,In_727,N_289);
nand U379 (N_379,In_443,In_105);
and U380 (N_380,In_267,N_100);
nand U381 (N_381,In_806,N_264);
nor U382 (N_382,N_259,In_890);
and U383 (N_383,In_257,N_122);
and U384 (N_384,In_219,In_117);
xor U385 (N_385,In_275,In_120);
or U386 (N_386,N_0,In_100);
or U387 (N_387,In_758,N_274);
xor U388 (N_388,N_224,N_283);
or U389 (N_389,In_95,In_509);
and U390 (N_390,In_98,In_469);
nor U391 (N_391,In_193,In_508);
nand U392 (N_392,N_191,In_936);
nand U393 (N_393,In_907,In_113);
nand U394 (N_394,In_709,In_335);
or U395 (N_395,N_142,In_705);
xor U396 (N_396,N_166,In_777);
and U397 (N_397,In_46,In_588);
nand U398 (N_398,In_812,In_686);
and U399 (N_399,In_418,In_213);
xor U400 (N_400,N_254,N_351);
xor U401 (N_401,N_363,In_726);
nor U402 (N_402,N_66,N_390);
nor U403 (N_403,N_300,N_326);
nand U404 (N_404,In_656,In_584);
or U405 (N_405,N_314,N_358);
xnor U406 (N_406,In_710,N_211);
or U407 (N_407,In_903,In_820);
or U408 (N_408,In_915,In_971);
nor U409 (N_409,In_953,In_990);
nand U410 (N_410,In_594,In_501);
nor U411 (N_411,In_205,N_221);
and U412 (N_412,In_185,N_155);
and U413 (N_413,N_179,N_323);
nor U414 (N_414,In_250,N_6);
or U415 (N_415,N_109,N_338);
nor U416 (N_416,In_296,In_202);
and U417 (N_417,In_192,N_136);
or U418 (N_418,N_180,N_220);
nand U419 (N_419,In_678,In_599);
and U420 (N_420,In_37,In_875);
nor U421 (N_421,In_338,N_304);
xnor U422 (N_422,N_320,In_517);
or U423 (N_423,In_916,N_244);
nand U424 (N_424,In_811,N_139);
nor U425 (N_425,N_104,N_163);
or U426 (N_426,N_378,N_342);
nor U427 (N_427,N_319,In_706);
xnor U428 (N_428,In_90,N_34);
xor U429 (N_429,In_986,N_353);
and U430 (N_430,In_665,N_25);
and U431 (N_431,In_393,In_365);
and U432 (N_432,In_534,N_379);
and U433 (N_433,In_324,N_73);
nor U434 (N_434,In_476,In_527);
and U435 (N_435,N_181,N_336);
nor U436 (N_436,N_328,N_188);
and U437 (N_437,In_331,N_102);
xnor U438 (N_438,In_772,In_623);
xor U439 (N_439,N_371,N_31);
and U440 (N_440,In_277,In_741);
xor U441 (N_441,In_19,N_200);
and U442 (N_442,In_36,In_646);
and U443 (N_443,N_235,N_396);
or U444 (N_444,N_61,N_315);
or U445 (N_445,In_237,N_373);
xor U446 (N_446,N_252,In_340);
xnor U447 (N_447,N_51,In_730);
xnor U448 (N_448,In_96,N_275);
or U449 (N_449,N_345,In_40);
xnor U450 (N_450,N_219,N_131);
and U451 (N_451,N_359,N_171);
nor U452 (N_452,N_84,In_77);
and U453 (N_453,In_769,In_12);
and U454 (N_454,In_451,N_40);
xor U455 (N_455,In_204,N_322);
or U456 (N_456,N_141,In_854);
or U457 (N_457,In_465,N_298);
nand U458 (N_458,N_341,In_554);
and U459 (N_459,N_337,In_0);
nor U460 (N_460,N_182,N_119);
nor U461 (N_461,In_615,N_307);
nand U462 (N_462,N_64,N_365);
xor U463 (N_463,N_388,N_384);
xnor U464 (N_464,In_931,N_230);
nor U465 (N_465,In_354,N_270);
xor U466 (N_466,N_387,N_389);
nor U467 (N_467,N_207,In_360);
nor U468 (N_468,N_92,N_305);
nand U469 (N_469,N_267,In_306);
xnor U470 (N_470,In_956,In_576);
xor U471 (N_471,In_217,In_830);
xnor U472 (N_472,N_13,In_516);
and U473 (N_473,N_313,N_347);
xor U474 (N_474,N_238,N_287);
nand U475 (N_475,In_156,In_5);
nand U476 (N_476,In_88,In_809);
xnor U477 (N_477,In_880,In_383);
and U478 (N_478,In_930,N_195);
nand U479 (N_479,In_979,N_213);
xor U480 (N_480,N_278,N_377);
and U481 (N_481,In_431,In_988);
or U482 (N_482,In_630,N_242);
nor U483 (N_483,In_79,N_271);
and U484 (N_484,N_137,N_308);
nand U485 (N_485,In_17,N_114);
nand U486 (N_486,In_151,In_717);
or U487 (N_487,In_981,N_145);
and U488 (N_488,In_610,N_397);
nand U489 (N_489,In_618,In_901);
or U490 (N_490,In_813,In_423);
nand U491 (N_491,In_985,In_422);
xor U492 (N_492,In_506,In_894);
nand U493 (N_493,In_91,N_236);
xor U494 (N_494,In_755,In_631);
xor U495 (N_495,In_612,N_46);
nand U496 (N_496,In_381,In_368);
nor U497 (N_497,In_31,N_89);
xnor U498 (N_498,N_214,In_625);
or U499 (N_499,In_864,In_964);
xor U500 (N_500,In_251,N_447);
nor U501 (N_501,In_613,N_258);
and U502 (N_502,N_110,In_734);
and U503 (N_503,N_393,In_209);
xnor U504 (N_504,N_203,N_432);
nand U505 (N_505,In_387,In_168);
or U506 (N_506,N_482,N_268);
and U507 (N_507,N_95,In_49);
xor U508 (N_508,N_448,N_439);
xnor U509 (N_509,In_488,N_247);
nor U510 (N_510,N_421,In_627);
or U511 (N_511,In_416,In_528);
xor U512 (N_512,N_391,N_21);
nor U513 (N_513,N_420,N_477);
or U514 (N_514,In_946,N_234);
nand U515 (N_515,In_13,N_286);
and U516 (N_516,N_303,N_459);
nand U517 (N_517,In_852,N_293);
and U518 (N_518,N_491,In_312);
nor U519 (N_519,N_57,In_579);
nor U520 (N_520,In_392,In_253);
or U521 (N_521,In_353,In_913);
xor U522 (N_522,N_407,In_148);
or U523 (N_523,In_765,N_115);
nand U524 (N_524,N_3,In_317);
and U525 (N_525,N_27,In_287);
xnor U526 (N_526,In_412,N_478);
nand U527 (N_527,In_831,N_463);
nand U528 (N_528,In_919,In_544);
nand U529 (N_529,N_118,N_291);
or U530 (N_530,N_446,N_330);
or U531 (N_531,N_437,In_963);
nand U532 (N_532,N_498,In_248);
or U533 (N_533,N_332,In_962);
and U534 (N_534,In_216,N_317);
and U535 (N_535,N_41,In_844);
xor U536 (N_536,N_277,N_457);
and U537 (N_537,In_798,N_451);
or U538 (N_538,In_788,N_488);
nand U539 (N_539,In_61,In_565);
or U540 (N_540,In_687,N_129);
and U541 (N_541,In_837,N_462);
xor U542 (N_542,N_245,N_405);
nor U543 (N_543,N_20,In_546);
or U544 (N_544,In_603,In_25);
or U545 (N_545,In_357,N_193);
xnor U546 (N_546,In_318,In_153);
nand U547 (N_547,N_324,In_133);
and U548 (N_548,N_279,In_633);
nand U549 (N_549,In_131,In_84);
and U550 (N_550,In_426,N_357);
xnor U551 (N_551,In_924,In_74);
nand U552 (N_552,In_609,In_114);
or U553 (N_553,N_292,N_366);
nor U554 (N_554,N_288,In_760);
or U555 (N_555,N_157,N_443);
xnor U556 (N_556,N_101,N_406);
or U557 (N_557,N_50,N_376);
xnor U558 (N_558,In_180,N_382);
xor U559 (N_559,N_350,N_90);
xnor U560 (N_560,N_408,N_256);
xor U561 (N_561,N_56,N_228);
or U562 (N_562,N_356,N_316);
xor U563 (N_563,N_148,N_299);
or U564 (N_564,N_239,N_339);
xnor U565 (N_565,In_22,In_75);
nand U566 (N_566,N_265,In_921);
or U567 (N_567,In_845,In_200);
nor U568 (N_568,In_63,N_434);
nand U569 (N_569,N_54,In_158);
nor U570 (N_570,N_403,N_444);
nor U571 (N_571,N_481,N_261);
and U572 (N_572,In_850,In_619);
or U573 (N_573,N_32,In_799);
nor U574 (N_574,N_81,In_937);
nand U575 (N_575,N_367,In_402);
xor U576 (N_576,N_440,N_466);
nor U577 (N_577,N_352,N_486);
nand U578 (N_578,N_372,In_784);
nand U579 (N_579,N_483,In_304);
nor U580 (N_580,N_184,In_992);
and U581 (N_581,N_346,N_210);
and U582 (N_582,In_140,N_302);
or U583 (N_583,In_266,In_290);
nand U584 (N_584,N_257,In_495);
nor U585 (N_585,In_781,N_301);
xnor U586 (N_586,N_424,In_391);
or U587 (N_587,N_475,N_321);
and U588 (N_588,N_402,In_861);
xor U589 (N_589,N_333,N_227);
nand U590 (N_590,In_933,N_479);
xnor U591 (N_591,N_496,In_596);
nand U592 (N_592,N_49,N_354);
or U593 (N_593,In_302,N_215);
and U594 (N_594,In_59,N_409);
xnor U595 (N_595,N_204,N_484);
nand U596 (N_596,In_288,N_98);
nand U597 (N_597,N_343,In_785);
nand U598 (N_598,N_52,In_838);
nand U599 (N_599,N_433,N_469);
nand U600 (N_600,N_558,In_895);
or U601 (N_601,N_455,N_426);
nor U602 (N_602,N_497,N_453);
or U603 (N_603,In_271,In_829);
nor U604 (N_604,In_234,N_465);
or U605 (N_605,N_500,N_461);
nor U606 (N_606,N_514,In_645);
or U607 (N_607,In_669,N_591);
xnor U608 (N_608,N_588,N_552);
nand U609 (N_609,N_165,In_658);
nor U610 (N_610,In_16,N_458);
nand U611 (N_611,In_797,N_492);
xnor U612 (N_612,N_553,In_949);
nor U613 (N_613,In_545,In_984);
nor U614 (N_614,N_564,In_679);
nor U615 (N_615,N_222,N_540);
xor U616 (N_616,In_834,N_593);
and U617 (N_617,N_42,N_505);
nand U618 (N_618,In_725,In_144);
nand U619 (N_619,In_11,In_722);
and U620 (N_620,N_494,N_577);
and U621 (N_621,N_161,In_307);
nand U622 (N_622,N_260,N_521);
nor U623 (N_623,N_183,N_471);
and U624 (N_624,N_306,N_233);
nor U625 (N_625,In_274,N_454);
and U626 (N_626,N_370,N_392);
or U627 (N_627,N_536,N_35);
or U628 (N_628,N_566,N_490);
xor U629 (N_629,N_107,In_513);
and U630 (N_630,N_547,In_766);
nand U631 (N_631,N_243,N_325);
and U632 (N_632,N_218,N_473);
nor U633 (N_633,In_155,In_352);
and U634 (N_634,In_419,N_18);
nand U635 (N_635,N_355,In_93);
or U636 (N_636,N_523,N_240);
xnor U637 (N_637,In_196,In_355);
and U638 (N_638,N_375,N_335);
nand U639 (N_639,N_563,N_160);
and U640 (N_640,In_884,N_551);
or U641 (N_641,In_448,In_731);
or U642 (N_642,N_232,In_42);
nand U643 (N_643,N_598,In_729);
nand U644 (N_644,In_21,In_51);
nor U645 (N_645,N_294,In_243);
and U646 (N_646,In_147,N_430);
and U647 (N_647,In_496,N_441);
or U648 (N_648,N_138,N_548);
nor U649 (N_649,N_310,N_562);
nand U650 (N_650,N_541,In_551);
and U651 (N_651,N_248,N_517);
xnor U652 (N_652,N_549,N_542);
and U653 (N_653,N_456,In_818);
xnor U654 (N_654,N_499,N_37);
xnor U655 (N_655,In_136,N_229);
xor U656 (N_656,N_450,In_329);
nor U657 (N_657,In_590,N_528);
xor U658 (N_658,N_546,N_507);
xnor U659 (N_659,In_638,N_125);
xor U660 (N_660,N_401,N_510);
xor U661 (N_661,N_334,N_196);
xor U662 (N_662,N_474,In_467);
or U663 (N_663,N_386,N_511);
nand U664 (N_664,In_399,N_597);
and U665 (N_665,N_282,N_249);
nand U666 (N_666,In_385,N_569);
or U667 (N_667,In_87,N_364);
nand U668 (N_668,N_572,N_385);
nand U669 (N_669,N_212,In_343);
or U670 (N_670,In_375,N_493);
and U671 (N_671,N_467,N_529);
nor U672 (N_672,N_197,In_948);
nor U673 (N_673,N_506,N_487);
and U674 (N_674,N_113,In_982);
xor U675 (N_675,N_208,In_172);
xor U676 (N_676,N_331,In_53);
and U677 (N_677,N_349,N_582);
or U678 (N_678,In_263,N_436);
nand U679 (N_679,In_24,N_512);
or U680 (N_680,In_635,N_587);
xnor U681 (N_681,N_568,In_910);
or U682 (N_682,In_568,In_482);
nand U683 (N_683,In_109,In_873);
or U684 (N_684,N_422,N_555);
or U685 (N_685,N_262,N_362);
xnor U686 (N_686,N_423,In_407);
xnor U687 (N_687,In_889,In_605);
or U688 (N_688,N_369,In_1);
or U689 (N_689,N_361,In_459);
and U690 (N_690,N_472,In_29);
nor U691 (N_691,N_296,In_858);
nor U692 (N_692,N_581,N_503);
nor U693 (N_693,N_83,N_554);
and U694 (N_694,In_822,N_47);
and U695 (N_695,N_445,In_720);
or U696 (N_696,N_594,N_522);
and U697 (N_697,In_768,In_441);
xor U698 (N_698,In_241,In_587);
nand U699 (N_699,N_255,N_539);
or U700 (N_700,N_67,N_266);
nand U701 (N_701,N_618,In_291);
nor U702 (N_702,N_624,N_652);
or U703 (N_703,N_476,In_247);
xor U704 (N_704,N_636,N_449);
xor U705 (N_705,N_130,N_550);
nor U706 (N_706,N_312,N_663);
nor U707 (N_707,N_578,N_610);
xor U708 (N_708,N_687,In_651);
nand U709 (N_709,N_631,N_576);
xnor U710 (N_710,N_655,N_638);
or U711 (N_711,N_516,In_560);
or U712 (N_712,N_669,N_489);
and U713 (N_713,N_668,N_646);
or U714 (N_714,N_480,N_431);
nand U715 (N_715,N_45,N_309);
nor U716 (N_716,N_605,N_590);
xnor U717 (N_717,N_659,N_621);
nand U718 (N_718,N_570,N_124);
and U719 (N_719,N_671,N_532);
and U720 (N_720,N_611,N_579);
xnor U721 (N_721,In_2,In_170);
nor U722 (N_722,In_228,N_685);
nor U723 (N_723,N_680,In_896);
nor U724 (N_724,N_635,N_344);
xor U725 (N_725,N_599,N_509);
xnor U726 (N_726,N_676,N_644);
or U727 (N_727,N_417,N_557);
xor U728 (N_728,N_205,N_664);
nand U729 (N_729,N_604,N_442);
nand U730 (N_730,In_346,N_383);
xnor U731 (N_731,N_625,In_491);
and U732 (N_732,N_156,N_360);
or U733 (N_733,N_400,N_592);
or U734 (N_734,N_318,N_75);
and U735 (N_735,N_639,N_609);
or U736 (N_736,N_689,N_574);
nor U737 (N_737,N_684,In_497);
nor U738 (N_738,In_358,N_628);
and U739 (N_739,N_595,N_535);
or U740 (N_740,N_295,N_543);
nor U741 (N_741,N_418,In_857);
or U742 (N_742,N_573,N_623);
and U743 (N_743,N_527,In_361);
xor U744 (N_744,N_620,N_533);
or U745 (N_745,N_530,N_225);
or U746 (N_746,N_584,N_633);
nand U747 (N_747,N_691,In_325);
or U748 (N_748,N_464,In_617);
xnor U749 (N_749,N_661,N_559);
nand U750 (N_750,N_368,N_134);
nand U751 (N_751,N_657,N_696);
nor U752 (N_752,N_374,In_999);
nand U753 (N_753,N_172,In_400);
and U754 (N_754,In_339,N_534);
or U755 (N_755,N_427,N_640);
xnor U756 (N_756,In_776,N_641);
nor U757 (N_757,N_580,In_178);
xnor U758 (N_758,N_525,N_470);
and U759 (N_759,N_537,N_688);
nor U760 (N_760,N_419,N_520);
nor U761 (N_761,N_99,N_538);
or U762 (N_762,N_560,In_666);
nand U763 (N_763,N_622,N_524);
or U764 (N_764,N_679,N_630);
xor U765 (N_765,N_348,In_929);
xor U766 (N_766,N_501,N_627);
nand U767 (N_767,N_226,N_606);
xnor U768 (N_768,N_690,N_460);
nand U769 (N_769,N_617,In_359);
xor U770 (N_770,In_487,N_607);
or U771 (N_771,N_485,N_602);
or U772 (N_772,N_146,In_268);
xnor U773 (N_773,N_48,In_89);
or U774 (N_774,N_697,In_698);
xnor U775 (N_775,N_653,In_72);
and U776 (N_776,N_176,N_515);
nand U777 (N_777,N_412,N_695);
nor U778 (N_778,N_632,N_544);
nor U779 (N_779,N_658,N_428);
xnor U780 (N_780,N_567,N_394);
or U781 (N_781,N_531,In_663);
nand U782 (N_782,N_178,N_616);
or U783 (N_783,N_650,In_292);
or U784 (N_784,N_411,N_201);
xnor U785 (N_785,N_589,N_656);
or U786 (N_786,In_188,In_611);
xnor U787 (N_787,N_675,N_612);
nor U788 (N_788,In_356,N_651);
nand U789 (N_789,N_678,N_575);
and U790 (N_790,N_673,N_600);
and U791 (N_791,N_629,N_416);
nand U792 (N_792,In_681,In_833);
nand U793 (N_793,N_438,N_672);
nand U794 (N_794,In_757,N_586);
nand U795 (N_795,N_217,N_290);
nand U796 (N_796,N_24,In_771);
nor U797 (N_797,N_666,N_410);
and U798 (N_798,N_649,N_381);
nor U799 (N_799,N_380,N_615);
xnor U800 (N_800,N_732,In_498);
nand U801 (N_801,N_735,N_662);
nor U802 (N_802,N_746,N_404);
or U803 (N_803,N_713,N_667);
or U804 (N_804,In_45,N_753);
and U805 (N_805,N_743,N_792);
nand U806 (N_806,N_681,N_782);
xor U807 (N_807,N_698,N_726);
xnor U808 (N_808,N_770,N_739);
nand U809 (N_809,N_761,N_413);
nand U810 (N_810,In_571,N_613);
nor U811 (N_811,N_755,N_767);
or U812 (N_812,In_149,In_135);
nor U813 (N_813,N_585,N_702);
or U814 (N_814,N_786,N_601);
and U815 (N_815,N_415,N_797);
xor U816 (N_816,In_902,N_791);
and U817 (N_817,N_395,N_683);
or U818 (N_818,N_705,In_52);
xnor U819 (N_819,In_670,N_762);
xor U820 (N_820,N_752,N_754);
xnor U821 (N_821,N_798,N_775);
and U822 (N_822,N_787,N_728);
xor U823 (N_823,N_251,N_759);
and U824 (N_824,N_495,N_565);
xor U825 (N_825,N_736,N_123);
or U826 (N_826,N_785,N_751);
nand U827 (N_827,N_704,N_508);
nand U828 (N_828,N_571,N_504);
xnor U829 (N_829,N_795,In_270);
nor U830 (N_830,N_734,N_596);
or U831 (N_831,N_778,N_729);
xor U832 (N_832,N_700,N_756);
xnor U833 (N_833,N_788,N_716);
xnor U834 (N_834,N_694,N_708);
and U835 (N_835,N_468,N_772);
nor U836 (N_836,N_769,N_398);
nand U837 (N_837,N_311,N_730);
xnor U838 (N_838,N_237,N_745);
nand U839 (N_839,N_727,N_692);
nor U840 (N_840,N_779,N_452);
nor U841 (N_841,N_794,N_518);
xnor U842 (N_842,N_686,N_502);
or U843 (N_843,N_748,In_435);
nand U844 (N_844,N_757,N_699);
and U845 (N_845,N_703,N_742);
nor U846 (N_846,N_693,N_682);
nor U847 (N_847,N_714,N_784);
and U848 (N_848,N_768,In_3);
nor U849 (N_849,N_718,In_836);
nand U850 (N_850,N_665,N_721);
nand U851 (N_851,N_771,N_747);
or U852 (N_852,N_763,N_725);
nor U853 (N_853,N_677,In_294);
xor U854 (N_854,N_707,N_647);
and U855 (N_855,N_660,N_619);
or U856 (N_856,N_429,N_719);
nand U857 (N_857,In_608,N_637);
and U858 (N_858,In_446,N_781);
and U859 (N_859,N_749,N_731);
and U860 (N_860,N_777,N_712);
nand U861 (N_861,N_733,N_720);
nand U862 (N_862,N_773,In_297);
xnor U863 (N_863,N_634,N_643);
and U864 (N_864,N_710,In_362);
xor U865 (N_865,N_513,N_723);
or U866 (N_866,N_519,In_736);
xor U867 (N_867,In_814,In_363);
xnor U868 (N_868,N_709,N_799);
xor U869 (N_869,N_202,N_796);
or U870 (N_870,N_783,N_545);
or U871 (N_871,N_760,In_782);
nor U872 (N_872,N_648,N_750);
or U873 (N_873,N_766,N_774);
and U874 (N_874,N_701,N_608);
nor U875 (N_875,In_602,N_715);
or U876 (N_876,In_742,In_792);
and U877 (N_877,N_556,N_758);
nor U878 (N_878,N_744,N_764);
xnor U879 (N_879,N_724,N_561);
or U880 (N_880,N_603,N_425);
nor U881 (N_881,In_252,N_583);
xnor U882 (N_882,N_740,N_399);
or U883 (N_883,N_717,N_526);
nand U884 (N_884,N_327,N_144);
and U885 (N_885,N_706,N_654);
nand U886 (N_886,N_790,In_293);
and U887 (N_887,N_780,N_737);
or U888 (N_888,N_626,In_207);
nand U889 (N_889,N_765,In_955);
nand U890 (N_890,N_614,N_741);
xor U891 (N_891,N_340,N_645);
nand U892 (N_892,In_34,N_776);
nor U893 (N_893,N_738,N_711);
nor U894 (N_894,In_132,N_435);
nor U895 (N_895,N_329,In_378);
or U896 (N_896,N_120,N_642);
nand U897 (N_897,N_670,N_674);
or U898 (N_898,N_789,N_722);
xnor U899 (N_899,N_414,N_793);
xnor U900 (N_900,N_839,N_889);
xnor U901 (N_901,N_878,N_812);
and U902 (N_902,N_897,N_873);
and U903 (N_903,N_838,N_823);
or U904 (N_904,N_824,N_880);
nand U905 (N_905,N_851,N_803);
or U906 (N_906,N_852,N_836);
and U907 (N_907,N_819,N_861);
or U908 (N_908,N_879,N_868);
or U909 (N_909,N_806,N_858);
nand U910 (N_910,N_869,N_863);
or U911 (N_911,N_827,N_860);
or U912 (N_912,N_887,N_804);
nor U913 (N_913,N_885,N_807);
xnor U914 (N_914,N_853,N_802);
and U915 (N_915,N_891,N_875);
nand U916 (N_916,N_888,N_817);
nor U917 (N_917,N_835,N_862);
or U918 (N_918,N_821,N_828);
xor U919 (N_919,N_884,N_811);
xor U920 (N_920,N_843,N_841);
nor U921 (N_921,N_896,N_857);
xor U922 (N_922,N_890,N_893);
xnor U923 (N_923,N_854,N_840);
xnor U924 (N_924,N_876,N_859);
or U925 (N_925,N_883,N_898);
and U926 (N_926,N_829,N_872);
xnor U927 (N_927,N_866,N_855);
or U928 (N_928,N_834,N_816);
nor U929 (N_929,N_848,N_849);
or U930 (N_930,N_886,N_895);
and U931 (N_931,N_822,N_844);
nor U932 (N_932,N_846,N_813);
or U933 (N_933,N_818,N_809);
xnor U934 (N_934,N_882,N_850);
or U935 (N_935,N_842,N_826);
and U936 (N_936,N_867,N_865);
and U937 (N_937,N_847,N_877);
nor U938 (N_938,N_864,N_845);
nor U939 (N_939,N_881,N_831);
nor U940 (N_940,N_830,N_894);
nand U941 (N_941,N_874,N_801);
nand U942 (N_942,N_856,N_832);
or U943 (N_943,N_833,N_892);
nand U944 (N_944,N_810,N_837);
nor U945 (N_945,N_808,N_870);
nand U946 (N_946,N_820,N_871);
or U947 (N_947,N_815,N_814);
or U948 (N_948,N_800,N_825);
nand U949 (N_949,N_899,N_805);
xnor U950 (N_950,N_803,N_819);
and U951 (N_951,N_844,N_827);
xor U952 (N_952,N_893,N_846);
nor U953 (N_953,N_839,N_891);
nand U954 (N_954,N_898,N_851);
nor U955 (N_955,N_889,N_872);
or U956 (N_956,N_874,N_851);
nand U957 (N_957,N_871,N_883);
nand U958 (N_958,N_875,N_817);
and U959 (N_959,N_858,N_868);
nor U960 (N_960,N_859,N_831);
nor U961 (N_961,N_894,N_813);
or U962 (N_962,N_851,N_871);
nor U963 (N_963,N_894,N_849);
xor U964 (N_964,N_890,N_894);
xor U965 (N_965,N_877,N_869);
and U966 (N_966,N_868,N_893);
xnor U967 (N_967,N_845,N_849);
nand U968 (N_968,N_818,N_806);
and U969 (N_969,N_894,N_868);
or U970 (N_970,N_877,N_894);
nor U971 (N_971,N_882,N_866);
xor U972 (N_972,N_873,N_887);
xor U973 (N_973,N_817,N_846);
nor U974 (N_974,N_807,N_835);
and U975 (N_975,N_829,N_859);
or U976 (N_976,N_809,N_845);
xor U977 (N_977,N_808,N_886);
nor U978 (N_978,N_875,N_805);
or U979 (N_979,N_824,N_804);
or U980 (N_980,N_840,N_825);
xor U981 (N_981,N_817,N_812);
and U982 (N_982,N_880,N_857);
nand U983 (N_983,N_898,N_808);
nand U984 (N_984,N_859,N_887);
xnor U985 (N_985,N_803,N_871);
or U986 (N_986,N_878,N_870);
or U987 (N_987,N_804,N_805);
nor U988 (N_988,N_805,N_845);
and U989 (N_989,N_824,N_837);
nand U990 (N_990,N_863,N_842);
nand U991 (N_991,N_866,N_836);
nor U992 (N_992,N_800,N_874);
xor U993 (N_993,N_850,N_849);
nand U994 (N_994,N_860,N_879);
nand U995 (N_995,N_816,N_820);
nor U996 (N_996,N_822,N_808);
nand U997 (N_997,N_892,N_816);
nor U998 (N_998,N_846,N_844);
xnor U999 (N_999,N_892,N_835);
xor U1000 (N_1000,N_902,N_935);
nor U1001 (N_1001,N_968,N_929);
or U1002 (N_1002,N_931,N_977);
nand U1003 (N_1003,N_966,N_982);
nand U1004 (N_1004,N_946,N_985);
xor U1005 (N_1005,N_979,N_920);
xnor U1006 (N_1006,N_911,N_932);
nand U1007 (N_1007,N_955,N_925);
nor U1008 (N_1008,N_908,N_998);
nand U1009 (N_1009,N_926,N_907);
or U1010 (N_1010,N_930,N_956);
xnor U1011 (N_1011,N_990,N_938);
nor U1012 (N_1012,N_904,N_976);
and U1013 (N_1013,N_948,N_942);
nand U1014 (N_1014,N_970,N_927);
xor U1015 (N_1015,N_958,N_959);
nand U1016 (N_1016,N_900,N_923);
and U1017 (N_1017,N_947,N_971);
nand U1018 (N_1018,N_995,N_962);
and U1019 (N_1019,N_919,N_949);
nand U1020 (N_1020,N_960,N_961);
nand U1021 (N_1021,N_967,N_980);
nand U1022 (N_1022,N_983,N_969);
xor U1023 (N_1023,N_939,N_972);
nor U1024 (N_1024,N_913,N_906);
nand U1025 (N_1025,N_975,N_934);
or U1026 (N_1026,N_963,N_915);
xor U1027 (N_1027,N_905,N_984);
and U1028 (N_1028,N_989,N_918);
and U1029 (N_1029,N_988,N_933);
nor U1030 (N_1030,N_992,N_903);
and U1031 (N_1031,N_996,N_950);
xnor U1032 (N_1032,N_936,N_922);
nand U1033 (N_1033,N_974,N_986);
or U1034 (N_1034,N_987,N_965);
and U1035 (N_1035,N_940,N_957);
nand U1036 (N_1036,N_951,N_964);
nand U1037 (N_1037,N_921,N_917);
xnor U1038 (N_1038,N_978,N_944);
and U1039 (N_1039,N_909,N_912);
nor U1040 (N_1040,N_916,N_910);
nor U1041 (N_1041,N_993,N_954);
nor U1042 (N_1042,N_999,N_994);
nand U1043 (N_1043,N_941,N_937);
and U1044 (N_1044,N_952,N_901);
and U1045 (N_1045,N_943,N_997);
xnor U1046 (N_1046,N_981,N_953);
nor U1047 (N_1047,N_924,N_914);
or U1048 (N_1048,N_945,N_991);
and U1049 (N_1049,N_928,N_973);
or U1050 (N_1050,N_938,N_904);
nor U1051 (N_1051,N_954,N_978);
xor U1052 (N_1052,N_937,N_911);
xnor U1053 (N_1053,N_978,N_951);
and U1054 (N_1054,N_959,N_953);
xor U1055 (N_1055,N_973,N_931);
xor U1056 (N_1056,N_913,N_961);
xor U1057 (N_1057,N_990,N_955);
or U1058 (N_1058,N_924,N_958);
or U1059 (N_1059,N_963,N_945);
and U1060 (N_1060,N_924,N_907);
xnor U1061 (N_1061,N_944,N_926);
xnor U1062 (N_1062,N_990,N_973);
or U1063 (N_1063,N_901,N_970);
or U1064 (N_1064,N_946,N_989);
nor U1065 (N_1065,N_918,N_967);
and U1066 (N_1066,N_947,N_985);
nor U1067 (N_1067,N_982,N_921);
or U1068 (N_1068,N_918,N_980);
or U1069 (N_1069,N_912,N_916);
and U1070 (N_1070,N_993,N_992);
and U1071 (N_1071,N_936,N_934);
and U1072 (N_1072,N_928,N_902);
or U1073 (N_1073,N_930,N_969);
nor U1074 (N_1074,N_988,N_919);
xnor U1075 (N_1075,N_933,N_937);
nand U1076 (N_1076,N_936,N_929);
xnor U1077 (N_1077,N_986,N_948);
xnor U1078 (N_1078,N_929,N_933);
and U1079 (N_1079,N_928,N_989);
nor U1080 (N_1080,N_901,N_988);
xor U1081 (N_1081,N_965,N_925);
xor U1082 (N_1082,N_984,N_943);
nor U1083 (N_1083,N_983,N_925);
nor U1084 (N_1084,N_950,N_919);
and U1085 (N_1085,N_915,N_999);
and U1086 (N_1086,N_906,N_967);
nor U1087 (N_1087,N_932,N_945);
nor U1088 (N_1088,N_942,N_913);
nand U1089 (N_1089,N_968,N_907);
or U1090 (N_1090,N_928,N_926);
nand U1091 (N_1091,N_949,N_996);
nand U1092 (N_1092,N_953,N_966);
nor U1093 (N_1093,N_910,N_923);
and U1094 (N_1094,N_939,N_915);
and U1095 (N_1095,N_960,N_913);
nor U1096 (N_1096,N_964,N_900);
nor U1097 (N_1097,N_920,N_985);
xor U1098 (N_1098,N_946,N_923);
or U1099 (N_1099,N_935,N_966);
or U1100 (N_1100,N_1026,N_1098);
xnor U1101 (N_1101,N_1047,N_1039);
xnor U1102 (N_1102,N_1037,N_1036);
xnor U1103 (N_1103,N_1029,N_1091);
or U1104 (N_1104,N_1020,N_1096);
nand U1105 (N_1105,N_1097,N_1072);
nor U1106 (N_1106,N_1068,N_1045);
and U1107 (N_1107,N_1009,N_1007);
nor U1108 (N_1108,N_1087,N_1074);
or U1109 (N_1109,N_1057,N_1006);
nor U1110 (N_1110,N_1065,N_1071);
or U1111 (N_1111,N_1076,N_1064);
or U1112 (N_1112,N_1059,N_1002);
xor U1113 (N_1113,N_1056,N_1034);
xnor U1114 (N_1114,N_1051,N_1035);
and U1115 (N_1115,N_1032,N_1080);
nor U1116 (N_1116,N_1073,N_1085);
xor U1117 (N_1117,N_1040,N_1077);
nor U1118 (N_1118,N_1003,N_1050);
and U1119 (N_1119,N_1000,N_1021);
or U1120 (N_1120,N_1054,N_1044);
xor U1121 (N_1121,N_1063,N_1022);
nor U1122 (N_1122,N_1001,N_1015);
nor U1123 (N_1123,N_1031,N_1053);
and U1124 (N_1124,N_1060,N_1083);
xor U1125 (N_1125,N_1033,N_1025);
or U1126 (N_1126,N_1090,N_1094);
and U1127 (N_1127,N_1019,N_1092);
and U1128 (N_1128,N_1046,N_1041);
xor U1129 (N_1129,N_1055,N_1093);
nand U1130 (N_1130,N_1084,N_1048);
nand U1131 (N_1131,N_1043,N_1016);
xor U1132 (N_1132,N_1049,N_1089);
nor U1133 (N_1133,N_1062,N_1067);
or U1134 (N_1134,N_1028,N_1066);
nor U1135 (N_1135,N_1012,N_1081);
and U1136 (N_1136,N_1027,N_1011);
xnor U1137 (N_1137,N_1058,N_1095);
nand U1138 (N_1138,N_1082,N_1017);
and U1139 (N_1139,N_1038,N_1075);
nand U1140 (N_1140,N_1013,N_1078);
nand U1141 (N_1141,N_1014,N_1030);
or U1142 (N_1142,N_1086,N_1052);
and U1143 (N_1143,N_1023,N_1099);
or U1144 (N_1144,N_1069,N_1004);
nand U1145 (N_1145,N_1042,N_1061);
xor U1146 (N_1146,N_1079,N_1088);
nand U1147 (N_1147,N_1008,N_1005);
nor U1148 (N_1148,N_1010,N_1070);
or U1149 (N_1149,N_1018,N_1024);
xor U1150 (N_1150,N_1019,N_1071);
nor U1151 (N_1151,N_1037,N_1052);
nand U1152 (N_1152,N_1078,N_1069);
or U1153 (N_1153,N_1063,N_1075);
nor U1154 (N_1154,N_1013,N_1076);
nand U1155 (N_1155,N_1037,N_1042);
and U1156 (N_1156,N_1059,N_1053);
and U1157 (N_1157,N_1043,N_1054);
nand U1158 (N_1158,N_1046,N_1018);
or U1159 (N_1159,N_1078,N_1004);
xnor U1160 (N_1160,N_1074,N_1019);
xor U1161 (N_1161,N_1034,N_1008);
and U1162 (N_1162,N_1004,N_1061);
nand U1163 (N_1163,N_1064,N_1019);
xnor U1164 (N_1164,N_1051,N_1039);
and U1165 (N_1165,N_1095,N_1094);
and U1166 (N_1166,N_1050,N_1020);
and U1167 (N_1167,N_1011,N_1019);
nand U1168 (N_1168,N_1019,N_1059);
xnor U1169 (N_1169,N_1009,N_1032);
or U1170 (N_1170,N_1053,N_1078);
and U1171 (N_1171,N_1054,N_1011);
and U1172 (N_1172,N_1017,N_1092);
or U1173 (N_1173,N_1010,N_1085);
xnor U1174 (N_1174,N_1003,N_1031);
and U1175 (N_1175,N_1002,N_1074);
nor U1176 (N_1176,N_1001,N_1085);
or U1177 (N_1177,N_1007,N_1042);
and U1178 (N_1178,N_1065,N_1088);
and U1179 (N_1179,N_1094,N_1045);
nand U1180 (N_1180,N_1053,N_1027);
or U1181 (N_1181,N_1055,N_1099);
nor U1182 (N_1182,N_1004,N_1067);
and U1183 (N_1183,N_1098,N_1003);
nand U1184 (N_1184,N_1037,N_1025);
nor U1185 (N_1185,N_1089,N_1040);
or U1186 (N_1186,N_1053,N_1097);
xor U1187 (N_1187,N_1033,N_1078);
nand U1188 (N_1188,N_1074,N_1049);
nor U1189 (N_1189,N_1069,N_1057);
nor U1190 (N_1190,N_1053,N_1064);
xor U1191 (N_1191,N_1086,N_1005);
xnor U1192 (N_1192,N_1059,N_1006);
xnor U1193 (N_1193,N_1070,N_1001);
nand U1194 (N_1194,N_1074,N_1070);
and U1195 (N_1195,N_1060,N_1082);
nand U1196 (N_1196,N_1071,N_1007);
nor U1197 (N_1197,N_1060,N_1039);
or U1198 (N_1198,N_1032,N_1047);
nor U1199 (N_1199,N_1017,N_1011);
xnor U1200 (N_1200,N_1101,N_1139);
and U1201 (N_1201,N_1106,N_1154);
and U1202 (N_1202,N_1193,N_1118);
nor U1203 (N_1203,N_1170,N_1115);
xnor U1204 (N_1204,N_1116,N_1132);
xor U1205 (N_1205,N_1188,N_1198);
nand U1206 (N_1206,N_1158,N_1144);
and U1207 (N_1207,N_1104,N_1180);
or U1208 (N_1208,N_1119,N_1146);
nand U1209 (N_1209,N_1124,N_1173);
nor U1210 (N_1210,N_1136,N_1159);
or U1211 (N_1211,N_1147,N_1176);
and U1212 (N_1212,N_1131,N_1164);
xnor U1213 (N_1213,N_1181,N_1126);
nor U1214 (N_1214,N_1122,N_1130);
xnor U1215 (N_1215,N_1168,N_1100);
and U1216 (N_1216,N_1184,N_1174);
xor U1217 (N_1217,N_1153,N_1121);
and U1218 (N_1218,N_1127,N_1150);
xnor U1219 (N_1219,N_1172,N_1111);
or U1220 (N_1220,N_1123,N_1149);
nand U1221 (N_1221,N_1199,N_1197);
nor U1222 (N_1222,N_1182,N_1125);
and U1223 (N_1223,N_1166,N_1129);
or U1224 (N_1224,N_1191,N_1128);
or U1225 (N_1225,N_1157,N_1108);
and U1226 (N_1226,N_1145,N_1151);
xor U1227 (N_1227,N_1163,N_1175);
nand U1228 (N_1228,N_1167,N_1156);
nand U1229 (N_1229,N_1171,N_1169);
nand U1230 (N_1230,N_1113,N_1189);
xor U1231 (N_1231,N_1196,N_1137);
nor U1232 (N_1232,N_1190,N_1138);
xor U1233 (N_1233,N_1152,N_1194);
xnor U1234 (N_1234,N_1109,N_1155);
nor U1235 (N_1235,N_1103,N_1134);
nand U1236 (N_1236,N_1140,N_1187);
nand U1237 (N_1237,N_1148,N_1160);
xor U1238 (N_1238,N_1107,N_1117);
nor U1239 (N_1239,N_1105,N_1183);
nor U1240 (N_1240,N_1112,N_1133);
nand U1241 (N_1241,N_1195,N_1135);
and U1242 (N_1242,N_1114,N_1141);
xnor U1243 (N_1243,N_1192,N_1185);
nor U1244 (N_1244,N_1179,N_1143);
nand U1245 (N_1245,N_1177,N_1162);
nor U1246 (N_1246,N_1165,N_1161);
nand U1247 (N_1247,N_1102,N_1110);
xnor U1248 (N_1248,N_1178,N_1142);
nand U1249 (N_1249,N_1120,N_1186);
and U1250 (N_1250,N_1115,N_1120);
nor U1251 (N_1251,N_1157,N_1169);
nor U1252 (N_1252,N_1132,N_1102);
and U1253 (N_1253,N_1189,N_1104);
nor U1254 (N_1254,N_1125,N_1195);
nor U1255 (N_1255,N_1137,N_1198);
xor U1256 (N_1256,N_1162,N_1124);
and U1257 (N_1257,N_1168,N_1163);
xnor U1258 (N_1258,N_1152,N_1168);
nand U1259 (N_1259,N_1109,N_1191);
xor U1260 (N_1260,N_1113,N_1136);
xor U1261 (N_1261,N_1160,N_1169);
and U1262 (N_1262,N_1119,N_1124);
nor U1263 (N_1263,N_1169,N_1161);
or U1264 (N_1264,N_1122,N_1190);
nand U1265 (N_1265,N_1140,N_1143);
or U1266 (N_1266,N_1119,N_1123);
and U1267 (N_1267,N_1125,N_1189);
or U1268 (N_1268,N_1166,N_1151);
or U1269 (N_1269,N_1168,N_1130);
or U1270 (N_1270,N_1180,N_1170);
or U1271 (N_1271,N_1119,N_1196);
nor U1272 (N_1272,N_1195,N_1146);
and U1273 (N_1273,N_1153,N_1160);
xor U1274 (N_1274,N_1177,N_1196);
nor U1275 (N_1275,N_1124,N_1188);
or U1276 (N_1276,N_1169,N_1101);
and U1277 (N_1277,N_1170,N_1171);
and U1278 (N_1278,N_1150,N_1187);
xor U1279 (N_1279,N_1126,N_1103);
xor U1280 (N_1280,N_1135,N_1124);
nor U1281 (N_1281,N_1169,N_1145);
nand U1282 (N_1282,N_1162,N_1127);
nor U1283 (N_1283,N_1137,N_1135);
nor U1284 (N_1284,N_1194,N_1136);
and U1285 (N_1285,N_1145,N_1166);
and U1286 (N_1286,N_1178,N_1124);
nor U1287 (N_1287,N_1146,N_1125);
and U1288 (N_1288,N_1165,N_1123);
xor U1289 (N_1289,N_1138,N_1146);
nand U1290 (N_1290,N_1177,N_1126);
nand U1291 (N_1291,N_1163,N_1173);
nor U1292 (N_1292,N_1152,N_1167);
nand U1293 (N_1293,N_1133,N_1148);
xnor U1294 (N_1294,N_1139,N_1107);
nand U1295 (N_1295,N_1159,N_1172);
nor U1296 (N_1296,N_1150,N_1138);
xnor U1297 (N_1297,N_1139,N_1178);
and U1298 (N_1298,N_1100,N_1192);
or U1299 (N_1299,N_1144,N_1143);
xnor U1300 (N_1300,N_1291,N_1236);
nand U1301 (N_1301,N_1204,N_1215);
nand U1302 (N_1302,N_1229,N_1235);
xnor U1303 (N_1303,N_1203,N_1240);
nand U1304 (N_1304,N_1208,N_1216);
nand U1305 (N_1305,N_1209,N_1259);
nand U1306 (N_1306,N_1275,N_1276);
or U1307 (N_1307,N_1232,N_1256);
or U1308 (N_1308,N_1233,N_1282);
xnor U1309 (N_1309,N_1299,N_1292);
xor U1310 (N_1310,N_1225,N_1254);
nand U1311 (N_1311,N_1205,N_1290);
nor U1312 (N_1312,N_1245,N_1287);
and U1313 (N_1313,N_1249,N_1202);
and U1314 (N_1314,N_1241,N_1220);
and U1315 (N_1315,N_1212,N_1253);
or U1316 (N_1316,N_1281,N_1234);
nor U1317 (N_1317,N_1297,N_1265);
xnor U1318 (N_1318,N_1255,N_1268);
xnor U1319 (N_1319,N_1207,N_1261);
xor U1320 (N_1320,N_1248,N_1266);
xor U1321 (N_1321,N_1201,N_1228);
nor U1322 (N_1322,N_1243,N_1277);
nand U1323 (N_1323,N_1267,N_1285);
nand U1324 (N_1324,N_1223,N_1284);
nor U1325 (N_1325,N_1280,N_1227);
and U1326 (N_1326,N_1238,N_1264);
or U1327 (N_1327,N_1226,N_1257);
and U1328 (N_1328,N_1237,N_1239);
and U1329 (N_1329,N_1288,N_1294);
nand U1330 (N_1330,N_1224,N_1263);
and U1331 (N_1331,N_1273,N_1279);
or U1332 (N_1332,N_1272,N_1222);
or U1333 (N_1333,N_1217,N_1247);
nand U1334 (N_1334,N_1251,N_1211);
and U1335 (N_1335,N_1298,N_1293);
or U1336 (N_1336,N_1286,N_1260);
xnor U1337 (N_1337,N_1221,N_1289);
and U1338 (N_1338,N_1271,N_1283);
nand U1339 (N_1339,N_1231,N_1250);
nand U1340 (N_1340,N_1295,N_1206);
xor U1341 (N_1341,N_1242,N_1213);
and U1342 (N_1342,N_1278,N_1269);
and U1343 (N_1343,N_1270,N_1219);
xor U1344 (N_1344,N_1218,N_1244);
and U1345 (N_1345,N_1200,N_1210);
nor U1346 (N_1346,N_1258,N_1214);
nand U1347 (N_1347,N_1296,N_1252);
and U1348 (N_1348,N_1274,N_1246);
and U1349 (N_1349,N_1230,N_1262);
xor U1350 (N_1350,N_1224,N_1285);
nand U1351 (N_1351,N_1279,N_1218);
xor U1352 (N_1352,N_1255,N_1286);
and U1353 (N_1353,N_1228,N_1240);
xor U1354 (N_1354,N_1254,N_1209);
xor U1355 (N_1355,N_1237,N_1209);
or U1356 (N_1356,N_1268,N_1211);
xor U1357 (N_1357,N_1279,N_1238);
xnor U1358 (N_1358,N_1215,N_1262);
xnor U1359 (N_1359,N_1280,N_1263);
nor U1360 (N_1360,N_1247,N_1273);
xnor U1361 (N_1361,N_1205,N_1267);
and U1362 (N_1362,N_1254,N_1202);
or U1363 (N_1363,N_1247,N_1219);
or U1364 (N_1364,N_1226,N_1243);
xor U1365 (N_1365,N_1211,N_1238);
xnor U1366 (N_1366,N_1266,N_1295);
nand U1367 (N_1367,N_1224,N_1280);
nand U1368 (N_1368,N_1224,N_1294);
xor U1369 (N_1369,N_1263,N_1265);
xor U1370 (N_1370,N_1261,N_1282);
nand U1371 (N_1371,N_1247,N_1237);
xor U1372 (N_1372,N_1204,N_1238);
nor U1373 (N_1373,N_1216,N_1254);
xor U1374 (N_1374,N_1267,N_1282);
nand U1375 (N_1375,N_1276,N_1232);
xnor U1376 (N_1376,N_1256,N_1234);
nor U1377 (N_1377,N_1279,N_1213);
and U1378 (N_1378,N_1241,N_1258);
nand U1379 (N_1379,N_1288,N_1204);
nand U1380 (N_1380,N_1233,N_1291);
xnor U1381 (N_1381,N_1283,N_1292);
and U1382 (N_1382,N_1292,N_1293);
xor U1383 (N_1383,N_1262,N_1269);
or U1384 (N_1384,N_1217,N_1273);
or U1385 (N_1385,N_1245,N_1267);
or U1386 (N_1386,N_1206,N_1265);
xor U1387 (N_1387,N_1278,N_1238);
nor U1388 (N_1388,N_1259,N_1279);
nor U1389 (N_1389,N_1259,N_1269);
and U1390 (N_1390,N_1255,N_1249);
and U1391 (N_1391,N_1248,N_1271);
and U1392 (N_1392,N_1270,N_1278);
and U1393 (N_1393,N_1258,N_1208);
or U1394 (N_1394,N_1271,N_1272);
or U1395 (N_1395,N_1275,N_1282);
nand U1396 (N_1396,N_1278,N_1281);
and U1397 (N_1397,N_1299,N_1287);
nand U1398 (N_1398,N_1256,N_1249);
or U1399 (N_1399,N_1258,N_1218);
nand U1400 (N_1400,N_1351,N_1314);
nand U1401 (N_1401,N_1374,N_1367);
xnor U1402 (N_1402,N_1303,N_1327);
and U1403 (N_1403,N_1317,N_1353);
nand U1404 (N_1404,N_1312,N_1399);
or U1405 (N_1405,N_1392,N_1373);
nand U1406 (N_1406,N_1338,N_1335);
and U1407 (N_1407,N_1326,N_1302);
nand U1408 (N_1408,N_1304,N_1390);
xor U1409 (N_1409,N_1319,N_1365);
nor U1410 (N_1410,N_1388,N_1358);
nand U1411 (N_1411,N_1386,N_1300);
and U1412 (N_1412,N_1389,N_1330);
nand U1413 (N_1413,N_1307,N_1380);
and U1414 (N_1414,N_1336,N_1339);
nor U1415 (N_1415,N_1345,N_1359);
xnor U1416 (N_1416,N_1379,N_1316);
or U1417 (N_1417,N_1342,N_1385);
nor U1418 (N_1418,N_1320,N_1352);
and U1419 (N_1419,N_1364,N_1310);
and U1420 (N_1420,N_1331,N_1377);
xnor U1421 (N_1421,N_1370,N_1332);
nand U1422 (N_1422,N_1362,N_1371);
nor U1423 (N_1423,N_1395,N_1381);
xnor U1424 (N_1424,N_1369,N_1325);
xnor U1425 (N_1425,N_1382,N_1321);
or U1426 (N_1426,N_1340,N_1383);
xnor U1427 (N_1427,N_1305,N_1355);
and U1428 (N_1428,N_1391,N_1356);
nand U1429 (N_1429,N_1396,N_1311);
or U1430 (N_1430,N_1322,N_1366);
and U1431 (N_1431,N_1368,N_1308);
nor U1432 (N_1432,N_1309,N_1376);
nor U1433 (N_1433,N_1384,N_1318);
and U1434 (N_1434,N_1346,N_1349);
nor U1435 (N_1435,N_1324,N_1357);
nand U1436 (N_1436,N_1306,N_1360);
and U1437 (N_1437,N_1387,N_1341);
xnor U1438 (N_1438,N_1323,N_1344);
or U1439 (N_1439,N_1363,N_1337);
nor U1440 (N_1440,N_1397,N_1354);
xnor U1441 (N_1441,N_1334,N_1347);
nand U1442 (N_1442,N_1372,N_1343);
and U1443 (N_1443,N_1333,N_1375);
or U1444 (N_1444,N_1393,N_1329);
xnor U1445 (N_1445,N_1350,N_1328);
nand U1446 (N_1446,N_1315,N_1348);
and U1447 (N_1447,N_1361,N_1398);
nand U1448 (N_1448,N_1313,N_1378);
or U1449 (N_1449,N_1301,N_1394);
or U1450 (N_1450,N_1370,N_1344);
and U1451 (N_1451,N_1328,N_1314);
nand U1452 (N_1452,N_1336,N_1390);
nand U1453 (N_1453,N_1325,N_1385);
and U1454 (N_1454,N_1381,N_1317);
nor U1455 (N_1455,N_1355,N_1398);
and U1456 (N_1456,N_1366,N_1304);
nand U1457 (N_1457,N_1364,N_1328);
nor U1458 (N_1458,N_1390,N_1314);
nor U1459 (N_1459,N_1370,N_1342);
xor U1460 (N_1460,N_1361,N_1345);
and U1461 (N_1461,N_1381,N_1365);
nor U1462 (N_1462,N_1301,N_1374);
and U1463 (N_1463,N_1372,N_1362);
nand U1464 (N_1464,N_1349,N_1308);
nand U1465 (N_1465,N_1350,N_1315);
xnor U1466 (N_1466,N_1361,N_1377);
xnor U1467 (N_1467,N_1326,N_1348);
nand U1468 (N_1468,N_1378,N_1319);
xnor U1469 (N_1469,N_1374,N_1306);
nand U1470 (N_1470,N_1334,N_1306);
xor U1471 (N_1471,N_1390,N_1348);
xor U1472 (N_1472,N_1382,N_1319);
nand U1473 (N_1473,N_1317,N_1303);
or U1474 (N_1474,N_1371,N_1345);
xnor U1475 (N_1475,N_1311,N_1346);
xor U1476 (N_1476,N_1387,N_1300);
nor U1477 (N_1477,N_1316,N_1385);
nand U1478 (N_1478,N_1393,N_1354);
nand U1479 (N_1479,N_1370,N_1334);
nor U1480 (N_1480,N_1337,N_1365);
and U1481 (N_1481,N_1382,N_1381);
or U1482 (N_1482,N_1381,N_1354);
or U1483 (N_1483,N_1390,N_1377);
and U1484 (N_1484,N_1353,N_1320);
nor U1485 (N_1485,N_1350,N_1391);
nor U1486 (N_1486,N_1323,N_1375);
and U1487 (N_1487,N_1386,N_1347);
and U1488 (N_1488,N_1393,N_1326);
nor U1489 (N_1489,N_1311,N_1356);
and U1490 (N_1490,N_1317,N_1307);
nor U1491 (N_1491,N_1330,N_1322);
and U1492 (N_1492,N_1300,N_1304);
xor U1493 (N_1493,N_1317,N_1344);
xor U1494 (N_1494,N_1320,N_1326);
xor U1495 (N_1495,N_1336,N_1363);
nor U1496 (N_1496,N_1377,N_1398);
and U1497 (N_1497,N_1371,N_1320);
nand U1498 (N_1498,N_1389,N_1399);
nor U1499 (N_1499,N_1381,N_1337);
xor U1500 (N_1500,N_1402,N_1419);
and U1501 (N_1501,N_1496,N_1476);
nor U1502 (N_1502,N_1406,N_1428);
and U1503 (N_1503,N_1450,N_1446);
nand U1504 (N_1504,N_1497,N_1417);
and U1505 (N_1505,N_1429,N_1480);
xnor U1506 (N_1506,N_1463,N_1412);
nand U1507 (N_1507,N_1478,N_1499);
xnor U1508 (N_1508,N_1473,N_1423);
nand U1509 (N_1509,N_1411,N_1483);
and U1510 (N_1510,N_1413,N_1467);
nand U1511 (N_1511,N_1453,N_1470);
and U1512 (N_1512,N_1471,N_1454);
nand U1513 (N_1513,N_1448,N_1439);
nand U1514 (N_1514,N_1420,N_1431);
and U1515 (N_1515,N_1445,N_1484);
xor U1516 (N_1516,N_1481,N_1493);
or U1517 (N_1517,N_1438,N_1447);
nor U1518 (N_1518,N_1422,N_1425);
and U1519 (N_1519,N_1440,N_1458);
nand U1520 (N_1520,N_1490,N_1430);
or U1521 (N_1521,N_1477,N_1415);
xor U1522 (N_1522,N_1407,N_1414);
xnor U1523 (N_1523,N_1427,N_1482);
nor U1524 (N_1524,N_1472,N_1469);
or U1525 (N_1525,N_1487,N_1442);
nand U1526 (N_1526,N_1491,N_1410);
xnor U1527 (N_1527,N_1461,N_1432);
or U1528 (N_1528,N_1409,N_1451);
nor U1529 (N_1529,N_1456,N_1441);
nor U1530 (N_1530,N_1489,N_1455);
or U1531 (N_1531,N_1449,N_1464);
or U1532 (N_1532,N_1479,N_1457);
nand U1533 (N_1533,N_1421,N_1460);
xor U1534 (N_1534,N_1494,N_1433);
or U1535 (N_1535,N_1486,N_1405);
xnor U1536 (N_1536,N_1434,N_1401);
nor U1537 (N_1537,N_1485,N_1474);
nor U1538 (N_1538,N_1475,N_1403);
and U1539 (N_1539,N_1424,N_1495);
and U1540 (N_1540,N_1465,N_1452);
nand U1541 (N_1541,N_1492,N_1408);
nand U1542 (N_1542,N_1404,N_1418);
or U1543 (N_1543,N_1468,N_1426);
xor U1544 (N_1544,N_1462,N_1437);
nand U1545 (N_1545,N_1466,N_1443);
and U1546 (N_1546,N_1416,N_1400);
and U1547 (N_1547,N_1459,N_1498);
nor U1548 (N_1548,N_1488,N_1444);
and U1549 (N_1549,N_1435,N_1436);
xor U1550 (N_1550,N_1471,N_1489);
nor U1551 (N_1551,N_1435,N_1496);
and U1552 (N_1552,N_1489,N_1454);
or U1553 (N_1553,N_1486,N_1494);
and U1554 (N_1554,N_1427,N_1432);
xor U1555 (N_1555,N_1401,N_1488);
or U1556 (N_1556,N_1456,N_1489);
or U1557 (N_1557,N_1465,N_1482);
nor U1558 (N_1558,N_1484,N_1482);
or U1559 (N_1559,N_1472,N_1492);
nand U1560 (N_1560,N_1445,N_1424);
xnor U1561 (N_1561,N_1481,N_1480);
nand U1562 (N_1562,N_1456,N_1445);
nor U1563 (N_1563,N_1409,N_1473);
nor U1564 (N_1564,N_1424,N_1449);
nand U1565 (N_1565,N_1473,N_1408);
or U1566 (N_1566,N_1481,N_1412);
xnor U1567 (N_1567,N_1410,N_1400);
or U1568 (N_1568,N_1485,N_1437);
or U1569 (N_1569,N_1421,N_1479);
xnor U1570 (N_1570,N_1478,N_1432);
and U1571 (N_1571,N_1456,N_1424);
nor U1572 (N_1572,N_1410,N_1426);
or U1573 (N_1573,N_1416,N_1425);
or U1574 (N_1574,N_1497,N_1458);
and U1575 (N_1575,N_1410,N_1444);
or U1576 (N_1576,N_1452,N_1496);
nor U1577 (N_1577,N_1494,N_1444);
nand U1578 (N_1578,N_1402,N_1434);
or U1579 (N_1579,N_1496,N_1420);
xor U1580 (N_1580,N_1466,N_1496);
xnor U1581 (N_1581,N_1432,N_1450);
and U1582 (N_1582,N_1430,N_1467);
and U1583 (N_1583,N_1445,N_1406);
xor U1584 (N_1584,N_1464,N_1453);
and U1585 (N_1585,N_1488,N_1414);
and U1586 (N_1586,N_1483,N_1462);
or U1587 (N_1587,N_1430,N_1461);
and U1588 (N_1588,N_1413,N_1408);
and U1589 (N_1589,N_1426,N_1417);
and U1590 (N_1590,N_1406,N_1478);
nor U1591 (N_1591,N_1476,N_1468);
nor U1592 (N_1592,N_1498,N_1484);
nand U1593 (N_1593,N_1468,N_1425);
nand U1594 (N_1594,N_1408,N_1486);
nor U1595 (N_1595,N_1466,N_1478);
or U1596 (N_1596,N_1424,N_1458);
or U1597 (N_1597,N_1428,N_1495);
nand U1598 (N_1598,N_1423,N_1446);
nor U1599 (N_1599,N_1417,N_1445);
nand U1600 (N_1600,N_1573,N_1507);
or U1601 (N_1601,N_1540,N_1593);
nor U1602 (N_1602,N_1519,N_1553);
or U1603 (N_1603,N_1574,N_1558);
or U1604 (N_1604,N_1568,N_1571);
xnor U1605 (N_1605,N_1564,N_1576);
nor U1606 (N_1606,N_1597,N_1542);
xnor U1607 (N_1607,N_1515,N_1534);
and U1608 (N_1608,N_1524,N_1520);
nor U1609 (N_1609,N_1548,N_1554);
nand U1610 (N_1610,N_1545,N_1580);
xor U1611 (N_1611,N_1594,N_1541);
nor U1612 (N_1612,N_1560,N_1591);
nand U1613 (N_1613,N_1508,N_1517);
nor U1614 (N_1614,N_1575,N_1533);
nor U1615 (N_1615,N_1543,N_1556);
nand U1616 (N_1616,N_1555,N_1501);
nor U1617 (N_1617,N_1536,N_1527);
nor U1618 (N_1618,N_1566,N_1522);
and U1619 (N_1619,N_1549,N_1595);
nor U1620 (N_1620,N_1559,N_1572);
xnor U1621 (N_1621,N_1510,N_1526);
xnor U1622 (N_1622,N_1562,N_1577);
and U1623 (N_1623,N_1539,N_1504);
nand U1624 (N_1624,N_1523,N_1537);
and U1625 (N_1625,N_1531,N_1582);
or U1626 (N_1626,N_1567,N_1563);
xor U1627 (N_1627,N_1599,N_1551);
xnor U1628 (N_1628,N_1506,N_1552);
nor U1629 (N_1629,N_1511,N_1502);
nand U1630 (N_1630,N_1544,N_1588);
xnor U1631 (N_1631,N_1592,N_1532);
nor U1632 (N_1632,N_1578,N_1561);
or U1633 (N_1633,N_1585,N_1535);
or U1634 (N_1634,N_1521,N_1518);
nand U1635 (N_1635,N_1529,N_1587);
and U1636 (N_1636,N_1528,N_1579);
xnor U1637 (N_1637,N_1589,N_1584);
or U1638 (N_1638,N_1503,N_1581);
nand U1639 (N_1639,N_1514,N_1513);
nand U1640 (N_1640,N_1590,N_1538);
nor U1641 (N_1641,N_1505,N_1500);
xnor U1642 (N_1642,N_1530,N_1546);
and U1643 (N_1643,N_1583,N_1516);
and U1644 (N_1644,N_1550,N_1586);
nor U1645 (N_1645,N_1569,N_1557);
nand U1646 (N_1646,N_1547,N_1509);
nor U1647 (N_1647,N_1570,N_1512);
xnor U1648 (N_1648,N_1596,N_1525);
and U1649 (N_1649,N_1598,N_1565);
nor U1650 (N_1650,N_1561,N_1562);
nor U1651 (N_1651,N_1531,N_1555);
nand U1652 (N_1652,N_1534,N_1532);
and U1653 (N_1653,N_1577,N_1518);
xor U1654 (N_1654,N_1562,N_1503);
or U1655 (N_1655,N_1586,N_1536);
or U1656 (N_1656,N_1549,N_1564);
xnor U1657 (N_1657,N_1505,N_1547);
nor U1658 (N_1658,N_1515,N_1599);
or U1659 (N_1659,N_1513,N_1506);
nand U1660 (N_1660,N_1583,N_1546);
nand U1661 (N_1661,N_1527,N_1552);
nor U1662 (N_1662,N_1595,N_1501);
or U1663 (N_1663,N_1594,N_1526);
xor U1664 (N_1664,N_1551,N_1555);
or U1665 (N_1665,N_1585,N_1508);
and U1666 (N_1666,N_1547,N_1560);
or U1667 (N_1667,N_1580,N_1525);
nor U1668 (N_1668,N_1568,N_1537);
nor U1669 (N_1669,N_1560,N_1525);
nor U1670 (N_1670,N_1573,N_1519);
nand U1671 (N_1671,N_1553,N_1582);
and U1672 (N_1672,N_1526,N_1592);
nand U1673 (N_1673,N_1598,N_1523);
xor U1674 (N_1674,N_1506,N_1594);
xnor U1675 (N_1675,N_1582,N_1523);
or U1676 (N_1676,N_1589,N_1523);
and U1677 (N_1677,N_1589,N_1548);
xor U1678 (N_1678,N_1588,N_1594);
or U1679 (N_1679,N_1594,N_1543);
nor U1680 (N_1680,N_1581,N_1512);
nor U1681 (N_1681,N_1550,N_1512);
nand U1682 (N_1682,N_1563,N_1542);
or U1683 (N_1683,N_1536,N_1535);
and U1684 (N_1684,N_1573,N_1528);
or U1685 (N_1685,N_1574,N_1538);
nor U1686 (N_1686,N_1503,N_1549);
nor U1687 (N_1687,N_1594,N_1524);
nor U1688 (N_1688,N_1551,N_1536);
nand U1689 (N_1689,N_1534,N_1554);
xnor U1690 (N_1690,N_1546,N_1513);
xnor U1691 (N_1691,N_1539,N_1568);
nand U1692 (N_1692,N_1539,N_1526);
xnor U1693 (N_1693,N_1557,N_1503);
and U1694 (N_1694,N_1529,N_1597);
xor U1695 (N_1695,N_1512,N_1561);
or U1696 (N_1696,N_1521,N_1505);
xnor U1697 (N_1697,N_1520,N_1518);
nand U1698 (N_1698,N_1583,N_1584);
xor U1699 (N_1699,N_1508,N_1593);
and U1700 (N_1700,N_1698,N_1609);
or U1701 (N_1701,N_1639,N_1648);
nand U1702 (N_1702,N_1663,N_1687);
nand U1703 (N_1703,N_1682,N_1679);
xor U1704 (N_1704,N_1652,N_1670);
nand U1705 (N_1705,N_1684,N_1661);
and U1706 (N_1706,N_1633,N_1653);
or U1707 (N_1707,N_1608,N_1631);
xnor U1708 (N_1708,N_1641,N_1655);
nand U1709 (N_1709,N_1656,N_1681);
or U1710 (N_1710,N_1634,N_1636);
or U1711 (N_1711,N_1632,N_1697);
xnor U1712 (N_1712,N_1692,N_1628);
and U1713 (N_1713,N_1635,N_1605);
or U1714 (N_1714,N_1696,N_1650);
nor U1715 (N_1715,N_1690,N_1668);
nand U1716 (N_1716,N_1676,N_1638);
or U1717 (N_1717,N_1699,N_1658);
xnor U1718 (N_1718,N_1610,N_1604);
nor U1719 (N_1719,N_1616,N_1654);
or U1720 (N_1720,N_1615,N_1691);
nor U1721 (N_1721,N_1671,N_1611);
nor U1722 (N_1722,N_1625,N_1665);
nor U1723 (N_1723,N_1620,N_1642);
and U1724 (N_1724,N_1600,N_1694);
nor U1725 (N_1725,N_1629,N_1680);
and U1726 (N_1726,N_1624,N_1622);
xnor U1727 (N_1727,N_1667,N_1607);
nand U1728 (N_1728,N_1657,N_1647);
nand U1729 (N_1729,N_1627,N_1602);
xor U1730 (N_1730,N_1664,N_1689);
or U1731 (N_1731,N_1659,N_1614);
nor U1732 (N_1732,N_1660,N_1677);
or U1733 (N_1733,N_1637,N_1603);
or U1734 (N_1734,N_1662,N_1651);
and U1735 (N_1735,N_1685,N_1618);
nand U1736 (N_1736,N_1649,N_1619);
or U1737 (N_1737,N_1675,N_1645);
nor U1738 (N_1738,N_1621,N_1646);
or U1739 (N_1739,N_1623,N_1606);
nor U1740 (N_1740,N_1669,N_1674);
and U1741 (N_1741,N_1686,N_1626);
nor U1742 (N_1742,N_1683,N_1693);
or U1743 (N_1743,N_1644,N_1673);
nand U1744 (N_1744,N_1666,N_1630);
nor U1745 (N_1745,N_1640,N_1643);
or U1746 (N_1746,N_1688,N_1613);
or U1747 (N_1747,N_1678,N_1617);
and U1748 (N_1748,N_1601,N_1672);
or U1749 (N_1749,N_1695,N_1612);
nand U1750 (N_1750,N_1657,N_1636);
xnor U1751 (N_1751,N_1614,N_1684);
or U1752 (N_1752,N_1622,N_1690);
and U1753 (N_1753,N_1601,N_1657);
and U1754 (N_1754,N_1674,N_1621);
xnor U1755 (N_1755,N_1626,N_1628);
and U1756 (N_1756,N_1693,N_1659);
nand U1757 (N_1757,N_1686,N_1660);
nand U1758 (N_1758,N_1606,N_1603);
and U1759 (N_1759,N_1647,N_1698);
and U1760 (N_1760,N_1683,N_1645);
nand U1761 (N_1761,N_1638,N_1620);
xnor U1762 (N_1762,N_1690,N_1611);
nor U1763 (N_1763,N_1696,N_1699);
or U1764 (N_1764,N_1644,N_1659);
xnor U1765 (N_1765,N_1616,N_1610);
or U1766 (N_1766,N_1627,N_1624);
xnor U1767 (N_1767,N_1618,N_1615);
xnor U1768 (N_1768,N_1635,N_1640);
xnor U1769 (N_1769,N_1610,N_1652);
nor U1770 (N_1770,N_1619,N_1633);
nor U1771 (N_1771,N_1602,N_1675);
xnor U1772 (N_1772,N_1600,N_1623);
or U1773 (N_1773,N_1600,N_1648);
xor U1774 (N_1774,N_1653,N_1687);
xor U1775 (N_1775,N_1661,N_1663);
nand U1776 (N_1776,N_1649,N_1625);
nand U1777 (N_1777,N_1606,N_1696);
nand U1778 (N_1778,N_1659,N_1664);
xor U1779 (N_1779,N_1693,N_1628);
or U1780 (N_1780,N_1632,N_1652);
or U1781 (N_1781,N_1606,N_1649);
nor U1782 (N_1782,N_1608,N_1642);
nand U1783 (N_1783,N_1652,N_1667);
and U1784 (N_1784,N_1651,N_1602);
and U1785 (N_1785,N_1689,N_1600);
and U1786 (N_1786,N_1606,N_1657);
or U1787 (N_1787,N_1600,N_1622);
xor U1788 (N_1788,N_1698,N_1641);
and U1789 (N_1789,N_1697,N_1694);
xnor U1790 (N_1790,N_1646,N_1644);
nand U1791 (N_1791,N_1643,N_1671);
and U1792 (N_1792,N_1614,N_1689);
xor U1793 (N_1793,N_1638,N_1621);
nor U1794 (N_1794,N_1604,N_1633);
nor U1795 (N_1795,N_1675,N_1670);
or U1796 (N_1796,N_1698,N_1639);
nor U1797 (N_1797,N_1602,N_1603);
and U1798 (N_1798,N_1606,N_1658);
nand U1799 (N_1799,N_1602,N_1632);
and U1800 (N_1800,N_1797,N_1702);
xnor U1801 (N_1801,N_1708,N_1748);
nand U1802 (N_1802,N_1795,N_1787);
and U1803 (N_1803,N_1779,N_1762);
nand U1804 (N_1804,N_1780,N_1730);
and U1805 (N_1805,N_1798,N_1754);
or U1806 (N_1806,N_1765,N_1746);
nor U1807 (N_1807,N_1706,N_1733);
or U1808 (N_1808,N_1727,N_1741);
nand U1809 (N_1809,N_1770,N_1731);
nand U1810 (N_1810,N_1734,N_1701);
and U1811 (N_1811,N_1724,N_1715);
xnor U1812 (N_1812,N_1768,N_1720);
or U1813 (N_1813,N_1705,N_1764);
and U1814 (N_1814,N_1703,N_1799);
and U1815 (N_1815,N_1794,N_1796);
nand U1816 (N_1816,N_1784,N_1788);
nor U1817 (N_1817,N_1712,N_1758);
nor U1818 (N_1818,N_1769,N_1700);
xor U1819 (N_1819,N_1726,N_1718);
nand U1820 (N_1820,N_1717,N_1767);
nand U1821 (N_1821,N_1725,N_1789);
nor U1822 (N_1822,N_1742,N_1793);
and U1823 (N_1823,N_1719,N_1778);
nand U1824 (N_1824,N_1745,N_1756);
xnor U1825 (N_1825,N_1721,N_1786);
xor U1826 (N_1826,N_1753,N_1760);
nand U1827 (N_1827,N_1713,N_1743);
or U1828 (N_1828,N_1776,N_1785);
nor U1829 (N_1829,N_1747,N_1729);
nand U1830 (N_1830,N_1736,N_1722);
or U1831 (N_1831,N_1750,N_1792);
and U1832 (N_1832,N_1766,N_1757);
nor U1833 (N_1833,N_1759,N_1755);
and U1834 (N_1834,N_1710,N_1709);
or U1835 (N_1835,N_1775,N_1751);
nand U1836 (N_1836,N_1704,N_1723);
xor U1837 (N_1837,N_1782,N_1737);
nor U1838 (N_1838,N_1771,N_1772);
nor U1839 (N_1839,N_1777,N_1716);
and U1840 (N_1840,N_1714,N_1711);
and U1841 (N_1841,N_1783,N_1761);
or U1842 (N_1842,N_1774,N_1773);
xnor U1843 (N_1843,N_1763,N_1790);
xnor U1844 (N_1844,N_1791,N_1781);
or U1845 (N_1845,N_1744,N_1740);
or U1846 (N_1846,N_1735,N_1728);
and U1847 (N_1847,N_1707,N_1752);
or U1848 (N_1848,N_1732,N_1738);
nor U1849 (N_1849,N_1749,N_1739);
or U1850 (N_1850,N_1793,N_1726);
nand U1851 (N_1851,N_1742,N_1752);
nor U1852 (N_1852,N_1743,N_1724);
nand U1853 (N_1853,N_1720,N_1744);
nand U1854 (N_1854,N_1774,N_1731);
nor U1855 (N_1855,N_1769,N_1747);
nor U1856 (N_1856,N_1787,N_1725);
or U1857 (N_1857,N_1758,N_1728);
nand U1858 (N_1858,N_1758,N_1788);
nand U1859 (N_1859,N_1722,N_1720);
and U1860 (N_1860,N_1797,N_1755);
xor U1861 (N_1861,N_1769,N_1755);
and U1862 (N_1862,N_1778,N_1727);
nor U1863 (N_1863,N_1765,N_1709);
nand U1864 (N_1864,N_1797,N_1740);
xor U1865 (N_1865,N_1781,N_1727);
nand U1866 (N_1866,N_1702,N_1775);
nor U1867 (N_1867,N_1755,N_1719);
and U1868 (N_1868,N_1793,N_1784);
xnor U1869 (N_1869,N_1728,N_1738);
nor U1870 (N_1870,N_1797,N_1752);
and U1871 (N_1871,N_1767,N_1796);
nor U1872 (N_1872,N_1740,N_1738);
nand U1873 (N_1873,N_1722,N_1743);
or U1874 (N_1874,N_1782,N_1767);
or U1875 (N_1875,N_1712,N_1709);
nor U1876 (N_1876,N_1751,N_1701);
and U1877 (N_1877,N_1706,N_1768);
nor U1878 (N_1878,N_1761,N_1750);
xnor U1879 (N_1879,N_1711,N_1731);
or U1880 (N_1880,N_1735,N_1768);
nand U1881 (N_1881,N_1738,N_1725);
nor U1882 (N_1882,N_1765,N_1710);
and U1883 (N_1883,N_1731,N_1763);
xnor U1884 (N_1884,N_1767,N_1726);
and U1885 (N_1885,N_1758,N_1718);
nor U1886 (N_1886,N_1790,N_1749);
nand U1887 (N_1887,N_1781,N_1758);
nor U1888 (N_1888,N_1725,N_1781);
nand U1889 (N_1889,N_1796,N_1789);
xnor U1890 (N_1890,N_1771,N_1742);
or U1891 (N_1891,N_1794,N_1771);
nor U1892 (N_1892,N_1729,N_1738);
nand U1893 (N_1893,N_1708,N_1774);
and U1894 (N_1894,N_1768,N_1751);
xnor U1895 (N_1895,N_1789,N_1729);
nor U1896 (N_1896,N_1701,N_1765);
xor U1897 (N_1897,N_1756,N_1764);
xor U1898 (N_1898,N_1779,N_1717);
xor U1899 (N_1899,N_1760,N_1793);
and U1900 (N_1900,N_1840,N_1820);
xor U1901 (N_1901,N_1835,N_1803);
or U1902 (N_1902,N_1823,N_1892);
or U1903 (N_1903,N_1811,N_1836);
and U1904 (N_1904,N_1813,N_1885);
or U1905 (N_1905,N_1893,N_1867);
nor U1906 (N_1906,N_1814,N_1805);
nor U1907 (N_1907,N_1852,N_1812);
xor U1908 (N_1908,N_1866,N_1858);
nand U1909 (N_1909,N_1828,N_1869);
xor U1910 (N_1910,N_1883,N_1861);
or U1911 (N_1911,N_1880,N_1879);
and U1912 (N_1912,N_1894,N_1872);
nand U1913 (N_1913,N_1897,N_1824);
or U1914 (N_1914,N_1864,N_1826);
xor U1915 (N_1915,N_1850,N_1833);
xnor U1916 (N_1916,N_1846,N_1874);
and U1917 (N_1917,N_1806,N_1856);
nor U1918 (N_1918,N_1888,N_1825);
xor U1919 (N_1919,N_1822,N_1863);
nand U1920 (N_1920,N_1878,N_1834);
and U1921 (N_1921,N_1807,N_1838);
nand U1922 (N_1922,N_1873,N_1890);
nor U1923 (N_1923,N_1875,N_1818);
or U1924 (N_1924,N_1821,N_1801);
nand U1925 (N_1925,N_1809,N_1886);
or U1926 (N_1926,N_1816,N_1857);
or U1927 (N_1927,N_1843,N_1815);
xnor U1928 (N_1928,N_1877,N_1804);
or U1929 (N_1929,N_1808,N_1881);
xnor U1930 (N_1930,N_1889,N_1845);
xor U1931 (N_1931,N_1896,N_1841);
xor U1932 (N_1932,N_1830,N_1895);
nand U1933 (N_1933,N_1839,N_1870);
nand U1934 (N_1934,N_1800,N_1898);
nor U1935 (N_1935,N_1860,N_1810);
nand U1936 (N_1936,N_1868,N_1899);
or U1937 (N_1937,N_1819,N_1848);
xor U1938 (N_1938,N_1851,N_1831);
and U1939 (N_1939,N_1855,N_1849);
nand U1940 (N_1940,N_1882,N_1802);
or U1941 (N_1941,N_1827,N_1817);
nor U1942 (N_1942,N_1842,N_1862);
and U1943 (N_1943,N_1837,N_1844);
or U1944 (N_1944,N_1854,N_1891);
or U1945 (N_1945,N_1865,N_1847);
or U1946 (N_1946,N_1871,N_1884);
or U1947 (N_1947,N_1859,N_1832);
and U1948 (N_1948,N_1829,N_1887);
nand U1949 (N_1949,N_1876,N_1853);
or U1950 (N_1950,N_1813,N_1809);
nand U1951 (N_1951,N_1877,N_1890);
nand U1952 (N_1952,N_1867,N_1848);
nand U1953 (N_1953,N_1816,N_1851);
nand U1954 (N_1954,N_1875,N_1880);
nand U1955 (N_1955,N_1822,N_1830);
and U1956 (N_1956,N_1815,N_1898);
and U1957 (N_1957,N_1872,N_1820);
nor U1958 (N_1958,N_1869,N_1887);
xor U1959 (N_1959,N_1890,N_1869);
or U1960 (N_1960,N_1809,N_1847);
nand U1961 (N_1961,N_1822,N_1856);
xor U1962 (N_1962,N_1885,N_1831);
xor U1963 (N_1963,N_1875,N_1891);
nand U1964 (N_1964,N_1829,N_1843);
xnor U1965 (N_1965,N_1839,N_1880);
xnor U1966 (N_1966,N_1800,N_1813);
nor U1967 (N_1967,N_1856,N_1889);
or U1968 (N_1968,N_1860,N_1832);
nand U1969 (N_1969,N_1854,N_1895);
nand U1970 (N_1970,N_1836,N_1889);
and U1971 (N_1971,N_1844,N_1888);
xor U1972 (N_1972,N_1801,N_1806);
nor U1973 (N_1973,N_1850,N_1886);
nor U1974 (N_1974,N_1874,N_1862);
nand U1975 (N_1975,N_1837,N_1861);
and U1976 (N_1976,N_1892,N_1816);
xnor U1977 (N_1977,N_1823,N_1805);
xnor U1978 (N_1978,N_1820,N_1821);
or U1979 (N_1979,N_1812,N_1819);
or U1980 (N_1980,N_1857,N_1870);
nor U1981 (N_1981,N_1845,N_1875);
nand U1982 (N_1982,N_1896,N_1872);
nand U1983 (N_1983,N_1803,N_1807);
nor U1984 (N_1984,N_1813,N_1847);
and U1985 (N_1985,N_1816,N_1898);
nand U1986 (N_1986,N_1842,N_1856);
and U1987 (N_1987,N_1855,N_1860);
and U1988 (N_1988,N_1860,N_1875);
nand U1989 (N_1989,N_1879,N_1860);
or U1990 (N_1990,N_1820,N_1851);
nand U1991 (N_1991,N_1836,N_1865);
nor U1992 (N_1992,N_1879,N_1843);
or U1993 (N_1993,N_1810,N_1836);
and U1994 (N_1994,N_1887,N_1839);
nor U1995 (N_1995,N_1859,N_1822);
xnor U1996 (N_1996,N_1837,N_1824);
and U1997 (N_1997,N_1864,N_1855);
xor U1998 (N_1998,N_1854,N_1821);
and U1999 (N_1999,N_1869,N_1862);
xnor U2000 (N_2000,N_1992,N_1914);
xor U2001 (N_2001,N_1926,N_1934);
nand U2002 (N_2002,N_1930,N_1956);
and U2003 (N_2003,N_1971,N_1940);
or U2004 (N_2004,N_1982,N_1901);
or U2005 (N_2005,N_1995,N_1953);
xor U2006 (N_2006,N_1962,N_1900);
nor U2007 (N_2007,N_1924,N_1958);
and U2008 (N_2008,N_1983,N_1975);
nand U2009 (N_2009,N_1970,N_1918);
nand U2010 (N_2010,N_1935,N_1965);
and U2011 (N_2011,N_1951,N_1972);
nor U2012 (N_2012,N_1976,N_1938);
nand U2013 (N_2013,N_1941,N_1966);
or U2014 (N_2014,N_1954,N_1917);
nor U2015 (N_2015,N_1952,N_1990);
and U2016 (N_2016,N_1928,N_1909);
nor U2017 (N_2017,N_1968,N_1932);
xnor U2018 (N_2018,N_1925,N_1997);
nand U2019 (N_2019,N_1937,N_1907);
xnor U2020 (N_2020,N_1994,N_1944);
nand U2021 (N_2021,N_1912,N_1989);
and U2022 (N_2022,N_1949,N_1984);
nor U2023 (N_2023,N_1963,N_1979);
or U2024 (N_2024,N_1945,N_1943);
or U2025 (N_2025,N_1959,N_1916);
and U2026 (N_2026,N_1947,N_1964);
or U2027 (N_2027,N_1920,N_1969);
nor U2028 (N_2028,N_1915,N_1978);
and U2029 (N_2029,N_1957,N_1933);
and U2030 (N_2030,N_1948,N_1911);
xnor U2031 (N_2031,N_1921,N_1927);
or U2032 (N_2032,N_1985,N_1987);
nor U2033 (N_2033,N_1923,N_1902);
nor U2034 (N_2034,N_1960,N_1967);
xor U2035 (N_2035,N_1906,N_1910);
nand U2036 (N_2036,N_1974,N_1905);
xor U2037 (N_2037,N_1908,N_1973);
nor U2038 (N_2038,N_1955,N_1913);
xor U2039 (N_2039,N_1991,N_1929);
and U2040 (N_2040,N_1936,N_1919);
nor U2041 (N_2041,N_1931,N_1988);
nand U2042 (N_2042,N_1942,N_1903);
and U2043 (N_2043,N_1999,N_1961);
or U2044 (N_2044,N_1986,N_1998);
or U2045 (N_2045,N_1981,N_1980);
xnor U2046 (N_2046,N_1950,N_1922);
nor U2047 (N_2047,N_1939,N_1993);
or U2048 (N_2048,N_1904,N_1996);
nor U2049 (N_2049,N_1946,N_1977);
xnor U2050 (N_2050,N_1999,N_1916);
nand U2051 (N_2051,N_1959,N_1996);
nor U2052 (N_2052,N_1994,N_1954);
nand U2053 (N_2053,N_1986,N_1900);
xnor U2054 (N_2054,N_1970,N_1964);
nor U2055 (N_2055,N_1911,N_1944);
or U2056 (N_2056,N_1922,N_1910);
and U2057 (N_2057,N_1933,N_1968);
nand U2058 (N_2058,N_1907,N_1968);
nand U2059 (N_2059,N_1910,N_1967);
and U2060 (N_2060,N_1939,N_1966);
nand U2061 (N_2061,N_1971,N_1969);
nand U2062 (N_2062,N_1972,N_1966);
nor U2063 (N_2063,N_1909,N_1947);
and U2064 (N_2064,N_1932,N_1954);
and U2065 (N_2065,N_1960,N_1989);
nand U2066 (N_2066,N_1982,N_1967);
and U2067 (N_2067,N_1989,N_1902);
xor U2068 (N_2068,N_1907,N_1902);
or U2069 (N_2069,N_1916,N_1947);
or U2070 (N_2070,N_1978,N_1966);
and U2071 (N_2071,N_1931,N_1975);
xor U2072 (N_2072,N_1969,N_1988);
nand U2073 (N_2073,N_1974,N_1934);
nor U2074 (N_2074,N_1937,N_1995);
and U2075 (N_2075,N_1953,N_1991);
nor U2076 (N_2076,N_1934,N_1952);
nand U2077 (N_2077,N_1922,N_1979);
xor U2078 (N_2078,N_1908,N_1931);
nor U2079 (N_2079,N_1905,N_1960);
nor U2080 (N_2080,N_1982,N_1960);
nand U2081 (N_2081,N_1998,N_1963);
or U2082 (N_2082,N_1983,N_1910);
nor U2083 (N_2083,N_1978,N_1910);
and U2084 (N_2084,N_1971,N_1945);
and U2085 (N_2085,N_1952,N_1938);
and U2086 (N_2086,N_1913,N_1941);
or U2087 (N_2087,N_1934,N_1949);
nor U2088 (N_2088,N_1995,N_1968);
or U2089 (N_2089,N_1966,N_1985);
and U2090 (N_2090,N_1901,N_1959);
nand U2091 (N_2091,N_1950,N_1952);
or U2092 (N_2092,N_1986,N_1964);
nand U2093 (N_2093,N_1973,N_1907);
nor U2094 (N_2094,N_1937,N_1986);
and U2095 (N_2095,N_1927,N_1973);
and U2096 (N_2096,N_1974,N_1941);
xor U2097 (N_2097,N_1992,N_1909);
nor U2098 (N_2098,N_1910,N_1926);
and U2099 (N_2099,N_1948,N_1995);
nor U2100 (N_2100,N_2098,N_2078);
xor U2101 (N_2101,N_2050,N_2006);
or U2102 (N_2102,N_2099,N_2029);
or U2103 (N_2103,N_2091,N_2012);
and U2104 (N_2104,N_2003,N_2037);
nand U2105 (N_2105,N_2022,N_2008);
or U2106 (N_2106,N_2084,N_2020);
nand U2107 (N_2107,N_2025,N_2088);
or U2108 (N_2108,N_2036,N_2079);
and U2109 (N_2109,N_2009,N_2030);
nand U2110 (N_2110,N_2073,N_2062);
xnor U2111 (N_2111,N_2066,N_2061);
nand U2112 (N_2112,N_2089,N_2070);
nand U2113 (N_2113,N_2014,N_2064);
or U2114 (N_2114,N_2095,N_2004);
xor U2115 (N_2115,N_2018,N_2086);
xor U2116 (N_2116,N_2067,N_2000);
and U2117 (N_2117,N_2082,N_2041);
xnor U2118 (N_2118,N_2087,N_2026);
xnor U2119 (N_2119,N_2071,N_2074);
nor U2120 (N_2120,N_2063,N_2001);
nor U2121 (N_2121,N_2038,N_2068);
nor U2122 (N_2122,N_2054,N_2044);
nand U2123 (N_2123,N_2015,N_2072);
or U2124 (N_2124,N_2080,N_2057);
or U2125 (N_2125,N_2094,N_2065);
xnor U2126 (N_2126,N_2047,N_2093);
nor U2127 (N_2127,N_2051,N_2035);
and U2128 (N_2128,N_2021,N_2060);
nand U2129 (N_2129,N_2090,N_2027);
xor U2130 (N_2130,N_2045,N_2046);
nand U2131 (N_2131,N_2043,N_2011);
and U2132 (N_2132,N_2023,N_2059);
xnor U2133 (N_2133,N_2024,N_2081);
nor U2134 (N_2134,N_2048,N_2076);
nand U2135 (N_2135,N_2040,N_2069);
or U2136 (N_2136,N_2039,N_2058);
nand U2137 (N_2137,N_2056,N_2007);
nand U2138 (N_2138,N_2034,N_2052);
and U2139 (N_2139,N_2032,N_2010);
or U2140 (N_2140,N_2033,N_2085);
xnor U2141 (N_2141,N_2016,N_2019);
nand U2142 (N_2142,N_2042,N_2002);
nand U2143 (N_2143,N_2049,N_2053);
and U2144 (N_2144,N_2028,N_2096);
or U2145 (N_2145,N_2097,N_2013);
nand U2146 (N_2146,N_2092,N_2055);
and U2147 (N_2147,N_2017,N_2075);
and U2148 (N_2148,N_2005,N_2031);
nor U2149 (N_2149,N_2077,N_2083);
or U2150 (N_2150,N_2080,N_2028);
or U2151 (N_2151,N_2083,N_2071);
xnor U2152 (N_2152,N_2072,N_2053);
or U2153 (N_2153,N_2068,N_2059);
nand U2154 (N_2154,N_2026,N_2046);
and U2155 (N_2155,N_2023,N_2006);
nand U2156 (N_2156,N_2073,N_2093);
nand U2157 (N_2157,N_2001,N_2093);
nor U2158 (N_2158,N_2092,N_2063);
and U2159 (N_2159,N_2008,N_2046);
nor U2160 (N_2160,N_2034,N_2050);
nand U2161 (N_2161,N_2036,N_2037);
xor U2162 (N_2162,N_2022,N_2040);
nand U2163 (N_2163,N_2079,N_2072);
and U2164 (N_2164,N_2042,N_2045);
and U2165 (N_2165,N_2016,N_2025);
and U2166 (N_2166,N_2059,N_2004);
or U2167 (N_2167,N_2098,N_2031);
or U2168 (N_2168,N_2017,N_2078);
nor U2169 (N_2169,N_2021,N_2077);
and U2170 (N_2170,N_2099,N_2041);
xor U2171 (N_2171,N_2020,N_2019);
and U2172 (N_2172,N_2018,N_2090);
and U2173 (N_2173,N_2015,N_2024);
nand U2174 (N_2174,N_2091,N_2073);
xnor U2175 (N_2175,N_2008,N_2002);
xor U2176 (N_2176,N_2099,N_2015);
or U2177 (N_2177,N_2020,N_2065);
xnor U2178 (N_2178,N_2027,N_2056);
and U2179 (N_2179,N_2040,N_2018);
nand U2180 (N_2180,N_2076,N_2016);
nand U2181 (N_2181,N_2006,N_2062);
nor U2182 (N_2182,N_2090,N_2095);
nor U2183 (N_2183,N_2039,N_2003);
and U2184 (N_2184,N_2053,N_2052);
or U2185 (N_2185,N_2070,N_2031);
and U2186 (N_2186,N_2015,N_2023);
nor U2187 (N_2187,N_2057,N_2011);
or U2188 (N_2188,N_2049,N_2085);
xor U2189 (N_2189,N_2066,N_2062);
xor U2190 (N_2190,N_2085,N_2005);
and U2191 (N_2191,N_2038,N_2012);
xor U2192 (N_2192,N_2055,N_2037);
and U2193 (N_2193,N_2033,N_2076);
and U2194 (N_2194,N_2011,N_2064);
and U2195 (N_2195,N_2055,N_2091);
or U2196 (N_2196,N_2099,N_2079);
xnor U2197 (N_2197,N_2003,N_2048);
and U2198 (N_2198,N_2060,N_2052);
nand U2199 (N_2199,N_2067,N_2085);
xor U2200 (N_2200,N_2170,N_2189);
and U2201 (N_2201,N_2130,N_2111);
or U2202 (N_2202,N_2124,N_2192);
xor U2203 (N_2203,N_2107,N_2157);
nor U2204 (N_2204,N_2118,N_2167);
and U2205 (N_2205,N_2193,N_2135);
nor U2206 (N_2206,N_2142,N_2176);
nand U2207 (N_2207,N_2146,N_2132);
nor U2208 (N_2208,N_2128,N_2154);
nor U2209 (N_2209,N_2168,N_2123);
nor U2210 (N_2210,N_2110,N_2191);
nand U2211 (N_2211,N_2121,N_2115);
and U2212 (N_2212,N_2156,N_2108);
or U2213 (N_2213,N_2126,N_2180);
or U2214 (N_2214,N_2188,N_2194);
nor U2215 (N_2215,N_2158,N_2174);
xor U2216 (N_2216,N_2143,N_2114);
or U2217 (N_2217,N_2184,N_2177);
xnor U2218 (N_2218,N_2181,N_2100);
or U2219 (N_2219,N_2179,N_2183);
nor U2220 (N_2220,N_2187,N_2197);
and U2221 (N_2221,N_2185,N_2163);
nor U2222 (N_2222,N_2104,N_2148);
nor U2223 (N_2223,N_2139,N_2116);
nand U2224 (N_2224,N_2145,N_2186);
nand U2225 (N_2225,N_2131,N_2196);
nor U2226 (N_2226,N_2103,N_2166);
nor U2227 (N_2227,N_2117,N_2105);
or U2228 (N_2228,N_2106,N_2112);
or U2229 (N_2229,N_2164,N_2113);
and U2230 (N_2230,N_2129,N_2141);
xor U2231 (N_2231,N_2160,N_2195);
nor U2232 (N_2232,N_2125,N_2172);
xnor U2233 (N_2233,N_2173,N_2102);
nor U2234 (N_2234,N_2138,N_2147);
and U2235 (N_2235,N_2162,N_2198);
nand U2236 (N_2236,N_2149,N_2199);
nand U2237 (N_2237,N_2159,N_2161);
or U2238 (N_2238,N_2144,N_2178);
and U2239 (N_2239,N_2150,N_2140);
nand U2240 (N_2240,N_2137,N_2136);
or U2241 (N_2241,N_2122,N_2165);
nand U2242 (N_2242,N_2120,N_2109);
nor U2243 (N_2243,N_2153,N_2169);
or U2244 (N_2244,N_2171,N_2152);
nand U2245 (N_2245,N_2101,N_2190);
nor U2246 (N_2246,N_2182,N_2134);
xnor U2247 (N_2247,N_2133,N_2151);
xnor U2248 (N_2248,N_2175,N_2155);
nand U2249 (N_2249,N_2127,N_2119);
nor U2250 (N_2250,N_2185,N_2166);
nor U2251 (N_2251,N_2115,N_2170);
xnor U2252 (N_2252,N_2179,N_2134);
and U2253 (N_2253,N_2132,N_2141);
xor U2254 (N_2254,N_2165,N_2150);
nor U2255 (N_2255,N_2156,N_2111);
xor U2256 (N_2256,N_2111,N_2128);
and U2257 (N_2257,N_2131,N_2152);
nand U2258 (N_2258,N_2121,N_2128);
xnor U2259 (N_2259,N_2198,N_2178);
and U2260 (N_2260,N_2132,N_2163);
and U2261 (N_2261,N_2158,N_2157);
xor U2262 (N_2262,N_2169,N_2127);
nand U2263 (N_2263,N_2159,N_2171);
nor U2264 (N_2264,N_2199,N_2168);
and U2265 (N_2265,N_2184,N_2138);
or U2266 (N_2266,N_2145,N_2166);
and U2267 (N_2267,N_2132,N_2166);
nand U2268 (N_2268,N_2131,N_2112);
xnor U2269 (N_2269,N_2139,N_2181);
xor U2270 (N_2270,N_2123,N_2139);
xnor U2271 (N_2271,N_2164,N_2197);
nor U2272 (N_2272,N_2165,N_2177);
nor U2273 (N_2273,N_2114,N_2158);
and U2274 (N_2274,N_2135,N_2180);
or U2275 (N_2275,N_2131,N_2120);
or U2276 (N_2276,N_2180,N_2148);
nand U2277 (N_2277,N_2161,N_2189);
nor U2278 (N_2278,N_2149,N_2153);
or U2279 (N_2279,N_2111,N_2163);
or U2280 (N_2280,N_2137,N_2154);
or U2281 (N_2281,N_2143,N_2111);
and U2282 (N_2282,N_2192,N_2101);
nor U2283 (N_2283,N_2157,N_2176);
xnor U2284 (N_2284,N_2150,N_2136);
xor U2285 (N_2285,N_2174,N_2198);
nand U2286 (N_2286,N_2120,N_2148);
nor U2287 (N_2287,N_2156,N_2110);
or U2288 (N_2288,N_2113,N_2178);
nor U2289 (N_2289,N_2156,N_2135);
and U2290 (N_2290,N_2103,N_2184);
nand U2291 (N_2291,N_2160,N_2142);
nor U2292 (N_2292,N_2110,N_2147);
nand U2293 (N_2293,N_2144,N_2171);
xor U2294 (N_2294,N_2123,N_2162);
and U2295 (N_2295,N_2113,N_2183);
xor U2296 (N_2296,N_2174,N_2166);
and U2297 (N_2297,N_2142,N_2182);
nor U2298 (N_2298,N_2197,N_2172);
and U2299 (N_2299,N_2156,N_2114);
nor U2300 (N_2300,N_2233,N_2241);
or U2301 (N_2301,N_2260,N_2204);
or U2302 (N_2302,N_2253,N_2259);
nor U2303 (N_2303,N_2208,N_2254);
xor U2304 (N_2304,N_2215,N_2210);
nor U2305 (N_2305,N_2263,N_2224);
or U2306 (N_2306,N_2202,N_2283);
nand U2307 (N_2307,N_2250,N_2279);
or U2308 (N_2308,N_2217,N_2205);
nand U2309 (N_2309,N_2247,N_2272);
nor U2310 (N_2310,N_2232,N_2293);
nand U2311 (N_2311,N_2256,N_2221);
nor U2312 (N_2312,N_2223,N_2258);
or U2313 (N_2313,N_2284,N_2248);
nor U2314 (N_2314,N_2238,N_2280);
or U2315 (N_2315,N_2207,N_2214);
nand U2316 (N_2316,N_2206,N_2255);
or U2317 (N_2317,N_2296,N_2235);
nor U2318 (N_2318,N_2228,N_2230);
and U2319 (N_2319,N_2229,N_2286);
or U2320 (N_2320,N_2264,N_2294);
nand U2321 (N_2321,N_2287,N_2242);
nor U2322 (N_2322,N_2265,N_2225);
xnor U2323 (N_2323,N_2244,N_2281);
nand U2324 (N_2324,N_2236,N_2220);
xnor U2325 (N_2325,N_2252,N_2222);
and U2326 (N_2326,N_2274,N_2227);
nor U2327 (N_2327,N_2285,N_2275);
and U2328 (N_2328,N_2231,N_2212);
nand U2329 (N_2329,N_2267,N_2237);
nand U2330 (N_2330,N_2269,N_2209);
or U2331 (N_2331,N_2201,N_2270);
nand U2332 (N_2332,N_2203,N_2200);
xnor U2333 (N_2333,N_2262,N_2234);
and U2334 (N_2334,N_2216,N_2251);
and U2335 (N_2335,N_2245,N_2276);
nand U2336 (N_2336,N_2213,N_2211);
nor U2337 (N_2337,N_2288,N_2271);
or U2338 (N_2338,N_2249,N_2243);
nand U2339 (N_2339,N_2261,N_2297);
xnor U2340 (N_2340,N_2273,N_2290);
nor U2341 (N_2341,N_2218,N_2289);
and U2342 (N_2342,N_2291,N_2295);
xor U2343 (N_2343,N_2292,N_2299);
nor U2344 (N_2344,N_2266,N_2277);
xor U2345 (N_2345,N_2239,N_2226);
nand U2346 (N_2346,N_2268,N_2282);
xnor U2347 (N_2347,N_2298,N_2219);
and U2348 (N_2348,N_2240,N_2246);
nand U2349 (N_2349,N_2278,N_2257);
nor U2350 (N_2350,N_2251,N_2227);
nor U2351 (N_2351,N_2236,N_2234);
and U2352 (N_2352,N_2219,N_2226);
nor U2353 (N_2353,N_2271,N_2216);
and U2354 (N_2354,N_2219,N_2293);
nor U2355 (N_2355,N_2251,N_2267);
or U2356 (N_2356,N_2238,N_2262);
or U2357 (N_2357,N_2203,N_2292);
nor U2358 (N_2358,N_2224,N_2211);
and U2359 (N_2359,N_2281,N_2291);
xnor U2360 (N_2360,N_2255,N_2238);
and U2361 (N_2361,N_2248,N_2226);
or U2362 (N_2362,N_2261,N_2236);
nor U2363 (N_2363,N_2261,N_2249);
nand U2364 (N_2364,N_2266,N_2250);
nand U2365 (N_2365,N_2207,N_2212);
or U2366 (N_2366,N_2250,N_2247);
and U2367 (N_2367,N_2298,N_2210);
or U2368 (N_2368,N_2264,N_2283);
and U2369 (N_2369,N_2237,N_2249);
nand U2370 (N_2370,N_2244,N_2295);
nor U2371 (N_2371,N_2207,N_2256);
and U2372 (N_2372,N_2239,N_2244);
nor U2373 (N_2373,N_2273,N_2267);
xnor U2374 (N_2374,N_2212,N_2213);
and U2375 (N_2375,N_2293,N_2226);
or U2376 (N_2376,N_2229,N_2239);
nand U2377 (N_2377,N_2215,N_2285);
and U2378 (N_2378,N_2269,N_2223);
xor U2379 (N_2379,N_2203,N_2238);
nand U2380 (N_2380,N_2217,N_2222);
and U2381 (N_2381,N_2273,N_2278);
or U2382 (N_2382,N_2298,N_2274);
or U2383 (N_2383,N_2234,N_2284);
xor U2384 (N_2384,N_2227,N_2299);
xor U2385 (N_2385,N_2240,N_2261);
nor U2386 (N_2386,N_2250,N_2291);
nand U2387 (N_2387,N_2266,N_2239);
nand U2388 (N_2388,N_2226,N_2289);
and U2389 (N_2389,N_2208,N_2266);
and U2390 (N_2390,N_2219,N_2276);
and U2391 (N_2391,N_2228,N_2213);
xnor U2392 (N_2392,N_2240,N_2278);
nand U2393 (N_2393,N_2293,N_2274);
nor U2394 (N_2394,N_2277,N_2206);
or U2395 (N_2395,N_2267,N_2293);
xor U2396 (N_2396,N_2253,N_2201);
xor U2397 (N_2397,N_2299,N_2206);
nand U2398 (N_2398,N_2239,N_2221);
nor U2399 (N_2399,N_2244,N_2269);
or U2400 (N_2400,N_2387,N_2340);
nand U2401 (N_2401,N_2308,N_2369);
nor U2402 (N_2402,N_2327,N_2304);
xnor U2403 (N_2403,N_2307,N_2311);
nor U2404 (N_2404,N_2386,N_2362);
or U2405 (N_2405,N_2350,N_2383);
nor U2406 (N_2406,N_2336,N_2352);
xnor U2407 (N_2407,N_2345,N_2329);
nand U2408 (N_2408,N_2391,N_2314);
xnor U2409 (N_2409,N_2343,N_2380);
nor U2410 (N_2410,N_2357,N_2339);
nor U2411 (N_2411,N_2319,N_2384);
or U2412 (N_2412,N_2334,N_2381);
xor U2413 (N_2413,N_2375,N_2302);
or U2414 (N_2414,N_2330,N_2373);
or U2415 (N_2415,N_2398,N_2365);
xnor U2416 (N_2416,N_2363,N_2360);
xor U2417 (N_2417,N_2315,N_2359);
nor U2418 (N_2418,N_2342,N_2349);
or U2419 (N_2419,N_2301,N_2300);
nand U2420 (N_2420,N_2379,N_2367);
or U2421 (N_2421,N_2346,N_2399);
xnor U2422 (N_2422,N_2323,N_2356);
xor U2423 (N_2423,N_2341,N_2344);
or U2424 (N_2424,N_2320,N_2348);
or U2425 (N_2425,N_2306,N_2309);
nor U2426 (N_2426,N_2332,N_2355);
or U2427 (N_2427,N_2376,N_2325);
nand U2428 (N_2428,N_2366,N_2353);
and U2429 (N_2429,N_2358,N_2371);
and U2430 (N_2430,N_2382,N_2338);
nor U2431 (N_2431,N_2374,N_2368);
and U2432 (N_2432,N_2394,N_2390);
nand U2433 (N_2433,N_2397,N_2335);
and U2434 (N_2434,N_2326,N_2396);
nor U2435 (N_2435,N_2305,N_2388);
nand U2436 (N_2436,N_2393,N_2303);
xnor U2437 (N_2437,N_2372,N_2317);
nand U2438 (N_2438,N_2312,N_2316);
nand U2439 (N_2439,N_2318,N_2364);
or U2440 (N_2440,N_2347,N_2310);
and U2441 (N_2441,N_2354,N_2377);
and U2442 (N_2442,N_2333,N_2331);
nand U2443 (N_2443,N_2324,N_2322);
nand U2444 (N_2444,N_2321,N_2351);
or U2445 (N_2445,N_2337,N_2370);
xor U2446 (N_2446,N_2389,N_2378);
nor U2447 (N_2447,N_2313,N_2385);
and U2448 (N_2448,N_2392,N_2328);
or U2449 (N_2449,N_2395,N_2361);
and U2450 (N_2450,N_2397,N_2332);
nand U2451 (N_2451,N_2338,N_2374);
nand U2452 (N_2452,N_2373,N_2319);
nor U2453 (N_2453,N_2324,N_2315);
or U2454 (N_2454,N_2382,N_2396);
and U2455 (N_2455,N_2355,N_2376);
nand U2456 (N_2456,N_2363,N_2311);
and U2457 (N_2457,N_2385,N_2389);
nor U2458 (N_2458,N_2365,N_2333);
or U2459 (N_2459,N_2342,N_2328);
and U2460 (N_2460,N_2314,N_2345);
and U2461 (N_2461,N_2313,N_2306);
and U2462 (N_2462,N_2305,N_2367);
or U2463 (N_2463,N_2325,N_2300);
and U2464 (N_2464,N_2310,N_2372);
nor U2465 (N_2465,N_2351,N_2389);
and U2466 (N_2466,N_2380,N_2356);
nand U2467 (N_2467,N_2376,N_2371);
xor U2468 (N_2468,N_2306,N_2321);
nor U2469 (N_2469,N_2387,N_2396);
and U2470 (N_2470,N_2342,N_2355);
nor U2471 (N_2471,N_2367,N_2301);
xnor U2472 (N_2472,N_2334,N_2319);
and U2473 (N_2473,N_2382,N_2304);
xor U2474 (N_2474,N_2305,N_2322);
and U2475 (N_2475,N_2317,N_2381);
nand U2476 (N_2476,N_2331,N_2323);
nor U2477 (N_2477,N_2333,N_2344);
xnor U2478 (N_2478,N_2367,N_2342);
or U2479 (N_2479,N_2366,N_2391);
xor U2480 (N_2480,N_2399,N_2378);
nor U2481 (N_2481,N_2312,N_2363);
nor U2482 (N_2482,N_2329,N_2307);
nand U2483 (N_2483,N_2310,N_2375);
or U2484 (N_2484,N_2384,N_2333);
nor U2485 (N_2485,N_2392,N_2336);
nand U2486 (N_2486,N_2304,N_2384);
or U2487 (N_2487,N_2370,N_2324);
nor U2488 (N_2488,N_2305,N_2390);
and U2489 (N_2489,N_2321,N_2382);
xor U2490 (N_2490,N_2333,N_2328);
xnor U2491 (N_2491,N_2301,N_2340);
or U2492 (N_2492,N_2370,N_2300);
nand U2493 (N_2493,N_2383,N_2316);
and U2494 (N_2494,N_2376,N_2309);
nand U2495 (N_2495,N_2322,N_2389);
or U2496 (N_2496,N_2307,N_2303);
or U2497 (N_2497,N_2380,N_2310);
xor U2498 (N_2498,N_2380,N_2325);
xnor U2499 (N_2499,N_2333,N_2360);
nor U2500 (N_2500,N_2488,N_2495);
and U2501 (N_2501,N_2412,N_2445);
and U2502 (N_2502,N_2408,N_2460);
and U2503 (N_2503,N_2400,N_2465);
and U2504 (N_2504,N_2406,N_2477);
and U2505 (N_2505,N_2455,N_2416);
nand U2506 (N_2506,N_2422,N_2437);
or U2507 (N_2507,N_2411,N_2403);
and U2508 (N_2508,N_2446,N_2438);
or U2509 (N_2509,N_2410,N_2458);
or U2510 (N_2510,N_2496,N_2407);
nand U2511 (N_2511,N_2467,N_2472);
xor U2512 (N_2512,N_2466,N_2491);
nor U2513 (N_2513,N_2469,N_2441);
and U2514 (N_2514,N_2413,N_2476);
xor U2515 (N_2515,N_2401,N_2485);
xor U2516 (N_2516,N_2490,N_2484);
and U2517 (N_2517,N_2417,N_2447);
or U2518 (N_2518,N_2402,N_2474);
nand U2519 (N_2519,N_2481,N_2498);
nor U2520 (N_2520,N_2448,N_2425);
nand U2521 (N_2521,N_2486,N_2420);
nor U2522 (N_2522,N_2449,N_2463);
xnor U2523 (N_2523,N_2475,N_2461);
xnor U2524 (N_2524,N_2473,N_2433);
xor U2525 (N_2525,N_2418,N_2409);
xor U2526 (N_2526,N_2497,N_2487);
or U2527 (N_2527,N_2444,N_2483);
xnor U2528 (N_2528,N_2430,N_2462);
nand U2529 (N_2529,N_2454,N_2482);
and U2530 (N_2530,N_2478,N_2489);
and U2531 (N_2531,N_2493,N_2499);
nand U2532 (N_2532,N_2450,N_2414);
nand U2533 (N_2533,N_2431,N_2443);
nand U2534 (N_2534,N_2451,N_2405);
nand U2535 (N_2535,N_2494,N_2442);
nand U2536 (N_2536,N_2464,N_2468);
nand U2537 (N_2537,N_2426,N_2457);
xor U2538 (N_2538,N_2453,N_2427);
nand U2539 (N_2539,N_2415,N_2459);
xnor U2540 (N_2540,N_2492,N_2439);
nor U2541 (N_2541,N_2424,N_2423);
nand U2542 (N_2542,N_2404,N_2419);
nand U2543 (N_2543,N_2434,N_2421);
nor U2544 (N_2544,N_2428,N_2429);
or U2545 (N_2545,N_2435,N_2432);
xnor U2546 (N_2546,N_2471,N_2456);
nand U2547 (N_2547,N_2480,N_2452);
nand U2548 (N_2548,N_2479,N_2436);
or U2549 (N_2549,N_2470,N_2440);
xnor U2550 (N_2550,N_2456,N_2405);
nor U2551 (N_2551,N_2420,N_2446);
or U2552 (N_2552,N_2444,N_2487);
nand U2553 (N_2553,N_2442,N_2481);
nor U2554 (N_2554,N_2470,N_2401);
nand U2555 (N_2555,N_2487,N_2421);
nand U2556 (N_2556,N_2489,N_2410);
nor U2557 (N_2557,N_2472,N_2419);
and U2558 (N_2558,N_2460,N_2493);
nor U2559 (N_2559,N_2442,N_2466);
nand U2560 (N_2560,N_2440,N_2468);
xor U2561 (N_2561,N_2490,N_2428);
nand U2562 (N_2562,N_2452,N_2431);
nor U2563 (N_2563,N_2459,N_2414);
nor U2564 (N_2564,N_2459,N_2455);
or U2565 (N_2565,N_2466,N_2496);
nand U2566 (N_2566,N_2448,N_2482);
and U2567 (N_2567,N_2443,N_2482);
xor U2568 (N_2568,N_2481,N_2405);
nor U2569 (N_2569,N_2458,N_2418);
nand U2570 (N_2570,N_2448,N_2451);
and U2571 (N_2571,N_2431,N_2457);
xnor U2572 (N_2572,N_2448,N_2424);
nand U2573 (N_2573,N_2436,N_2452);
and U2574 (N_2574,N_2447,N_2436);
or U2575 (N_2575,N_2471,N_2447);
nand U2576 (N_2576,N_2428,N_2459);
and U2577 (N_2577,N_2472,N_2483);
and U2578 (N_2578,N_2425,N_2446);
or U2579 (N_2579,N_2433,N_2425);
xor U2580 (N_2580,N_2425,N_2404);
nor U2581 (N_2581,N_2452,N_2447);
nand U2582 (N_2582,N_2477,N_2400);
or U2583 (N_2583,N_2479,N_2488);
xnor U2584 (N_2584,N_2490,N_2483);
nand U2585 (N_2585,N_2476,N_2493);
nor U2586 (N_2586,N_2498,N_2495);
nor U2587 (N_2587,N_2455,N_2456);
and U2588 (N_2588,N_2471,N_2479);
nor U2589 (N_2589,N_2453,N_2408);
nand U2590 (N_2590,N_2484,N_2461);
nor U2591 (N_2591,N_2486,N_2432);
nand U2592 (N_2592,N_2400,N_2460);
nand U2593 (N_2593,N_2494,N_2479);
nor U2594 (N_2594,N_2428,N_2434);
or U2595 (N_2595,N_2464,N_2478);
or U2596 (N_2596,N_2426,N_2427);
xnor U2597 (N_2597,N_2477,N_2428);
xor U2598 (N_2598,N_2423,N_2498);
nor U2599 (N_2599,N_2473,N_2435);
xnor U2600 (N_2600,N_2504,N_2502);
or U2601 (N_2601,N_2541,N_2558);
xor U2602 (N_2602,N_2578,N_2545);
and U2603 (N_2603,N_2533,N_2573);
xor U2604 (N_2604,N_2569,N_2508);
nand U2605 (N_2605,N_2572,N_2581);
nor U2606 (N_2606,N_2597,N_2537);
nor U2607 (N_2607,N_2554,N_2568);
nand U2608 (N_2608,N_2565,N_2593);
or U2609 (N_2609,N_2548,N_2539);
nand U2610 (N_2610,N_2589,N_2510);
nor U2611 (N_2611,N_2531,N_2560);
or U2612 (N_2612,N_2575,N_2579);
and U2613 (N_2613,N_2574,N_2566);
nand U2614 (N_2614,N_2535,N_2523);
xnor U2615 (N_2615,N_2598,N_2529);
nor U2616 (N_2616,N_2519,N_2577);
and U2617 (N_2617,N_2570,N_2564);
nor U2618 (N_2618,N_2592,N_2596);
and U2619 (N_2619,N_2513,N_2524);
nand U2620 (N_2620,N_2542,N_2516);
nand U2621 (N_2621,N_2571,N_2520);
nand U2622 (N_2622,N_2595,N_2522);
or U2623 (N_2623,N_2587,N_2546);
and U2624 (N_2624,N_2549,N_2521);
xnor U2625 (N_2625,N_2538,N_2530);
nand U2626 (N_2626,N_2576,N_2547);
nor U2627 (N_2627,N_2526,N_2507);
nor U2628 (N_2628,N_2584,N_2559);
and U2629 (N_2629,N_2511,N_2525);
xor U2630 (N_2630,N_2553,N_2591);
nand U2631 (N_2631,N_2599,N_2563);
and U2632 (N_2632,N_2580,N_2582);
nor U2633 (N_2633,N_2567,N_2551);
nand U2634 (N_2634,N_2544,N_2534);
or U2635 (N_2635,N_2583,N_2588);
nor U2636 (N_2636,N_2586,N_2512);
nand U2637 (N_2637,N_2506,N_2552);
nand U2638 (N_2638,N_2515,N_2505);
nand U2639 (N_2639,N_2532,N_2543);
nand U2640 (N_2640,N_2527,N_2503);
nand U2641 (N_2641,N_2590,N_2500);
or U2642 (N_2642,N_2561,N_2540);
nor U2643 (N_2643,N_2501,N_2509);
and U2644 (N_2644,N_2585,N_2514);
nand U2645 (N_2645,N_2557,N_2562);
and U2646 (N_2646,N_2594,N_2550);
nand U2647 (N_2647,N_2536,N_2528);
or U2648 (N_2648,N_2518,N_2517);
and U2649 (N_2649,N_2556,N_2555);
xor U2650 (N_2650,N_2590,N_2592);
nor U2651 (N_2651,N_2560,N_2579);
nor U2652 (N_2652,N_2542,N_2560);
nand U2653 (N_2653,N_2510,N_2597);
nand U2654 (N_2654,N_2568,N_2580);
and U2655 (N_2655,N_2533,N_2503);
nor U2656 (N_2656,N_2549,N_2511);
nand U2657 (N_2657,N_2559,N_2568);
nor U2658 (N_2658,N_2588,N_2566);
and U2659 (N_2659,N_2597,N_2593);
nand U2660 (N_2660,N_2531,N_2587);
or U2661 (N_2661,N_2536,N_2533);
and U2662 (N_2662,N_2588,N_2596);
nand U2663 (N_2663,N_2584,N_2582);
nor U2664 (N_2664,N_2542,N_2531);
or U2665 (N_2665,N_2504,N_2541);
nor U2666 (N_2666,N_2589,N_2522);
and U2667 (N_2667,N_2568,N_2519);
nand U2668 (N_2668,N_2531,N_2569);
nor U2669 (N_2669,N_2514,N_2562);
xor U2670 (N_2670,N_2545,N_2513);
nand U2671 (N_2671,N_2561,N_2575);
nand U2672 (N_2672,N_2584,N_2523);
nand U2673 (N_2673,N_2538,N_2594);
nand U2674 (N_2674,N_2502,N_2585);
nor U2675 (N_2675,N_2568,N_2567);
nor U2676 (N_2676,N_2535,N_2517);
nor U2677 (N_2677,N_2532,N_2563);
nand U2678 (N_2678,N_2545,N_2555);
nand U2679 (N_2679,N_2516,N_2584);
xor U2680 (N_2680,N_2587,N_2563);
nor U2681 (N_2681,N_2572,N_2526);
nor U2682 (N_2682,N_2599,N_2521);
xnor U2683 (N_2683,N_2526,N_2520);
or U2684 (N_2684,N_2547,N_2532);
nand U2685 (N_2685,N_2578,N_2532);
and U2686 (N_2686,N_2506,N_2502);
xor U2687 (N_2687,N_2539,N_2575);
nor U2688 (N_2688,N_2578,N_2561);
nand U2689 (N_2689,N_2517,N_2512);
nand U2690 (N_2690,N_2569,N_2518);
xor U2691 (N_2691,N_2588,N_2569);
nor U2692 (N_2692,N_2578,N_2570);
and U2693 (N_2693,N_2540,N_2523);
nor U2694 (N_2694,N_2514,N_2584);
or U2695 (N_2695,N_2502,N_2567);
nand U2696 (N_2696,N_2599,N_2551);
nor U2697 (N_2697,N_2517,N_2573);
nor U2698 (N_2698,N_2521,N_2509);
nor U2699 (N_2699,N_2513,N_2549);
nor U2700 (N_2700,N_2637,N_2684);
xor U2701 (N_2701,N_2636,N_2697);
xnor U2702 (N_2702,N_2631,N_2622);
and U2703 (N_2703,N_2604,N_2640);
nor U2704 (N_2704,N_2625,N_2687);
or U2705 (N_2705,N_2693,N_2668);
xor U2706 (N_2706,N_2662,N_2629);
xnor U2707 (N_2707,N_2603,N_2614);
nand U2708 (N_2708,N_2674,N_2671);
xor U2709 (N_2709,N_2689,N_2649);
nand U2710 (N_2710,N_2665,N_2619);
and U2711 (N_2711,N_2663,N_2677);
nand U2712 (N_2712,N_2606,N_2611);
or U2713 (N_2713,N_2676,N_2659);
nand U2714 (N_2714,N_2630,N_2688);
nand U2715 (N_2715,N_2681,N_2673);
nand U2716 (N_2716,N_2610,N_2605);
xor U2717 (N_2717,N_2645,N_2618);
nand U2718 (N_2718,N_2638,N_2691);
nor U2719 (N_2719,N_2639,N_2621);
or U2720 (N_2720,N_2602,N_2682);
xnor U2721 (N_2721,N_2613,N_2634);
nand U2722 (N_2722,N_2664,N_2623);
xnor U2723 (N_2723,N_2657,N_2648);
and U2724 (N_2724,N_2695,N_2694);
nor U2725 (N_2725,N_2652,N_2685);
xnor U2726 (N_2726,N_2643,N_2655);
nand U2727 (N_2727,N_2680,N_2658);
nand U2728 (N_2728,N_2612,N_2690);
and U2729 (N_2729,N_2609,N_2666);
and U2730 (N_2730,N_2620,N_2683);
xor U2731 (N_2731,N_2650,N_2651);
or U2732 (N_2732,N_2646,N_2632);
and U2733 (N_2733,N_2692,N_2686);
xor U2734 (N_2734,N_2669,N_2672);
xor U2735 (N_2735,N_2616,N_2653);
or U2736 (N_2736,N_2627,N_2661);
nand U2737 (N_2737,N_2641,N_2607);
nand U2738 (N_2738,N_2656,N_2654);
nor U2739 (N_2739,N_2678,N_2600);
xnor U2740 (N_2740,N_2626,N_2635);
nor U2741 (N_2741,N_2617,N_2667);
and U2742 (N_2742,N_2628,N_2647);
nand U2743 (N_2743,N_2679,N_2699);
nor U2744 (N_2744,N_2675,N_2642);
or U2745 (N_2745,N_2608,N_2633);
and U2746 (N_2746,N_2696,N_2601);
nand U2747 (N_2747,N_2624,N_2698);
nand U2748 (N_2748,N_2615,N_2660);
xnor U2749 (N_2749,N_2670,N_2644);
or U2750 (N_2750,N_2687,N_2609);
nor U2751 (N_2751,N_2696,N_2610);
nor U2752 (N_2752,N_2611,N_2625);
nand U2753 (N_2753,N_2609,N_2623);
nor U2754 (N_2754,N_2690,N_2650);
nand U2755 (N_2755,N_2648,N_2667);
nand U2756 (N_2756,N_2622,N_2600);
nor U2757 (N_2757,N_2697,N_2604);
xor U2758 (N_2758,N_2643,N_2622);
or U2759 (N_2759,N_2632,N_2600);
xnor U2760 (N_2760,N_2611,N_2605);
or U2761 (N_2761,N_2643,N_2621);
nand U2762 (N_2762,N_2630,N_2634);
nor U2763 (N_2763,N_2646,N_2612);
xor U2764 (N_2764,N_2623,N_2607);
nand U2765 (N_2765,N_2698,N_2678);
nor U2766 (N_2766,N_2663,N_2639);
nor U2767 (N_2767,N_2627,N_2613);
and U2768 (N_2768,N_2696,N_2603);
xnor U2769 (N_2769,N_2646,N_2625);
nand U2770 (N_2770,N_2629,N_2604);
xor U2771 (N_2771,N_2612,N_2637);
nand U2772 (N_2772,N_2601,N_2697);
and U2773 (N_2773,N_2607,N_2678);
xnor U2774 (N_2774,N_2692,N_2620);
nand U2775 (N_2775,N_2680,N_2670);
or U2776 (N_2776,N_2672,N_2630);
nand U2777 (N_2777,N_2602,N_2639);
xor U2778 (N_2778,N_2686,N_2626);
nand U2779 (N_2779,N_2660,N_2616);
or U2780 (N_2780,N_2622,N_2680);
nand U2781 (N_2781,N_2633,N_2635);
and U2782 (N_2782,N_2628,N_2698);
nor U2783 (N_2783,N_2629,N_2600);
nor U2784 (N_2784,N_2665,N_2647);
xor U2785 (N_2785,N_2612,N_2683);
or U2786 (N_2786,N_2629,N_2646);
and U2787 (N_2787,N_2635,N_2675);
nand U2788 (N_2788,N_2699,N_2687);
or U2789 (N_2789,N_2615,N_2682);
nand U2790 (N_2790,N_2680,N_2601);
xnor U2791 (N_2791,N_2616,N_2664);
or U2792 (N_2792,N_2629,N_2697);
and U2793 (N_2793,N_2694,N_2657);
nand U2794 (N_2794,N_2644,N_2698);
nand U2795 (N_2795,N_2623,N_2669);
or U2796 (N_2796,N_2686,N_2638);
nor U2797 (N_2797,N_2629,N_2628);
xnor U2798 (N_2798,N_2681,N_2695);
or U2799 (N_2799,N_2672,N_2645);
and U2800 (N_2800,N_2717,N_2738);
and U2801 (N_2801,N_2760,N_2700);
or U2802 (N_2802,N_2736,N_2750);
and U2803 (N_2803,N_2724,N_2777);
nor U2804 (N_2804,N_2749,N_2723);
nand U2805 (N_2805,N_2711,N_2798);
and U2806 (N_2806,N_2752,N_2747);
nor U2807 (N_2807,N_2794,N_2734);
and U2808 (N_2808,N_2789,N_2708);
or U2809 (N_2809,N_2709,N_2786);
and U2810 (N_2810,N_2725,N_2742);
and U2811 (N_2811,N_2737,N_2722);
and U2812 (N_2812,N_2755,N_2799);
or U2813 (N_2813,N_2727,N_2705);
xor U2814 (N_2814,N_2767,N_2769);
and U2815 (N_2815,N_2772,N_2771);
and U2816 (N_2816,N_2729,N_2721);
xor U2817 (N_2817,N_2781,N_2710);
or U2818 (N_2818,N_2714,N_2785);
nor U2819 (N_2819,N_2707,N_2741);
xor U2820 (N_2820,N_2715,N_2762);
xor U2821 (N_2821,N_2743,N_2788);
nand U2822 (N_2822,N_2766,N_2764);
or U2823 (N_2823,N_2735,N_2745);
and U2824 (N_2824,N_2701,N_2779);
nand U2825 (N_2825,N_2702,N_2751);
nand U2826 (N_2826,N_2719,N_2775);
or U2827 (N_2827,N_2739,N_2763);
or U2828 (N_2828,N_2778,N_2773);
and U2829 (N_2829,N_2780,N_2792);
and U2830 (N_2830,N_2754,N_2761);
nand U2831 (N_2831,N_2758,N_2706);
nand U2832 (N_2832,N_2703,N_2759);
nor U2833 (N_2833,N_2740,N_2753);
or U2834 (N_2834,N_2765,N_2796);
nor U2835 (N_2835,N_2712,N_2720);
or U2836 (N_2836,N_2768,N_2776);
or U2837 (N_2837,N_2784,N_2731);
xor U2838 (N_2838,N_2748,N_2791);
nand U2839 (N_2839,N_2746,N_2782);
nor U2840 (N_2840,N_2756,N_2770);
or U2841 (N_2841,N_2732,N_2718);
or U2842 (N_2842,N_2726,N_2793);
nand U2843 (N_2843,N_2730,N_2797);
and U2844 (N_2844,N_2783,N_2716);
xor U2845 (N_2845,N_2744,N_2704);
xnor U2846 (N_2846,N_2733,N_2774);
or U2847 (N_2847,N_2790,N_2713);
and U2848 (N_2848,N_2757,N_2728);
nand U2849 (N_2849,N_2795,N_2787);
or U2850 (N_2850,N_2761,N_2790);
or U2851 (N_2851,N_2773,N_2734);
nor U2852 (N_2852,N_2779,N_2714);
nor U2853 (N_2853,N_2703,N_2710);
or U2854 (N_2854,N_2784,N_2725);
nor U2855 (N_2855,N_2754,N_2751);
and U2856 (N_2856,N_2720,N_2792);
nand U2857 (N_2857,N_2767,N_2703);
nand U2858 (N_2858,N_2798,N_2704);
xnor U2859 (N_2859,N_2746,N_2711);
nand U2860 (N_2860,N_2779,N_2722);
nand U2861 (N_2861,N_2717,N_2795);
and U2862 (N_2862,N_2737,N_2796);
or U2863 (N_2863,N_2787,N_2773);
nor U2864 (N_2864,N_2740,N_2793);
or U2865 (N_2865,N_2796,N_2744);
or U2866 (N_2866,N_2730,N_2716);
nand U2867 (N_2867,N_2728,N_2786);
xnor U2868 (N_2868,N_2758,N_2753);
xor U2869 (N_2869,N_2730,N_2710);
xor U2870 (N_2870,N_2702,N_2769);
nor U2871 (N_2871,N_2740,N_2780);
nand U2872 (N_2872,N_2718,N_2705);
nor U2873 (N_2873,N_2706,N_2775);
or U2874 (N_2874,N_2766,N_2701);
nor U2875 (N_2875,N_2722,N_2700);
xnor U2876 (N_2876,N_2723,N_2796);
or U2877 (N_2877,N_2702,N_2729);
xor U2878 (N_2878,N_2793,N_2730);
xor U2879 (N_2879,N_2742,N_2762);
or U2880 (N_2880,N_2742,N_2798);
and U2881 (N_2881,N_2757,N_2755);
or U2882 (N_2882,N_2753,N_2732);
nand U2883 (N_2883,N_2792,N_2718);
and U2884 (N_2884,N_2741,N_2703);
or U2885 (N_2885,N_2792,N_2753);
xor U2886 (N_2886,N_2730,N_2707);
xor U2887 (N_2887,N_2714,N_2798);
nor U2888 (N_2888,N_2758,N_2748);
xor U2889 (N_2889,N_2772,N_2763);
or U2890 (N_2890,N_2727,N_2740);
nand U2891 (N_2891,N_2759,N_2773);
nor U2892 (N_2892,N_2755,N_2722);
xor U2893 (N_2893,N_2754,N_2741);
and U2894 (N_2894,N_2729,N_2769);
nor U2895 (N_2895,N_2773,N_2707);
nand U2896 (N_2896,N_2721,N_2775);
nor U2897 (N_2897,N_2776,N_2730);
or U2898 (N_2898,N_2727,N_2776);
or U2899 (N_2899,N_2749,N_2740);
xnor U2900 (N_2900,N_2877,N_2896);
nand U2901 (N_2901,N_2866,N_2876);
and U2902 (N_2902,N_2881,N_2887);
and U2903 (N_2903,N_2847,N_2818);
and U2904 (N_2904,N_2875,N_2823);
xor U2905 (N_2905,N_2848,N_2800);
nor U2906 (N_2906,N_2849,N_2822);
nand U2907 (N_2907,N_2825,N_2809);
and U2908 (N_2908,N_2826,N_2840);
or U2909 (N_2909,N_2839,N_2846);
and U2910 (N_2910,N_2869,N_2804);
or U2911 (N_2911,N_2855,N_2835);
nor U2912 (N_2912,N_2864,N_2891);
and U2913 (N_2913,N_2874,N_2817);
nor U2914 (N_2914,N_2850,N_2859);
nor U2915 (N_2915,N_2813,N_2808);
nand U2916 (N_2916,N_2888,N_2851);
nand U2917 (N_2917,N_2811,N_2838);
nor U2918 (N_2918,N_2815,N_2820);
xnor U2919 (N_2919,N_2878,N_2897);
nand U2920 (N_2920,N_2833,N_2803);
or U2921 (N_2921,N_2858,N_2895);
nor U2922 (N_2922,N_2883,N_2837);
and U2923 (N_2923,N_2865,N_2898);
xor U2924 (N_2924,N_2894,N_2899);
nand U2925 (N_2925,N_2893,N_2802);
and U2926 (N_2926,N_2867,N_2828);
and U2927 (N_2927,N_2836,N_2830);
xnor U2928 (N_2928,N_2807,N_2816);
xor U2929 (N_2929,N_2844,N_2821);
and U2930 (N_2930,N_2806,N_2824);
xor U2931 (N_2931,N_2854,N_2863);
or U2932 (N_2932,N_2834,N_2841);
xor U2933 (N_2933,N_2814,N_2845);
nand U2934 (N_2934,N_2885,N_2890);
nand U2935 (N_2935,N_2862,N_2810);
nand U2936 (N_2936,N_2805,N_2861);
or U2937 (N_2937,N_2872,N_2880);
nand U2938 (N_2938,N_2871,N_2886);
nand U2939 (N_2939,N_2892,N_2843);
and U2940 (N_2940,N_2857,N_2879);
xor U2941 (N_2941,N_2856,N_2870);
nor U2942 (N_2942,N_2801,N_2873);
nand U2943 (N_2943,N_2812,N_2884);
or U2944 (N_2944,N_2831,N_2827);
xor U2945 (N_2945,N_2852,N_2832);
nor U2946 (N_2946,N_2842,N_2882);
or U2947 (N_2947,N_2868,N_2819);
nand U2948 (N_2948,N_2829,N_2860);
nand U2949 (N_2949,N_2853,N_2889);
and U2950 (N_2950,N_2890,N_2854);
xor U2951 (N_2951,N_2881,N_2821);
and U2952 (N_2952,N_2847,N_2890);
nor U2953 (N_2953,N_2810,N_2886);
xor U2954 (N_2954,N_2821,N_2861);
xnor U2955 (N_2955,N_2841,N_2851);
or U2956 (N_2956,N_2896,N_2844);
and U2957 (N_2957,N_2852,N_2808);
or U2958 (N_2958,N_2891,N_2807);
xor U2959 (N_2959,N_2827,N_2868);
and U2960 (N_2960,N_2855,N_2882);
and U2961 (N_2961,N_2846,N_2808);
xor U2962 (N_2962,N_2857,N_2846);
and U2963 (N_2963,N_2870,N_2862);
and U2964 (N_2964,N_2812,N_2878);
nor U2965 (N_2965,N_2864,N_2833);
xnor U2966 (N_2966,N_2898,N_2888);
xnor U2967 (N_2967,N_2825,N_2863);
nand U2968 (N_2968,N_2892,N_2881);
or U2969 (N_2969,N_2806,N_2802);
or U2970 (N_2970,N_2815,N_2870);
nor U2971 (N_2971,N_2812,N_2877);
nand U2972 (N_2972,N_2851,N_2873);
or U2973 (N_2973,N_2833,N_2895);
and U2974 (N_2974,N_2867,N_2889);
or U2975 (N_2975,N_2872,N_2840);
or U2976 (N_2976,N_2848,N_2852);
and U2977 (N_2977,N_2840,N_2820);
and U2978 (N_2978,N_2842,N_2898);
nor U2979 (N_2979,N_2889,N_2885);
nand U2980 (N_2980,N_2862,N_2888);
nor U2981 (N_2981,N_2812,N_2860);
and U2982 (N_2982,N_2847,N_2877);
xnor U2983 (N_2983,N_2851,N_2826);
nand U2984 (N_2984,N_2865,N_2840);
xor U2985 (N_2985,N_2809,N_2880);
and U2986 (N_2986,N_2808,N_2800);
and U2987 (N_2987,N_2859,N_2868);
nand U2988 (N_2988,N_2812,N_2842);
nor U2989 (N_2989,N_2818,N_2880);
nor U2990 (N_2990,N_2853,N_2883);
or U2991 (N_2991,N_2853,N_2817);
nor U2992 (N_2992,N_2868,N_2889);
nor U2993 (N_2993,N_2898,N_2815);
xnor U2994 (N_2994,N_2845,N_2836);
nor U2995 (N_2995,N_2810,N_2858);
and U2996 (N_2996,N_2863,N_2860);
or U2997 (N_2997,N_2897,N_2834);
nor U2998 (N_2998,N_2817,N_2821);
xor U2999 (N_2999,N_2873,N_2806);
xor U3000 (N_3000,N_2901,N_2919);
nor U3001 (N_3001,N_2939,N_2929);
xnor U3002 (N_3002,N_2995,N_2930);
nor U3003 (N_3003,N_2955,N_2963);
and U3004 (N_3004,N_2926,N_2970);
and U3005 (N_3005,N_2946,N_2973);
and U3006 (N_3006,N_2942,N_2947);
nand U3007 (N_3007,N_2981,N_2903);
and U3008 (N_3008,N_2917,N_2991);
and U3009 (N_3009,N_2993,N_2948);
or U3010 (N_3010,N_2971,N_2977);
or U3011 (N_3011,N_2956,N_2998);
and U3012 (N_3012,N_2923,N_2905);
nand U3013 (N_3013,N_2937,N_2997);
nor U3014 (N_3014,N_2925,N_2960);
xnor U3015 (N_3015,N_2913,N_2931);
nand U3016 (N_3016,N_2974,N_2982);
nand U3017 (N_3017,N_2967,N_2984);
nand U3018 (N_3018,N_2988,N_2987);
nor U3019 (N_3019,N_2924,N_2934);
nand U3020 (N_3020,N_2944,N_2914);
nand U3021 (N_3021,N_2933,N_2932);
or U3022 (N_3022,N_2910,N_2943);
or U3023 (N_3023,N_2927,N_2940);
nor U3024 (N_3024,N_2968,N_2950);
and U3025 (N_3025,N_2915,N_2904);
nand U3026 (N_3026,N_2941,N_2918);
nor U3027 (N_3027,N_2902,N_2920);
nand U3028 (N_3028,N_2965,N_2962);
xnor U3029 (N_3029,N_2909,N_2908);
and U3030 (N_3030,N_2922,N_2900);
or U3031 (N_3031,N_2979,N_2959);
nand U3032 (N_3032,N_2999,N_2976);
or U3033 (N_3033,N_2994,N_2907);
xnor U3034 (N_3034,N_2906,N_2961);
xor U3035 (N_3035,N_2972,N_2938);
and U3036 (N_3036,N_2986,N_2952);
and U3037 (N_3037,N_2921,N_2928);
and U3038 (N_3038,N_2916,N_2990);
nand U3039 (N_3039,N_2983,N_2966);
or U3040 (N_3040,N_2953,N_2957);
or U3041 (N_3041,N_2989,N_2945);
xnor U3042 (N_3042,N_2975,N_2935);
xnor U3043 (N_3043,N_2964,N_2954);
xnor U3044 (N_3044,N_2912,N_2969);
nand U3045 (N_3045,N_2911,N_2949);
nor U3046 (N_3046,N_2992,N_2958);
xor U3047 (N_3047,N_2980,N_2936);
xnor U3048 (N_3048,N_2978,N_2985);
and U3049 (N_3049,N_2951,N_2996);
xnor U3050 (N_3050,N_2900,N_2966);
nor U3051 (N_3051,N_2940,N_2937);
xnor U3052 (N_3052,N_2956,N_2975);
or U3053 (N_3053,N_2959,N_2998);
nand U3054 (N_3054,N_2927,N_2968);
nand U3055 (N_3055,N_2957,N_2905);
and U3056 (N_3056,N_2928,N_2958);
xnor U3057 (N_3057,N_2988,N_2979);
nor U3058 (N_3058,N_2931,N_2956);
nand U3059 (N_3059,N_2944,N_2975);
nand U3060 (N_3060,N_2901,N_2942);
and U3061 (N_3061,N_2926,N_2906);
nor U3062 (N_3062,N_2952,N_2946);
xor U3063 (N_3063,N_2924,N_2997);
or U3064 (N_3064,N_2951,N_2972);
and U3065 (N_3065,N_2912,N_2920);
or U3066 (N_3066,N_2911,N_2915);
nor U3067 (N_3067,N_2923,N_2982);
nor U3068 (N_3068,N_2976,N_2947);
and U3069 (N_3069,N_2954,N_2922);
nor U3070 (N_3070,N_2933,N_2931);
and U3071 (N_3071,N_2988,N_2938);
nand U3072 (N_3072,N_2986,N_2967);
and U3073 (N_3073,N_2943,N_2960);
xnor U3074 (N_3074,N_2965,N_2977);
nor U3075 (N_3075,N_2955,N_2950);
xor U3076 (N_3076,N_2972,N_2973);
nor U3077 (N_3077,N_2988,N_2923);
nor U3078 (N_3078,N_2912,N_2942);
or U3079 (N_3079,N_2954,N_2965);
nor U3080 (N_3080,N_2969,N_2926);
nand U3081 (N_3081,N_2989,N_2927);
xor U3082 (N_3082,N_2923,N_2952);
nand U3083 (N_3083,N_2948,N_2924);
or U3084 (N_3084,N_2914,N_2998);
nor U3085 (N_3085,N_2990,N_2913);
xnor U3086 (N_3086,N_2923,N_2957);
and U3087 (N_3087,N_2946,N_2958);
nor U3088 (N_3088,N_2929,N_2923);
xor U3089 (N_3089,N_2923,N_2997);
xnor U3090 (N_3090,N_2914,N_2929);
nand U3091 (N_3091,N_2956,N_2994);
and U3092 (N_3092,N_2968,N_2993);
xnor U3093 (N_3093,N_2943,N_2952);
xor U3094 (N_3094,N_2929,N_2987);
nor U3095 (N_3095,N_2964,N_2912);
nand U3096 (N_3096,N_2910,N_2930);
nand U3097 (N_3097,N_2936,N_2987);
nand U3098 (N_3098,N_2939,N_2993);
nand U3099 (N_3099,N_2948,N_2992);
nor U3100 (N_3100,N_3007,N_3045);
or U3101 (N_3101,N_3065,N_3055);
or U3102 (N_3102,N_3024,N_3079);
xnor U3103 (N_3103,N_3026,N_3083);
and U3104 (N_3104,N_3095,N_3028);
nand U3105 (N_3105,N_3014,N_3009);
or U3106 (N_3106,N_3098,N_3025);
xnor U3107 (N_3107,N_3004,N_3043);
and U3108 (N_3108,N_3048,N_3088);
or U3109 (N_3109,N_3061,N_3094);
xnor U3110 (N_3110,N_3080,N_3020);
nand U3111 (N_3111,N_3089,N_3013);
nor U3112 (N_3112,N_3068,N_3008);
nand U3113 (N_3113,N_3097,N_3066);
or U3114 (N_3114,N_3047,N_3050);
nor U3115 (N_3115,N_3021,N_3067);
or U3116 (N_3116,N_3042,N_3000);
or U3117 (N_3117,N_3032,N_3086);
xnor U3118 (N_3118,N_3073,N_3006);
xor U3119 (N_3119,N_3075,N_3082);
and U3120 (N_3120,N_3041,N_3038);
and U3121 (N_3121,N_3034,N_3063);
xnor U3122 (N_3122,N_3027,N_3062);
xor U3123 (N_3123,N_3031,N_3054);
nand U3124 (N_3124,N_3081,N_3010);
nor U3125 (N_3125,N_3052,N_3060);
nor U3126 (N_3126,N_3092,N_3046);
nor U3127 (N_3127,N_3019,N_3022);
and U3128 (N_3128,N_3096,N_3023);
nor U3129 (N_3129,N_3069,N_3093);
nand U3130 (N_3130,N_3018,N_3053);
or U3131 (N_3131,N_3030,N_3017);
nor U3132 (N_3132,N_3035,N_3074);
xor U3133 (N_3133,N_3002,N_3051);
xor U3134 (N_3134,N_3037,N_3084);
xor U3135 (N_3135,N_3049,N_3016);
nor U3136 (N_3136,N_3057,N_3040);
xor U3137 (N_3137,N_3011,N_3001);
or U3138 (N_3138,N_3003,N_3015);
and U3139 (N_3139,N_3029,N_3076);
or U3140 (N_3140,N_3099,N_3087);
or U3141 (N_3141,N_3036,N_3012);
and U3142 (N_3142,N_3005,N_3091);
nand U3143 (N_3143,N_3064,N_3085);
or U3144 (N_3144,N_3072,N_3056);
or U3145 (N_3145,N_3071,N_3039);
xor U3146 (N_3146,N_3058,N_3044);
xor U3147 (N_3147,N_3059,N_3078);
nor U3148 (N_3148,N_3070,N_3077);
nor U3149 (N_3149,N_3033,N_3090);
and U3150 (N_3150,N_3077,N_3089);
and U3151 (N_3151,N_3093,N_3049);
and U3152 (N_3152,N_3052,N_3054);
xor U3153 (N_3153,N_3029,N_3003);
nand U3154 (N_3154,N_3005,N_3027);
and U3155 (N_3155,N_3077,N_3041);
nand U3156 (N_3156,N_3074,N_3005);
nand U3157 (N_3157,N_3085,N_3089);
and U3158 (N_3158,N_3027,N_3028);
or U3159 (N_3159,N_3086,N_3038);
or U3160 (N_3160,N_3061,N_3014);
and U3161 (N_3161,N_3067,N_3006);
nor U3162 (N_3162,N_3052,N_3010);
or U3163 (N_3163,N_3058,N_3097);
nor U3164 (N_3164,N_3043,N_3063);
nand U3165 (N_3165,N_3062,N_3040);
xnor U3166 (N_3166,N_3087,N_3011);
xnor U3167 (N_3167,N_3043,N_3022);
nand U3168 (N_3168,N_3088,N_3002);
or U3169 (N_3169,N_3046,N_3080);
nand U3170 (N_3170,N_3038,N_3081);
or U3171 (N_3171,N_3017,N_3003);
xor U3172 (N_3172,N_3005,N_3043);
and U3173 (N_3173,N_3020,N_3031);
nand U3174 (N_3174,N_3090,N_3084);
or U3175 (N_3175,N_3051,N_3048);
nand U3176 (N_3176,N_3061,N_3030);
or U3177 (N_3177,N_3037,N_3054);
and U3178 (N_3178,N_3088,N_3049);
or U3179 (N_3179,N_3037,N_3034);
nor U3180 (N_3180,N_3084,N_3044);
and U3181 (N_3181,N_3047,N_3081);
nand U3182 (N_3182,N_3041,N_3018);
and U3183 (N_3183,N_3067,N_3059);
and U3184 (N_3184,N_3024,N_3031);
xnor U3185 (N_3185,N_3042,N_3002);
and U3186 (N_3186,N_3020,N_3008);
and U3187 (N_3187,N_3089,N_3093);
xor U3188 (N_3188,N_3085,N_3001);
nor U3189 (N_3189,N_3069,N_3017);
xnor U3190 (N_3190,N_3061,N_3056);
xnor U3191 (N_3191,N_3020,N_3062);
nand U3192 (N_3192,N_3075,N_3050);
xor U3193 (N_3193,N_3061,N_3059);
and U3194 (N_3194,N_3002,N_3069);
nand U3195 (N_3195,N_3079,N_3000);
nand U3196 (N_3196,N_3065,N_3083);
nand U3197 (N_3197,N_3083,N_3050);
nor U3198 (N_3198,N_3062,N_3076);
or U3199 (N_3199,N_3065,N_3069);
xor U3200 (N_3200,N_3169,N_3113);
xor U3201 (N_3201,N_3196,N_3171);
xor U3202 (N_3202,N_3127,N_3143);
and U3203 (N_3203,N_3111,N_3187);
nand U3204 (N_3204,N_3106,N_3178);
and U3205 (N_3205,N_3133,N_3193);
xor U3206 (N_3206,N_3190,N_3149);
nand U3207 (N_3207,N_3160,N_3131);
xnor U3208 (N_3208,N_3129,N_3174);
xnor U3209 (N_3209,N_3155,N_3162);
xor U3210 (N_3210,N_3163,N_3104);
nor U3211 (N_3211,N_3109,N_3168);
nand U3212 (N_3212,N_3191,N_3144);
nor U3213 (N_3213,N_3119,N_3115);
nand U3214 (N_3214,N_3146,N_3153);
and U3215 (N_3215,N_3125,N_3124);
or U3216 (N_3216,N_3122,N_3185);
xor U3217 (N_3217,N_3197,N_3136);
xnor U3218 (N_3218,N_3114,N_3139);
nor U3219 (N_3219,N_3105,N_3177);
or U3220 (N_3220,N_3100,N_3135);
or U3221 (N_3221,N_3145,N_3181);
nor U3222 (N_3222,N_3118,N_3134);
nand U3223 (N_3223,N_3140,N_3154);
nand U3224 (N_3224,N_3102,N_3188);
or U3225 (N_3225,N_3107,N_3138);
or U3226 (N_3226,N_3172,N_3198);
or U3227 (N_3227,N_3165,N_3148);
nand U3228 (N_3228,N_3126,N_3112);
nor U3229 (N_3229,N_3117,N_3183);
nor U3230 (N_3230,N_3184,N_3195);
and U3231 (N_3231,N_3186,N_3147);
or U3232 (N_3232,N_3164,N_3128);
nor U3233 (N_3233,N_3176,N_3142);
nor U3234 (N_3234,N_3179,N_3175);
xor U3235 (N_3235,N_3161,N_3103);
xnor U3236 (N_3236,N_3123,N_3182);
xor U3237 (N_3237,N_3157,N_3158);
nand U3238 (N_3238,N_3199,N_3189);
nand U3239 (N_3239,N_3116,N_3150);
nor U3240 (N_3240,N_3159,N_3132);
or U3241 (N_3241,N_3120,N_3167);
nor U3242 (N_3242,N_3192,N_3180);
and U3243 (N_3243,N_3166,N_3130);
nand U3244 (N_3244,N_3110,N_3156);
nor U3245 (N_3245,N_3108,N_3194);
xor U3246 (N_3246,N_3151,N_3137);
nand U3247 (N_3247,N_3101,N_3170);
nand U3248 (N_3248,N_3152,N_3121);
nand U3249 (N_3249,N_3141,N_3173);
xnor U3250 (N_3250,N_3112,N_3175);
or U3251 (N_3251,N_3156,N_3176);
or U3252 (N_3252,N_3191,N_3122);
nor U3253 (N_3253,N_3186,N_3109);
and U3254 (N_3254,N_3199,N_3192);
nand U3255 (N_3255,N_3173,N_3140);
nand U3256 (N_3256,N_3170,N_3185);
nand U3257 (N_3257,N_3196,N_3136);
nor U3258 (N_3258,N_3190,N_3111);
and U3259 (N_3259,N_3179,N_3101);
xor U3260 (N_3260,N_3135,N_3143);
nand U3261 (N_3261,N_3147,N_3158);
xnor U3262 (N_3262,N_3133,N_3149);
xor U3263 (N_3263,N_3198,N_3150);
or U3264 (N_3264,N_3146,N_3108);
nand U3265 (N_3265,N_3191,N_3161);
xnor U3266 (N_3266,N_3131,N_3158);
xnor U3267 (N_3267,N_3126,N_3174);
nor U3268 (N_3268,N_3184,N_3172);
or U3269 (N_3269,N_3169,N_3138);
and U3270 (N_3270,N_3186,N_3176);
nor U3271 (N_3271,N_3147,N_3166);
nand U3272 (N_3272,N_3162,N_3145);
or U3273 (N_3273,N_3164,N_3156);
xnor U3274 (N_3274,N_3112,N_3142);
xnor U3275 (N_3275,N_3120,N_3143);
and U3276 (N_3276,N_3191,N_3180);
xor U3277 (N_3277,N_3155,N_3121);
and U3278 (N_3278,N_3193,N_3111);
or U3279 (N_3279,N_3138,N_3180);
nand U3280 (N_3280,N_3131,N_3147);
and U3281 (N_3281,N_3197,N_3190);
or U3282 (N_3282,N_3128,N_3151);
or U3283 (N_3283,N_3166,N_3146);
xor U3284 (N_3284,N_3197,N_3124);
nor U3285 (N_3285,N_3112,N_3128);
or U3286 (N_3286,N_3198,N_3142);
nor U3287 (N_3287,N_3184,N_3181);
xor U3288 (N_3288,N_3104,N_3149);
and U3289 (N_3289,N_3121,N_3195);
xnor U3290 (N_3290,N_3152,N_3154);
or U3291 (N_3291,N_3177,N_3164);
nor U3292 (N_3292,N_3130,N_3198);
nor U3293 (N_3293,N_3134,N_3132);
nor U3294 (N_3294,N_3160,N_3121);
and U3295 (N_3295,N_3186,N_3113);
xor U3296 (N_3296,N_3176,N_3101);
nor U3297 (N_3297,N_3126,N_3199);
nor U3298 (N_3298,N_3156,N_3187);
and U3299 (N_3299,N_3118,N_3158);
or U3300 (N_3300,N_3200,N_3244);
or U3301 (N_3301,N_3289,N_3252);
nand U3302 (N_3302,N_3235,N_3259);
xnor U3303 (N_3303,N_3233,N_3232);
and U3304 (N_3304,N_3215,N_3249);
and U3305 (N_3305,N_3216,N_3238);
nor U3306 (N_3306,N_3204,N_3245);
nor U3307 (N_3307,N_3278,N_3254);
xor U3308 (N_3308,N_3286,N_3251);
nand U3309 (N_3309,N_3229,N_3208);
xor U3310 (N_3310,N_3230,N_3258);
or U3311 (N_3311,N_3222,N_3219);
xnor U3312 (N_3312,N_3294,N_3243);
and U3313 (N_3313,N_3205,N_3247);
or U3314 (N_3314,N_3296,N_3265);
or U3315 (N_3315,N_3210,N_3227);
or U3316 (N_3316,N_3272,N_3277);
and U3317 (N_3317,N_3285,N_3260);
or U3318 (N_3318,N_3280,N_3250);
or U3319 (N_3319,N_3269,N_3220);
and U3320 (N_3320,N_3207,N_3299);
and U3321 (N_3321,N_3275,N_3214);
or U3322 (N_3322,N_3242,N_3279);
nor U3323 (N_3323,N_3268,N_3255);
nand U3324 (N_3324,N_3224,N_3203);
or U3325 (N_3325,N_3281,N_3282);
xor U3326 (N_3326,N_3246,N_3228);
xnor U3327 (N_3327,N_3241,N_3288);
nand U3328 (N_3328,N_3226,N_3264);
xnor U3329 (N_3329,N_3273,N_3284);
nor U3330 (N_3330,N_3262,N_3276);
xor U3331 (N_3331,N_3274,N_3221);
nor U3332 (N_3332,N_3266,N_3231);
xor U3333 (N_3333,N_3283,N_3263);
and U3334 (N_3334,N_3209,N_3223);
xnor U3335 (N_3335,N_3297,N_3290);
xnor U3336 (N_3336,N_3270,N_3261);
and U3337 (N_3337,N_3256,N_3211);
or U3338 (N_3338,N_3271,N_3218);
or U3339 (N_3339,N_3237,N_3292);
nor U3340 (N_3340,N_3248,N_3225);
nand U3341 (N_3341,N_3293,N_3239);
or U3342 (N_3342,N_3298,N_3257);
nand U3343 (N_3343,N_3201,N_3236);
xor U3344 (N_3344,N_3295,N_3212);
xnor U3345 (N_3345,N_3253,N_3213);
and U3346 (N_3346,N_3287,N_3234);
and U3347 (N_3347,N_3291,N_3240);
or U3348 (N_3348,N_3267,N_3206);
or U3349 (N_3349,N_3217,N_3202);
nand U3350 (N_3350,N_3291,N_3251);
nor U3351 (N_3351,N_3278,N_3290);
nor U3352 (N_3352,N_3298,N_3288);
or U3353 (N_3353,N_3280,N_3259);
nand U3354 (N_3354,N_3268,N_3264);
nand U3355 (N_3355,N_3210,N_3270);
xnor U3356 (N_3356,N_3256,N_3289);
or U3357 (N_3357,N_3296,N_3278);
nor U3358 (N_3358,N_3264,N_3288);
and U3359 (N_3359,N_3214,N_3245);
and U3360 (N_3360,N_3218,N_3239);
nor U3361 (N_3361,N_3265,N_3272);
nor U3362 (N_3362,N_3280,N_3272);
and U3363 (N_3363,N_3284,N_3258);
and U3364 (N_3364,N_3280,N_3278);
or U3365 (N_3365,N_3268,N_3269);
nand U3366 (N_3366,N_3203,N_3279);
or U3367 (N_3367,N_3280,N_3261);
nand U3368 (N_3368,N_3222,N_3252);
nand U3369 (N_3369,N_3299,N_3236);
nor U3370 (N_3370,N_3292,N_3299);
and U3371 (N_3371,N_3277,N_3241);
nor U3372 (N_3372,N_3287,N_3258);
nand U3373 (N_3373,N_3273,N_3272);
or U3374 (N_3374,N_3297,N_3206);
and U3375 (N_3375,N_3217,N_3273);
xnor U3376 (N_3376,N_3252,N_3255);
or U3377 (N_3377,N_3243,N_3200);
nand U3378 (N_3378,N_3224,N_3288);
xor U3379 (N_3379,N_3267,N_3241);
nand U3380 (N_3380,N_3211,N_3209);
xnor U3381 (N_3381,N_3226,N_3247);
xnor U3382 (N_3382,N_3216,N_3211);
or U3383 (N_3383,N_3296,N_3232);
or U3384 (N_3384,N_3261,N_3272);
and U3385 (N_3385,N_3262,N_3226);
or U3386 (N_3386,N_3223,N_3204);
and U3387 (N_3387,N_3259,N_3220);
nor U3388 (N_3388,N_3287,N_3273);
xnor U3389 (N_3389,N_3251,N_3290);
nor U3390 (N_3390,N_3261,N_3235);
nand U3391 (N_3391,N_3243,N_3227);
and U3392 (N_3392,N_3216,N_3226);
xor U3393 (N_3393,N_3220,N_3282);
nand U3394 (N_3394,N_3279,N_3212);
nand U3395 (N_3395,N_3216,N_3284);
nor U3396 (N_3396,N_3204,N_3289);
nor U3397 (N_3397,N_3244,N_3269);
nor U3398 (N_3398,N_3251,N_3234);
xnor U3399 (N_3399,N_3238,N_3236);
xnor U3400 (N_3400,N_3383,N_3382);
or U3401 (N_3401,N_3315,N_3309);
nand U3402 (N_3402,N_3386,N_3325);
xor U3403 (N_3403,N_3317,N_3304);
nor U3404 (N_3404,N_3320,N_3324);
nor U3405 (N_3405,N_3326,N_3323);
xnor U3406 (N_3406,N_3350,N_3376);
nand U3407 (N_3407,N_3316,N_3305);
nand U3408 (N_3408,N_3336,N_3360);
xor U3409 (N_3409,N_3308,N_3385);
nor U3410 (N_3410,N_3348,N_3380);
and U3411 (N_3411,N_3372,N_3369);
and U3412 (N_3412,N_3341,N_3359);
nor U3413 (N_3413,N_3391,N_3330);
xor U3414 (N_3414,N_3354,N_3353);
nand U3415 (N_3415,N_3390,N_3349);
or U3416 (N_3416,N_3374,N_3388);
nor U3417 (N_3417,N_3337,N_3399);
xnor U3418 (N_3418,N_3364,N_3394);
and U3419 (N_3419,N_3361,N_3310);
xnor U3420 (N_3420,N_3392,N_3312);
nand U3421 (N_3421,N_3377,N_3378);
and U3422 (N_3422,N_3357,N_3375);
nor U3423 (N_3423,N_3334,N_3342);
or U3424 (N_3424,N_3347,N_3366);
nor U3425 (N_3425,N_3352,N_3301);
xor U3426 (N_3426,N_3351,N_3344);
nand U3427 (N_3427,N_3319,N_3370);
or U3428 (N_3428,N_3397,N_3381);
nor U3429 (N_3429,N_3321,N_3368);
and U3430 (N_3430,N_3340,N_3356);
and U3431 (N_3431,N_3327,N_3393);
nor U3432 (N_3432,N_3306,N_3303);
xor U3433 (N_3433,N_3345,N_3329);
nand U3434 (N_3434,N_3363,N_3300);
nor U3435 (N_3435,N_3387,N_3313);
nor U3436 (N_3436,N_3395,N_3389);
and U3437 (N_3437,N_3328,N_3355);
nor U3438 (N_3438,N_3311,N_3333);
nor U3439 (N_3439,N_3358,N_3371);
xor U3440 (N_3440,N_3373,N_3332);
xor U3441 (N_3441,N_3302,N_3365);
and U3442 (N_3442,N_3318,N_3339);
and U3443 (N_3443,N_3322,N_3367);
and U3444 (N_3444,N_3396,N_3338);
and U3445 (N_3445,N_3331,N_3362);
nor U3446 (N_3446,N_3346,N_3384);
and U3447 (N_3447,N_3307,N_3379);
xor U3448 (N_3448,N_3398,N_3314);
and U3449 (N_3449,N_3335,N_3343);
xnor U3450 (N_3450,N_3381,N_3318);
nor U3451 (N_3451,N_3375,N_3306);
nor U3452 (N_3452,N_3301,N_3386);
nor U3453 (N_3453,N_3348,N_3317);
and U3454 (N_3454,N_3321,N_3391);
nand U3455 (N_3455,N_3334,N_3309);
nand U3456 (N_3456,N_3390,N_3385);
and U3457 (N_3457,N_3342,N_3382);
and U3458 (N_3458,N_3317,N_3360);
nand U3459 (N_3459,N_3325,N_3321);
nand U3460 (N_3460,N_3320,N_3358);
nand U3461 (N_3461,N_3336,N_3307);
and U3462 (N_3462,N_3331,N_3357);
and U3463 (N_3463,N_3308,N_3378);
nand U3464 (N_3464,N_3388,N_3331);
nor U3465 (N_3465,N_3315,N_3366);
and U3466 (N_3466,N_3351,N_3383);
xnor U3467 (N_3467,N_3304,N_3383);
and U3468 (N_3468,N_3301,N_3334);
xnor U3469 (N_3469,N_3350,N_3348);
nand U3470 (N_3470,N_3350,N_3398);
and U3471 (N_3471,N_3341,N_3390);
or U3472 (N_3472,N_3398,N_3372);
or U3473 (N_3473,N_3353,N_3374);
nand U3474 (N_3474,N_3360,N_3310);
nor U3475 (N_3475,N_3395,N_3326);
nand U3476 (N_3476,N_3371,N_3354);
xnor U3477 (N_3477,N_3331,N_3368);
xnor U3478 (N_3478,N_3346,N_3365);
or U3479 (N_3479,N_3323,N_3383);
xnor U3480 (N_3480,N_3321,N_3308);
xor U3481 (N_3481,N_3393,N_3385);
and U3482 (N_3482,N_3325,N_3364);
or U3483 (N_3483,N_3352,N_3373);
xnor U3484 (N_3484,N_3358,N_3307);
or U3485 (N_3485,N_3387,N_3331);
xnor U3486 (N_3486,N_3313,N_3388);
nand U3487 (N_3487,N_3322,N_3309);
nor U3488 (N_3488,N_3363,N_3325);
xor U3489 (N_3489,N_3301,N_3349);
nand U3490 (N_3490,N_3328,N_3377);
nor U3491 (N_3491,N_3382,N_3329);
and U3492 (N_3492,N_3346,N_3318);
nand U3493 (N_3493,N_3383,N_3318);
xnor U3494 (N_3494,N_3317,N_3355);
or U3495 (N_3495,N_3343,N_3359);
and U3496 (N_3496,N_3349,N_3329);
or U3497 (N_3497,N_3392,N_3342);
nor U3498 (N_3498,N_3337,N_3361);
and U3499 (N_3499,N_3392,N_3337);
or U3500 (N_3500,N_3468,N_3451);
nor U3501 (N_3501,N_3443,N_3409);
xnor U3502 (N_3502,N_3498,N_3480);
and U3503 (N_3503,N_3420,N_3450);
or U3504 (N_3504,N_3446,N_3457);
xnor U3505 (N_3505,N_3418,N_3427);
nand U3506 (N_3506,N_3441,N_3472);
nand U3507 (N_3507,N_3401,N_3463);
nor U3508 (N_3508,N_3469,N_3402);
and U3509 (N_3509,N_3466,N_3416);
or U3510 (N_3510,N_3477,N_3404);
and U3511 (N_3511,N_3434,N_3429);
or U3512 (N_3512,N_3448,N_3482);
nand U3513 (N_3513,N_3485,N_3479);
or U3514 (N_3514,N_3474,N_3496);
xnor U3515 (N_3515,N_3491,N_3413);
nand U3516 (N_3516,N_3481,N_3436);
and U3517 (N_3517,N_3497,N_3464);
and U3518 (N_3518,N_3453,N_3470);
or U3519 (N_3519,N_3447,N_3428);
nor U3520 (N_3520,N_3421,N_3486);
nor U3521 (N_3521,N_3493,N_3440);
xnor U3522 (N_3522,N_3417,N_3495);
or U3523 (N_3523,N_3419,N_3490);
xnor U3524 (N_3524,N_3433,N_3484);
and U3525 (N_3525,N_3431,N_3488);
and U3526 (N_3526,N_3437,N_3449);
or U3527 (N_3527,N_3492,N_3435);
xor U3528 (N_3528,N_3458,N_3411);
xor U3529 (N_3529,N_3455,N_3499);
xnor U3530 (N_3530,N_3444,N_3406);
or U3531 (N_3531,N_3471,N_3425);
nand U3532 (N_3532,N_3422,N_3461);
nor U3533 (N_3533,N_3407,N_3454);
nand U3534 (N_3534,N_3494,N_3473);
nand U3535 (N_3535,N_3438,N_3487);
nand U3536 (N_3536,N_3412,N_3414);
or U3537 (N_3537,N_3459,N_3445);
nand U3538 (N_3538,N_3462,N_3415);
xor U3539 (N_3539,N_3483,N_3442);
and U3540 (N_3540,N_3465,N_3423);
xor U3541 (N_3541,N_3400,N_3426);
nand U3542 (N_3542,N_3478,N_3460);
or U3543 (N_3543,N_3403,N_3405);
xor U3544 (N_3544,N_3452,N_3467);
nand U3545 (N_3545,N_3476,N_3430);
nand U3546 (N_3546,N_3439,N_3489);
or U3547 (N_3547,N_3475,N_3424);
nand U3548 (N_3548,N_3432,N_3410);
nand U3549 (N_3549,N_3456,N_3408);
or U3550 (N_3550,N_3489,N_3467);
nand U3551 (N_3551,N_3425,N_3416);
or U3552 (N_3552,N_3456,N_3454);
nor U3553 (N_3553,N_3460,N_3492);
nand U3554 (N_3554,N_3480,N_3457);
nand U3555 (N_3555,N_3447,N_3462);
or U3556 (N_3556,N_3468,N_3439);
or U3557 (N_3557,N_3421,N_3434);
and U3558 (N_3558,N_3436,N_3406);
or U3559 (N_3559,N_3402,N_3423);
xor U3560 (N_3560,N_3454,N_3443);
xnor U3561 (N_3561,N_3481,N_3424);
or U3562 (N_3562,N_3477,N_3403);
xor U3563 (N_3563,N_3406,N_3422);
nor U3564 (N_3564,N_3483,N_3496);
xnor U3565 (N_3565,N_3434,N_3462);
nand U3566 (N_3566,N_3489,N_3490);
or U3567 (N_3567,N_3496,N_3401);
or U3568 (N_3568,N_3473,N_3499);
xnor U3569 (N_3569,N_3492,N_3407);
xnor U3570 (N_3570,N_3453,N_3441);
or U3571 (N_3571,N_3475,N_3429);
and U3572 (N_3572,N_3446,N_3419);
and U3573 (N_3573,N_3481,N_3459);
nand U3574 (N_3574,N_3426,N_3440);
nor U3575 (N_3575,N_3460,N_3431);
nor U3576 (N_3576,N_3454,N_3462);
or U3577 (N_3577,N_3441,N_3490);
xnor U3578 (N_3578,N_3444,N_3494);
and U3579 (N_3579,N_3486,N_3495);
nor U3580 (N_3580,N_3474,N_3449);
nand U3581 (N_3581,N_3445,N_3405);
or U3582 (N_3582,N_3424,N_3488);
and U3583 (N_3583,N_3460,N_3428);
nand U3584 (N_3584,N_3439,N_3435);
xor U3585 (N_3585,N_3498,N_3437);
nand U3586 (N_3586,N_3489,N_3475);
or U3587 (N_3587,N_3455,N_3490);
and U3588 (N_3588,N_3499,N_3446);
and U3589 (N_3589,N_3448,N_3427);
or U3590 (N_3590,N_3425,N_3412);
or U3591 (N_3591,N_3496,N_3402);
or U3592 (N_3592,N_3456,N_3478);
nand U3593 (N_3593,N_3471,N_3458);
and U3594 (N_3594,N_3404,N_3474);
and U3595 (N_3595,N_3444,N_3408);
and U3596 (N_3596,N_3405,N_3436);
and U3597 (N_3597,N_3428,N_3427);
nor U3598 (N_3598,N_3490,N_3442);
nand U3599 (N_3599,N_3451,N_3472);
nand U3600 (N_3600,N_3535,N_3571);
xnor U3601 (N_3601,N_3583,N_3527);
nor U3602 (N_3602,N_3526,N_3543);
or U3603 (N_3603,N_3591,N_3585);
and U3604 (N_3604,N_3532,N_3509);
and U3605 (N_3605,N_3514,N_3573);
or U3606 (N_3606,N_3540,N_3516);
nor U3607 (N_3607,N_3563,N_3556);
or U3608 (N_3608,N_3512,N_3522);
or U3609 (N_3609,N_3531,N_3567);
xor U3610 (N_3610,N_3520,N_3548);
nor U3611 (N_3611,N_3578,N_3570);
xnor U3612 (N_3612,N_3506,N_3557);
and U3613 (N_3613,N_3545,N_3559);
or U3614 (N_3614,N_3576,N_3550);
and U3615 (N_3615,N_3595,N_3566);
and U3616 (N_3616,N_3503,N_3581);
and U3617 (N_3617,N_3541,N_3500);
or U3618 (N_3618,N_3546,N_3517);
xnor U3619 (N_3619,N_3552,N_3577);
xor U3620 (N_3620,N_3580,N_3560);
or U3621 (N_3621,N_3539,N_3530);
nand U3622 (N_3622,N_3558,N_3524);
xor U3623 (N_3623,N_3528,N_3533);
or U3624 (N_3624,N_3588,N_3587);
or U3625 (N_3625,N_3505,N_3547);
or U3626 (N_3626,N_3592,N_3574);
and U3627 (N_3627,N_3529,N_3593);
or U3628 (N_3628,N_3513,N_3569);
or U3629 (N_3629,N_3572,N_3502);
xnor U3630 (N_3630,N_3553,N_3501);
and U3631 (N_3631,N_3594,N_3561);
nor U3632 (N_3632,N_3554,N_3544);
or U3633 (N_3633,N_3521,N_3575);
nand U3634 (N_3634,N_3579,N_3582);
nor U3635 (N_3635,N_3538,N_3542);
nor U3636 (N_3636,N_3537,N_3511);
nor U3637 (N_3637,N_3523,N_3525);
and U3638 (N_3638,N_3507,N_3504);
or U3639 (N_3639,N_3597,N_3599);
nand U3640 (N_3640,N_3565,N_3596);
or U3641 (N_3641,N_3555,N_3534);
or U3642 (N_3642,N_3568,N_3586);
or U3643 (N_3643,N_3518,N_3584);
xor U3644 (N_3644,N_3590,N_3598);
nor U3645 (N_3645,N_3508,N_3562);
xnor U3646 (N_3646,N_3515,N_3589);
or U3647 (N_3647,N_3551,N_3549);
and U3648 (N_3648,N_3564,N_3519);
or U3649 (N_3649,N_3536,N_3510);
or U3650 (N_3650,N_3573,N_3587);
nand U3651 (N_3651,N_3514,N_3531);
and U3652 (N_3652,N_3597,N_3546);
xnor U3653 (N_3653,N_3523,N_3595);
nor U3654 (N_3654,N_3521,N_3588);
nor U3655 (N_3655,N_3530,N_3599);
and U3656 (N_3656,N_3548,N_3541);
nand U3657 (N_3657,N_3515,N_3502);
nand U3658 (N_3658,N_3547,N_3516);
nand U3659 (N_3659,N_3598,N_3504);
or U3660 (N_3660,N_3521,N_3533);
xnor U3661 (N_3661,N_3558,N_3563);
xnor U3662 (N_3662,N_3552,N_3571);
nor U3663 (N_3663,N_3524,N_3544);
nand U3664 (N_3664,N_3503,N_3556);
xor U3665 (N_3665,N_3515,N_3565);
and U3666 (N_3666,N_3506,N_3504);
nand U3667 (N_3667,N_3565,N_3513);
xnor U3668 (N_3668,N_3540,N_3530);
xor U3669 (N_3669,N_3586,N_3592);
xnor U3670 (N_3670,N_3541,N_3536);
and U3671 (N_3671,N_3566,N_3532);
xnor U3672 (N_3672,N_3508,N_3567);
or U3673 (N_3673,N_3552,N_3541);
nor U3674 (N_3674,N_3528,N_3527);
nor U3675 (N_3675,N_3568,N_3562);
xor U3676 (N_3676,N_3530,N_3558);
nand U3677 (N_3677,N_3503,N_3570);
nor U3678 (N_3678,N_3535,N_3512);
or U3679 (N_3679,N_3564,N_3520);
nand U3680 (N_3680,N_3576,N_3565);
or U3681 (N_3681,N_3548,N_3581);
nor U3682 (N_3682,N_3507,N_3538);
nor U3683 (N_3683,N_3537,N_3525);
xnor U3684 (N_3684,N_3501,N_3509);
nor U3685 (N_3685,N_3589,N_3557);
nand U3686 (N_3686,N_3506,N_3528);
or U3687 (N_3687,N_3531,N_3527);
nand U3688 (N_3688,N_3506,N_3516);
nor U3689 (N_3689,N_3543,N_3580);
xnor U3690 (N_3690,N_3575,N_3585);
nor U3691 (N_3691,N_3518,N_3520);
nor U3692 (N_3692,N_3588,N_3543);
xnor U3693 (N_3693,N_3563,N_3515);
or U3694 (N_3694,N_3547,N_3512);
and U3695 (N_3695,N_3545,N_3537);
or U3696 (N_3696,N_3573,N_3500);
nand U3697 (N_3697,N_3516,N_3599);
nor U3698 (N_3698,N_3526,N_3507);
or U3699 (N_3699,N_3552,N_3546);
nor U3700 (N_3700,N_3636,N_3649);
xnor U3701 (N_3701,N_3611,N_3600);
xor U3702 (N_3702,N_3665,N_3628);
xnor U3703 (N_3703,N_3654,N_3624);
nand U3704 (N_3704,N_3662,N_3696);
or U3705 (N_3705,N_3677,N_3653);
and U3706 (N_3706,N_3699,N_3661);
nand U3707 (N_3707,N_3660,N_3610);
nand U3708 (N_3708,N_3646,N_3604);
and U3709 (N_3709,N_3695,N_3618);
or U3710 (N_3710,N_3656,N_3688);
nor U3711 (N_3711,N_3619,N_3697);
nor U3712 (N_3712,N_3674,N_3664);
nor U3713 (N_3713,N_3622,N_3672);
nand U3714 (N_3714,N_3640,N_3657);
nor U3715 (N_3715,N_3643,N_3633);
nand U3716 (N_3716,N_3647,N_3607);
nand U3717 (N_3717,N_3602,N_3679);
nand U3718 (N_3718,N_3666,N_3641);
and U3719 (N_3719,N_3675,N_3634);
nand U3720 (N_3720,N_3663,N_3684);
nand U3721 (N_3721,N_3627,N_3608);
nand U3722 (N_3722,N_3686,N_3615);
or U3723 (N_3723,N_3639,N_3651);
or U3724 (N_3724,N_3637,N_3630);
nor U3725 (N_3725,N_3616,N_3601);
or U3726 (N_3726,N_3678,N_3670);
or U3727 (N_3727,N_3676,N_3681);
or U3728 (N_3728,N_3614,N_3689);
or U3729 (N_3729,N_3680,N_3606);
xor U3730 (N_3730,N_3655,N_3652);
or U3731 (N_3731,N_3693,N_3621);
nor U3732 (N_3732,N_3623,N_3694);
or U3733 (N_3733,N_3667,N_3673);
or U3734 (N_3734,N_3659,N_3698);
nor U3735 (N_3735,N_3617,N_3648);
nand U3736 (N_3736,N_3658,N_3635);
xor U3737 (N_3737,N_3613,N_3645);
and U3738 (N_3738,N_3612,N_3687);
and U3739 (N_3739,N_3671,N_3644);
nor U3740 (N_3740,N_3609,N_3669);
and U3741 (N_3741,N_3691,N_3682);
and U3742 (N_3742,N_3620,N_3683);
nor U3743 (N_3743,N_3625,N_3629);
xor U3744 (N_3744,N_3692,N_3690);
or U3745 (N_3745,N_3631,N_3603);
or U3746 (N_3746,N_3638,N_3632);
xnor U3747 (N_3747,N_3642,N_3668);
xnor U3748 (N_3748,N_3685,N_3626);
xor U3749 (N_3749,N_3650,N_3605);
nor U3750 (N_3750,N_3636,N_3693);
or U3751 (N_3751,N_3698,N_3654);
nor U3752 (N_3752,N_3611,N_3669);
nor U3753 (N_3753,N_3682,N_3601);
nor U3754 (N_3754,N_3678,N_3697);
xor U3755 (N_3755,N_3679,N_3680);
and U3756 (N_3756,N_3633,N_3668);
nand U3757 (N_3757,N_3692,N_3655);
and U3758 (N_3758,N_3608,N_3670);
nor U3759 (N_3759,N_3602,N_3647);
nor U3760 (N_3760,N_3640,N_3673);
xnor U3761 (N_3761,N_3665,N_3675);
nand U3762 (N_3762,N_3629,N_3609);
or U3763 (N_3763,N_3677,N_3636);
xor U3764 (N_3764,N_3690,N_3616);
nand U3765 (N_3765,N_3638,N_3614);
and U3766 (N_3766,N_3628,N_3688);
and U3767 (N_3767,N_3638,N_3664);
nor U3768 (N_3768,N_3645,N_3642);
or U3769 (N_3769,N_3606,N_3638);
nand U3770 (N_3770,N_3686,N_3643);
and U3771 (N_3771,N_3689,N_3691);
nor U3772 (N_3772,N_3621,N_3647);
xor U3773 (N_3773,N_3698,N_3685);
or U3774 (N_3774,N_3646,N_3680);
or U3775 (N_3775,N_3624,N_3689);
nor U3776 (N_3776,N_3608,N_3616);
nand U3777 (N_3777,N_3601,N_3618);
nand U3778 (N_3778,N_3679,N_3675);
and U3779 (N_3779,N_3688,N_3607);
xor U3780 (N_3780,N_3652,N_3699);
xnor U3781 (N_3781,N_3674,N_3693);
or U3782 (N_3782,N_3616,N_3667);
nor U3783 (N_3783,N_3653,N_3603);
or U3784 (N_3784,N_3631,N_3662);
xor U3785 (N_3785,N_3647,N_3698);
or U3786 (N_3786,N_3611,N_3637);
or U3787 (N_3787,N_3676,N_3632);
nand U3788 (N_3788,N_3657,N_3637);
nor U3789 (N_3789,N_3634,N_3614);
nor U3790 (N_3790,N_3601,N_3611);
nor U3791 (N_3791,N_3695,N_3686);
or U3792 (N_3792,N_3664,N_3672);
and U3793 (N_3793,N_3613,N_3660);
nand U3794 (N_3794,N_3673,N_3693);
xor U3795 (N_3795,N_3687,N_3619);
or U3796 (N_3796,N_3645,N_3659);
xnor U3797 (N_3797,N_3644,N_3606);
or U3798 (N_3798,N_3697,N_3666);
nor U3799 (N_3799,N_3627,N_3636);
and U3800 (N_3800,N_3724,N_3717);
and U3801 (N_3801,N_3713,N_3702);
nor U3802 (N_3802,N_3765,N_3785);
nand U3803 (N_3803,N_3755,N_3783);
xor U3804 (N_3804,N_3794,N_3709);
nor U3805 (N_3805,N_3745,N_3737);
and U3806 (N_3806,N_3776,N_3784);
and U3807 (N_3807,N_3750,N_3733);
nor U3808 (N_3808,N_3731,N_3754);
nand U3809 (N_3809,N_3780,N_3704);
and U3810 (N_3810,N_3712,N_3798);
and U3811 (N_3811,N_3739,N_3795);
nor U3812 (N_3812,N_3793,N_3727);
and U3813 (N_3813,N_3720,N_3722);
or U3814 (N_3814,N_3759,N_3714);
and U3815 (N_3815,N_3772,N_3769);
xor U3816 (N_3816,N_3799,N_3746);
nor U3817 (N_3817,N_3770,N_3753);
xor U3818 (N_3818,N_3701,N_3742);
nor U3819 (N_3819,N_3760,N_3775);
nor U3820 (N_3820,N_3758,N_3741);
nor U3821 (N_3821,N_3728,N_3716);
nand U3822 (N_3822,N_3751,N_3744);
nand U3823 (N_3823,N_3787,N_3721);
nand U3824 (N_3824,N_3706,N_3763);
xor U3825 (N_3825,N_3779,N_3729);
nor U3826 (N_3826,N_3747,N_3797);
nor U3827 (N_3827,N_3764,N_3719);
xor U3828 (N_3828,N_3752,N_3718);
or U3829 (N_3829,N_3761,N_3715);
xnor U3830 (N_3830,N_3734,N_3796);
and U3831 (N_3831,N_3762,N_3756);
and U3832 (N_3832,N_3792,N_3708);
nor U3833 (N_3833,N_3723,N_3738);
nor U3834 (N_3834,N_3748,N_3711);
or U3835 (N_3835,N_3743,N_3790);
nor U3836 (N_3836,N_3782,N_3768);
or U3837 (N_3837,N_3766,N_3757);
nand U3838 (N_3838,N_3749,N_3705);
xor U3839 (N_3839,N_3740,N_3791);
nor U3840 (N_3840,N_3732,N_3710);
xor U3841 (N_3841,N_3786,N_3700);
xnor U3842 (N_3842,N_3788,N_3789);
or U3843 (N_3843,N_3735,N_3774);
nand U3844 (N_3844,N_3773,N_3703);
nor U3845 (N_3845,N_3725,N_3726);
nor U3846 (N_3846,N_3767,N_3707);
nand U3847 (N_3847,N_3778,N_3736);
xor U3848 (N_3848,N_3777,N_3730);
nor U3849 (N_3849,N_3781,N_3771);
xnor U3850 (N_3850,N_3707,N_3777);
or U3851 (N_3851,N_3758,N_3710);
xnor U3852 (N_3852,N_3700,N_3797);
and U3853 (N_3853,N_3762,N_3779);
nand U3854 (N_3854,N_3786,N_3740);
nor U3855 (N_3855,N_3714,N_3791);
nand U3856 (N_3856,N_3742,N_3730);
or U3857 (N_3857,N_3731,N_3715);
nor U3858 (N_3858,N_3792,N_3738);
and U3859 (N_3859,N_3717,N_3749);
nand U3860 (N_3860,N_3781,N_3772);
nand U3861 (N_3861,N_3729,N_3725);
nand U3862 (N_3862,N_3709,N_3707);
nor U3863 (N_3863,N_3770,N_3757);
nand U3864 (N_3864,N_3727,N_3761);
nor U3865 (N_3865,N_3767,N_3791);
nor U3866 (N_3866,N_3773,N_3735);
and U3867 (N_3867,N_3736,N_3750);
xnor U3868 (N_3868,N_3796,N_3713);
and U3869 (N_3869,N_3770,N_3738);
and U3870 (N_3870,N_3740,N_3752);
and U3871 (N_3871,N_3773,N_3788);
nor U3872 (N_3872,N_3710,N_3753);
or U3873 (N_3873,N_3733,N_3752);
xor U3874 (N_3874,N_3716,N_3797);
or U3875 (N_3875,N_3771,N_3709);
and U3876 (N_3876,N_3707,N_3737);
or U3877 (N_3877,N_3729,N_3721);
or U3878 (N_3878,N_3727,N_3720);
or U3879 (N_3879,N_3772,N_3700);
and U3880 (N_3880,N_3720,N_3796);
nand U3881 (N_3881,N_3772,N_3799);
nor U3882 (N_3882,N_3719,N_3769);
nor U3883 (N_3883,N_3722,N_3784);
and U3884 (N_3884,N_3732,N_3773);
nand U3885 (N_3885,N_3754,N_3726);
and U3886 (N_3886,N_3744,N_3749);
nor U3887 (N_3887,N_3741,N_3712);
xor U3888 (N_3888,N_3756,N_3702);
nand U3889 (N_3889,N_3764,N_3777);
xor U3890 (N_3890,N_3777,N_3774);
xnor U3891 (N_3891,N_3770,N_3723);
or U3892 (N_3892,N_3764,N_3772);
nand U3893 (N_3893,N_3700,N_3702);
nand U3894 (N_3894,N_3792,N_3759);
and U3895 (N_3895,N_3734,N_3728);
xnor U3896 (N_3896,N_3796,N_3711);
or U3897 (N_3897,N_3747,N_3728);
xnor U3898 (N_3898,N_3742,N_3778);
nand U3899 (N_3899,N_3752,N_3742);
nor U3900 (N_3900,N_3825,N_3887);
nand U3901 (N_3901,N_3832,N_3816);
xor U3902 (N_3902,N_3871,N_3860);
nand U3903 (N_3903,N_3801,N_3879);
and U3904 (N_3904,N_3820,N_3851);
xor U3905 (N_3905,N_3848,N_3859);
and U3906 (N_3906,N_3850,N_3823);
and U3907 (N_3907,N_3803,N_3873);
xnor U3908 (N_3908,N_3835,N_3828);
or U3909 (N_3909,N_3889,N_3824);
and U3910 (N_3910,N_3857,N_3853);
and U3911 (N_3911,N_3834,N_3845);
nand U3912 (N_3912,N_3822,N_3842);
or U3913 (N_3913,N_3882,N_3839);
nand U3914 (N_3914,N_3812,N_3868);
nand U3915 (N_3915,N_3833,N_3897);
nand U3916 (N_3916,N_3894,N_3826);
nor U3917 (N_3917,N_3844,N_3890);
or U3918 (N_3918,N_3831,N_3819);
nor U3919 (N_3919,N_3856,N_3864);
nor U3920 (N_3920,N_3862,N_3808);
xor U3921 (N_3921,N_3837,N_3896);
nand U3922 (N_3922,N_3867,N_3883);
nand U3923 (N_3923,N_3885,N_3892);
nor U3924 (N_3924,N_3806,N_3817);
and U3925 (N_3925,N_3854,N_3814);
or U3926 (N_3926,N_3855,N_3807);
xnor U3927 (N_3927,N_3893,N_3841);
and U3928 (N_3928,N_3876,N_3895);
nand U3929 (N_3929,N_3836,N_3840);
or U3930 (N_3930,N_3869,N_3827);
and U3931 (N_3931,N_3872,N_3846);
xnor U3932 (N_3932,N_3870,N_3858);
and U3933 (N_3933,N_3800,N_3878);
and U3934 (N_3934,N_3888,N_3852);
or U3935 (N_3935,N_3805,N_3843);
and U3936 (N_3936,N_3899,N_3861);
and U3937 (N_3937,N_3811,N_3813);
nand U3938 (N_3938,N_3877,N_3829);
nand U3939 (N_3939,N_3810,N_3898);
nor U3940 (N_3940,N_3802,N_3804);
and U3941 (N_3941,N_3891,N_3815);
xnor U3942 (N_3942,N_3863,N_3881);
or U3943 (N_3943,N_3830,N_3847);
nand U3944 (N_3944,N_3865,N_3880);
nor U3945 (N_3945,N_3809,N_3875);
nor U3946 (N_3946,N_3874,N_3866);
xor U3947 (N_3947,N_3818,N_3838);
and U3948 (N_3948,N_3849,N_3884);
or U3949 (N_3949,N_3821,N_3886);
nor U3950 (N_3950,N_3875,N_3896);
nand U3951 (N_3951,N_3868,N_3840);
xnor U3952 (N_3952,N_3894,N_3856);
xor U3953 (N_3953,N_3865,N_3836);
and U3954 (N_3954,N_3877,N_3869);
nand U3955 (N_3955,N_3893,N_3891);
and U3956 (N_3956,N_3891,N_3892);
xor U3957 (N_3957,N_3829,N_3864);
nand U3958 (N_3958,N_3896,N_3836);
or U3959 (N_3959,N_3845,N_3867);
and U3960 (N_3960,N_3872,N_3833);
nor U3961 (N_3961,N_3840,N_3844);
or U3962 (N_3962,N_3893,N_3806);
xor U3963 (N_3963,N_3816,N_3865);
nand U3964 (N_3964,N_3845,N_3833);
nand U3965 (N_3965,N_3801,N_3883);
and U3966 (N_3966,N_3856,N_3862);
nor U3967 (N_3967,N_3859,N_3818);
nor U3968 (N_3968,N_3822,N_3871);
nor U3969 (N_3969,N_3805,N_3839);
nor U3970 (N_3970,N_3818,N_3856);
or U3971 (N_3971,N_3843,N_3831);
and U3972 (N_3972,N_3809,N_3832);
nor U3973 (N_3973,N_3811,N_3854);
nand U3974 (N_3974,N_3848,N_3837);
nor U3975 (N_3975,N_3870,N_3835);
nand U3976 (N_3976,N_3802,N_3891);
and U3977 (N_3977,N_3891,N_3839);
or U3978 (N_3978,N_3832,N_3872);
nor U3979 (N_3979,N_3844,N_3805);
or U3980 (N_3980,N_3894,N_3853);
or U3981 (N_3981,N_3833,N_3825);
nor U3982 (N_3982,N_3895,N_3832);
nor U3983 (N_3983,N_3837,N_3816);
nand U3984 (N_3984,N_3888,N_3822);
nand U3985 (N_3985,N_3832,N_3807);
nand U3986 (N_3986,N_3834,N_3838);
nand U3987 (N_3987,N_3815,N_3821);
nor U3988 (N_3988,N_3839,N_3826);
nor U3989 (N_3989,N_3868,N_3829);
and U3990 (N_3990,N_3872,N_3863);
and U3991 (N_3991,N_3852,N_3801);
nor U3992 (N_3992,N_3869,N_3829);
nand U3993 (N_3993,N_3808,N_3816);
xnor U3994 (N_3994,N_3851,N_3817);
xnor U3995 (N_3995,N_3851,N_3805);
nor U3996 (N_3996,N_3847,N_3880);
or U3997 (N_3997,N_3884,N_3845);
or U3998 (N_3998,N_3856,N_3879);
nand U3999 (N_3999,N_3837,N_3859);
xnor U4000 (N_4000,N_3913,N_3990);
or U4001 (N_4001,N_3987,N_3986);
and U4002 (N_4002,N_3957,N_3964);
and U4003 (N_4003,N_3959,N_3996);
or U4004 (N_4004,N_3912,N_3968);
and U4005 (N_4005,N_3908,N_3917);
nor U4006 (N_4006,N_3947,N_3971);
nand U4007 (N_4007,N_3958,N_3906);
nor U4008 (N_4008,N_3978,N_3929);
or U4009 (N_4009,N_3966,N_3902);
or U4010 (N_4010,N_3932,N_3937);
nor U4011 (N_4011,N_3948,N_3994);
nor U4012 (N_4012,N_3928,N_3900);
nor U4013 (N_4013,N_3962,N_3924);
or U4014 (N_4014,N_3931,N_3950);
or U4015 (N_4015,N_3972,N_3998);
and U4016 (N_4016,N_3997,N_3923);
xnor U4017 (N_4017,N_3988,N_3933);
xnor U4018 (N_4018,N_3989,N_3943);
or U4019 (N_4019,N_3979,N_3935);
xor U4020 (N_4020,N_3904,N_3946);
and U4021 (N_4021,N_3903,N_3909);
nor U4022 (N_4022,N_3918,N_3999);
and U4023 (N_4023,N_3963,N_3907);
and U4024 (N_4024,N_3938,N_3955);
or U4025 (N_4025,N_3952,N_3956);
nand U4026 (N_4026,N_3910,N_3981);
nand U4027 (N_4027,N_3991,N_3940);
nor U4028 (N_4028,N_3969,N_3945);
xor U4029 (N_4029,N_3934,N_3965);
or U4030 (N_4030,N_3967,N_3926);
and U4031 (N_4031,N_3980,N_3973);
and U4032 (N_4032,N_3944,N_3914);
nand U4033 (N_4033,N_3954,N_3995);
xor U4034 (N_4034,N_3942,N_3939);
xor U4035 (N_4035,N_3911,N_3919);
nor U4036 (N_4036,N_3925,N_3960);
nor U4037 (N_4037,N_3976,N_3951);
and U4038 (N_4038,N_3941,N_3949);
xnor U4039 (N_4039,N_3927,N_3920);
xnor U4040 (N_4040,N_3984,N_3953);
nand U4041 (N_4041,N_3970,N_3901);
nor U4042 (N_4042,N_3915,N_3974);
nor U4043 (N_4043,N_3936,N_3985);
and U4044 (N_4044,N_3983,N_3916);
and U4045 (N_4045,N_3993,N_3977);
xnor U4046 (N_4046,N_3921,N_3922);
xor U4047 (N_4047,N_3961,N_3992);
nand U4048 (N_4048,N_3905,N_3930);
and U4049 (N_4049,N_3975,N_3982);
nor U4050 (N_4050,N_3946,N_3977);
and U4051 (N_4051,N_3915,N_3920);
nand U4052 (N_4052,N_3966,N_3972);
xor U4053 (N_4053,N_3905,N_3955);
nor U4054 (N_4054,N_3909,N_3992);
and U4055 (N_4055,N_3905,N_3954);
nand U4056 (N_4056,N_3941,N_3994);
xnor U4057 (N_4057,N_3958,N_3945);
and U4058 (N_4058,N_3900,N_3959);
nor U4059 (N_4059,N_3925,N_3921);
and U4060 (N_4060,N_3906,N_3927);
nor U4061 (N_4061,N_3964,N_3978);
xnor U4062 (N_4062,N_3953,N_3964);
xor U4063 (N_4063,N_3908,N_3990);
and U4064 (N_4064,N_3978,N_3980);
or U4065 (N_4065,N_3922,N_3978);
nor U4066 (N_4066,N_3943,N_3944);
or U4067 (N_4067,N_3988,N_3982);
xnor U4068 (N_4068,N_3919,N_3917);
and U4069 (N_4069,N_3989,N_3977);
or U4070 (N_4070,N_3959,N_3987);
nand U4071 (N_4071,N_3965,N_3902);
nor U4072 (N_4072,N_3994,N_3984);
nand U4073 (N_4073,N_3944,N_3901);
nand U4074 (N_4074,N_3996,N_3901);
and U4075 (N_4075,N_3968,N_3929);
nor U4076 (N_4076,N_3946,N_3997);
xnor U4077 (N_4077,N_3904,N_3917);
nand U4078 (N_4078,N_3958,N_3925);
or U4079 (N_4079,N_3986,N_3910);
nor U4080 (N_4080,N_3907,N_3998);
or U4081 (N_4081,N_3952,N_3947);
nor U4082 (N_4082,N_3971,N_3953);
nor U4083 (N_4083,N_3945,N_3939);
nor U4084 (N_4084,N_3974,N_3956);
nand U4085 (N_4085,N_3941,N_3944);
or U4086 (N_4086,N_3900,N_3979);
and U4087 (N_4087,N_3971,N_3941);
or U4088 (N_4088,N_3918,N_3970);
xnor U4089 (N_4089,N_3922,N_3910);
or U4090 (N_4090,N_3983,N_3906);
xor U4091 (N_4091,N_3976,N_3941);
or U4092 (N_4092,N_3924,N_3915);
and U4093 (N_4093,N_3906,N_3940);
xor U4094 (N_4094,N_3926,N_3971);
nand U4095 (N_4095,N_3998,N_3905);
or U4096 (N_4096,N_3917,N_3997);
xor U4097 (N_4097,N_3996,N_3994);
and U4098 (N_4098,N_3970,N_3929);
nor U4099 (N_4099,N_3916,N_3992);
nor U4100 (N_4100,N_4057,N_4066);
or U4101 (N_4101,N_4052,N_4031);
or U4102 (N_4102,N_4019,N_4047);
or U4103 (N_4103,N_4053,N_4004);
and U4104 (N_4104,N_4006,N_4002);
nand U4105 (N_4105,N_4075,N_4060);
and U4106 (N_4106,N_4099,N_4078);
and U4107 (N_4107,N_4042,N_4003);
nand U4108 (N_4108,N_4056,N_4070);
nor U4109 (N_4109,N_4079,N_4067);
nor U4110 (N_4110,N_4008,N_4096);
and U4111 (N_4111,N_4030,N_4058);
or U4112 (N_4112,N_4054,N_4069);
xor U4113 (N_4113,N_4081,N_4029);
or U4114 (N_4114,N_4046,N_4026);
xnor U4115 (N_4115,N_4037,N_4064);
nand U4116 (N_4116,N_4032,N_4010);
or U4117 (N_4117,N_4089,N_4015);
xnor U4118 (N_4118,N_4080,N_4044);
or U4119 (N_4119,N_4041,N_4065);
nor U4120 (N_4120,N_4036,N_4097);
or U4121 (N_4121,N_4023,N_4073);
nand U4122 (N_4122,N_4007,N_4039);
or U4123 (N_4123,N_4033,N_4048);
nand U4124 (N_4124,N_4062,N_4040);
or U4125 (N_4125,N_4074,N_4076);
nor U4126 (N_4126,N_4092,N_4001);
and U4127 (N_4127,N_4024,N_4017);
and U4128 (N_4128,N_4028,N_4011);
nand U4129 (N_4129,N_4025,N_4043);
or U4130 (N_4130,N_4000,N_4093);
nand U4131 (N_4131,N_4071,N_4018);
and U4132 (N_4132,N_4051,N_4049);
nand U4133 (N_4133,N_4055,N_4027);
and U4134 (N_4134,N_4012,N_4072);
or U4135 (N_4135,N_4013,N_4086);
and U4136 (N_4136,N_4085,N_4045);
xor U4137 (N_4137,N_4005,N_4022);
nand U4138 (N_4138,N_4084,N_4020);
nand U4139 (N_4139,N_4090,N_4038);
xor U4140 (N_4140,N_4088,N_4098);
or U4141 (N_4141,N_4014,N_4035);
or U4142 (N_4142,N_4068,N_4059);
and U4143 (N_4143,N_4034,N_4061);
or U4144 (N_4144,N_4095,N_4063);
and U4145 (N_4145,N_4016,N_4091);
nor U4146 (N_4146,N_4009,N_4050);
and U4147 (N_4147,N_4083,N_4082);
xor U4148 (N_4148,N_4077,N_4094);
and U4149 (N_4149,N_4021,N_4087);
nand U4150 (N_4150,N_4055,N_4039);
xor U4151 (N_4151,N_4014,N_4022);
nor U4152 (N_4152,N_4069,N_4045);
xor U4153 (N_4153,N_4066,N_4083);
nor U4154 (N_4154,N_4045,N_4095);
nand U4155 (N_4155,N_4046,N_4068);
nand U4156 (N_4156,N_4071,N_4068);
xor U4157 (N_4157,N_4069,N_4051);
xnor U4158 (N_4158,N_4094,N_4051);
and U4159 (N_4159,N_4064,N_4035);
xnor U4160 (N_4160,N_4077,N_4006);
or U4161 (N_4161,N_4078,N_4076);
nor U4162 (N_4162,N_4082,N_4017);
nor U4163 (N_4163,N_4059,N_4019);
nor U4164 (N_4164,N_4089,N_4072);
nor U4165 (N_4165,N_4010,N_4088);
and U4166 (N_4166,N_4026,N_4087);
and U4167 (N_4167,N_4061,N_4054);
nor U4168 (N_4168,N_4031,N_4014);
nor U4169 (N_4169,N_4063,N_4045);
xnor U4170 (N_4170,N_4057,N_4042);
or U4171 (N_4171,N_4073,N_4020);
nor U4172 (N_4172,N_4096,N_4015);
xor U4173 (N_4173,N_4041,N_4022);
nor U4174 (N_4174,N_4067,N_4069);
nand U4175 (N_4175,N_4038,N_4002);
nor U4176 (N_4176,N_4030,N_4084);
or U4177 (N_4177,N_4084,N_4032);
xnor U4178 (N_4178,N_4081,N_4066);
nor U4179 (N_4179,N_4097,N_4044);
nor U4180 (N_4180,N_4004,N_4011);
nand U4181 (N_4181,N_4064,N_4046);
and U4182 (N_4182,N_4066,N_4092);
and U4183 (N_4183,N_4019,N_4062);
or U4184 (N_4184,N_4043,N_4095);
xnor U4185 (N_4185,N_4018,N_4021);
xnor U4186 (N_4186,N_4083,N_4005);
or U4187 (N_4187,N_4049,N_4034);
nor U4188 (N_4188,N_4040,N_4084);
and U4189 (N_4189,N_4032,N_4087);
nand U4190 (N_4190,N_4079,N_4096);
nor U4191 (N_4191,N_4055,N_4049);
nor U4192 (N_4192,N_4086,N_4037);
nand U4193 (N_4193,N_4000,N_4002);
nand U4194 (N_4194,N_4083,N_4038);
and U4195 (N_4195,N_4036,N_4081);
nor U4196 (N_4196,N_4002,N_4001);
xnor U4197 (N_4197,N_4015,N_4064);
nor U4198 (N_4198,N_4026,N_4040);
and U4199 (N_4199,N_4028,N_4025);
and U4200 (N_4200,N_4166,N_4132);
xnor U4201 (N_4201,N_4106,N_4181);
and U4202 (N_4202,N_4104,N_4133);
and U4203 (N_4203,N_4177,N_4127);
nand U4204 (N_4204,N_4100,N_4175);
xor U4205 (N_4205,N_4123,N_4163);
and U4206 (N_4206,N_4179,N_4178);
nand U4207 (N_4207,N_4151,N_4190);
nor U4208 (N_4208,N_4108,N_4182);
xnor U4209 (N_4209,N_4116,N_4176);
nor U4210 (N_4210,N_4172,N_4120);
and U4211 (N_4211,N_4168,N_4145);
xnor U4212 (N_4212,N_4126,N_4118);
or U4213 (N_4213,N_4156,N_4189);
nand U4214 (N_4214,N_4186,N_4131);
nor U4215 (N_4215,N_4192,N_4152);
or U4216 (N_4216,N_4187,N_4102);
nand U4217 (N_4217,N_4155,N_4184);
nor U4218 (N_4218,N_4160,N_4142);
nand U4219 (N_4219,N_4173,N_4135);
nand U4220 (N_4220,N_4134,N_4113);
xnor U4221 (N_4221,N_4146,N_4196);
or U4222 (N_4222,N_4169,N_4107);
and U4223 (N_4223,N_4147,N_4101);
nor U4224 (N_4224,N_4194,N_4115);
nand U4225 (N_4225,N_4124,N_4125);
xor U4226 (N_4226,N_4140,N_4138);
xnor U4227 (N_4227,N_4150,N_4162);
and U4228 (N_4228,N_4170,N_4191);
or U4229 (N_4229,N_4171,N_4141);
nand U4230 (N_4230,N_4159,N_4109);
nor U4231 (N_4231,N_4185,N_4157);
and U4232 (N_4232,N_4158,N_4129);
and U4233 (N_4233,N_4105,N_4154);
xor U4234 (N_4234,N_4183,N_4122);
nor U4235 (N_4235,N_4193,N_4117);
nor U4236 (N_4236,N_4165,N_4139);
nor U4237 (N_4237,N_4103,N_4111);
and U4238 (N_4238,N_4128,N_4153);
xnor U4239 (N_4239,N_4119,N_4114);
xnor U4240 (N_4240,N_4180,N_4121);
and U4241 (N_4241,N_4197,N_4199);
or U4242 (N_4242,N_4149,N_4195);
xor U4243 (N_4243,N_4167,N_4112);
or U4244 (N_4244,N_4130,N_4161);
nand U4245 (N_4245,N_4143,N_4110);
nor U4246 (N_4246,N_4164,N_4136);
or U4247 (N_4247,N_4137,N_4198);
nand U4248 (N_4248,N_4144,N_4174);
nor U4249 (N_4249,N_4148,N_4188);
and U4250 (N_4250,N_4175,N_4171);
and U4251 (N_4251,N_4167,N_4152);
nor U4252 (N_4252,N_4167,N_4119);
and U4253 (N_4253,N_4170,N_4125);
or U4254 (N_4254,N_4140,N_4164);
xor U4255 (N_4255,N_4119,N_4109);
nor U4256 (N_4256,N_4145,N_4187);
nand U4257 (N_4257,N_4119,N_4123);
xor U4258 (N_4258,N_4152,N_4151);
nor U4259 (N_4259,N_4145,N_4165);
or U4260 (N_4260,N_4198,N_4167);
or U4261 (N_4261,N_4178,N_4183);
or U4262 (N_4262,N_4157,N_4179);
or U4263 (N_4263,N_4131,N_4130);
nand U4264 (N_4264,N_4175,N_4103);
or U4265 (N_4265,N_4100,N_4165);
nor U4266 (N_4266,N_4168,N_4108);
or U4267 (N_4267,N_4182,N_4162);
or U4268 (N_4268,N_4155,N_4119);
nor U4269 (N_4269,N_4125,N_4139);
xnor U4270 (N_4270,N_4170,N_4143);
nand U4271 (N_4271,N_4140,N_4176);
xnor U4272 (N_4272,N_4107,N_4130);
xor U4273 (N_4273,N_4180,N_4142);
xor U4274 (N_4274,N_4158,N_4143);
nand U4275 (N_4275,N_4127,N_4114);
or U4276 (N_4276,N_4103,N_4198);
or U4277 (N_4277,N_4122,N_4156);
nand U4278 (N_4278,N_4178,N_4131);
and U4279 (N_4279,N_4119,N_4170);
and U4280 (N_4280,N_4192,N_4129);
nand U4281 (N_4281,N_4171,N_4179);
xor U4282 (N_4282,N_4118,N_4134);
nor U4283 (N_4283,N_4190,N_4179);
nand U4284 (N_4284,N_4185,N_4199);
nor U4285 (N_4285,N_4141,N_4132);
nand U4286 (N_4286,N_4195,N_4155);
xnor U4287 (N_4287,N_4122,N_4111);
nor U4288 (N_4288,N_4132,N_4124);
xnor U4289 (N_4289,N_4125,N_4123);
xor U4290 (N_4290,N_4174,N_4125);
xor U4291 (N_4291,N_4168,N_4176);
nand U4292 (N_4292,N_4137,N_4101);
nor U4293 (N_4293,N_4133,N_4170);
xnor U4294 (N_4294,N_4157,N_4163);
and U4295 (N_4295,N_4194,N_4193);
and U4296 (N_4296,N_4126,N_4197);
xor U4297 (N_4297,N_4134,N_4123);
xor U4298 (N_4298,N_4162,N_4184);
xnor U4299 (N_4299,N_4154,N_4192);
xor U4300 (N_4300,N_4211,N_4200);
nor U4301 (N_4301,N_4239,N_4285);
nor U4302 (N_4302,N_4246,N_4268);
nor U4303 (N_4303,N_4298,N_4267);
xnor U4304 (N_4304,N_4234,N_4244);
xnor U4305 (N_4305,N_4254,N_4229);
or U4306 (N_4306,N_4208,N_4210);
nand U4307 (N_4307,N_4209,N_4262);
xnor U4308 (N_4308,N_4201,N_4226);
and U4309 (N_4309,N_4271,N_4214);
xor U4310 (N_4310,N_4274,N_4205);
xor U4311 (N_4311,N_4222,N_4223);
nand U4312 (N_4312,N_4240,N_4250);
xor U4313 (N_4313,N_4213,N_4238);
nor U4314 (N_4314,N_4230,N_4237);
and U4315 (N_4315,N_4277,N_4259);
xnor U4316 (N_4316,N_4272,N_4288);
nor U4317 (N_4317,N_4241,N_4235);
nor U4318 (N_4318,N_4290,N_4270);
or U4319 (N_4319,N_4257,N_4261);
and U4320 (N_4320,N_4212,N_4275);
nand U4321 (N_4321,N_4282,N_4218);
nand U4322 (N_4322,N_4292,N_4203);
nor U4323 (N_4323,N_4278,N_4221);
nor U4324 (N_4324,N_4242,N_4202);
nand U4325 (N_4325,N_4264,N_4291);
nor U4326 (N_4326,N_4299,N_4258);
nor U4327 (N_4327,N_4248,N_4279);
and U4328 (N_4328,N_4289,N_4269);
xor U4329 (N_4329,N_4219,N_4287);
or U4330 (N_4330,N_4228,N_4255);
and U4331 (N_4331,N_4245,N_4243);
nand U4332 (N_4332,N_4232,N_4293);
nor U4333 (N_4333,N_4236,N_4296);
xor U4334 (N_4334,N_4294,N_4247);
nand U4335 (N_4335,N_4207,N_4280);
and U4336 (N_4336,N_4260,N_4216);
and U4337 (N_4337,N_4252,N_4224);
and U4338 (N_4338,N_4215,N_4295);
and U4339 (N_4339,N_4283,N_4227);
nor U4340 (N_4340,N_4206,N_4276);
and U4341 (N_4341,N_4249,N_4286);
nand U4342 (N_4342,N_4263,N_4297);
and U4343 (N_4343,N_4266,N_4253);
or U4344 (N_4344,N_4251,N_4233);
nor U4345 (N_4345,N_4220,N_4284);
and U4346 (N_4346,N_4273,N_4256);
or U4347 (N_4347,N_4265,N_4204);
and U4348 (N_4348,N_4225,N_4217);
and U4349 (N_4349,N_4281,N_4231);
nand U4350 (N_4350,N_4222,N_4289);
and U4351 (N_4351,N_4281,N_4292);
nand U4352 (N_4352,N_4276,N_4292);
nand U4353 (N_4353,N_4261,N_4208);
nor U4354 (N_4354,N_4292,N_4230);
xor U4355 (N_4355,N_4231,N_4206);
nor U4356 (N_4356,N_4246,N_4201);
xor U4357 (N_4357,N_4296,N_4207);
nor U4358 (N_4358,N_4271,N_4239);
nand U4359 (N_4359,N_4295,N_4259);
nand U4360 (N_4360,N_4267,N_4295);
nor U4361 (N_4361,N_4280,N_4264);
nor U4362 (N_4362,N_4234,N_4293);
and U4363 (N_4363,N_4269,N_4280);
xor U4364 (N_4364,N_4227,N_4272);
nor U4365 (N_4365,N_4218,N_4293);
nor U4366 (N_4366,N_4243,N_4276);
nor U4367 (N_4367,N_4234,N_4205);
and U4368 (N_4368,N_4280,N_4218);
nor U4369 (N_4369,N_4278,N_4260);
xor U4370 (N_4370,N_4267,N_4241);
nor U4371 (N_4371,N_4208,N_4277);
nor U4372 (N_4372,N_4222,N_4234);
nor U4373 (N_4373,N_4296,N_4239);
xnor U4374 (N_4374,N_4255,N_4219);
nand U4375 (N_4375,N_4207,N_4279);
and U4376 (N_4376,N_4217,N_4212);
or U4377 (N_4377,N_4225,N_4269);
nand U4378 (N_4378,N_4201,N_4212);
nor U4379 (N_4379,N_4235,N_4216);
and U4380 (N_4380,N_4242,N_4241);
xnor U4381 (N_4381,N_4259,N_4245);
xnor U4382 (N_4382,N_4202,N_4298);
and U4383 (N_4383,N_4216,N_4275);
nor U4384 (N_4384,N_4294,N_4279);
or U4385 (N_4385,N_4294,N_4211);
or U4386 (N_4386,N_4206,N_4224);
nand U4387 (N_4387,N_4221,N_4255);
xnor U4388 (N_4388,N_4234,N_4211);
nor U4389 (N_4389,N_4230,N_4253);
nor U4390 (N_4390,N_4275,N_4251);
nor U4391 (N_4391,N_4253,N_4286);
xnor U4392 (N_4392,N_4231,N_4209);
nor U4393 (N_4393,N_4255,N_4258);
xor U4394 (N_4394,N_4246,N_4230);
nand U4395 (N_4395,N_4220,N_4230);
or U4396 (N_4396,N_4240,N_4212);
nand U4397 (N_4397,N_4204,N_4224);
or U4398 (N_4398,N_4263,N_4226);
or U4399 (N_4399,N_4285,N_4203);
nor U4400 (N_4400,N_4374,N_4310);
nand U4401 (N_4401,N_4349,N_4323);
nand U4402 (N_4402,N_4370,N_4367);
xor U4403 (N_4403,N_4368,N_4381);
nand U4404 (N_4404,N_4319,N_4372);
nand U4405 (N_4405,N_4309,N_4377);
nand U4406 (N_4406,N_4376,N_4341);
and U4407 (N_4407,N_4340,N_4383);
nor U4408 (N_4408,N_4318,N_4311);
nand U4409 (N_4409,N_4327,N_4396);
nor U4410 (N_4410,N_4388,N_4354);
nand U4411 (N_4411,N_4325,N_4355);
xor U4412 (N_4412,N_4317,N_4342);
xor U4413 (N_4413,N_4352,N_4316);
xnor U4414 (N_4414,N_4324,N_4387);
and U4415 (N_4415,N_4303,N_4330);
and U4416 (N_4416,N_4307,N_4305);
and U4417 (N_4417,N_4371,N_4380);
xor U4418 (N_4418,N_4399,N_4395);
nand U4419 (N_4419,N_4382,N_4326);
nand U4420 (N_4420,N_4300,N_4308);
nor U4421 (N_4421,N_4321,N_4302);
or U4422 (N_4422,N_4333,N_4373);
and U4423 (N_4423,N_4358,N_4356);
xor U4424 (N_4424,N_4391,N_4362);
nand U4425 (N_4425,N_4312,N_4347);
and U4426 (N_4426,N_4304,N_4301);
or U4427 (N_4427,N_4331,N_4345);
or U4428 (N_4428,N_4379,N_4329);
nor U4429 (N_4429,N_4366,N_4365);
xnor U4430 (N_4430,N_4397,N_4306);
nor U4431 (N_4431,N_4313,N_4328);
nor U4432 (N_4432,N_4359,N_4353);
nor U4433 (N_4433,N_4363,N_4393);
and U4434 (N_4434,N_4378,N_4351);
xor U4435 (N_4435,N_4369,N_4338);
nand U4436 (N_4436,N_4392,N_4364);
nand U4437 (N_4437,N_4315,N_4337);
nor U4438 (N_4438,N_4336,N_4361);
nor U4439 (N_4439,N_4386,N_4398);
or U4440 (N_4440,N_4389,N_4314);
nand U4441 (N_4441,N_4322,N_4339);
nand U4442 (N_4442,N_4394,N_4320);
or U4443 (N_4443,N_4334,N_4344);
xor U4444 (N_4444,N_4346,N_4348);
xnor U4445 (N_4445,N_4384,N_4375);
and U4446 (N_4446,N_4332,N_4385);
xor U4447 (N_4447,N_4343,N_4350);
and U4448 (N_4448,N_4360,N_4357);
nor U4449 (N_4449,N_4390,N_4335);
nand U4450 (N_4450,N_4326,N_4367);
or U4451 (N_4451,N_4369,N_4314);
xor U4452 (N_4452,N_4365,N_4372);
nor U4453 (N_4453,N_4396,N_4306);
nor U4454 (N_4454,N_4385,N_4374);
xnor U4455 (N_4455,N_4395,N_4362);
and U4456 (N_4456,N_4399,N_4369);
and U4457 (N_4457,N_4349,N_4359);
and U4458 (N_4458,N_4361,N_4320);
nor U4459 (N_4459,N_4396,N_4344);
nor U4460 (N_4460,N_4321,N_4351);
or U4461 (N_4461,N_4320,N_4316);
or U4462 (N_4462,N_4352,N_4349);
nor U4463 (N_4463,N_4367,N_4316);
nand U4464 (N_4464,N_4312,N_4355);
and U4465 (N_4465,N_4329,N_4301);
nor U4466 (N_4466,N_4325,N_4326);
nor U4467 (N_4467,N_4311,N_4364);
xnor U4468 (N_4468,N_4383,N_4302);
and U4469 (N_4469,N_4388,N_4396);
or U4470 (N_4470,N_4316,N_4390);
and U4471 (N_4471,N_4359,N_4379);
and U4472 (N_4472,N_4353,N_4322);
or U4473 (N_4473,N_4362,N_4328);
xnor U4474 (N_4474,N_4305,N_4365);
and U4475 (N_4475,N_4387,N_4392);
or U4476 (N_4476,N_4303,N_4331);
nand U4477 (N_4477,N_4352,N_4353);
xor U4478 (N_4478,N_4330,N_4332);
xnor U4479 (N_4479,N_4385,N_4366);
and U4480 (N_4480,N_4353,N_4306);
and U4481 (N_4481,N_4391,N_4331);
or U4482 (N_4482,N_4320,N_4389);
nand U4483 (N_4483,N_4304,N_4313);
and U4484 (N_4484,N_4316,N_4355);
nand U4485 (N_4485,N_4304,N_4355);
nand U4486 (N_4486,N_4381,N_4313);
xnor U4487 (N_4487,N_4327,N_4306);
nand U4488 (N_4488,N_4364,N_4388);
and U4489 (N_4489,N_4388,N_4351);
nand U4490 (N_4490,N_4323,N_4322);
nor U4491 (N_4491,N_4301,N_4382);
xnor U4492 (N_4492,N_4305,N_4373);
nor U4493 (N_4493,N_4301,N_4376);
xnor U4494 (N_4494,N_4372,N_4395);
and U4495 (N_4495,N_4383,N_4328);
xnor U4496 (N_4496,N_4306,N_4322);
xnor U4497 (N_4497,N_4339,N_4316);
xnor U4498 (N_4498,N_4391,N_4324);
nand U4499 (N_4499,N_4300,N_4313);
xnor U4500 (N_4500,N_4439,N_4440);
xor U4501 (N_4501,N_4436,N_4491);
or U4502 (N_4502,N_4463,N_4461);
nand U4503 (N_4503,N_4464,N_4422);
nand U4504 (N_4504,N_4465,N_4434);
or U4505 (N_4505,N_4495,N_4477);
nand U4506 (N_4506,N_4494,N_4424);
or U4507 (N_4507,N_4487,N_4474);
nor U4508 (N_4508,N_4414,N_4453);
and U4509 (N_4509,N_4431,N_4409);
nand U4510 (N_4510,N_4444,N_4475);
nand U4511 (N_4511,N_4407,N_4432);
nor U4512 (N_4512,N_4468,N_4498);
or U4513 (N_4513,N_4411,N_4427);
nor U4514 (N_4514,N_4441,N_4403);
xor U4515 (N_4515,N_4447,N_4460);
or U4516 (N_4516,N_4479,N_4466);
nor U4517 (N_4517,N_4406,N_4459);
nor U4518 (N_4518,N_4493,N_4421);
and U4519 (N_4519,N_4428,N_4476);
or U4520 (N_4520,N_4449,N_4419);
nand U4521 (N_4521,N_4426,N_4442);
nor U4522 (N_4522,N_4412,N_4492);
xnor U4523 (N_4523,N_4481,N_4413);
and U4524 (N_4524,N_4482,N_4451);
or U4525 (N_4525,N_4445,N_4490);
xor U4526 (N_4526,N_4472,N_4408);
nor U4527 (N_4527,N_4401,N_4454);
xor U4528 (N_4528,N_4471,N_4448);
xor U4529 (N_4529,N_4499,N_4497);
or U4530 (N_4530,N_4450,N_4417);
nand U4531 (N_4531,N_4470,N_4433);
xor U4532 (N_4532,N_4402,N_4437);
and U4533 (N_4533,N_4473,N_4452);
nand U4534 (N_4534,N_4404,N_4446);
xnor U4535 (N_4535,N_4400,N_4423);
xnor U4536 (N_4536,N_4480,N_4429);
xor U4537 (N_4537,N_4458,N_4410);
nor U4538 (N_4538,N_4469,N_4405);
nor U4539 (N_4539,N_4486,N_4455);
nor U4540 (N_4540,N_4467,N_4415);
nor U4541 (N_4541,N_4484,N_4425);
xor U4542 (N_4542,N_4457,N_4478);
and U4543 (N_4543,N_4485,N_4418);
xnor U4544 (N_4544,N_4489,N_4443);
and U4545 (N_4545,N_4488,N_4435);
or U4546 (N_4546,N_4483,N_4430);
or U4547 (N_4547,N_4416,N_4456);
nand U4548 (N_4548,N_4438,N_4420);
nand U4549 (N_4549,N_4462,N_4496);
xor U4550 (N_4550,N_4443,N_4475);
and U4551 (N_4551,N_4495,N_4448);
or U4552 (N_4552,N_4488,N_4402);
or U4553 (N_4553,N_4486,N_4420);
and U4554 (N_4554,N_4437,N_4471);
nor U4555 (N_4555,N_4458,N_4423);
xnor U4556 (N_4556,N_4419,N_4483);
or U4557 (N_4557,N_4446,N_4487);
xor U4558 (N_4558,N_4445,N_4467);
nor U4559 (N_4559,N_4460,N_4404);
or U4560 (N_4560,N_4437,N_4410);
xor U4561 (N_4561,N_4468,N_4426);
xor U4562 (N_4562,N_4411,N_4424);
nor U4563 (N_4563,N_4490,N_4405);
or U4564 (N_4564,N_4401,N_4427);
nor U4565 (N_4565,N_4436,N_4445);
nor U4566 (N_4566,N_4417,N_4471);
and U4567 (N_4567,N_4434,N_4442);
nand U4568 (N_4568,N_4439,N_4409);
and U4569 (N_4569,N_4444,N_4459);
xor U4570 (N_4570,N_4475,N_4479);
nand U4571 (N_4571,N_4413,N_4477);
and U4572 (N_4572,N_4481,N_4485);
xor U4573 (N_4573,N_4467,N_4433);
or U4574 (N_4574,N_4405,N_4444);
nand U4575 (N_4575,N_4446,N_4449);
nand U4576 (N_4576,N_4402,N_4493);
nand U4577 (N_4577,N_4457,N_4417);
nor U4578 (N_4578,N_4409,N_4468);
xnor U4579 (N_4579,N_4491,N_4435);
or U4580 (N_4580,N_4452,N_4488);
xnor U4581 (N_4581,N_4401,N_4475);
nand U4582 (N_4582,N_4425,N_4492);
or U4583 (N_4583,N_4481,N_4456);
nor U4584 (N_4584,N_4478,N_4469);
nor U4585 (N_4585,N_4413,N_4496);
or U4586 (N_4586,N_4457,N_4406);
nor U4587 (N_4587,N_4457,N_4439);
xor U4588 (N_4588,N_4459,N_4422);
nor U4589 (N_4589,N_4450,N_4433);
nand U4590 (N_4590,N_4489,N_4480);
and U4591 (N_4591,N_4450,N_4476);
nor U4592 (N_4592,N_4471,N_4436);
or U4593 (N_4593,N_4430,N_4464);
nor U4594 (N_4594,N_4413,N_4425);
xnor U4595 (N_4595,N_4470,N_4429);
xor U4596 (N_4596,N_4437,N_4416);
or U4597 (N_4597,N_4477,N_4498);
xor U4598 (N_4598,N_4492,N_4453);
nor U4599 (N_4599,N_4489,N_4449);
and U4600 (N_4600,N_4559,N_4580);
nand U4601 (N_4601,N_4586,N_4528);
nor U4602 (N_4602,N_4508,N_4506);
or U4603 (N_4603,N_4544,N_4573);
and U4604 (N_4604,N_4530,N_4569);
or U4605 (N_4605,N_4519,N_4572);
xor U4606 (N_4606,N_4574,N_4517);
xor U4607 (N_4607,N_4533,N_4501);
xor U4608 (N_4608,N_4550,N_4598);
xnor U4609 (N_4609,N_4513,N_4520);
and U4610 (N_4610,N_4595,N_4583);
and U4611 (N_4611,N_4525,N_4576);
xnor U4612 (N_4612,N_4581,N_4518);
xnor U4613 (N_4613,N_4557,N_4534);
nand U4614 (N_4614,N_4511,N_4547);
and U4615 (N_4615,N_4582,N_4535);
nor U4616 (N_4616,N_4561,N_4510);
nor U4617 (N_4617,N_4546,N_4504);
and U4618 (N_4618,N_4579,N_4521);
nand U4619 (N_4619,N_4577,N_4512);
nand U4620 (N_4620,N_4503,N_4560);
or U4621 (N_4621,N_4555,N_4541);
and U4622 (N_4622,N_4543,N_4502);
nand U4623 (N_4623,N_4570,N_4542);
or U4624 (N_4624,N_4523,N_4509);
or U4625 (N_4625,N_4532,N_4522);
xor U4626 (N_4626,N_4526,N_4558);
xnor U4627 (N_4627,N_4578,N_4539);
nand U4628 (N_4628,N_4568,N_4537);
nor U4629 (N_4629,N_4590,N_4500);
and U4630 (N_4630,N_4571,N_4548);
nand U4631 (N_4631,N_4584,N_4566);
or U4632 (N_4632,N_4552,N_4593);
and U4633 (N_4633,N_4575,N_4554);
or U4634 (N_4634,N_4591,N_4563);
xnor U4635 (N_4635,N_4592,N_4538);
nand U4636 (N_4636,N_4556,N_4587);
or U4637 (N_4637,N_4527,N_4588);
nor U4638 (N_4638,N_4540,N_4516);
or U4639 (N_4639,N_4549,N_4545);
and U4640 (N_4640,N_4585,N_4514);
xnor U4641 (N_4641,N_4524,N_4536);
nand U4642 (N_4642,N_4507,N_4599);
nor U4643 (N_4643,N_4515,N_4562);
nor U4644 (N_4644,N_4551,N_4589);
nor U4645 (N_4645,N_4531,N_4553);
nor U4646 (N_4646,N_4567,N_4564);
and U4647 (N_4647,N_4505,N_4597);
or U4648 (N_4648,N_4596,N_4594);
or U4649 (N_4649,N_4529,N_4565);
and U4650 (N_4650,N_4570,N_4578);
or U4651 (N_4651,N_4596,N_4530);
and U4652 (N_4652,N_4593,N_4573);
xnor U4653 (N_4653,N_4563,N_4519);
xor U4654 (N_4654,N_4513,N_4516);
xor U4655 (N_4655,N_4564,N_4538);
xor U4656 (N_4656,N_4533,N_4550);
or U4657 (N_4657,N_4514,N_4506);
nand U4658 (N_4658,N_4540,N_4505);
or U4659 (N_4659,N_4572,N_4555);
or U4660 (N_4660,N_4581,N_4511);
nand U4661 (N_4661,N_4590,N_4575);
nand U4662 (N_4662,N_4500,N_4533);
nor U4663 (N_4663,N_4505,N_4551);
nand U4664 (N_4664,N_4527,N_4584);
nand U4665 (N_4665,N_4564,N_4529);
nor U4666 (N_4666,N_4565,N_4595);
nand U4667 (N_4667,N_4584,N_4544);
nor U4668 (N_4668,N_4590,N_4556);
and U4669 (N_4669,N_4550,N_4581);
nand U4670 (N_4670,N_4507,N_4540);
or U4671 (N_4671,N_4580,N_4577);
and U4672 (N_4672,N_4568,N_4501);
and U4673 (N_4673,N_4513,N_4555);
and U4674 (N_4674,N_4543,N_4527);
and U4675 (N_4675,N_4586,N_4547);
nand U4676 (N_4676,N_4549,N_4598);
or U4677 (N_4677,N_4532,N_4570);
nor U4678 (N_4678,N_4546,N_4581);
and U4679 (N_4679,N_4588,N_4524);
and U4680 (N_4680,N_4540,N_4524);
and U4681 (N_4681,N_4561,N_4558);
and U4682 (N_4682,N_4520,N_4555);
and U4683 (N_4683,N_4510,N_4542);
xor U4684 (N_4684,N_4573,N_4580);
nor U4685 (N_4685,N_4516,N_4508);
xor U4686 (N_4686,N_4519,N_4504);
or U4687 (N_4687,N_4581,N_4591);
nand U4688 (N_4688,N_4521,N_4527);
xnor U4689 (N_4689,N_4590,N_4539);
or U4690 (N_4690,N_4598,N_4574);
nand U4691 (N_4691,N_4555,N_4525);
xnor U4692 (N_4692,N_4545,N_4561);
or U4693 (N_4693,N_4572,N_4501);
xnor U4694 (N_4694,N_4542,N_4547);
xor U4695 (N_4695,N_4557,N_4518);
or U4696 (N_4696,N_4527,N_4559);
nor U4697 (N_4697,N_4554,N_4597);
nand U4698 (N_4698,N_4591,N_4558);
nor U4699 (N_4699,N_4529,N_4514);
nand U4700 (N_4700,N_4654,N_4636);
and U4701 (N_4701,N_4645,N_4646);
or U4702 (N_4702,N_4621,N_4675);
nor U4703 (N_4703,N_4660,N_4626);
and U4704 (N_4704,N_4663,N_4624);
nand U4705 (N_4705,N_4604,N_4616);
and U4706 (N_4706,N_4631,N_4644);
or U4707 (N_4707,N_4694,N_4659);
nor U4708 (N_4708,N_4674,N_4602);
and U4709 (N_4709,N_4685,N_4651);
nand U4710 (N_4710,N_4656,N_4672);
and U4711 (N_4711,N_4669,N_4606);
xnor U4712 (N_4712,N_4601,N_4623);
and U4713 (N_4713,N_4658,N_4670);
or U4714 (N_4714,N_4600,N_4680);
nor U4715 (N_4715,N_4633,N_4643);
nand U4716 (N_4716,N_4691,N_4678);
and U4717 (N_4717,N_4639,N_4648);
nand U4718 (N_4718,N_4650,N_4619);
and U4719 (N_4719,N_4695,N_4668);
nand U4720 (N_4720,N_4611,N_4687);
nand U4721 (N_4721,N_4622,N_4618);
xor U4722 (N_4722,N_4613,N_4630);
and U4723 (N_4723,N_4665,N_4693);
xnor U4724 (N_4724,N_4649,N_4677);
or U4725 (N_4725,N_4664,N_4676);
nand U4726 (N_4726,N_4666,N_4615);
and U4727 (N_4727,N_4608,N_4684);
xor U4728 (N_4728,N_4653,N_4667);
xor U4729 (N_4729,N_4699,N_4697);
nand U4730 (N_4730,N_4657,N_4610);
and U4731 (N_4731,N_4637,N_4632);
or U4732 (N_4732,N_4688,N_4692);
nor U4733 (N_4733,N_4661,N_4690);
nand U4734 (N_4734,N_4641,N_4605);
or U4735 (N_4735,N_4635,N_4629);
xnor U4736 (N_4736,N_4698,N_4683);
and U4737 (N_4737,N_4620,N_4673);
nand U4738 (N_4738,N_4603,N_4607);
and U4739 (N_4739,N_4640,N_4682);
or U4740 (N_4740,N_4679,N_4627);
or U4741 (N_4741,N_4612,N_4625);
and U4742 (N_4742,N_4662,N_4696);
and U4743 (N_4743,N_4628,N_4609);
nor U4744 (N_4744,N_4686,N_4634);
nor U4745 (N_4745,N_4671,N_4681);
nand U4746 (N_4746,N_4689,N_4647);
nand U4747 (N_4747,N_4614,N_4655);
nor U4748 (N_4748,N_4642,N_4617);
nand U4749 (N_4749,N_4638,N_4652);
nor U4750 (N_4750,N_4693,N_4611);
xnor U4751 (N_4751,N_4614,N_4644);
nand U4752 (N_4752,N_4629,N_4642);
xnor U4753 (N_4753,N_4634,N_4671);
xnor U4754 (N_4754,N_4656,N_4602);
or U4755 (N_4755,N_4657,N_4645);
nor U4756 (N_4756,N_4619,N_4656);
xor U4757 (N_4757,N_4667,N_4657);
nor U4758 (N_4758,N_4644,N_4695);
or U4759 (N_4759,N_4636,N_4685);
nor U4760 (N_4760,N_4657,N_4677);
or U4761 (N_4761,N_4611,N_4627);
nor U4762 (N_4762,N_4689,N_4617);
nor U4763 (N_4763,N_4649,N_4662);
nand U4764 (N_4764,N_4605,N_4647);
xnor U4765 (N_4765,N_4630,N_4659);
nand U4766 (N_4766,N_4614,N_4627);
nand U4767 (N_4767,N_4654,N_4664);
or U4768 (N_4768,N_4615,N_4622);
xnor U4769 (N_4769,N_4606,N_4680);
xnor U4770 (N_4770,N_4674,N_4683);
xnor U4771 (N_4771,N_4693,N_4675);
and U4772 (N_4772,N_4699,N_4607);
and U4773 (N_4773,N_4624,N_4620);
and U4774 (N_4774,N_4685,N_4697);
and U4775 (N_4775,N_4645,N_4671);
or U4776 (N_4776,N_4682,N_4681);
nand U4777 (N_4777,N_4664,N_4611);
xor U4778 (N_4778,N_4692,N_4630);
nor U4779 (N_4779,N_4661,N_4643);
and U4780 (N_4780,N_4676,N_4606);
and U4781 (N_4781,N_4633,N_4682);
and U4782 (N_4782,N_4672,N_4664);
or U4783 (N_4783,N_4629,N_4621);
nand U4784 (N_4784,N_4681,N_4676);
and U4785 (N_4785,N_4601,N_4618);
xnor U4786 (N_4786,N_4633,N_4639);
or U4787 (N_4787,N_4679,N_4660);
nand U4788 (N_4788,N_4674,N_4672);
nand U4789 (N_4789,N_4675,N_4668);
nor U4790 (N_4790,N_4610,N_4660);
nand U4791 (N_4791,N_4687,N_4641);
xor U4792 (N_4792,N_4615,N_4605);
and U4793 (N_4793,N_4627,N_4629);
xnor U4794 (N_4794,N_4678,N_4631);
and U4795 (N_4795,N_4667,N_4618);
nand U4796 (N_4796,N_4697,N_4677);
nand U4797 (N_4797,N_4650,N_4690);
or U4798 (N_4798,N_4616,N_4621);
nor U4799 (N_4799,N_4685,N_4609);
and U4800 (N_4800,N_4755,N_4746);
nor U4801 (N_4801,N_4791,N_4738);
or U4802 (N_4802,N_4756,N_4704);
and U4803 (N_4803,N_4757,N_4781);
or U4804 (N_4804,N_4785,N_4705);
nand U4805 (N_4805,N_4772,N_4742);
nor U4806 (N_4806,N_4725,N_4797);
and U4807 (N_4807,N_4749,N_4744);
nor U4808 (N_4808,N_4778,N_4761);
and U4809 (N_4809,N_4707,N_4721);
xnor U4810 (N_4810,N_4736,N_4776);
and U4811 (N_4811,N_4711,N_4771);
xnor U4812 (N_4812,N_4799,N_4795);
nor U4813 (N_4813,N_4766,N_4775);
and U4814 (N_4814,N_4726,N_4793);
and U4815 (N_4815,N_4794,N_4729);
and U4816 (N_4816,N_4740,N_4722);
or U4817 (N_4817,N_4782,N_4724);
xnor U4818 (N_4818,N_4703,N_4706);
and U4819 (N_4819,N_4768,N_4759);
or U4820 (N_4820,N_4741,N_4714);
nand U4821 (N_4821,N_4700,N_4734);
and U4822 (N_4822,N_4730,N_4787);
nand U4823 (N_4823,N_4709,N_4710);
nand U4824 (N_4824,N_4779,N_4780);
and U4825 (N_4825,N_4777,N_4789);
nand U4826 (N_4826,N_4760,N_4701);
xor U4827 (N_4827,N_4753,N_4718);
nor U4828 (N_4828,N_4735,N_4720);
xor U4829 (N_4829,N_4765,N_4716);
xor U4830 (N_4830,N_4712,N_4739);
nand U4831 (N_4831,N_4737,N_4748);
xor U4832 (N_4832,N_4732,N_4790);
and U4833 (N_4833,N_4796,N_4702);
and U4834 (N_4834,N_4727,N_4728);
xnor U4835 (N_4835,N_4786,N_4763);
nand U4836 (N_4836,N_4715,N_4750);
and U4837 (N_4837,N_4798,N_4773);
and U4838 (N_4838,N_4752,N_4764);
or U4839 (N_4839,N_4719,N_4770);
and U4840 (N_4840,N_4751,N_4758);
or U4841 (N_4841,N_4792,N_4769);
nand U4842 (N_4842,N_4745,N_4754);
nand U4843 (N_4843,N_4784,N_4783);
xnor U4844 (N_4844,N_4774,N_4733);
xnor U4845 (N_4845,N_4731,N_4743);
and U4846 (N_4846,N_4747,N_4708);
nor U4847 (N_4847,N_4788,N_4713);
xnor U4848 (N_4848,N_4723,N_4762);
and U4849 (N_4849,N_4717,N_4767);
nor U4850 (N_4850,N_4740,N_4716);
xnor U4851 (N_4851,N_4785,N_4783);
and U4852 (N_4852,N_4746,N_4728);
xor U4853 (N_4853,N_4758,N_4721);
nand U4854 (N_4854,N_4794,N_4703);
nand U4855 (N_4855,N_4768,N_4712);
or U4856 (N_4856,N_4771,N_4706);
or U4857 (N_4857,N_4725,N_4700);
nand U4858 (N_4858,N_4772,N_4746);
xnor U4859 (N_4859,N_4717,N_4749);
or U4860 (N_4860,N_4742,N_4757);
nand U4861 (N_4861,N_4721,N_4710);
and U4862 (N_4862,N_4767,N_4787);
nand U4863 (N_4863,N_4714,N_4710);
or U4864 (N_4864,N_4762,N_4708);
and U4865 (N_4865,N_4774,N_4787);
nor U4866 (N_4866,N_4759,N_4791);
or U4867 (N_4867,N_4715,N_4738);
or U4868 (N_4868,N_4704,N_4762);
nand U4869 (N_4869,N_4701,N_4717);
and U4870 (N_4870,N_4760,N_4756);
nand U4871 (N_4871,N_4757,N_4701);
and U4872 (N_4872,N_4787,N_4736);
or U4873 (N_4873,N_4747,N_4785);
and U4874 (N_4874,N_4702,N_4703);
nor U4875 (N_4875,N_4790,N_4797);
nand U4876 (N_4876,N_4730,N_4775);
and U4877 (N_4877,N_4754,N_4753);
nor U4878 (N_4878,N_4789,N_4795);
xor U4879 (N_4879,N_4718,N_4762);
nand U4880 (N_4880,N_4700,N_4783);
nor U4881 (N_4881,N_4782,N_4771);
nor U4882 (N_4882,N_4745,N_4748);
or U4883 (N_4883,N_4746,N_4794);
and U4884 (N_4884,N_4707,N_4760);
and U4885 (N_4885,N_4784,N_4720);
or U4886 (N_4886,N_4710,N_4769);
and U4887 (N_4887,N_4761,N_4788);
nand U4888 (N_4888,N_4723,N_4741);
nand U4889 (N_4889,N_4752,N_4713);
nor U4890 (N_4890,N_4797,N_4747);
nand U4891 (N_4891,N_4725,N_4704);
nand U4892 (N_4892,N_4704,N_4736);
or U4893 (N_4893,N_4781,N_4763);
nor U4894 (N_4894,N_4772,N_4752);
and U4895 (N_4895,N_4760,N_4776);
xnor U4896 (N_4896,N_4788,N_4747);
and U4897 (N_4897,N_4776,N_4783);
and U4898 (N_4898,N_4724,N_4797);
nor U4899 (N_4899,N_4754,N_4797);
or U4900 (N_4900,N_4804,N_4875);
nor U4901 (N_4901,N_4825,N_4861);
xor U4902 (N_4902,N_4808,N_4836);
xor U4903 (N_4903,N_4894,N_4864);
and U4904 (N_4904,N_4820,N_4822);
nor U4905 (N_4905,N_4815,N_4872);
xor U4906 (N_4906,N_4838,N_4890);
nand U4907 (N_4907,N_4889,N_4824);
nand U4908 (N_4908,N_4867,N_4848);
and U4909 (N_4909,N_4854,N_4865);
and U4910 (N_4910,N_4852,N_4829);
nand U4911 (N_4911,N_4814,N_4839);
xor U4912 (N_4912,N_4845,N_4897);
nor U4913 (N_4913,N_4802,N_4881);
or U4914 (N_4914,N_4862,N_4850);
nor U4915 (N_4915,N_4866,N_4880);
or U4916 (N_4916,N_4888,N_4874);
nor U4917 (N_4917,N_4813,N_4819);
xor U4918 (N_4918,N_4870,N_4809);
or U4919 (N_4919,N_4843,N_4857);
and U4920 (N_4920,N_4834,N_4841);
xnor U4921 (N_4921,N_4858,N_4878);
xnor U4922 (N_4922,N_4883,N_4810);
xor U4923 (N_4923,N_4859,N_4882);
or U4924 (N_4924,N_4831,N_4833);
and U4925 (N_4925,N_4860,N_4801);
xor U4926 (N_4926,N_4847,N_4828);
or U4927 (N_4927,N_4895,N_4812);
nand U4928 (N_4928,N_4869,N_4871);
nand U4929 (N_4929,N_4805,N_4899);
nand U4930 (N_4930,N_4877,N_4853);
or U4931 (N_4931,N_4816,N_4876);
and U4932 (N_4932,N_4846,N_4803);
or U4933 (N_4933,N_4806,N_4879);
nand U4934 (N_4934,N_4817,N_4885);
or U4935 (N_4935,N_4891,N_4818);
nand U4936 (N_4936,N_4855,N_4826);
or U4937 (N_4937,N_4842,N_4868);
xor U4938 (N_4938,N_4849,N_4873);
or U4939 (N_4939,N_4827,N_4896);
nor U4940 (N_4940,N_4884,N_4832);
nor U4941 (N_4941,N_4835,N_4807);
nor U4942 (N_4942,N_4830,N_4887);
nor U4943 (N_4943,N_4844,N_4821);
nor U4944 (N_4944,N_4823,N_4886);
nor U4945 (N_4945,N_4840,N_4898);
nor U4946 (N_4946,N_4811,N_4800);
or U4947 (N_4947,N_4851,N_4856);
and U4948 (N_4948,N_4863,N_4892);
xor U4949 (N_4949,N_4893,N_4837);
xor U4950 (N_4950,N_4807,N_4806);
xor U4951 (N_4951,N_4889,N_4880);
or U4952 (N_4952,N_4866,N_4862);
or U4953 (N_4953,N_4885,N_4816);
nand U4954 (N_4954,N_4839,N_4859);
nor U4955 (N_4955,N_4870,N_4833);
nor U4956 (N_4956,N_4898,N_4868);
xnor U4957 (N_4957,N_4842,N_4814);
nand U4958 (N_4958,N_4889,N_4877);
xor U4959 (N_4959,N_4889,N_4862);
xnor U4960 (N_4960,N_4865,N_4884);
nand U4961 (N_4961,N_4877,N_4881);
xnor U4962 (N_4962,N_4838,N_4892);
nand U4963 (N_4963,N_4849,N_4841);
xnor U4964 (N_4964,N_4841,N_4802);
xnor U4965 (N_4965,N_4846,N_4819);
xor U4966 (N_4966,N_4887,N_4820);
and U4967 (N_4967,N_4896,N_4881);
and U4968 (N_4968,N_4842,N_4816);
nor U4969 (N_4969,N_4838,N_4846);
nor U4970 (N_4970,N_4808,N_4819);
nor U4971 (N_4971,N_4895,N_4864);
or U4972 (N_4972,N_4836,N_4877);
nand U4973 (N_4973,N_4801,N_4811);
and U4974 (N_4974,N_4846,N_4868);
and U4975 (N_4975,N_4823,N_4879);
nand U4976 (N_4976,N_4822,N_4824);
nand U4977 (N_4977,N_4804,N_4813);
and U4978 (N_4978,N_4877,N_4826);
xor U4979 (N_4979,N_4818,N_4821);
nor U4980 (N_4980,N_4809,N_4812);
xor U4981 (N_4981,N_4852,N_4879);
or U4982 (N_4982,N_4825,N_4832);
and U4983 (N_4983,N_4877,N_4810);
or U4984 (N_4984,N_4851,N_4839);
nand U4985 (N_4985,N_4868,N_4814);
xor U4986 (N_4986,N_4843,N_4863);
or U4987 (N_4987,N_4828,N_4846);
xnor U4988 (N_4988,N_4875,N_4822);
nor U4989 (N_4989,N_4853,N_4814);
nor U4990 (N_4990,N_4847,N_4801);
and U4991 (N_4991,N_4864,N_4883);
or U4992 (N_4992,N_4810,N_4856);
and U4993 (N_4993,N_4899,N_4806);
and U4994 (N_4994,N_4819,N_4852);
xor U4995 (N_4995,N_4880,N_4839);
xnor U4996 (N_4996,N_4816,N_4846);
nor U4997 (N_4997,N_4872,N_4857);
xnor U4998 (N_4998,N_4839,N_4874);
and U4999 (N_4999,N_4876,N_4823);
nand U5000 (N_5000,N_4934,N_4939);
xnor U5001 (N_5001,N_4943,N_4935);
xor U5002 (N_5002,N_4949,N_4948);
and U5003 (N_5003,N_4905,N_4912);
nor U5004 (N_5004,N_4911,N_4956);
nor U5005 (N_5005,N_4980,N_4920);
nor U5006 (N_5006,N_4903,N_4906);
and U5007 (N_5007,N_4910,N_4963);
xnor U5008 (N_5008,N_4914,N_4946);
nand U5009 (N_5009,N_4974,N_4998);
xor U5010 (N_5010,N_4926,N_4960);
xor U5011 (N_5011,N_4990,N_4908);
xor U5012 (N_5012,N_4950,N_4944);
nor U5013 (N_5013,N_4957,N_4987);
and U5014 (N_5014,N_4937,N_4927);
and U5015 (N_5015,N_4999,N_4904);
nor U5016 (N_5016,N_4989,N_4933);
nand U5017 (N_5017,N_4991,N_4975);
or U5018 (N_5018,N_4977,N_4971);
xnor U5019 (N_5019,N_4947,N_4996);
and U5020 (N_5020,N_4900,N_4917);
and U5021 (N_5021,N_4907,N_4968);
nand U5022 (N_5022,N_4924,N_4966);
nor U5023 (N_5023,N_4992,N_4985);
and U5024 (N_5024,N_4915,N_4921);
nand U5025 (N_5025,N_4954,N_4988);
xnor U5026 (N_5026,N_4955,N_4922);
or U5027 (N_5027,N_4961,N_4913);
or U5028 (N_5028,N_4994,N_4918);
xnor U5029 (N_5029,N_4958,N_4967);
nand U5030 (N_5030,N_4965,N_4945);
or U5031 (N_5031,N_4936,N_4938);
and U5032 (N_5032,N_4951,N_4932);
or U5033 (N_5033,N_4942,N_4984);
xnor U5034 (N_5034,N_4981,N_4972);
nor U5035 (N_5035,N_4976,N_4962);
nand U5036 (N_5036,N_4982,N_4986);
and U5037 (N_5037,N_4929,N_4941);
nand U5038 (N_5038,N_4931,N_4953);
nor U5039 (N_5039,N_4959,N_4993);
nor U5040 (N_5040,N_4952,N_4983);
and U5041 (N_5041,N_4979,N_4928);
or U5042 (N_5042,N_4919,N_4978);
xor U5043 (N_5043,N_4973,N_4909);
and U5044 (N_5044,N_4940,N_4969);
and U5045 (N_5045,N_4901,N_4902);
nand U5046 (N_5046,N_4995,N_4964);
and U5047 (N_5047,N_4930,N_4997);
nor U5048 (N_5048,N_4923,N_4925);
xnor U5049 (N_5049,N_4916,N_4970);
nor U5050 (N_5050,N_4975,N_4998);
or U5051 (N_5051,N_4920,N_4911);
xnor U5052 (N_5052,N_4942,N_4937);
or U5053 (N_5053,N_4944,N_4968);
xor U5054 (N_5054,N_4901,N_4963);
and U5055 (N_5055,N_4952,N_4988);
xnor U5056 (N_5056,N_4985,N_4923);
and U5057 (N_5057,N_4970,N_4965);
or U5058 (N_5058,N_4967,N_4993);
nand U5059 (N_5059,N_4985,N_4940);
nand U5060 (N_5060,N_4905,N_4973);
nor U5061 (N_5061,N_4995,N_4934);
or U5062 (N_5062,N_4990,N_4911);
xnor U5063 (N_5063,N_4904,N_4901);
and U5064 (N_5064,N_4916,N_4919);
or U5065 (N_5065,N_4986,N_4950);
xor U5066 (N_5066,N_4903,N_4930);
or U5067 (N_5067,N_4995,N_4924);
nor U5068 (N_5068,N_4977,N_4954);
and U5069 (N_5069,N_4919,N_4963);
and U5070 (N_5070,N_4983,N_4979);
nand U5071 (N_5071,N_4965,N_4923);
and U5072 (N_5072,N_4990,N_4945);
nor U5073 (N_5073,N_4987,N_4901);
xnor U5074 (N_5074,N_4983,N_4919);
nand U5075 (N_5075,N_4927,N_4986);
nor U5076 (N_5076,N_4965,N_4946);
nor U5077 (N_5077,N_4916,N_4978);
or U5078 (N_5078,N_4948,N_4976);
nand U5079 (N_5079,N_4943,N_4969);
and U5080 (N_5080,N_4912,N_4906);
xor U5081 (N_5081,N_4933,N_4927);
xor U5082 (N_5082,N_4958,N_4971);
nor U5083 (N_5083,N_4932,N_4994);
or U5084 (N_5084,N_4997,N_4950);
xnor U5085 (N_5085,N_4980,N_4953);
nor U5086 (N_5086,N_4993,N_4994);
xnor U5087 (N_5087,N_4967,N_4982);
xor U5088 (N_5088,N_4941,N_4924);
nor U5089 (N_5089,N_4953,N_4934);
nor U5090 (N_5090,N_4977,N_4970);
nand U5091 (N_5091,N_4943,N_4923);
or U5092 (N_5092,N_4910,N_4927);
nor U5093 (N_5093,N_4959,N_4927);
or U5094 (N_5094,N_4996,N_4934);
nor U5095 (N_5095,N_4976,N_4938);
nor U5096 (N_5096,N_4926,N_4918);
xnor U5097 (N_5097,N_4949,N_4939);
nor U5098 (N_5098,N_4935,N_4968);
xor U5099 (N_5099,N_4930,N_4965);
nand U5100 (N_5100,N_5025,N_5009);
and U5101 (N_5101,N_5027,N_5072);
and U5102 (N_5102,N_5041,N_5081);
nor U5103 (N_5103,N_5088,N_5005);
nor U5104 (N_5104,N_5099,N_5051);
and U5105 (N_5105,N_5060,N_5002);
or U5106 (N_5106,N_5033,N_5008);
xnor U5107 (N_5107,N_5054,N_5004);
and U5108 (N_5108,N_5074,N_5065);
nor U5109 (N_5109,N_5073,N_5012);
nand U5110 (N_5110,N_5010,N_5076);
and U5111 (N_5111,N_5092,N_5063);
xnor U5112 (N_5112,N_5082,N_5069);
xnor U5113 (N_5113,N_5038,N_5006);
nor U5114 (N_5114,N_5048,N_5044);
nor U5115 (N_5115,N_5011,N_5037);
nor U5116 (N_5116,N_5079,N_5095);
nor U5117 (N_5117,N_5078,N_5058);
nand U5118 (N_5118,N_5014,N_5080);
xnor U5119 (N_5119,N_5096,N_5042);
xnor U5120 (N_5120,N_5097,N_5035);
nand U5121 (N_5121,N_5003,N_5064);
and U5122 (N_5122,N_5046,N_5031);
or U5123 (N_5123,N_5085,N_5024);
xnor U5124 (N_5124,N_5084,N_5043);
nor U5125 (N_5125,N_5018,N_5053);
nand U5126 (N_5126,N_5070,N_5050);
nand U5127 (N_5127,N_5021,N_5062);
nor U5128 (N_5128,N_5023,N_5040);
or U5129 (N_5129,N_5093,N_5047);
or U5130 (N_5130,N_5017,N_5056);
nor U5131 (N_5131,N_5020,N_5032);
nor U5132 (N_5132,N_5015,N_5086);
and U5133 (N_5133,N_5055,N_5090);
nand U5134 (N_5134,N_5001,N_5052);
xnor U5135 (N_5135,N_5026,N_5067);
or U5136 (N_5136,N_5059,N_5016);
and U5137 (N_5137,N_5030,N_5089);
and U5138 (N_5138,N_5083,N_5077);
or U5139 (N_5139,N_5022,N_5098);
xor U5140 (N_5140,N_5071,N_5075);
and U5141 (N_5141,N_5094,N_5029);
or U5142 (N_5142,N_5034,N_5066);
nor U5143 (N_5143,N_5061,N_5045);
nor U5144 (N_5144,N_5028,N_5039);
xnor U5145 (N_5145,N_5049,N_5087);
xor U5146 (N_5146,N_5007,N_5068);
nor U5147 (N_5147,N_5036,N_5019);
and U5148 (N_5148,N_5091,N_5057);
nor U5149 (N_5149,N_5000,N_5013);
and U5150 (N_5150,N_5035,N_5074);
and U5151 (N_5151,N_5004,N_5072);
or U5152 (N_5152,N_5055,N_5003);
xor U5153 (N_5153,N_5026,N_5084);
nand U5154 (N_5154,N_5052,N_5051);
nand U5155 (N_5155,N_5067,N_5077);
nor U5156 (N_5156,N_5039,N_5016);
or U5157 (N_5157,N_5036,N_5041);
xor U5158 (N_5158,N_5047,N_5037);
xnor U5159 (N_5159,N_5006,N_5013);
nor U5160 (N_5160,N_5029,N_5025);
nand U5161 (N_5161,N_5056,N_5088);
nor U5162 (N_5162,N_5069,N_5068);
nor U5163 (N_5163,N_5052,N_5013);
nor U5164 (N_5164,N_5042,N_5011);
xnor U5165 (N_5165,N_5079,N_5071);
nand U5166 (N_5166,N_5081,N_5001);
or U5167 (N_5167,N_5007,N_5077);
or U5168 (N_5168,N_5091,N_5042);
nor U5169 (N_5169,N_5050,N_5097);
xnor U5170 (N_5170,N_5091,N_5052);
or U5171 (N_5171,N_5038,N_5031);
or U5172 (N_5172,N_5057,N_5093);
or U5173 (N_5173,N_5089,N_5042);
xnor U5174 (N_5174,N_5011,N_5084);
nand U5175 (N_5175,N_5071,N_5086);
nor U5176 (N_5176,N_5054,N_5019);
or U5177 (N_5177,N_5031,N_5012);
and U5178 (N_5178,N_5060,N_5075);
and U5179 (N_5179,N_5082,N_5025);
nand U5180 (N_5180,N_5052,N_5034);
xnor U5181 (N_5181,N_5007,N_5096);
nand U5182 (N_5182,N_5000,N_5055);
xnor U5183 (N_5183,N_5087,N_5029);
or U5184 (N_5184,N_5056,N_5078);
or U5185 (N_5185,N_5032,N_5030);
xor U5186 (N_5186,N_5041,N_5015);
and U5187 (N_5187,N_5052,N_5039);
or U5188 (N_5188,N_5005,N_5009);
nor U5189 (N_5189,N_5010,N_5024);
and U5190 (N_5190,N_5055,N_5066);
nand U5191 (N_5191,N_5076,N_5037);
or U5192 (N_5192,N_5080,N_5084);
nand U5193 (N_5193,N_5051,N_5000);
or U5194 (N_5194,N_5036,N_5085);
or U5195 (N_5195,N_5017,N_5000);
and U5196 (N_5196,N_5043,N_5096);
or U5197 (N_5197,N_5029,N_5044);
xnor U5198 (N_5198,N_5071,N_5055);
nor U5199 (N_5199,N_5067,N_5013);
and U5200 (N_5200,N_5164,N_5146);
xnor U5201 (N_5201,N_5111,N_5186);
nor U5202 (N_5202,N_5134,N_5185);
nand U5203 (N_5203,N_5149,N_5197);
nor U5204 (N_5204,N_5198,N_5177);
xor U5205 (N_5205,N_5113,N_5166);
xnor U5206 (N_5206,N_5153,N_5138);
xor U5207 (N_5207,N_5139,N_5136);
nor U5208 (N_5208,N_5174,N_5100);
and U5209 (N_5209,N_5182,N_5123);
and U5210 (N_5210,N_5176,N_5148);
and U5211 (N_5211,N_5161,N_5163);
and U5212 (N_5212,N_5151,N_5160);
nand U5213 (N_5213,N_5143,N_5105);
xor U5214 (N_5214,N_5135,N_5114);
or U5215 (N_5215,N_5171,N_5156);
or U5216 (N_5216,N_5118,N_5124);
xnor U5217 (N_5217,N_5152,N_5121);
and U5218 (N_5218,N_5181,N_5120);
and U5219 (N_5219,N_5108,N_5142);
xnor U5220 (N_5220,N_5184,N_5119);
nand U5221 (N_5221,N_5173,N_5127);
and U5222 (N_5222,N_5147,N_5116);
and U5223 (N_5223,N_5101,N_5175);
or U5224 (N_5224,N_5183,N_5188);
xor U5225 (N_5225,N_5126,N_5189);
nand U5226 (N_5226,N_5196,N_5187);
nor U5227 (N_5227,N_5129,N_5180);
nor U5228 (N_5228,N_5132,N_5190);
and U5229 (N_5229,N_5170,N_5150);
nand U5230 (N_5230,N_5192,N_5194);
xnor U5231 (N_5231,N_5168,N_5131);
and U5232 (N_5232,N_5140,N_5154);
and U5233 (N_5233,N_5158,N_5167);
xor U5234 (N_5234,N_5178,N_5199);
nand U5235 (N_5235,N_5162,N_5155);
and U5236 (N_5236,N_5195,N_5159);
and U5237 (N_5237,N_5193,N_5117);
xnor U5238 (N_5238,N_5133,N_5107);
xnor U5239 (N_5239,N_5104,N_5102);
nand U5240 (N_5240,N_5179,N_5106);
or U5241 (N_5241,N_5144,N_5110);
and U5242 (N_5242,N_5112,N_5122);
nand U5243 (N_5243,N_5157,N_5137);
and U5244 (N_5244,N_5172,N_5145);
nand U5245 (N_5245,N_5141,N_5165);
nand U5246 (N_5246,N_5191,N_5125);
xnor U5247 (N_5247,N_5128,N_5130);
nand U5248 (N_5248,N_5109,N_5115);
or U5249 (N_5249,N_5103,N_5169);
and U5250 (N_5250,N_5135,N_5149);
nand U5251 (N_5251,N_5156,N_5177);
nand U5252 (N_5252,N_5147,N_5171);
nand U5253 (N_5253,N_5139,N_5131);
or U5254 (N_5254,N_5189,N_5190);
or U5255 (N_5255,N_5122,N_5115);
or U5256 (N_5256,N_5158,N_5178);
nand U5257 (N_5257,N_5107,N_5126);
or U5258 (N_5258,N_5154,N_5137);
nand U5259 (N_5259,N_5171,N_5173);
xor U5260 (N_5260,N_5104,N_5101);
nand U5261 (N_5261,N_5163,N_5109);
and U5262 (N_5262,N_5120,N_5191);
xor U5263 (N_5263,N_5110,N_5124);
nand U5264 (N_5264,N_5129,N_5154);
xnor U5265 (N_5265,N_5111,N_5136);
xnor U5266 (N_5266,N_5142,N_5159);
and U5267 (N_5267,N_5131,N_5104);
or U5268 (N_5268,N_5120,N_5152);
nand U5269 (N_5269,N_5139,N_5168);
xnor U5270 (N_5270,N_5145,N_5173);
or U5271 (N_5271,N_5177,N_5140);
nor U5272 (N_5272,N_5157,N_5135);
nand U5273 (N_5273,N_5197,N_5110);
or U5274 (N_5274,N_5180,N_5137);
or U5275 (N_5275,N_5163,N_5113);
nor U5276 (N_5276,N_5199,N_5185);
and U5277 (N_5277,N_5131,N_5172);
and U5278 (N_5278,N_5198,N_5133);
xor U5279 (N_5279,N_5185,N_5113);
or U5280 (N_5280,N_5171,N_5131);
xnor U5281 (N_5281,N_5131,N_5119);
nand U5282 (N_5282,N_5118,N_5190);
and U5283 (N_5283,N_5143,N_5171);
and U5284 (N_5284,N_5135,N_5165);
and U5285 (N_5285,N_5122,N_5149);
xnor U5286 (N_5286,N_5147,N_5103);
nand U5287 (N_5287,N_5100,N_5125);
nor U5288 (N_5288,N_5179,N_5133);
and U5289 (N_5289,N_5140,N_5190);
nand U5290 (N_5290,N_5130,N_5195);
nand U5291 (N_5291,N_5198,N_5151);
nor U5292 (N_5292,N_5199,N_5120);
nand U5293 (N_5293,N_5176,N_5113);
xor U5294 (N_5294,N_5192,N_5136);
nor U5295 (N_5295,N_5168,N_5123);
nand U5296 (N_5296,N_5159,N_5149);
xor U5297 (N_5297,N_5152,N_5189);
nand U5298 (N_5298,N_5143,N_5189);
nor U5299 (N_5299,N_5194,N_5179);
xnor U5300 (N_5300,N_5286,N_5289);
nor U5301 (N_5301,N_5247,N_5216);
and U5302 (N_5302,N_5274,N_5242);
nand U5303 (N_5303,N_5254,N_5280);
and U5304 (N_5304,N_5210,N_5201);
nand U5305 (N_5305,N_5208,N_5257);
xnor U5306 (N_5306,N_5285,N_5209);
nand U5307 (N_5307,N_5200,N_5211);
xnor U5308 (N_5308,N_5298,N_5267);
nor U5309 (N_5309,N_5225,N_5299);
xnor U5310 (N_5310,N_5262,N_5213);
or U5311 (N_5311,N_5268,N_5217);
nand U5312 (N_5312,N_5252,N_5249);
and U5313 (N_5313,N_5261,N_5233);
nand U5314 (N_5314,N_5236,N_5256);
or U5315 (N_5315,N_5296,N_5205);
or U5316 (N_5316,N_5229,N_5259);
or U5317 (N_5317,N_5230,N_5204);
nor U5318 (N_5318,N_5292,N_5237);
or U5319 (N_5319,N_5269,N_5207);
or U5320 (N_5320,N_5297,N_5253);
nor U5321 (N_5321,N_5287,N_5221);
nor U5322 (N_5322,N_5234,N_5270);
or U5323 (N_5323,N_5284,N_5240);
nand U5324 (N_5324,N_5224,N_5202);
or U5325 (N_5325,N_5222,N_5203);
and U5326 (N_5326,N_5251,N_5232);
nor U5327 (N_5327,N_5250,N_5214);
nor U5328 (N_5328,N_5212,N_5263);
nor U5329 (N_5329,N_5265,N_5243);
xor U5330 (N_5330,N_5294,N_5228);
nand U5331 (N_5331,N_5226,N_5276);
xor U5332 (N_5332,N_5206,N_5278);
and U5333 (N_5333,N_5264,N_5218);
nand U5334 (N_5334,N_5219,N_5275);
xor U5335 (N_5335,N_5231,N_5238);
or U5336 (N_5336,N_5245,N_5248);
xor U5337 (N_5337,N_5244,N_5246);
nand U5338 (N_5338,N_5239,N_5227);
and U5339 (N_5339,N_5273,N_5241);
xnor U5340 (N_5340,N_5282,N_5291);
xnor U5341 (N_5341,N_5293,N_5255);
xnor U5342 (N_5342,N_5277,N_5272);
xor U5343 (N_5343,N_5288,N_5266);
or U5344 (N_5344,N_5215,N_5271);
nand U5345 (N_5345,N_5220,N_5295);
nor U5346 (N_5346,N_5258,N_5281);
xnor U5347 (N_5347,N_5283,N_5290);
xor U5348 (N_5348,N_5223,N_5260);
nand U5349 (N_5349,N_5279,N_5235);
nand U5350 (N_5350,N_5229,N_5292);
nor U5351 (N_5351,N_5266,N_5291);
nand U5352 (N_5352,N_5232,N_5278);
nand U5353 (N_5353,N_5201,N_5231);
or U5354 (N_5354,N_5257,N_5247);
nand U5355 (N_5355,N_5247,N_5209);
or U5356 (N_5356,N_5263,N_5258);
xor U5357 (N_5357,N_5297,N_5205);
or U5358 (N_5358,N_5271,N_5211);
and U5359 (N_5359,N_5298,N_5284);
or U5360 (N_5360,N_5272,N_5240);
xor U5361 (N_5361,N_5212,N_5230);
nor U5362 (N_5362,N_5220,N_5250);
and U5363 (N_5363,N_5270,N_5238);
nand U5364 (N_5364,N_5222,N_5259);
nand U5365 (N_5365,N_5285,N_5216);
nand U5366 (N_5366,N_5251,N_5262);
and U5367 (N_5367,N_5240,N_5215);
and U5368 (N_5368,N_5239,N_5263);
nor U5369 (N_5369,N_5250,N_5272);
and U5370 (N_5370,N_5260,N_5268);
and U5371 (N_5371,N_5249,N_5282);
xnor U5372 (N_5372,N_5229,N_5220);
or U5373 (N_5373,N_5271,N_5209);
and U5374 (N_5374,N_5213,N_5266);
or U5375 (N_5375,N_5262,N_5272);
nor U5376 (N_5376,N_5259,N_5212);
xor U5377 (N_5377,N_5294,N_5263);
and U5378 (N_5378,N_5205,N_5238);
xor U5379 (N_5379,N_5231,N_5240);
or U5380 (N_5380,N_5294,N_5281);
nand U5381 (N_5381,N_5247,N_5204);
xor U5382 (N_5382,N_5288,N_5295);
xnor U5383 (N_5383,N_5225,N_5209);
and U5384 (N_5384,N_5284,N_5243);
nor U5385 (N_5385,N_5242,N_5215);
or U5386 (N_5386,N_5221,N_5268);
and U5387 (N_5387,N_5249,N_5215);
and U5388 (N_5388,N_5279,N_5242);
and U5389 (N_5389,N_5281,N_5296);
or U5390 (N_5390,N_5208,N_5241);
or U5391 (N_5391,N_5210,N_5262);
nor U5392 (N_5392,N_5295,N_5254);
or U5393 (N_5393,N_5219,N_5201);
or U5394 (N_5394,N_5258,N_5231);
xor U5395 (N_5395,N_5299,N_5221);
or U5396 (N_5396,N_5267,N_5206);
xnor U5397 (N_5397,N_5248,N_5278);
nor U5398 (N_5398,N_5250,N_5283);
nor U5399 (N_5399,N_5233,N_5296);
nand U5400 (N_5400,N_5358,N_5339);
or U5401 (N_5401,N_5343,N_5317);
and U5402 (N_5402,N_5395,N_5330);
and U5403 (N_5403,N_5349,N_5388);
nor U5404 (N_5404,N_5353,N_5377);
or U5405 (N_5405,N_5380,N_5303);
and U5406 (N_5406,N_5382,N_5338);
xnor U5407 (N_5407,N_5348,N_5311);
and U5408 (N_5408,N_5399,N_5325);
xnor U5409 (N_5409,N_5393,N_5373);
xor U5410 (N_5410,N_5376,N_5385);
and U5411 (N_5411,N_5334,N_5352);
nor U5412 (N_5412,N_5367,N_5346);
nand U5413 (N_5413,N_5300,N_5362);
and U5414 (N_5414,N_5350,N_5328);
or U5415 (N_5415,N_5342,N_5360);
and U5416 (N_5416,N_5397,N_5312);
nor U5417 (N_5417,N_5324,N_5331);
nand U5418 (N_5418,N_5351,N_5394);
xnor U5419 (N_5419,N_5337,N_5369);
xnor U5420 (N_5420,N_5354,N_5384);
and U5421 (N_5421,N_5316,N_5313);
nor U5422 (N_5422,N_5381,N_5301);
nor U5423 (N_5423,N_5389,N_5310);
xor U5424 (N_5424,N_5309,N_5319);
nand U5425 (N_5425,N_5374,N_5340);
nand U5426 (N_5426,N_5327,N_5356);
or U5427 (N_5427,N_5307,N_5305);
or U5428 (N_5428,N_5357,N_5322);
and U5429 (N_5429,N_5370,N_5306);
xnor U5430 (N_5430,N_5323,N_5363);
or U5431 (N_5431,N_5341,N_5308);
or U5432 (N_5432,N_5372,N_5335);
and U5433 (N_5433,N_5318,N_5396);
xor U5434 (N_5434,N_5387,N_5320);
nor U5435 (N_5435,N_5332,N_5344);
nand U5436 (N_5436,N_5386,N_5336);
xnor U5437 (N_5437,N_5361,N_5355);
nand U5438 (N_5438,N_5333,N_5345);
or U5439 (N_5439,N_5368,N_5371);
nand U5440 (N_5440,N_5375,N_5364);
and U5441 (N_5441,N_5365,N_5329);
xnor U5442 (N_5442,N_5302,N_5304);
nor U5443 (N_5443,N_5392,N_5321);
nor U5444 (N_5444,N_5314,N_5359);
nand U5445 (N_5445,N_5315,N_5378);
or U5446 (N_5446,N_5390,N_5398);
nand U5447 (N_5447,N_5379,N_5326);
xnor U5448 (N_5448,N_5391,N_5347);
or U5449 (N_5449,N_5383,N_5366);
or U5450 (N_5450,N_5379,N_5331);
xor U5451 (N_5451,N_5304,N_5369);
xor U5452 (N_5452,N_5339,N_5343);
nand U5453 (N_5453,N_5356,N_5368);
xnor U5454 (N_5454,N_5388,N_5318);
or U5455 (N_5455,N_5321,N_5339);
and U5456 (N_5456,N_5366,N_5384);
nand U5457 (N_5457,N_5322,N_5324);
xor U5458 (N_5458,N_5315,N_5341);
nand U5459 (N_5459,N_5310,N_5363);
nor U5460 (N_5460,N_5307,N_5321);
or U5461 (N_5461,N_5391,N_5342);
or U5462 (N_5462,N_5301,N_5388);
and U5463 (N_5463,N_5308,N_5302);
or U5464 (N_5464,N_5381,N_5362);
nand U5465 (N_5465,N_5300,N_5357);
nor U5466 (N_5466,N_5325,N_5364);
or U5467 (N_5467,N_5392,N_5329);
or U5468 (N_5468,N_5377,N_5321);
and U5469 (N_5469,N_5300,N_5342);
xor U5470 (N_5470,N_5325,N_5358);
and U5471 (N_5471,N_5383,N_5367);
nor U5472 (N_5472,N_5316,N_5308);
or U5473 (N_5473,N_5305,N_5369);
xnor U5474 (N_5474,N_5323,N_5345);
or U5475 (N_5475,N_5344,N_5343);
xnor U5476 (N_5476,N_5344,N_5388);
xor U5477 (N_5477,N_5335,N_5382);
nor U5478 (N_5478,N_5339,N_5336);
nand U5479 (N_5479,N_5394,N_5383);
and U5480 (N_5480,N_5324,N_5388);
nand U5481 (N_5481,N_5319,N_5312);
and U5482 (N_5482,N_5361,N_5376);
or U5483 (N_5483,N_5359,N_5337);
and U5484 (N_5484,N_5372,N_5322);
xor U5485 (N_5485,N_5397,N_5319);
and U5486 (N_5486,N_5396,N_5334);
nor U5487 (N_5487,N_5329,N_5374);
or U5488 (N_5488,N_5359,N_5387);
nor U5489 (N_5489,N_5353,N_5325);
nor U5490 (N_5490,N_5347,N_5303);
xor U5491 (N_5491,N_5305,N_5387);
and U5492 (N_5492,N_5318,N_5339);
or U5493 (N_5493,N_5377,N_5329);
xor U5494 (N_5494,N_5389,N_5386);
or U5495 (N_5495,N_5379,N_5378);
or U5496 (N_5496,N_5395,N_5343);
nand U5497 (N_5497,N_5329,N_5313);
nor U5498 (N_5498,N_5317,N_5385);
xor U5499 (N_5499,N_5389,N_5381);
xor U5500 (N_5500,N_5472,N_5414);
or U5501 (N_5501,N_5410,N_5474);
or U5502 (N_5502,N_5425,N_5457);
xnor U5503 (N_5503,N_5421,N_5468);
or U5504 (N_5504,N_5405,N_5411);
and U5505 (N_5505,N_5456,N_5452);
nor U5506 (N_5506,N_5431,N_5418);
nand U5507 (N_5507,N_5404,N_5491);
nor U5508 (N_5508,N_5471,N_5429);
xor U5509 (N_5509,N_5486,N_5437);
and U5510 (N_5510,N_5493,N_5482);
or U5511 (N_5511,N_5440,N_5408);
or U5512 (N_5512,N_5454,N_5481);
xor U5513 (N_5513,N_5444,N_5467);
and U5514 (N_5514,N_5446,N_5455);
or U5515 (N_5515,N_5434,N_5443);
nor U5516 (N_5516,N_5498,N_5415);
xnor U5517 (N_5517,N_5439,N_5476);
nor U5518 (N_5518,N_5413,N_5499);
and U5519 (N_5519,N_5460,N_5445);
xnor U5520 (N_5520,N_5447,N_5419);
xnor U5521 (N_5521,N_5403,N_5424);
xor U5522 (N_5522,N_5409,N_5464);
nor U5523 (N_5523,N_5478,N_5432);
or U5524 (N_5524,N_5492,N_5459);
and U5525 (N_5525,N_5490,N_5469);
or U5526 (N_5526,N_5402,N_5433);
xnor U5527 (N_5527,N_5400,N_5453);
or U5528 (N_5528,N_5401,N_5477);
xnor U5529 (N_5529,N_5487,N_5412);
nand U5530 (N_5530,N_5416,N_5458);
nor U5531 (N_5531,N_5427,N_5479);
or U5532 (N_5532,N_5450,N_5485);
xnor U5533 (N_5533,N_5494,N_5497);
or U5534 (N_5534,N_5480,N_5441);
xnor U5535 (N_5535,N_5488,N_5430);
and U5536 (N_5536,N_5470,N_5407);
xor U5537 (N_5537,N_5420,N_5462);
or U5538 (N_5538,N_5423,N_5484);
or U5539 (N_5539,N_5448,N_5466);
or U5540 (N_5540,N_5463,N_5489);
xnor U5541 (N_5541,N_5428,N_5442);
nor U5542 (N_5542,N_5406,N_5435);
and U5543 (N_5543,N_5496,N_5483);
nand U5544 (N_5544,N_5449,N_5451);
nand U5545 (N_5545,N_5473,N_5436);
nand U5546 (N_5546,N_5495,N_5461);
nor U5547 (N_5547,N_5422,N_5426);
or U5548 (N_5548,N_5438,N_5417);
and U5549 (N_5549,N_5475,N_5465);
xnor U5550 (N_5550,N_5418,N_5458);
or U5551 (N_5551,N_5416,N_5441);
xnor U5552 (N_5552,N_5403,N_5452);
or U5553 (N_5553,N_5450,N_5498);
and U5554 (N_5554,N_5416,N_5478);
and U5555 (N_5555,N_5456,N_5464);
or U5556 (N_5556,N_5498,N_5490);
nand U5557 (N_5557,N_5411,N_5420);
or U5558 (N_5558,N_5416,N_5453);
nor U5559 (N_5559,N_5464,N_5433);
xor U5560 (N_5560,N_5488,N_5489);
xor U5561 (N_5561,N_5477,N_5440);
nand U5562 (N_5562,N_5425,N_5478);
nor U5563 (N_5563,N_5401,N_5410);
or U5564 (N_5564,N_5463,N_5412);
xor U5565 (N_5565,N_5402,N_5483);
or U5566 (N_5566,N_5462,N_5472);
nand U5567 (N_5567,N_5426,N_5464);
nor U5568 (N_5568,N_5445,N_5484);
or U5569 (N_5569,N_5416,N_5431);
and U5570 (N_5570,N_5487,N_5435);
xor U5571 (N_5571,N_5487,N_5429);
nor U5572 (N_5572,N_5458,N_5415);
nand U5573 (N_5573,N_5400,N_5481);
nand U5574 (N_5574,N_5409,N_5486);
xnor U5575 (N_5575,N_5483,N_5421);
xnor U5576 (N_5576,N_5465,N_5479);
xnor U5577 (N_5577,N_5495,N_5497);
nand U5578 (N_5578,N_5494,N_5420);
nor U5579 (N_5579,N_5424,N_5400);
xor U5580 (N_5580,N_5440,N_5426);
or U5581 (N_5581,N_5469,N_5496);
and U5582 (N_5582,N_5413,N_5419);
nor U5583 (N_5583,N_5464,N_5420);
and U5584 (N_5584,N_5444,N_5434);
nor U5585 (N_5585,N_5406,N_5484);
and U5586 (N_5586,N_5449,N_5426);
or U5587 (N_5587,N_5476,N_5436);
nor U5588 (N_5588,N_5431,N_5486);
and U5589 (N_5589,N_5410,N_5430);
xor U5590 (N_5590,N_5480,N_5451);
or U5591 (N_5591,N_5432,N_5468);
and U5592 (N_5592,N_5426,N_5494);
or U5593 (N_5593,N_5463,N_5453);
nand U5594 (N_5594,N_5437,N_5489);
nand U5595 (N_5595,N_5435,N_5456);
or U5596 (N_5596,N_5464,N_5488);
nand U5597 (N_5597,N_5485,N_5497);
xnor U5598 (N_5598,N_5403,N_5425);
xor U5599 (N_5599,N_5450,N_5484);
nand U5600 (N_5600,N_5545,N_5552);
nor U5601 (N_5601,N_5571,N_5588);
xor U5602 (N_5602,N_5528,N_5553);
nand U5603 (N_5603,N_5590,N_5544);
nand U5604 (N_5604,N_5512,N_5515);
nor U5605 (N_5605,N_5579,N_5573);
nand U5606 (N_5606,N_5551,N_5570);
and U5607 (N_5607,N_5586,N_5568);
nor U5608 (N_5608,N_5538,N_5557);
xnor U5609 (N_5609,N_5530,N_5597);
or U5610 (N_5610,N_5589,N_5523);
nor U5611 (N_5611,N_5527,N_5549);
nor U5612 (N_5612,N_5591,N_5598);
nand U5613 (N_5613,N_5563,N_5599);
nand U5614 (N_5614,N_5558,N_5520);
or U5615 (N_5615,N_5518,N_5509);
and U5616 (N_5616,N_5565,N_5540);
xnor U5617 (N_5617,N_5572,N_5560);
xnor U5618 (N_5618,N_5500,N_5535);
xor U5619 (N_5619,N_5542,N_5504);
xor U5620 (N_5620,N_5584,N_5546);
nand U5621 (N_5621,N_5577,N_5519);
xor U5622 (N_5622,N_5511,N_5576);
nand U5623 (N_5623,N_5593,N_5548);
or U5624 (N_5624,N_5524,N_5525);
xnor U5625 (N_5625,N_5567,N_5534);
xor U5626 (N_5626,N_5587,N_5501);
nand U5627 (N_5627,N_5505,N_5516);
or U5628 (N_5628,N_5582,N_5539);
nand U5629 (N_5629,N_5543,N_5594);
nor U5630 (N_5630,N_5575,N_5537);
nor U5631 (N_5631,N_5556,N_5502);
nor U5632 (N_5632,N_5580,N_5529);
xnor U5633 (N_5633,N_5532,N_5536);
nand U5634 (N_5634,N_5569,N_5513);
nand U5635 (N_5635,N_5581,N_5562);
or U5636 (N_5636,N_5506,N_5510);
nand U5637 (N_5637,N_5585,N_5514);
xnor U5638 (N_5638,N_5526,N_5595);
nand U5639 (N_5639,N_5566,N_5533);
and U5640 (N_5640,N_5521,N_5554);
nor U5641 (N_5641,N_5547,N_5596);
and U5642 (N_5642,N_5503,N_5574);
or U5643 (N_5643,N_5583,N_5508);
xor U5644 (N_5644,N_5559,N_5541);
nor U5645 (N_5645,N_5592,N_5561);
xnor U5646 (N_5646,N_5555,N_5578);
and U5647 (N_5647,N_5550,N_5522);
or U5648 (N_5648,N_5517,N_5531);
xnor U5649 (N_5649,N_5507,N_5564);
nand U5650 (N_5650,N_5589,N_5501);
nand U5651 (N_5651,N_5518,N_5559);
or U5652 (N_5652,N_5513,N_5558);
and U5653 (N_5653,N_5504,N_5522);
nor U5654 (N_5654,N_5526,N_5533);
or U5655 (N_5655,N_5543,N_5500);
nor U5656 (N_5656,N_5513,N_5571);
nand U5657 (N_5657,N_5529,N_5574);
or U5658 (N_5658,N_5540,N_5561);
and U5659 (N_5659,N_5557,N_5545);
and U5660 (N_5660,N_5583,N_5594);
nor U5661 (N_5661,N_5506,N_5597);
or U5662 (N_5662,N_5571,N_5582);
or U5663 (N_5663,N_5552,N_5554);
nand U5664 (N_5664,N_5539,N_5553);
and U5665 (N_5665,N_5556,N_5529);
or U5666 (N_5666,N_5524,N_5548);
xnor U5667 (N_5667,N_5575,N_5518);
or U5668 (N_5668,N_5586,N_5588);
xnor U5669 (N_5669,N_5564,N_5588);
or U5670 (N_5670,N_5570,N_5542);
and U5671 (N_5671,N_5597,N_5525);
nor U5672 (N_5672,N_5566,N_5553);
xnor U5673 (N_5673,N_5517,N_5528);
nand U5674 (N_5674,N_5546,N_5551);
nand U5675 (N_5675,N_5525,N_5526);
or U5676 (N_5676,N_5509,N_5557);
or U5677 (N_5677,N_5513,N_5548);
nor U5678 (N_5678,N_5594,N_5544);
or U5679 (N_5679,N_5595,N_5549);
and U5680 (N_5680,N_5581,N_5545);
nor U5681 (N_5681,N_5558,N_5539);
nor U5682 (N_5682,N_5551,N_5518);
or U5683 (N_5683,N_5591,N_5504);
nand U5684 (N_5684,N_5567,N_5582);
and U5685 (N_5685,N_5567,N_5535);
nor U5686 (N_5686,N_5573,N_5504);
nand U5687 (N_5687,N_5521,N_5583);
nor U5688 (N_5688,N_5565,N_5560);
nor U5689 (N_5689,N_5558,N_5599);
and U5690 (N_5690,N_5569,N_5558);
xnor U5691 (N_5691,N_5547,N_5576);
xnor U5692 (N_5692,N_5552,N_5520);
nor U5693 (N_5693,N_5592,N_5587);
xnor U5694 (N_5694,N_5530,N_5566);
nand U5695 (N_5695,N_5573,N_5590);
nand U5696 (N_5696,N_5552,N_5538);
or U5697 (N_5697,N_5562,N_5515);
nor U5698 (N_5698,N_5533,N_5578);
nand U5699 (N_5699,N_5568,N_5575);
xor U5700 (N_5700,N_5676,N_5670);
and U5701 (N_5701,N_5694,N_5657);
or U5702 (N_5702,N_5613,N_5665);
or U5703 (N_5703,N_5647,N_5658);
nor U5704 (N_5704,N_5644,N_5673);
nand U5705 (N_5705,N_5661,N_5690);
and U5706 (N_5706,N_5693,N_5696);
or U5707 (N_5707,N_5675,N_5626);
nor U5708 (N_5708,N_5629,N_5648);
nand U5709 (N_5709,N_5680,N_5643);
xnor U5710 (N_5710,N_5667,N_5636);
nor U5711 (N_5711,N_5668,N_5641);
xor U5712 (N_5712,N_5642,N_5682);
nand U5713 (N_5713,N_5607,N_5630);
or U5714 (N_5714,N_5650,N_5600);
nor U5715 (N_5715,N_5663,N_5632);
xor U5716 (N_5716,N_5691,N_5604);
xnor U5717 (N_5717,N_5654,N_5698);
nand U5718 (N_5718,N_5679,N_5603);
or U5719 (N_5719,N_5606,N_5646);
nand U5720 (N_5720,N_5683,N_5627);
nor U5721 (N_5721,N_5678,N_5635);
and U5722 (N_5722,N_5669,N_5621);
and U5723 (N_5723,N_5601,N_5686);
nand U5724 (N_5724,N_5656,N_5649);
xnor U5725 (N_5725,N_5674,N_5645);
xnor U5726 (N_5726,N_5625,N_5618);
nor U5727 (N_5727,N_5611,N_5628);
nor U5728 (N_5728,N_5659,N_5660);
nand U5729 (N_5729,N_5697,N_5640);
nand U5730 (N_5730,N_5681,N_5652);
or U5731 (N_5731,N_5605,N_5609);
nor U5732 (N_5732,N_5633,N_5602);
nand U5733 (N_5733,N_5638,N_5620);
xor U5734 (N_5734,N_5608,N_5623);
or U5735 (N_5735,N_5685,N_5631);
and U5736 (N_5736,N_5637,N_5617);
nand U5737 (N_5737,N_5653,N_5684);
or U5738 (N_5738,N_5639,N_5688);
and U5739 (N_5739,N_5634,N_5610);
nand U5740 (N_5740,N_5671,N_5666);
and U5741 (N_5741,N_5672,N_5612);
and U5742 (N_5742,N_5622,N_5662);
or U5743 (N_5743,N_5624,N_5689);
nor U5744 (N_5744,N_5687,N_5695);
or U5745 (N_5745,N_5655,N_5664);
xnor U5746 (N_5746,N_5619,N_5614);
nand U5747 (N_5747,N_5699,N_5651);
and U5748 (N_5748,N_5615,N_5616);
and U5749 (N_5749,N_5692,N_5677);
and U5750 (N_5750,N_5692,N_5638);
and U5751 (N_5751,N_5695,N_5686);
nor U5752 (N_5752,N_5602,N_5623);
nand U5753 (N_5753,N_5651,N_5697);
nor U5754 (N_5754,N_5654,N_5681);
nor U5755 (N_5755,N_5619,N_5602);
or U5756 (N_5756,N_5656,N_5690);
nor U5757 (N_5757,N_5634,N_5638);
xor U5758 (N_5758,N_5617,N_5663);
and U5759 (N_5759,N_5689,N_5631);
and U5760 (N_5760,N_5678,N_5604);
and U5761 (N_5761,N_5668,N_5639);
nand U5762 (N_5762,N_5601,N_5644);
nand U5763 (N_5763,N_5622,N_5654);
nor U5764 (N_5764,N_5648,N_5625);
and U5765 (N_5765,N_5622,N_5657);
nor U5766 (N_5766,N_5604,N_5650);
nand U5767 (N_5767,N_5608,N_5683);
and U5768 (N_5768,N_5641,N_5649);
or U5769 (N_5769,N_5614,N_5633);
xnor U5770 (N_5770,N_5621,N_5650);
nand U5771 (N_5771,N_5635,N_5608);
and U5772 (N_5772,N_5639,N_5647);
or U5773 (N_5773,N_5622,N_5656);
xnor U5774 (N_5774,N_5639,N_5662);
xor U5775 (N_5775,N_5631,N_5600);
and U5776 (N_5776,N_5651,N_5644);
and U5777 (N_5777,N_5615,N_5651);
nor U5778 (N_5778,N_5660,N_5630);
or U5779 (N_5779,N_5670,N_5654);
and U5780 (N_5780,N_5615,N_5690);
xnor U5781 (N_5781,N_5675,N_5613);
or U5782 (N_5782,N_5680,N_5656);
nor U5783 (N_5783,N_5674,N_5634);
xnor U5784 (N_5784,N_5666,N_5694);
nand U5785 (N_5785,N_5665,N_5684);
and U5786 (N_5786,N_5603,N_5616);
xnor U5787 (N_5787,N_5686,N_5672);
xor U5788 (N_5788,N_5646,N_5684);
xor U5789 (N_5789,N_5689,N_5630);
or U5790 (N_5790,N_5695,N_5614);
xor U5791 (N_5791,N_5651,N_5605);
nand U5792 (N_5792,N_5678,N_5618);
xnor U5793 (N_5793,N_5621,N_5692);
and U5794 (N_5794,N_5604,N_5676);
nand U5795 (N_5795,N_5676,N_5641);
nand U5796 (N_5796,N_5688,N_5660);
nand U5797 (N_5797,N_5658,N_5622);
or U5798 (N_5798,N_5639,N_5627);
nor U5799 (N_5799,N_5695,N_5642);
and U5800 (N_5800,N_5748,N_5799);
and U5801 (N_5801,N_5798,N_5727);
xor U5802 (N_5802,N_5701,N_5704);
xnor U5803 (N_5803,N_5715,N_5746);
nand U5804 (N_5804,N_5794,N_5756);
nor U5805 (N_5805,N_5767,N_5789);
or U5806 (N_5806,N_5710,N_5790);
or U5807 (N_5807,N_5791,N_5788);
nand U5808 (N_5808,N_5784,N_5730);
or U5809 (N_5809,N_5753,N_5703);
nand U5810 (N_5810,N_5757,N_5754);
nor U5811 (N_5811,N_5713,N_5786);
and U5812 (N_5812,N_5708,N_5705);
and U5813 (N_5813,N_5772,N_5702);
and U5814 (N_5814,N_5711,N_5751);
nor U5815 (N_5815,N_5734,N_5783);
and U5816 (N_5816,N_5774,N_5712);
nor U5817 (N_5817,N_5747,N_5777);
nand U5818 (N_5818,N_5796,N_5787);
or U5819 (N_5819,N_5760,N_5755);
or U5820 (N_5820,N_5732,N_5762);
and U5821 (N_5821,N_5773,N_5735);
nand U5822 (N_5822,N_5766,N_5771);
xnor U5823 (N_5823,N_5758,N_5706);
nor U5824 (N_5824,N_5728,N_5700);
nor U5825 (N_5825,N_5793,N_5724);
nand U5826 (N_5826,N_5733,N_5779);
and U5827 (N_5827,N_5721,N_5720);
or U5828 (N_5828,N_5719,N_5775);
nand U5829 (N_5829,N_5776,N_5723);
nor U5830 (N_5830,N_5741,N_5749);
and U5831 (N_5831,N_5765,N_5739);
xnor U5832 (N_5832,N_5792,N_5778);
nor U5833 (N_5833,N_5743,N_5738);
nand U5834 (N_5834,N_5785,N_5737);
and U5835 (N_5835,N_5740,N_5731);
xor U5836 (N_5836,N_5717,N_5714);
nand U5837 (N_5837,N_5742,N_5725);
or U5838 (N_5838,N_5726,N_5745);
nor U5839 (N_5839,N_5781,N_5716);
and U5840 (N_5840,N_5718,N_5752);
and U5841 (N_5841,N_5782,N_5770);
or U5842 (N_5842,N_5759,N_5768);
nor U5843 (N_5843,N_5729,N_5707);
and U5844 (N_5844,N_5761,N_5750);
xor U5845 (N_5845,N_5744,N_5763);
xor U5846 (N_5846,N_5769,N_5795);
nor U5847 (N_5847,N_5797,N_5722);
or U5848 (N_5848,N_5736,N_5780);
xor U5849 (N_5849,N_5764,N_5709);
xor U5850 (N_5850,N_5728,N_5746);
or U5851 (N_5851,N_5766,N_5745);
xnor U5852 (N_5852,N_5728,N_5701);
nand U5853 (N_5853,N_5725,N_5798);
xnor U5854 (N_5854,N_5746,N_5754);
nand U5855 (N_5855,N_5793,N_5768);
and U5856 (N_5856,N_5739,N_5705);
nor U5857 (N_5857,N_5783,N_5763);
and U5858 (N_5858,N_5707,N_5770);
nor U5859 (N_5859,N_5713,N_5710);
xnor U5860 (N_5860,N_5724,N_5797);
nor U5861 (N_5861,N_5759,N_5706);
xnor U5862 (N_5862,N_5762,N_5745);
xor U5863 (N_5863,N_5766,N_5755);
nand U5864 (N_5864,N_5709,N_5734);
and U5865 (N_5865,N_5796,N_5702);
or U5866 (N_5866,N_5798,N_5779);
and U5867 (N_5867,N_5703,N_5739);
and U5868 (N_5868,N_5722,N_5729);
and U5869 (N_5869,N_5731,N_5797);
nor U5870 (N_5870,N_5708,N_5754);
and U5871 (N_5871,N_5776,N_5728);
nor U5872 (N_5872,N_5763,N_5757);
and U5873 (N_5873,N_5747,N_5727);
and U5874 (N_5874,N_5722,N_5775);
nand U5875 (N_5875,N_5770,N_5716);
nor U5876 (N_5876,N_5763,N_5717);
or U5877 (N_5877,N_5791,N_5767);
or U5878 (N_5878,N_5724,N_5772);
and U5879 (N_5879,N_5779,N_5708);
nand U5880 (N_5880,N_5737,N_5753);
nor U5881 (N_5881,N_5745,N_5706);
and U5882 (N_5882,N_5709,N_5784);
or U5883 (N_5883,N_5762,N_5759);
nor U5884 (N_5884,N_5767,N_5793);
nor U5885 (N_5885,N_5747,N_5733);
xor U5886 (N_5886,N_5714,N_5748);
and U5887 (N_5887,N_5707,N_5740);
nand U5888 (N_5888,N_5703,N_5720);
nand U5889 (N_5889,N_5736,N_5792);
nor U5890 (N_5890,N_5703,N_5727);
xor U5891 (N_5891,N_5749,N_5729);
nand U5892 (N_5892,N_5797,N_5728);
nand U5893 (N_5893,N_5782,N_5732);
or U5894 (N_5894,N_5722,N_5799);
xnor U5895 (N_5895,N_5733,N_5719);
and U5896 (N_5896,N_5719,N_5765);
nor U5897 (N_5897,N_5725,N_5750);
nor U5898 (N_5898,N_5758,N_5717);
nand U5899 (N_5899,N_5720,N_5775);
nand U5900 (N_5900,N_5897,N_5863);
or U5901 (N_5901,N_5816,N_5809);
and U5902 (N_5902,N_5815,N_5827);
or U5903 (N_5903,N_5831,N_5867);
xor U5904 (N_5904,N_5825,N_5830);
nor U5905 (N_5905,N_5852,N_5886);
nand U5906 (N_5906,N_5849,N_5874);
nand U5907 (N_5907,N_5870,N_5884);
xnor U5908 (N_5908,N_5848,N_5839);
or U5909 (N_5909,N_5808,N_5892);
and U5910 (N_5910,N_5823,N_5860);
or U5911 (N_5911,N_5856,N_5889);
xnor U5912 (N_5912,N_5851,N_5829);
nand U5913 (N_5913,N_5803,N_5869);
nor U5914 (N_5914,N_5838,N_5850);
and U5915 (N_5915,N_5800,N_5842);
nor U5916 (N_5916,N_5887,N_5840);
nor U5917 (N_5917,N_5841,N_5833);
nor U5918 (N_5918,N_5855,N_5805);
or U5919 (N_5919,N_5821,N_5801);
nand U5920 (N_5920,N_5806,N_5822);
and U5921 (N_5921,N_5812,N_5802);
and U5922 (N_5922,N_5862,N_5824);
nor U5923 (N_5923,N_5868,N_5895);
nor U5924 (N_5924,N_5807,N_5883);
nor U5925 (N_5925,N_5875,N_5837);
nor U5926 (N_5926,N_5873,N_5836);
or U5927 (N_5927,N_5858,N_5846);
and U5928 (N_5928,N_5832,N_5891);
xnor U5929 (N_5929,N_5804,N_5854);
xor U5930 (N_5930,N_5845,N_5820);
xnor U5931 (N_5931,N_5826,N_5885);
nor U5932 (N_5932,N_5882,N_5810);
xor U5933 (N_5933,N_5890,N_5879);
and U5934 (N_5934,N_5893,N_5864);
nand U5935 (N_5935,N_5817,N_5866);
and U5936 (N_5936,N_5877,N_5818);
and U5937 (N_5937,N_5828,N_5888);
and U5938 (N_5938,N_5834,N_5896);
and U5939 (N_5939,N_5872,N_5876);
and U5940 (N_5940,N_5853,N_5881);
nor U5941 (N_5941,N_5835,N_5813);
nor U5942 (N_5942,N_5898,N_5811);
nand U5943 (N_5943,N_5844,N_5880);
nand U5944 (N_5944,N_5861,N_5814);
or U5945 (N_5945,N_5894,N_5857);
or U5946 (N_5946,N_5865,N_5843);
nor U5947 (N_5947,N_5878,N_5871);
or U5948 (N_5948,N_5859,N_5899);
xor U5949 (N_5949,N_5819,N_5847);
nand U5950 (N_5950,N_5801,N_5818);
or U5951 (N_5951,N_5856,N_5817);
nor U5952 (N_5952,N_5802,N_5881);
and U5953 (N_5953,N_5882,N_5884);
xor U5954 (N_5954,N_5857,N_5808);
nor U5955 (N_5955,N_5848,N_5813);
xnor U5956 (N_5956,N_5810,N_5808);
xor U5957 (N_5957,N_5834,N_5893);
nor U5958 (N_5958,N_5873,N_5881);
or U5959 (N_5959,N_5885,N_5832);
xor U5960 (N_5960,N_5838,N_5871);
xor U5961 (N_5961,N_5853,N_5823);
nor U5962 (N_5962,N_5877,N_5852);
xnor U5963 (N_5963,N_5820,N_5834);
xor U5964 (N_5964,N_5846,N_5828);
nand U5965 (N_5965,N_5833,N_5899);
nor U5966 (N_5966,N_5897,N_5849);
nor U5967 (N_5967,N_5868,N_5887);
nor U5968 (N_5968,N_5845,N_5852);
or U5969 (N_5969,N_5886,N_5896);
nand U5970 (N_5970,N_5805,N_5827);
nor U5971 (N_5971,N_5868,N_5826);
nor U5972 (N_5972,N_5892,N_5842);
and U5973 (N_5973,N_5849,N_5882);
nor U5974 (N_5974,N_5899,N_5884);
nand U5975 (N_5975,N_5843,N_5800);
and U5976 (N_5976,N_5842,N_5801);
nor U5977 (N_5977,N_5870,N_5857);
xor U5978 (N_5978,N_5821,N_5831);
xor U5979 (N_5979,N_5814,N_5890);
and U5980 (N_5980,N_5825,N_5844);
or U5981 (N_5981,N_5822,N_5871);
and U5982 (N_5982,N_5868,N_5823);
and U5983 (N_5983,N_5802,N_5844);
and U5984 (N_5984,N_5830,N_5842);
and U5985 (N_5985,N_5805,N_5869);
or U5986 (N_5986,N_5851,N_5844);
nand U5987 (N_5987,N_5875,N_5827);
and U5988 (N_5988,N_5800,N_5866);
xnor U5989 (N_5989,N_5853,N_5860);
nor U5990 (N_5990,N_5874,N_5807);
and U5991 (N_5991,N_5859,N_5849);
nand U5992 (N_5992,N_5875,N_5858);
or U5993 (N_5993,N_5840,N_5861);
and U5994 (N_5994,N_5883,N_5850);
and U5995 (N_5995,N_5899,N_5880);
nor U5996 (N_5996,N_5838,N_5851);
and U5997 (N_5997,N_5860,N_5829);
nor U5998 (N_5998,N_5809,N_5805);
or U5999 (N_5999,N_5879,N_5851);
and U6000 (N_6000,N_5933,N_5994);
and U6001 (N_6001,N_5900,N_5939);
or U6002 (N_6002,N_5951,N_5967);
or U6003 (N_6003,N_5905,N_5927);
or U6004 (N_6004,N_5907,N_5993);
nand U6005 (N_6005,N_5942,N_5990);
and U6006 (N_6006,N_5964,N_5949);
and U6007 (N_6007,N_5986,N_5911);
and U6008 (N_6008,N_5935,N_5973);
and U6009 (N_6009,N_5981,N_5966);
and U6010 (N_6010,N_5956,N_5945);
nor U6011 (N_6011,N_5932,N_5955);
nand U6012 (N_6012,N_5915,N_5902);
or U6013 (N_6013,N_5906,N_5953);
xnor U6014 (N_6014,N_5926,N_5919);
nand U6015 (N_6015,N_5974,N_5987);
or U6016 (N_6016,N_5909,N_5952);
and U6017 (N_6017,N_5920,N_5989);
nor U6018 (N_6018,N_5929,N_5924);
or U6019 (N_6019,N_5961,N_5957);
xor U6020 (N_6020,N_5910,N_5997);
or U6021 (N_6021,N_5934,N_5930);
nor U6022 (N_6022,N_5980,N_5903);
xnor U6023 (N_6023,N_5959,N_5936);
xnor U6024 (N_6024,N_5962,N_5976);
nor U6025 (N_6025,N_5999,N_5960);
or U6026 (N_6026,N_5925,N_5963);
xor U6027 (N_6027,N_5977,N_5992);
xor U6028 (N_6028,N_5917,N_5904);
and U6029 (N_6029,N_5908,N_5913);
nor U6030 (N_6030,N_5916,N_5931);
xnor U6031 (N_6031,N_5995,N_5948);
nor U6032 (N_6032,N_5979,N_5914);
xor U6033 (N_6033,N_5944,N_5991);
nand U6034 (N_6034,N_5950,N_5965);
nand U6035 (N_6035,N_5937,N_5972);
and U6036 (N_6036,N_5943,N_5938);
or U6037 (N_6037,N_5928,N_5921);
nand U6038 (N_6038,N_5968,N_5922);
nor U6039 (N_6039,N_5918,N_5984);
xor U6040 (N_6040,N_5969,N_5998);
nor U6041 (N_6041,N_5983,N_5940);
or U6042 (N_6042,N_5982,N_5912);
nand U6043 (N_6043,N_5978,N_5985);
nor U6044 (N_6044,N_5954,N_5958);
xnor U6045 (N_6045,N_5996,N_5970);
and U6046 (N_6046,N_5946,N_5947);
xor U6047 (N_6047,N_5971,N_5988);
nor U6048 (N_6048,N_5923,N_5941);
nand U6049 (N_6049,N_5975,N_5901);
xor U6050 (N_6050,N_5959,N_5944);
nor U6051 (N_6051,N_5957,N_5979);
or U6052 (N_6052,N_5919,N_5963);
and U6053 (N_6053,N_5969,N_5981);
or U6054 (N_6054,N_5921,N_5976);
and U6055 (N_6055,N_5929,N_5985);
and U6056 (N_6056,N_5909,N_5945);
and U6057 (N_6057,N_5986,N_5993);
or U6058 (N_6058,N_5977,N_5959);
xor U6059 (N_6059,N_5954,N_5965);
xor U6060 (N_6060,N_5900,N_5985);
and U6061 (N_6061,N_5935,N_5902);
nand U6062 (N_6062,N_5946,N_5982);
and U6063 (N_6063,N_5948,N_5943);
nand U6064 (N_6064,N_5995,N_5943);
and U6065 (N_6065,N_5917,N_5959);
nor U6066 (N_6066,N_5955,N_5935);
or U6067 (N_6067,N_5921,N_5975);
nor U6068 (N_6068,N_5933,N_5980);
and U6069 (N_6069,N_5970,N_5929);
or U6070 (N_6070,N_5902,N_5942);
nor U6071 (N_6071,N_5960,N_5906);
nor U6072 (N_6072,N_5968,N_5992);
xnor U6073 (N_6073,N_5908,N_5950);
and U6074 (N_6074,N_5949,N_5994);
nand U6075 (N_6075,N_5918,N_5994);
nor U6076 (N_6076,N_5966,N_5998);
xnor U6077 (N_6077,N_5996,N_5983);
nor U6078 (N_6078,N_5979,N_5986);
and U6079 (N_6079,N_5999,N_5916);
xor U6080 (N_6080,N_5952,N_5965);
and U6081 (N_6081,N_5931,N_5999);
or U6082 (N_6082,N_5946,N_5973);
nor U6083 (N_6083,N_5910,N_5953);
xnor U6084 (N_6084,N_5904,N_5914);
xor U6085 (N_6085,N_5906,N_5973);
nand U6086 (N_6086,N_5908,N_5994);
nor U6087 (N_6087,N_5978,N_5940);
or U6088 (N_6088,N_5938,N_5921);
nand U6089 (N_6089,N_5925,N_5901);
nand U6090 (N_6090,N_5973,N_5912);
nor U6091 (N_6091,N_5978,N_5941);
nor U6092 (N_6092,N_5977,N_5926);
or U6093 (N_6093,N_5904,N_5927);
nand U6094 (N_6094,N_5910,N_5915);
nor U6095 (N_6095,N_5962,N_5979);
nor U6096 (N_6096,N_5941,N_5971);
nand U6097 (N_6097,N_5963,N_5992);
and U6098 (N_6098,N_5900,N_5978);
xor U6099 (N_6099,N_5982,N_5972);
xnor U6100 (N_6100,N_6002,N_6067);
nand U6101 (N_6101,N_6061,N_6048);
nor U6102 (N_6102,N_6009,N_6071);
xor U6103 (N_6103,N_6030,N_6017);
nand U6104 (N_6104,N_6095,N_6052);
nor U6105 (N_6105,N_6053,N_6097);
xnor U6106 (N_6106,N_6084,N_6059);
and U6107 (N_6107,N_6043,N_6062);
xnor U6108 (N_6108,N_6019,N_6023);
nor U6109 (N_6109,N_6070,N_6031);
or U6110 (N_6110,N_6081,N_6013);
xnor U6111 (N_6111,N_6049,N_6054);
and U6112 (N_6112,N_6088,N_6069);
xor U6113 (N_6113,N_6055,N_6010);
nor U6114 (N_6114,N_6068,N_6000);
xor U6115 (N_6115,N_6011,N_6079);
xor U6116 (N_6116,N_6027,N_6087);
xor U6117 (N_6117,N_6096,N_6001);
nand U6118 (N_6118,N_6036,N_6066);
xor U6119 (N_6119,N_6012,N_6051);
and U6120 (N_6120,N_6037,N_6014);
nand U6121 (N_6121,N_6057,N_6029);
and U6122 (N_6122,N_6025,N_6083);
nor U6123 (N_6123,N_6038,N_6047);
xor U6124 (N_6124,N_6045,N_6040);
and U6125 (N_6125,N_6039,N_6042);
nand U6126 (N_6126,N_6021,N_6065);
xor U6127 (N_6127,N_6015,N_6074);
nand U6128 (N_6128,N_6077,N_6032);
or U6129 (N_6129,N_6033,N_6018);
or U6130 (N_6130,N_6034,N_6024);
nand U6131 (N_6131,N_6075,N_6080);
and U6132 (N_6132,N_6056,N_6007);
and U6133 (N_6133,N_6003,N_6086);
xnor U6134 (N_6134,N_6092,N_6098);
nor U6135 (N_6135,N_6060,N_6035);
nor U6136 (N_6136,N_6016,N_6064);
nor U6137 (N_6137,N_6078,N_6006);
nor U6138 (N_6138,N_6041,N_6076);
nand U6139 (N_6139,N_6073,N_6058);
xnor U6140 (N_6140,N_6090,N_6020);
nand U6141 (N_6141,N_6093,N_6085);
and U6142 (N_6142,N_6026,N_6046);
nand U6143 (N_6143,N_6022,N_6063);
and U6144 (N_6144,N_6008,N_6094);
and U6145 (N_6145,N_6089,N_6028);
and U6146 (N_6146,N_6072,N_6005);
or U6147 (N_6147,N_6050,N_6082);
and U6148 (N_6148,N_6091,N_6004);
nand U6149 (N_6149,N_6099,N_6044);
or U6150 (N_6150,N_6088,N_6028);
or U6151 (N_6151,N_6072,N_6008);
xnor U6152 (N_6152,N_6060,N_6061);
or U6153 (N_6153,N_6070,N_6059);
or U6154 (N_6154,N_6071,N_6040);
nand U6155 (N_6155,N_6070,N_6029);
nor U6156 (N_6156,N_6028,N_6023);
or U6157 (N_6157,N_6093,N_6008);
or U6158 (N_6158,N_6010,N_6031);
or U6159 (N_6159,N_6061,N_6083);
nand U6160 (N_6160,N_6026,N_6067);
xnor U6161 (N_6161,N_6063,N_6061);
nand U6162 (N_6162,N_6043,N_6019);
or U6163 (N_6163,N_6045,N_6003);
or U6164 (N_6164,N_6020,N_6010);
or U6165 (N_6165,N_6034,N_6013);
and U6166 (N_6166,N_6070,N_6008);
or U6167 (N_6167,N_6016,N_6073);
and U6168 (N_6168,N_6035,N_6033);
or U6169 (N_6169,N_6079,N_6077);
xor U6170 (N_6170,N_6070,N_6087);
or U6171 (N_6171,N_6088,N_6089);
and U6172 (N_6172,N_6054,N_6004);
xnor U6173 (N_6173,N_6069,N_6065);
nand U6174 (N_6174,N_6077,N_6041);
and U6175 (N_6175,N_6086,N_6019);
xor U6176 (N_6176,N_6084,N_6046);
xor U6177 (N_6177,N_6035,N_6012);
xnor U6178 (N_6178,N_6039,N_6057);
or U6179 (N_6179,N_6000,N_6053);
nor U6180 (N_6180,N_6049,N_6004);
or U6181 (N_6181,N_6094,N_6061);
nor U6182 (N_6182,N_6096,N_6055);
nor U6183 (N_6183,N_6020,N_6011);
nor U6184 (N_6184,N_6037,N_6018);
xnor U6185 (N_6185,N_6073,N_6031);
nor U6186 (N_6186,N_6099,N_6072);
nand U6187 (N_6187,N_6037,N_6082);
nand U6188 (N_6188,N_6061,N_6097);
xnor U6189 (N_6189,N_6009,N_6030);
or U6190 (N_6190,N_6097,N_6040);
and U6191 (N_6191,N_6093,N_6088);
xnor U6192 (N_6192,N_6019,N_6092);
or U6193 (N_6193,N_6040,N_6069);
xnor U6194 (N_6194,N_6019,N_6091);
or U6195 (N_6195,N_6061,N_6084);
nand U6196 (N_6196,N_6016,N_6033);
or U6197 (N_6197,N_6012,N_6092);
nand U6198 (N_6198,N_6062,N_6088);
and U6199 (N_6199,N_6026,N_6014);
nand U6200 (N_6200,N_6108,N_6123);
xnor U6201 (N_6201,N_6145,N_6106);
xor U6202 (N_6202,N_6137,N_6150);
nand U6203 (N_6203,N_6158,N_6181);
nor U6204 (N_6204,N_6154,N_6174);
nand U6205 (N_6205,N_6111,N_6199);
nand U6206 (N_6206,N_6172,N_6122);
and U6207 (N_6207,N_6162,N_6104);
nand U6208 (N_6208,N_6125,N_6135);
nor U6209 (N_6209,N_6148,N_6159);
nor U6210 (N_6210,N_6192,N_6140);
nor U6211 (N_6211,N_6151,N_6179);
or U6212 (N_6212,N_6149,N_6129);
nand U6213 (N_6213,N_6198,N_6147);
xnor U6214 (N_6214,N_6102,N_6136);
xor U6215 (N_6215,N_6146,N_6113);
nand U6216 (N_6216,N_6141,N_6163);
and U6217 (N_6217,N_6117,N_6124);
and U6218 (N_6218,N_6166,N_6171);
nor U6219 (N_6219,N_6127,N_6153);
nor U6220 (N_6220,N_6160,N_6112);
nand U6221 (N_6221,N_6116,N_6196);
xnor U6222 (N_6222,N_6169,N_6119);
xnor U6223 (N_6223,N_6131,N_6175);
or U6224 (N_6224,N_6186,N_6189);
and U6225 (N_6225,N_6164,N_6110);
nor U6226 (N_6226,N_6118,N_6178);
nor U6227 (N_6227,N_6143,N_6190);
and U6228 (N_6228,N_6121,N_6168);
xnor U6229 (N_6229,N_6115,N_6182);
nand U6230 (N_6230,N_6173,N_6139);
or U6231 (N_6231,N_6130,N_6194);
and U6232 (N_6232,N_6180,N_6193);
nor U6233 (N_6233,N_6133,N_6144);
nor U6234 (N_6234,N_6165,N_6167);
or U6235 (N_6235,N_6156,N_6185);
and U6236 (N_6236,N_6126,N_6177);
and U6237 (N_6237,N_6195,N_6187);
xor U6238 (N_6238,N_6183,N_6184);
or U6239 (N_6239,N_6152,N_6157);
nor U6240 (N_6240,N_6120,N_6101);
nand U6241 (N_6241,N_6197,N_6176);
nor U6242 (N_6242,N_6191,N_6132);
nand U6243 (N_6243,N_6155,N_6107);
and U6244 (N_6244,N_6114,N_6138);
or U6245 (N_6245,N_6161,N_6109);
and U6246 (N_6246,N_6128,N_6142);
or U6247 (N_6247,N_6134,N_6103);
or U6248 (N_6248,N_6170,N_6105);
xor U6249 (N_6249,N_6188,N_6100);
nand U6250 (N_6250,N_6138,N_6110);
or U6251 (N_6251,N_6143,N_6165);
nand U6252 (N_6252,N_6170,N_6136);
and U6253 (N_6253,N_6154,N_6173);
or U6254 (N_6254,N_6108,N_6132);
xnor U6255 (N_6255,N_6131,N_6102);
nor U6256 (N_6256,N_6191,N_6161);
and U6257 (N_6257,N_6166,N_6138);
nand U6258 (N_6258,N_6199,N_6160);
and U6259 (N_6259,N_6120,N_6151);
nand U6260 (N_6260,N_6114,N_6182);
nor U6261 (N_6261,N_6192,N_6146);
nand U6262 (N_6262,N_6135,N_6173);
nand U6263 (N_6263,N_6151,N_6106);
nand U6264 (N_6264,N_6140,N_6102);
nand U6265 (N_6265,N_6105,N_6157);
or U6266 (N_6266,N_6154,N_6198);
nand U6267 (N_6267,N_6111,N_6131);
nor U6268 (N_6268,N_6199,N_6103);
nand U6269 (N_6269,N_6149,N_6158);
or U6270 (N_6270,N_6120,N_6185);
nand U6271 (N_6271,N_6176,N_6120);
nand U6272 (N_6272,N_6141,N_6135);
xnor U6273 (N_6273,N_6175,N_6174);
nor U6274 (N_6274,N_6170,N_6145);
or U6275 (N_6275,N_6127,N_6198);
xor U6276 (N_6276,N_6126,N_6138);
xnor U6277 (N_6277,N_6102,N_6199);
or U6278 (N_6278,N_6199,N_6135);
xnor U6279 (N_6279,N_6124,N_6114);
nor U6280 (N_6280,N_6188,N_6149);
nor U6281 (N_6281,N_6141,N_6192);
nand U6282 (N_6282,N_6167,N_6137);
nand U6283 (N_6283,N_6182,N_6154);
or U6284 (N_6284,N_6169,N_6189);
or U6285 (N_6285,N_6119,N_6131);
nor U6286 (N_6286,N_6169,N_6138);
nand U6287 (N_6287,N_6171,N_6141);
nand U6288 (N_6288,N_6140,N_6131);
or U6289 (N_6289,N_6172,N_6167);
or U6290 (N_6290,N_6103,N_6190);
and U6291 (N_6291,N_6163,N_6120);
and U6292 (N_6292,N_6100,N_6122);
xnor U6293 (N_6293,N_6170,N_6139);
xnor U6294 (N_6294,N_6172,N_6181);
or U6295 (N_6295,N_6130,N_6133);
xor U6296 (N_6296,N_6155,N_6122);
nand U6297 (N_6297,N_6145,N_6104);
or U6298 (N_6298,N_6178,N_6194);
and U6299 (N_6299,N_6193,N_6147);
nor U6300 (N_6300,N_6227,N_6217);
nand U6301 (N_6301,N_6289,N_6230);
nor U6302 (N_6302,N_6271,N_6236);
nand U6303 (N_6303,N_6263,N_6282);
nand U6304 (N_6304,N_6202,N_6291);
nand U6305 (N_6305,N_6226,N_6212);
or U6306 (N_6306,N_6222,N_6242);
and U6307 (N_6307,N_6209,N_6255);
and U6308 (N_6308,N_6211,N_6286);
xor U6309 (N_6309,N_6228,N_6231);
or U6310 (N_6310,N_6200,N_6294);
and U6311 (N_6311,N_6262,N_6293);
or U6312 (N_6312,N_6279,N_6266);
or U6313 (N_6313,N_6229,N_6288);
and U6314 (N_6314,N_6216,N_6265);
xor U6315 (N_6315,N_6270,N_6237);
and U6316 (N_6316,N_6247,N_6278);
and U6317 (N_6317,N_6243,N_6277);
or U6318 (N_6318,N_6287,N_6240);
xor U6319 (N_6319,N_6281,N_6239);
nor U6320 (N_6320,N_6208,N_6276);
and U6321 (N_6321,N_6207,N_6256);
or U6322 (N_6322,N_6248,N_6296);
nor U6323 (N_6323,N_6213,N_6215);
or U6324 (N_6324,N_6221,N_6290);
nor U6325 (N_6325,N_6232,N_6260);
xor U6326 (N_6326,N_6284,N_6223);
nor U6327 (N_6327,N_6267,N_6275);
or U6328 (N_6328,N_6285,N_6258);
xnor U6329 (N_6329,N_6225,N_6203);
nand U6330 (N_6330,N_6254,N_6218);
xnor U6331 (N_6331,N_6299,N_6206);
xor U6332 (N_6332,N_6257,N_6214);
xor U6333 (N_6333,N_6272,N_6252);
nor U6334 (N_6334,N_6210,N_6233);
or U6335 (N_6335,N_6224,N_6244);
and U6336 (N_6336,N_6269,N_6268);
or U6337 (N_6337,N_6246,N_6251);
xor U6338 (N_6338,N_6201,N_6264);
and U6339 (N_6339,N_6273,N_6249);
xnor U6340 (N_6340,N_6283,N_6235);
xnor U6341 (N_6341,N_6297,N_6245);
or U6342 (N_6342,N_6205,N_6280);
nand U6343 (N_6343,N_6253,N_6292);
and U6344 (N_6344,N_6274,N_6259);
nand U6345 (N_6345,N_6261,N_6238);
xor U6346 (N_6346,N_6250,N_6219);
nand U6347 (N_6347,N_6295,N_6204);
xnor U6348 (N_6348,N_6220,N_6234);
nor U6349 (N_6349,N_6298,N_6241);
xnor U6350 (N_6350,N_6249,N_6258);
or U6351 (N_6351,N_6221,N_6280);
nand U6352 (N_6352,N_6213,N_6296);
nor U6353 (N_6353,N_6266,N_6207);
xor U6354 (N_6354,N_6206,N_6221);
nand U6355 (N_6355,N_6290,N_6206);
nand U6356 (N_6356,N_6239,N_6237);
xor U6357 (N_6357,N_6241,N_6284);
xnor U6358 (N_6358,N_6217,N_6201);
or U6359 (N_6359,N_6243,N_6228);
or U6360 (N_6360,N_6204,N_6272);
or U6361 (N_6361,N_6237,N_6238);
nor U6362 (N_6362,N_6283,N_6232);
xor U6363 (N_6363,N_6200,N_6230);
nand U6364 (N_6364,N_6295,N_6289);
and U6365 (N_6365,N_6275,N_6208);
nand U6366 (N_6366,N_6228,N_6254);
and U6367 (N_6367,N_6252,N_6255);
nor U6368 (N_6368,N_6226,N_6295);
or U6369 (N_6369,N_6259,N_6224);
and U6370 (N_6370,N_6282,N_6244);
or U6371 (N_6371,N_6296,N_6249);
or U6372 (N_6372,N_6291,N_6246);
and U6373 (N_6373,N_6227,N_6209);
and U6374 (N_6374,N_6207,N_6205);
xor U6375 (N_6375,N_6214,N_6248);
and U6376 (N_6376,N_6264,N_6211);
nand U6377 (N_6377,N_6274,N_6280);
or U6378 (N_6378,N_6269,N_6209);
nand U6379 (N_6379,N_6205,N_6219);
xor U6380 (N_6380,N_6225,N_6238);
and U6381 (N_6381,N_6217,N_6251);
nor U6382 (N_6382,N_6288,N_6220);
nor U6383 (N_6383,N_6251,N_6202);
or U6384 (N_6384,N_6222,N_6250);
nor U6385 (N_6385,N_6250,N_6214);
nor U6386 (N_6386,N_6298,N_6230);
or U6387 (N_6387,N_6213,N_6246);
xor U6388 (N_6388,N_6249,N_6245);
nor U6389 (N_6389,N_6243,N_6260);
and U6390 (N_6390,N_6207,N_6203);
nand U6391 (N_6391,N_6231,N_6266);
nand U6392 (N_6392,N_6233,N_6203);
or U6393 (N_6393,N_6276,N_6297);
and U6394 (N_6394,N_6205,N_6291);
nor U6395 (N_6395,N_6221,N_6256);
and U6396 (N_6396,N_6210,N_6280);
or U6397 (N_6397,N_6202,N_6264);
or U6398 (N_6398,N_6252,N_6295);
or U6399 (N_6399,N_6267,N_6226);
or U6400 (N_6400,N_6339,N_6338);
xor U6401 (N_6401,N_6395,N_6345);
nor U6402 (N_6402,N_6306,N_6389);
and U6403 (N_6403,N_6387,N_6320);
nor U6404 (N_6404,N_6322,N_6353);
xor U6405 (N_6405,N_6359,N_6383);
or U6406 (N_6406,N_6388,N_6343);
nor U6407 (N_6407,N_6311,N_6368);
nor U6408 (N_6408,N_6370,N_6386);
and U6409 (N_6409,N_6332,N_6391);
and U6410 (N_6410,N_6327,N_6392);
and U6411 (N_6411,N_6363,N_6364);
xor U6412 (N_6412,N_6309,N_6361);
nand U6413 (N_6413,N_6371,N_6308);
xnor U6414 (N_6414,N_6385,N_6372);
and U6415 (N_6415,N_6367,N_6330);
or U6416 (N_6416,N_6334,N_6346);
or U6417 (N_6417,N_6328,N_6394);
nand U6418 (N_6418,N_6382,N_6300);
nor U6419 (N_6419,N_6356,N_6398);
and U6420 (N_6420,N_6378,N_6399);
nor U6421 (N_6421,N_6342,N_6369);
nand U6422 (N_6422,N_6303,N_6314);
and U6423 (N_6423,N_6373,N_6335);
nand U6424 (N_6424,N_6318,N_6393);
or U6425 (N_6425,N_6331,N_6329);
and U6426 (N_6426,N_6313,N_6305);
xor U6427 (N_6427,N_6319,N_6366);
xor U6428 (N_6428,N_6384,N_6397);
and U6429 (N_6429,N_6350,N_6312);
or U6430 (N_6430,N_6317,N_6362);
nor U6431 (N_6431,N_6316,N_6360);
or U6432 (N_6432,N_6376,N_6377);
nor U6433 (N_6433,N_6380,N_6340);
nor U6434 (N_6434,N_6304,N_6354);
or U6435 (N_6435,N_6315,N_6344);
nand U6436 (N_6436,N_6374,N_6396);
xnor U6437 (N_6437,N_6302,N_6337);
xor U6438 (N_6438,N_6381,N_6324);
or U6439 (N_6439,N_6352,N_6390);
nand U6440 (N_6440,N_6325,N_6326);
nand U6441 (N_6441,N_6310,N_6365);
and U6442 (N_6442,N_6351,N_6336);
nand U6443 (N_6443,N_6348,N_6321);
or U6444 (N_6444,N_6323,N_6341);
and U6445 (N_6445,N_6379,N_6358);
and U6446 (N_6446,N_6375,N_6307);
nor U6447 (N_6447,N_6349,N_6347);
xnor U6448 (N_6448,N_6355,N_6333);
nor U6449 (N_6449,N_6357,N_6301);
nand U6450 (N_6450,N_6364,N_6355);
or U6451 (N_6451,N_6322,N_6324);
or U6452 (N_6452,N_6396,N_6326);
nand U6453 (N_6453,N_6330,N_6331);
or U6454 (N_6454,N_6310,N_6381);
or U6455 (N_6455,N_6301,N_6316);
or U6456 (N_6456,N_6378,N_6389);
nand U6457 (N_6457,N_6373,N_6393);
nor U6458 (N_6458,N_6336,N_6360);
xor U6459 (N_6459,N_6313,N_6352);
and U6460 (N_6460,N_6382,N_6352);
or U6461 (N_6461,N_6309,N_6359);
nand U6462 (N_6462,N_6319,N_6324);
or U6463 (N_6463,N_6378,N_6325);
and U6464 (N_6464,N_6361,N_6349);
nor U6465 (N_6465,N_6365,N_6372);
and U6466 (N_6466,N_6397,N_6374);
nand U6467 (N_6467,N_6365,N_6357);
nor U6468 (N_6468,N_6305,N_6377);
nor U6469 (N_6469,N_6306,N_6345);
xor U6470 (N_6470,N_6318,N_6309);
and U6471 (N_6471,N_6355,N_6366);
nor U6472 (N_6472,N_6391,N_6365);
xor U6473 (N_6473,N_6322,N_6342);
or U6474 (N_6474,N_6382,N_6313);
nand U6475 (N_6475,N_6342,N_6399);
or U6476 (N_6476,N_6375,N_6361);
nand U6477 (N_6477,N_6350,N_6380);
nand U6478 (N_6478,N_6398,N_6342);
xnor U6479 (N_6479,N_6331,N_6327);
and U6480 (N_6480,N_6364,N_6310);
and U6481 (N_6481,N_6307,N_6378);
nor U6482 (N_6482,N_6311,N_6384);
nand U6483 (N_6483,N_6353,N_6347);
nand U6484 (N_6484,N_6349,N_6355);
nand U6485 (N_6485,N_6302,N_6323);
xnor U6486 (N_6486,N_6319,N_6316);
or U6487 (N_6487,N_6343,N_6359);
xor U6488 (N_6488,N_6382,N_6351);
nor U6489 (N_6489,N_6369,N_6387);
and U6490 (N_6490,N_6366,N_6392);
nand U6491 (N_6491,N_6331,N_6358);
xor U6492 (N_6492,N_6355,N_6385);
nor U6493 (N_6493,N_6387,N_6389);
xor U6494 (N_6494,N_6325,N_6394);
xor U6495 (N_6495,N_6305,N_6331);
xnor U6496 (N_6496,N_6386,N_6351);
nor U6497 (N_6497,N_6379,N_6349);
xor U6498 (N_6498,N_6305,N_6337);
or U6499 (N_6499,N_6346,N_6342);
and U6500 (N_6500,N_6486,N_6445);
or U6501 (N_6501,N_6412,N_6484);
nand U6502 (N_6502,N_6404,N_6456);
or U6503 (N_6503,N_6491,N_6488);
and U6504 (N_6504,N_6417,N_6424);
and U6505 (N_6505,N_6494,N_6423);
nand U6506 (N_6506,N_6482,N_6475);
or U6507 (N_6507,N_6439,N_6463);
nor U6508 (N_6508,N_6460,N_6490);
and U6509 (N_6509,N_6419,N_6450);
nand U6510 (N_6510,N_6473,N_6485);
nor U6511 (N_6511,N_6402,N_6405);
xnor U6512 (N_6512,N_6478,N_6479);
nor U6513 (N_6513,N_6410,N_6452);
or U6514 (N_6514,N_6474,N_6407);
or U6515 (N_6515,N_6477,N_6422);
and U6516 (N_6516,N_6489,N_6470);
or U6517 (N_6517,N_6420,N_6472);
and U6518 (N_6518,N_6468,N_6443);
or U6519 (N_6519,N_6480,N_6454);
and U6520 (N_6520,N_6430,N_6498);
nor U6521 (N_6521,N_6457,N_6401);
and U6522 (N_6522,N_6492,N_6448);
or U6523 (N_6523,N_6435,N_6449);
xor U6524 (N_6524,N_6427,N_6444);
nand U6525 (N_6525,N_6432,N_6464);
xnor U6526 (N_6526,N_6496,N_6428);
nor U6527 (N_6527,N_6413,N_6487);
or U6528 (N_6528,N_6416,N_6411);
nand U6529 (N_6529,N_6471,N_6469);
and U6530 (N_6530,N_6453,N_6499);
nor U6531 (N_6531,N_6447,N_6467);
and U6532 (N_6532,N_6483,N_6414);
nand U6533 (N_6533,N_6438,N_6406);
or U6534 (N_6534,N_6461,N_6403);
xnor U6535 (N_6535,N_6434,N_6462);
nand U6536 (N_6536,N_6481,N_6421);
xor U6537 (N_6537,N_6497,N_6408);
or U6538 (N_6538,N_6466,N_6458);
xnor U6539 (N_6539,N_6441,N_6400);
nor U6540 (N_6540,N_6442,N_6418);
nand U6541 (N_6541,N_6440,N_6493);
or U6542 (N_6542,N_6426,N_6455);
xor U6543 (N_6543,N_6431,N_6446);
or U6544 (N_6544,N_6433,N_6409);
or U6545 (N_6545,N_6476,N_6436);
nor U6546 (N_6546,N_6415,N_6465);
nor U6547 (N_6547,N_6451,N_6437);
nand U6548 (N_6548,N_6429,N_6425);
xnor U6549 (N_6549,N_6495,N_6459);
nand U6550 (N_6550,N_6472,N_6436);
or U6551 (N_6551,N_6407,N_6467);
or U6552 (N_6552,N_6452,N_6428);
nor U6553 (N_6553,N_6433,N_6465);
and U6554 (N_6554,N_6432,N_6488);
and U6555 (N_6555,N_6427,N_6426);
or U6556 (N_6556,N_6467,N_6486);
xnor U6557 (N_6557,N_6443,N_6456);
and U6558 (N_6558,N_6400,N_6402);
nand U6559 (N_6559,N_6441,N_6459);
xor U6560 (N_6560,N_6494,N_6435);
nand U6561 (N_6561,N_6433,N_6442);
nand U6562 (N_6562,N_6445,N_6450);
nor U6563 (N_6563,N_6441,N_6454);
xor U6564 (N_6564,N_6485,N_6448);
or U6565 (N_6565,N_6495,N_6437);
xor U6566 (N_6566,N_6466,N_6424);
or U6567 (N_6567,N_6463,N_6441);
or U6568 (N_6568,N_6489,N_6420);
xor U6569 (N_6569,N_6437,N_6469);
or U6570 (N_6570,N_6450,N_6455);
and U6571 (N_6571,N_6430,N_6406);
xor U6572 (N_6572,N_6423,N_6420);
and U6573 (N_6573,N_6447,N_6436);
xor U6574 (N_6574,N_6438,N_6475);
and U6575 (N_6575,N_6449,N_6420);
and U6576 (N_6576,N_6498,N_6441);
and U6577 (N_6577,N_6413,N_6425);
nor U6578 (N_6578,N_6485,N_6474);
or U6579 (N_6579,N_6487,N_6447);
nand U6580 (N_6580,N_6491,N_6418);
nand U6581 (N_6581,N_6458,N_6447);
nand U6582 (N_6582,N_6430,N_6489);
nand U6583 (N_6583,N_6422,N_6481);
and U6584 (N_6584,N_6484,N_6498);
xor U6585 (N_6585,N_6404,N_6421);
nor U6586 (N_6586,N_6490,N_6466);
nor U6587 (N_6587,N_6422,N_6441);
nand U6588 (N_6588,N_6498,N_6400);
nor U6589 (N_6589,N_6442,N_6439);
or U6590 (N_6590,N_6451,N_6482);
or U6591 (N_6591,N_6478,N_6447);
nor U6592 (N_6592,N_6453,N_6456);
nand U6593 (N_6593,N_6428,N_6468);
or U6594 (N_6594,N_6468,N_6456);
nor U6595 (N_6595,N_6492,N_6423);
nand U6596 (N_6596,N_6429,N_6475);
nand U6597 (N_6597,N_6483,N_6470);
nand U6598 (N_6598,N_6430,N_6478);
xnor U6599 (N_6599,N_6431,N_6450);
or U6600 (N_6600,N_6500,N_6596);
and U6601 (N_6601,N_6559,N_6552);
nor U6602 (N_6602,N_6549,N_6582);
and U6603 (N_6603,N_6541,N_6594);
nor U6604 (N_6604,N_6512,N_6550);
nor U6605 (N_6605,N_6590,N_6543);
xor U6606 (N_6606,N_6530,N_6551);
nor U6607 (N_6607,N_6562,N_6586);
xnor U6608 (N_6608,N_6569,N_6518);
and U6609 (N_6609,N_6517,N_6565);
and U6610 (N_6610,N_6507,N_6591);
or U6611 (N_6611,N_6520,N_6521);
nand U6612 (N_6612,N_6580,N_6598);
nand U6613 (N_6613,N_6575,N_6597);
nor U6614 (N_6614,N_6514,N_6510);
nor U6615 (N_6615,N_6599,N_6576);
xnor U6616 (N_6616,N_6529,N_6557);
nand U6617 (N_6617,N_6563,N_6534);
nand U6618 (N_6618,N_6584,N_6544);
nor U6619 (N_6619,N_6502,N_6513);
or U6620 (N_6620,N_6509,N_6595);
nor U6621 (N_6621,N_6539,N_6573);
and U6622 (N_6622,N_6504,N_6538);
and U6623 (N_6623,N_6525,N_6564);
xor U6624 (N_6624,N_6532,N_6501);
xor U6625 (N_6625,N_6548,N_6556);
nand U6626 (N_6626,N_6593,N_6542);
xnor U6627 (N_6627,N_6545,N_6589);
and U6628 (N_6628,N_6572,N_6527);
or U6629 (N_6629,N_6588,N_6536);
and U6630 (N_6630,N_6511,N_6567);
nand U6631 (N_6631,N_6523,N_6528);
nand U6632 (N_6632,N_6540,N_6579);
and U6633 (N_6633,N_6560,N_6546);
nand U6634 (N_6634,N_6531,N_6571);
or U6635 (N_6635,N_6516,N_6554);
nor U6636 (N_6636,N_6561,N_6583);
xnor U6637 (N_6637,N_6537,N_6574);
or U6638 (N_6638,N_6519,N_6581);
or U6639 (N_6639,N_6524,N_6522);
nand U6640 (N_6640,N_6578,N_6547);
nand U6641 (N_6641,N_6526,N_6553);
nand U6642 (N_6642,N_6555,N_6558);
and U6643 (N_6643,N_6577,N_6508);
xnor U6644 (N_6644,N_6566,N_6533);
nand U6645 (N_6645,N_6585,N_6506);
nand U6646 (N_6646,N_6570,N_6515);
or U6647 (N_6647,N_6503,N_6592);
or U6648 (N_6648,N_6505,N_6535);
and U6649 (N_6649,N_6587,N_6568);
nor U6650 (N_6650,N_6501,N_6589);
nand U6651 (N_6651,N_6585,N_6568);
nand U6652 (N_6652,N_6594,N_6596);
nand U6653 (N_6653,N_6526,N_6514);
and U6654 (N_6654,N_6558,N_6548);
xnor U6655 (N_6655,N_6501,N_6560);
or U6656 (N_6656,N_6564,N_6534);
nor U6657 (N_6657,N_6521,N_6500);
nor U6658 (N_6658,N_6591,N_6581);
and U6659 (N_6659,N_6501,N_6542);
or U6660 (N_6660,N_6549,N_6501);
and U6661 (N_6661,N_6525,N_6579);
nor U6662 (N_6662,N_6507,N_6567);
or U6663 (N_6663,N_6574,N_6519);
nand U6664 (N_6664,N_6563,N_6528);
nand U6665 (N_6665,N_6555,N_6517);
and U6666 (N_6666,N_6556,N_6507);
nand U6667 (N_6667,N_6582,N_6541);
nor U6668 (N_6668,N_6523,N_6511);
nand U6669 (N_6669,N_6523,N_6591);
or U6670 (N_6670,N_6592,N_6586);
xnor U6671 (N_6671,N_6551,N_6529);
nor U6672 (N_6672,N_6543,N_6581);
and U6673 (N_6673,N_6567,N_6579);
xor U6674 (N_6674,N_6507,N_6540);
xor U6675 (N_6675,N_6550,N_6571);
or U6676 (N_6676,N_6539,N_6587);
nand U6677 (N_6677,N_6536,N_6535);
and U6678 (N_6678,N_6522,N_6541);
and U6679 (N_6679,N_6525,N_6594);
xnor U6680 (N_6680,N_6566,N_6585);
nand U6681 (N_6681,N_6541,N_6587);
xnor U6682 (N_6682,N_6519,N_6527);
nor U6683 (N_6683,N_6566,N_6557);
nand U6684 (N_6684,N_6533,N_6575);
nor U6685 (N_6685,N_6521,N_6545);
xor U6686 (N_6686,N_6577,N_6561);
or U6687 (N_6687,N_6546,N_6547);
and U6688 (N_6688,N_6573,N_6574);
and U6689 (N_6689,N_6531,N_6594);
or U6690 (N_6690,N_6544,N_6534);
nand U6691 (N_6691,N_6597,N_6532);
nor U6692 (N_6692,N_6596,N_6574);
xnor U6693 (N_6693,N_6532,N_6545);
and U6694 (N_6694,N_6596,N_6565);
nand U6695 (N_6695,N_6578,N_6522);
nor U6696 (N_6696,N_6518,N_6511);
nand U6697 (N_6697,N_6503,N_6543);
and U6698 (N_6698,N_6511,N_6571);
and U6699 (N_6699,N_6549,N_6530);
nor U6700 (N_6700,N_6673,N_6696);
xnor U6701 (N_6701,N_6678,N_6610);
nand U6702 (N_6702,N_6655,N_6605);
nor U6703 (N_6703,N_6653,N_6659);
nor U6704 (N_6704,N_6625,N_6671);
and U6705 (N_6705,N_6674,N_6656);
and U6706 (N_6706,N_6691,N_6603);
or U6707 (N_6707,N_6684,N_6629);
nand U6708 (N_6708,N_6635,N_6651);
xor U6709 (N_6709,N_6645,N_6658);
nand U6710 (N_6710,N_6617,N_6611);
nand U6711 (N_6711,N_6663,N_6650);
xnor U6712 (N_6712,N_6604,N_6690);
nor U6713 (N_6713,N_6638,N_6685);
xnor U6714 (N_6714,N_6633,N_6680);
or U6715 (N_6715,N_6649,N_6676);
xor U6716 (N_6716,N_6679,N_6698);
or U6717 (N_6717,N_6600,N_6682);
nand U6718 (N_6718,N_6646,N_6697);
and U6719 (N_6719,N_6699,N_6692);
nand U6720 (N_6720,N_6601,N_6677);
nor U6721 (N_6721,N_6606,N_6660);
nor U6722 (N_6722,N_6647,N_6608);
nor U6723 (N_6723,N_6669,N_6687);
or U6724 (N_6724,N_6632,N_6637);
nor U6725 (N_6725,N_6627,N_6641);
or U6726 (N_6726,N_6686,N_6683);
or U6727 (N_6727,N_6672,N_6631);
and U6728 (N_6728,N_6618,N_6642);
or U6729 (N_6729,N_6630,N_6657);
xor U6730 (N_6730,N_6689,N_6664);
nor U6731 (N_6731,N_6621,N_6612);
and U6732 (N_6732,N_6643,N_6607);
nand U6733 (N_6733,N_6654,N_6619);
xnor U6734 (N_6734,N_6616,N_6624);
or U6735 (N_6735,N_6652,N_6662);
xor U6736 (N_6736,N_6668,N_6626);
nand U6737 (N_6737,N_6675,N_6639);
or U6738 (N_6738,N_6623,N_6693);
nand U6739 (N_6739,N_6620,N_6695);
nor U6740 (N_6740,N_6622,N_6640);
nor U6741 (N_6741,N_6670,N_6609);
nor U6742 (N_6742,N_6648,N_6667);
and U6743 (N_6743,N_6688,N_6694);
nor U6744 (N_6744,N_6644,N_6636);
and U6745 (N_6745,N_6628,N_6665);
and U6746 (N_6746,N_6634,N_6661);
or U6747 (N_6747,N_6614,N_6666);
nor U6748 (N_6748,N_6615,N_6602);
nand U6749 (N_6749,N_6613,N_6681);
and U6750 (N_6750,N_6694,N_6682);
nor U6751 (N_6751,N_6614,N_6669);
xnor U6752 (N_6752,N_6681,N_6632);
and U6753 (N_6753,N_6644,N_6672);
xor U6754 (N_6754,N_6609,N_6620);
and U6755 (N_6755,N_6637,N_6678);
and U6756 (N_6756,N_6649,N_6636);
or U6757 (N_6757,N_6636,N_6679);
xnor U6758 (N_6758,N_6611,N_6607);
xor U6759 (N_6759,N_6610,N_6664);
or U6760 (N_6760,N_6620,N_6646);
or U6761 (N_6761,N_6649,N_6664);
nor U6762 (N_6762,N_6669,N_6675);
and U6763 (N_6763,N_6621,N_6697);
and U6764 (N_6764,N_6675,N_6662);
or U6765 (N_6765,N_6608,N_6644);
nor U6766 (N_6766,N_6639,N_6647);
or U6767 (N_6767,N_6612,N_6658);
xnor U6768 (N_6768,N_6685,N_6601);
nand U6769 (N_6769,N_6673,N_6686);
xnor U6770 (N_6770,N_6662,N_6626);
xor U6771 (N_6771,N_6659,N_6638);
or U6772 (N_6772,N_6652,N_6648);
nor U6773 (N_6773,N_6684,N_6606);
xor U6774 (N_6774,N_6657,N_6663);
and U6775 (N_6775,N_6652,N_6619);
and U6776 (N_6776,N_6637,N_6630);
or U6777 (N_6777,N_6680,N_6696);
nor U6778 (N_6778,N_6607,N_6681);
and U6779 (N_6779,N_6608,N_6648);
and U6780 (N_6780,N_6696,N_6695);
xor U6781 (N_6781,N_6664,N_6644);
and U6782 (N_6782,N_6693,N_6692);
or U6783 (N_6783,N_6670,N_6610);
nor U6784 (N_6784,N_6609,N_6611);
nand U6785 (N_6785,N_6637,N_6663);
xor U6786 (N_6786,N_6686,N_6619);
and U6787 (N_6787,N_6604,N_6674);
nand U6788 (N_6788,N_6645,N_6668);
xor U6789 (N_6789,N_6617,N_6612);
nor U6790 (N_6790,N_6650,N_6620);
or U6791 (N_6791,N_6694,N_6609);
and U6792 (N_6792,N_6606,N_6627);
xor U6793 (N_6793,N_6646,N_6657);
and U6794 (N_6794,N_6624,N_6666);
nor U6795 (N_6795,N_6647,N_6698);
nand U6796 (N_6796,N_6649,N_6623);
or U6797 (N_6797,N_6643,N_6629);
and U6798 (N_6798,N_6652,N_6601);
and U6799 (N_6799,N_6639,N_6645);
or U6800 (N_6800,N_6735,N_6790);
nand U6801 (N_6801,N_6798,N_6772);
xor U6802 (N_6802,N_6703,N_6788);
nor U6803 (N_6803,N_6708,N_6747);
or U6804 (N_6804,N_6778,N_6756);
or U6805 (N_6805,N_6757,N_6721);
and U6806 (N_6806,N_6722,N_6780);
or U6807 (N_6807,N_6740,N_6781);
nand U6808 (N_6808,N_6724,N_6746);
and U6809 (N_6809,N_6745,N_6711);
xnor U6810 (N_6810,N_6725,N_6771);
or U6811 (N_6811,N_6718,N_6749);
or U6812 (N_6812,N_6764,N_6794);
nand U6813 (N_6813,N_6753,N_6701);
or U6814 (N_6814,N_6762,N_6752);
xor U6815 (N_6815,N_6720,N_6719);
xor U6816 (N_6816,N_6734,N_6737);
and U6817 (N_6817,N_6732,N_6750);
and U6818 (N_6818,N_6715,N_6786);
or U6819 (N_6819,N_6754,N_6710);
nor U6820 (N_6820,N_6793,N_6712);
nand U6821 (N_6821,N_6792,N_6742);
xor U6822 (N_6822,N_6787,N_6748);
and U6823 (N_6823,N_6799,N_6796);
nor U6824 (N_6824,N_6759,N_6723);
nor U6825 (N_6825,N_6707,N_6702);
nand U6826 (N_6826,N_6782,N_6768);
nand U6827 (N_6827,N_6760,N_6770);
or U6828 (N_6828,N_6726,N_6785);
nand U6829 (N_6829,N_6789,N_6765);
nand U6830 (N_6830,N_6761,N_6767);
xnor U6831 (N_6831,N_6751,N_6705);
nand U6832 (N_6832,N_6727,N_6769);
nand U6833 (N_6833,N_6758,N_6730);
nor U6834 (N_6834,N_6743,N_6777);
or U6835 (N_6835,N_6728,N_6766);
nor U6836 (N_6836,N_6776,N_6733);
or U6837 (N_6837,N_6706,N_6709);
nand U6838 (N_6838,N_6773,N_6736);
nand U6839 (N_6839,N_6741,N_6714);
xor U6840 (N_6840,N_6791,N_6716);
or U6841 (N_6841,N_6755,N_6763);
nand U6842 (N_6842,N_6744,N_6775);
and U6843 (N_6843,N_6795,N_6713);
and U6844 (N_6844,N_6774,N_6729);
nand U6845 (N_6845,N_6797,N_6704);
nor U6846 (N_6846,N_6779,N_6700);
or U6847 (N_6847,N_6738,N_6739);
and U6848 (N_6848,N_6731,N_6784);
nand U6849 (N_6849,N_6717,N_6783);
nor U6850 (N_6850,N_6765,N_6769);
and U6851 (N_6851,N_6735,N_6761);
nand U6852 (N_6852,N_6727,N_6721);
or U6853 (N_6853,N_6701,N_6724);
xnor U6854 (N_6854,N_6734,N_6752);
nor U6855 (N_6855,N_6794,N_6772);
nor U6856 (N_6856,N_6783,N_6781);
and U6857 (N_6857,N_6717,N_6786);
xnor U6858 (N_6858,N_6744,N_6753);
and U6859 (N_6859,N_6748,N_6788);
nor U6860 (N_6860,N_6778,N_6753);
and U6861 (N_6861,N_6733,N_6761);
or U6862 (N_6862,N_6757,N_6716);
nor U6863 (N_6863,N_6768,N_6705);
nand U6864 (N_6864,N_6721,N_6758);
and U6865 (N_6865,N_6703,N_6781);
nor U6866 (N_6866,N_6746,N_6704);
and U6867 (N_6867,N_6725,N_6752);
or U6868 (N_6868,N_6766,N_6763);
nand U6869 (N_6869,N_6722,N_6747);
or U6870 (N_6870,N_6740,N_6782);
nand U6871 (N_6871,N_6756,N_6743);
nand U6872 (N_6872,N_6731,N_6726);
nand U6873 (N_6873,N_6722,N_6776);
nor U6874 (N_6874,N_6706,N_6778);
xnor U6875 (N_6875,N_6728,N_6737);
and U6876 (N_6876,N_6780,N_6750);
nor U6877 (N_6877,N_6798,N_6701);
nand U6878 (N_6878,N_6743,N_6765);
xnor U6879 (N_6879,N_6730,N_6776);
and U6880 (N_6880,N_6752,N_6747);
or U6881 (N_6881,N_6739,N_6712);
or U6882 (N_6882,N_6729,N_6706);
nor U6883 (N_6883,N_6743,N_6737);
xor U6884 (N_6884,N_6759,N_6733);
nand U6885 (N_6885,N_6760,N_6780);
or U6886 (N_6886,N_6799,N_6752);
and U6887 (N_6887,N_6740,N_6737);
xnor U6888 (N_6888,N_6748,N_6720);
xnor U6889 (N_6889,N_6792,N_6747);
or U6890 (N_6890,N_6711,N_6753);
or U6891 (N_6891,N_6720,N_6710);
nor U6892 (N_6892,N_6769,N_6734);
or U6893 (N_6893,N_6792,N_6749);
or U6894 (N_6894,N_6706,N_6775);
and U6895 (N_6895,N_6702,N_6729);
xor U6896 (N_6896,N_6740,N_6774);
or U6897 (N_6897,N_6782,N_6749);
xor U6898 (N_6898,N_6781,N_6710);
nand U6899 (N_6899,N_6794,N_6793);
nor U6900 (N_6900,N_6849,N_6873);
xor U6901 (N_6901,N_6829,N_6817);
or U6902 (N_6902,N_6878,N_6898);
nand U6903 (N_6903,N_6850,N_6876);
nand U6904 (N_6904,N_6802,N_6807);
nor U6905 (N_6905,N_6869,N_6841);
nor U6906 (N_6906,N_6825,N_6835);
or U6907 (N_6907,N_6853,N_6846);
nand U6908 (N_6908,N_6811,N_6805);
or U6909 (N_6909,N_6847,N_6894);
xnor U6910 (N_6910,N_6877,N_6862);
xnor U6911 (N_6911,N_6855,N_6823);
nand U6912 (N_6912,N_6856,N_6834);
or U6913 (N_6913,N_6837,N_6887);
nand U6914 (N_6914,N_6891,N_6806);
nor U6915 (N_6915,N_6871,N_6892);
nand U6916 (N_6916,N_6860,N_6863);
xor U6917 (N_6917,N_6831,N_6833);
or U6918 (N_6918,N_6838,N_6895);
nor U6919 (N_6919,N_6804,N_6840);
xor U6920 (N_6920,N_6879,N_6866);
nor U6921 (N_6921,N_6867,N_6842);
nand U6922 (N_6922,N_6858,N_6821);
nor U6923 (N_6923,N_6865,N_6864);
or U6924 (N_6924,N_6828,N_6819);
xnor U6925 (N_6925,N_6816,N_6803);
and U6926 (N_6926,N_6886,N_6814);
or U6927 (N_6927,N_6896,N_6832);
xnor U6928 (N_6928,N_6827,N_6885);
and U6929 (N_6929,N_6818,N_6888);
xor U6930 (N_6930,N_6890,N_6801);
nor U6931 (N_6931,N_6881,N_6868);
or U6932 (N_6932,N_6800,N_6882);
nand U6933 (N_6933,N_6851,N_6874);
nor U6934 (N_6934,N_6810,N_6848);
nand U6935 (N_6935,N_6883,N_6893);
or U6936 (N_6936,N_6830,N_6859);
and U6937 (N_6937,N_6897,N_6826);
nor U6938 (N_6938,N_6813,N_6854);
nor U6939 (N_6939,N_6815,N_6824);
nand U6940 (N_6940,N_6880,N_6861);
or U6941 (N_6941,N_6809,N_6875);
and U6942 (N_6942,N_6812,N_6822);
and U6943 (N_6943,N_6844,N_6899);
xor U6944 (N_6944,N_6852,N_6820);
or U6945 (N_6945,N_6839,N_6836);
xnor U6946 (N_6946,N_6872,N_6889);
nor U6947 (N_6947,N_6857,N_6808);
xor U6948 (N_6948,N_6870,N_6884);
nor U6949 (N_6949,N_6845,N_6843);
xnor U6950 (N_6950,N_6860,N_6882);
nand U6951 (N_6951,N_6827,N_6872);
and U6952 (N_6952,N_6887,N_6893);
xor U6953 (N_6953,N_6866,N_6887);
and U6954 (N_6954,N_6817,N_6899);
nand U6955 (N_6955,N_6871,N_6852);
and U6956 (N_6956,N_6802,N_6876);
or U6957 (N_6957,N_6833,N_6898);
or U6958 (N_6958,N_6887,N_6858);
xnor U6959 (N_6959,N_6865,N_6896);
nand U6960 (N_6960,N_6833,N_6892);
nor U6961 (N_6961,N_6836,N_6845);
nor U6962 (N_6962,N_6888,N_6887);
and U6963 (N_6963,N_6861,N_6896);
and U6964 (N_6964,N_6865,N_6858);
or U6965 (N_6965,N_6880,N_6891);
or U6966 (N_6966,N_6896,N_6879);
nand U6967 (N_6967,N_6812,N_6807);
or U6968 (N_6968,N_6801,N_6816);
or U6969 (N_6969,N_6845,N_6879);
or U6970 (N_6970,N_6837,N_6891);
nor U6971 (N_6971,N_6830,N_6843);
or U6972 (N_6972,N_6898,N_6834);
nand U6973 (N_6973,N_6836,N_6859);
xnor U6974 (N_6974,N_6873,N_6816);
nor U6975 (N_6975,N_6800,N_6850);
nand U6976 (N_6976,N_6811,N_6851);
and U6977 (N_6977,N_6836,N_6881);
and U6978 (N_6978,N_6880,N_6846);
nor U6979 (N_6979,N_6874,N_6857);
xnor U6980 (N_6980,N_6825,N_6807);
nand U6981 (N_6981,N_6865,N_6868);
nor U6982 (N_6982,N_6855,N_6814);
or U6983 (N_6983,N_6833,N_6806);
and U6984 (N_6984,N_6888,N_6819);
and U6985 (N_6985,N_6822,N_6835);
xnor U6986 (N_6986,N_6891,N_6812);
xnor U6987 (N_6987,N_6806,N_6892);
nand U6988 (N_6988,N_6869,N_6896);
and U6989 (N_6989,N_6813,N_6890);
xor U6990 (N_6990,N_6896,N_6890);
or U6991 (N_6991,N_6856,N_6840);
and U6992 (N_6992,N_6852,N_6804);
nor U6993 (N_6993,N_6816,N_6821);
and U6994 (N_6994,N_6805,N_6808);
nand U6995 (N_6995,N_6813,N_6810);
xnor U6996 (N_6996,N_6826,N_6862);
xor U6997 (N_6997,N_6880,N_6829);
xnor U6998 (N_6998,N_6894,N_6880);
and U6999 (N_6999,N_6805,N_6862);
or U7000 (N_7000,N_6980,N_6954);
and U7001 (N_7001,N_6904,N_6905);
nand U7002 (N_7002,N_6960,N_6919);
or U7003 (N_7003,N_6973,N_6946);
xor U7004 (N_7004,N_6942,N_6948);
nand U7005 (N_7005,N_6950,N_6955);
nand U7006 (N_7006,N_6978,N_6977);
nor U7007 (N_7007,N_6910,N_6961);
xor U7008 (N_7008,N_6997,N_6972);
nor U7009 (N_7009,N_6911,N_6983);
xor U7010 (N_7010,N_6965,N_6974);
or U7011 (N_7011,N_6913,N_6981);
or U7012 (N_7012,N_6941,N_6970);
nor U7013 (N_7013,N_6992,N_6985);
xnor U7014 (N_7014,N_6968,N_6934);
and U7015 (N_7015,N_6902,N_6924);
or U7016 (N_7016,N_6926,N_6999);
nand U7017 (N_7017,N_6909,N_6929);
xnor U7018 (N_7018,N_6971,N_6994);
and U7019 (N_7019,N_6979,N_6949);
nand U7020 (N_7020,N_6903,N_6900);
xor U7021 (N_7021,N_6906,N_6989);
xnor U7022 (N_7022,N_6953,N_6921);
nor U7023 (N_7023,N_6923,N_6957);
nand U7024 (N_7024,N_6986,N_6935);
nand U7025 (N_7025,N_6963,N_6930);
nand U7026 (N_7026,N_6933,N_6995);
and U7027 (N_7027,N_6958,N_6931);
and U7028 (N_7028,N_6916,N_6945);
or U7029 (N_7029,N_6947,N_6915);
xnor U7030 (N_7030,N_6917,N_6984);
and U7031 (N_7031,N_6922,N_6990);
or U7032 (N_7032,N_6925,N_6937);
or U7033 (N_7033,N_6998,N_6988);
or U7034 (N_7034,N_6952,N_6938);
nor U7035 (N_7035,N_6928,N_6912);
xor U7036 (N_7036,N_6944,N_6918);
nand U7037 (N_7037,N_6991,N_6927);
nand U7038 (N_7038,N_6996,N_6943);
xor U7039 (N_7039,N_6967,N_6914);
and U7040 (N_7040,N_6920,N_6940);
or U7041 (N_7041,N_6975,N_6936);
nor U7042 (N_7042,N_6901,N_6962);
nor U7043 (N_7043,N_6969,N_6987);
xor U7044 (N_7044,N_6939,N_6964);
nor U7045 (N_7045,N_6982,N_6908);
or U7046 (N_7046,N_6966,N_6951);
or U7047 (N_7047,N_6932,N_6956);
xnor U7048 (N_7048,N_6976,N_6907);
xnor U7049 (N_7049,N_6993,N_6959);
or U7050 (N_7050,N_6940,N_6934);
and U7051 (N_7051,N_6964,N_6979);
or U7052 (N_7052,N_6955,N_6957);
and U7053 (N_7053,N_6929,N_6924);
nor U7054 (N_7054,N_6914,N_6995);
and U7055 (N_7055,N_6924,N_6954);
or U7056 (N_7056,N_6937,N_6918);
or U7057 (N_7057,N_6978,N_6980);
and U7058 (N_7058,N_6972,N_6942);
or U7059 (N_7059,N_6983,N_6971);
or U7060 (N_7060,N_6952,N_6980);
nand U7061 (N_7061,N_6972,N_6926);
xnor U7062 (N_7062,N_6987,N_6942);
nor U7063 (N_7063,N_6911,N_6976);
nand U7064 (N_7064,N_6901,N_6963);
or U7065 (N_7065,N_6989,N_6949);
xnor U7066 (N_7066,N_6941,N_6994);
or U7067 (N_7067,N_6977,N_6994);
nor U7068 (N_7068,N_6985,N_6974);
and U7069 (N_7069,N_6996,N_6970);
nand U7070 (N_7070,N_6957,N_6985);
or U7071 (N_7071,N_6944,N_6907);
nand U7072 (N_7072,N_6930,N_6931);
nor U7073 (N_7073,N_6999,N_6939);
xor U7074 (N_7074,N_6973,N_6990);
nor U7075 (N_7075,N_6978,N_6928);
and U7076 (N_7076,N_6930,N_6979);
and U7077 (N_7077,N_6980,N_6919);
xnor U7078 (N_7078,N_6923,N_6932);
and U7079 (N_7079,N_6910,N_6939);
or U7080 (N_7080,N_6921,N_6976);
or U7081 (N_7081,N_6900,N_6987);
nand U7082 (N_7082,N_6945,N_6989);
nand U7083 (N_7083,N_6978,N_6903);
xnor U7084 (N_7084,N_6979,N_6985);
xor U7085 (N_7085,N_6979,N_6940);
nor U7086 (N_7086,N_6970,N_6969);
or U7087 (N_7087,N_6949,N_6915);
xnor U7088 (N_7088,N_6928,N_6904);
xor U7089 (N_7089,N_6945,N_6902);
nand U7090 (N_7090,N_6904,N_6985);
nor U7091 (N_7091,N_6906,N_6986);
nor U7092 (N_7092,N_6954,N_6986);
xnor U7093 (N_7093,N_6968,N_6985);
nand U7094 (N_7094,N_6988,N_6906);
nor U7095 (N_7095,N_6955,N_6930);
and U7096 (N_7096,N_6906,N_6950);
nand U7097 (N_7097,N_6982,N_6911);
and U7098 (N_7098,N_6978,N_6918);
or U7099 (N_7099,N_6972,N_6989);
nor U7100 (N_7100,N_7089,N_7047);
and U7101 (N_7101,N_7059,N_7049);
or U7102 (N_7102,N_7053,N_7006);
or U7103 (N_7103,N_7084,N_7090);
nand U7104 (N_7104,N_7095,N_7030);
or U7105 (N_7105,N_7069,N_7011);
nor U7106 (N_7106,N_7033,N_7046);
or U7107 (N_7107,N_7062,N_7036);
nand U7108 (N_7108,N_7094,N_7099);
nand U7109 (N_7109,N_7082,N_7032);
nand U7110 (N_7110,N_7063,N_7067);
nand U7111 (N_7111,N_7042,N_7091);
nand U7112 (N_7112,N_7077,N_7061);
xor U7113 (N_7113,N_7041,N_7000);
nor U7114 (N_7114,N_7086,N_7074);
xnor U7115 (N_7115,N_7092,N_7019);
xor U7116 (N_7116,N_7017,N_7064);
and U7117 (N_7117,N_7037,N_7088);
or U7118 (N_7118,N_7010,N_7001);
and U7119 (N_7119,N_7005,N_7079);
nand U7120 (N_7120,N_7040,N_7075);
or U7121 (N_7121,N_7039,N_7022);
or U7122 (N_7122,N_7013,N_7078);
or U7123 (N_7123,N_7081,N_7003);
or U7124 (N_7124,N_7065,N_7050);
nor U7125 (N_7125,N_7051,N_7021);
xor U7126 (N_7126,N_7070,N_7087);
or U7127 (N_7127,N_7016,N_7066);
nor U7128 (N_7128,N_7024,N_7055);
or U7129 (N_7129,N_7012,N_7080);
xnor U7130 (N_7130,N_7038,N_7007);
xor U7131 (N_7131,N_7073,N_7052);
xor U7132 (N_7132,N_7058,N_7097);
nand U7133 (N_7133,N_7085,N_7096);
xnor U7134 (N_7134,N_7076,N_7020);
xnor U7135 (N_7135,N_7026,N_7028);
nand U7136 (N_7136,N_7093,N_7035);
nand U7137 (N_7137,N_7002,N_7068);
and U7138 (N_7138,N_7014,N_7008);
nor U7139 (N_7139,N_7015,N_7071);
and U7140 (N_7140,N_7048,N_7045);
and U7141 (N_7141,N_7023,N_7072);
nand U7142 (N_7142,N_7044,N_7009);
and U7143 (N_7143,N_7056,N_7043);
or U7144 (N_7144,N_7054,N_7034);
and U7145 (N_7145,N_7004,N_7029);
xor U7146 (N_7146,N_7027,N_7098);
and U7147 (N_7147,N_7083,N_7025);
nor U7148 (N_7148,N_7031,N_7057);
nand U7149 (N_7149,N_7060,N_7018);
xnor U7150 (N_7150,N_7003,N_7078);
xor U7151 (N_7151,N_7050,N_7016);
nand U7152 (N_7152,N_7017,N_7077);
or U7153 (N_7153,N_7035,N_7043);
nand U7154 (N_7154,N_7092,N_7001);
nand U7155 (N_7155,N_7066,N_7093);
nor U7156 (N_7156,N_7050,N_7062);
nand U7157 (N_7157,N_7019,N_7032);
xnor U7158 (N_7158,N_7056,N_7060);
and U7159 (N_7159,N_7018,N_7082);
or U7160 (N_7160,N_7016,N_7089);
and U7161 (N_7161,N_7000,N_7028);
nand U7162 (N_7162,N_7072,N_7011);
nor U7163 (N_7163,N_7021,N_7042);
xnor U7164 (N_7164,N_7097,N_7096);
nand U7165 (N_7165,N_7028,N_7091);
nor U7166 (N_7166,N_7071,N_7059);
or U7167 (N_7167,N_7011,N_7007);
nor U7168 (N_7168,N_7096,N_7041);
nand U7169 (N_7169,N_7005,N_7070);
nand U7170 (N_7170,N_7081,N_7063);
xnor U7171 (N_7171,N_7002,N_7038);
or U7172 (N_7172,N_7010,N_7025);
nand U7173 (N_7173,N_7062,N_7047);
xor U7174 (N_7174,N_7080,N_7060);
nor U7175 (N_7175,N_7074,N_7062);
or U7176 (N_7176,N_7063,N_7071);
xor U7177 (N_7177,N_7018,N_7068);
or U7178 (N_7178,N_7099,N_7088);
or U7179 (N_7179,N_7032,N_7061);
or U7180 (N_7180,N_7082,N_7035);
nand U7181 (N_7181,N_7093,N_7071);
or U7182 (N_7182,N_7076,N_7052);
xnor U7183 (N_7183,N_7065,N_7057);
xor U7184 (N_7184,N_7029,N_7068);
or U7185 (N_7185,N_7087,N_7037);
or U7186 (N_7186,N_7021,N_7090);
nand U7187 (N_7187,N_7008,N_7068);
and U7188 (N_7188,N_7097,N_7007);
or U7189 (N_7189,N_7068,N_7099);
nand U7190 (N_7190,N_7084,N_7094);
nand U7191 (N_7191,N_7023,N_7051);
xor U7192 (N_7192,N_7084,N_7027);
nand U7193 (N_7193,N_7025,N_7008);
or U7194 (N_7194,N_7092,N_7037);
xnor U7195 (N_7195,N_7007,N_7005);
nor U7196 (N_7196,N_7000,N_7060);
nor U7197 (N_7197,N_7049,N_7026);
and U7198 (N_7198,N_7004,N_7035);
and U7199 (N_7199,N_7068,N_7007);
xnor U7200 (N_7200,N_7162,N_7189);
xnor U7201 (N_7201,N_7139,N_7158);
or U7202 (N_7202,N_7104,N_7100);
xor U7203 (N_7203,N_7134,N_7184);
xor U7204 (N_7204,N_7164,N_7153);
and U7205 (N_7205,N_7151,N_7144);
nand U7206 (N_7206,N_7108,N_7119);
nor U7207 (N_7207,N_7143,N_7176);
nor U7208 (N_7208,N_7117,N_7113);
nor U7209 (N_7209,N_7102,N_7112);
nor U7210 (N_7210,N_7181,N_7179);
nand U7211 (N_7211,N_7167,N_7110);
and U7212 (N_7212,N_7115,N_7118);
xor U7213 (N_7213,N_7160,N_7126);
nand U7214 (N_7214,N_7137,N_7141);
xor U7215 (N_7215,N_7136,N_7196);
and U7216 (N_7216,N_7155,N_7183);
or U7217 (N_7217,N_7170,N_7116);
xor U7218 (N_7218,N_7171,N_7191);
and U7219 (N_7219,N_7123,N_7128);
nor U7220 (N_7220,N_7121,N_7193);
nand U7221 (N_7221,N_7157,N_7105);
xnor U7222 (N_7222,N_7142,N_7197);
nor U7223 (N_7223,N_7175,N_7178);
nor U7224 (N_7224,N_7186,N_7152);
or U7225 (N_7225,N_7146,N_7103);
nor U7226 (N_7226,N_7188,N_7154);
nor U7227 (N_7227,N_7190,N_7187);
or U7228 (N_7228,N_7182,N_7125);
nor U7229 (N_7229,N_7169,N_7122);
nand U7230 (N_7230,N_7129,N_7132);
nand U7231 (N_7231,N_7174,N_7114);
xor U7232 (N_7232,N_7173,N_7195);
and U7233 (N_7233,N_7111,N_7180);
or U7234 (N_7234,N_7107,N_7130);
or U7235 (N_7235,N_7140,N_7138);
and U7236 (N_7236,N_7147,N_7131);
nor U7237 (N_7237,N_7145,N_7168);
and U7238 (N_7238,N_7120,N_7198);
and U7239 (N_7239,N_7192,N_7185);
nand U7240 (N_7240,N_7165,N_7148);
or U7241 (N_7241,N_7109,N_7106);
nand U7242 (N_7242,N_7149,N_7150);
or U7243 (N_7243,N_7124,N_7177);
nand U7244 (N_7244,N_7156,N_7135);
nor U7245 (N_7245,N_7166,N_7194);
xnor U7246 (N_7246,N_7101,N_7163);
xnor U7247 (N_7247,N_7127,N_7172);
nand U7248 (N_7248,N_7133,N_7159);
and U7249 (N_7249,N_7161,N_7199);
xor U7250 (N_7250,N_7112,N_7186);
or U7251 (N_7251,N_7136,N_7121);
or U7252 (N_7252,N_7107,N_7124);
xor U7253 (N_7253,N_7145,N_7118);
nand U7254 (N_7254,N_7100,N_7173);
nor U7255 (N_7255,N_7184,N_7116);
nor U7256 (N_7256,N_7177,N_7132);
nand U7257 (N_7257,N_7195,N_7119);
and U7258 (N_7258,N_7132,N_7122);
nor U7259 (N_7259,N_7144,N_7161);
nand U7260 (N_7260,N_7187,N_7149);
and U7261 (N_7261,N_7148,N_7178);
xor U7262 (N_7262,N_7113,N_7154);
and U7263 (N_7263,N_7108,N_7178);
nor U7264 (N_7264,N_7175,N_7191);
or U7265 (N_7265,N_7123,N_7168);
or U7266 (N_7266,N_7127,N_7119);
xor U7267 (N_7267,N_7179,N_7127);
nor U7268 (N_7268,N_7170,N_7151);
or U7269 (N_7269,N_7125,N_7176);
nand U7270 (N_7270,N_7134,N_7185);
or U7271 (N_7271,N_7121,N_7131);
and U7272 (N_7272,N_7159,N_7162);
or U7273 (N_7273,N_7128,N_7129);
nor U7274 (N_7274,N_7199,N_7198);
and U7275 (N_7275,N_7108,N_7126);
xor U7276 (N_7276,N_7140,N_7168);
nor U7277 (N_7277,N_7185,N_7169);
xnor U7278 (N_7278,N_7143,N_7115);
nor U7279 (N_7279,N_7116,N_7190);
and U7280 (N_7280,N_7138,N_7181);
nand U7281 (N_7281,N_7184,N_7180);
and U7282 (N_7282,N_7161,N_7166);
or U7283 (N_7283,N_7106,N_7189);
and U7284 (N_7284,N_7107,N_7190);
or U7285 (N_7285,N_7172,N_7156);
nand U7286 (N_7286,N_7186,N_7157);
and U7287 (N_7287,N_7196,N_7160);
nand U7288 (N_7288,N_7198,N_7181);
nor U7289 (N_7289,N_7141,N_7170);
nand U7290 (N_7290,N_7142,N_7144);
or U7291 (N_7291,N_7143,N_7135);
or U7292 (N_7292,N_7183,N_7136);
and U7293 (N_7293,N_7125,N_7156);
and U7294 (N_7294,N_7133,N_7125);
and U7295 (N_7295,N_7135,N_7146);
and U7296 (N_7296,N_7177,N_7155);
nand U7297 (N_7297,N_7155,N_7187);
xnor U7298 (N_7298,N_7158,N_7197);
or U7299 (N_7299,N_7193,N_7155);
nand U7300 (N_7300,N_7219,N_7271);
nand U7301 (N_7301,N_7226,N_7206);
and U7302 (N_7302,N_7218,N_7205);
nand U7303 (N_7303,N_7284,N_7279);
xor U7304 (N_7304,N_7277,N_7222);
nor U7305 (N_7305,N_7262,N_7253);
nor U7306 (N_7306,N_7290,N_7227);
or U7307 (N_7307,N_7255,N_7223);
nor U7308 (N_7308,N_7274,N_7268);
nand U7309 (N_7309,N_7294,N_7202);
nor U7310 (N_7310,N_7269,N_7288);
and U7311 (N_7311,N_7237,N_7282);
nand U7312 (N_7312,N_7280,N_7215);
nor U7313 (N_7313,N_7258,N_7272);
nor U7314 (N_7314,N_7221,N_7281);
and U7315 (N_7315,N_7298,N_7213);
and U7316 (N_7316,N_7217,N_7263);
or U7317 (N_7317,N_7239,N_7278);
xnor U7318 (N_7318,N_7216,N_7295);
or U7319 (N_7319,N_7211,N_7233);
xor U7320 (N_7320,N_7275,N_7209);
nand U7321 (N_7321,N_7273,N_7260);
and U7322 (N_7322,N_7292,N_7235);
nor U7323 (N_7323,N_7203,N_7244);
or U7324 (N_7324,N_7240,N_7250);
xor U7325 (N_7325,N_7204,N_7289);
nor U7326 (N_7326,N_7236,N_7224);
nand U7327 (N_7327,N_7212,N_7231);
xnor U7328 (N_7328,N_7259,N_7200);
and U7329 (N_7329,N_7287,N_7229);
xor U7330 (N_7330,N_7241,N_7248);
xor U7331 (N_7331,N_7220,N_7297);
xor U7332 (N_7332,N_7251,N_7232);
and U7333 (N_7333,N_7245,N_7299);
and U7334 (N_7334,N_7270,N_7208);
xnor U7335 (N_7335,N_7265,N_7252);
nor U7336 (N_7336,N_7254,N_7201);
and U7337 (N_7337,N_7261,N_7210);
nand U7338 (N_7338,N_7286,N_7246);
nor U7339 (N_7339,N_7243,N_7207);
or U7340 (N_7340,N_7249,N_7256);
nand U7341 (N_7341,N_7234,N_7264);
or U7342 (N_7342,N_7238,N_7228);
nor U7343 (N_7343,N_7266,N_7285);
xnor U7344 (N_7344,N_7296,N_7230);
nand U7345 (N_7345,N_7283,N_7293);
nand U7346 (N_7346,N_7267,N_7214);
xor U7347 (N_7347,N_7276,N_7247);
xnor U7348 (N_7348,N_7291,N_7225);
or U7349 (N_7349,N_7257,N_7242);
and U7350 (N_7350,N_7257,N_7282);
nor U7351 (N_7351,N_7283,N_7270);
nand U7352 (N_7352,N_7231,N_7274);
nor U7353 (N_7353,N_7247,N_7294);
or U7354 (N_7354,N_7265,N_7220);
and U7355 (N_7355,N_7263,N_7292);
xnor U7356 (N_7356,N_7220,N_7249);
or U7357 (N_7357,N_7201,N_7297);
and U7358 (N_7358,N_7231,N_7207);
xor U7359 (N_7359,N_7281,N_7298);
xor U7360 (N_7360,N_7269,N_7230);
or U7361 (N_7361,N_7241,N_7268);
or U7362 (N_7362,N_7250,N_7284);
nand U7363 (N_7363,N_7233,N_7238);
xor U7364 (N_7364,N_7296,N_7274);
xor U7365 (N_7365,N_7247,N_7233);
nor U7366 (N_7366,N_7269,N_7257);
nand U7367 (N_7367,N_7266,N_7251);
xor U7368 (N_7368,N_7293,N_7210);
and U7369 (N_7369,N_7219,N_7215);
xor U7370 (N_7370,N_7206,N_7247);
or U7371 (N_7371,N_7232,N_7213);
xnor U7372 (N_7372,N_7291,N_7283);
nor U7373 (N_7373,N_7265,N_7231);
and U7374 (N_7374,N_7253,N_7241);
or U7375 (N_7375,N_7298,N_7244);
nand U7376 (N_7376,N_7264,N_7219);
and U7377 (N_7377,N_7280,N_7229);
or U7378 (N_7378,N_7285,N_7201);
or U7379 (N_7379,N_7217,N_7258);
xor U7380 (N_7380,N_7279,N_7268);
nand U7381 (N_7381,N_7222,N_7279);
nand U7382 (N_7382,N_7223,N_7219);
and U7383 (N_7383,N_7275,N_7234);
or U7384 (N_7384,N_7211,N_7253);
or U7385 (N_7385,N_7248,N_7278);
or U7386 (N_7386,N_7274,N_7222);
or U7387 (N_7387,N_7260,N_7266);
and U7388 (N_7388,N_7285,N_7241);
or U7389 (N_7389,N_7210,N_7262);
xnor U7390 (N_7390,N_7288,N_7260);
and U7391 (N_7391,N_7259,N_7229);
xnor U7392 (N_7392,N_7296,N_7275);
xor U7393 (N_7393,N_7233,N_7214);
nor U7394 (N_7394,N_7266,N_7292);
xnor U7395 (N_7395,N_7228,N_7292);
xnor U7396 (N_7396,N_7256,N_7218);
nand U7397 (N_7397,N_7280,N_7242);
or U7398 (N_7398,N_7235,N_7201);
nand U7399 (N_7399,N_7298,N_7271);
nor U7400 (N_7400,N_7366,N_7339);
xor U7401 (N_7401,N_7333,N_7304);
nor U7402 (N_7402,N_7313,N_7377);
and U7403 (N_7403,N_7396,N_7381);
nor U7404 (N_7404,N_7318,N_7370);
nand U7405 (N_7405,N_7358,N_7390);
xor U7406 (N_7406,N_7306,N_7322);
nand U7407 (N_7407,N_7320,N_7331);
nand U7408 (N_7408,N_7392,N_7338);
or U7409 (N_7409,N_7316,N_7343);
and U7410 (N_7410,N_7372,N_7336);
or U7411 (N_7411,N_7386,N_7352);
nand U7412 (N_7412,N_7341,N_7382);
nor U7413 (N_7413,N_7310,N_7345);
xnor U7414 (N_7414,N_7354,N_7362);
nor U7415 (N_7415,N_7367,N_7347);
nor U7416 (N_7416,N_7394,N_7359);
and U7417 (N_7417,N_7303,N_7335);
nor U7418 (N_7418,N_7348,N_7369);
xnor U7419 (N_7419,N_7324,N_7334);
xnor U7420 (N_7420,N_7393,N_7328);
and U7421 (N_7421,N_7388,N_7317);
or U7422 (N_7422,N_7340,N_7344);
and U7423 (N_7423,N_7351,N_7361);
or U7424 (N_7424,N_7389,N_7379);
xor U7425 (N_7425,N_7374,N_7373);
xnor U7426 (N_7426,N_7307,N_7342);
nand U7427 (N_7427,N_7346,N_7380);
and U7428 (N_7428,N_7327,N_7395);
and U7429 (N_7429,N_7326,N_7385);
nand U7430 (N_7430,N_7378,N_7319);
nand U7431 (N_7431,N_7364,N_7365);
xnor U7432 (N_7432,N_7355,N_7350);
and U7433 (N_7433,N_7363,N_7399);
or U7434 (N_7434,N_7309,N_7371);
xnor U7435 (N_7435,N_7301,N_7360);
nand U7436 (N_7436,N_7315,N_7376);
nor U7437 (N_7437,N_7311,N_7356);
and U7438 (N_7438,N_7375,N_7325);
xnor U7439 (N_7439,N_7332,N_7368);
nor U7440 (N_7440,N_7323,N_7357);
or U7441 (N_7441,N_7308,N_7383);
or U7442 (N_7442,N_7330,N_7397);
or U7443 (N_7443,N_7349,N_7387);
nor U7444 (N_7444,N_7305,N_7300);
xor U7445 (N_7445,N_7321,N_7312);
xor U7446 (N_7446,N_7391,N_7353);
nand U7447 (N_7447,N_7398,N_7329);
and U7448 (N_7448,N_7337,N_7302);
nand U7449 (N_7449,N_7314,N_7384);
and U7450 (N_7450,N_7361,N_7372);
nand U7451 (N_7451,N_7359,N_7364);
xnor U7452 (N_7452,N_7347,N_7313);
and U7453 (N_7453,N_7356,N_7362);
nor U7454 (N_7454,N_7311,N_7300);
nor U7455 (N_7455,N_7398,N_7396);
and U7456 (N_7456,N_7312,N_7322);
nor U7457 (N_7457,N_7337,N_7386);
xor U7458 (N_7458,N_7333,N_7359);
nand U7459 (N_7459,N_7378,N_7307);
nor U7460 (N_7460,N_7362,N_7348);
or U7461 (N_7461,N_7318,N_7333);
or U7462 (N_7462,N_7310,N_7329);
nand U7463 (N_7463,N_7343,N_7340);
or U7464 (N_7464,N_7360,N_7391);
and U7465 (N_7465,N_7357,N_7334);
nand U7466 (N_7466,N_7358,N_7397);
and U7467 (N_7467,N_7391,N_7380);
or U7468 (N_7468,N_7384,N_7309);
and U7469 (N_7469,N_7367,N_7380);
or U7470 (N_7470,N_7366,N_7399);
or U7471 (N_7471,N_7367,N_7350);
nor U7472 (N_7472,N_7393,N_7326);
and U7473 (N_7473,N_7302,N_7356);
nand U7474 (N_7474,N_7323,N_7382);
nor U7475 (N_7475,N_7319,N_7387);
and U7476 (N_7476,N_7320,N_7387);
nand U7477 (N_7477,N_7374,N_7376);
and U7478 (N_7478,N_7375,N_7309);
xnor U7479 (N_7479,N_7378,N_7368);
or U7480 (N_7480,N_7381,N_7336);
xnor U7481 (N_7481,N_7387,N_7331);
xor U7482 (N_7482,N_7300,N_7391);
or U7483 (N_7483,N_7383,N_7300);
or U7484 (N_7484,N_7374,N_7356);
nor U7485 (N_7485,N_7378,N_7336);
or U7486 (N_7486,N_7378,N_7345);
or U7487 (N_7487,N_7325,N_7382);
nor U7488 (N_7488,N_7314,N_7309);
or U7489 (N_7489,N_7301,N_7389);
nand U7490 (N_7490,N_7334,N_7351);
or U7491 (N_7491,N_7332,N_7356);
nor U7492 (N_7492,N_7334,N_7396);
or U7493 (N_7493,N_7339,N_7348);
nand U7494 (N_7494,N_7314,N_7324);
xnor U7495 (N_7495,N_7366,N_7383);
nand U7496 (N_7496,N_7300,N_7385);
and U7497 (N_7497,N_7365,N_7307);
and U7498 (N_7498,N_7352,N_7321);
and U7499 (N_7499,N_7397,N_7370);
nand U7500 (N_7500,N_7486,N_7425);
or U7501 (N_7501,N_7497,N_7495);
xor U7502 (N_7502,N_7448,N_7418);
nor U7503 (N_7503,N_7403,N_7462);
and U7504 (N_7504,N_7421,N_7400);
nand U7505 (N_7505,N_7447,N_7423);
nor U7506 (N_7506,N_7455,N_7489);
or U7507 (N_7507,N_7444,N_7463);
nor U7508 (N_7508,N_7493,N_7433);
and U7509 (N_7509,N_7458,N_7443);
xor U7510 (N_7510,N_7450,N_7454);
and U7511 (N_7511,N_7404,N_7446);
and U7512 (N_7512,N_7496,N_7402);
and U7513 (N_7513,N_7456,N_7451);
nand U7514 (N_7514,N_7499,N_7436);
and U7515 (N_7515,N_7409,N_7498);
and U7516 (N_7516,N_7437,N_7467);
nand U7517 (N_7517,N_7466,N_7474);
or U7518 (N_7518,N_7420,N_7483);
nand U7519 (N_7519,N_7413,N_7439);
nor U7520 (N_7520,N_7432,N_7430);
or U7521 (N_7521,N_7482,N_7410);
xnor U7522 (N_7522,N_7469,N_7484);
xnor U7523 (N_7523,N_7475,N_7416);
nand U7524 (N_7524,N_7494,N_7487);
xnor U7525 (N_7525,N_7401,N_7480);
and U7526 (N_7526,N_7434,N_7492);
nor U7527 (N_7527,N_7424,N_7461);
nand U7528 (N_7528,N_7471,N_7460);
or U7529 (N_7529,N_7431,N_7473);
nor U7530 (N_7530,N_7453,N_7427);
nand U7531 (N_7531,N_7452,N_7414);
nand U7532 (N_7532,N_7411,N_7457);
or U7533 (N_7533,N_7415,N_7490);
or U7534 (N_7534,N_7445,N_7472);
nor U7535 (N_7535,N_7479,N_7441);
nor U7536 (N_7536,N_7426,N_7459);
nor U7537 (N_7537,N_7449,N_7405);
and U7538 (N_7538,N_7477,N_7429);
nor U7539 (N_7539,N_7417,N_7491);
or U7540 (N_7540,N_7442,N_7407);
xnor U7541 (N_7541,N_7435,N_7481);
xnor U7542 (N_7542,N_7465,N_7438);
xnor U7543 (N_7543,N_7422,N_7488);
and U7544 (N_7544,N_7408,N_7428);
xnor U7545 (N_7545,N_7468,N_7406);
xnor U7546 (N_7546,N_7440,N_7470);
nand U7547 (N_7547,N_7412,N_7485);
and U7548 (N_7548,N_7478,N_7476);
nand U7549 (N_7549,N_7464,N_7419);
nor U7550 (N_7550,N_7462,N_7485);
nor U7551 (N_7551,N_7443,N_7466);
nor U7552 (N_7552,N_7455,N_7481);
xor U7553 (N_7553,N_7474,N_7480);
or U7554 (N_7554,N_7469,N_7406);
nand U7555 (N_7555,N_7480,N_7417);
nor U7556 (N_7556,N_7479,N_7463);
nor U7557 (N_7557,N_7471,N_7485);
nand U7558 (N_7558,N_7438,N_7478);
or U7559 (N_7559,N_7428,N_7400);
nor U7560 (N_7560,N_7447,N_7421);
or U7561 (N_7561,N_7440,N_7441);
xnor U7562 (N_7562,N_7487,N_7462);
or U7563 (N_7563,N_7452,N_7437);
nand U7564 (N_7564,N_7455,N_7466);
nand U7565 (N_7565,N_7452,N_7419);
or U7566 (N_7566,N_7422,N_7408);
xnor U7567 (N_7567,N_7487,N_7457);
nand U7568 (N_7568,N_7493,N_7445);
nor U7569 (N_7569,N_7450,N_7437);
nand U7570 (N_7570,N_7448,N_7478);
and U7571 (N_7571,N_7422,N_7433);
xor U7572 (N_7572,N_7489,N_7473);
nand U7573 (N_7573,N_7456,N_7449);
nor U7574 (N_7574,N_7455,N_7479);
nand U7575 (N_7575,N_7455,N_7411);
and U7576 (N_7576,N_7498,N_7434);
nor U7577 (N_7577,N_7455,N_7442);
or U7578 (N_7578,N_7440,N_7484);
xor U7579 (N_7579,N_7480,N_7436);
nand U7580 (N_7580,N_7406,N_7476);
nor U7581 (N_7581,N_7453,N_7406);
and U7582 (N_7582,N_7461,N_7495);
and U7583 (N_7583,N_7454,N_7460);
or U7584 (N_7584,N_7458,N_7479);
nand U7585 (N_7585,N_7495,N_7401);
nor U7586 (N_7586,N_7471,N_7430);
xor U7587 (N_7587,N_7403,N_7449);
nor U7588 (N_7588,N_7479,N_7469);
nor U7589 (N_7589,N_7454,N_7438);
and U7590 (N_7590,N_7499,N_7418);
nand U7591 (N_7591,N_7492,N_7491);
nand U7592 (N_7592,N_7444,N_7439);
or U7593 (N_7593,N_7483,N_7499);
and U7594 (N_7594,N_7494,N_7499);
or U7595 (N_7595,N_7468,N_7444);
or U7596 (N_7596,N_7469,N_7451);
nor U7597 (N_7597,N_7419,N_7497);
or U7598 (N_7598,N_7465,N_7499);
or U7599 (N_7599,N_7429,N_7410);
and U7600 (N_7600,N_7587,N_7565);
xor U7601 (N_7601,N_7537,N_7571);
nor U7602 (N_7602,N_7590,N_7533);
or U7603 (N_7603,N_7597,N_7592);
nor U7604 (N_7604,N_7575,N_7521);
or U7605 (N_7605,N_7545,N_7531);
nand U7606 (N_7606,N_7555,N_7568);
nor U7607 (N_7607,N_7596,N_7548);
xor U7608 (N_7608,N_7525,N_7543);
or U7609 (N_7609,N_7570,N_7559);
and U7610 (N_7610,N_7557,N_7578);
nor U7611 (N_7611,N_7551,N_7562);
nor U7612 (N_7612,N_7519,N_7529);
nor U7613 (N_7613,N_7561,N_7509);
nor U7614 (N_7614,N_7591,N_7532);
and U7615 (N_7615,N_7573,N_7508);
and U7616 (N_7616,N_7583,N_7540);
xor U7617 (N_7617,N_7515,N_7550);
or U7618 (N_7618,N_7585,N_7511);
or U7619 (N_7619,N_7502,N_7546);
or U7620 (N_7620,N_7520,N_7514);
and U7621 (N_7621,N_7541,N_7505);
nand U7622 (N_7622,N_7589,N_7598);
and U7623 (N_7623,N_7588,N_7593);
or U7624 (N_7624,N_7535,N_7563);
nand U7625 (N_7625,N_7594,N_7524);
and U7626 (N_7626,N_7558,N_7544);
nor U7627 (N_7627,N_7518,N_7526);
nand U7628 (N_7628,N_7523,N_7516);
xnor U7629 (N_7629,N_7534,N_7504);
and U7630 (N_7630,N_7599,N_7507);
nor U7631 (N_7631,N_7510,N_7595);
nand U7632 (N_7632,N_7552,N_7527);
nor U7633 (N_7633,N_7564,N_7503);
or U7634 (N_7634,N_7528,N_7567);
and U7635 (N_7635,N_7549,N_7556);
xnor U7636 (N_7636,N_7569,N_7500);
xor U7637 (N_7637,N_7560,N_7566);
nand U7638 (N_7638,N_7553,N_7522);
nor U7639 (N_7639,N_7547,N_7582);
or U7640 (N_7640,N_7580,N_7512);
or U7641 (N_7641,N_7579,N_7584);
or U7642 (N_7642,N_7542,N_7506);
and U7643 (N_7643,N_7501,N_7554);
nor U7644 (N_7644,N_7574,N_7536);
nor U7645 (N_7645,N_7517,N_7513);
and U7646 (N_7646,N_7581,N_7530);
nor U7647 (N_7647,N_7586,N_7539);
nor U7648 (N_7648,N_7572,N_7576);
xnor U7649 (N_7649,N_7577,N_7538);
or U7650 (N_7650,N_7542,N_7558);
and U7651 (N_7651,N_7563,N_7547);
nand U7652 (N_7652,N_7589,N_7548);
nand U7653 (N_7653,N_7592,N_7560);
nor U7654 (N_7654,N_7512,N_7590);
nand U7655 (N_7655,N_7562,N_7594);
or U7656 (N_7656,N_7535,N_7558);
nand U7657 (N_7657,N_7551,N_7539);
xnor U7658 (N_7658,N_7518,N_7557);
xor U7659 (N_7659,N_7542,N_7574);
or U7660 (N_7660,N_7548,N_7508);
nand U7661 (N_7661,N_7566,N_7522);
nor U7662 (N_7662,N_7505,N_7576);
xor U7663 (N_7663,N_7512,N_7502);
nor U7664 (N_7664,N_7541,N_7549);
or U7665 (N_7665,N_7578,N_7583);
nand U7666 (N_7666,N_7535,N_7537);
nand U7667 (N_7667,N_7551,N_7513);
xor U7668 (N_7668,N_7597,N_7563);
and U7669 (N_7669,N_7538,N_7563);
nor U7670 (N_7670,N_7580,N_7516);
xor U7671 (N_7671,N_7520,N_7589);
or U7672 (N_7672,N_7594,N_7511);
or U7673 (N_7673,N_7568,N_7530);
and U7674 (N_7674,N_7517,N_7554);
xor U7675 (N_7675,N_7556,N_7501);
xnor U7676 (N_7676,N_7547,N_7562);
nor U7677 (N_7677,N_7531,N_7513);
xor U7678 (N_7678,N_7561,N_7518);
nor U7679 (N_7679,N_7563,N_7545);
and U7680 (N_7680,N_7508,N_7581);
nand U7681 (N_7681,N_7501,N_7558);
or U7682 (N_7682,N_7543,N_7509);
and U7683 (N_7683,N_7573,N_7572);
nor U7684 (N_7684,N_7533,N_7571);
nor U7685 (N_7685,N_7514,N_7572);
nand U7686 (N_7686,N_7581,N_7599);
and U7687 (N_7687,N_7519,N_7595);
nand U7688 (N_7688,N_7594,N_7592);
or U7689 (N_7689,N_7565,N_7566);
or U7690 (N_7690,N_7521,N_7565);
or U7691 (N_7691,N_7515,N_7577);
xnor U7692 (N_7692,N_7580,N_7549);
nand U7693 (N_7693,N_7585,N_7527);
nor U7694 (N_7694,N_7546,N_7563);
xor U7695 (N_7695,N_7537,N_7534);
xnor U7696 (N_7696,N_7501,N_7583);
nor U7697 (N_7697,N_7557,N_7594);
and U7698 (N_7698,N_7551,N_7556);
nor U7699 (N_7699,N_7589,N_7572);
and U7700 (N_7700,N_7611,N_7638);
and U7701 (N_7701,N_7631,N_7607);
or U7702 (N_7702,N_7699,N_7616);
or U7703 (N_7703,N_7680,N_7670);
nor U7704 (N_7704,N_7664,N_7612);
nor U7705 (N_7705,N_7698,N_7665);
nor U7706 (N_7706,N_7621,N_7656);
nor U7707 (N_7707,N_7624,N_7660);
nor U7708 (N_7708,N_7625,N_7618);
xnor U7709 (N_7709,N_7609,N_7667);
and U7710 (N_7710,N_7688,N_7692);
nor U7711 (N_7711,N_7654,N_7641);
xor U7712 (N_7712,N_7623,N_7682);
and U7713 (N_7713,N_7633,N_7666);
and U7714 (N_7714,N_7683,N_7635);
or U7715 (N_7715,N_7658,N_7672);
or U7716 (N_7716,N_7649,N_7678);
or U7717 (N_7717,N_7668,N_7684);
or U7718 (N_7718,N_7690,N_7691);
and U7719 (N_7719,N_7622,N_7663);
nand U7720 (N_7720,N_7669,N_7655);
nor U7721 (N_7721,N_7613,N_7687);
xnor U7722 (N_7722,N_7608,N_7640);
and U7723 (N_7723,N_7643,N_7662);
nand U7724 (N_7724,N_7628,N_7610);
and U7725 (N_7725,N_7601,N_7671);
nand U7726 (N_7726,N_7606,N_7626);
and U7727 (N_7727,N_7652,N_7629);
or U7728 (N_7728,N_7604,N_7644);
and U7729 (N_7729,N_7632,N_7645);
nor U7730 (N_7730,N_7657,N_7651);
nand U7731 (N_7731,N_7639,N_7603);
nor U7732 (N_7732,N_7695,N_7634);
or U7733 (N_7733,N_7673,N_7681);
or U7734 (N_7734,N_7602,N_7677);
or U7735 (N_7735,N_7685,N_7679);
nand U7736 (N_7736,N_7676,N_7646);
nand U7737 (N_7737,N_7600,N_7615);
nand U7738 (N_7738,N_7619,N_7648);
xor U7739 (N_7739,N_7694,N_7630);
nand U7740 (N_7740,N_7647,N_7627);
nand U7741 (N_7741,N_7650,N_7620);
or U7742 (N_7742,N_7617,N_7653);
and U7743 (N_7743,N_7661,N_7659);
and U7744 (N_7744,N_7689,N_7696);
nand U7745 (N_7745,N_7637,N_7697);
nor U7746 (N_7746,N_7636,N_7686);
or U7747 (N_7747,N_7642,N_7674);
nand U7748 (N_7748,N_7675,N_7605);
and U7749 (N_7749,N_7693,N_7614);
nand U7750 (N_7750,N_7695,N_7612);
or U7751 (N_7751,N_7613,N_7610);
nand U7752 (N_7752,N_7665,N_7642);
nand U7753 (N_7753,N_7645,N_7612);
nor U7754 (N_7754,N_7656,N_7605);
and U7755 (N_7755,N_7658,N_7691);
nor U7756 (N_7756,N_7601,N_7616);
nor U7757 (N_7757,N_7693,N_7665);
xor U7758 (N_7758,N_7628,N_7663);
xor U7759 (N_7759,N_7640,N_7650);
nor U7760 (N_7760,N_7617,N_7698);
or U7761 (N_7761,N_7673,N_7621);
xnor U7762 (N_7762,N_7676,N_7674);
nor U7763 (N_7763,N_7638,N_7647);
xor U7764 (N_7764,N_7683,N_7626);
and U7765 (N_7765,N_7657,N_7626);
nor U7766 (N_7766,N_7601,N_7648);
nor U7767 (N_7767,N_7604,N_7666);
xor U7768 (N_7768,N_7640,N_7642);
and U7769 (N_7769,N_7695,N_7646);
nand U7770 (N_7770,N_7663,N_7602);
xor U7771 (N_7771,N_7697,N_7640);
xnor U7772 (N_7772,N_7642,N_7604);
nand U7773 (N_7773,N_7615,N_7659);
nor U7774 (N_7774,N_7601,N_7664);
nand U7775 (N_7775,N_7608,N_7615);
xor U7776 (N_7776,N_7647,N_7624);
or U7777 (N_7777,N_7636,N_7684);
and U7778 (N_7778,N_7647,N_7674);
and U7779 (N_7779,N_7604,N_7657);
xnor U7780 (N_7780,N_7626,N_7640);
nor U7781 (N_7781,N_7610,N_7671);
and U7782 (N_7782,N_7615,N_7618);
or U7783 (N_7783,N_7651,N_7656);
nand U7784 (N_7784,N_7690,N_7689);
and U7785 (N_7785,N_7660,N_7621);
and U7786 (N_7786,N_7688,N_7633);
nand U7787 (N_7787,N_7641,N_7672);
or U7788 (N_7788,N_7671,N_7651);
nand U7789 (N_7789,N_7616,N_7632);
and U7790 (N_7790,N_7625,N_7612);
xor U7791 (N_7791,N_7624,N_7663);
and U7792 (N_7792,N_7675,N_7626);
and U7793 (N_7793,N_7606,N_7693);
nand U7794 (N_7794,N_7664,N_7639);
nor U7795 (N_7795,N_7650,N_7606);
nor U7796 (N_7796,N_7672,N_7673);
nand U7797 (N_7797,N_7622,N_7605);
nand U7798 (N_7798,N_7699,N_7614);
xor U7799 (N_7799,N_7604,N_7627);
nor U7800 (N_7800,N_7784,N_7772);
xor U7801 (N_7801,N_7751,N_7741);
xor U7802 (N_7802,N_7747,N_7738);
nand U7803 (N_7803,N_7718,N_7771);
nor U7804 (N_7804,N_7742,N_7703);
xnor U7805 (N_7805,N_7743,N_7752);
and U7806 (N_7806,N_7734,N_7728);
and U7807 (N_7807,N_7786,N_7705);
xnor U7808 (N_7808,N_7704,N_7744);
and U7809 (N_7809,N_7735,N_7711);
nor U7810 (N_7810,N_7702,N_7774);
nand U7811 (N_7811,N_7783,N_7789);
or U7812 (N_7812,N_7730,N_7756);
xnor U7813 (N_7813,N_7709,N_7717);
nand U7814 (N_7814,N_7732,N_7722);
nor U7815 (N_7815,N_7733,N_7746);
xnor U7816 (N_7816,N_7765,N_7712);
and U7817 (N_7817,N_7768,N_7788);
or U7818 (N_7818,N_7764,N_7782);
xor U7819 (N_7819,N_7713,N_7787);
nor U7820 (N_7820,N_7769,N_7716);
and U7821 (N_7821,N_7737,N_7758);
nand U7822 (N_7822,N_7727,N_7721);
or U7823 (N_7823,N_7798,N_7777);
nand U7824 (N_7824,N_7729,N_7757);
nand U7825 (N_7825,N_7770,N_7766);
nor U7826 (N_7826,N_7739,N_7773);
nand U7827 (N_7827,N_7749,N_7720);
and U7828 (N_7828,N_7759,N_7776);
nor U7829 (N_7829,N_7700,N_7715);
or U7830 (N_7830,N_7799,N_7785);
nor U7831 (N_7831,N_7791,N_7707);
xnor U7832 (N_7832,N_7714,N_7794);
or U7833 (N_7833,N_7706,N_7792);
xor U7834 (N_7834,N_7779,N_7719);
or U7835 (N_7835,N_7753,N_7761);
and U7836 (N_7836,N_7796,N_7778);
nand U7837 (N_7837,N_7795,N_7781);
nand U7838 (N_7838,N_7763,N_7726);
nand U7839 (N_7839,N_7723,N_7760);
nor U7840 (N_7840,N_7780,N_7775);
xnor U7841 (N_7841,N_7736,N_7797);
or U7842 (N_7842,N_7748,N_7745);
or U7843 (N_7843,N_7731,N_7701);
nor U7844 (N_7844,N_7767,N_7754);
and U7845 (N_7845,N_7750,N_7740);
nand U7846 (N_7846,N_7755,N_7724);
nand U7847 (N_7847,N_7762,N_7793);
nand U7848 (N_7848,N_7710,N_7708);
nor U7849 (N_7849,N_7790,N_7725);
or U7850 (N_7850,N_7783,N_7732);
nor U7851 (N_7851,N_7793,N_7742);
xnor U7852 (N_7852,N_7739,N_7788);
or U7853 (N_7853,N_7736,N_7739);
nand U7854 (N_7854,N_7762,N_7701);
and U7855 (N_7855,N_7767,N_7707);
and U7856 (N_7856,N_7739,N_7767);
nor U7857 (N_7857,N_7744,N_7739);
nand U7858 (N_7858,N_7773,N_7771);
and U7859 (N_7859,N_7773,N_7756);
xor U7860 (N_7860,N_7757,N_7799);
or U7861 (N_7861,N_7714,N_7736);
nand U7862 (N_7862,N_7762,N_7771);
xnor U7863 (N_7863,N_7706,N_7784);
and U7864 (N_7864,N_7734,N_7725);
and U7865 (N_7865,N_7714,N_7767);
and U7866 (N_7866,N_7725,N_7736);
nor U7867 (N_7867,N_7730,N_7736);
xnor U7868 (N_7868,N_7747,N_7784);
xnor U7869 (N_7869,N_7754,N_7722);
and U7870 (N_7870,N_7767,N_7725);
nor U7871 (N_7871,N_7763,N_7718);
and U7872 (N_7872,N_7747,N_7755);
or U7873 (N_7873,N_7794,N_7757);
and U7874 (N_7874,N_7784,N_7755);
xor U7875 (N_7875,N_7777,N_7705);
and U7876 (N_7876,N_7716,N_7784);
or U7877 (N_7877,N_7734,N_7764);
and U7878 (N_7878,N_7746,N_7738);
nand U7879 (N_7879,N_7778,N_7761);
xnor U7880 (N_7880,N_7778,N_7709);
and U7881 (N_7881,N_7770,N_7717);
and U7882 (N_7882,N_7732,N_7757);
or U7883 (N_7883,N_7714,N_7704);
xnor U7884 (N_7884,N_7725,N_7759);
and U7885 (N_7885,N_7770,N_7798);
and U7886 (N_7886,N_7776,N_7774);
xnor U7887 (N_7887,N_7763,N_7793);
and U7888 (N_7888,N_7751,N_7777);
and U7889 (N_7889,N_7775,N_7796);
xnor U7890 (N_7890,N_7783,N_7763);
xnor U7891 (N_7891,N_7767,N_7780);
nor U7892 (N_7892,N_7741,N_7720);
and U7893 (N_7893,N_7743,N_7734);
nor U7894 (N_7894,N_7748,N_7776);
nand U7895 (N_7895,N_7736,N_7712);
nand U7896 (N_7896,N_7758,N_7757);
xor U7897 (N_7897,N_7742,N_7725);
nor U7898 (N_7898,N_7707,N_7739);
nand U7899 (N_7899,N_7733,N_7798);
nand U7900 (N_7900,N_7827,N_7871);
nor U7901 (N_7901,N_7860,N_7876);
xnor U7902 (N_7902,N_7821,N_7862);
nand U7903 (N_7903,N_7885,N_7837);
and U7904 (N_7904,N_7823,N_7896);
and U7905 (N_7905,N_7810,N_7845);
nor U7906 (N_7906,N_7864,N_7802);
xnor U7907 (N_7907,N_7804,N_7883);
nor U7908 (N_7908,N_7859,N_7879);
nand U7909 (N_7909,N_7872,N_7809);
nor U7910 (N_7910,N_7881,N_7882);
or U7911 (N_7911,N_7824,N_7841);
and U7912 (N_7912,N_7816,N_7892);
and U7913 (N_7913,N_7858,N_7898);
nor U7914 (N_7914,N_7806,N_7866);
nand U7915 (N_7915,N_7843,N_7829);
or U7916 (N_7916,N_7884,N_7831);
nand U7917 (N_7917,N_7851,N_7855);
xor U7918 (N_7918,N_7826,N_7875);
xor U7919 (N_7919,N_7853,N_7814);
xnor U7920 (N_7920,N_7847,N_7800);
xnor U7921 (N_7921,N_7852,N_7886);
nand U7922 (N_7922,N_7870,N_7897);
nand U7923 (N_7923,N_7840,N_7891);
xnor U7924 (N_7924,N_7839,N_7880);
and U7925 (N_7925,N_7873,N_7822);
xor U7926 (N_7926,N_7893,N_7894);
nand U7927 (N_7927,N_7819,N_7857);
or U7928 (N_7928,N_7895,N_7812);
and U7929 (N_7929,N_7867,N_7801);
or U7930 (N_7930,N_7878,N_7854);
or U7931 (N_7931,N_7846,N_7869);
nor U7932 (N_7932,N_7817,N_7818);
nand U7933 (N_7933,N_7820,N_7856);
nand U7934 (N_7934,N_7861,N_7833);
or U7935 (N_7935,N_7890,N_7805);
and U7936 (N_7936,N_7844,N_7848);
xor U7937 (N_7937,N_7811,N_7808);
or U7938 (N_7938,N_7874,N_7838);
nor U7939 (N_7939,N_7834,N_7899);
nand U7940 (N_7940,N_7832,N_7835);
and U7941 (N_7941,N_7865,N_7825);
xor U7942 (N_7942,N_7830,N_7849);
xnor U7943 (N_7943,N_7813,N_7863);
xnor U7944 (N_7944,N_7850,N_7807);
nor U7945 (N_7945,N_7815,N_7803);
nand U7946 (N_7946,N_7836,N_7828);
or U7947 (N_7947,N_7877,N_7868);
nor U7948 (N_7948,N_7888,N_7889);
and U7949 (N_7949,N_7887,N_7842);
or U7950 (N_7950,N_7893,N_7812);
or U7951 (N_7951,N_7857,N_7887);
xnor U7952 (N_7952,N_7811,N_7862);
nor U7953 (N_7953,N_7826,N_7800);
or U7954 (N_7954,N_7884,N_7800);
xnor U7955 (N_7955,N_7804,N_7827);
or U7956 (N_7956,N_7885,N_7828);
or U7957 (N_7957,N_7842,N_7811);
nand U7958 (N_7958,N_7847,N_7832);
or U7959 (N_7959,N_7862,N_7872);
nand U7960 (N_7960,N_7834,N_7898);
xnor U7961 (N_7961,N_7883,N_7862);
nand U7962 (N_7962,N_7811,N_7818);
and U7963 (N_7963,N_7826,N_7876);
and U7964 (N_7964,N_7899,N_7895);
nor U7965 (N_7965,N_7866,N_7867);
nand U7966 (N_7966,N_7815,N_7874);
or U7967 (N_7967,N_7816,N_7866);
or U7968 (N_7968,N_7812,N_7836);
and U7969 (N_7969,N_7873,N_7828);
nand U7970 (N_7970,N_7894,N_7829);
xor U7971 (N_7971,N_7820,N_7879);
and U7972 (N_7972,N_7859,N_7876);
nand U7973 (N_7973,N_7875,N_7804);
xor U7974 (N_7974,N_7888,N_7857);
and U7975 (N_7975,N_7835,N_7844);
xnor U7976 (N_7976,N_7859,N_7835);
xnor U7977 (N_7977,N_7829,N_7801);
nand U7978 (N_7978,N_7816,N_7860);
and U7979 (N_7979,N_7812,N_7834);
nor U7980 (N_7980,N_7805,N_7883);
or U7981 (N_7981,N_7868,N_7843);
and U7982 (N_7982,N_7823,N_7870);
or U7983 (N_7983,N_7841,N_7884);
or U7984 (N_7984,N_7897,N_7825);
xnor U7985 (N_7985,N_7803,N_7804);
or U7986 (N_7986,N_7846,N_7842);
or U7987 (N_7987,N_7859,N_7888);
and U7988 (N_7988,N_7883,N_7877);
nor U7989 (N_7989,N_7875,N_7852);
xor U7990 (N_7990,N_7890,N_7802);
and U7991 (N_7991,N_7884,N_7846);
xnor U7992 (N_7992,N_7865,N_7808);
or U7993 (N_7993,N_7888,N_7826);
xnor U7994 (N_7994,N_7816,N_7890);
xnor U7995 (N_7995,N_7812,N_7840);
and U7996 (N_7996,N_7867,N_7853);
nand U7997 (N_7997,N_7891,N_7881);
xor U7998 (N_7998,N_7840,N_7832);
nor U7999 (N_7999,N_7829,N_7827);
nor U8000 (N_8000,N_7936,N_7998);
or U8001 (N_8001,N_7987,N_7953);
xor U8002 (N_8002,N_7928,N_7955);
nand U8003 (N_8003,N_7933,N_7916);
or U8004 (N_8004,N_7926,N_7924);
nand U8005 (N_8005,N_7989,N_7994);
nand U8006 (N_8006,N_7913,N_7935);
nor U8007 (N_8007,N_7969,N_7918);
xor U8008 (N_8008,N_7995,N_7929);
and U8009 (N_8009,N_7981,N_7971);
and U8010 (N_8010,N_7992,N_7993);
or U8011 (N_8011,N_7947,N_7965);
nor U8012 (N_8012,N_7914,N_7973);
xor U8013 (N_8013,N_7906,N_7963);
nor U8014 (N_8014,N_7960,N_7937);
nand U8015 (N_8015,N_7911,N_7975);
and U8016 (N_8016,N_7991,N_7983);
xnor U8017 (N_8017,N_7938,N_7925);
xnor U8018 (N_8018,N_7988,N_7903);
and U8019 (N_8019,N_7917,N_7978);
nand U8020 (N_8020,N_7901,N_7967);
and U8021 (N_8021,N_7922,N_7970);
xnor U8022 (N_8022,N_7920,N_7908);
or U8023 (N_8023,N_7959,N_7980);
and U8024 (N_8024,N_7990,N_7964);
nor U8025 (N_8025,N_7958,N_7907);
nor U8026 (N_8026,N_7968,N_7909);
or U8027 (N_8027,N_7979,N_7910);
or U8028 (N_8028,N_7986,N_7984);
or U8029 (N_8029,N_7932,N_7950);
nor U8030 (N_8030,N_7997,N_7974);
or U8031 (N_8031,N_7957,N_7921);
and U8032 (N_8032,N_7900,N_7934);
xnor U8033 (N_8033,N_7912,N_7951);
nand U8034 (N_8034,N_7902,N_7948);
nor U8035 (N_8035,N_7927,N_7904);
nor U8036 (N_8036,N_7952,N_7946);
nor U8037 (N_8037,N_7966,N_7962);
xnor U8038 (N_8038,N_7943,N_7941);
nor U8039 (N_8039,N_7919,N_7954);
and U8040 (N_8040,N_7977,N_7923);
xor U8041 (N_8041,N_7939,N_7944);
xor U8042 (N_8042,N_7985,N_7942);
xnor U8043 (N_8043,N_7949,N_7961);
and U8044 (N_8044,N_7976,N_7931);
or U8045 (N_8045,N_7956,N_7915);
and U8046 (N_8046,N_7945,N_7905);
and U8047 (N_8047,N_7982,N_7996);
nand U8048 (N_8048,N_7972,N_7999);
nor U8049 (N_8049,N_7930,N_7940);
nor U8050 (N_8050,N_7912,N_7972);
and U8051 (N_8051,N_7951,N_7920);
xor U8052 (N_8052,N_7940,N_7968);
nand U8053 (N_8053,N_7908,N_7927);
nor U8054 (N_8054,N_7991,N_7926);
nor U8055 (N_8055,N_7918,N_7937);
and U8056 (N_8056,N_7966,N_7960);
nand U8057 (N_8057,N_7967,N_7966);
and U8058 (N_8058,N_7936,N_7939);
and U8059 (N_8059,N_7967,N_7964);
nand U8060 (N_8060,N_7911,N_7998);
nand U8061 (N_8061,N_7999,N_7941);
nand U8062 (N_8062,N_7946,N_7923);
xor U8063 (N_8063,N_7976,N_7913);
xnor U8064 (N_8064,N_7988,N_7975);
nor U8065 (N_8065,N_7968,N_7972);
nor U8066 (N_8066,N_7988,N_7931);
nor U8067 (N_8067,N_7965,N_7942);
or U8068 (N_8068,N_7946,N_7909);
or U8069 (N_8069,N_7910,N_7924);
nand U8070 (N_8070,N_7924,N_7977);
xnor U8071 (N_8071,N_7942,N_7934);
and U8072 (N_8072,N_7954,N_7908);
nand U8073 (N_8073,N_7945,N_7966);
xnor U8074 (N_8074,N_7970,N_7924);
xor U8075 (N_8075,N_7914,N_7987);
and U8076 (N_8076,N_7905,N_7923);
and U8077 (N_8077,N_7962,N_7952);
nor U8078 (N_8078,N_7901,N_7902);
and U8079 (N_8079,N_7923,N_7991);
and U8080 (N_8080,N_7933,N_7936);
or U8081 (N_8081,N_7977,N_7946);
xor U8082 (N_8082,N_7974,N_7978);
xor U8083 (N_8083,N_7970,N_7940);
xnor U8084 (N_8084,N_7934,N_7952);
and U8085 (N_8085,N_7906,N_7935);
or U8086 (N_8086,N_7904,N_7934);
nand U8087 (N_8087,N_7957,N_7969);
or U8088 (N_8088,N_7933,N_7914);
xor U8089 (N_8089,N_7920,N_7990);
nand U8090 (N_8090,N_7961,N_7964);
nand U8091 (N_8091,N_7920,N_7947);
and U8092 (N_8092,N_7960,N_7994);
and U8093 (N_8093,N_7983,N_7963);
nand U8094 (N_8094,N_7999,N_7967);
nor U8095 (N_8095,N_7901,N_7930);
and U8096 (N_8096,N_7942,N_7989);
nor U8097 (N_8097,N_7930,N_7957);
nand U8098 (N_8098,N_7963,N_7956);
nor U8099 (N_8099,N_7968,N_7943);
and U8100 (N_8100,N_8016,N_8046);
nor U8101 (N_8101,N_8085,N_8082);
or U8102 (N_8102,N_8033,N_8036);
and U8103 (N_8103,N_8031,N_8063);
xnor U8104 (N_8104,N_8070,N_8026);
xor U8105 (N_8105,N_8079,N_8062);
xor U8106 (N_8106,N_8096,N_8099);
or U8107 (N_8107,N_8009,N_8048);
nor U8108 (N_8108,N_8004,N_8003);
nor U8109 (N_8109,N_8090,N_8015);
xor U8110 (N_8110,N_8022,N_8011);
nor U8111 (N_8111,N_8053,N_8089);
nand U8112 (N_8112,N_8094,N_8068);
nand U8113 (N_8113,N_8006,N_8043);
nor U8114 (N_8114,N_8058,N_8092);
and U8115 (N_8115,N_8042,N_8086);
xnor U8116 (N_8116,N_8027,N_8038);
nand U8117 (N_8117,N_8071,N_8064);
nor U8118 (N_8118,N_8061,N_8047);
or U8119 (N_8119,N_8080,N_8052);
xnor U8120 (N_8120,N_8039,N_8037);
nand U8121 (N_8121,N_8057,N_8044);
and U8122 (N_8122,N_8075,N_8023);
or U8123 (N_8123,N_8069,N_8014);
and U8124 (N_8124,N_8017,N_8049);
xnor U8125 (N_8125,N_8073,N_8008);
nor U8126 (N_8126,N_8034,N_8012);
xnor U8127 (N_8127,N_8030,N_8081);
and U8128 (N_8128,N_8056,N_8084);
xnor U8129 (N_8129,N_8001,N_8007);
xor U8130 (N_8130,N_8041,N_8066);
and U8131 (N_8131,N_8060,N_8025);
nor U8132 (N_8132,N_8040,N_8013);
or U8133 (N_8133,N_8002,N_8051);
or U8134 (N_8134,N_8005,N_8029);
and U8135 (N_8135,N_8024,N_8072);
and U8136 (N_8136,N_8035,N_8021);
xor U8137 (N_8137,N_8098,N_8028);
nand U8138 (N_8138,N_8078,N_8074);
or U8139 (N_8139,N_8010,N_8045);
nand U8140 (N_8140,N_8093,N_8055);
and U8141 (N_8141,N_8087,N_8067);
nand U8142 (N_8142,N_8000,N_8083);
or U8143 (N_8143,N_8018,N_8054);
nand U8144 (N_8144,N_8059,N_8088);
nor U8145 (N_8145,N_8076,N_8091);
nor U8146 (N_8146,N_8095,N_8050);
xor U8147 (N_8147,N_8032,N_8097);
nor U8148 (N_8148,N_8077,N_8065);
nand U8149 (N_8149,N_8020,N_8019);
and U8150 (N_8150,N_8032,N_8056);
xor U8151 (N_8151,N_8049,N_8057);
or U8152 (N_8152,N_8027,N_8062);
and U8153 (N_8153,N_8012,N_8020);
nand U8154 (N_8154,N_8059,N_8023);
xnor U8155 (N_8155,N_8055,N_8007);
xnor U8156 (N_8156,N_8095,N_8072);
nand U8157 (N_8157,N_8079,N_8028);
nand U8158 (N_8158,N_8037,N_8075);
nor U8159 (N_8159,N_8040,N_8010);
or U8160 (N_8160,N_8053,N_8085);
and U8161 (N_8161,N_8076,N_8053);
or U8162 (N_8162,N_8024,N_8076);
xor U8163 (N_8163,N_8000,N_8075);
or U8164 (N_8164,N_8068,N_8079);
nand U8165 (N_8165,N_8051,N_8071);
nor U8166 (N_8166,N_8031,N_8017);
nand U8167 (N_8167,N_8022,N_8050);
xor U8168 (N_8168,N_8021,N_8085);
or U8169 (N_8169,N_8012,N_8094);
and U8170 (N_8170,N_8018,N_8070);
and U8171 (N_8171,N_8092,N_8053);
or U8172 (N_8172,N_8009,N_8041);
and U8173 (N_8173,N_8090,N_8018);
nor U8174 (N_8174,N_8008,N_8082);
nand U8175 (N_8175,N_8041,N_8043);
nand U8176 (N_8176,N_8026,N_8065);
nor U8177 (N_8177,N_8075,N_8019);
xor U8178 (N_8178,N_8072,N_8091);
nor U8179 (N_8179,N_8086,N_8055);
or U8180 (N_8180,N_8049,N_8032);
xor U8181 (N_8181,N_8003,N_8052);
and U8182 (N_8182,N_8028,N_8050);
xnor U8183 (N_8183,N_8017,N_8038);
xor U8184 (N_8184,N_8047,N_8004);
and U8185 (N_8185,N_8045,N_8011);
nor U8186 (N_8186,N_8006,N_8052);
or U8187 (N_8187,N_8068,N_8099);
and U8188 (N_8188,N_8053,N_8082);
xnor U8189 (N_8189,N_8016,N_8090);
and U8190 (N_8190,N_8059,N_8063);
and U8191 (N_8191,N_8064,N_8060);
and U8192 (N_8192,N_8000,N_8053);
nor U8193 (N_8193,N_8058,N_8028);
nand U8194 (N_8194,N_8012,N_8083);
xnor U8195 (N_8195,N_8050,N_8053);
or U8196 (N_8196,N_8005,N_8048);
nand U8197 (N_8197,N_8044,N_8070);
and U8198 (N_8198,N_8072,N_8075);
nor U8199 (N_8199,N_8078,N_8025);
or U8200 (N_8200,N_8121,N_8164);
and U8201 (N_8201,N_8196,N_8117);
nand U8202 (N_8202,N_8147,N_8149);
and U8203 (N_8203,N_8175,N_8158);
or U8204 (N_8204,N_8104,N_8124);
xor U8205 (N_8205,N_8167,N_8188);
or U8206 (N_8206,N_8179,N_8108);
and U8207 (N_8207,N_8152,N_8112);
nand U8208 (N_8208,N_8166,N_8142);
xor U8209 (N_8209,N_8105,N_8102);
nand U8210 (N_8210,N_8138,N_8132);
or U8211 (N_8211,N_8148,N_8194);
or U8212 (N_8212,N_8101,N_8192);
or U8213 (N_8213,N_8177,N_8125);
and U8214 (N_8214,N_8131,N_8155);
and U8215 (N_8215,N_8190,N_8172);
xor U8216 (N_8216,N_8186,N_8134);
xor U8217 (N_8217,N_8157,N_8116);
xor U8218 (N_8218,N_8174,N_8106);
or U8219 (N_8219,N_8137,N_8187);
nor U8220 (N_8220,N_8173,N_8144);
or U8221 (N_8221,N_8113,N_8176);
and U8222 (N_8222,N_8170,N_8133);
or U8223 (N_8223,N_8110,N_8111);
xor U8224 (N_8224,N_8139,N_8146);
xnor U8225 (N_8225,N_8150,N_8129);
nand U8226 (N_8226,N_8136,N_8160);
or U8227 (N_8227,N_8171,N_8159);
nand U8228 (N_8228,N_8199,N_8143);
nand U8229 (N_8229,N_8128,N_8191);
or U8230 (N_8230,N_8193,N_8130);
xor U8231 (N_8231,N_8156,N_8122);
nor U8232 (N_8232,N_8169,N_8161);
and U8233 (N_8233,N_8163,N_8118);
xor U8234 (N_8234,N_8151,N_8197);
xnor U8235 (N_8235,N_8119,N_8120);
xnor U8236 (N_8236,N_8107,N_8168);
and U8237 (N_8237,N_8103,N_8165);
and U8238 (N_8238,N_8114,N_8182);
xor U8239 (N_8239,N_8189,N_8183);
nor U8240 (N_8240,N_8145,N_8127);
or U8241 (N_8241,N_8115,N_8154);
nor U8242 (N_8242,N_8178,N_8126);
nand U8243 (N_8243,N_8140,N_8181);
xnor U8244 (N_8244,N_8185,N_8184);
nand U8245 (N_8245,N_8109,N_8195);
nor U8246 (N_8246,N_8162,N_8123);
nor U8247 (N_8247,N_8100,N_8153);
nand U8248 (N_8248,N_8135,N_8180);
nand U8249 (N_8249,N_8198,N_8141);
nor U8250 (N_8250,N_8145,N_8141);
and U8251 (N_8251,N_8164,N_8166);
or U8252 (N_8252,N_8154,N_8110);
xor U8253 (N_8253,N_8136,N_8194);
nand U8254 (N_8254,N_8135,N_8120);
or U8255 (N_8255,N_8105,N_8186);
xnor U8256 (N_8256,N_8157,N_8184);
and U8257 (N_8257,N_8131,N_8121);
nand U8258 (N_8258,N_8132,N_8179);
and U8259 (N_8259,N_8105,N_8177);
nor U8260 (N_8260,N_8195,N_8134);
xnor U8261 (N_8261,N_8129,N_8118);
and U8262 (N_8262,N_8174,N_8191);
and U8263 (N_8263,N_8122,N_8184);
and U8264 (N_8264,N_8168,N_8100);
or U8265 (N_8265,N_8136,N_8199);
nand U8266 (N_8266,N_8105,N_8150);
nor U8267 (N_8267,N_8173,N_8148);
nor U8268 (N_8268,N_8158,N_8187);
or U8269 (N_8269,N_8180,N_8185);
nand U8270 (N_8270,N_8128,N_8139);
or U8271 (N_8271,N_8192,N_8184);
nand U8272 (N_8272,N_8151,N_8190);
nor U8273 (N_8273,N_8107,N_8144);
nor U8274 (N_8274,N_8127,N_8104);
xnor U8275 (N_8275,N_8125,N_8194);
and U8276 (N_8276,N_8198,N_8107);
or U8277 (N_8277,N_8117,N_8182);
nor U8278 (N_8278,N_8146,N_8138);
nor U8279 (N_8279,N_8100,N_8132);
or U8280 (N_8280,N_8111,N_8103);
xor U8281 (N_8281,N_8184,N_8180);
and U8282 (N_8282,N_8180,N_8159);
or U8283 (N_8283,N_8107,N_8175);
nand U8284 (N_8284,N_8119,N_8146);
xor U8285 (N_8285,N_8173,N_8104);
and U8286 (N_8286,N_8104,N_8107);
xor U8287 (N_8287,N_8157,N_8166);
nand U8288 (N_8288,N_8179,N_8117);
or U8289 (N_8289,N_8123,N_8108);
and U8290 (N_8290,N_8160,N_8176);
nor U8291 (N_8291,N_8186,N_8148);
nor U8292 (N_8292,N_8152,N_8166);
nor U8293 (N_8293,N_8106,N_8165);
or U8294 (N_8294,N_8165,N_8132);
or U8295 (N_8295,N_8195,N_8197);
and U8296 (N_8296,N_8174,N_8169);
or U8297 (N_8297,N_8120,N_8162);
nand U8298 (N_8298,N_8129,N_8103);
nor U8299 (N_8299,N_8113,N_8165);
xor U8300 (N_8300,N_8233,N_8259);
and U8301 (N_8301,N_8260,N_8289);
and U8302 (N_8302,N_8215,N_8298);
nor U8303 (N_8303,N_8239,N_8299);
xnor U8304 (N_8304,N_8203,N_8235);
or U8305 (N_8305,N_8223,N_8224);
or U8306 (N_8306,N_8237,N_8227);
xor U8307 (N_8307,N_8232,N_8278);
nand U8308 (N_8308,N_8231,N_8202);
nor U8309 (N_8309,N_8252,N_8207);
and U8310 (N_8310,N_8256,N_8201);
or U8311 (N_8311,N_8247,N_8269);
xor U8312 (N_8312,N_8273,N_8220);
xnor U8313 (N_8313,N_8216,N_8234);
nand U8314 (N_8314,N_8257,N_8288);
or U8315 (N_8315,N_8229,N_8261);
xnor U8316 (N_8316,N_8205,N_8292);
nand U8317 (N_8317,N_8217,N_8226);
or U8318 (N_8318,N_8214,N_8254);
and U8319 (N_8319,N_8284,N_8244);
xnor U8320 (N_8320,N_8277,N_8212);
or U8321 (N_8321,N_8282,N_8287);
or U8322 (N_8322,N_8251,N_8296);
xor U8323 (N_8323,N_8267,N_8280);
xnor U8324 (N_8324,N_8290,N_8240);
nand U8325 (N_8325,N_8230,N_8211);
and U8326 (N_8326,N_8243,N_8218);
and U8327 (N_8327,N_8291,N_8249);
or U8328 (N_8328,N_8264,N_8294);
nand U8329 (N_8329,N_8255,N_8295);
and U8330 (N_8330,N_8285,N_8246);
and U8331 (N_8331,N_8209,N_8265);
and U8332 (N_8332,N_8204,N_8221);
nor U8333 (N_8333,N_8297,N_8208);
nor U8334 (N_8334,N_8248,N_8262);
xor U8335 (N_8335,N_8276,N_8253);
nor U8336 (N_8336,N_8222,N_8245);
xnor U8337 (N_8337,N_8286,N_8279);
nand U8338 (N_8338,N_8236,N_8270);
or U8339 (N_8339,N_8213,N_8225);
nand U8340 (N_8340,N_8274,N_8228);
xor U8341 (N_8341,N_8268,N_8241);
nand U8342 (N_8342,N_8271,N_8283);
nand U8343 (N_8343,N_8250,N_8206);
or U8344 (N_8344,N_8275,N_8238);
nand U8345 (N_8345,N_8200,N_8258);
and U8346 (N_8346,N_8219,N_8210);
and U8347 (N_8347,N_8293,N_8281);
nand U8348 (N_8348,N_8242,N_8263);
nor U8349 (N_8349,N_8272,N_8266);
xnor U8350 (N_8350,N_8235,N_8278);
and U8351 (N_8351,N_8267,N_8220);
or U8352 (N_8352,N_8205,N_8214);
xnor U8353 (N_8353,N_8228,N_8219);
or U8354 (N_8354,N_8299,N_8234);
or U8355 (N_8355,N_8251,N_8273);
nor U8356 (N_8356,N_8274,N_8208);
or U8357 (N_8357,N_8240,N_8210);
nand U8358 (N_8358,N_8273,N_8265);
nor U8359 (N_8359,N_8250,N_8269);
nand U8360 (N_8360,N_8259,N_8269);
nor U8361 (N_8361,N_8240,N_8297);
nor U8362 (N_8362,N_8279,N_8225);
or U8363 (N_8363,N_8204,N_8255);
and U8364 (N_8364,N_8280,N_8265);
and U8365 (N_8365,N_8266,N_8256);
nor U8366 (N_8366,N_8290,N_8278);
or U8367 (N_8367,N_8255,N_8228);
and U8368 (N_8368,N_8270,N_8212);
nor U8369 (N_8369,N_8244,N_8296);
or U8370 (N_8370,N_8257,N_8203);
and U8371 (N_8371,N_8270,N_8209);
or U8372 (N_8372,N_8218,N_8200);
nand U8373 (N_8373,N_8203,N_8209);
nor U8374 (N_8374,N_8216,N_8266);
or U8375 (N_8375,N_8284,N_8234);
and U8376 (N_8376,N_8216,N_8211);
and U8377 (N_8377,N_8249,N_8297);
nand U8378 (N_8378,N_8201,N_8257);
nor U8379 (N_8379,N_8273,N_8212);
nor U8380 (N_8380,N_8290,N_8216);
or U8381 (N_8381,N_8228,N_8253);
nor U8382 (N_8382,N_8214,N_8211);
xor U8383 (N_8383,N_8203,N_8206);
or U8384 (N_8384,N_8298,N_8214);
nand U8385 (N_8385,N_8263,N_8288);
or U8386 (N_8386,N_8227,N_8264);
or U8387 (N_8387,N_8209,N_8200);
or U8388 (N_8388,N_8275,N_8244);
nor U8389 (N_8389,N_8202,N_8274);
nand U8390 (N_8390,N_8262,N_8204);
nor U8391 (N_8391,N_8239,N_8233);
nand U8392 (N_8392,N_8265,N_8252);
nor U8393 (N_8393,N_8233,N_8250);
nor U8394 (N_8394,N_8216,N_8274);
nor U8395 (N_8395,N_8277,N_8227);
or U8396 (N_8396,N_8203,N_8287);
and U8397 (N_8397,N_8296,N_8203);
and U8398 (N_8398,N_8286,N_8227);
nor U8399 (N_8399,N_8278,N_8241);
nand U8400 (N_8400,N_8371,N_8344);
and U8401 (N_8401,N_8355,N_8380);
xor U8402 (N_8402,N_8396,N_8310);
and U8403 (N_8403,N_8386,N_8381);
xnor U8404 (N_8404,N_8327,N_8383);
or U8405 (N_8405,N_8394,N_8398);
or U8406 (N_8406,N_8370,N_8300);
nand U8407 (N_8407,N_8389,N_8397);
nor U8408 (N_8408,N_8393,N_8328);
and U8409 (N_8409,N_8365,N_8347);
and U8410 (N_8410,N_8313,N_8321);
and U8411 (N_8411,N_8353,N_8319);
xnor U8412 (N_8412,N_8356,N_8363);
and U8413 (N_8413,N_8316,N_8318);
nand U8414 (N_8414,N_8304,N_8366);
and U8415 (N_8415,N_8308,N_8341);
nor U8416 (N_8416,N_8358,N_8314);
or U8417 (N_8417,N_8331,N_8338);
nand U8418 (N_8418,N_8359,N_8361);
and U8419 (N_8419,N_8354,N_8306);
or U8420 (N_8420,N_8372,N_8326);
nor U8421 (N_8421,N_8364,N_8348);
nand U8422 (N_8422,N_8362,N_8312);
xnor U8423 (N_8423,N_8388,N_8350);
nand U8424 (N_8424,N_8367,N_8343);
nor U8425 (N_8425,N_8333,N_8307);
nor U8426 (N_8426,N_8334,N_8369);
nor U8427 (N_8427,N_8322,N_8390);
and U8428 (N_8428,N_8382,N_8373);
and U8429 (N_8429,N_8315,N_8339);
xor U8430 (N_8430,N_8305,N_8352);
xor U8431 (N_8431,N_8378,N_8346);
nand U8432 (N_8432,N_8387,N_8399);
xor U8433 (N_8433,N_8302,N_8360);
nor U8434 (N_8434,N_8332,N_8323);
or U8435 (N_8435,N_8309,N_8384);
xnor U8436 (N_8436,N_8391,N_8320);
or U8437 (N_8437,N_8336,N_8340);
or U8438 (N_8438,N_8311,N_8379);
nand U8439 (N_8439,N_8329,N_8375);
or U8440 (N_8440,N_8325,N_8317);
or U8441 (N_8441,N_8301,N_8349);
or U8442 (N_8442,N_8377,N_8357);
and U8443 (N_8443,N_8324,N_8376);
or U8444 (N_8444,N_8335,N_8368);
and U8445 (N_8445,N_8351,N_8345);
or U8446 (N_8446,N_8374,N_8385);
and U8447 (N_8447,N_8392,N_8337);
and U8448 (N_8448,N_8395,N_8342);
nor U8449 (N_8449,N_8330,N_8303);
nand U8450 (N_8450,N_8307,N_8320);
nand U8451 (N_8451,N_8374,N_8332);
nor U8452 (N_8452,N_8357,N_8315);
nand U8453 (N_8453,N_8361,N_8396);
xnor U8454 (N_8454,N_8364,N_8357);
and U8455 (N_8455,N_8367,N_8318);
or U8456 (N_8456,N_8311,N_8349);
xor U8457 (N_8457,N_8322,N_8378);
nor U8458 (N_8458,N_8309,N_8357);
and U8459 (N_8459,N_8339,N_8382);
or U8460 (N_8460,N_8351,N_8372);
nor U8461 (N_8461,N_8351,N_8341);
nor U8462 (N_8462,N_8337,N_8390);
or U8463 (N_8463,N_8310,N_8353);
xnor U8464 (N_8464,N_8349,N_8381);
nor U8465 (N_8465,N_8304,N_8330);
or U8466 (N_8466,N_8334,N_8361);
nand U8467 (N_8467,N_8325,N_8376);
or U8468 (N_8468,N_8351,N_8332);
xnor U8469 (N_8469,N_8364,N_8313);
or U8470 (N_8470,N_8359,N_8398);
nand U8471 (N_8471,N_8373,N_8340);
nand U8472 (N_8472,N_8365,N_8302);
xor U8473 (N_8473,N_8376,N_8316);
xor U8474 (N_8474,N_8372,N_8341);
nor U8475 (N_8475,N_8312,N_8395);
xor U8476 (N_8476,N_8385,N_8320);
or U8477 (N_8477,N_8311,N_8312);
nand U8478 (N_8478,N_8375,N_8326);
nand U8479 (N_8479,N_8351,N_8324);
xnor U8480 (N_8480,N_8301,N_8307);
nor U8481 (N_8481,N_8384,N_8376);
xor U8482 (N_8482,N_8336,N_8398);
xnor U8483 (N_8483,N_8398,N_8318);
and U8484 (N_8484,N_8362,N_8310);
and U8485 (N_8485,N_8330,N_8385);
nand U8486 (N_8486,N_8331,N_8314);
and U8487 (N_8487,N_8364,N_8376);
nand U8488 (N_8488,N_8359,N_8383);
xor U8489 (N_8489,N_8312,N_8344);
xor U8490 (N_8490,N_8360,N_8367);
and U8491 (N_8491,N_8307,N_8337);
and U8492 (N_8492,N_8365,N_8384);
or U8493 (N_8493,N_8346,N_8365);
nand U8494 (N_8494,N_8361,N_8381);
nor U8495 (N_8495,N_8395,N_8321);
nor U8496 (N_8496,N_8385,N_8357);
or U8497 (N_8497,N_8371,N_8312);
xor U8498 (N_8498,N_8332,N_8324);
xnor U8499 (N_8499,N_8388,N_8303);
or U8500 (N_8500,N_8437,N_8424);
nand U8501 (N_8501,N_8498,N_8404);
nand U8502 (N_8502,N_8401,N_8458);
xor U8503 (N_8503,N_8492,N_8417);
or U8504 (N_8504,N_8440,N_8407);
nand U8505 (N_8505,N_8484,N_8447);
and U8506 (N_8506,N_8410,N_8466);
nor U8507 (N_8507,N_8405,N_8496);
nand U8508 (N_8508,N_8469,N_8464);
and U8509 (N_8509,N_8448,N_8433);
nand U8510 (N_8510,N_8429,N_8455);
nand U8511 (N_8511,N_8478,N_8444);
xor U8512 (N_8512,N_8419,N_8415);
nand U8513 (N_8513,N_8480,N_8465);
and U8514 (N_8514,N_8445,N_8436);
nor U8515 (N_8515,N_8434,N_8477);
nand U8516 (N_8516,N_8406,N_8463);
nor U8517 (N_8517,N_8487,N_8425);
or U8518 (N_8518,N_8453,N_8499);
nand U8519 (N_8519,N_8493,N_8426);
nor U8520 (N_8520,N_8488,N_8411);
nor U8521 (N_8521,N_8471,N_8443);
xnor U8522 (N_8522,N_8486,N_8489);
or U8523 (N_8523,N_8467,N_8446);
and U8524 (N_8524,N_8402,N_8451);
nand U8525 (N_8525,N_8457,N_8412);
and U8526 (N_8526,N_8423,N_8470);
nand U8527 (N_8527,N_8416,N_8475);
nand U8528 (N_8528,N_8422,N_8460);
nor U8529 (N_8529,N_8441,N_8456);
and U8530 (N_8530,N_8418,N_8430);
and U8531 (N_8531,N_8431,N_8483);
nand U8532 (N_8532,N_8461,N_8491);
nand U8533 (N_8533,N_8485,N_8468);
or U8534 (N_8534,N_8473,N_8400);
nor U8535 (N_8535,N_8428,N_8474);
or U8536 (N_8536,N_8432,N_8459);
nand U8537 (N_8537,N_8450,N_8438);
nor U8538 (N_8538,N_8452,N_8449);
nand U8539 (N_8539,N_8494,N_8462);
xor U8540 (N_8540,N_8435,N_8408);
or U8541 (N_8541,N_8479,N_8420);
nand U8542 (N_8542,N_8421,N_8472);
nand U8543 (N_8543,N_8409,N_8495);
xor U8544 (N_8544,N_8413,N_8476);
xnor U8545 (N_8545,N_8427,N_8439);
and U8546 (N_8546,N_8490,N_8482);
or U8547 (N_8547,N_8454,N_8497);
nor U8548 (N_8548,N_8442,N_8414);
or U8549 (N_8549,N_8481,N_8403);
nand U8550 (N_8550,N_8440,N_8419);
xor U8551 (N_8551,N_8490,N_8450);
nor U8552 (N_8552,N_8492,N_8476);
nand U8553 (N_8553,N_8449,N_8413);
nor U8554 (N_8554,N_8426,N_8416);
or U8555 (N_8555,N_8437,N_8408);
nor U8556 (N_8556,N_8445,N_8405);
xnor U8557 (N_8557,N_8479,N_8400);
nand U8558 (N_8558,N_8405,N_8451);
nand U8559 (N_8559,N_8407,N_8458);
or U8560 (N_8560,N_8419,N_8438);
or U8561 (N_8561,N_8491,N_8456);
nand U8562 (N_8562,N_8448,N_8410);
or U8563 (N_8563,N_8457,N_8466);
nor U8564 (N_8564,N_8468,N_8426);
nand U8565 (N_8565,N_8415,N_8427);
nand U8566 (N_8566,N_8413,N_8414);
or U8567 (N_8567,N_8497,N_8447);
nand U8568 (N_8568,N_8476,N_8478);
nand U8569 (N_8569,N_8408,N_8430);
nand U8570 (N_8570,N_8444,N_8442);
nand U8571 (N_8571,N_8459,N_8442);
or U8572 (N_8572,N_8497,N_8489);
xnor U8573 (N_8573,N_8443,N_8419);
and U8574 (N_8574,N_8490,N_8445);
nand U8575 (N_8575,N_8455,N_8469);
nor U8576 (N_8576,N_8475,N_8428);
nor U8577 (N_8577,N_8421,N_8469);
or U8578 (N_8578,N_8407,N_8439);
and U8579 (N_8579,N_8434,N_8457);
and U8580 (N_8580,N_8449,N_8470);
nand U8581 (N_8581,N_8474,N_8418);
nor U8582 (N_8582,N_8414,N_8417);
nor U8583 (N_8583,N_8488,N_8413);
or U8584 (N_8584,N_8479,N_8424);
xor U8585 (N_8585,N_8461,N_8459);
nand U8586 (N_8586,N_8482,N_8488);
nor U8587 (N_8587,N_8484,N_8440);
and U8588 (N_8588,N_8466,N_8405);
nor U8589 (N_8589,N_8469,N_8493);
or U8590 (N_8590,N_8428,N_8441);
or U8591 (N_8591,N_8486,N_8471);
and U8592 (N_8592,N_8421,N_8437);
and U8593 (N_8593,N_8495,N_8461);
nor U8594 (N_8594,N_8401,N_8419);
xor U8595 (N_8595,N_8439,N_8416);
nand U8596 (N_8596,N_8460,N_8445);
nand U8597 (N_8597,N_8438,N_8470);
and U8598 (N_8598,N_8446,N_8401);
nand U8599 (N_8599,N_8446,N_8483);
xor U8600 (N_8600,N_8595,N_8558);
nor U8601 (N_8601,N_8589,N_8500);
and U8602 (N_8602,N_8516,N_8526);
or U8603 (N_8603,N_8586,N_8573);
or U8604 (N_8604,N_8531,N_8539);
nor U8605 (N_8605,N_8540,N_8552);
xor U8606 (N_8606,N_8533,N_8518);
xor U8607 (N_8607,N_8559,N_8582);
and U8608 (N_8608,N_8503,N_8564);
or U8609 (N_8609,N_8572,N_8515);
nand U8610 (N_8610,N_8545,N_8527);
and U8611 (N_8611,N_8512,N_8565);
nor U8612 (N_8612,N_8513,N_8594);
or U8613 (N_8613,N_8568,N_8535);
xor U8614 (N_8614,N_8560,N_8548);
or U8615 (N_8615,N_8549,N_8562);
nor U8616 (N_8616,N_8514,N_8566);
or U8617 (N_8617,N_8563,N_8561);
nand U8618 (N_8618,N_8576,N_8521);
nor U8619 (N_8619,N_8543,N_8583);
nand U8620 (N_8620,N_8569,N_8553);
nor U8621 (N_8621,N_8587,N_8599);
nor U8622 (N_8622,N_8551,N_8520);
xor U8623 (N_8623,N_8577,N_8550);
xnor U8624 (N_8624,N_8590,N_8554);
nor U8625 (N_8625,N_8597,N_8530);
nor U8626 (N_8626,N_8525,N_8502);
xor U8627 (N_8627,N_8593,N_8506);
and U8628 (N_8628,N_8546,N_8567);
or U8629 (N_8629,N_8532,N_8541);
xnor U8630 (N_8630,N_8547,N_8578);
xor U8631 (N_8631,N_8523,N_8517);
xor U8632 (N_8632,N_8528,N_8575);
or U8633 (N_8633,N_8529,N_8591);
and U8634 (N_8634,N_8579,N_8570);
xor U8635 (N_8635,N_8596,N_8504);
nand U8636 (N_8636,N_8507,N_8584);
nor U8637 (N_8637,N_8519,N_8580);
and U8638 (N_8638,N_8557,N_8524);
or U8639 (N_8639,N_8510,N_8592);
or U8640 (N_8640,N_8581,N_8509);
and U8641 (N_8641,N_8511,N_8505);
and U8642 (N_8642,N_8571,N_8534);
nor U8643 (N_8643,N_8585,N_8501);
nor U8644 (N_8644,N_8556,N_8522);
or U8645 (N_8645,N_8542,N_8508);
or U8646 (N_8646,N_8544,N_8538);
nand U8647 (N_8647,N_8555,N_8588);
nor U8648 (N_8648,N_8536,N_8598);
or U8649 (N_8649,N_8574,N_8537);
nor U8650 (N_8650,N_8503,N_8573);
or U8651 (N_8651,N_8513,N_8517);
and U8652 (N_8652,N_8528,N_8590);
and U8653 (N_8653,N_8517,N_8567);
xnor U8654 (N_8654,N_8502,N_8596);
xnor U8655 (N_8655,N_8596,N_8588);
or U8656 (N_8656,N_8532,N_8517);
and U8657 (N_8657,N_8547,N_8536);
nand U8658 (N_8658,N_8519,N_8536);
and U8659 (N_8659,N_8570,N_8568);
or U8660 (N_8660,N_8502,N_8530);
or U8661 (N_8661,N_8535,N_8565);
xnor U8662 (N_8662,N_8578,N_8522);
nor U8663 (N_8663,N_8545,N_8538);
and U8664 (N_8664,N_8594,N_8543);
or U8665 (N_8665,N_8549,N_8552);
and U8666 (N_8666,N_8580,N_8542);
or U8667 (N_8667,N_8587,N_8543);
xor U8668 (N_8668,N_8517,N_8522);
or U8669 (N_8669,N_8507,N_8532);
xor U8670 (N_8670,N_8597,N_8592);
or U8671 (N_8671,N_8547,N_8516);
or U8672 (N_8672,N_8585,N_8566);
xnor U8673 (N_8673,N_8556,N_8548);
nor U8674 (N_8674,N_8567,N_8582);
nor U8675 (N_8675,N_8539,N_8581);
or U8676 (N_8676,N_8599,N_8532);
and U8677 (N_8677,N_8512,N_8572);
or U8678 (N_8678,N_8523,N_8598);
nand U8679 (N_8679,N_8537,N_8551);
and U8680 (N_8680,N_8530,N_8546);
xnor U8681 (N_8681,N_8516,N_8501);
or U8682 (N_8682,N_8528,N_8525);
or U8683 (N_8683,N_8546,N_8572);
or U8684 (N_8684,N_8507,N_8580);
xor U8685 (N_8685,N_8545,N_8520);
nor U8686 (N_8686,N_8526,N_8590);
or U8687 (N_8687,N_8540,N_8565);
and U8688 (N_8688,N_8547,N_8584);
xor U8689 (N_8689,N_8511,N_8501);
xnor U8690 (N_8690,N_8542,N_8515);
or U8691 (N_8691,N_8503,N_8532);
or U8692 (N_8692,N_8506,N_8599);
nand U8693 (N_8693,N_8575,N_8531);
nor U8694 (N_8694,N_8527,N_8543);
and U8695 (N_8695,N_8506,N_8502);
nand U8696 (N_8696,N_8500,N_8597);
or U8697 (N_8697,N_8588,N_8531);
nand U8698 (N_8698,N_8501,N_8500);
or U8699 (N_8699,N_8563,N_8560);
xnor U8700 (N_8700,N_8633,N_8663);
or U8701 (N_8701,N_8635,N_8694);
and U8702 (N_8702,N_8664,N_8668);
or U8703 (N_8703,N_8613,N_8648);
xor U8704 (N_8704,N_8655,N_8665);
nand U8705 (N_8705,N_8634,N_8617);
xnor U8706 (N_8706,N_8653,N_8658);
nor U8707 (N_8707,N_8626,N_8632);
xnor U8708 (N_8708,N_8609,N_8639);
xor U8709 (N_8709,N_8611,N_8676);
and U8710 (N_8710,N_8678,N_8644);
or U8711 (N_8711,N_8691,N_8685);
or U8712 (N_8712,N_8607,N_8687);
nor U8713 (N_8713,N_8621,N_8647);
or U8714 (N_8714,N_8681,N_8637);
or U8715 (N_8715,N_8624,N_8698);
nand U8716 (N_8716,N_8628,N_8640);
xnor U8717 (N_8717,N_8686,N_8659);
nor U8718 (N_8718,N_8649,N_8604);
and U8719 (N_8719,N_8669,N_8684);
nand U8720 (N_8720,N_8638,N_8616);
and U8721 (N_8721,N_8661,N_8606);
nand U8722 (N_8722,N_8682,N_8654);
and U8723 (N_8723,N_8651,N_8615);
nor U8724 (N_8724,N_8693,N_8630);
and U8725 (N_8725,N_8667,N_8619);
nor U8726 (N_8726,N_8618,N_8697);
nand U8727 (N_8727,N_8673,N_8672);
nor U8728 (N_8728,N_8696,N_8614);
or U8729 (N_8729,N_8603,N_8652);
nor U8730 (N_8730,N_8623,N_8692);
nor U8731 (N_8731,N_8662,N_8660);
xor U8732 (N_8732,N_8679,N_8602);
and U8733 (N_8733,N_8625,N_8656);
or U8734 (N_8734,N_8650,N_8643);
nor U8735 (N_8735,N_8671,N_8629);
nor U8736 (N_8736,N_8675,N_8645);
and U8737 (N_8737,N_8627,N_8605);
and U8738 (N_8738,N_8636,N_8657);
or U8739 (N_8739,N_8610,N_8674);
or U8740 (N_8740,N_8631,N_8622);
nor U8741 (N_8741,N_8677,N_8699);
nor U8742 (N_8742,N_8666,N_8601);
nor U8743 (N_8743,N_8642,N_8688);
nor U8744 (N_8744,N_8612,N_8600);
nand U8745 (N_8745,N_8680,N_8608);
or U8746 (N_8746,N_8695,N_8689);
nor U8747 (N_8747,N_8646,N_8690);
nand U8748 (N_8748,N_8620,N_8641);
nand U8749 (N_8749,N_8683,N_8670);
nor U8750 (N_8750,N_8650,N_8620);
xnor U8751 (N_8751,N_8621,N_8661);
nor U8752 (N_8752,N_8686,N_8674);
xor U8753 (N_8753,N_8684,N_8697);
and U8754 (N_8754,N_8663,N_8635);
or U8755 (N_8755,N_8666,N_8643);
xnor U8756 (N_8756,N_8677,N_8610);
xor U8757 (N_8757,N_8646,N_8614);
and U8758 (N_8758,N_8699,N_8661);
nand U8759 (N_8759,N_8686,N_8634);
and U8760 (N_8760,N_8633,N_8666);
nor U8761 (N_8761,N_8685,N_8600);
xnor U8762 (N_8762,N_8646,N_8643);
or U8763 (N_8763,N_8636,N_8671);
nor U8764 (N_8764,N_8663,N_8670);
xnor U8765 (N_8765,N_8652,N_8651);
nand U8766 (N_8766,N_8614,N_8628);
nor U8767 (N_8767,N_8658,N_8602);
nand U8768 (N_8768,N_8658,N_8682);
or U8769 (N_8769,N_8674,N_8678);
or U8770 (N_8770,N_8666,N_8664);
or U8771 (N_8771,N_8643,N_8677);
xnor U8772 (N_8772,N_8683,N_8658);
nor U8773 (N_8773,N_8609,N_8606);
or U8774 (N_8774,N_8649,N_8620);
nand U8775 (N_8775,N_8643,N_8632);
nor U8776 (N_8776,N_8617,N_8667);
or U8777 (N_8777,N_8664,N_8682);
and U8778 (N_8778,N_8623,N_8657);
nor U8779 (N_8779,N_8603,N_8694);
nand U8780 (N_8780,N_8698,N_8637);
xor U8781 (N_8781,N_8632,N_8657);
or U8782 (N_8782,N_8679,N_8654);
xor U8783 (N_8783,N_8677,N_8625);
nor U8784 (N_8784,N_8679,N_8622);
xnor U8785 (N_8785,N_8650,N_8673);
nand U8786 (N_8786,N_8683,N_8624);
nor U8787 (N_8787,N_8668,N_8630);
and U8788 (N_8788,N_8667,N_8681);
or U8789 (N_8789,N_8673,N_8666);
xnor U8790 (N_8790,N_8617,N_8662);
or U8791 (N_8791,N_8679,N_8620);
xnor U8792 (N_8792,N_8646,N_8695);
nand U8793 (N_8793,N_8666,N_8656);
nand U8794 (N_8794,N_8614,N_8676);
nor U8795 (N_8795,N_8644,N_8608);
or U8796 (N_8796,N_8606,N_8689);
nor U8797 (N_8797,N_8645,N_8670);
nor U8798 (N_8798,N_8676,N_8609);
nand U8799 (N_8799,N_8691,N_8629);
xnor U8800 (N_8800,N_8733,N_8700);
xnor U8801 (N_8801,N_8766,N_8714);
nor U8802 (N_8802,N_8723,N_8734);
nor U8803 (N_8803,N_8779,N_8755);
nor U8804 (N_8804,N_8710,N_8768);
xor U8805 (N_8805,N_8712,N_8754);
nor U8806 (N_8806,N_8706,N_8717);
and U8807 (N_8807,N_8713,N_8780);
and U8808 (N_8808,N_8789,N_8751);
nand U8809 (N_8809,N_8720,N_8764);
or U8810 (N_8810,N_8790,N_8739);
xor U8811 (N_8811,N_8781,N_8722);
nor U8812 (N_8812,N_8731,N_8741);
or U8813 (N_8813,N_8775,N_8743);
nand U8814 (N_8814,N_8784,N_8787);
nor U8815 (N_8815,N_8763,N_8715);
nor U8816 (N_8816,N_8718,N_8707);
nand U8817 (N_8817,N_8794,N_8736);
or U8818 (N_8818,N_8742,N_8758);
nor U8819 (N_8819,N_8747,N_8785);
nor U8820 (N_8820,N_8765,N_8708);
nor U8821 (N_8821,N_8767,N_8778);
xnor U8822 (N_8822,N_8735,N_8797);
nor U8823 (N_8823,N_8705,N_8725);
and U8824 (N_8824,N_8732,N_8709);
and U8825 (N_8825,N_8738,N_8729);
and U8826 (N_8826,N_8791,N_8748);
or U8827 (N_8827,N_8724,N_8737);
xor U8828 (N_8828,N_8752,N_8796);
nand U8829 (N_8829,N_8711,N_8798);
and U8830 (N_8830,N_8745,N_8740);
and U8831 (N_8831,N_8793,N_8772);
xor U8832 (N_8832,N_8770,N_8769);
nand U8833 (N_8833,N_8757,N_8762);
xnor U8834 (N_8834,N_8759,N_8702);
nand U8835 (N_8835,N_8777,N_8776);
or U8836 (N_8836,N_8786,N_8792);
and U8837 (N_8837,N_8749,N_8704);
and U8838 (N_8838,N_8771,N_8774);
nor U8839 (N_8839,N_8756,N_8726);
nor U8840 (N_8840,N_8703,N_8744);
nor U8841 (N_8841,N_8716,N_8746);
nand U8842 (N_8842,N_8728,N_8773);
or U8843 (N_8843,N_8760,N_8753);
xnor U8844 (N_8844,N_8761,N_8701);
nor U8845 (N_8845,N_8795,N_8799);
nor U8846 (N_8846,N_8721,N_8783);
xor U8847 (N_8847,N_8719,N_8782);
and U8848 (N_8848,N_8750,N_8730);
nor U8849 (N_8849,N_8788,N_8727);
nand U8850 (N_8850,N_8738,N_8791);
nand U8851 (N_8851,N_8720,N_8725);
nor U8852 (N_8852,N_8718,N_8703);
nor U8853 (N_8853,N_8757,N_8743);
and U8854 (N_8854,N_8731,N_8723);
and U8855 (N_8855,N_8715,N_8722);
nor U8856 (N_8856,N_8792,N_8799);
xor U8857 (N_8857,N_8715,N_8705);
xor U8858 (N_8858,N_8729,N_8774);
nor U8859 (N_8859,N_8773,N_8710);
or U8860 (N_8860,N_8707,N_8798);
and U8861 (N_8861,N_8701,N_8789);
nand U8862 (N_8862,N_8749,N_8768);
xnor U8863 (N_8863,N_8772,N_8778);
nand U8864 (N_8864,N_8722,N_8732);
nand U8865 (N_8865,N_8785,N_8757);
and U8866 (N_8866,N_8735,N_8774);
nor U8867 (N_8867,N_8717,N_8744);
nand U8868 (N_8868,N_8715,N_8766);
xnor U8869 (N_8869,N_8706,N_8710);
xor U8870 (N_8870,N_8753,N_8700);
and U8871 (N_8871,N_8756,N_8706);
xnor U8872 (N_8872,N_8724,N_8784);
nand U8873 (N_8873,N_8777,N_8736);
nand U8874 (N_8874,N_8792,N_8751);
nand U8875 (N_8875,N_8748,N_8794);
nand U8876 (N_8876,N_8788,N_8730);
nor U8877 (N_8877,N_8718,N_8786);
nand U8878 (N_8878,N_8722,N_8730);
nor U8879 (N_8879,N_8708,N_8747);
xnor U8880 (N_8880,N_8747,N_8786);
or U8881 (N_8881,N_8758,N_8774);
nand U8882 (N_8882,N_8742,N_8785);
xnor U8883 (N_8883,N_8721,N_8774);
nor U8884 (N_8884,N_8791,N_8706);
xnor U8885 (N_8885,N_8739,N_8793);
xor U8886 (N_8886,N_8772,N_8798);
and U8887 (N_8887,N_8724,N_8792);
or U8888 (N_8888,N_8707,N_8774);
nor U8889 (N_8889,N_8776,N_8739);
or U8890 (N_8890,N_8734,N_8710);
nand U8891 (N_8891,N_8748,N_8754);
nor U8892 (N_8892,N_8763,N_8724);
nor U8893 (N_8893,N_8739,N_8705);
or U8894 (N_8894,N_8760,N_8706);
or U8895 (N_8895,N_8777,N_8722);
or U8896 (N_8896,N_8747,N_8766);
and U8897 (N_8897,N_8726,N_8754);
xor U8898 (N_8898,N_8793,N_8767);
or U8899 (N_8899,N_8795,N_8759);
or U8900 (N_8900,N_8846,N_8890);
and U8901 (N_8901,N_8885,N_8860);
and U8902 (N_8902,N_8865,N_8843);
nor U8903 (N_8903,N_8802,N_8883);
or U8904 (N_8904,N_8880,N_8874);
nor U8905 (N_8905,N_8822,N_8857);
nor U8906 (N_8906,N_8800,N_8878);
nor U8907 (N_8907,N_8816,N_8868);
nand U8908 (N_8908,N_8813,N_8819);
nand U8909 (N_8909,N_8882,N_8830);
or U8910 (N_8910,N_8814,N_8825);
xor U8911 (N_8911,N_8806,N_8867);
xnor U8912 (N_8912,N_8840,N_8848);
and U8913 (N_8913,N_8851,N_8892);
and U8914 (N_8914,N_8881,N_8844);
nor U8915 (N_8915,N_8828,N_8864);
and U8916 (N_8916,N_8872,N_8884);
xnor U8917 (N_8917,N_8899,N_8858);
or U8918 (N_8918,N_8836,N_8850);
and U8919 (N_8919,N_8854,N_8877);
or U8920 (N_8920,N_8801,N_8886);
or U8921 (N_8921,N_8862,N_8827);
xor U8922 (N_8922,N_8845,N_8863);
nor U8923 (N_8923,N_8834,N_8841);
nor U8924 (N_8924,N_8837,N_8897);
nand U8925 (N_8925,N_8812,N_8817);
nand U8926 (N_8926,N_8804,N_8898);
xor U8927 (N_8927,N_8831,N_8809);
nand U8928 (N_8928,N_8871,N_8808);
nor U8929 (N_8929,N_8824,N_8810);
or U8930 (N_8930,N_8866,N_8889);
nor U8931 (N_8931,N_8873,N_8896);
or U8932 (N_8932,N_8823,N_8856);
nor U8933 (N_8933,N_8859,N_8833);
xnor U8934 (N_8934,N_8805,N_8838);
xor U8935 (N_8935,N_8879,N_8835);
nand U8936 (N_8936,N_8869,N_8842);
nor U8937 (N_8937,N_8888,N_8893);
xor U8938 (N_8938,N_8891,N_8811);
and U8939 (N_8939,N_8818,N_8847);
nor U8940 (N_8940,N_8832,N_8826);
or U8941 (N_8941,N_8895,N_8807);
and U8942 (N_8942,N_8853,N_8894);
or U8943 (N_8943,N_8829,N_8870);
and U8944 (N_8944,N_8887,N_8849);
and U8945 (N_8945,N_8855,N_8821);
nand U8946 (N_8946,N_8875,N_8820);
nor U8947 (N_8947,N_8803,N_8815);
nand U8948 (N_8948,N_8876,N_8852);
nand U8949 (N_8949,N_8861,N_8839);
or U8950 (N_8950,N_8816,N_8890);
xnor U8951 (N_8951,N_8891,N_8806);
or U8952 (N_8952,N_8801,N_8865);
nor U8953 (N_8953,N_8831,N_8875);
nand U8954 (N_8954,N_8850,N_8824);
nor U8955 (N_8955,N_8803,N_8811);
or U8956 (N_8956,N_8827,N_8813);
and U8957 (N_8957,N_8821,N_8801);
nor U8958 (N_8958,N_8892,N_8821);
nor U8959 (N_8959,N_8898,N_8819);
and U8960 (N_8960,N_8890,N_8836);
and U8961 (N_8961,N_8885,N_8853);
xor U8962 (N_8962,N_8844,N_8849);
or U8963 (N_8963,N_8887,N_8806);
and U8964 (N_8964,N_8867,N_8879);
nand U8965 (N_8965,N_8875,N_8858);
nor U8966 (N_8966,N_8882,N_8823);
and U8967 (N_8967,N_8845,N_8806);
or U8968 (N_8968,N_8826,N_8871);
or U8969 (N_8969,N_8805,N_8850);
xor U8970 (N_8970,N_8851,N_8895);
or U8971 (N_8971,N_8845,N_8822);
nor U8972 (N_8972,N_8867,N_8857);
nor U8973 (N_8973,N_8819,N_8815);
and U8974 (N_8974,N_8886,N_8871);
or U8975 (N_8975,N_8826,N_8828);
nand U8976 (N_8976,N_8853,N_8800);
or U8977 (N_8977,N_8860,N_8803);
xnor U8978 (N_8978,N_8826,N_8892);
nor U8979 (N_8979,N_8895,N_8823);
xor U8980 (N_8980,N_8839,N_8811);
nand U8981 (N_8981,N_8879,N_8884);
nand U8982 (N_8982,N_8886,N_8894);
xnor U8983 (N_8983,N_8859,N_8875);
or U8984 (N_8984,N_8880,N_8817);
or U8985 (N_8985,N_8882,N_8811);
or U8986 (N_8986,N_8860,N_8800);
nand U8987 (N_8987,N_8804,N_8832);
xor U8988 (N_8988,N_8843,N_8808);
nand U8989 (N_8989,N_8854,N_8899);
nor U8990 (N_8990,N_8899,N_8807);
nor U8991 (N_8991,N_8862,N_8815);
and U8992 (N_8992,N_8868,N_8800);
and U8993 (N_8993,N_8809,N_8865);
and U8994 (N_8994,N_8834,N_8842);
nor U8995 (N_8995,N_8848,N_8884);
xnor U8996 (N_8996,N_8855,N_8894);
nand U8997 (N_8997,N_8845,N_8856);
or U8998 (N_8998,N_8885,N_8875);
nor U8999 (N_8999,N_8894,N_8832);
xor U9000 (N_9000,N_8967,N_8902);
or U9001 (N_9001,N_8998,N_8921);
and U9002 (N_9002,N_8985,N_8959);
nand U9003 (N_9003,N_8980,N_8907);
nor U9004 (N_9004,N_8957,N_8971);
and U9005 (N_9005,N_8984,N_8900);
nor U9006 (N_9006,N_8938,N_8905);
nor U9007 (N_9007,N_8910,N_8963);
or U9008 (N_9008,N_8974,N_8964);
and U9009 (N_9009,N_8925,N_8932);
nand U9010 (N_9010,N_8966,N_8996);
or U9011 (N_9011,N_8968,N_8989);
xor U9012 (N_9012,N_8955,N_8906);
nor U9013 (N_9013,N_8937,N_8960);
nand U9014 (N_9014,N_8927,N_8934);
xnor U9015 (N_9015,N_8991,N_8986);
xor U9016 (N_9016,N_8935,N_8928);
nand U9017 (N_9017,N_8983,N_8987);
nand U9018 (N_9018,N_8915,N_8930);
xor U9019 (N_9019,N_8949,N_8982);
nor U9020 (N_9020,N_8943,N_8948);
or U9021 (N_9021,N_8961,N_8919);
xor U9022 (N_9022,N_8976,N_8901);
xnor U9023 (N_9023,N_8941,N_8994);
or U9024 (N_9024,N_8947,N_8920);
nand U9025 (N_9025,N_8926,N_8979);
nand U9026 (N_9026,N_8946,N_8954);
and U9027 (N_9027,N_8956,N_8981);
xor U9028 (N_9028,N_8903,N_8978);
nand U9029 (N_9029,N_8988,N_8951);
or U9030 (N_9030,N_8972,N_8965);
nand U9031 (N_9031,N_8962,N_8913);
nor U9032 (N_9032,N_8952,N_8939);
and U9033 (N_9033,N_8993,N_8922);
nor U9034 (N_9034,N_8916,N_8992);
nand U9035 (N_9035,N_8969,N_8911);
and U9036 (N_9036,N_8917,N_8936);
and U9037 (N_9037,N_8909,N_8944);
xnor U9038 (N_9038,N_8908,N_8923);
xnor U9039 (N_9039,N_8958,N_8929);
and U9040 (N_9040,N_8975,N_8977);
nor U9041 (N_9041,N_8953,N_8970);
xor U9042 (N_9042,N_8973,N_8945);
nand U9043 (N_9043,N_8918,N_8914);
and U9044 (N_9044,N_8950,N_8995);
or U9045 (N_9045,N_8912,N_8931);
nand U9046 (N_9046,N_8999,N_8933);
nand U9047 (N_9047,N_8924,N_8990);
and U9048 (N_9048,N_8942,N_8997);
nand U9049 (N_9049,N_8940,N_8904);
and U9050 (N_9050,N_8992,N_8941);
and U9051 (N_9051,N_8928,N_8991);
nor U9052 (N_9052,N_8975,N_8983);
nor U9053 (N_9053,N_8909,N_8997);
nor U9054 (N_9054,N_8919,N_8938);
nand U9055 (N_9055,N_8904,N_8914);
and U9056 (N_9056,N_8902,N_8947);
or U9057 (N_9057,N_8980,N_8999);
and U9058 (N_9058,N_8956,N_8961);
nand U9059 (N_9059,N_8992,N_8900);
and U9060 (N_9060,N_8919,N_8900);
and U9061 (N_9061,N_8924,N_8950);
or U9062 (N_9062,N_8997,N_8946);
xor U9063 (N_9063,N_8998,N_8956);
xnor U9064 (N_9064,N_8963,N_8990);
nand U9065 (N_9065,N_8934,N_8905);
nor U9066 (N_9066,N_8953,N_8949);
or U9067 (N_9067,N_8987,N_8978);
or U9068 (N_9068,N_8980,N_8933);
nor U9069 (N_9069,N_8923,N_8947);
and U9070 (N_9070,N_8941,N_8951);
nor U9071 (N_9071,N_8912,N_8977);
or U9072 (N_9072,N_8985,N_8964);
nor U9073 (N_9073,N_8936,N_8965);
nand U9074 (N_9074,N_8917,N_8926);
nor U9075 (N_9075,N_8981,N_8932);
nand U9076 (N_9076,N_8934,N_8974);
nand U9077 (N_9077,N_8913,N_8967);
and U9078 (N_9078,N_8931,N_8970);
or U9079 (N_9079,N_8960,N_8901);
xnor U9080 (N_9080,N_8972,N_8993);
xnor U9081 (N_9081,N_8930,N_8975);
nor U9082 (N_9082,N_8941,N_8940);
and U9083 (N_9083,N_8943,N_8991);
xor U9084 (N_9084,N_8913,N_8989);
and U9085 (N_9085,N_8922,N_8912);
nor U9086 (N_9086,N_8943,N_8978);
or U9087 (N_9087,N_8926,N_8936);
or U9088 (N_9088,N_8910,N_8986);
or U9089 (N_9089,N_8934,N_8954);
nand U9090 (N_9090,N_8933,N_8968);
nand U9091 (N_9091,N_8998,N_8901);
xnor U9092 (N_9092,N_8958,N_8993);
nand U9093 (N_9093,N_8999,N_8987);
xor U9094 (N_9094,N_8960,N_8947);
or U9095 (N_9095,N_8976,N_8935);
and U9096 (N_9096,N_8900,N_8955);
nor U9097 (N_9097,N_8914,N_8915);
xor U9098 (N_9098,N_8935,N_8923);
nand U9099 (N_9099,N_8935,N_8960);
or U9100 (N_9100,N_9019,N_9039);
or U9101 (N_9101,N_9099,N_9073);
xnor U9102 (N_9102,N_9083,N_9015);
xor U9103 (N_9103,N_9036,N_9060);
and U9104 (N_9104,N_9066,N_9041);
nor U9105 (N_9105,N_9009,N_9017);
nor U9106 (N_9106,N_9046,N_9059);
or U9107 (N_9107,N_9054,N_9023);
or U9108 (N_9108,N_9026,N_9033);
nand U9109 (N_9109,N_9000,N_9052);
nand U9110 (N_9110,N_9035,N_9038);
and U9111 (N_9111,N_9088,N_9032);
or U9112 (N_9112,N_9040,N_9013);
nand U9113 (N_9113,N_9006,N_9055);
xor U9114 (N_9114,N_9048,N_9016);
and U9115 (N_9115,N_9081,N_9091);
and U9116 (N_9116,N_9062,N_9098);
nor U9117 (N_9117,N_9008,N_9064);
or U9118 (N_9118,N_9012,N_9043);
nand U9119 (N_9119,N_9082,N_9056);
and U9120 (N_9120,N_9020,N_9049);
or U9121 (N_9121,N_9086,N_9045);
nand U9122 (N_9122,N_9002,N_9094);
nor U9123 (N_9123,N_9097,N_9072);
xor U9124 (N_9124,N_9010,N_9079);
or U9125 (N_9125,N_9004,N_9077);
or U9126 (N_9126,N_9057,N_9018);
nand U9127 (N_9127,N_9031,N_9075);
or U9128 (N_9128,N_9076,N_9037);
or U9129 (N_9129,N_9047,N_9061);
xnor U9130 (N_9130,N_9070,N_9001);
nor U9131 (N_9131,N_9005,N_9065);
and U9132 (N_9132,N_9014,N_9024);
or U9133 (N_9133,N_9027,N_9050);
nand U9134 (N_9134,N_9029,N_9051);
nor U9135 (N_9135,N_9028,N_9058);
nor U9136 (N_9136,N_9093,N_9085);
nor U9137 (N_9137,N_9021,N_9074);
and U9138 (N_9138,N_9080,N_9022);
and U9139 (N_9139,N_9068,N_9084);
xor U9140 (N_9140,N_9090,N_9011);
nor U9141 (N_9141,N_9030,N_9069);
nand U9142 (N_9142,N_9071,N_9096);
nand U9143 (N_9143,N_9087,N_9042);
nor U9144 (N_9144,N_9007,N_9089);
nor U9145 (N_9145,N_9003,N_9063);
and U9146 (N_9146,N_9092,N_9025);
or U9147 (N_9147,N_9034,N_9078);
or U9148 (N_9148,N_9053,N_9095);
and U9149 (N_9149,N_9044,N_9067);
or U9150 (N_9150,N_9031,N_9049);
xor U9151 (N_9151,N_9099,N_9039);
or U9152 (N_9152,N_9032,N_9089);
nand U9153 (N_9153,N_9045,N_9083);
nor U9154 (N_9154,N_9043,N_9017);
nand U9155 (N_9155,N_9010,N_9005);
or U9156 (N_9156,N_9053,N_9047);
nand U9157 (N_9157,N_9024,N_9079);
nor U9158 (N_9158,N_9078,N_9075);
and U9159 (N_9159,N_9096,N_9022);
nand U9160 (N_9160,N_9077,N_9089);
and U9161 (N_9161,N_9008,N_9028);
xnor U9162 (N_9162,N_9020,N_9079);
nand U9163 (N_9163,N_9090,N_9014);
or U9164 (N_9164,N_9003,N_9044);
xnor U9165 (N_9165,N_9025,N_9035);
and U9166 (N_9166,N_9025,N_9099);
and U9167 (N_9167,N_9094,N_9089);
xnor U9168 (N_9168,N_9032,N_9099);
nand U9169 (N_9169,N_9072,N_9014);
or U9170 (N_9170,N_9000,N_9071);
and U9171 (N_9171,N_9006,N_9020);
xor U9172 (N_9172,N_9019,N_9060);
nand U9173 (N_9173,N_9061,N_9089);
and U9174 (N_9174,N_9050,N_9002);
or U9175 (N_9175,N_9015,N_9072);
nand U9176 (N_9176,N_9018,N_9005);
nand U9177 (N_9177,N_9017,N_9085);
nand U9178 (N_9178,N_9004,N_9085);
and U9179 (N_9179,N_9090,N_9081);
nand U9180 (N_9180,N_9043,N_9083);
or U9181 (N_9181,N_9072,N_9076);
and U9182 (N_9182,N_9055,N_9010);
or U9183 (N_9183,N_9008,N_9088);
and U9184 (N_9184,N_9017,N_9042);
and U9185 (N_9185,N_9042,N_9099);
and U9186 (N_9186,N_9088,N_9028);
or U9187 (N_9187,N_9059,N_9023);
and U9188 (N_9188,N_9020,N_9060);
nand U9189 (N_9189,N_9040,N_9008);
and U9190 (N_9190,N_9044,N_9029);
nand U9191 (N_9191,N_9030,N_9020);
nand U9192 (N_9192,N_9049,N_9051);
nor U9193 (N_9193,N_9042,N_9055);
or U9194 (N_9194,N_9031,N_9024);
and U9195 (N_9195,N_9016,N_9095);
nand U9196 (N_9196,N_9047,N_9056);
and U9197 (N_9197,N_9067,N_9031);
xor U9198 (N_9198,N_9031,N_9028);
nor U9199 (N_9199,N_9006,N_9083);
nor U9200 (N_9200,N_9168,N_9194);
xor U9201 (N_9201,N_9122,N_9149);
nand U9202 (N_9202,N_9176,N_9189);
nand U9203 (N_9203,N_9119,N_9187);
nand U9204 (N_9204,N_9184,N_9137);
and U9205 (N_9205,N_9197,N_9144);
nand U9206 (N_9206,N_9132,N_9188);
nand U9207 (N_9207,N_9198,N_9164);
nand U9208 (N_9208,N_9139,N_9131);
and U9209 (N_9209,N_9151,N_9127);
and U9210 (N_9210,N_9104,N_9192);
or U9211 (N_9211,N_9123,N_9160);
nor U9212 (N_9212,N_9113,N_9117);
nor U9213 (N_9213,N_9153,N_9180);
nand U9214 (N_9214,N_9100,N_9102);
and U9215 (N_9215,N_9141,N_9185);
nor U9216 (N_9216,N_9145,N_9173);
nor U9217 (N_9217,N_9165,N_9118);
and U9218 (N_9218,N_9107,N_9142);
nor U9219 (N_9219,N_9106,N_9174);
and U9220 (N_9220,N_9154,N_9163);
nand U9221 (N_9221,N_9179,N_9121);
and U9222 (N_9222,N_9191,N_9186);
or U9223 (N_9223,N_9109,N_9134);
xor U9224 (N_9224,N_9182,N_9148);
nor U9225 (N_9225,N_9167,N_9115);
xor U9226 (N_9226,N_9105,N_9169);
xnor U9227 (N_9227,N_9177,N_9103);
or U9228 (N_9228,N_9124,N_9126);
xor U9229 (N_9229,N_9190,N_9125);
nor U9230 (N_9230,N_9140,N_9158);
xor U9231 (N_9231,N_9120,N_9181);
and U9232 (N_9232,N_9195,N_9112);
nand U9233 (N_9233,N_9150,N_9199);
or U9234 (N_9234,N_9161,N_9111);
or U9235 (N_9235,N_9172,N_9162);
nand U9236 (N_9236,N_9196,N_9101);
and U9237 (N_9237,N_9146,N_9157);
nor U9238 (N_9238,N_9166,N_9170);
nand U9239 (N_9239,N_9155,N_9159);
nand U9240 (N_9240,N_9147,N_9143);
nand U9241 (N_9241,N_9133,N_9114);
or U9242 (N_9242,N_9175,N_9138);
xnor U9243 (N_9243,N_9129,N_9171);
nor U9244 (N_9244,N_9110,N_9108);
and U9245 (N_9245,N_9128,N_9116);
xnor U9246 (N_9246,N_9183,N_9193);
xnor U9247 (N_9247,N_9130,N_9136);
or U9248 (N_9248,N_9135,N_9156);
xnor U9249 (N_9249,N_9178,N_9152);
or U9250 (N_9250,N_9183,N_9116);
nand U9251 (N_9251,N_9160,N_9122);
nor U9252 (N_9252,N_9181,N_9106);
and U9253 (N_9253,N_9199,N_9103);
and U9254 (N_9254,N_9129,N_9167);
and U9255 (N_9255,N_9128,N_9122);
or U9256 (N_9256,N_9166,N_9138);
nand U9257 (N_9257,N_9177,N_9168);
nor U9258 (N_9258,N_9193,N_9157);
xor U9259 (N_9259,N_9193,N_9105);
and U9260 (N_9260,N_9110,N_9153);
nor U9261 (N_9261,N_9110,N_9198);
or U9262 (N_9262,N_9122,N_9123);
xnor U9263 (N_9263,N_9125,N_9170);
or U9264 (N_9264,N_9111,N_9105);
nand U9265 (N_9265,N_9186,N_9166);
nor U9266 (N_9266,N_9144,N_9155);
xor U9267 (N_9267,N_9141,N_9144);
xor U9268 (N_9268,N_9158,N_9150);
nor U9269 (N_9269,N_9120,N_9150);
and U9270 (N_9270,N_9180,N_9170);
xor U9271 (N_9271,N_9181,N_9140);
and U9272 (N_9272,N_9104,N_9133);
or U9273 (N_9273,N_9194,N_9130);
nor U9274 (N_9274,N_9105,N_9107);
nand U9275 (N_9275,N_9137,N_9115);
nand U9276 (N_9276,N_9104,N_9121);
and U9277 (N_9277,N_9113,N_9148);
nand U9278 (N_9278,N_9127,N_9135);
and U9279 (N_9279,N_9178,N_9177);
and U9280 (N_9280,N_9113,N_9115);
nor U9281 (N_9281,N_9148,N_9106);
and U9282 (N_9282,N_9125,N_9198);
nor U9283 (N_9283,N_9131,N_9193);
nor U9284 (N_9284,N_9178,N_9128);
nor U9285 (N_9285,N_9195,N_9191);
and U9286 (N_9286,N_9149,N_9184);
nor U9287 (N_9287,N_9182,N_9115);
nand U9288 (N_9288,N_9165,N_9169);
or U9289 (N_9289,N_9135,N_9104);
and U9290 (N_9290,N_9159,N_9191);
or U9291 (N_9291,N_9151,N_9184);
xor U9292 (N_9292,N_9117,N_9101);
xor U9293 (N_9293,N_9155,N_9162);
and U9294 (N_9294,N_9129,N_9189);
nor U9295 (N_9295,N_9125,N_9143);
nand U9296 (N_9296,N_9158,N_9106);
or U9297 (N_9297,N_9162,N_9109);
or U9298 (N_9298,N_9132,N_9184);
nand U9299 (N_9299,N_9190,N_9195);
nor U9300 (N_9300,N_9201,N_9293);
and U9301 (N_9301,N_9294,N_9275);
nor U9302 (N_9302,N_9258,N_9256);
nor U9303 (N_9303,N_9209,N_9208);
nor U9304 (N_9304,N_9273,N_9265);
or U9305 (N_9305,N_9299,N_9277);
nand U9306 (N_9306,N_9288,N_9251);
nand U9307 (N_9307,N_9284,N_9266);
and U9308 (N_9308,N_9264,N_9255);
xnor U9309 (N_9309,N_9214,N_9263);
or U9310 (N_9310,N_9238,N_9267);
or U9311 (N_9311,N_9272,N_9206);
nand U9312 (N_9312,N_9235,N_9210);
xor U9313 (N_9313,N_9213,N_9205);
nand U9314 (N_9314,N_9260,N_9215);
nor U9315 (N_9315,N_9268,N_9236);
nand U9316 (N_9316,N_9218,N_9229);
and U9317 (N_9317,N_9270,N_9237);
nor U9318 (N_9318,N_9287,N_9249);
and U9319 (N_9319,N_9242,N_9219);
nor U9320 (N_9320,N_9289,N_9217);
and U9321 (N_9321,N_9261,N_9222);
nand U9322 (N_9322,N_9231,N_9274);
xnor U9323 (N_9323,N_9234,N_9281);
xor U9324 (N_9324,N_9250,N_9228);
xnor U9325 (N_9325,N_9241,N_9279);
xor U9326 (N_9326,N_9282,N_9297);
or U9327 (N_9327,N_9292,N_9232);
or U9328 (N_9328,N_9245,N_9204);
or U9329 (N_9329,N_9262,N_9226);
nor U9330 (N_9330,N_9203,N_9247);
nand U9331 (N_9331,N_9295,N_9221);
nor U9332 (N_9332,N_9202,N_9271);
nor U9333 (N_9333,N_9257,N_9216);
or U9334 (N_9334,N_9291,N_9286);
or U9335 (N_9335,N_9246,N_9240);
xnor U9336 (N_9336,N_9296,N_9290);
nor U9337 (N_9337,N_9225,N_9233);
nand U9338 (N_9338,N_9211,N_9276);
xnor U9339 (N_9339,N_9252,N_9244);
and U9340 (N_9340,N_9269,N_9285);
and U9341 (N_9341,N_9254,N_9220);
xor U9342 (N_9342,N_9253,N_9227);
nor U9343 (N_9343,N_9207,N_9230);
xor U9344 (N_9344,N_9212,N_9200);
xnor U9345 (N_9345,N_9224,N_9248);
nand U9346 (N_9346,N_9243,N_9298);
and U9347 (N_9347,N_9223,N_9259);
nand U9348 (N_9348,N_9283,N_9239);
xor U9349 (N_9349,N_9278,N_9280);
xnor U9350 (N_9350,N_9208,N_9286);
nor U9351 (N_9351,N_9205,N_9290);
and U9352 (N_9352,N_9225,N_9281);
and U9353 (N_9353,N_9224,N_9271);
nor U9354 (N_9354,N_9208,N_9257);
xor U9355 (N_9355,N_9244,N_9264);
nand U9356 (N_9356,N_9251,N_9230);
or U9357 (N_9357,N_9260,N_9274);
xor U9358 (N_9358,N_9296,N_9243);
nor U9359 (N_9359,N_9271,N_9258);
nand U9360 (N_9360,N_9238,N_9299);
or U9361 (N_9361,N_9256,N_9222);
nor U9362 (N_9362,N_9248,N_9273);
xor U9363 (N_9363,N_9210,N_9243);
and U9364 (N_9364,N_9215,N_9219);
or U9365 (N_9365,N_9244,N_9204);
or U9366 (N_9366,N_9267,N_9296);
nand U9367 (N_9367,N_9256,N_9271);
nand U9368 (N_9368,N_9209,N_9247);
nor U9369 (N_9369,N_9238,N_9203);
or U9370 (N_9370,N_9270,N_9299);
and U9371 (N_9371,N_9260,N_9227);
or U9372 (N_9372,N_9223,N_9228);
or U9373 (N_9373,N_9279,N_9233);
nand U9374 (N_9374,N_9263,N_9205);
nand U9375 (N_9375,N_9240,N_9293);
or U9376 (N_9376,N_9296,N_9257);
or U9377 (N_9377,N_9255,N_9222);
or U9378 (N_9378,N_9233,N_9221);
nor U9379 (N_9379,N_9278,N_9296);
nand U9380 (N_9380,N_9211,N_9244);
nand U9381 (N_9381,N_9230,N_9274);
nor U9382 (N_9382,N_9298,N_9269);
nand U9383 (N_9383,N_9286,N_9237);
or U9384 (N_9384,N_9253,N_9219);
nand U9385 (N_9385,N_9234,N_9294);
nor U9386 (N_9386,N_9220,N_9203);
or U9387 (N_9387,N_9244,N_9282);
or U9388 (N_9388,N_9274,N_9276);
nor U9389 (N_9389,N_9239,N_9220);
or U9390 (N_9390,N_9259,N_9256);
nand U9391 (N_9391,N_9239,N_9232);
nor U9392 (N_9392,N_9266,N_9246);
or U9393 (N_9393,N_9218,N_9208);
and U9394 (N_9394,N_9232,N_9205);
nor U9395 (N_9395,N_9299,N_9245);
and U9396 (N_9396,N_9284,N_9275);
xnor U9397 (N_9397,N_9221,N_9260);
nand U9398 (N_9398,N_9239,N_9285);
nand U9399 (N_9399,N_9295,N_9230);
or U9400 (N_9400,N_9370,N_9320);
nand U9401 (N_9401,N_9360,N_9399);
nand U9402 (N_9402,N_9343,N_9335);
nand U9403 (N_9403,N_9324,N_9388);
nor U9404 (N_9404,N_9310,N_9323);
xor U9405 (N_9405,N_9303,N_9347);
or U9406 (N_9406,N_9318,N_9352);
nor U9407 (N_9407,N_9336,N_9348);
and U9408 (N_9408,N_9321,N_9357);
or U9409 (N_9409,N_9385,N_9376);
nand U9410 (N_9410,N_9380,N_9314);
xor U9411 (N_9411,N_9389,N_9350);
xnor U9412 (N_9412,N_9308,N_9369);
nand U9413 (N_9413,N_9337,N_9395);
nand U9414 (N_9414,N_9377,N_9306);
nand U9415 (N_9415,N_9382,N_9351);
and U9416 (N_9416,N_9315,N_9309);
or U9417 (N_9417,N_9312,N_9349);
nand U9418 (N_9418,N_9361,N_9331);
nand U9419 (N_9419,N_9301,N_9375);
nor U9420 (N_9420,N_9332,N_9387);
xnor U9421 (N_9421,N_9358,N_9354);
or U9422 (N_9422,N_9355,N_9339);
nand U9423 (N_9423,N_9392,N_9373);
nor U9424 (N_9424,N_9328,N_9304);
xor U9425 (N_9425,N_9364,N_9390);
or U9426 (N_9426,N_9316,N_9397);
nand U9427 (N_9427,N_9341,N_9300);
and U9428 (N_9428,N_9311,N_9384);
and U9429 (N_9429,N_9374,N_9398);
nor U9430 (N_9430,N_9345,N_9359);
or U9431 (N_9431,N_9379,N_9383);
nand U9432 (N_9432,N_9330,N_9307);
nand U9433 (N_9433,N_9366,N_9372);
nor U9434 (N_9434,N_9346,N_9367);
and U9435 (N_9435,N_9326,N_9340);
or U9436 (N_9436,N_9365,N_9342);
nor U9437 (N_9437,N_9302,N_9319);
nand U9438 (N_9438,N_9327,N_9394);
nor U9439 (N_9439,N_9391,N_9325);
and U9440 (N_9440,N_9305,N_9353);
xor U9441 (N_9441,N_9393,N_9362);
or U9442 (N_9442,N_9368,N_9356);
or U9443 (N_9443,N_9333,N_9329);
or U9444 (N_9444,N_9322,N_9344);
nand U9445 (N_9445,N_9386,N_9371);
nand U9446 (N_9446,N_9334,N_9363);
nor U9447 (N_9447,N_9396,N_9317);
or U9448 (N_9448,N_9381,N_9338);
xnor U9449 (N_9449,N_9313,N_9378);
and U9450 (N_9450,N_9353,N_9388);
xnor U9451 (N_9451,N_9368,N_9338);
nor U9452 (N_9452,N_9352,N_9321);
xnor U9453 (N_9453,N_9369,N_9357);
and U9454 (N_9454,N_9358,N_9351);
nor U9455 (N_9455,N_9355,N_9326);
or U9456 (N_9456,N_9324,N_9365);
xor U9457 (N_9457,N_9324,N_9316);
nand U9458 (N_9458,N_9306,N_9330);
and U9459 (N_9459,N_9305,N_9310);
xnor U9460 (N_9460,N_9332,N_9378);
xor U9461 (N_9461,N_9327,N_9376);
nand U9462 (N_9462,N_9350,N_9320);
xor U9463 (N_9463,N_9338,N_9386);
and U9464 (N_9464,N_9314,N_9302);
xor U9465 (N_9465,N_9366,N_9387);
xor U9466 (N_9466,N_9347,N_9353);
or U9467 (N_9467,N_9309,N_9377);
nand U9468 (N_9468,N_9393,N_9303);
nand U9469 (N_9469,N_9362,N_9390);
nand U9470 (N_9470,N_9316,N_9326);
or U9471 (N_9471,N_9358,N_9367);
xnor U9472 (N_9472,N_9309,N_9362);
nor U9473 (N_9473,N_9359,N_9337);
nor U9474 (N_9474,N_9385,N_9398);
or U9475 (N_9475,N_9302,N_9397);
and U9476 (N_9476,N_9322,N_9381);
xnor U9477 (N_9477,N_9300,N_9306);
and U9478 (N_9478,N_9356,N_9300);
nor U9479 (N_9479,N_9335,N_9320);
and U9480 (N_9480,N_9355,N_9386);
nand U9481 (N_9481,N_9307,N_9325);
nand U9482 (N_9482,N_9307,N_9319);
nor U9483 (N_9483,N_9352,N_9327);
nand U9484 (N_9484,N_9300,N_9320);
nand U9485 (N_9485,N_9364,N_9352);
xnor U9486 (N_9486,N_9399,N_9381);
xnor U9487 (N_9487,N_9312,N_9330);
or U9488 (N_9488,N_9343,N_9366);
or U9489 (N_9489,N_9304,N_9390);
xnor U9490 (N_9490,N_9359,N_9339);
or U9491 (N_9491,N_9322,N_9306);
xor U9492 (N_9492,N_9311,N_9389);
nand U9493 (N_9493,N_9346,N_9366);
or U9494 (N_9494,N_9366,N_9392);
nand U9495 (N_9495,N_9322,N_9302);
xnor U9496 (N_9496,N_9394,N_9333);
and U9497 (N_9497,N_9368,N_9315);
nand U9498 (N_9498,N_9373,N_9398);
and U9499 (N_9499,N_9335,N_9321);
xor U9500 (N_9500,N_9461,N_9496);
nor U9501 (N_9501,N_9423,N_9427);
and U9502 (N_9502,N_9419,N_9463);
or U9503 (N_9503,N_9464,N_9462);
xor U9504 (N_9504,N_9403,N_9472);
or U9505 (N_9505,N_9484,N_9418);
xor U9506 (N_9506,N_9465,N_9428);
nor U9507 (N_9507,N_9448,N_9438);
xor U9508 (N_9508,N_9439,N_9412);
nor U9509 (N_9509,N_9410,N_9453);
nand U9510 (N_9510,N_9432,N_9407);
nand U9511 (N_9511,N_9479,N_9493);
xor U9512 (N_9512,N_9422,N_9455);
and U9513 (N_9513,N_9494,N_9430);
or U9514 (N_9514,N_9415,N_9442);
and U9515 (N_9515,N_9478,N_9490);
nand U9516 (N_9516,N_9431,N_9404);
or U9517 (N_9517,N_9483,N_9446);
or U9518 (N_9518,N_9459,N_9454);
and U9519 (N_9519,N_9402,N_9441);
xnor U9520 (N_9520,N_9466,N_9452);
xor U9521 (N_9521,N_9401,N_9495);
and U9522 (N_9522,N_9414,N_9482);
or U9523 (N_9523,N_9409,N_9469);
and U9524 (N_9524,N_9434,N_9429);
nand U9525 (N_9525,N_9498,N_9425);
xor U9526 (N_9526,N_9499,N_9445);
nor U9527 (N_9527,N_9450,N_9477);
xor U9528 (N_9528,N_9421,N_9433);
nand U9529 (N_9529,N_9406,N_9411);
or U9530 (N_9530,N_9485,N_9481);
nand U9531 (N_9531,N_9420,N_9458);
xor U9532 (N_9532,N_9416,N_9475);
nor U9533 (N_9533,N_9460,N_9476);
xor U9534 (N_9534,N_9497,N_9451);
or U9535 (N_9535,N_9413,N_9405);
xnor U9536 (N_9536,N_9488,N_9456);
nor U9537 (N_9537,N_9486,N_9436);
xor U9538 (N_9538,N_9480,N_9449);
or U9539 (N_9539,N_9491,N_9468);
or U9540 (N_9540,N_9408,N_9443);
xnor U9541 (N_9541,N_9489,N_9471);
and U9542 (N_9542,N_9473,N_9424);
nand U9543 (N_9543,N_9457,N_9487);
nand U9544 (N_9544,N_9426,N_9470);
nand U9545 (N_9545,N_9474,N_9444);
nand U9546 (N_9546,N_9492,N_9417);
nand U9547 (N_9547,N_9447,N_9440);
nand U9548 (N_9548,N_9467,N_9435);
xor U9549 (N_9549,N_9400,N_9437);
nand U9550 (N_9550,N_9404,N_9452);
xor U9551 (N_9551,N_9442,N_9457);
nand U9552 (N_9552,N_9420,N_9417);
nor U9553 (N_9553,N_9484,N_9422);
and U9554 (N_9554,N_9487,N_9410);
nor U9555 (N_9555,N_9403,N_9402);
and U9556 (N_9556,N_9425,N_9437);
nand U9557 (N_9557,N_9415,N_9498);
nor U9558 (N_9558,N_9411,N_9423);
xor U9559 (N_9559,N_9441,N_9470);
nor U9560 (N_9560,N_9409,N_9431);
nor U9561 (N_9561,N_9496,N_9407);
xor U9562 (N_9562,N_9483,N_9443);
or U9563 (N_9563,N_9421,N_9475);
nand U9564 (N_9564,N_9436,N_9427);
and U9565 (N_9565,N_9429,N_9482);
xnor U9566 (N_9566,N_9421,N_9483);
nor U9567 (N_9567,N_9451,N_9462);
nor U9568 (N_9568,N_9436,N_9490);
or U9569 (N_9569,N_9406,N_9450);
and U9570 (N_9570,N_9432,N_9420);
xor U9571 (N_9571,N_9491,N_9499);
or U9572 (N_9572,N_9483,N_9425);
xnor U9573 (N_9573,N_9411,N_9460);
xnor U9574 (N_9574,N_9448,N_9405);
and U9575 (N_9575,N_9442,N_9456);
or U9576 (N_9576,N_9407,N_9480);
or U9577 (N_9577,N_9410,N_9440);
or U9578 (N_9578,N_9452,N_9481);
nor U9579 (N_9579,N_9423,N_9430);
or U9580 (N_9580,N_9451,N_9442);
and U9581 (N_9581,N_9447,N_9411);
xnor U9582 (N_9582,N_9402,N_9404);
or U9583 (N_9583,N_9496,N_9457);
nor U9584 (N_9584,N_9484,N_9490);
nor U9585 (N_9585,N_9455,N_9449);
nor U9586 (N_9586,N_9428,N_9436);
and U9587 (N_9587,N_9424,N_9407);
nand U9588 (N_9588,N_9482,N_9464);
and U9589 (N_9589,N_9446,N_9445);
nor U9590 (N_9590,N_9405,N_9463);
and U9591 (N_9591,N_9412,N_9479);
and U9592 (N_9592,N_9455,N_9493);
nand U9593 (N_9593,N_9454,N_9439);
nand U9594 (N_9594,N_9451,N_9403);
nand U9595 (N_9595,N_9497,N_9485);
nor U9596 (N_9596,N_9449,N_9491);
xnor U9597 (N_9597,N_9417,N_9474);
xnor U9598 (N_9598,N_9458,N_9460);
and U9599 (N_9599,N_9438,N_9444);
nand U9600 (N_9600,N_9526,N_9516);
xnor U9601 (N_9601,N_9588,N_9532);
or U9602 (N_9602,N_9552,N_9593);
nand U9603 (N_9603,N_9534,N_9533);
and U9604 (N_9604,N_9539,N_9529);
nor U9605 (N_9605,N_9581,N_9506);
and U9606 (N_9606,N_9551,N_9503);
and U9607 (N_9607,N_9518,N_9510);
and U9608 (N_9608,N_9543,N_9511);
or U9609 (N_9609,N_9571,N_9577);
xnor U9610 (N_9610,N_9512,N_9514);
or U9611 (N_9611,N_9587,N_9542);
xor U9612 (N_9612,N_9523,N_9553);
xor U9613 (N_9613,N_9555,N_9595);
or U9614 (N_9614,N_9508,N_9569);
nand U9615 (N_9615,N_9579,N_9548);
xnor U9616 (N_9616,N_9565,N_9550);
nor U9617 (N_9617,N_9568,N_9504);
and U9618 (N_9618,N_9580,N_9598);
or U9619 (N_9619,N_9599,N_9528);
nand U9620 (N_9620,N_9505,N_9502);
nand U9621 (N_9621,N_9538,N_9583);
xor U9622 (N_9622,N_9540,N_9575);
nand U9623 (N_9623,N_9592,N_9560);
nand U9624 (N_9624,N_9536,N_9544);
or U9625 (N_9625,N_9573,N_9556);
and U9626 (N_9626,N_9578,N_9586);
and U9627 (N_9627,N_9564,N_9576);
xnor U9628 (N_9628,N_9584,N_9527);
nand U9629 (N_9629,N_9525,N_9562);
nand U9630 (N_9630,N_9541,N_9545);
and U9631 (N_9631,N_9517,N_9547);
xnor U9632 (N_9632,N_9561,N_9589);
or U9633 (N_9633,N_9522,N_9554);
or U9634 (N_9634,N_9521,N_9549);
nor U9635 (N_9635,N_9513,N_9524);
and U9636 (N_9636,N_9530,N_9515);
nor U9637 (N_9637,N_9520,N_9563);
and U9638 (N_9638,N_9558,N_9597);
nand U9639 (N_9639,N_9594,N_9596);
nand U9640 (N_9640,N_9590,N_9546);
or U9641 (N_9641,N_9501,N_9591);
and U9642 (N_9642,N_9574,N_9582);
or U9643 (N_9643,N_9570,N_9537);
or U9644 (N_9644,N_9500,N_9559);
nor U9645 (N_9645,N_9535,N_9567);
nand U9646 (N_9646,N_9531,N_9519);
or U9647 (N_9647,N_9566,N_9557);
nand U9648 (N_9648,N_9507,N_9585);
xor U9649 (N_9649,N_9572,N_9509);
nor U9650 (N_9650,N_9551,N_9592);
xnor U9651 (N_9651,N_9534,N_9568);
nor U9652 (N_9652,N_9554,N_9541);
or U9653 (N_9653,N_9566,N_9561);
and U9654 (N_9654,N_9574,N_9567);
nand U9655 (N_9655,N_9586,N_9531);
or U9656 (N_9656,N_9584,N_9500);
or U9657 (N_9657,N_9578,N_9509);
or U9658 (N_9658,N_9530,N_9573);
nor U9659 (N_9659,N_9529,N_9534);
xnor U9660 (N_9660,N_9555,N_9520);
or U9661 (N_9661,N_9569,N_9545);
and U9662 (N_9662,N_9590,N_9535);
xor U9663 (N_9663,N_9589,N_9509);
xnor U9664 (N_9664,N_9569,N_9503);
nor U9665 (N_9665,N_9527,N_9514);
and U9666 (N_9666,N_9525,N_9566);
nor U9667 (N_9667,N_9590,N_9564);
xnor U9668 (N_9668,N_9508,N_9532);
nor U9669 (N_9669,N_9567,N_9508);
nand U9670 (N_9670,N_9556,N_9580);
and U9671 (N_9671,N_9589,N_9593);
nand U9672 (N_9672,N_9512,N_9583);
xor U9673 (N_9673,N_9558,N_9586);
nand U9674 (N_9674,N_9554,N_9567);
nor U9675 (N_9675,N_9577,N_9598);
xnor U9676 (N_9676,N_9554,N_9537);
xor U9677 (N_9677,N_9564,N_9584);
nand U9678 (N_9678,N_9526,N_9562);
nand U9679 (N_9679,N_9571,N_9597);
xnor U9680 (N_9680,N_9588,N_9559);
nor U9681 (N_9681,N_9563,N_9510);
nor U9682 (N_9682,N_9547,N_9597);
and U9683 (N_9683,N_9565,N_9581);
and U9684 (N_9684,N_9565,N_9536);
xor U9685 (N_9685,N_9570,N_9561);
or U9686 (N_9686,N_9533,N_9527);
nor U9687 (N_9687,N_9551,N_9526);
nand U9688 (N_9688,N_9589,N_9550);
nand U9689 (N_9689,N_9526,N_9576);
or U9690 (N_9690,N_9544,N_9519);
nor U9691 (N_9691,N_9595,N_9527);
xnor U9692 (N_9692,N_9528,N_9577);
and U9693 (N_9693,N_9521,N_9591);
and U9694 (N_9694,N_9535,N_9582);
nand U9695 (N_9695,N_9558,N_9594);
and U9696 (N_9696,N_9599,N_9561);
xnor U9697 (N_9697,N_9564,N_9518);
and U9698 (N_9698,N_9531,N_9545);
or U9699 (N_9699,N_9504,N_9566);
and U9700 (N_9700,N_9691,N_9678);
xor U9701 (N_9701,N_9668,N_9633);
xor U9702 (N_9702,N_9663,N_9606);
nor U9703 (N_9703,N_9605,N_9601);
or U9704 (N_9704,N_9620,N_9607);
nor U9705 (N_9705,N_9674,N_9694);
and U9706 (N_9706,N_9635,N_9669);
nand U9707 (N_9707,N_9661,N_9699);
or U9708 (N_9708,N_9617,N_9693);
xor U9709 (N_9709,N_9637,N_9641);
and U9710 (N_9710,N_9632,N_9684);
or U9711 (N_9711,N_9656,N_9628);
xor U9712 (N_9712,N_9638,N_9697);
and U9713 (N_9713,N_9631,N_9615);
or U9714 (N_9714,N_9680,N_9683);
xnor U9715 (N_9715,N_9686,N_9621);
and U9716 (N_9716,N_9640,N_9630);
and U9717 (N_9717,N_9653,N_9658);
or U9718 (N_9718,N_9650,N_9657);
nor U9719 (N_9719,N_9698,N_9647);
and U9720 (N_9720,N_9660,N_9609);
xor U9721 (N_9721,N_9665,N_9692);
xor U9722 (N_9722,N_9625,N_9624);
and U9723 (N_9723,N_9616,N_9600);
and U9724 (N_9724,N_9652,N_9689);
and U9725 (N_9725,N_9672,N_9618);
nand U9726 (N_9726,N_9690,N_9648);
and U9727 (N_9727,N_9627,N_9671);
nand U9728 (N_9728,N_9626,N_9612);
xor U9729 (N_9729,N_9646,N_9610);
and U9730 (N_9730,N_9682,N_9695);
nor U9731 (N_9731,N_9611,N_9654);
xor U9732 (N_9732,N_9666,N_9645);
nand U9733 (N_9733,N_9613,N_9634);
nor U9734 (N_9734,N_9670,N_9614);
nor U9735 (N_9735,N_9679,N_9623);
and U9736 (N_9736,N_9677,N_9619);
nand U9737 (N_9737,N_9636,N_9696);
or U9738 (N_9738,N_9659,N_9655);
nand U9739 (N_9739,N_9673,N_9608);
nand U9740 (N_9740,N_9667,N_9643);
or U9741 (N_9741,N_9651,N_9642);
nand U9742 (N_9742,N_9687,N_9675);
and U9743 (N_9743,N_9662,N_9676);
nor U9744 (N_9744,N_9681,N_9644);
or U9745 (N_9745,N_9664,N_9603);
xnor U9746 (N_9746,N_9622,N_9649);
nand U9747 (N_9747,N_9639,N_9604);
or U9748 (N_9748,N_9688,N_9602);
nor U9749 (N_9749,N_9629,N_9685);
xnor U9750 (N_9750,N_9686,N_9666);
and U9751 (N_9751,N_9661,N_9630);
nor U9752 (N_9752,N_9656,N_9669);
xor U9753 (N_9753,N_9619,N_9689);
and U9754 (N_9754,N_9671,N_9620);
nand U9755 (N_9755,N_9696,N_9628);
xor U9756 (N_9756,N_9629,N_9633);
or U9757 (N_9757,N_9600,N_9671);
or U9758 (N_9758,N_9670,N_9684);
and U9759 (N_9759,N_9648,N_9663);
or U9760 (N_9760,N_9673,N_9604);
or U9761 (N_9761,N_9699,N_9616);
nor U9762 (N_9762,N_9642,N_9671);
nand U9763 (N_9763,N_9638,N_9685);
or U9764 (N_9764,N_9604,N_9647);
and U9765 (N_9765,N_9676,N_9620);
xnor U9766 (N_9766,N_9640,N_9654);
or U9767 (N_9767,N_9651,N_9692);
nor U9768 (N_9768,N_9639,N_9642);
xnor U9769 (N_9769,N_9672,N_9633);
nand U9770 (N_9770,N_9681,N_9663);
or U9771 (N_9771,N_9602,N_9687);
xor U9772 (N_9772,N_9695,N_9648);
xnor U9773 (N_9773,N_9650,N_9639);
xor U9774 (N_9774,N_9661,N_9684);
xor U9775 (N_9775,N_9601,N_9619);
nand U9776 (N_9776,N_9603,N_9670);
and U9777 (N_9777,N_9696,N_9659);
and U9778 (N_9778,N_9693,N_9673);
nor U9779 (N_9779,N_9609,N_9641);
nor U9780 (N_9780,N_9690,N_9646);
or U9781 (N_9781,N_9680,N_9687);
nand U9782 (N_9782,N_9633,N_9686);
and U9783 (N_9783,N_9697,N_9621);
nor U9784 (N_9784,N_9673,N_9633);
and U9785 (N_9785,N_9642,N_9676);
nor U9786 (N_9786,N_9669,N_9619);
xor U9787 (N_9787,N_9621,N_9636);
nand U9788 (N_9788,N_9685,N_9613);
and U9789 (N_9789,N_9601,N_9661);
or U9790 (N_9790,N_9657,N_9614);
nor U9791 (N_9791,N_9695,N_9628);
or U9792 (N_9792,N_9681,N_9635);
nor U9793 (N_9793,N_9611,N_9623);
and U9794 (N_9794,N_9605,N_9632);
xnor U9795 (N_9795,N_9626,N_9618);
xor U9796 (N_9796,N_9629,N_9660);
or U9797 (N_9797,N_9618,N_9678);
xnor U9798 (N_9798,N_9654,N_9645);
nor U9799 (N_9799,N_9640,N_9611);
nand U9800 (N_9800,N_9784,N_9710);
or U9801 (N_9801,N_9776,N_9763);
nand U9802 (N_9802,N_9709,N_9798);
and U9803 (N_9803,N_9769,N_9713);
nand U9804 (N_9804,N_9797,N_9706);
and U9805 (N_9805,N_9701,N_9793);
or U9806 (N_9806,N_9745,N_9748);
nor U9807 (N_9807,N_9747,N_9773);
and U9808 (N_9808,N_9762,N_9730);
or U9809 (N_9809,N_9708,N_9724);
xnor U9810 (N_9810,N_9765,N_9744);
and U9811 (N_9811,N_9759,N_9772);
or U9812 (N_9812,N_9790,N_9742);
or U9813 (N_9813,N_9796,N_9782);
nand U9814 (N_9814,N_9729,N_9707);
nor U9815 (N_9815,N_9780,N_9743);
nor U9816 (N_9816,N_9733,N_9702);
or U9817 (N_9817,N_9716,N_9768);
or U9818 (N_9818,N_9771,N_9705);
nand U9819 (N_9819,N_9767,N_9720);
nand U9820 (N_9820,N_9766,N_9718);
xnor U9821 (N_9821,N_9726,N_9789);
xor U9822 (N_9822,N_9794,N_9755);
and U9823 (N_9823,N_9750,N_9722);
nor U9824 (N_9824,N_9736,N_9731);
nor U9825 (N_9825,N_9787,N_9727);
or U9826 (N_9826,N_9712,N_9764);
or U9827 (N_9827,N_9711,N_9740);
nor U9828 (N_9828,N_9781,N_9786);
nand U9829 (N_9829,N_9778,N_9717);
nor U9830 (N_9830,N_9751,N_9785);
xor U9831 (N_9831,N_9775,N_9715);
nand U9832 (N_9832,N_9704,N_9719);
nand U9833 (N_9833,N_9760,N_9774);
and U9834 (N_9834,N_9737,N_9728);
nand U9835 (N_9835,N_9777,N_9741);
nor U9836 (N_9836,N_9700,N_9757);
or U9837 (N_9837,N_9792,N_9732);
xnor U9838 (N_9838,N_9738,N_9753);
nor U9839 (N_9839,N_9788,N_9783);
nand U9840 (N_9840,N_9734,N_9749);
nor U9841 (N_9841,N_9735,N_9703);
nand U9842 (N_9842,N_9791,N_9725);
xor U9843 (N_9843,N_9714,N_9723);
or U9844 (N_9844,N_9746,N_9795);
nor U9845 (N_9845,N_9779,N_9721);
nand U9846 (N_9846,N_9770,N_9761);
nand U9847 (N_9847,N_9756,N_9752);
xor U9848 (N_9848,N_9799,N_9758);
xnor U9849 (N_9849,N_9739,N_9754);
nand U9850 (N_9850,N_9777,N_9739);
nor U9851 (N_9851,N_9751,N_9722);
nand U9852 (N_9852,N_9724,N_9789);
nor U9853 (N_9853,N_9702,N_9763);
and U9854 (N_9854,N_9737,N_9740);
nor U9855 (N_9855,N_9798,N_9727);
nand U9856 (N_9856,N_9717,N_9752);
or U9857 (N_9857,N_9765,N_9771);
nor U9858 (N_9858,N_9764,N_9714);
or U9859 (N_9859,N_9748,N_9765);
xnor U9860 (N_9860,N_9797,N_9705);
or U9861 (N_9861,N_9703,N_9776);
and U9862 (N_9862,N_9720,N_9731);
or U9863 (N_9863,N_9733,N_9756);
xor U9864 (N_9864,N_9785,N_9718);
nor U9865 (N_9865,N_9754,N_9770);
and U9866 (N_9866,N_9739,N_9741);
and U9867 (N_9867,N_9752,N_9788);
nor U9868 (N_9868,N_9798,N_9783);
and U9869 (N_9869,N_9785,N_9779);
nor U9870 (N_9870,N_9704,N_9770);
nor U9871 (N_9871,N_9773,N_9735);
xor U9872 (N_9872,N_9768,N_9744);
xor U9873 (N_9873,N_9727,N_9732);
or U9874 (N_9874,N_9747,N_9714);
xnor U9875 (N_9875,N_9749,N_9716);
xor U9876 (N_9876,N_9710,N_9767);
or U9877 (N_9877,N_9788,N_9772);
or U9878 (N_9878,N_9765,N_9766);
nor U9879 (N_9879,N_9781,N_9768);
and U9880 (N_9880,N_9791,N_9723);
or U9881 (N_9881,N_9707,N_9782);
or U9882 (N_9882,N_9752,N_9712);
and U9883 (N_9883,N_9795,N_9798);
or U9884 (N_9884,N_9752,N_9736);
nand U9885 (N_9885,N_9701,N_9757);
or U9886 (N_9886,N_9770,N_9701);
xor U9887 (N_9887,N_9752,N_9760);
xnor U9888 (N_9888,N_9758,N_9752);
nor U9889 (N_9889,N_9770,N_9741);
xnor U9890 (N_9890,N_9777,N_9798);
or U9891 (N_9891,N_9737,N_9765);
and U9892 (N_9892,N_9701,N_9719);
and U9893 (N_9893,N_9718,N_9757);
nand U9894 (N_9894,N_9794,N_9730);
or U9895 (N_9895,N_9744,N_9722);
nand U9896 (N_9896,N_9739,N_9727);
and U9897 (N_9897,N_9766,N_9797);
xnor U9898 (N_9898,N_9791,N_9753);
nor U9899 (N_9899,N_9739,N_9756);
nor U9900 (N_9900,N_9826,N_9813);
or U9901 (N_9901,N_9855,N_9859);
and U9902 (N_9902,N_9882,N_9806);
or U9903 (N_9903,N_9839,N_9866);
nand U9904 (N_9904,N_9848,N_9876);
nor U9905 (N_9905,N_9886,N_9893);
nand U9906 (N_9906,N_9894,N_9858);
nand U9907 (N_9907,N_9879,N_9849);
xor U9908 (N_9908,N_9843,N_9804);
and U9909 (N_9909,N_9825,N_9851);
or U9910 (N_9910,N_9836,N_9892);
nor U9911 (N_9911,N_9885,N_9824);
xnor U9912 (N_9912,N_9829,N_9878);
or U9913 (N_9913,N_9842,N_9846);
xor U9914 (N_9914,N_9820,N_9823);
or U9915 (N_9915,N_9898,N_9850);
and U9916 (N_9916,N_9840,N_9800);
nor U9917 (N_9917,N_9887,N_9870);
and U9918 (N_9918,N_9828,N_9812);
nor U9919 (N_9919,N_9809,N_9830);
or U9920 (N_9920,N_9897,N_9890);
or U9921 (N_9921,N_9872,N_9854);
and U9922 (N_9922,N_9873,N_9807);
and U9923 (N_9923,N_9853,N_9803);
nor U9924 (N_9924,N_9875,N_9860);
nand U9925 (N_9925,N_9847,N_9883);
xor U9926 (N_9926,N_9844,N_9838);
or U9927 (N_9927,N_9896,N_9817);
nand U9928 (N_9928,N_9895,N_9862);
nor U9929 (N_9929,N_9899,N_9880);
xnor U9930 (N_9930,N_9871,N_9877);
and U9931 (N_9931,N_9864,N_9827);
nor U9932 (N_9932,N_9884,N_9816);
and U9933 (N_9933,N_9834,N_9808);
or U9934 (N_9934,N_9841,N_9865);
or U9935 (N_9935,N_9881,N_9863);
nand U9936 (N_9936,N_9837,N_9822);
nor U9937 (N_9937,N_9819,N_9891);
nor U9938 (N_9938,N_9889,N_9801);
nand U9939 (N_9939,N_9856,N_9821);
nor U9940 (N_9940,N_9861,N_9869);
xor U9941 (N_9941,N_9832,N_9852);
and U9942 (N_9942,N_9874,N_9805);
and U9943 (N_9943,N_9818,N_9835);
nor U9944 (N_9944,N_9810,N_9811);
nand U9945 (N_9945,N_9857,N_9831);
nand U9946 (N_9946,N_9802,N_9845);
xor U9947 (N_9947,N_9868,N_9833);
xnor U9948 (N_9948,N_9867,N_9888);
nand U9949 (N_9949,N_9815,N_9814);
or U9950 (N_9950,N_9820,N_9853);
and U9951 (N_9951,N_9894,N_9860);
or U9952 (N_9952,N_9860,N_9848);
or U9953 (N_9953,N_9816,N_9865);
and U9954 (N_9954,N_9892,N_9823);
nand U9955 (N_9955,N_9846,N_9838);
and U9956 (N_9956,N_9899,N_9877);
nor U9957 (N_9957,N_9821,N_9877);
nand U9958 (N_9958,N_9850,N_9858);
nor U9959 (N_9959,N_9858,N_9842);
nand U9960 (N_9960,N_9824,N_9823);
xor U9961 (N_9961,N_9803,N_9854);
and U9962 (N_9962,N_9883,N_9832);
or U9963 (N_9963,N_9804,N_9870);
or U9964 (N_9964,N_9819,N_9854);
nand U9965 (N_9965,N_9899,N_9839);
nor U9966 (N_9966,N_9806,N_9860);
nand U9967 (N_9967,N_9894,N_9869);
and U9968 (N_9968,N_9889,N_9838);
xnor U9969 (N_9969,N_9829,N_9846);
and U9970 (N_9970,N_9846,N_9870);
xor U9971 (N_9971,N_9835,N_9800);
nor U9972 (N_9972,N_9838,N_9823);
or U9973 (N_9973,N_9898,N_9832);
and U9974 (N_9974,N_9844,N_9882);
xor U9975 (N_9975,N_9817,N_9825);
nand U9976 (N_9976,N_9813,N_9886);
xor U9977 (N_9977,N_9888,N_9829);
xnor U9978 (N_9978,N_9899,N_9859);
nand U9979 (N_9979,N_9818,N_9810);
and U9980 (N_9980,N_9889,N_9850);
xor U9981 (N_9981,N_9829,N_9850);
and U9982 (N_9982,N_9875,N_9881);
xnor U9983 (N_9983,N_9810,N_9886);
nor U9984 (N_9984,N_9836,N_9802);
or U9985 (N_9985,N_9835,N_9881);
and U9986 (N_9986,N_9833,N_9888);
or U9987 (N_9987,N_9894,N_9812);
nand U9988 (N_9988,N_9880,N_9892);
xnor U9989 (N_9989,N_9837,N_9804);
nand U9990 (N_9990,N_9886,N_9802);
nor U9991 (N_9991,N_9889,N_9895);
xor U9992 (N_9992,N_9863,N_9870);
nand U9993 (N_9993,N_9805,N_9884);
xor U9994 (N_9994,N_9897,N_9837);
xor U9995 (N_9995,N_9892,N_9886);
and U9996 (N_9996,N_9846,N_9875);
nand U9997 (N_9997,N_9810,N_9877);
xnor U9998 (N_9998,N_9877,N_9819);
nor U9999 (N_9999,N_9821,N_9836);
and UO_0 (O_0,N_9906,N_9931);
and UO_1 (O_1,N_9930,N_9979);
nand UO_2 (O_2,N_9919,N_9985);
xnor UO_3 (O_3,N_9972,N_9968);
xor UO_4 (O_4,N_9993,N_9937);
or UO_5 (O_5,N_9922,N_9923);
nand UO_6 (O_6,N_9996,N_9916);
xor UO_7 (O_7,N_9986,N_9984);
xnor UO_8 (O_8,N_9947,N_9920);
nand UO_9 (O_9,N_9904,N_9955);
xor UO_10 (O_10,N_9949,N_9981);
nor UO_11 (O_11,N_9946,N_9905);
or UO_12 (O_12,N_9969,N_9913);
nand UO_13 (O_13,N_9957,N_9990);
and UO_14 (O_14,N_9974,N_9907);
nand UO_15 (O_15,N_9939,N_9938);
and UO_16 (O_16,N_9911,N_9978);
nor UO_17 (O_17,N_9940,N_9964);
or UO_18 (O_18,N_9901,N_9970);
nand UO_19 (O_19,N_9991,N_9954);
nand UO_20 (O_20,N_9988,N_9925);
and UO_21 (O_21,N_9951,N_9944);
or UO_22 (O_22,N_9932,N_9997);
and UO_23 (O_23,N_9953,N_9921);
or UO_24 (O_24,N_9983,N_9914);
xnor UO_25 (O_25,N_9987,N_9994);
nor UO_26 (O_26,N_9965,N_9910);
nor UO_27 (O_27,N_9924,N_9902);
nor UO_28 (O_28,N_9927,N_9963);
or UO_29 (O_29,N_9950,N_9948);
and UO_30 (O_30,N_9918,N_9973);
xor UO_31 (O_31,N_9915,N_9917);
xnor UO_32 (O_32,N_9941,N_9958);
or UO_33 (O_33,N_9943,N_9945);
and UO_34 (O_34,N_9912,N_9929);
xnor UO_35 (O_35,N_9909,N_9962);
nor UO_36 (O_36,N_9980,N_9976);
nand UO_37 (O_37,N_9933,N_9935);
nand UO_38 (O_38,N_9959,N_9975);
nand UO_39 (O_39,N_9998,N_9982);
or UO_40 (O_40,N_9961,N_9926);
nand UO_41 (O_41,N_9995,N_9900);
and UO_42 (O_42,N_9971,N_9999);
nor UO_43 (O_43,N_9992,N_9977);
nand UO_44 (O_44,N_9966,N_9967);
and UO_45 (O_45,N_9956,N_9934);
and UO_46 (O_46,N_9960,N_9908);
nand UO_47 (O_47,N_9903,N_9952);
and UO_48 (O_48,N_9936,N_9989);
nand UO_49 (O_49,N_9942,N_9928);
nor UO_50 (O_50,N_9948,N_9911);
xor UO_51 (O_51,N_9998,N_9902);
or UO_52 (O_52,N_9986,N_9911);
or UO_53 (O_53,N_9974,N_9979);
nand UO_54 (O_54,N_9974,N_9968);
nor UO_55 (O_55,N_9948,N_9964);
nor UO_56 (O_56,N_9922,N_9967);
xnor UO_57 (O_57,N_9918,N_9952);
nand UO_58 (O_58,N_9980,N_9958);
xor UO_59 (O_59,N_9910,N_9932);
nor UO_60 (O_60,N_9996,N_9977);
nor UO_61 (O_61,N_9990,N_9986);
nand UO_62 (O_62,N_9952,N_9962);
nand UO_63 (O_63,N_9978,N_9924);
nand UO_64 (O_64,N_9995,N_9904);
nor UO_65 (O_65,N_9938,N_9900);
or UO_66 (O_66,N_9957,N_9925);
nand UO_67 (O_67,N_9912,N_9963);
nand UO_68 (O_68,N_9919,N_9927);
nand UO_69 (O_69,N_9954,N_9988);
or UO_70 (O_70,N_9957,N_9999);
nor UO_71 (O_71,N_9915,N_9987);
nand UO_72 (O_72,N_9901,N_9977);
nor UO_73 (O_73,N_9963,N_9929);
nor UO_74 (O_74,N_9972,N_9979);
and UO_75 (O_75,N_9917,N_9941);
or UO_76 (O_76,N_9957,N_9946);
nor UO_77 (O_77,N_9978,N_9920);
xnor UO_78 (O_78,N_9906,N_9989);
nor UO_79 (O_79,N_9958,N_9984);
nor UO_80 (O_80,N_9948,N_9966);
or UO_81 (O_81,N_9968,N_9919);
or UO_82 (O_82,N_9907,N_9928);
nand UO_83 (O_83,N_9930,N_9923);
or UO_84 (O_84,N_9916,N_9921);
nor UO_85 (O_85,N_9975,N_9941);
xnor UO_86 (O_86,N_9944,N_9927);
xnor UO_87 (O_87,N_9994,N_9938);
nor UO_88 (O_88,N_9954,N_9916);
xnor UO_89 (O_89,N_9969,N_9995);
nand UO_90 (O_90,N_9986,N_9941);
and UO_91 (O_91,N_9924,N_9986);
nor UO_92 (O_92,N_9985,N_9933);
xor UO_93 (O_93,N_9982,N_9904);
nor UO_94 (O_94,N_9969,N_9937);
or UO_95 (O_95,N_9965,N_9908);
and UO_96 (O_96,N_9910,N_9916);
nand UO_97 (O_97,N_9987,N_9904);
nand UO_98 (O_98,N_9963,N_9990);
or UO_99 (O_99,N_9949,N_9956);
nand UO_100 (O_100,N_9993,N_9964);
nor UO_101 (O_101,N_9918,N_9903);
and UO_102 (O_102,N_9955,N_9980);
and UO_103 (O_103,N_9928,N_9981);
nand UO_104 (O_104,N_9974,N_9913);
and UO_105 (O_105,N_9998,N_9920);
or UO_106 (O_106,N_9945,N_9928);
nand UO_107 (O_107,N_9982,N_9905);
nor UO_108 (O_108,N_9925,N_9920);
nand UO_109 (O_109,N_9979,N_9926);
or UO_110 (O_110,N_9987,N_9909);
nand UO_111 (O_111,N_9937,N_9900);
xnor UO_112 (O_112,N_9965,N_9937);
xnor UO_113 (O_113,N_9981,N_9960);
xor UO_114 (O_114,N_9998,N_9917);
nand UO_115 (O_115,N_9999,N_9944);
xor UO_116 (O_116,N_9965,N_9964);
xor UO_117 (O_117,N_9907,N_9982);
and UO_118 (O_118,N_9965,N_9935);
xnor UO_119 (O_119,N_9942,N_9903);
nor UO_120 (O_120,N_9934,N_9965);
nor UO_121 (O_121,N_9997,N_9907);
nor UO_122 (O_122,N_9970,N_9986);
nand UO_123 (O_123,N_9959,N_9914);
and UO_124 (O_124,N_9915,N_9927);
nand UO_125 (O_125,N_9973,N_9912);
nand UO_126 (O_126,N_9904,N_9921);
or UO_127 (O_127,N_9916,N_9969);
nand UO_128 (O_128,N_9905,N_9976);
nand UO_129 (O_129,N_9956,N_9913);
nor UO_130 (O_130,N_9920,N_9904);
or UO_131 (O_131,N_9986,N_9989);
or UO_132 (O_132,N_9991,N_9949);
nand UO_133 (O_133,N_9938,N_9910);
nor UO_134 (O_134,N_9986,N_9966);
and UO_135 (O_135,N_9909,N_9929);
nor UO_136 (O_136,N_9961,N_9998);
and UO_137 (O_137,N_9954,N_9911);
and UO_138 (O_138,N_9926,N_9983);
and UO_139 (O_139,N_9907,N_9993);
or UO_140 (O_140,N_9957,N_9904);
and UO_141 (O_141,N_9940,N_9937);
or UO_142 (O_142,N_9985,N_9978);
or UO_143 (O_143,N_9901,N_9962);
nand UO_144 (O_144,N_9990,N_9927);
nand UO_145 (O_145,N_9977,N_9943);
and UO_146 (O_146,N_9949,N_9953);
xor UO_147 (O_147,N_9955,N_9916);
xor UO_148 (O_148,N_9963,N_9940);
and UO_149 (O_149,N_9921,N_9919);
nor UO_150 (O_150,N_9988,N_9910);
nand UO_151 (O_151,N_9922,N_9980);
nand UO_152 (O_152,N_9908,N_9984);
or UO_153 (O_153,N_9940,N_9987);
xnor UO_154 (O_154,N_9931,N_9965);
xnor UO_155 (O_155,N_9914,N_9943);
nor UO_156 (O_156,N_9916,N_9911);
xor UO_157 (O_157,N_9941,N_9998);
nor UO_158 (O_158,N_9925,N_9934);
or UO_159 (O_159,N_9995,N_9980);
nand UO_160 (O_160,N_9987,N_9947);
or UO_161 (O_161,N_9911,N_9909);
or UO_162 (O_162,N_9918,N_9999);
nand UO_163 (O_163,N_9983,N_9903);
nor UO_164 (O_164,N_9917,N_9928);
nor UO_165 (O_165,N_9927,N_9971);
xnor UO_166 (O_166,N_9965,N_9976);
or UO_167 (O_167,N_9985,N_9971);
nor UO_168 (O_168,N_9956,N_9968);
and UO_169 (O_169,N_9995,N_9917);
and UO_170 (O_170,N_9906,N_9916);
and UO_171 (O_171,N_9903,N_9981);
nor UO_172 (O_172,N_9970,N_9916);
and UO_173 (O_173,N_9953,N_9936);
nand UO_174 (O_174,N_9922,N_9979);
and UO_175 (O_175,N_9982,N_9976);
xnor UO_176 (O_176,N_9925,N_9937);
or UO_177 (O_177,N_9923,N_9920);
or UO_178 (O_178,N_9908,N_9919);
and UO_179 (O_179,N_9904,N_9949);
nand UO_180 (O_180,N_9900,N_9912);
nand UO_181 (O_181,N_9940,N_9984);
or UO_182 (O_182,N_9930,N_9966);
xor UO_183 (O_183,N_9988,N_9960);
xor UO_184 (O_184,N_9964,N_9929);
nor UO_185 (O_185,N_9953,N_9911);
nor UO_186 (O_186,N_9948,N_9919);
nor UO_187 (O_187,N_9901,N_9921);
xnor UO_188 (O_188,N_9963,N_9956);
nand UO_189 (O_189,N_9996,N_9991);
or UO_190 (O_190,N_9982,N_9949);
nor UO_191 (O_191,N_9971,N_9944);
or UO_192 (O_192,N_9900,N_9959);
and UO_193 (O_193,N_9948,N_9977);
xnor UO_194 (O_194,N_9920,N_9960);
or UO_195 (O_195,N_9999,N_9964);
or UO_196 (O_196,N_9914,N_9906);
and UO_197 (O_197,N_9984,N_9930);
nand UO_198 (O_198,N_9959,N_9984);
and UO_199 (O_199,N_9934,N_9916);
and UO_200 (O_200,N_9905,N_9930);
nor UO_201 (O_201,N_9994,N_9988);
xnor UO_202 (O_202,N_9964,N_9944);
nand UO_203 (O_203,N_9998,N_9925);
nor UO_204 (O_204,N_9956,N_9998);
nor UO_205 (O_205,N_9926,N_9987);
nand UO_206 (O_206,N_9957,N_9964);
xnor UO_207 (O_207,N_9961,N_9902);
and UO_208 (O_208,N_9979,N_9962);
xor UO_209 (O_209,N_9974,N_9923);
xnor UO_210 (O_210,N_9997,N_9943);
or UO_211 (O_211,N_9943,N_9907);
nand UO_212 (O_212,N_9947,N_9980);
nor UO_213 (O_213,N_9949,N_9995);
and UO_214 (O_214,N_9989,N_9909);
and UO_215 (O_215,N_9900,N_9934);
nand UO_216 (O_216,N_9949,N_9974);
or UO_217 (O_217,N_9966,N_9957);
nand UO_218 (O_218,N_9926,N_9995);
xor UO_219 (O_219,N_9911,N_9922);
xnor UO_220 (O_220,N_9944,N_9941);
nand UO_221 (O_221,N_9908,N_9917);
xor UO_222 (O_222,N_9914,N_9928);
nor UO_223 (O_223,N_9914,N_9947);
and UO_224 (O_224,N_9909,N_9900);
nand UO_225 (O_225,N_9987,N_9957);
or UO_226 (O_226,N_9976,N_9988);
nand UO_227 (O_227,N_9977,N_9937);
nor UO_228 (O_228,N_9906,N_9956);
xnor UO_229 (O_229,N_9945,N_9950);
xnor UO_230 (O_230,N_9948,N_9903);
xor UO_231 (O_231,N_9938,N_9941);
nand UO_232 (O_232,N_9945,N_9994);
nor UO_233 (O_233,N_9971,N_9925);
nand UO_234 (O_234,N_9967,N_9992);
or UO_235 (O_235,N_9979,N_9997);
xnor UO_236 (O_236,N_9900,N_9955);
xnor UO_237 (O_237,N_9957,N_9986);
xnor UO_238 (O_238,N_9946,N_9903);
and UO_239 (O_239,N_9990,N_9991);
nand UO_240 (O_240,N_9905,N_9965);
nor UO_241 (O_241,N_9956,N_9938);
or UO_242 (O_242,N_9951,N_9957);
nand UO_243 (O_243,N_9984,N_9914);
nor UO_244 (O_244,N_9980,N_9966);
and UO_245 (O_245,N_9998,N_9957);
nand UO_246 (O_246,N_9918,N_9990);
nand UO_247 (O_247,N_9922,N_9931);
nand UO_248 (O_248,N_9934,N_9983);
nand UO_249 (O_249,N_9996,N_9903);
xor UO_250 (O_250,N_9953,N_9904);
and UO_251 (O_251,N_9920,N_9967);
nor UO_252 (O_252,N_9992,N_9914);
nand UO_253 (O_253,N_9960,N_9986);
nor UO_254 (O_254,N_9992,N_9903);
or UO_255 (O_255,N_9994,N_9943);
nand UO_256 (O_256,N_9928,N_9910);
or UO_257 (O_257,N_9915,N_9956);
nand UO_258 (O_258,N_9937,N_9902);
nor UO_259 (O_259,N_9970,N_9980);
and UO_260 (O_260,N_9991,N_9911);
nor UO_261 (O_261,N_9961,N_9976);
or UO_262 (O_262,N_9984,N_9966);
and UO_263 (O_263,N_9982,N_9967);
nor UO_264 (O_264,N_9963,N_9920);
or UO_265 (O_265,N_9938,N_9954);
or UO_266 (O_266,N_9976,N_9955);
and UO_267 (O_267,N_9938,N_9907);
or UO_268 (O_268,N_9949,N_9986);
xor UO_269 (O_269,N_9939,N_9906);
xor UO_270 (O_270,N_9970,N_9945);
and UO_271 (O_271,N_9913,N_9948);
and UO_272 (O_272,N_9966,N_9931);
xor UO_273 (O_273,N_9996,N_9953);
and UO_274 (O_274,N_9984,N_9916);
nor UO_275 (O_275,N_9949,N_9933);
or UO_276 (O_276,N_9966,N_9999);
and UO_277 (O_277,N_9904,N_9906);
nand UO_278 (O_278,N_9973,N_9925);
nand UO_279 (O_279,N_9938,N_9975);
or UO_280 (O_280,N_9978,N_9990);
xnor UO_281 (O_281,N_9941,N_9900);
nand UO_282 (O_282,N_9925,N_9981);
nand UO_283 (O_283,N_9933,N_9937);
or UO_284 (O_284,N_9987,N_9929);
xor UO_285 (O_285,N_9938,N_9903);
nand UO_286 (O_286,N_9927,N_9928);
nand UO_287 (O_287,N_9954,N_9964);
or UO_288 (O_288,N_9996,N_9959);
nor UO_289 (O_289,N_9960,N_9905);
nor UO_290 (O_290,N_9955,N_9961);
and UO_291 (O_291,N_9957,N_9934);
xor UO_292 (O_292,N_9999,N_9934);
nand UO_293 (O_293,N_9949,N_9960);
xnor UO_294 (O_294,N_9938,N_9961);
xnor UO_295 (O_295,N_9980,N_9986);
or UO_296 (O_296,N_9969,N_9997);
or UO_297 (O_297,N_9962,N_9914);
or UO_298 (O_298,N_9915,N_9990);
or UO_299 (O_299,N_9900,N_9965);
or UO_300 (O_300,N_9944,N_9931);
xor UO_301 (O_301,N_9975,N_9900);
and UO_302 (O_302,N_9968,N_9991);
or UO_303 (O_303,N_9940,N_9925);
nor UO_304 (O_304,N_9924,N_9953);
nor UO_305 (O_305,N_9933,N_9926);
nand UO_306 (O_306,N_9938,N_9984);
xor UO_307 (O_307,N_9909,N_9971);
nor UO_308 (O_308,N_9958,N_9957);
xor UO_309 (O_309,N_9934,N_9980);
nand UO_310 (O_310,N_9948,N_9901);
xor UO_311 (O_311,N_9924,N_9960);
nand UO_312 (O_312,N_9977,N_9900);
nor UO_313 (O_313,N_9930,N_9998);
or UO_314 (O_314,N_9955,N_9928);
or UO_315 (O_315,N_9934,N_9990);
xnor UO_316 (O_316,N_9991,N_9938);
nor UO_317 (O_317,N_9959,N_9934);
or UO_318 (O_318,N_9905,N_9919);
or UO_319 (O_319,N_9973,N_9926);
nand UO_320 (O_320,N_9928,N_9930);
and UO_321 (O_321,N_9927,N_9966);
xnor UO_322 (O_322,N_9991,N_9921);
and UO_323 (O_323,N_9984,N_9952);
xor UO_324 (O_324,N_9946,N_9988);
nor UO_325 (O_325,N_9932,N_9900);
and UO_326 (O_326,N_9925,N_9975);
xnor UO_327 (O_327,N_9999,N_9960);
nor UO_328 (O_328,N_9907,N_9905);
and UO_329 (O_329,N_9902,N_9971);
nand UO_330 (O_330,N_9904,N_9924);
or UO_331 (O_331,N_9944,N_9915);
nor UO_332 (O_332,N_9928,N_9939);
nand UO_333 (O_333,N_9997,N_9992);
xor UO_334 (O_334,N_9944,N_9972);
xor UO_335 (O_335,N_9999,N_9969);
and UO_336 (O_336,N_9941,N_9914);
xnor UO_337 (O_337,N_9960,N_9902);
or UO_338 (O_338,N_9900,N_9907);
and UO_339 (O_339,N_9980,N_9900);
nand UO_340 (O_340,N_9941,N_9963);
and UO_341 (O_341,N_9956,N_9933);
nor UO_342 (O_342,N_9995,N_9941);
xnor UO_343 (O_343,N_9994,N_9971);
xor UO_344 (O_344,N_9916,N_9994);
and UO_345 (O_345,N_9948,N_9940);
xnor UO_346 (O_346,N_9900,N_9978);
xor UO_347 (O_347,N_9945,N_9929);
nand UO_348 (O_348,N_9982,N_9971);
xnor UO_349 (O_349,N_9912,N_9924);
or UO_350 (O_350,N_9950,N_9974);
or UO_351 (O_351,N_9905,N_9921);
nand UO_352 (O_352,N_9980,N_9917);
xor UO_353 (O_353,N_9939,N_9978);
or UO_354 (O_354,N_9948,N_9970);
xnor UO_355 (O_355,N_9952,N_9929);
and UO_356 (O_356,N_9945,N_9975);
or UO_357 (O_357,N_9957,N_9921);
xnor UO_358 (O_358,N_9907,N_9912);
and UO_359 (O_359,N_9943,N_9958);
nand UO_360 (O_360,N_9933,N_9909);
or UO_361 (O_361,N_9972,N_9913);
or UO_362 (O_362,N_9922,N_9969);
nand UO_363 (O_363,N_9960,N_9995);
xor UO_364 (O_364,N_9990,N_9911);
or UO_365 (O_365,N_9983,N_9928);
nand UO_366 (O_366,N_9926,N_9944);
or UO_367 (O_367,N_9975,N_9971);
nor UO_368 (O_368,N_9906,N_9949);
or UO_369 (O_369,N_9964,N_9972);
or UO_370 (O_370,N_9936,N_9933);
nor UO_371 (O_371,N_9928,N_9975);
or UO_372 (O_372,N_9991,N_9989);
xnor UO_373 (O_373,N_9961,N_9968);
and UO_374 (O_374,N_9955,N_9940);
and UO_375 (O_375,N_9940,N_9922);
nand UO_376 (O_376,N_9924,N_9964);
or UO_377 (O_377,N_9914,N_9905);
and UO_378 (O_378,N_9973,N_9933);
or UO_379 (O_379,N_9975,N_9919);
xnor UO_380 (O_380,N_9914,N_9964);
or UO_381 (O_381,N_9920,N_9924);
or UO_382 (O_382,N_9914,N_9955);
and UO_383 (O_383,N_9980,N_9912);
or UO_384 (O_384,N_9969,N_9908);
xnor UO_385 (O_385,N_9906,N_9929);
xnor UO_386 (O_386,N_9930,N_9952);
xor UO_387 (O_387,N_9903,N_9904);
xnor UO_388 (O_388,N_9922,N_9905);
xor UO_389 (O_389,N_9945,N_9965);
nor UO_390 (O_390,N_9940,N_9905);
xnor UO_391 (O_391,N_9999,N_9981);
and UO_392 (O_392,N_9979,N_9908);
nor UO_393 (O_393,N_9976,N_9998);
nand UO_394 (O_394,N_9999,N_9923);
nand UO_395 (O_395,N_9976,N_9999);
and UO_396 (O_396,N_9917,N_9938);
nor UO_397 (O_397,N_9984,N_9962);
nand UO_398 (O_398,N_9910,N_9911);
and UO_399 (O_399,N_9964,N_9947);
xor UO_400 (O_400,N_9996,N_9905);
xor UO_401 (O_401,N_9989,N_9979);
nand UO_402 (O_402,N_9994,N_9928);
nand UO_403 (O_403,N_9996,N_9944);
nor UO_404 (O_404,N_9904,N_9997);
xor UO_405 (O_405,N_9996,N_9974);
and UO_406 (O_406,N_9919,N_9904);
nand UO_407 (O_407,N_9954,N_9963);
or UO_408 (O_408,N_9954,N_9902);
nand UO_409 (O_409,N_9912,N_9955);
xnor UO_410 (O_410,N_9990,N_9936);
nor UO_411 (O_411,N_9975,N_9902);
and UO_412 (O_412,N_9983,N_9932);
nor UO_413 (O_413,N_9915,N_9995);
and UO_414 (O_414,N_9903,N_9935);
xnor UO_415 (O_415,N_9962,N_9933);
nand UO_416 (O_416,N_9954,N_9965);
xnor UO_417 (O_417,N_9947,N_9941);
and UO_418 (O_418,N_9976,N_9912);
nor UO_419 (O_419,N_9963,N_9906);
xor UO_420 (O_420,N_9956,N_9954);
nand UO_421 (O_421,N_9918,N_9944);
nand UO_422 (O_422,N_9933,N_9964);
or UO_423 (O_423,N_9992,N_9949);
and UO_424 (O_424,N_9900,N_9972);
nand UO_425 (O_425,N_9909,N_9939);
xor UO_426 (O_426,N_9969,N_9953);
xnor UO_427 (O_427,N_9918,N_9913);
xnor UO_428 (O_428,N_9925,N_9913);
or UO_429 (O_429,N_9962,N_9915);
nand UO_430 (O_430,N_9980,N_9938);
or UO_431 (O_431,N_9969,N_9952);
and UO_432 (O_432,N_9924,N_9923);
or UO_433 (O_433,N_9961,N_9965);
nor UO_434 (O_434,N_9958,N_9961);
nand UO_435 (O_435,N_9956,N_9996);
xor UO_436 (O_436,N_9974,N_9970);
nor UO_437 (O_437,N_9907,N_9940);
and UO_438 (O_438,N_9975,N_9986);
nor UO_439 (O_439,N_9940,N_9978);
or UO_440 (O_440,N_9933,N_9969);
nand UO_441 (O_441,N_9906,N_9932);
xor UO_442 (O_442,N_9913,N_9962);
nand UO_443 (O_443,N_9937,N_9988);
or UO_444 (O_444,N_9996,N_9972);
nand UO_445 (O_445,N_9988,N_9945);
xor UO_446 (O_446,N_9948,N_9908);
and UO_447 (O_447,N_9981,N_9945);
and UO_448 (O_448,N_9958,N_9989);
nand UO_449 (O_449,N_9992,N_9987);
nand UO_450 (O_450,N_9939,N_9985);
xor UO_451 (O_451,N_9940,N_9959);
and UO_452 (O_452,N_9915,N_9960);
nand UO_453 (O_453,N_9929,N_9962);
and UO_454 (O_454,N_9906,N_9964);
and UO_455 (O_455,N_9946,N_9963);
nand UO_456 (O_456,N_9921,N_9956);
xnor UO_457 (O_457,N_9902,N_9905);
and UO_458 (O_458,N_9958,N_9924);
or UO_459 (O_459,N_9955,N_9970);
nand UO_460 (O_460,N_9915,N_9976);
nor UO_461 (O_461,N_9986,N_9931);
and UO_462 (O_462,N_9904,N_9999);
nor UO_463 (O_463,N_9927,N_9937);
and UO_464 (O_464,N_9922,N_9974);
or UO_465 (O_465,N_9982,N_9915);
or UO_466 (O_466,N_9933,N_9923);
nor UO_467 (O_467,N_9971,N_9995);
or UO_468 (O_468,N_9970,N_9913);
and UO_469 (O_469,N_9928,N_9948);
or UO_470 (O_470,N_9968,N_9953);
nand UO_471 (O_471,N_9907,N_9919);
xnor UO_472 (O_472,N_9906,N_9965);
nor UO_473 (O_473,N_9919,N_9957);
xor UO_474 (O_474,N_9925,N_9977);
nor UO_475 (O_475,N_9943,N_9962);
nand UO_476 (O_476,N_9914,N_9971);
and UO_477 (O_477,N_9976,N_9971);
or UO_478 (O_478,N_9949,N_9913);
nand UO_479 (O_479,N_9924,N_9995);
and UO_480 (O_480,N_9901,N_9931);
and UO_481 (O_481,N_9991,N_9943);
nand UO_482 (O_482,N_9949,N_9903);
nand UO_483 (O_483,N_9975,N_9952);
and UO_484 (O_484,N_9912,N_9944);
nand UO_485 (O_485,N_9970,N_9996);
nor UO_486 (O_486,N_9926,N_9925);
nand UO_487 (O_487,N_9908,N_9930);
nand UO_488 (O_488,N_9953,N_9934);
nand UO_489 (O_489,N_9958,N_9930);
xor UO_490 (O_490,N_9966,N_9946);
or UO_491 (O_491,N_9979,N_9994);
xnor UO_492 (O_492,N_9958,N_9931);
xnor UO_493 (O_493,N_9950,N_9904);
nor UO_494 (O_494,N_9927,N_9992);
nand UO_495 (O_495,N_9961,N_9907);
and UO_496 (O_496,N_9936,N_9934);
xnor UO_497 (O_497,N_9991,N_9931);
nor UO_498 (O_498,N_9907,N_9904);
or UO_499 (O_499,N_9970,N_9992);
nand UO_500 (O_500,N_9996,N_9982);
and UO_501 (O_501,N_9917,N_9975);
nor UO_502 (O_502,N_9912,N_9993);
xnor UO_503 (O_503,N_9913,N_9900);
or UO_504 (O_504,N_9955,N_9923);
and UO_505 (O_505,N_9969,N_9956);
and UO_506 (O_506,N_9967,N_9963);
and UO_507 (O_507,N_9994,N_9919);
or UO_508 (O_508,N_9959,N_9980);
and UO_509 (O_509,N_9943,N_9900);
or UO_510 (O_510,N_9987,N_9931);
xnor UO_511 (O_511,N_9948,N_9915);
nor UO_512 (O_512,N_9996,N_9964);
and UO_513 (O_513,N_9971,N_9993);
or UO_514 (O_514,N_9954,N_9995);
nor UO_515 (O_515,N_9967,N_9947);
nor UO_516 (O_516,N_9944,N_9979);
and UO_517 (O_517,N_9974,N_9917);
or UO_518 (O_518,N_9923,N_9972);
nor UO_519 (O_519,N_9939,N_9989);
nand UO_520 (O_520,N_9949,N_9961);
xor UO_521 (O_521,N_9978,N_9947);
and UO_522 (O_522,N_9942,N_9990);
nor UO_523 (O_523,N_9960,N_9947);
nor UO_524 (O_524,N_9950,N_9998);
nand UO_525 (O_525,N_9991,N_9964);
xnor UO_526 (O_526,N_9958,N_9935);
or UO_527 (O_527,N_9971,N_9900);
and UO_528 (O_528,N_9959,N_9971);
or UO_529 (O_529,N_9925,N_9909);
nand UO_530 (O_530,N_9956,N_9931);
and UO_531 (O_531,N_9947,N_9938);
nor UO_532 (O_532,N_9982,N_9925);
nor UO_533 (O_533,N_9918,N_9974);
nand UO_534 (O_534,N_9980,N_9943);
and UO_535 (O_535,N_9990,N_9932);
or UO_536 (O_536,N_9937,N_9958);
and UO_537 (O_537,N_9983,N_9981);
nand UO_538 (O_538,N_9982,N_9950);
xor UO_539 (O_539,N_9918,N_9948);
nand UO_540 (O_540,N_9917,N_9929);
nand UO_541 (O_541,N_9945,N_9900);
or UO_542 (O_542,N_9914,N_9916);
nor UO_543 (O_543,N_9916,N_9925);
xnor UO_544 (O_544,N_9955,N_9946);
nor UO_545 (O_545,N_9974,N_9956);
nor UO_546 (O_546,N_9968,N_9914);
and UO_547 (O_547,N_9913,N_9985);
nor UO_548 (O_548,N_9944,N_9961);
nor UO_549 (O_549,N_9921,N_9992);
nand UO_550 (O_550,N_9915,N_9920);
nand UO_551 (O_551,N_9981,N_9959);
nor UO_552 (O_552,N_9947,N_9931);
and UO_553 (O_553,N_9972,N_9942);
or UO_554 (O_554,N_9939,N_9936);
and UO_555 (O_555,N_9914,N_9996);
xnor UO_556 (O_556,N_9944,N_9960);
nor UO_557 (O_557,N_9911,N_9906);
xnor UO_558 (O_558,N_9944,N_9998);
xor UO_559 (O_559,N_9951,N_9985);
nor UO_560 (O_560,N_9973,N_9966);
xnor UO_561 (O_561,N_9988,N_9929);
nor UO_562 (O_562,N_9923,N_9945);
nor UO_563 (O_563,N_9919,N_9972);
xor UO_564 (O_564,N_9900,N_9915);
nor UO_565 (O_565,N_9912,N_9972);
or UO_566 (O_566,N_9981,N_9941);
and UO_567 (O_567,N_9913,N_9938);
and UO_568 (O_568,N_9900,N_9948);
and UO_569 (O_569,N_9908,N_9920);
nor UO_570 (O_570,N_9963,N_9950);
or UO_571 (O_571,N_9946,N_9989);
nor UO_572 (O_572,N_9927,N_9938);
xnor UO_573 (O_573,N_9960,N_9970);
and UO_574 (O_574,N_9984,N_9985);
and UO_575 (O_575,N_9946,N_9985);
nand UO_576 (O_576,N_9902,N_9995);
xor UO_577 (O_577,N_9931,N_9963);
xnor UO_578 (O_578,N_9969,N_9975);
xnor UO_579 (O_579,N_9986,N_9981);
nand UO_580 (O_580,N_9935,N_9957);
xor UO_581 (O_581,N_9993,N_9909);
nand UO_582 (O_582,N_9962,N_9964);
nand UO_583 (O_583,N_9921,N_9910);
nor UO_584 (O_584,N_9952,N_9960);
or UO_585 (O_585,N_9929,N_9934);
or UO_586 (O_586,N_9972,N_9995);
nand UO_587 (O_587,N_9908,N_9907);
or UO_588 (O_588,N_9927,N_9978);
nand UO_589 (O_589,N_9994,N_9952);
or UO_590 (O_590,N_9917,N_9919);
and UO_591 (O_591,N_9953,N_9947);
nor UO_592 (O_592,N_9941,N_9916);
xor UO_593 (O_593,N_9953,N_9903);
and UO_594 (O_594,N_9967,N_9987);
xor UO_595 (O_595,N_9932,N_9992);
nor UO_596 (O_596,N_9995,N_9956);
nor UO_597 (O_597,N_9955,N_9934);
or UO_598 (O_598,N_9998,N_9986);
nand UO_599 (O_599,N_9956,N_9958);
and UO_600 (O_600,N_9955,N_9964);
or UO_601 (O_601,N_9922,N_9943);
or UO_602 (O_602,N_9950,N_9934);
xnor UO_603 (O_603,N_9951,N_9907);
xor UO_604 (O_604,N_9958,N_9940);
xor UO_605 (O_605,N_9988,N_9958);
or UO_606 (O_606,N_9959,N_9942);
or UO_607 (O_607,N_9983,N_9956);
nor UO_608 (O_608,N_9936,N_9931);
and UO_609 (O_609,N_9910,N_9903);
nand UO_610 (O_610,N_9987,N_9902);
nand UO_611 (O_611,N_9942,N_9922);
xnor UO_612 (O_612,N_9920,N_9901);
and UO_613 (O_613,N_9968,N_9998);
or UO_614 (O_614,N_9970,N_9912);
or UO_615 (O_615,N_9918,N_9950);
nand UO_616 (O_616,N_9937,N_9976);
or UO_617 (O_617,N_9934,N_9988);
xor UO_618 (O_618,N_9952,N_9965);
xor UO_619 (O_619,N_9991,N_9979);
or UO_620 (O_620,N_9908,N_9985);
xnor UO_621 (O_621,N_9998,N_9988);
nand UO_622 (O_622,N_9930,N_9900);
xor UO_623 (O_623,N_9959,N_9925);
or UO_624 (O_624,N_9923,N_9990);
nor UO_625 (O_625,N_9908,N_9941);
and UO_626 (O_626,N_9989,N_9987);
or UO_627 (O_627,N_9923,N_9939);
and UO_628 (O_628,N_9954,N_9984);
xnor UO_629 (O_629,N_9959,N_9998);
xor UO_630 (O_630,N_9942,N_9970);
and UO_631 (O_631,N_9986,N_9965);
xor UO_632 (O_632,N_9989,N_9953);
and UO_633 (O_633,N_9936,N_9966);
xor UO_634 (O_634,N_9923,N_9950);
xor UO_635 (O_635,N_9925,N_9974);
nor UO_636 (O_636,N_9974,N_9957);
or UO_637 (O_637,N_9941,N_9962);
xor UO_638 (O_638,N_9921,N_9982);
xnor UO_639 (O_639,N_9937,N_9950);
nand UO_640 (O_640,N_9924,N_9938);
or UO_641 (O_641,N_9936,N_9941);
nor UO_642 (O_642,N_9936,N_9974);
and UO_643 (O_643,N_9962,N_9926);
nand UO_644 (O_644,N_9904,N_9913);
nand UO_645 (O_645,N_9910,N_9983);
or UO_646 (O_646,N_9950,N_9922);
nor UO_647 (O_647,N_9957,N_9980);
and UO_648 (O_648,N_9930,N_9935);
xor UO_649 (O_649,N_9982,N_9988);
and UO_650 (O_650,N_9906,N_9983);
nand UO_651 (O_651,N_9949,N_9976);
nor UO_652 (O_652,N_9965,N_9948);
nor UO_653 (O_653,N_9906,N_9993);
or UO_654 (O_654,N_9926,N_9952);
nand UO_655 (O_655,N_9973,N_9908);
nor UO_656 (O_656,N_9931,N_9974);
xor UO_657 (O_657,N_9905,N_9925);
or UO_658 (O_658,N_9904,N_9945);
xor UO_659 (O_659,N_9915,N_9931);
xnor UO_660 (O_660,N_9987,N_9962);
nor UO_661 (O_661,N_9912,N_9978);
xnor UO_662 (O_662,N_9906,N_9995);
and UO_663 (O_663,N_9958,N_9949);
nand UO_664 (O_664,N_9951,N_9929);
nand UO_665 (O_665,N_9917,N_9964);
or UO_666 (O_666,N_9920,N_9993);
and UO_667 (O_667,N_9917,N_9972);
nand UO_668 (O_668,N_9979,N_9960);
nor UO_669 (O_669,N_9974,N_9915);
and UO_670 (O_670,N_9941,N_9920);
or UO_671 (O_671,N_9947,N_9940);
and UO_672 (O_672,N_9958,N_9906);
nor UO_673 (O_673,N_9996,N_9938);
nor UO_674 (O_674,N_9957,N_9965);
xor UO_675 (O_675,N_9976,N_9944);
nand UO_676 (O_676,N_9958,N_9986);
nor UO_677 (O_677,N_9970,N_9968);
xor UO_678 (O_678,N_9992,N_9912);
nand UO_679 (O_679,N_9956,N_9909);
xnor UO_680 (O_680,N_9981,N_9902);
xor UO_681 (O_681,N_9992,N_9990);
xor UO_682 (O_682,N_9918,N_9986);
xnor UO_683 (O_683,N_9901,N_9957);
and UO_684 (O_684,N_9940,N_9903);
or UO_685 (O_685,N_9934,N_9948);
or UO_686 (O_686,N_9970,N_9936);
and UO_687 (O_687,N_9932,N_9988);
and UO_688 (O_688,N_9920,N_9921);
or UO_689 (O_689,N_9970,N_9925);
nor UO_690 (O_690,N_9938,N_9935);
nor UO_691 (O_691,N_9911,N_9971);
nand UO_692 (O_692,N_9978,N_9949);
nand UO_693 (O_693,N_9979,N_9952);
nor UO_694 (O_694,N_9918,N_9953);
and UO_695 (O_695,N_9930,N_9929);
nand UO_696 (O_696,N_9982,N_9955);
xnor UO_697 (O_697,N_9909,N_9958);
nand UO_698 (O_698,N_9998,N_9991);
nand UO_699 (O_699,N_9997,N_9970);
and UO_700 (O_700,N_9995,N_9967);
nor UO_701 (O_701,N_9967,N_9909);
and UO_702 (O_702,N_9955,N_9996);
nor UO_703 (O_703,N_9989,N_9951);
or UO_704 (O_704,N_9944,N_9983);
xor UO_705 (O_705,N_9936,N_9976);
xor UO_706 (O_706,N_9946,N_9992);
or UO_707 (O_707,N_9972,N_9971);
or UO_708 (O_708,N_9976,N_9933);
xor UO_709 (O_709,N_9986,N_9979);
xor UO_710 (O_710,N_9932,N_9944);
nand UO_711 (O_711,N_9940,N_9988);
nand UO_712 (O_712,N_9924,N_9918);
nand UO_713 (O_713,N_9970,N_9947);
nor UO_714 (O_714,N_9948,N_9945);
or UO_715 (O_715,N_9956,N_9952);
nor UO_716 (O_716,N_9953,N_9925);
xor UO_717 (O_717,N_9982,N_9956);
or UO_718 (O_718,N_9980,N_9945);
nor UO_719 (O_719,N_9979,N_9988);
nand UO_720 (O_720,N_9934,N_9979);
or UO_721 (O_721,N_9907,N_9971);
and UO_722 (O_722,N_9939,N_9924);
nor UO_723 (O_723,N_9956,N_9976);
and UO_724 (O_724,N_9934,N_9937);
and UO_725 (O_725,N_9931,N_9923);
xnor UO_726 (O_726,N_9983,N_9991);
or UO_727 (O_727,N_9989,N_9926);
or UO_728 (O_728,N_9949,N_9979);
nor UO_729 (O_729,N_9974,N_9955);
nor UO_730 (O_730,N_9973,N_9909);
nand UO_731 (O_731,N_9904,N_9915);
nor UO_732 (O_732,N_9912,N_9919);
xnor UO_733 (O_733,N_9999,N_9911);
or UO_734 (O_734,N_9927,N_9945);
nor UO_735 (O_735,N_9940,N_9931);
and UO_736 (O_736,N_9961,N_9948);
nor UO_737 (O_737,N_9982,N_9958);
and UO_738 (O_738,N_9947,N_9999);
nor UO_739 (O_739,N_9971,N_9901);
and UO_740 (O_740,N_9923,N_9966);
and UO_741 (O_741,N_9967,N_9927);
and UO_742 (O_742,N_9939,N_9967);
and UO_743 (O_743,N_9930,N_9951);
nand UO_744 (O_744,N_9917,N_9940);
xor UO_745 (O_745,N_9917,N_9930);
xnor UO_746 (O_746,N_9908,N_9982);
nand UO_747 (O_747,N_9934,N_9981);
and UO_748 (O_748,N_9952,N_9920);
or UO_749 (O_749,N_9940,N_9913);
nor UO_750 (O_750,N_9927,N_9924);
nor UO_751 (O_751,N_9916,N_9939);
or UO_752 (O_752,N_9922,N_9954);
nand UO_753 (O_753,N_9903,N_9922);
xnor UO_754 (O_754,N_9934,N_9931);
or UO_755 (O_755,N_9922,N_9909);
nand UO_756 (O_756,N_9918,N_9925);
and UO_757 (O_757,N_9956,N_9930);
nor UO_758 (O_758,N_9974,N_9951);
nand UO_759 (O_759,N_9966,N_9998);
nand UO_760 (O_760,N_9942,N_9943);
or UO_761 (O_761,N_9943,N_9949);
or UO_762 (O_762,N_9930,N_9934);
nand UO_763 (O_763,N_9941,N_9994);
nand UO_764 (O_764,N_9920,N_9988);
nor UO_765 (O_765,N_9984,N_9922);
xnor UO_766 (O_766,N_9984,N_9904);
or UO_767 (O_767,N_9996,N_9931);
or UO_768 (O_768,N_9939,N_9965);
or UO_769 (O_769,N_9955,N_9977);
nor UO_770 (O_770,N_9934,N_9972);
nor UO_771 (O_771,N_9993,N_9949);
and UO_772 (O_772,N_9922,N_9996);
nand UO_773 (O_773,N_9902,N_9939);
and UO_774 (O_774,N_9928,N_9980);
nand UO_775 (O_775,N_9901,N_9926);
nand UO_776 (O_776,N_9904,N_9998);
xnor UO_777 (O_777,N_9933,N_9920);
or UO_778 (O_778,N_9946,N_9917);
nor UO_779 (O_779,N_9983,N_9975);
or UO_780 (O_780,N_9998,N_9989);
xnor UO_781 (O_781,N_9926,N_9966);
and UO_782 (O_782,N_9901,N_9916);
and UO_783 (O_783,N_9948,N_9956);
nor UO_784 (O_784,N_9905,N_9992);
and UO_785 (O_785,N_9938,N_9995);
and UO_786 (O_786,N_9933,N_9944);
or UO_787 (O_787,N_9909,N_9937);
nor UO_788 (O_788,N_9997,N_9977);
or UO_789 (O_789,N_9999,N_9903);
or UO_790 (O_790,N_9920,N_9946);
or UO_791 (O_791,N_9982,N_9940);
xnor UO_792 (O_792,N_9917,N_9992);
xor UO_793 (O_793,N_9903,N_9966);
nor UO_794 (O_794,N_9912,N_9938);
xor UO_795 (O_795,N_9970,N_9959);
nand UO_796 (O_796,N_9972,N_9983);
and UO_797 (O_797,N_9911,N_9998);
and UO_798 (O_798,N_9906,N_9975);
and UO_799 (O_799,N_9962,N_9989);
and UO_800 (O_800,N_9982,N_9997);
or UO_801 (O_801,N_9944,N_9965);
or UO_802 (O_802,N_9927,N_9932);
nor UO_803 (O_803,N_9911,N_9929);
xnor UO_804 (O_804,N_9919,N_9932);
xnor UO_805 (O_805,N_9934,N_9985);
nor UO_806 (O_806,N_9994,N_9902);
nor UO_807 (O_807,N_9957,N_9983);
xor UO_808 (O_808,N_9907,N_9939);
nor UO_809 (O_809,N_9956,N_9981);
nand UO_810 (O_810,N_9959,N_9920);
or UO_811 (O_811,N_9975,N_9958);
and UO_812 (O_812,N_9903,N_9951);
xor UO_813 (O_813,N_9935,N_9912);
nand UO_814 (O_814,N_9960,N_9906);
nor UO_815 (O_815,N_9916,N_9966);
and UO_816 (O_816,N_9934,N_9964);
or UO_817 (O_817,N_9940,N_9993);
and UO_818 (O_818,N_9900,N_9925);
or UO_819 (O_819,N_9994,N_9969);
nor UO_820 (O_820,N_9908,N_9928);
nand UO_821 (O_821,N_9971,N_9931);
nor UO_822 (O_822,N_9985,N_9976);
and UO_823 (O_823,N_9998,N_9970);
or UO_824 (O_824,N_9974,N_9937);
nor UO_825 (O_825,N_9939,N_9918);
nand UO_826 (O_826,N_9976,N_9911);
nand UO_827 (O_827,N_9971,N_9992);
or UO_828 (O_828,N_9958,N_9962);
nor UO_829 (O_829,N_9904,N_9928);
or UO_830 (O_830,N_9932,N_9961);
or UO_831 (O_831,N_9956,N_9903);
nor UO_832 (O_832,N_9937,N_9995);
xor UO_833 (O_833,N_9926,N_9964);
or UO_834 (O_834,N_9935,N_9944);
and UO_835 (O_835,N_9999,N_9997);
xor UO_836 (O_836,N_9976,N_9992);
and UO_837 (O_837,N_9986,N_9991);
and UO_838 (O_838,N_9994,N_9906);
or UO_839 (O_839,N_9953,N_9913);
xor UO_840 (O_840,N_9992,N_9965);
nor UO_841 (O_841,N_9908,N_9909);
and UO_842 (O_842,N_9924,N_9903);
and UO_843 (O_843,N_9971,N_9954);
or UO_844 (O_844,N_9920,N_9936);
nand UO_845 (O_845,N_9983,N_9969);
nand UO_846 (O_846,N_9970,N_9915);
or UO_847 (O_847,N_9928,N_9932);
nor UO_848 (O_848,N_9929,N_9982);
nand UO_849 (O_849,N_9962,N_9950);
nand UO_850 (O_850,N_9995,N_9936);
and UO_851 (O_851,N_9910,N_9991);
nand UO_852 (O_852,N_9946,N_9921);
nand UO_853 (O_853,N_9958,N_9985);
nand UO_854 (O_854,N_9937,N_9948);
or UO_855 (O_855,N_9908,N_9972);
and UO_856 (O_856,N_9967,N_9900);
nand UO_857 (O_857,N_9904,N_9935);
and UO_858 (O_858,N_9917,N_9981);
xor UO_859 (O_859,N_9985,N_9904);
and UO_860 (O_860,N_9977,N_9980);
nor UO_861 (O_861,N_9990,N_9971);
or UO_862 (O_862,N_9926,N_9909);
nand UO_863 (O_863,N_9917,N_9983);
xor UO_864 (O_864,N_9948,N_9971);
nand UO_865 (O_865,N_9975,N_9956);
or UO_866 (O_866,N_9954,N_9997);
xor UO_867 (O_867,N_9942,N_9955);
nand UO_868 (O_868,N_9985,N_9912);
nor UO_869 (O_869,N_9906,N_9901);
nand UO_870 (O_870,N_9999,N_9994);
or UO_871 (O_871,N_9907,N_9960);
nor UO_872 (O_872,N_9996,N_9941);
or UO_873 (O_873,N_9984,N_9941);
nor UO_874 (O_874,N_9901,N_9983);
and UO_875 (O_875,N_9912,N_9974);
or UO_876 (O_876,N_9951,N_9978);
xnor UO_877 (O_877,N_9923,N_9997);
nand UO_878 (O_878,N_9963,N_9902);
or UO_879 (O_879,N_9961,N_9928);
xnor UO_880 (O_880,N_9967,N_9917);
or UO_881 (O_881,N_9926,N_9902);
nand UO_882 (O_882,N_9921,N_9907);
xor UO_883 (O_883,N_9993,N_9967);
or UO_884 (O_884,N_9907,N_9964);
xor UO_885 (O_885,N_9931,N_9985);
xor UO_886 (O_886,N_9966,N_9905);
nor UO_887 (O_887,N_9993,N_9944);
and UO_888 (O_888,N_9998,N_9907);
and UO_889 (O_889,N_9988,N_9972);
nor UO_890 (O_890,N_9955,N_9952);
and UO_891 (O_891,N_9978,N_9921);
xor UO_892 (O_892,N_9929,N_9972);
nand UO_893 (O_893,N_9907,N_9909);
nand UO_894 (O_894,N_9977,N_9910);
nor UO_895 (O_895,N_9900,N_9926);
and UO_896 (O_896,N_9910,N_9900);
xnor UO_897 (O_897,N_9909,N_9938);
nand UO_898 (O_898,N_9986,N_9937);
xor UO_899 (O_899,N_9959,N_9931);
xor UO_900 (O_900,N_9939,N_9930);
or UO_901 (O_901,N_9912,N_9977);
nor UO_902 (O_902,N_9973,N_9953);
or UO_903 (O_903,N_9924,N_9929);
or UO_904 (O_904,N_9921,N_9950);
or UO_905 (O_905,N_9926,N_9914);
xor UO_906 (O_906,N_9904,N_9976);
and UO_907 (O_907,N_9950,N_9925);
nand UO_908 (O_908,N_9916,N_9945);
nand UO_909 (O_909,N_9980,N_9915);
xor UO_910 (O_910,N_9924,N_9951);
and UO_911 (O_911,N_9986,N_9927);
and UO_912 (O_912,N_9995,N_9973);
nand UO_913 (O_913,N_9951,N_9911);
nand UO_914 (O_914,N_9996,N_9990);
nor UO_915 (O_915,N_9951,N_9988);
and UO_916 (O_916,N_9951,N_9984);
nand UO_917 (O_917,N_9901,N_9918);
nor UO_918 (O_918,N_9919,N_9924);
xnor UO_919 (O_919,N_9923,N_9959);
xnor UO_920 (O_920,N_9958,N_9954);
nor UO_921 (O_921,N_9949,N_9990);
nand UO_922 (O_922,N_9931,N_9967);
nor UO_923 (O_923,N_9921,N_9995);
and UO_924 (O_924,N_9992,N_9991);
nor UO_925 (O_925,N_9913,N_9923);
xnor UO_926 (O_926,N_9910,N_9961);
nor UO_927 (O_927,N_9925,N_9997);
or UO_928 (O_928,N_9906,N_9936);
nor UO_929 (O_929,N_9916,N_9978);
nand UO_930 (O_930,N_9953,N_9993);
xnor UO_931 (O_931,N_9927,N_9950);
nor UO_932 (O_932,N_9932,N_9942);
nor UO_933 (O_933,N_9915,N_9966);
or UO_934 (O_934,N_9918,N_9946);
nand UO_935 (O_935,N_9968,N_9929);
and UO_936 (O_936,N_9975,N_9962);
xor UO_937 (O_937,N_9929,N_9977);
nor UO_938 (O_938,N_9937,N_9906);
or UO_939 (O_939,N_9962,N_9939);
nand UO_940 (O_940,N_9972,N_9902);
nand UO_941 (O_941,N_9939,N_9961);
or UO_942 (O_942,N_9986,N_9916);
nand UO_943 (O_943,N_9984,N_9995);
nand UO_944 (O_944,N_9982,N_9974);
nor UO_945 (O_945,N_9995,N_9931);
xnor UO_946 (O_946,N_9970,N_9944);
and UO_947 (O_947,N_9983,N_9939);
and UO_948 (O_948,N_9944,N_9943);
or UO_949 (O_949,N_9933,N_9958);
nor UO_950 (O_950,N_9946,N_9916);
nor UO_951 (O_951,N_9920,N_9971);
nand UO_952 (O_952,N_9944,N_9990);
or UO_953 (O_953,N_9978,N_9907);
nand UO_954 (O_954,N_9937,N_9990);
nand UO_955 (O_955,N_9994,N_9918);
nand UO_956 (O_956,N_9976,N_9957);
or UO_957 (O_957,N_9974,N_9929);
nor UO_958 (O_958,N_9951,N_9921);
and UO_959 (O_959,N_9990,N_9977);
and UO_960 (O_960,N_9912,N_9934);
xnor UO_961 (O_961,N_9981,N_9935);
and UO_962 (O_962,N_9921,N_9994);
and UO_963 (O_963,N_9955,N_9981);
or UO_964 (O_964,N_9920,N_9973);
nor UO_965 (O_965,N_9921,N_9999);
and UO_966 (O_966,N_9930,N_9975);
and UO_967 (O_967,N_9981,N_9908);
nor UO_968 (O_968,N_9900,N_9963);
nor UO_969 (O_969,N_9995,N_9978);
and UO_970 (O_970,N_9931,N_9999);
and UO_971 (O_971,N_9949,N_9940);
or UO_972 (O_972,N_9948,N_9926);
nand UO_973 (O_973,N_9977,N_9968);
and UO_974 (O_974,N_9966,N_9982);
nor UO_975 (O_975,N_9934,N_9994);
or UO_976 (O_976,N_9984,N_9977);
nor UO_977 (O_977,N_9937,N_9981);
and UO_978 (O_978,N_9946,N_9980);
or UO_979 (O_979,N_9999,N_9927);
nand UO_980 (O_980,N_9982,N_9918);
nand UO_981 (O_981,N_9933,N_9945);
nor UO_982 (O_982,N_9921,N_9986);
nand UO_983 (O_983,N_9913,N_9941);
nor UO_984 (O_984,N_9927,N_9977);
nand UO_985 (O_985,N_9969,N_9957);
nor UO_986 (O_986,N_9950,N_9961);
xnor UO_987 (O_987,N_9919,N_9926);
nor UO_988 (O_988,N_9965,N_9947);
nor UO_989 (O_989,N_9912,N_9952);
nand UO_990 (O_990,N_9924,N_9936);
or UO_991 (O_991,N_9939,N_9970);
and UO_992 (O_992,N_9937,N_9984);
nand UO_993 (O_993,N_9936,N_9959);
xor UO_994 (O_994,N_9920,N_9909);
xnor UO_995 (O_995,N_9990,N_9959);
nor UO_996 (O_996,N_9945,N_9939);
xor UO_997 (O_997,N_9944,N_9995);
and UO_998 (O_998,N_9983,N_9930);
nand UO_999 (O_999,N_9983,N_9993);
nand UO_1000 (O_1000,N_9949,N_9994);
nor UO_1001 (O_1001,N_9928,N_9926);
or UO_1002 (O_1002,N_9996,N_9933);
and UO_1003 (O_1003,N_9997,N_9946);
xor UO_1004 (O_1004,N_9999,N_9916);
xor UO_1005 (O_1005,N_9920,N_9954);
and UO_1006 (O_1006,N_9908,N_9918);
and UO_1007 (O_1007,N_9939,N_9952);
and UO_1008 (O_1008,N_9919,N_9955);
and UO_1009 (O_1009,N_9944,N_9919);
and UO_1010 (O_1010,N_9976,N_9940);
nand UO_1011 (O_1011,N_9970,N_9935);
and UO_1012 (O_1012,N_9987,N_9956);
nand UO_1013 (O_1013,N_9945,N_9962);
xnor UO_1014 (O_1014,N_9931,N_9981);
nor UO_1015 (O_1015,N_9938,N_9974);
nand UO_1016 (O_1016,N_9900,N_9999);
xor UO_1017 (O_1017,N_9994,N_9920);
or UO_1018 (O_1018,N_9967,N_9911);
nor UO_1019 (O_1019,N_9909,N_9977);
or UO_1020 (O_1020,N_9902,N_9916);
nor UO_1021 (O_1021,N_9935,N_9934);
nand UO_1022 (O_1022,N_9937,N_9913);
or UO_1023 (O_1023,N_9988,N_9903);
nand UO_1024 (O_1024,N_9940,N_9906);
nand UO_1025 (O_1025,N_9981,N_9979);
or UO_1026 (O_1026,N_9914,N_9985);
and UO_1027 (O_1027,N_9937,N_9928);
and UO_1028 (O_1028,N_9962,N_9949);
nand UO_1029 (O_1029,N_9948,N_9996);
nand UO_1030 (O_1030,N_9923,N_9915);
nand UO_1031 (O_1031,N_9985,N_9927);
xor UO_1032 (O_1032,N_9935,N_9969);
or UO_1033 (O_1033,N_9918,N_9916);
and UO_1034 (O_1034,N_9994,N_9931);
nand UO_1035 (O_1035,N_9962,N_9954);
nor UO_1036 (O_1036,N_9988,N_9962);
or UO_1037 (O_1037,N_9965,N_9923);
or UO_1038 (O_1038,N_9941,N_9976);
or UO_1039 (O_1039,N_9901,N_9952);
or UO_1040 (O_1040,N_9960,N_9983);
and UO_1041 (O_1041,N_9916,N_9932);
or UO_1042 (O_1042,N_9967,N_9912);
nor UO_1043 (O_1043,N_9973,N_9938);
and UO_1044 (O_1044,N_9938,N_9962);
xnor UO_1045 (O_1045,N_9947,N_9910);
nor UO_1046 (O_1046,N_9931,N_9912);
xor UO_1047 (O_1047,N_9962,N_9971);
or UO_1048 (O_1048,N_9971,N_9981);
and UO_1049 (O_1049,N_9964,N_9984);
nand UO_1050 (O_1050,N_9946,N_9948);
and UO_1051 (O_1051,N_9980,N_9994);
nor UO_1052 (O_1052,N_9970,N_9923);
xor UO_1053 (O_1053,N_9973,N_9981);
nor UO_1054 (O_1054,N_9971,N_9984);
and UO_1055 (O_1055,N_9912,N_9908);
xor UO_1056 (O_1056,N_9966,N_9912);
or UO_1057 (O_1057,N_9989,N_9914);
nand UO_1058 (O_1058,N_9959,N_9977);
nand UO_1059 (O_1059,N_9902,N_9969);
xnor UO_1060 (O_1060,N_9972,N_9959);
nor UO_1061 (O_1061,N_9932,N_9922);
xor UO_1062 (O_1062,N_9938,N_9931);
or UO_1063 (O_1063,N_9959,N_9979);
or UO_1064 (O_1064,N_9951,N_9948);
and UO_1065 (O_1065,N_9939,N_9946);
and UO_1066 (O_1066,N_9914,N_9948);
xor UO_1067 (O_1067,N_9925,N_9948);
or UO_1068 (O_1068,N_9979,N_9977);
nand UO_1069 (O_1069,N_9985,N_9997);
or UO_1070 (O_1070,N_9938,N_9906);
nor UO_1071 (O_1071,N_9980,N_9954);
or UO_1072 (O_1072,N_9997,N_9973);
or UO_1073 (O_1073,N_9904,N_9917);
or UO_1074 (O_1074,N_9974,N_9900);
xnor UO_1075 (O_1075,N_9921,N_9925);
and UO_1076 (O_1076,N_9973,N_9991);
nand UO_1077 (O_1077,N_9972,N_9954);
or UO_1078 (O_1078,N_9956,N_9993);
and UO_1079 (O_1079,N_9992,N_9951);
nand UO_1080 (O_1080,N_9919,N_9959);
or UO_1081 (O_1081,N_9903,N_9925);
nor UO_1082 (O_1082,N_9972,N_9977);
or UO_1083 (O_1083,N_9994,N_9991);
or UO_1084 (O_1084,N_9976,N_9993);
nand UO_1085 (O_1085,N_9992,N_9937);
or UO_1086 (O_1086,N_9924,N_9970);
and UO_1087 (O_1087,N_9914,N_9972);
or UO_1088 (O_1088,N_9995,N_9977);
and UO_1089 (O_1089,N_9914,N_9936);
nor UO_1090 (O_1090,N_9991,N_9939);
or UO_1091 (O_1091,N_9988,N_9950);
nand UO_1092 (O_1092,N_9973,N_9901);
and UO_1093 (O_1093,N_9999,N_9978);
and UO_1094 (O_1094,N_9944,N_9901);
and UO_1095 (O_1095,N_9998,N_9922);
or UO_1096 (O_1096,N_9910,N_9959);
nand UO_1097 (O_1097,N_9903,N_9905);
nand UO_1098 (O_1098,N_9969,N_9919);
xnor UO_1099 (O_1099,N_9954,N_9900);
nor UO_1100 (O_1100,N_9965,N_9918);
and UO_1101 (O_1101,N_9993,N_9945);
nor UO_1102 (O_1102,N_9939,N_9990);
nand UO_1103 (O_1103,N_9974,N_9944);
and UO_1104 (O_1104,N_9990,N_9933);
xnor UO_1105 (O_1105,N_9908,N_9950);
and UO_1106 (O_1106,N_9973,N_9957);
or UO_1107 (O_1107,N_9908,N_9970);
nor UO_1108 (O_1108,N_9991,N_9952);
and UO_1109 (O_1109,N_9952,N_9946);
xnor UO_1110 (O_1110,N_9960,N_9946);
nor UO_1111 (O_1111,N_9981,N_9965);
nor UO_1112 (O_1112,N_9984,N_9998);
nand UO_1113 (O_1113,N_9922,N_9912);
xnor UO_1114 (O_1114,N_9965,N_9950);
xnor UO_1115 (O_1115,N_9948,N_9936);
or UO_1116 (O_1116,N_9995,N_9990);
or UO_1117 (O_1117,N_9944,N_9988);
and UO_1118 (O_1118,N_9940,N_9960);
nor UO_1119 (O_1119,N_9920,N_9996);
nand UO_1120 (O_1120,N_9927,N_9979);
nand UO_1121 (O_1121,N_9924,N_9922);
xor UO_1122 (O_1122,N_9915,N_9901);
nand UO_1123 (O_1123,N_9987,N_9938);
nand UO_1124 (O_1124,N_9983,N_9999);
nand UO_1125 (O_1125,N_9964,N_9910);
or UO_1126 (O_1126,N_9949,N_9911);
xnor UO_1127 (O_1127,N_9982,N_9953);
nand UO_1128 (O_1128,N_9945,N_9957);
and UO_1129 (O_1129,N_9990,N_9905);
xnor UO_1130 (O_1130,N_9944,N_9997);
and UO_1131 (O_1131,N_9940,N_9936);
xnor UO_1132 (O_1132,N_9957,N_9928);
xor UO_1133 (O_1133,N_9961,N_9901);
or UO_1134 (O_1134,N_9989,N_9947);
and UO_1135 (O_1135,N_9950,N_9980);
xnor UO_1136 (O_1136,N_9932,N_9998);
or UO_1137 (O_1137,N_9908,N_9943);
or UO_1138 (O_1138,N_9919,N_9941);
nor UO_1139 (O_1139,N_9910,N_9962);
nand UO_1140 (O_1140,N_9948,N_9909);
or UO_1141 (O_1141,N_9993,N_9914);
and UO_1142 (O_1142,N_9911,N_9975);
and UO_1143 (O_1143,N_9977,N_9965);
xnor UO_1144 (O_1144,N_9943,N_9932);
nor UO_1145 (O_1145,N_9936,N_9957);
nand UO_1146 (O_1146,N_9923,N_9926);
nand UO_1147 (O_1147,N_9933,N_9924);
and UO_1148 (O_1148,N_9955,N_9937);
xor UO_1149 (O_1149,N_9946,N_9970);
nand UO_1150 (O_1150,N_9989,N_9961);
and UO_1151 (O_1151,N_9978,N_9982);
or UO_1152 (O_1152,N_9956,N_9917);
or UO_1153 (O_1153,N_9931,N_9929);
nand UO_1154 (O_1154,N_9908,N_9952);
or UO_1155 (O_1155,N_9983,N_9937);
and UO_1156 (O_1156,N_9997,N_9901);
nand UO_1157 (O_1157,N_9987,N_9900);
nor UO_1158 (O_1158,N_9915,N_9924);
nor UO_1159 (O_1159,N_9914,N_9958);
and UO_1160 (O_1160,N_9999,N_9902);
or UO_1161 (O_1161,N_9937,N_9996);
xnor UO_1162 (O_1162,N_9968,N_9955);
nand UO_1163 (O_1163,N_9948,N_9992);
xor UO_1164 (O_1164,N_9971,N_9904);
nor UO_1165 (O_1165,N_9969,N_9959);
and UO_1166 (O_1166,N_9957,N_9926);
nor UO_1167 (O_1167,N_9938,N_9960);
nand UO_1168 (O_1168,N_9924,N_9952);
nand UO_1169 (O_1169,N_9928,N_9934);
nand UO_1170 (O_1170,N_9966,N_9941);
nor UO_1171 (O_1171,N_9983,N_9961);
and UO_1172 (O_1172,N_9997,N_9961);
or UO_1173 (O_1173,N_9922,N_9933);
or UO_1174 (O_1174,N_9980,N_9905);
nor UO_1175 (O_1175,N_9942,N_9946);
nand UO_1176 (O_1176,N_9928,N_9915);
nand UO_1177 (O_1177,N_9926,N_9920);
and UO_1178 (O_1178,N_9969,N_9947);
nand UO_1179 (O_1179,N_9984,N_9987);
or UO_1180 (O_1180,N_9930,N_9978);
or UO_1181 (O_1181,N_9928,N_9966);
or UO_1182 (O_1182,N_9907,N_9936);
xor UO_1183 (O_1183,N_9942,N_9935);
and UO_1184 (O_1184,N_9949,N_9964);
nor UO_1185 (O_1185,N_9939,N_9966);
or UO_1186 (O_1186,N_9949,N_9925);
nand UO_1187 (O_1187,N_9912,N_9946);
nand UO_1188 (O_1188,N_9974,N_9980);
nor UO_1189 (O_1189,N_9948,N_9973);
nor UO_1190 (O_1190,N_9927,N_9958);
or UO_1191 (O_1191,N_9984,N_9903);
or UO_1192 (O_1192,N_9920,N_9927);
or UO_1193 (O_1193,N_9932,N_9902);
or UO_1194 (O_1194,N_9921,N_9906);
nor UO_1195 (O_1195,N_9951,N_9912);
nor UO_1196 (O_1196,N_9971,N_9935);
and UO_1197 (O_1197,N_9960,N_9957);
xor UO_1198 (O_1198,N_9918,N_9945);
or UO_1199 (O_1199,N_9910,N_9960);
or UO_1200 (O_1200,N_9976,N_9989);
nor UO_1201 (O_1201,N_9994,N_9989);
and UO_1202 (O_1202,N_9916,N_9962);
and UO_1203 (O_1203,N_9976,N_9967);
nand UO_1204 (O_1204,N_9974,N_9989);
nor UO_1205 (O_1205,N_9909,N_9981);
and UO_1206 (O_1206,N_9977,N_9964);
or UO_1207 (O_1207,N_9992,N_9935);
or UO_1208 (O_1208,N_9939,N_9979);
xnor UO_1209 (O_1209,N_9988,N_9924);
and UO_1210 (O_1210,N_9928,N_9968);
nand UO_1211 (O_1211,N_9944,N_9968);
and UO_1212 (O_1212,N_9942,N_9979);
xnor UO_1213 (O_1213,N_9939,N_9943);
nor UO_1214 (O_1214,N_9950,N_9995);
xnor UO_1215 (O_1215,N_9936,N_9975);
and UO_1216 (O_1216,N_9905,N_9920);
or UO_1217 (O_1217,N_9922,N_9906);
nor UO_1218 (O_1218,N_9937,N_9949);
and UO_1219 (O_1219,N_9943,N_9938);
xnor UO_1220 (O_1220,N_9970,N_9989);
or UO_1221 (O_1221,N_9965,N_9938);
nor UO_1222 (O_1222,N_9955,N_9909);
nor UO_1223 (O_1223,N_9916,N_9905);
xor UO_1224 (O_1224,N_9911,N_9925);
nand UO_1225 (O_1225,N_9965,N_9915);
xnor UO_1226 (O_1226,N_9918,N_9951);
nand UO_1227 (O_1227,N_9908,N_9905);
xnor UO_1228 (O_1228,N_9993,N_9930);
nand UO_1229 (O_1229,N_9966,N_9981);
nor UO_1230 (O_1230,N_9959,N_9902);
xnor UO_1231 (O_1231,N_9997,N_9903);
xor UO_1232 (O_1232,N_9989,N_9933);
nor UO_1233 (O_1233,N_9966,N_9970);
nand UO_1234 (O_1234,N_9951,N_9952);
xor UO_1235 (O_1235,N_9914,N_9909);
nand UO_1236 (O_1236,N_9933,N_9911);
nor UO_1237 (O_1237,N_9903,N_9945);
nor UO_1238 (O_1238,N_9953,N_9990);
or UO_1239 (O_1239,N_9950,N_9949);
nand UO_1240 (O_1240,N_9972,N_9963);
nand UO_1241 (O_1241,N_9911,N_9955);
nor UO_1242 (O_1242,N_9973,N_9932);
and UO_1243 (O_1243,N_9913,N_9926);
xor UO_1244 (O_1244,N_9986,N_9932);
or UO_1245 (O_1245,N_9958,N_9942);
and UO_1246 (O_1246,N_9942,N_9952);
nand UO_1247 (O_1247,N_9911,N_9926);
nand UO_1248 (O_1248,N_9944,N_9992);
or UO_1249 (O_1249,N_9945,N_9989);
or UO_1250 (O_1250,N_9948,N_9984);
or UO_1251 (O_1251,N_9974,N_9995);
and UO_1252 (O_1252,N_9971,N_9937);
nor UO_1253 (O_1253,N_9991,N_9934);
xor UO_1254 (O_1254,N_9954,N_9993);
and UO_1255 (O_1255,N_9977,N_9940);
xnor UO_1256 (O_1256,N_9936,N_9971);
and UO_1257 (O_1257,N_9918,N_9947);
nor UO_1258 (O_1258,N_9910,N_9956);
xnor UO_1259 (O_1259,N_9915,N_9954);
nor UO_1260 (O_1260,N_9924,N_9973);
xor UO_1261 (O_1261,N_9969,N_9984);
nor UO_1262 (O_1262,N_9943,N_9955);
nor UO_1263 (O_1263,N_9966,N_9958);
nor UO_1264 (O_1264,N_9966,N_9944);
and UO_1265 (O_1265,N_9974,N_9945);
nand UO_1266 (O_1266,N_9979,N_9996);
and UO_1267 (O_1267,N_9917,N_9997);
and UO_1268 (O_1268,N_9914,N_9919);
nand UO_1269 (O_1269,N_9979,N_9953);
or UO_1270 (O_1270,N_9979,N_9973);
xnor UO_1271 (O_1271,N_9908,N_9924);
and UO_1272 (O_1272,N_9979,N_9917);
or UO_1273 (O_1273,N_9983,N_9942);
nor UO_1274 (O_1274,N_9977,N_9998);
nor UO_1275 (O_1275,N_9912,N_9975);
nor UO_1276 (O_1276,N_9947,N_9937);
or UO_1277 (O_1277,N_9964,N_9974);
nand UO_1278 (O_1278,N_9963,N_9984);
xnor UO_1279 (O_1279,N_9926,N_9924);
and UO_1280 (O_1280,N_9941,N_9987);
nand UO_1281 (O_1281,N_9972,N_9962);
xnor UO_1282 (O_1282,N_9928,N_9991);
xor UO_1283 (O_1283,N_9957,N_9953);
and UO_1284 (O_1284,N_9948,N_9949);
and UO_1285 (O_1285,N_9928,N_9970);
xor UO_1286 (O_1286,N_9968,N_9971);
xnor UO_1287 (O_1287,N_9928,N_9978);
xnor UO_1288 (O_1288,N_9967,N_9984);
nor UO_1289 (O_1289,N_9913,N_9952);
xor UO_1290 (O_1290,N_9946,N_9993);
nor UO_1291 (O_1291,N_9968,N_9950);
nand UO_1292 (O_1292,N_9920,N_9975);
or UO_1293 (O_1293,N_9903,N_9926);
nand UO_1294 (O_1294,N_9952,N_9998);
xor UO_1295 (O_1295,N_9931,N_9993);
nand UO_1296 (O_1296,N_9911,N_9942);
nand UO_1297 (O_1297,N_9916,N_9960);
or UO_1298 (O_1298,N_9989,N_9907);
or UO_1299 (O_1299,N_9953,N_9978);
nand UO_1300 (O_1300,N_9911,N_9919);
nand UO_1301 (O_1301,N_9987,N_9946);
xnor UO_1302 (O_1302,N_9911,N_9935);
or UO_1303 (O_1303,N_9996,N_9962);
nand UO_1304 (O_1304,N_9976,N_9963);
or UO_1305 (O_1305,N_9968,N_9913);
nand UO_1306 (O_1306,N_9988,N_9933);
and UO_1307 (O_1307,N_9937,N_9926);
nor UO_1308 (O_1308,N_9964,N_9930);
nor UO_1309 (O_1309,N_9988,N_9905);
or UO_1310 (O_1310,N_9926,N_9976);
xor UO_1311 (O_1311,N_9927,N_9903);
or UO_1312 (O_1312,N_9920,N_9951);
nor UO_1313 (O_1313,N_9918,N_9968);
nand UO_1314 (O_1314,N_9916,N_9998);
or UO_1315 (O_1315,N_9960,N_9978);
and UO_1316 (O_1316,N_9983,N_9953);
and UO_1317 (O_1317,N_9975,N_9908);
nand UO_1318 (O_1318,N_9943,N_9971);
nand UO_1319 (O_1319,N_9953,N_9910);
and UO_1320 (O_1320,N_9904,N_9981);
or UO_1321 (O_1321,N_9975,N_9977);
and UO_1322 (O_1322,N_9999,N_9912);
xnor UO_1323 (O_1323,N_9953,N_9977);
or UO_1324 (O_1324,N_9948,N_9998);
nor UO_1325 (O_1325,N_9947,N_9909);
or UO_1326 (O_1326,N_9912,N_9953);
xor UO_1327 (O_1327,N_9900,N_9922);
and UO_1328 (O_1328,N_9934,N_9989);
nand UO_1329 (O_1329,N_9954,N_9998);
nor UO_1330 (O_1330,N_9984,N_9989);
nand UO_1331 (O_1331,N_9964,N_9918);
and UO_1332 (O_1332,N_9950,N_9969);
nand UO_1333 (O_1333,N_9901,N_9995);
nor UO_1334 (O_1334,N_9968,N_9938);
xnor UO_1335 (O_1335,N_9912,N_9994);
xor UO_1336 (O_1336,N_9959,N_9967);
nand UO_1337 (O_1337,N_9935,N_9943);
xnor UO_1338 (O_1338,N_9924,N_9963);
nor UO_1339 (O_1339,N_9944,N_9928);
nand UO_1340 (O_1340,N_9934,N_9911);
or UO_1341 (O_1341,N_9921,N_9942);
nor UO_1342 (O_1342,N_9932,N_9968);
xnor UO_1343 (O_1343,N_9940,N_9985);
xnor UO_1344 (O_1344,N_9932,N_9965);
or UO_1345 (O_1345,N_9991,N_9916);
or UO_1346 (O_1346,N_9926,N_9992);
nand UO_1347 (O_1347,N_9959,N_9916);
xnor UO_1348 (O_1348,N_9901,N_9911);
xor UO_1349 (O_1349,N_9997,N_9986);
xnor UO_1350 (O_1350,N_9967,N_9906);
and UO_1351 (O_1351,N_9941,N_9980);
xor UO_1352 (O_1352,N_9940,N_9999);
or UO_1353 (O_1353,N_9936,N_9962);
and UO_1354 (O_1354,N_9914,N_9921);
nor UO_1355 (O_1355,N_9960,N_9964);
and UO_1356 (O_1356,N_9935,N_9917);
or UO_1357 (O_1357,N_9992,N_9906);
nand UO_1358 (O_1358,N_9937,N_9920);
and UO_1359 (O_1359,N_9967,N_9999);
nor UO_1360 (O_1360,N_9951,N_9996);
xor UO_1361 (O_1361,N_9993,N_9984);
xnor UO_1362 (O_1362,N_9904,N_9923);
nand UO_1363 (O_1363,N_9913,N_9995);
or UO_1364 (O_1364,N_9962,N_9935);
nand UO_1365 (O_1365,N_9991,N_9915);
nor UO_1366 (O_1366,N_9977,N_9902);
and UO_1367 (O_1367,N_9923,N_9967);
or UO_1368 (O_1368,N_9945,N_9983);
and UO_1369 (O_1369,N_9935,N_9902);
nand UO_1370 (O_1370,N_9999,N_9910);
or UO_1371 (O_1371,N_9995,N_9959);
xor UO_1372 (O_1372,N_9984,N_9927);
xor UO_1373 (O_1373,N_9928,N_9947);
nor UO_1374 (O_1374,N_9919,N_9993);
nor UO_1375 (O_1375,N_9961,N_9962);
nand UO_1376 (O_1376,N_9943,N_9920);
nand UO_1377 (O_1377,N_9917,N_9949);
nor UO_1378 (O_1378,N_9999,N_9922);
nor UO_1379 (O_1379,N_9986,N_9902);
and UO_1380 (O_1380,N_9992,N_9901);
nor UO_1381 (O_1381,N_9987,N_9999);
and UO_1382 (O_1382,N_9918,N_9993);
nor UO_1383 (O_1383,N_9940,N_9935);
or UO_1384 (O_1384,N_9989,N_9943);
and UO_1385 (O_1385,N_9913,N_9957);
xor UO_1386 (O_1386,N_9968,N_9949);
or UO_1387 (O_1387,N_9923,N_9960);
nor UO_1388 (O_1388,N_9936,N_9945);
and UO_1389 (O_1389,N_9920,N_9939);
or UO_1390 (O_1390,N_9998,N_9908);
xnor UO_1391 (O_1391,N_9997,N_9913);
and UO_1392 (O_1392,N_9968,N_9920);
nor UO_1393 (O_1393,N_9960,N_9932);
or UO_1394 (O_1394,N_9967,N_9977);
or UO_1395 (O_1395,N_9958,N_9993);
nor UO_1396 (O_1396,N_9958,N_9945);
and UO_1397 (O_1397,N_9989,N_9932);
nand UO_1398 (O_1398,N_9975,N_9968);
nand UO_1399 (O_1399,N_9942,N_9938);
nand UO_1400 (O_1400,N_9999,N_9975);
xnor UO_1401 (O_1401,N_9954,N_9950);
xor UO_1402 (O_1402,N_9946,N_9928);
or UO_1403 (O_1403,N_9901,N_9917);
nor UO_1404 (O_1404,N_9977,N_9935);
nand UO_1405 (O_1405,N_9903,N_9954);
nor UO_1406 (O_1406,N_9973,N_9950);
xnor UO_1407 (O_1407,N_9900,N_9993);
nand UO_1408 (O_1408,N_9965,N_9997);
nor UO_1409 (O_1409,N_9907,N_9970);
or UO_1410 (O_1410,N_9947,N_9944);
nand UO_1411 (O_1411,N_9953,N_9919);
and UO_1412 (O_1412,N_9959,N_9963);
and UO_1413 (O_1413,N_9920,N_9958);
nor UO_1414 (O_1414,N_9932,N_9962);
and UO_1415 (O_1415,N_9914,N_9979);
xor UO_1416 (O_1416,N_9970,N_9961);
nor UO_1417 (O_1417,N_9963,N_9917);
and UO_1418 (O_1418,N_9936,N_9900);
nor UO_1419 (O_1419,N_9952,N_9981);
and UO_1420 (O_1420,N_9920,N_9955);
nand UO_1421 (O_1421,N_9986,N_9983);
or UO_1422 (O_1422,N_9918,N_9989);
or UO_1423 (O_1423,N_9967,N_9986);
nand UO_1424 (O_1424,N_9961,N_9916);
and UO_1425 (O_1425,N_9978,N_9963);
nor UO_1426 (O_1426,N_9949,N_9999);
xnor UO_1427 (O_1427,N_9918,N_9975);
xnor UO_1428 (O_1428,N_9991,N_9967);
nand UO_1429 (O_1429,N_9979,N_9916);
and UO_1430 (O_1430,N_9941,N_9993);
or UO_1431 (O_1431,N_9930,N_9960);
or UO_1432 (O_1432,N_9944,N_9937);
xor UO_1433 (O_1433,N_9989,N_9995);
xnor UO_1434 (O_1434,N_9955,N_9950);
xnor UO_1435 (O_1435,N_9983,N_9946);
xnor UO_1436 (O_1436,N_9974,N_9933);
or UO_1437 (O_1437,N_9977,N_9976);
nor UO_1438 (O_1438,N_9907,N_9913);
nand UO_1439 (O_1439,N_9965,N_9967);
nor UO_1440 (O_1440,N_9918,N_9921);
or UO_1441 (O_1441,N_9947,N_9935);
nand UO_1442 (O_1442,N_9924,N_9989);
xnor UO_1443 (O_1443,N_9924,N_9917);
and UO_1444 (O_1444,N_9993,N_9989);
and UO_1445 (O_1445,N_9937,N_9904);
xor UO_1446 (O_1446,N_9929,N_9938);
nor UO_1447 (O_1447,N_9916,N_9951);
or UO_1448 (O_1448,N_9937,N_9959);
nand UO_1449 (O_1449,N_9972,N_9990);
or UO_1450 (O_1450,N_9984,N_9905);
xor UO_1451 (O_1451,N_9966,N_9904);
or UO_1452 (O_1452,N_9939,N_9975);
xnor UO_1453 (O_1453,N_9918,N_9917);
or UO_1454 (O_1454,N_9919,N_9910);
nand UO_1455 (O_1455,N_9954,N_9961);
and UO_1456 (O_1456,N_9901,N_9950);
xnor UO_1457 (O_1457,N_9980,N_9948);
xnor UO_1458 (O_1458,N_9966,N_9985);
and UO_1459 (O_1459,N_9961,N_9959);
nor UO_1460 (O_1460,N_9907,N_9952);
xor UO_1461 (O_1461,N_9900,N_9935);
nor UO_1462 (O_1462,N_9936,N_9917);
or UO_1463 (O_1463,N_9956,N_9937);
nand UO_1464 (O_1464,N_9955,N_9938);
xor UO_1465 (O_1465,N_9970,N_9977);
nand UO_1466 (O_1466,N_9920,N_9999);
nor UO_1467 (O_1467,N_9943,N_9941);
or UO_1468 (O_1468,N_9907,N_9945);
nand UO_1469 (O_1469,N_9928,N_9979);
nor UO_1470 (O_1470,N_9942,N_9927);
xor UO_1471 (O_1471,N_9960,N_9904);
or UO_1472 (O_1472,N_9919,N_9902);
and UO_1473 (O_1473,N_9944,N_9900);
or UO_1474 (O_1474,N_9959,N_9983);
and UO_1475 (O_1475,N_9968,N_9962);
nand UO_1476 (O_1476,N_9978,N_9984);
nand UO_1477 (O_1477,N_9982,N_9968);
or UO_1478 (O_1478,N_9977,N_9945);
nor UO_1479 (O_1479,N_9961,N_9925);
or UO_1480 (O_1480,N_9979,N_9965);
or UO_1481 (O_1481,N_9957,N_9947);
nand UO_1482 (O_1482,N_9969,N_9910);
or UO_1483 (O_1483,N_9993,N_9901);
or UO_1484 (O_1484,N_9953,N_9951);
or UO_1485 (O_1485,N_9901,N_9986);
or UO_1486 (O_1486,N_9980,N_9916);
nand UO_1487 (O_1487,N_9978,N_9987);
nor UO_1488 (O_1488,N_9992,N_9978);
nor UO_1489 (O_1489,N_9918,N_9962);
nor UO_1490 (O_1490,N_9917,N_9912);
nor UO_1491 (O_1491,N_9902,N_9984);
or UO_1492 (O_1492,N_9909,N_9916);
or UO_1493 (O_1493,N_9907,N_9991);
nand UO_1494 (O_1494,N_9980,N_9978);
or UO_1495 (O_1495,N_9977,N_9950);
nand UO_1496 (O_1496,N_9984,N_9945);
nand UO_1497 (O_1497,N_9972,N_9951);
xor UO_1498 (O_1498,N_9927,N_9969);
and UO_1499 (O_1499,N_9913,N_9964);
endmodule