module basic_500_3000_500_40_levels_2xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
or U0 (N_0,In_467,In_236);
or U1 (N_1,In_93,In_374);
nand U2 (N_2,In_382,In_5);
nor U3 (N_3,In_183,In_181);
nand U4 (N_4,In_334,In_395);
nor U5 (N_5,In_323,In_404);
nor U6 (N_6,In_25,In_65);
or U7 (N_7,In_310,In_384);
nand U8 (N_8,In_268,In_473);
or U9 (N_9,In_238,In_254);
nor U10 (N_10,In_78,In_159);
nand U11 (N_11,In_222,In_237);
nand U12 (N_12,In_193,In_249);
or U13 (N_13,In_21,In_312);
nand U14 (N_14,In_357,In_250);
and U15 (N_15,In_35,In_278);
and U16 (N_16,In_8,In_100);
xnor U17 (N_17,In_485,In_273);
nand U18 (N_18,In_387,In_296);
nand U19 (N_19,In_179,In_147);
or U20 (N_20,In_62,In_319);
nor U21 (N_21,In_487,In_212);
nand U22 (N_22,In_205,In_256);
and U23 (N_23,In_74,In_88);
xor U24 (N_24,In_418,In_82);
nor U25 (N_25,In_325,In_469);
nor U26 (N_26,In_414,In_182);
or U27 (N_27,In_162,In_191);
nor U28 (N_28,In_57,In_172);
and U29 (N_29,In_341,In_290);
nor U30 (N_30,In_379,In_40);
and U31 (N_31,In_129,In_184);
nor U32 (N_32,In_208,In_386);
and U33 (N_33,In_192,In_491);
and U34 (N_34,In_330,In_335);
nor U35 (N_35,In_381,In_200);
nor U36 (N_36,In_114,In_13);
nor U37 (N_37,In_291,In_429);
nand U38 (N_38,In_391,In_36);
nand U39 (N_39,In_318,In_456);
and U40 (N_40,In_136,In_143);
and U41 (N_41,In_402,In_116);
or U42 (N_42,In_400,In_112);
nand U43 (N_43,In_284,In_393);
or U44 (N_44,In_17,In_71);
or U45 (N_45,In_288,In_23);
nor U46 (N_46,In_104,In_92);
and U47 (N_47,In_347,In_107);
nand U48 (N_48,In_331,In_377);
and U49 (N_49,In_432,In_232);
nor U50 (N_50,In_175,In_102);
and U51 (N_51,In_252,In_297);
or U52 (N_52,In_287,In_239);
nand U53 (N_53,In_26,In_144);
or U54 (N_54,In_195,In_321);
or U55 (N_55,In_446,In_1);
or U56 (N_56,In_210,In_439);
xnor U57 (N_57,In_369,In_316);
or U58 (N_58,In_242,In_241);
nand U59 (N_59,In_224,In_443);
or U60 (N_60,In_96,In_203);
nand U61 (N_61,In_348,In_405);
nand U62 (N_62,In_226,In_324);
nor U63 (N_63,In_190,In_176);
and U64 (N_64,In_263,In_59);
nor U65 (N_65,In_265,In_362);
nand U66 (N_66,In_320,In_251);
nor U67 (N_67,In_279,In_86);
and U68 (N_68,In_180,In_213);
or U69 (N_69,In_34,In_15);
and U70 (N_70,In_11,In_73);
and U71 (N_71,In_217,In_253);
or U72 (N_72,In_255,In_465);
or U73 (N_73,In_267,In_480);
nand U74 (N_74,In_458,In_177);
and U75 (N_75,In_422,In_257);
nor U76 (N_76,In_295,In_264);
or U77 (N_77,In_18,In_122);
and U78 (N_78,In_132,In_77);
nand U79 (N_79,In_332,In_160);
xnor U80 (N_80,N_15,In_152);
or U81 (N_81,In_135,N_0);
nor U82 (N_82,In_29,In_139);
nor U83 (N_83,In_276,In_428);
nor U84 (N_84,In_338,In_219);
nor U85 (N_85,In_388,In_294);
or U86 (N_86,In_486,In_120);
nor U87 (N_87,In_399,In_365);
nand U88 (N_88,In_140,N_21);
or U89 (N_89,In_427,In_466);
or U90 (N_90,In_42,N_27);
or U91 (N_91,In_186,In_234);
nand U92 (N_92,In_451,In_385);
and U93 (N_93,In_63,In_138);
nand U94 (N_94,N_22,In_484);
or U95 (N_95,In_281,In_389);
or U96 (N_96,N_26,In_328);
nand U97 (N_97,In_302,In_336);
or U98 (N_98,N_74,In_2);
nor U99 (N_99,In_390,In_482);
nand U100 (N_100,In_157,In_499);
or U101 (N_101,In_342,In_375);
nand U102 (N_102,N_19,In_353);
nand U103 (N_103,In_364,N_42);
nand U104 (N_104,In_12,In_449);
xor U105 (N_105,N_8,In_309);
and U106 (N_106,In_0,In_174);
nand U107 (N_107,In_475,In_53);
nand U108 (N_108,In_105,N_51);
and U109 (N_109,In_277,N_59);
or U110 (N_110,In_194,In_289);
and U111 (N_111,In_206,N_17);
nand U112 (N_112,In_271,In_45);
xnor U113 (N_113,In_413,In_245);
and U114 (N_114,In_10,In_344);
nand U115 (N_115,N_31,In_398);
or U116 (N_116,In_60,In_424);
nand U117 (N_117,In_43,In_37);
and U118 (N_118,In_83,In_202);
nor U119 (N_119,In_119,In_161);
and U120 (N_120,In_343,In_275);
nor U121 (N_121,In_261,In_141);
or U122 (N_122,N_45,In_260);
or U123 (N_123,In_483,In_233);
nand U124 (N_124,In_168,In_81);
or U125 (N_125,In_305,In_470);
and U126 (N_126,In_113,In_149);
nor U127 (N_127,N_30,In_87);
nor U128 (N_128,In_372,N_46);
nand U129 (N_129,In_489,In_22);
and U130 (N_130,In_409,In_445);
nand U131 (N_131,In_125,N_67);
and U132 (N_132,In_340,N_25);
nor U133 (N_133,In_196,In_95);
nor U134 (N_134,In_490,In_401);
or U135 (N_135,In_356,N_3);
nor U136 (N_136,In_410,In_201);
nand U137 (N_137,In_154,In_51);
nand U138 (N_138,In_229,In_438);
nand U139 (N_139,N_38,In_69);
nor U140 (N_140,N_23,In_454);
nand U141 (N_141,In_231,In_142);
nor U142 (N_142,In_207,In_376);
nor U143 (N_143,In_58,In_150);
and U144 (N_144,In_464,N_63);
nand U145 (N_145,In_94,In_370);
nor U146 (N_146,In_270,N_58);
or U147 (N_147,In_70,In_198);
and U148 (N_148,N_72,In_283);
or U149 (N_149,In_492,In_27);
nand U150 (N_150,In_121,N_83);
nor U151 (N_151,N_97,N_141);
or U152 (N_152,N_81,N_35);
or U153 (N_153,N_85,In_303);
or U154 (N_154,In_165,N_57);
and U155 (N_155,In_478,In_280);
nor U156 (N_156,In_156,In_378);
nand U157 (N_157,N_13,In_227);
or U158 (N_158,N_28,N_99);
and U159 (N_159,In_108,In_89);
nor U160 (N_160,N_79,In_355);
or U161 (N_161,In_115,In_298);
or U162 (N_162,In_339,In_97);
nor U163 (N_163,In_423,In_462);
or U164 (N_164,N_91,N_89);
and U165 (N_165,In_9,In_488);
nor U166 (N_166,N_41,In_118);
nor U167 (N_167,In_98,N_7);
and U168 (N_168,In_272,In_461);
and U169 (N_169,In_3,N_44);
or U170 (N_170,In_425,In_313);
xor U171 (N_171,In_479,N_146);
or U172 (N_172,In_75,In_247);
nor U173 (N_173,N_129,In_373);
or U174 (N_174,N_43,In_197);
nand U175 (N_175,In_444,In_285);
nor U176 (N_176,In_493,In_359);
nand U177 (N_177,In_472,In_56);
nand U178 (N_178,N_87,In_223);
nand U179 (N_179,In_350,In_54);
nor U180 (N_180,N_86,N_70);
nand U181 (N_181,N_62,In_292);
nand U182 (N_182,N_110,In_333);
or U183 (N_183,N_16,N_73);
nor U184 (N_184,N_12,In_240);
nand U185 (N_185,In_228,In_366);
and U186 (N_186,N_112,N_128);
nor U187 (N_187,N_78,In_433);
nor U188 (N_188,In_266,In_419);
or U189 (N_189,N_11,In_170);
and U190 (N_190,In_55,In_435);
nand U191 (N_191,In_392,In_477);
nand U192 (N_192,N_36,N_80);
or U193 (N_193,In_322,In_109);
or U194 (N_194,N_94,N_20);
and U195 (N_195,In_440,In_178);
nand U196 (N_196,In_243,In_166);
nor U197 (N_197,In_131,In_468);
and U198 (N_198,In_308,In_117);
and U199 (N_199,N_56,N_5);
and U200 (N_200,In_24,In_337);
or U201 (N_201,In_354,In_358);
nand U202 (N_202,In_158,In_430);
and U203 (N_203,N_148,In_155);
and U204 (N_204,N_68,In_188);
nor U205 (N_205,N_149,In_85);
and U206 (N_206,In_99,N_145);
nand U207 (N_207,In_7,N_64);
nor U208 (N_208,N_133,In_361);
and U209 (N_209,In_420,N_144);
and U210 (N_210,N_106,In_412);
and U211 (N_211,In_304,N_134);
nand U212 (N_212,In_90,In_367);
and U213 (N_213,In_14,In_19);
nor U214 (N_214,In_459,In_408);
nand U215 (N_215,In_153,In_244);
and U216 (N_216,In_471,N_71);
or U217 (N_217,In_259,N_98);
and U218 (N_218,In_199,In_146);
or U219 (N_219,In_49,N_32);
and U220 (N_220,In_103,N_130);
or U221 (N_221,In_415,N_37);
nand U222 (N_222,N_120,N_10);
nor U223 (N_223,In_476,N_108);
nor U224 (N_224,In_106,In_216);
or U225 (N_225,N_224,In_126);
nand U226 (N_226,N_102,In_167);
or U227 (N_227,N_118,In_52);
nor U228 (N_228,N_131,N_139);
nand U229 (N_229,In_326,In_383);
nor U230 (N_230,N_171,In_80);
nand U231 (N_231,In_286,In_417);
xor U232 (N_232,N_138,In_453);
or U233 (N_233,In_163,N_150);
and U234 (N_234,N_180,In_28);
nor U235 (N_235,In_16,In_442);
and U236 (N_236,In_235,In_41);
nand U237 (N_237,N_135,In_148);
nor U238 (N_238,N_153,N_193);
and U239 (N_239,In_185,In_474);
or U240 (N_240,N_209,In_30);
or U241 (N_241,N_105,In_460);
or U242 (N_242,N_104,N_175);
nor U243 (N_243,N_196,In_301);
nand U244 (N_244,N_117,N_220);
nand U245 (N_245,N_214,N_140);
nor U246 (N_246,In_434,In_351);
xnor U247 (N_247,N_113,N_121);
or U248 (N_248,N_198,In_211);
or U249 (N_249,In_421,N_93);
and U250 (N_250,N_127,In_431);
nor U251 (N_251,In_368,In_416);
or U252 (N_252,N_189,In_91);
nand U253 (N_253,In_300,In_327);
xor U254 (N_254,In_457,In_110);
nor U255 (N_255,In_495,In_215);
and U256 (N_256,In_494,N_49);
or U257 (N_257,In_352,N_188);
nor U258 (N_258,N_191,In_38);
nor U259 (N_259,N_200,N_219);
or U260 (N_260,N_197,In_220);
and U261 (N_261,N_164,In_246);
xnor U262 (N_262,N_65,In_317);
and U263 (N_263,In_189,In_307);
or U264 (N_264,N_33,In_371);
or U265 (N_265,In_455,N_9);
nand U266 (N_266,In_130,N_223);
nand U267 (N_267,In_463,In_345);
or U268 (N_268,N_159,In_214);
nand U269 (N_269,N_173,N_143);
and U270 (N_270,N_152,N_77);
and U271 (N_271,N_207,N_82);
or U272 (N_272,In_221,In_218);
nor U273 (N_273,In_496,N_2);
nand U274 (N_274,In_269,N_199);
nor U275 (N_275,N_96,N_14);
nor U276 (N_276,In_329,N_109);
nor U277 (N_277,N_204,In_396);
nand U278 (N_278,N_185,In_299);
nor U279 (N_279,In_84,In_123);
nor U280 (N_280,N_176,N_151);
nor U281 (N_281,N_48,N_160);
nor U282 (N_282,In_481,N_54);
nand U283 (N_283,N_177,In_447);
nand U284 (N_284,N_95,In_436);
nand U285 (N_285,N_4,N_221);
nor U286 (N_286,In_258,In_64);
and U287 (N_287,In_111,N_170);
and U288 (N_288,In_248,In_33);
and U289 (N_289,In_293,In_44);
and U290 (N_290,In_209,In_50);
or U291 (N_291,In_46,N_217);
nor U292 (N_292,In_282,N_213);
or U293 (N_293,N_116,N_222);
nor U294 (N_294,N_34,In_128);
or U295 (N_295,In_315,In_31);
nand U296 (N_296,N_47,In_145);
xor U297 (N_297,N_29,N_202);
or U298 (N_298,N_39,In_68);
and U299 (N_299,In_204,N_162);
nor U300 (N_300,N_259,N_256);
nor U301 (N_301,N_181,In_48);
or U302 (N_302,N_61,N_161);
nand U303 (N_303,In_133,In_406);
and U304 (N_304,N_84,N_294);
xnor U305 (N_305,N_289,In_47);
nand U306 (N_306,N_107,N_211);
nor U307 (N_307,In_169,In_151);
and U308 (N_308,N_276,In_230);
and U309 (N_309,N_292,In_6);
nand U310 (N_310,N_119,N_92);
nand U311 (N_311,N_258,N_53);
or U312 (N_312,N_242,In_173);
nand U313 (N_313,In_441,N_69);
nor U314 (N_314,N_285,In_450);
nand U315 (N_315,N_228,N_243);
nand U316 (N_316,N_293,In_314);
nand U317 (N_317,N_186,In_20);
or U318 (N_318,N_55,N_206);
nand U319 (N_319,N_190,N_247);
or U320 (N_320,N_167,N_257);
nor U321 (N_321,N_178,N_218);
nor U322 (N_322,N_157,In_4);
nand U323 (N_323,N_136,N_52);
nor U324 (N_324,N_234,In_262);
and U325 (N_325,N_279,N_194);
nor U326 (N_326,N_122,N_142);
and U327 (N_327,In_363,N_66);
nor U328 (N_328,N_248,N_272);
nand U329 (N_329,N_290,N_169);
or U330 (N_330,N_271,N_179);
nor U331 (N_331,N_165,N_268);
or U332 (N_332,N_205,N_158);
or U333 (N_333,N_264,N_168);
and U334 (N_334,In_403,N_246);
or U335 (N_335,N_261,N_210);
or U336 (N_336,N_182,N_286);
and U337 (N_337,In_349,N_269);
or U338 (N_338,In_311,In_124);
nand U339 (N_339,N_282,N_299);
nand U340 (N_340,In_394,N_238);
or U341 (N_341,N_277,N_230);
and U342 (N_342,In_137,N_75);
nor U343 (N_343,N_296,In_225);
nor U344 (N_344,N_291,N_1);
or U345 (N_345,N_250,N_172);
nand U346 (N_346,In_346,In_134);
nor U347 (N_347,N_280,N_288);
nand U348 (N_348,N_244,N_226);
or U349 (N_349,In_76,N_260);
xor U350 (N_350,N_274,N_227);
nor U351 (N_351,N_156,N_50);
and U352 (N_352,N_187,N_225);
and U353 (N_353,N_267,N_283);
and U354 (N_354,N_295,N_184);
or U355 (N_355,N_298,N_137);
and U356 (N_356,N_270,N_125);
or U357 (N_357,N_101,N_253);
xor U358 (N_358,In_452,N_40);
nor U359 (N_359,N_100,N_233);
or U360 (N_360,N_215,N_132);
nand U361 (N_361,In_411,N_266);
or U362 (N_362,In_360,N_241);
nor U363 (N_363,In_79,N_249);
and U364 (N_364,N_60,N_251);
nor U365 (N_365,N_278,In_407);
xor U366 (N_366,N_76,N_208);
and U367 (N_367,N_166,In_171);
and U368 (N_368,In_164,N_195);
nor U369 (N_369,N_262,N_6);
nor U370 (N_370,N_154,N_201);
or U371 (N_371,N_273,N_240);
and U372 (N_372,In_72,N_231);
or U373 (N_373,In_497,N_255);
nand U374 (N_374,N_275,N_281);
nand U375 (N_375,N_301,N_346);
nand U376 (N_376,N_340,N_315);
xnor U377 (N_377,N_174,N_350);
nand U378 (N_378,N_124,N_103);
or U379 (N_379,In_67,N_317);
nand U380 (N_380,N_367,N_326);
nand U381 (N_381,N_343,In_274);
and U382 (N_382,N_329,N_322);
or U383 (N_383,N_368,In_187);
and U384 (N_384,N_313,N_338);
and U385 (N_385,N_366,N_358);
nor U386 (N_386,N_351,N_353);
nand U387 (N_387,N_359,N_354);
and U388 (N_388,In_39,N_341);
or U389 (N_389,N_370,N_327);
nand U390 (N_390,N_318,N_111);
nand U391 (N_391,N_328,N_374);
or U392 (N_392,N_335,N_362);
and U393 (N_393,N_316,N_365);
or U394 (N_394,N_321,N_320);
nand U395 (N_395,N_245,N_373);
nand U396 (N_396,N_307,N_342);
nand U397 (N_397,In_380,N_356);
or U398 (N_398,N_237,N_309);
nand U399 (N_399,N_308,In_127);
nand U400 (N_400,N_265,N_254);
nand U401 (N_401,N_126,N_163);
and U402 (N_402,N_352,N_155);
or U403 (N_403,In_426,N_305);
and U404 (N_404,N_361,N_311);
nor U405 (N_405,N_347,In_437);
nand U406 (N_406,N_344,In_397);
or U407 (N_407,N_239,N_300);
and U408 (N_408,N_235,N_302);
or U409 (N_409,In_448,N_360);
or U410 (N_410,N_331,N_330);
nand U411 (N_411,N_24,In_306);
or U412 (N_412,N_371,N_349);
and U413 (N_413,In_498,N_252);
or U414 (N_414,N_345,In_101);
or U415 (N_415,N_90,N_306);
nor U416 (N_416,N_333,N_363);
and U417 (N_417,N_115,In_32);
and U418 (N_418,N_263,N_303);
or U419 (N_419,N_18,N_236);
nand U420 (N_420,N_216,In_66);
nand U421 (N_421,N_88,N_339);
and U422 (N_422,N_323,N_314);
xnor U423 (N_423,N_203,N_183);
nand U424 (N_424,N_332,N_364);
nand U425 (N_425,N_297,N_355);
or U426 (N_426,N_312,In_61);
and U427 (N_427,N_324,N_147);
nor U428 (N_428,N_357,N_232);
xor U429 (N_429,N_284,N_325);
nor U430 (N_430,N_114,N_369);
nor U431 (N_431,N_287,N_337);
nand U432 (N_432,N_123,N_334);
or U433 (N_433,N_229,N_304);
nor U434 (N_434,N_348,N_336);
nor U435 (N_435,N_310,N_372);
or U436 (N_436,N_192,N_319);
or U437 (N_437,N_212,N_331);
nor U438 (N_438,N_360,In_67);
nor U439 (N_439,N_370,N_123);
or U440 (N_440,N_335,In_274);
and U441 (N_441,N_312,N_88);
and U442 (N_442,N_370,In_66);
and U443 (N_443,N_372,N_350);
nand U444 (N_444,N_103,N_183);
nand U445 (N_445,N_192,N_124);
nand U446 (N_446,N_124,N_343);
and U447 (N_447,N_326,In_127);
nor U448 (N_448,N_252,N_315);
or U449 (N_449,N_245,N_297);
xnor U450 (N_450,N_378,N_387);
nor U451 (N_451,N_393,N_444);
and U452 (N_452,N_375,N_416);
and U453 (N_453,N_431,N_397);
nor U454 (N_454,N_408,N_384);
nor U455 (N_455,N_422,N_398);
or U456 (N_456,N_390,N_406);
nor U457 (N_457,N_412,N_441);
nor U458 (N_458,N_429,N_445);
nand U459 (N_459,N_386,N_426);
or U460 (N_460,N_415,N_427);
nor U461 (N_461,N_379,N_381);
nor U462 (N_462,N_382,N_418);
or U463 (N_463,N_443,N_423);
and U464 (N_464,N_405,N_401);
nor U465 (N_465,N_402,N_428);
and U466 (N_466,N_414,N_432);
or U467 (N_467,N_439,N_442);
and U468 (N_468,N_395,N_419);
nor U469 (N_469,N_403,N_446);
or U470 (N_470,N_383,N_411);
nor U471 (N_471,N_449,N_388);
nand U472 (N_472,N_421,N_440);
nor U473 (N_473,N_420,N_389);
and U474 (N_474,N_436,N_396);
or U475 (N_475,N_385,N_433);
nor U476 (N_476,N_376,N_448);
and U477 (N_477,N_434,N_380);
or U478 (N_478,N_430,N_447);
nor U479 (N_479,N_391,N_400);
and U480 (N_480,N_407,N_392);
nor U481 (N_481,N_438,N_435);
or U482 (N_482,N_410,N_413);
or U483 (N_483,N_377,N_394);
nand U484 (N_484,N_425,N_424);
or U485 (N_485,N_404,N_437);
and U486 (N_486,N_399,N_409);
and U487 (N_487,N_417,N_387);
nor U488 (N_488,N_447,N_420);
nor U489 (N_489,N_408,N_386);
xor U490 (N_490,N_436,N_432);
nand U491 (N_491,N_392,N_378);
and U492 (N_492,N_392,N_376);
nor U493 (N_493,N_390,N_410);
nor U494 (N_494,N_441,N_445);
nor U495 (N_495,N_435,N_397);
and U496 (N_496,N_398,N_423);
nand U497 (N_497,N_379,N_424);
nand U498 (N_498,N_382,N_443);
and U499 (N_499,N_418,N_444);
and U500 (N_500,N_433,N_413);
nand U501 (N_501,N_415,N_407);
nor U502 (N_502,N_420,N_426);
nand U503 (N_503,N_425,N_441);
and U504 (N_504,N_449,N_424);
or U505 (N_505,N_392,N_403);
nor U506 (N_506,N_438,N_394);
or U507 (N_507,N_381,N_420);
nor U508 (N_508,N_397,N_395);
and U509 (N_509,N_423,N_396);
and U510 (N_510,N_413,N_376);
or U511 (N_511,N_448,N_444);
nor U512 (N_512,N_442,N_403);
or U513 (N_513,N_416,N_422);
nand U514 (N_514,N_392,N_443);
and U515 (N_515,N_409,N_382);
or U516 (N_516,N_414,N_388);
and U517 (N_517,N_392,N_437);
and U518 (N_518,N_427,N_437);
and U519 (N_519,N_423,N_385);
or U520 (N_520,N_429,N_447);
nor U521 (N_521,N_388,N_443);
nor U522 (N_522,N_389,N_414);
and U523 (N_523,N_419,N_423);
or U524 (N_524,N_388,N_444);
and U525 (N_525,N_524,N_485);
nand U526 (N_526,N_493,N_517);
nor U527 (N_527,N_464,N_501);
and U528 (N_528,N_461,N_456);
or U529 (N_529,N_515,N_518);
and U530 (N_530,N_505,N_516);
nand U531 (N_531,N_497,N_522);
nand U532 (N_532,N_473,N_460);
and U533 (N_533,N_487,N_452);
or U534 (N_534,N_451,N_506);
and U535 (N_535,N_511,N_512);
and U536 (N_536,N_508,N_488);
and U537 (N_537,N_465,N_519);
nand U538 (N_538,N_457,N_498);
or U539 (N_539,N_521,N_478);
nand U540 (N_540,N_474,N_507);
nand U541 (N_541,N_490,N_467);
nand U542 (N_542,N_484,N_475);
and U543 (N_543,N_491,N_489);
nor U544 (N_544,N_500,N_492);
or U545 (N_545,N_504,N_455);
and U546 (N_546,N_496,N_494);
nor U547 (N_547,N_458,N_514);
xor U548 (N_548,N_450,N_499);
nand U549 (N_549,N_513,N_481);
or U550 (N_550,N_495,N_471);
or U551 (N_551,N_502,N_453);
nand U552 (N_552,N_459,N_468);
nor U553 (N_553,N_470,N_523);
and U554 (N_554,N_466,N_469);
nand U555 (N_555,N_509,N_472);
nor U556 (N_556,N_482,N_510);
xor U557 (N_557,N_486,N_463);
and U558 (N_558,N_480,N_503);
nand U559 (N_559,N_483,N_476);
nor U560 (N_560,N_479,N_462);
or U561 (N_561,N_454,N_477);
nand U562 (N_562,N_520,N_507);
or U563 (N_563,N_501,N_502);
nand U564 (N_564,N_466,N_521);
or U565 (N_565,N_491,N_496);
or U566 (N_566,N_488,N_514);
nand U567 (N_567,N_472,N_507);
or U568 (N_568,N_516,N_469);
and U569 (N_569,N_495,N_513);
and U570 (N_570,N_458,N_502);
or U571 (N_571,N_473,N_484);
nand U572 (N_572,N_477,N_495);
or U573 (N_573,N_467,N_488);
nor U574 (N_574,N_489,N_468);
nand U575 (N_575,N_486,N_462);
nand U576 (N_576,N_508,N_500);
xnor U577 (N_577,N_520,N_475);
nand U578 (N_578,N_463,N_495);
nor U579 (N_579,N_500,N_518);
nand U580 (N_580,N_499,N_498);
or U581 (N_581,N_515,N_451);
xnor U582 (N_582,N_466,N_484);
xor U583 (N_583,N_501,N_519);
or U584 (N_584,N_523,N_472);
nand U585 (N_585,N_517,N_474);
nand U586 (N_586,N_521,N_476);
or U587 (N_587,N_456,N_491);
and U588 (N_588,N_512,N_517);
or U589 (N_589,N_496,N_479);
or U590 (N_590,N_473,N_456);
nor U591 (N_591,N_490,N_504);
nand U592 (N_592,N_489,N_521);
or U593 (N_593,N_520,N_502);
and U594 (N_594,N_454,N_507);
or U595 (N_595,N_500,N_477);
nand U596 (N_596,N_490,N_461);
and U597 (N_597,N_460,N_493);
and U598 (N_598,N_470,N_462);
nand U599 (N_599,N_468,N_462);
or U600 (N_600,N_588,N_549);
and U601 (N_601,N_575,N_547);
nor U602 (N_602,N_553,N_538);
or U603 (N_603,N_541,N_569);
nor U604 (N_604,N_579,N_552);
nor U605 (N_605,N_544,N_576);
or U606 (N_606,N_559,N_581);
and U607 (N_607,N_561,N_591);
nor U608 (N_608,N_599,N_545);
or U609 (N_609,N_537,N_551);
or U610 (N_610,N_596,N_528);
xnor U611 (N_611,N_539,N_595);
nand U612 (N_612,N_585,N_555);
and U613 (N_613,N_587,N_556);
nand U614 (N_614,N_540,N_583);
and U615 (N_615,N_527,N_570);
or U616 (N_616,N_546,N_574);
or U617 (N_617,N_568,N_542);
and U618 (N_618,N_598,N_560);
and U619 (N_619,N_526,N_531);
nand U620 (N_620,N_550,N_525);
nor U621 (N_621,N_597,N_586);
nand U622 (N_622,N_562,N_532);
nand U623 (N_623,N_557,N_543);
and U624 (N_624,N_582,N_584);
nor U625 (N_625,N_572,N_573);
and U626 (N_626,N_565,N_580);
nand U627 (N_627,N_534,N_577);
or U628 (N_628,N_536,N_530);
or U629 (N_629,N_558,N_533);
and U630 (N_630,N_594,N_564);
nor U631 (N_631,N_590,N_563);
and U632 (N_632,N_589,N_571);
or U633 (N_633,N_535,N_578);
or U634 (N_634,N_529,N_592);
and U635 (N_635,N_548,N_566);
nor U636 (N_636,N_567,N_554);
or U637 (N_637,N_593,N_535);
nand U638 (N_638,N_572,N_598);
nor U639 (N_639,N_590,N_593);
nor U640 (N_640,N_541,N_573);
nand U641 (N_641,N_590,N_564);
xnor U642 (N_642,N_567,N_565);
nand U643 (N_643,N_526,N_574);
nand U644 (N_644,N_569,N_534);
nand U645 (N_645,N_536,N_543);
nand U646 (N_646,N_540,N_594);
or U647 (N_647,N_545,N_547);
and U648 (N_648,N_560,N_536);
and U649 (N_649,N_531,N_567);
nand U650 (N_650,N_566,N_597);
nor U651 (N_651,N_548,N_599);
nor U652 (N_652,N_579,N_562);
nand U653 (N_653,N_538,N_589);
nor U654 (N_654,N_585,N_568);
or U655 (N_655,N_567,N_575);
nor U656 (N_656,N_595,N_544);
and U657 (N_657,N_579,N_554);
and U658 (N_658,N_541,N_533);
or U659 (N_659,N_532,N_599);
nor U660 (N_660,N_553,N_563);
or U661 (N_661,N_527,N_580);
nand U662 (N_662,N_598,N_569);
and U663 (N_663,N_534,N_557);
or U664 (N_664,N_537,N_555);
nor U665 (N_665,N_538,N_574);
or U666 (N_666,N_585,N_550);
nand U667 (N_667,N_570,N_573);
nand U668 (N_668,N_588,N_540);
nand U669 (N_669,N_541,N_585);
or U670 (N_670,N_579,N_556);
nand U671 (N_671,N_598,N_565);
nand U672 (N_672,N_549,N_560);
nand U673 (N_673,N_541,N_581);
and U674 (N_674,N_540,N_599);
nor U675 (N_675,N_611,N_673);
nand U676 (N_676,N_627,N_653);
or U677 (N_677,N_624,N_615);
or U678 (N_678,N_648,N_650);
nor U679 (N_679,N_618,N_643);
and U680 (N_680,N_667,N_633);
nand U681 (N_681,N_610,N_614);
or U682 (N_682,N_634,N_606);
or U683 (N_683,N_602,N_639);
nor U684 (N_684,N_670,N_630);
and U685 (N_685,N_654,N_638);
nand U686 (N_686,N_647,N_623);
nand U687 (N_687,N_626,N_669);
nor U688 (N_688,N_604,N_635);
or U689 (N_689,N_636,N_620);
nor U690 (N_690,N_663,N_655);
nor U691 (N_691,N_652,N_666);
or U692 (N_692,N_605,N_645);
or U693 (N_693,N_600,N_612);
or U694 (N_694,N_658,N_674);
or U695 (N_695,N_661,N_603);
nand U696 (N_696,N_660,N_613);
nor U697 (N_697,N_601,N_631);
nand U698 (N_698,N_659,N_616);
and U699 (N_699,N_651,N_642);
xnor U700 (N_700,N_632,N_668);
nand U701 (N_701,N_664,N_640);
nor U702 (N_702,N_672,N_649);
or U703 (N_703,N_662,N_637);
nand U704 (N_704,N_621,N_617);
and U705 (N_705,N_628,N_629);
nor U706 (N_706,N_646,N_665);
nor U707 (N_707,N_607,N_657);
nand U708 (N_708,N_608,N_622);
nand U709 (N_709,N_609,N_644);
nor U710 (N_710,N_671,N_619);
and U711 (N_711,N_656,N_625);
nor U712 (N_712,N_641,N_609);
and U713 (N_713,N_625,N_672);
or U714 (N_714,N_669,N_635);
xnor U715 (N_715,N_614,N_666);
nor U716 (N_716,N_637,N_630);
or U717 (N_717,N_650,N_667);
or U718 (N_718,N_604,N_660);
or U719 (N_719,N_635,N_600);
nor U720 (N_720,N_637,N_609);
and U721 (N_721,N_670,N_659);
and U722 (N_722,N_667,N_661);
nand U723 (N_723,N_609,N_612);
or U724 (N_724,N_674,N_629);
nand U725 (N_725,N_670,N_650);
or U726 (N_726,N_600,N_602);
nand U727 (N_727,N_613,N_609);
or U728 (N_728,N_673,N_640);
nand U729 (N_729,N_614,N_634);
or U730 (N_730,N_662,N_625);
and U731 (N_731,N_618,N_636);
nand U732 (N_732,N_663,N_603);
nand U733 (N_733,N_620,N_641);
nand U734 (N_734,N_668,N_649);
and U735 (N_735,N_667,N_654);
or U736 (N_736,N_625,N_604);
and U737 (N_737,N_666,N_621);
and U738 (N_738,N_669,N_621);
nor U739 (N_739,N_619,N_639);
or U740 (N_740,N_636,N_634);
and U741 (N_741,N_659,N_625);
or U742 (N_742,N_649,N_631);
nor U743 (N_743,N_625,N_623);
nand U744 (N_744,N_663,N_641);
nor U745 (N_745,N_630,N_610);
and U746 (N_746,N_649,N_600);
nor U747 (N_747,N_622,N_628);
nor U748 (N_748,N_629,N_655);
or U749 (N_749,N_622,N_607);
and U750 (N_750,N_686,N_727);
and U751 (N_751,N_695,N_729);
or U752 (N_752,N_737,N_676);
and U753 (N_753,N_678,N_723);
nor U754 (N_754,N_707,N_748);
and U755 (N_755,N_725,N_742);
and U756 (N_756,N_680,N_714);
and U757 (N_757,N_743,N_710);
nand U758 (N_758,N_708,N_717);
nand U759 (N_759,N_704,N_682);
or U760 (N_760,N_681,N_689);
nor U761 (N_761,N_687,N_694);
and U762 (N_762,N_745,N_684);
and U763 (N_763,N_732,N_702);
and U764 (N_764,N_711,N_736);
nor U765 (N_765,N_744,N_738);
nand U766 (N_766,N_697,N_740);
and U767 (N_767,N_709,N_685);
nor U768 (N_768,N_715,N_749);
or U769 (N_769,N_730,N_683);
nor U770 (N_770,N_735,N_741);
nand U771 (N_771,N_690,N_719);
nor U772 (N_772,N_747,N_679);
nand U773 (N_773,N_700,N_718);
nor U774 (N_774,N_731,N_706);
nor U775 (N_775,N_705,N_728);
or U776 (N_776,N_720,N_722);
or U777 (N_777,N_746,N_712);
and U778 (N_778,N_691,N_726);
nand U779 (N_779,N_688,N_701);
and U780 (N_780,N_699,N_692);
nor U781 (N_781,N_696,N_739);
or U782 (N_782,N_677,N_698);
or U783 (N_783,N_721,N_675);
and U784 (N_784,N_693,N_716);
nand U785 (N_785,N_724,N_733);
nor U786 (N_786,N_713,N_703);
nand U787 (N_787,N_734,N_730);
nand U788 (N_788,N_722,N_698);
nor U789 (N_789,N_693,N_709);
and U790 (N_790,N_745,N_689);
nor U791 (N_791,N_740,N_707);
nand U792 (N_792,N_701,N_680);
nand U793 (N_793,N_705,N_688);
nor U794 (N_794,N_728,N_682);
or U795 (N_795,N_695,N_733);
nor U796 (N_796,N_721,N_682);
or U797 (N_797,N_745,N_678);
or U798 (N_798,N_737,N_709);
or U799 (N_799,N_719,N_721);
nand U800 (N_800,N_691,N_729);
and U801 (N_801,N_735,N_698);
nand U802 (N_802,N_698,N_718);
and U803 (N_803,N_729,N_722);
and U804 (N_804,N_679,N_701);
nand U805 (N_805,N_731,N_689);
nor U806 (N_806,N_727,N_749);
nor U807 (N_807,N_740,N_688);
or U808 (N_808,N_689,N_704);
nor U809 (N_809,N_686,N_740);
or U810 (N_810,N_746,N_718);
nor U811 (N_811,N_698,N_743);
or U812 (N_812,N_729,N_732);
nor U813 (N_813,N_742,N_685);
nand U814 (N_814,N_702,N_738);
nor U815 (N_815,N_693,N_721);
or U816 (N_816,N_710,N_698);
xnor U817 (N_817,N_696,N_744);
and U818 (N_818,N_732,N_723);
nand U819 (N_819,N_726,N_701);
or U820 (N_820,N_717,N_735);
and U821 (N_821,N_685,N_708);
or U822 (N_822,N_714,N_719);
nand U823 (N_823,N_749,N_729);
and U824 (N_824,N_729,N_678);
and U825 (N_825,N_796,N_758);
or U826 (N_826,N_823,N_802);
or U827 (N_827,N_819,N_790);
nor U828 (N_828,N_811,N_767);
nor U829 (N_829,N_773,N_763);
or U830 (N_830,N_751,N_768);
nor U831 (N_831,N_762,N_822);
or U832 (N_832,N_769,N_775);
nor U833 (N_833,N_760,N_753);
and U834 (N_834,N_815,N_817);
nor U835 (N_835,N_777,N_772);
nand U836 (N_836,N_810,N_788);
nor U837 (N_837,N_774,N_752);
or U838 (N_838,N_809,N_807);
nand U839 (N_839,N_771,N_795);
or U840 (N_840,N_800,N_770);
nand U841 (N_841,N_820,N_818);
or U842 (N_842,N_798,N_761);
or U843 (N_843,N_814,N_801);
or U844 (N_844,N_757,N_797);
nand U845 (N_845,N_759,N_776);
and U846 (N_846,N_766,N_750);
and U847 (N_847,N_787,N_803);
nor U848 (N_848,N_813,N_824);
nor U849 (N_849,N_754,N_808);
and U850 (N_850,N_816,N_778);
nor U851 (N_851,N_765,N_821);
nand U852 (N_852,N_806,N_755);
or U853 (N_853,N_791,N_785);
xor U854 (N_854,N_805,N_812);
or U855 (N_855,N_756,N_794);
and U856 (N_856,N_789,N_786);
nor U857 (N_857,N_782,N_764);
nand U858 (N_858,N_779,N_780);
and U859 (N_859,N_799,N_792);
or U860 (N_860,N_781,N_804);
nand U861 (N_861,N_783,N_784);
or U862 (N_862,N_793,N_809);
and U863 (N_863,N_811,N_787);
and U864 (N_864,N_801,N_781);
nor U865 (N_865,N_798,N_779);
or U866 (N_866,N_778,N_784);
nand U867 (N_867,N_776,N_753);
and U868 (N_868,N_819,N_775);
nor U869 (N_869,N_800,N_769);
and U870 (N_870,N_798,N_769);
nor U871 (N_871,N_782,N_812);
or U872 (N_872,N_763,N_802);
nor U873 (N_873,N_784,N_776);
or U874 (N_874,N_777,N_819);
nor U875 (N_875,N_755,N_823);
nor U876 (N_876,N_811,N_758);
nor U877 (N_877,N_814,N_771);
nor U878 (N_878,N_824,N_751);
and U879 (N_879,N_813,N_765);
nand U880 (N_880,N_808,N_758);
nand U881 (N_881,N_811,N_772);
nand U882 (N_882,N_751,N_808);
and U883 (N_883,N_751,N_805);
nor U884 (N_884,N_798,N_817);
nand U885 (N_885,N_782,N_787);
nor U886 (N_886,N_824,N_759);
nand U887 (N_887,N_772,N_805);
or U888 (N_888,N_764,N_789);
nand U889 (N_889,N_751,N_815);
nor U890 (N_890,N_774,N_794);
nand U891 (N_891,N_794,N_784);
nand U892 (N_892,N_755,N_797);
and U893 (N_893,N_787,N_777);
nand U894 (N_894,N_778,N_785);
nor U895 (N_895,N_788,N_804);
or U896 (N_896,N_752,N_807);
or U897 (N_897,N_799,N_797);
and U898 (N_898,N_750,N_776);
nor U899 (N_899,N_818,N_766);
nand U900 (N_900,N_860,N_873);
and U901 (N_901,N_870,N_849);
nor U902 (N_902,N_874,N_837);
or U903 (N_903,N_883,N_838);
and U904 (N_904,N_827,N_836);
nor U905 (N_905,N_884,N_862);
nand U906 (N_906,N_834,N_841);
and U907 (N_907,N_851,N_839);
xnor U908 (N_908,N_840,N_845);
or U909 (N_909,N_868,N_833);
nor U910 (N_910,N_867,N_855);
or U911 (N_911,N_881,N_826);
and U912 (N_912,N_858,N_897);
or U913 (N_913,N_877,N_842);
or U914 (N_914,N_888,N_843);
nor U915 (N_915,N_852,N_890);
nand U916 (N_916,N_898,N_848);
nor U917 (N_917,N_859,N_831);
nand U918 (N_918,N_895,N_871);
and U919 (N_919,N_879,N_861);
nor U920 (N_920,N_893,N_894);
or U921 (N_921,N_850,N_828);
and U922 (N_922,N_892,N_825);
and U923 (N_923,N_872,N_835);
or U924 (N_924,N_882,N_886);
nor U925 (N_925,N_847,N_891);
nand U926 (N_926,N_846,N_896);
and U927 (N_927,N_856,N_854);
nand U928 (N_928,N_864,N_880);
and U929 (N_929,N_853,N_863);
nor U930 (N_930,N_889,N_885);
nor U931 (N_931,N_878,N_830);
nor U932 (N_932,N_869,N_887);
nand U933 (N_933,N_876,N_899);
or U934 (N_934,N_875,N_829);
xor U935 (N_935,N_866,N_865);
nor U936 (N_936,N_857,N_844);
nor U937 (N_937,N_832,N_844);
and U938 (N_938,N_848,N_864);
nor U939 (N_939,N_862,N_871);
nand U940 (N_940,N_860,N_847);
xnor U941 (N_941,N_854,N_881);
or U942 (N_942,N_851,N_899);
nand U943 (N_943,N_825,N_873);
nor U944 (N_944,N_825,N_886);
nor U945 (N_945,N_829,N_899);
and U946 (N_946,N_874,N_829);
nand U947 (N_947,N_868,N_871);
nor U948 (N_948,N_855,N_895);
and U949 (N_949,N_898,N_893);
and U950 (N_950,N_894,N_873);
or U951 (N_951,N_828,N_888);
and U952 (N_952,N_868,N_884);
and U953 (N_953,N_825,N_845);
nor U954 (N_954,N_830,N_870);
nor U955 (N_955,N_837,N_863);
nor U956 (N_956,N_852,N_838);
nand U957 (N_957,N_869,N_866);
xor U958 (N_958,N_838,N_894);
nand U959 (N_959,N_887,N_842);
nand U960 (N_960,N_889,N_834);
nor U961 (N_961,N_842,N_850);
nand U962 (N_962,N_883,N_875);
or U963 (N_963,N_870,N_835);
and U964 (N_964,N_853,N_828);
nor U965 (N_965,N_843,N_855);
or U966 (N_966,N_871,N_894);
nand U967 (N_967,N_883,N_826);
and U968 (N_968,N_882,N_875);
or U969 (N_969,N_880,N_865);
and U970 (N_970,N_843,N_847);
or U971 (N_971,N_836,N_864);
or U972 (N_972,N_883,N_867);
nand U973 (N_973,N_835,N_862);
nor U974 (N_974,N_880,N_857);
and U975 (N_975,N_964,N_941);
nor U976 (N_976,N_970,N_926);
and U977 (N_977,N_912,N_911);
and U978 (N_978,N_917,N_960);
nor U979 (N_979,N_919,N_958);
nor U980 (N_980,N_973,N_938);
nor U981 (N_981,N_910,N_901);
or U982 (N_982,N_929,N_965);
and U983 (N_983,N_933,N_904);
and U984 (N_984,N_920,N_953);
or U985 (N_985,N_915,N_968);
or U986 (N_986,N_966,N_918);
nand U987 (N_987,N_907,N_913);
and U988 (N_988,N_930,N_932);
and U989 (N_989,N_944,N_936);
nand U990 (N_990,N_928,N_921);
and U991 (N_991,N_963,N_902);
nor U992 (N_992,N_948,N_952);
nor U993 (N_993,N_950,N_955);
nor U994 (N_994,N_931,N_906);
or U995 (N_995,N_914,N_934);
nand U996 (N_996,N_908,N_903);
nor U997 (N_997,N_945,N_909);
and U998 (N_998,N_961,N_967);
and U999 (N_999,N_916,N_949);
nand U1000 (N_1000,N_937,N_905);
or U1001 (N_1001,N_962,N_900);
or U1002 (N_1002,N_942,N_922);
or U1003 (N_1003,N_972,N_954);
nand U1004 (N_1004,N_925,N_974);
or U1005 (N_1005,N_971,N_947);
nor U1006 (N_1006,N_939,N_927);
xor U1007 (N_1007,N_957,N_943);
nand U1008 (N_1008,N_946,N_923);
or U1009 (N_1009,N_935,N_956);
nor U1010 (N_1010,N_951,N_924);
nor U1011 (N_1011,N_959,N_969);
nor U1012 (N_1012,N_940,N_970);
nand U1013 (N_1013,N_929,N_959);
and U1014 (N_1014,N_919,N_927);
or U1015 (N_1015,N_901,N_971);
nand U1016 (N_1016,N_955,N_923);
or U1017 (N_1017,N_956,N_946);
xnor U1018 (N_1018,N_961,N_902);
or U1019 (N_1019,N_953,N_930);
or U1020 (N_1020,N_944,N_926);
and U1021 (N_1021,N_932,N_952);
or U1022 (N_1022,N_967,N_969);
or U1023 (N_1023,N_932,N_968);
nor U1024 (N_1024,N_972,N_928);
or U1025 (N_1025,N_922,N_903);
or U1026 (N_1026,N_959,N_970);
and U1027 (N_1027,N_918,N_948);
or U1028 (N_1028,N_920,N_955);
or U1029 (N_1029,N_969,N_928);
nand U1030 (N_1030,N_905,N_929);
or U1031 (N_1031,N_913,N_952);
nand U1032 (N_1032,N_929,N_939);
nand U1033 (N_1033,N_963,N_931);
and U1034 (N_1034,N_939,N_915);
or U1035 (N_1035,N_917,N_937);
nor U1036 (N_1036,N_969,N_955);
xor U1037 (N_1037,N_923,N_951);
or U1038 (N_1038,N_928,N_965);
or U1039 (N_1039,N_973,N_910);
nor U1040 (N_1040,N_944,N_970);
nor U1041 (N_1041,N_940,N_947);
nand U1042 (N_1042,N_942,N_970);
nand U1043 (N_1043,N_952,N_936);
or U1044 (N_1044,N_955,N_953);
nor U1045 (N_1045,N_963,N_954);
nor U1046 (N_1046,N_901,N_943);
or U1047 (N_1047,N_959,N_902);
nand U1048 (N_1048,N_938,N_945);
or U1049 (N_1049,N_934,N_905);
xnor U1050 (N_1050,N_1030,N_1031);
or U1051 (N_1051,N_996,N_990);
nand U1052 (N_1052,N_1041,N_1023);
nand U1053 (N_1053,N_1021,N_1018);
nand U1054 (N_1054,N_978,N_976);
nor U1055 (N_1055,N_983,N_1045);
nor U1056 (N_1056,N_1014,N_1034);
nor U1057 (N_1057,N_1007,N_1039);
nand U1058 (N_1058,N_1024,N_1044);
and U1059 (N_1059,N_992,N_1025);
nand U1060 (N_1060,N_988,N_977);
nor U1061 (N_1061,N_982,N_1012);
and U1062 (N_1062,N_1011,N_1038);
and U1063 (N_1063,N_1005,N_1022);
nor U1064 (N_1064,N_993,N_1032);
or U1065 (N_1065,N_1010,N_1026);
nand U1066 (N_1066,N_1029,N_1002);
nor U1067 (N_1067,N_980,N_1049);
nor U1068 (N_1068,N_1013,N_1008);
and U1069 (N_1069,N_1016,N_994);
nor U1070 (N_1070,N_1048,N_1017);
nor U1071 (N_1071,N_1042,N_1015);
nand U1072 (N_1072,N_1000,N_1020);
nor U1073 (N_1073,N_1027,N_1009);
nand U1074 (N_1074,N_1004,N_1035);
and U1075 (N_1075,N_997,N_979);
and U1076 (N_1076,N_1040,N_1037);
nand U1077 (N_1077,N_1047,N_985);
nor U1078 (N_1078,N_975,N_1028);
or U1079 (N_1079,N_1046,N_995);
nand U1080 (N_1080,N_1006,N_981);
nand U1081 (N_1081,N_989,N_1036);
or U1082 (N_1082,N_986,N_1003);
nand U1083 (N_1083,N_999,N_998);
nand U1084 (N_1084,N_1001,N_991);
or U1085 (N_1085,N_1019,N_1043);
or U1086 (N_1086,N_1033,N_984);
nor U1087 (N_1087,N_987,N_1000);
nand U1088 (N_1088,N_1007,N_1045);
nand U1089 (N_1089,N_992,N_1033);
or U1090 (N_1090,N_1018,N_975);
nor U1091 (N_1091,N_1012,N_975);
nor U1092 (N_1092,N_982,N_986);
nor U1093 (N_1093,N_1001,N_997);
nand U1094 (N_1094,N_1004,N_991);
nand U1095 (N_1095,N_975,N_994);
or U1096 (N_1096,N_1044,N_1005);
or U1097 (N_1097,N_1044,N_983);
and U1098 (N_1098,N_995,N_993);
nand U1099 (N_1099,N_996,N_989);
nor U1100 (N_1100,N_995,N_1041);
or U1101 (N_1101,N_1025,N_999);
nand U1102 (N_1102,N_1041,N_1035);
nand U1103 (N_1103,N_978,N_1019);
or U1104 (N_1104,N_1031,N_1008);
or U1105 (N_1105,N_1044,N_998);
nor U1106 (N_1106,N_983,N_979);
nand U1107 (N_1107,N_1001,N_1018);
and U1108 (N_1108,N_993,N_1009);
nand U1109 (N_1109,N_1044,N_1030);
or U1110 (N_1110,N_1043,N_1022);
or U1111 (N_1111,N_1013,N_987);
nand U1112 (N_1112,N_977,N_1039);
nand U1113 (N_1113,N_1027,N_1010);
or U1114 (N_1114,N_1044,N_1010);
nor U1115 (N_1115,N_1016,N_1011);
and U1116 (N_1116,N_1038,N_1004);
or U1117 (N_1117,N_1007,N_1015);
or U1118 (N_1118,N_975,N_999);
and U1119 (N_1119,N_989,N_1018);
nor U1120 (N_1120,N_980,N_1023);
nor U1121 (N_1121,N_1001,N_978);
nand U1122 (N_1122,N_1038,N_1027);
xor U1123 (N_1123,N_981,N_1032);
xnor U1124 (N_1124,N_1036,N_1017);
and U1125 (N_1125,N_1114,N_1073);
nor U1126 (N_1126,N_1091,N_1102);
nand U1127 (N_1127,N_1074,N_1086);
or U1128 (N_1128,N_1084,N_1077);
nand U1129 (N_1129,N_1080,N_1053);
xnor U1130 (N_1130,N_1069,N_1093);
nor U1131 (N_1131,N_1097,N_1050);
nor U1132 (N_1132,N_1098,N_1120);
nor U1133 (N_1133,N_1063,N_1079);
nand U1134 (N_1134,N_1115,N_1111);
nand U1135 (N_1135,N_1068,N_1075);
nor U1136 (N_1136,N_1110,N_1090);
xnor U1137 (N_1137,N_1119,N_1101);
nor U1138 (N_1138,N_1055,N_1103);
nor U1139 (N_1139,N_1122,N_1118);
or U1140 (N_1140,N_1059,N_1051);
and U1141 (N_1141,N_1052,N_1082);
xor U1142 (N_1142,N_1070,N_1100);
and U1143 (N_1143,N_1076,N_1067);
or U1144 (N_1144,N_1078,N_1108);
and U1145 (N_1145,N_1089,N_1105);
and U1146 (N_1146,N_1057,N_1088);
nand U1147 (N_1147,N_1065,N_1061);
nor U1148 (N_1148,N_1094,N_1062);
or U1149 (N_1149,N_1058,N_1071);
nand U1150 (N_1150,N_1095,N_1104);
nor U1151 (N_1151,N_1121,N_1107);
nand U1152 (N_1152,N_1060,N_1085);
nor U1153 (N_1153,N_1113,N_1072);
nand U1154 (N_1154,N_1106,N_1092);
and U1155 (N_1155,N_1066,N_1081);
nor U1156 (N_1156,N_1096,N_1087);
and U1157 (N_1157,N_1112,N_1064);
nor U1158 (N_1158,N_1123,N_1117);
nor U1159 (N_1159,N_1054,N_1056);
nor U1160 (N_1160,N_1124,N_1109);
or U1161 (N_1161,N_1083,N_1116);
and U1162 (N_1162,N_1099,N_1123);
or U1163 (N_1163,N_1118,N_1103);
nand U1164 (N_1164,N_1094,N_1075);
nand U1165 (N_1165,N_1104,N_1101);
and U1166 (N_1166,N_1109,N_1113);
and U1167 (N_1167,N_1104,N_1066);
xnor U1168 (N_1168,N_1089,N_1056);
and U1169 (N_1169,N_1053,N_1102);
and U1170 (N_1170,N_1068,N_1101);
nor U1171 (N_1171,N_1110,N_1112);
nor U1172 (N_1172,N_1122,N_1061);
or U1173 (N_1173,N_1079,N_1062);
nor U1174 (N_1174,N_1124,N_1070);
and U1175 (N_1175,N_1116,N_1089);
nor U1176 (N_1176,N_1104,N_1074);
nor U1177 (N_1177,N_1094,N_1108);
nand U1178 (N_1178,N_1085,N_1120);
and U1179 (N_1179,N_1119,N_1055);
nor U1180 (N_1180,N_1087,N_1069);
or U1181 (N_1181,N_1087,N_1078);
or U1182 (N_1182,N_1112,N_1124);
or U1183 (N_1183,N_1080,N_1116);
or U1184 (N_1184,N_1112,N_1059);
nor U1185 (N_1185,N_1066,N_1122);
or U1186 (N_1186,N_1123,N_1106);
and U1187 (N_1187,N_1076,N_1088);
and U1188 (N_1188,N_1102,N_1052);
nand U1189 (N_1189,N_1082,N_1057);
nand U1190 (N_1190,N_1091,N_1058);
and U1191 (N_1191,N_1093,N_1099);
nand U1192 (N_1192,N_1084,N_1101);
and U1193 (N_1193,N_1118,N_1059);
or U1194 (N_1194,N_1085,N_1062);
xnor U1195 (N_1195,N_1102,N_1121);
nand U1196 (N_1196,N_1079,N_1122);
and U1197 (N_1197,N_1086,N_1093);
and U1198 (N_1198,N_1096,N_1062);
and U1199 (N_1199,N_1052,N_1077);
and U1200 (N_1200,N_1153,N_1169);
nor U1201 (N_1201,N_1143,N_1150);
and U1202 (N_1202,N_1171,N_1130);
and U1203 (N_1203,N_1176,N_1151);
and U1204 (N_1204,N_1175,N_1196);
nor U1205 (N_1205,N_1134,N_1132);
and U1206 (N_1206,N_1145,N_1154);
nor U1207 (N_1207,N_1165,N_1177);
or U1208 (N_1208,N_1136,N_1187);
xnor U1209 (N_1209,N_1185,N_1199);
and U1210 (N_1210,N_1139,N_1197);
and U1211 (N_1211,N_1180,N_1191);
xnor U1212 (N_1212,N_1174,N_1127);
nand U1213 (N_1213,N_1193,N_1182);
nor U1214 (N_1214,N_1157,N_1198);
nor U1215 (N_1215,N_1152,N_1162);
and U1216 (N_1216,N_1146,N_1163);
and U1217 (N_1217,N_1156,N_1161);
xnor U1218 (N_1218,N_1147,N_1184);
nand U1219 (N_1219,N_1144,N_1140);
nand U1220 (N_1220,N_1188,N_1138);
nand U1221 (N_1221,N_1186,N_1192);
and U1222 (N_1222,N_1131,N_1189);
or U1223 (N_1223,N_1195,N_1155);
nor U1224 (N_1224,N_1170,N_1135);
nand U1225 (N_1225,N_1128,N_1178);
and U1226 (N_1226,N_1190,N_1168);
nor U1227 (N_1227,N_1172,N_1125);
or U1228 (N_1228,N_1194,N_1129);
and U1229 (N_1229,N_1159,N_1183);
nor U1230 (N_1230,N_1166,N_1148);
nor U1231 (N_1231,N_1141,N_1158);
nor U1232 (N_1232,N_1160,N_1181);
nand U1233 (N_1233,N_1173,N_1137);
or U1234 (N_1234,N_1126,N_1142);
or U1235 (N_1235,N_1133,N_1164);
nor U1236 (N_1236,N_1167,N_1179);
or U1237 (N_1237,N_1149,N_1198);
nor U1238 (N_1238,N_1198,N_1184);
nor U1239 (N_1239,N_1178,N_1131);
nor U1240 (N_1240,N_1136,N_1125);
nor U1241 (N_1241,N_1173,N_1145);
nor U1242 (N_1242,N_1159,N_1195);
nand U1243 (N_1243,N_1140,N_1128);
nor U1244 (N_1244,N_1184,N_1175);
nand U1245 (N_1245,N_1133,N_1134);
or U1246 (N_1246,N_1184,N_1130);
xor U1247 (N_1247,N_1155,N_1197);
or U1248 (N_1248,N_1179,N_1182);
or U1249 (N_1249,N_1149,N_1128);
nor U1250 (N_1250,N_1157,N_1156);
or U1251 (N_1251,N_1181,N_1194);
or U1252 (N_1252,N_1156,N_1149);
or U1253 (N_1253,N_1155,N_1177);
nand U1254 (N_1254,N_1161,N_1151);
nand U1255 (N_1255,N_1140,N_1168);
nor U1256 (N_1256,N_1185,N_1191);
nand U1257 (N_1257,N_1158,N_1180);
or U1258 (N_1258,N_1145,N_1142);
nand U1259 (N_1259,N_1129,N_1162);
nor U1260 (N_1260,N_1163,N_1187);
nor U1261 (N_1261,N_1153,N_1183);
nand U1262 (N_1262,N_1137,N_1188);
nand U1263 (N_1263,N_1141,N_1152);
nand U1264 (N_1264,N_1186,N_1144);
or U1265 (N_1265,N_1145,N_1188);
or U1266 (N_1266,N_1146,N_1129);
and U1267 (N_1267,N_1138,N_1189);
and U1268 (N_1268,N_1165,N_1196);
nor U1269 (N_1269,N_1140,N_1141);
nand U1270 (N_1270,N_1137,N_1185);
nand U1271 (N_1271,N_1179,N_1156);
nand U1272 (N_1272,N_1196,N_1137);
or U1273 (N_1273,N_1145,N_1133);
and U1274 (N_1274,N_1166,N_1179);
or U1275 (N_1275,N_1229,N_1208);
nand U1276 (N_1276,N_1239,N_1260);
nor U1277 (N_1277,N_1270,N_1217);
or U1278 (N_1278,N_1272,N_1241);
and U1279 (N_1279,N_1228,N_1248);
and U1280 (N_1280,N_1243,N_1268);
nor U1281 (N_1281,N_1212,N_1221);
and U1282 (N_1282,N_1230,N_1265);
nand U1283 (N_1283,N_1262,N_1240);
or U1284 (N_1284,N_1252,N_1271);
nand U1285 (N_1285,N_1210,N_1201);
nor U1286 (N_1286,N_1238,N_1220);
nor U1287 (N_1287,N_1257,N_1224);
nor U1288 (N_1288,N_1273,N_1269);
or U1289 (N_1289,N_1261,N_1200);
nor U1290 (N_1290,N_1225,N_1207);
nand U1291 (N_1291,N_1250,N_1247);
or U1292 (N_1292,N_1244,N_1254);
nor U1293 (N_1293,N_1205,N_1226);
nand U1294 (N_1294,N_1234,N_1267);
or U1295 (N_1295,N_1258,N_1249);
or U1296 (N_1296,N_1203,N_1211);
and U1297 (N_1297,N_1235,N_1233);
and U1298 (N_1298,N_1259,N_1204);
nand U1299 (N_1299,N_1256,N_1218);
or U1300 (N_1300,N_1237,N_1231);
nand U1301 (N_1301,N_1214,N_1216);
and U1302 (N_1302,N_1253,N_1264);
or U1303 (N_1303,N_1223,N_1206);
and U1304 (N_1304,N_1219,N_1215);
or U1305 (N_1305,N_1274,N_1263);
or U1306 (N_1306,N_1213,N_1202);
nor U1307 (N_1307,N_1227,N_1232);
nand U1308 (N_1308,N_1209,N_1245);
and U1309 (N_1309,N_1255,N_1236);
or U1310 (N_1310,N_1251,N_1222);
or U1311 (N_1311,N_1266,N_1246);
or U1312 (N_1312,N_1242,N_1227);
or U1313 (N_1313,N_1237,N_1251);
or U1314 (N_1314,N_1233,N_1223);
nor U1315 (N_1315,N_1230,N_1249);
nand U1316 (N_1316,N_1244,N_1227);
nor U1317 (N_1317,N_1229,N_1263);
nand U1318 (N_1318,N_1222,N_1258);
and U1319 (N_1319,N_1249,N_1252);
nand U1320 (N_1320,N_1232,N_1258);
or U1321 (N_1321,N_1258,N_1224);
or U1322 (N_1322,N_1274,N_1240);
or U1323 (N_1323,N_1270,N_1222);
and U1324 (N_1324,N_1267,N_1259);
nand U1325 (N_1325,N_1234,N_1222);
nand U1326 (N_1326,N_1220,N_1202);
nor U1327 (N_1327,N_1236,N_1254);
nor U1328 (N_1328,N_1220,N_1250);
nand U1329 (N_1329,N_1273,N_1231);
nor U1330 (N_1330,N_1216,N_1228);
nand U1331 (N_1331,N_1222,N_1229);
nand U1332 (N_1332,N_1235,N_1201);
and U1333 (N_1333,N_1241,N_1244);
and U1334 (N_1334,N_1265,N_1273);
nand U1335 (N_1335,N_1272,N_1212);
or U1336 (N_1336,N_1251,N_1216);
xor U1337 (N_1337,N_1259,N_1211);
nand U1338 (N_1338,N_1200,N_1237);
xor U1339 (N_1339,N_1252,N_1227);
nor U1340 (N_1340,N_1216,N_1270);
or U1341 (N_1341,N_1242,N_1217);
nand U1342 (N_1342,N_1252,N_1229);
or U1343 (N_1343,N_1241,N_1212);
and U1344 (N_1344,N_1273,N_1244);
and U1345 (N_1345,N_1265,N_1204);
xor U1346 (N_1346,N_1238,N_1247);
nor U1347 (N_1347,N_1269,N_1272);
and U1348 (N_1348,N_1224,N_1214);
and U1349 (N_1349,N_1226,N_1206);
nand U1350 (N_1350,N_1304,N_1300);
nor U1351 (N_1351,N_1345,N_1284);
or U1352 (N_1352,N_1340,N_1299);
or U1353 (N_1353,N_1296,N_1335);
and U1354 (N_1354,N_1337,N_1326);
nor U1355 (N_1355,N_1292,N_1280);
or U1356 (N_1356,N_1324,N_1283);
or U1357 (N_1357,N_1276,N_1305);
nor U1358 (N_1358,N_1291,N_1302);
nand U1359 (N_1359,N_1329,N_1348);
or U1360 (N_1360,N_1334,N_1287);
nand U1361 (N_1361,N_1285,N_1311);
or U1362 (N_1362,N_1313,N_1306);
nand U1363 (N_1363,N_1327,N_1342);
or U1364 (N_1364,N_1316,N_1279);
nor U1365 (N_1365,N_1294,N_1318);
and U1366 (N_1366,N_1282,N_1330);
nand U1367 (N_1367,N_1312,N_1297);
or U1368 (N_1368,N_1320,N_1331);
nor U1369 (N_1369,N_1295,N_1310);
and U1370 (N_1370,N_1275,N_1290);
nor U1371 (N_1371,N_1303,N_1286);
nand U1372 (N_1372,N_1338,N_1315);
or U1373 (N_1373,N_1341,N_1346);
and U1374 (N_1374,N_1317,N_1301);
nor U1375 (N_1375,N_1321,N_1281);
or U1376 (N_1376,N_1309,N_1288);
nand U1377 (N_1377,N_1314,N_1332);
nor U1378 (N_1378,N_1328,N_1278);
and U1379 (N_1379,N_1347,N_1289);
nand U1380 (N_1380,N_1333,N_1298);
and U1381 (N_1381,N_1325,N_1307);
nor U1382 (N_1382,N_1344,N_1277);
and U1383 (N_1383,N_1322,N_1339);
nand U1384 (N_1384,N_1336,N_1349);
nand U1385 (N_1385,N_1343,N_1319);
nor U1386 (N_1386,N_1308,N_1293);
and U1387 (N_1387,N_1323,N_1327);
nand U1388 (N_1388,N_1296,N_1275);
nand U1389 (N_1389,N_1289,N_1312);
and U1390 (N_1390,N_1340,N_1343);
and U1391 (N_1391,N_1329,N_1335);
and U1392 (N_1392,N_1318,N_1302);
or U1393 (N_1393,N_1333,N_1339);
xor U1394 (N_1394,N_1275,N_1276);
or U1395 (N_1395,N_1275,N_1281);
or U1396 (N_1396,N_1281,N_1287);
nand U1397 (N_1397,N_1329,N_1349);
or U1398 (N_1398,N_1329,N_1299);
and U1399 (N_1399,N_1308,N_1294);
or U1400 (N_1400,N_1340,N_1331);
nor U1401 (N_1401,N_1308,N_1325);
and U1402 (N_1402,N_1317,N_1283);
nand U1403 (N_1403,N_1276,N_1310);
nor U1404 (N_1404,N_1325,N_1285);
and U1405 (N_1405,N_1276,N_1300);
or U1406 (N_1406,N_1276,N_1347);
or U1407 (N_1407,N_1324,N_1322);
nor U1408 (N_1408,N_1325,N_1295);
nand U1409 (N_1409,N_1344,N_1320);
or U1410 (N_1410,N_1321,N_1302);
nor U1411 (N_1411,N_1290,N_1323);
or U1412 (N_1412,N_1342,N_1298);
xnor U1413 (N_1413,N_1278,N_1316);
nor U1414 (N_1414,N_1345,N_1341);
and U1415 (N_1415,N_1321,N_1328);
nor U1416 (N_1416,N_1308,N_1323);
and U1417 (N_1417,N_1314,N_1308);
and U1418 (N_1418,N_1286,N_1329);
nand U1419 (N_1419,N_1319,N_1337);
and U1420 (N_1420,N_1279,N_1326);
nand U1421 (N_1421,N_1345,N_1333);
nor U1422 (N_1422,N_1277,N_1335);
nor U1423 (N_1423,N_1344,N_1302);
nand U1424 (N_1424,N_1304,N_1291);
xor U1425 (N_1425,N_1355,N_1383);
nor U1426 (N_1426,N_1413,N_1365);
or U1427 (N_1427,N_1404,N_1374);
nor U1428 (N_1428,N_1354,N_1376);
nor U1429 (N_1429,N_1380,N_1421);
and U1430 (N_1430,N_1361,N_1403);
and U1431 (N_1431,N_1424,N_1402);
and U1432 (N_1432,N_1381,N_1394);
nor U1433 (N_1433,N_1371,N_1399);
and U1434 (N_1434,N_1370,N_1360);
nor U1435 (N_1435,N_1351,N_1389);
or U1436 (N_1436,N_1411,N_1390);
nor U1437 (N_1437,N_1372,N_1418);
nor U1438 (N_1438,N_1419,N_1385);
nand U1439 (N_1439,N_1420,N_1416);
xnor U1440 (N_1440,N_1379,N_1368);
and U1441 (N_1441,N_1409,N_1414);
nand U1442 (N_1442,N_1364,N_1353);
nor U1443 (N_1443,N_1358,N_1408);
or U1444 (N_1444,N_1400,N_1369);
nor U1445 (N_1445,N_1412,N_1363);
and U1446 (N_1446,N_1392,N_1393);
nor U1447 (N_1447,N_1357,N_1366);
and U1448 (N_1448,N_1405,N_1396);
nand U1449 (N_1449,N_1417,N_1391);
nor U1450 (N_1450,N_1362,N_1378);
nor U1451 (N_1451,N_1386,N_1367);
nor U1452 (N_1452,N_1377,N_1387);
and U1453 (N_1453,N_1401,N_1422);
xor U1454 (N_1454,N_1382,N_1373);
or U1455 (N_1455,N_1352,N_1398);
nor U1456 (N_1456,N_1407,N_1350);
nor U1457 (N_1457,N_1410,N_1406);
nor U1458 (N_1458,N_1388,N_1359);
nand U1459 (N_1459,N_1384,N_1356);
nor U1460 (N_1460,N_1397,N_1415);
or U1461 (N_1461,N_1423,N_1375);
and U1462 (N_1462,N_1395,N_1386);
nand U1463 (N_1463,N_1390,N_1408);
and U1464 (N_1464,N_1398,N_1416);
nand U1465 (N_1465,N_1397,N_1416);
nand U1466 (N_1466,N_1395,N_1374);
nor U1467 (N_1467,N_1356,N_1367);
or U1468 (N_1468,N_1350,N_1358);
nor U1469 (N_1469,N_1367,N_1396);
nor U1470 (N_1470,N_1423,N_1424);
and U1471 (N_1471,N_1359,N_1354);
and U1472 (N_1472,N_1364,N_1402);
nor U1473 (N_1473,N_1411,N_1394);
nor U1474 (N_1474,N_1399,N_1418);
or U1475 (N_1475,N_1409,N_1422);
nor U1476 (N_1476,N_1362,N_1366);
nand U1477 (N_1477,N_1394,N_1424);
nor U1478 (N_1478,N_1356,N_1390);
and U1479 (N_1479,N_1355,N_1419);
nor U1480 (N_1480,N_1355,N_1371);
nor U1481 (N_1481,N_1372,N_1368);
or U1482 (N_1482,N_1407,N_1362);
or U1483 (N_1483,N_1398,N_1377);
nand U1484 (N_1484,N_1396,N_1351);
nor U1485 (N_1485,N_1376,N_1389);
nand U1486 (N_1486,N_1396,N_1411);
and U1487 (N_1487,N_1384,N_1424);
and U1488 (N_1488,N_1371,N_1368);
or U1489 (N_1489,N_1389,N_1368);
and U1490 (N_1490,N_1381,N_1404);
xor U1491 (N_1491,N_1378,N_1420);
or U1492 (N_1492,N_1406,N_1391);
nor U1493 (N_1493,N_1364,N_1362);
nor U1494 (N_1494,N_1415,N_1371);
or U1495 (N_1495,N_1416,N_1403);
nor U1496 (N_1496,N_1421,N_1371);
nor U1497 (N_1497,N_1395,N_1401);
nand U1498 (N_1498,N_1363,N_1385);
nand U1499 (N_1499,N_1381,N_1408);
nor U1500 (N_1500,N_1497,N_1429);
nand U1501 (N_1501,N_1465,N_1469);
or U1502 (N_1502,N_1425,N_1494);
and U1503 (N_1503,N_1478,N_1464);
or U1504 (N_1504,N_1484,N_1479);
or U1505 (N_1505,N_1434,N_1486);
and U1506 (N_1506,N_1450,N_1485);
and U1507 (N_1507,N_1431,N_1452);
nand U1508 (N_1508,N_1438,N_1490);
and U1509 (N_1509,N_1448,N_1493);
and U1510 (N_1510,N_1488,N_1468);
and U1511 (N_1511,N_1447,N_1461);
or U1512 (N_1512,N_1445,N_1428);
nor U1513 (N_1513,N_1474,N_1483);
or U1514 (N_1514,N_1454,N_1499);
or U1515 (N_1515,N_1432,N_1487);
or U1516 (N_1516,N_1457,N_1440);
xor U1517 (N_1517,N_1456,N_1459);
or U1518 (N_1518,N_1430,N_1463);
and U1519 (N_1519,N_1427,N_1426);
or U1520 (N_1520,N_1489,N_1491);
nor U1521 (N_1521,N_1453,N_1441);
and U1522 (N_1522,N_1442,N_1498);
nor U1523 (N_1523,N_1467,N_1496);
nand U1524 (N_1524,N_1475,N_1471);
and U1525 (N_1525,N_1492,N_1477);
nor U1526 (N_1526,N_1472,N_1495);
and U1527 (N_1527,N_1443,N_1451);
and U1528 (N_1528,N_1460,N_1444);
nand U1529 (N_1529,N_1476,N_1482);
nor U1530 (N_1530,N_1473,N_1458);
and U1531 (N_1531,N_1455,N_1466);
nand U1532 (N_1532,N_1433,N_1446);
and U1533 (N_1533,N_1436,N_1437);
and U1534 (N_1534,N_1439,N_1480);
nand U1535 (N_1535,N_1449,N_1470);
nor U1536 (N_1536,N_1435,N_1462);
or U1537 (N_1537,N_1481,N_1453);
nor U1538 (N_1538,N_1499,N_1463);
nand U1539 (N_1539,N_1431,N_1494);
or U1540 (N_1540,N_1496,N_1440);
and U1541 (N_1541,N_1460,N_1499);
nor U1542 (N_1542,N_1435,N_1448);
or U1543 (N_1543,N_1458,N_1466);
xnor U1544 (N_1544,N_1478,N_1458);
nand U1545 (N_1545,N_1488,N_1479);
nor U1546 (N_1546,N_1463,N_1495);
and U1547 (N_1547,N_1447,N_1444);
or U1548 (N_1548,N_1469,N_1449);
nor U1549 (N_1549,N_1476,N_1459);
and U1550 (N_1550,N_1430,N_1445);
and U1551 (N_1551,N_1497,N_1430);
and U1552 (N_1552,N_1486,N_1488);
nand U1553 (N_1553,N_1477,N_1491);
or U1554 (N_1554,N_1475,N_1438);
nor U1555 (N_1555,N_1463,N_1447);
or U1556 (N_1556,N_1439,N_1464);
or U1557 (N_1557,N_1449,N_1448);
xnor U1558 (N_1558,N_1459,N_1488);
nand U1559 (N_1559,N_1496,N_1443);
nor U1560 (N_1560,N_1498,N_1428);
and U1561 (N_1561,N_1446,N_1481);
and U1562 (N_1562,N_1446,N_1480);
nand U1563 (N_1563,N_1427,N_1463);
nor U1564 (N_1564,N_1464,N_1491);
nand U1565 (N_1565,N_1448,N_1494);
and U1566 (N_1566,N_1459,N_1497);
or U1567 (N_1567,N_1425,N_1440);
nand U1568 (N_1568,N_1451,N_1466);
nand U1569 (N_1569,N_1426,N_1457);
or U1570 (N_1570,N_1434,N_1495);
and U1571 (N_1571,N_1432,N_1473);
nor U1572 (N_1572,N_1469,N_1478);
or U1573 (N_1573,N_1476,N_1493);
nand U1574 (N_1574,N_1433,N_1469);
nand U1575 (N_1575,N_1514,N_1550);
nand U1576 (N_1576,N_1563,N_1552);
and U1577 (N_1577,N_1512,N_1541);
and U1578 (N_1578,N_1569,N_1533);
nor U1579 (N_1579,N_1502,N_1527);
nand U1580 (N_1580,N_1556,N_1510);
nand U1581 (N_1581,N_1543,N_1534);
and U1582 (N_1582,N_1562,N_1547);
or U1583 (N_1583,N_1515,N_1546);
and U1584 (N_1584,N_1509,N_1518);
xor U1585 (N_1585,N_1507,N_1549);
nand U1586 (N_1586,N_1525,N_1532);
and U1587 (N_1587,N_1523,N_1528);
nor U1588 (N_1588,N_1542,N_1567);
nor U1589 (N_1589,N_1568,N_1572);
nand U1590 (N_1590,N_1560,N_1548);
xor U1591 (N_1591,N_1536,N_1551);
and U1592 (N_1592,N_1516,N_1503);
or U1593 (N_1593,N_1565,N_1555);
nor U1594 (N_1594,N_1530,N_1564);
and U1595 (N_1595,N_1561,N_1539);
nand U1596 (N_1596,N_1521,N_1501);
nor U1597 (N_1597,N_1540,N_1570);
nand U1598 (N_1598,N_1537,N_1506);
nor U1599 (N_1599,N_1544,N_1500);
and U1600 (N_1600,N_1538,N_1526);
nand U1601 (N_1601,N_1511,N_1553);
and U1602 (N_1602,N_1535,N_1558);
and U1603 (N_1603,N_1566,N_1524);
nor U1604 (N_1604,N_1545,N_1557);
or U1605 (N_1605,N_1504,N_1573);
and U1606 (N_1606,N_1522,N_1531);
or U1607 (N_1607,N_1517,N_1519);
or U1608 (N_1608,N_1559,N_1554);
xnor U1609 (N_1609,N_1520,N_1571);
nor U1610 (N_1610,N_1508,N_1505);
nand U1611 (N_1611,N_1513,N_1529);
nor U1612 (N_1612,N_1574,N_1550);
nor U1613 (N_1613,N_1549,N_1540);
nor U1614 (N_1614,N_1545,N_1569);
or U1615 (N_1615,N_1565,N_1542);
nor U1616 (N_1616,N_1556,N_1507);
nand U1617 (N_1617,N_1500,N_1533);
or U1618 (N_1618,N_1571,N_1516);
nor U1619 (N_1619,N_1560,N_1510);
and U1620 (N_1620,N_1554,N_1522);
and U1621 (N_1621,N_1558,N_1528);
or U1622 (N_1622,N_1540,N_1572);
and U1623 (N_1623,N_1559,N_1533);
nand U1624 (N_1624,N_1552,N_1556);
nand U1625 (N_1625,N_1562,N_1501);
or U1626 (N_1626,N_1540,N_1562);
or U1627 (N_1627,N_1532,N_1573);
and U1628 (N_1628,N_1533,N_1562);
nor U1629 (N_1629,N_1558,N_1531);
nor U1630 (N_1630,N_1559,N_1537);
or U1631 (N_1631,N_1521,N_1509);
and U1632 (N_1632,N_1513,N_1528);
or U1633 (N_1633,N_1574,N_1559);
nand U1634 (N_1634,N_1554,N_1520);
nor U1635 (N_1635,N_1557,N_1507);
and U1636 (N_1636,N_1503,N_1524);
or U1637 (N_1637,N_1544,N_1521);
nand U1638 (N_1638,N_1549,N_1506);
or U1639 (N_1639,N_1501,N_1506);
nor U1640 (N_1640,N_1540,N_1522);
or U1641 (N_1641,N_1574,N_1566);
or U1642 (N_1642,N_1555,N_1543);
nand U1643 (N_1643,N_1568,N_1557);
nor U1644 (N_1644,N_1555,N_1541);
nand U1645 (N_1645,N_1566,N_1504);
nand U1646 (N_1646,N_1539,N_1500);
nand U1647 (N_1647,N_1562,N_1539);
and U1648 (N_1648,N_1510,N_1544);
and U1649 (N_1649,N_1540,N_1569);
or U1650 (N_1650,N_1626,N_1636);
nor U1651 (N_1651,N_1646,N_1648);
or U1652 (N_1652,N_1589,N_1598);
nor U1653 (N_1653,N_1588,N_1639);
nor U1654 (N_1654,N_1624,N_1611);
and U1655 (N_1655,N_1647,N_1620);
or U1656 (N_1656,N_1605,N_1590);
and U1657 (N_1657,N_1618,N_1621);
or U1658 (N_1658,N_1633,N_1641);
nor U1659 (N_1659,N_1616,N_1630);
nor U1660 (N_1660,N_1577,N_1643);
and U1661 (N_1661,N_1600,N_1603);
or U1662 (N_1662,N_1596,N_1649);
and U1663 (N_1663,N_1593,N_1617);
nand U1664 (N_1664,N_1608,N_1613);
nand U1665 (N_1665,N_1595,N_1585);
and U1666 (N_1666,N_1586,N_1582);
nand U1667 (N_1667,N_1602,N_1599);
or U1668 (N_1668,N_1592,N_1637);
and U1669 (N_1669,N_1612,N_1629);
or U1670 (N_1670,N_1578,N_1607);
and U1671 (N_1671,N_1622,N_1623);
nor U1672 (N_1672,N_1581,N_1583);
nor U1673 (N_1673,N_1619,N_1587);
or U1674 (N_1674,N_1601,N_1597);
nor U1675 (N_1675,N_1632,N_1604);
xor U1676 (N_1676,N_1635,N_1614);
nor U1677 (N_1677,N_1628,N_1625);
or U1678 (N_1678,N_1640,N_1638);
or U1679 (N_1679,N_1584,N_1645);
nand U1680 (N_1680,N_1606,N_1634);
and U1681 (N_1681,N_1615,N_1642);
nor U1682 (N_1682,N_1627,N_1609);
nor U1683 (N_1683,N_1579,N_1591);
nand U1684 (N_1684,N_1580,N_1610);
or U1685 (N_1685,N_1575,N_1631);
nor U1686 (N_1686,N_1644,N_1594);
nand U1687 (N_1687,N_1576,N_1594);
nor U1688 (N_1688,N_1636,N_1629);
or U1689 (N_1689,N_1619,N_1618);
nor U1690 (N_1690,N_1586,N_1600);
or U1691 (N_1691,N_1592,N_1610);
and U1692 (N_1692,N_1635,N_1634);
and U1693 (N_1693,N_1607,N_1591);
or U1694 (N_1694,N_1612,N_1645);
or U1695 (N_1695,N_1645,N_1647);
nor U1696 (N_1696,N_1642,N_1586);
nand U1697 (N_1697,N_1618,N_1577);
or U1698 (N_1698,N_1625,N_1592);
or U1699 (N_1699,N_1605,N_1635);
nor U1700 (N_1700,N_1597,N_1635);
nand U1701 (N_1701,N_1640,N_1602);
nand U1702 (N_1702,N_1628,N_1588);
and U1703 (N_1703,N_1646,N_1622);
or U1704 (N_1704,N_1623,N_1575);
xor U1705 (N_1705,N_1596,N_1591);
and U1706 (N_1706,N_1613,N_1584);
nand U1707 (N_1707,N_1586,N_1639);
nand U1708 (N_1708,N_1628,N_1629);
nand U1709 (N_1709,N_1575,N_1594);
nor U1710 (N_1710,N_1621,N_1649);
nand U1711 (N_1711,N_1596,N_1637);
nand U1712 (N_1712,N_1615,N_1619);
nor U1713 (N_1713,N_1619,N_1632);
or U1714 (N_1714,N_1649,N_1578);
or U1715 (N_1715,N_1625,N_1582);
nand U1716 (N_1716,N_1616,N_1637);
and U1717 (N_1717,N_1589,N_1595);
or U1718 (N_1718,N_1642,N_1645);
or U1719 (N_1719,N_1606,N_1627);
nand U1720 (N_1720,N_1610,N_1603);
or U1721 (N_1721,N_1623,N_1579);
nand U1722 (N_1722,N_1620,N_1600);
nand U1723 (N_1723,N_1607,N_1601);
or U1724 (N_1724,N_1576,N_1598);
and U1725 (N_1725,N_1663,N_1652);
or U1726 (N_1726,N_1661,N_1676);
and U1727 (N_1727,N_1656,N_1677);
nor U1728 (N_1728,N_1658,N_1702);
nor U1729 (N_1729,N_1693,N_1651);
and U1730 (N_1730,N_1691,N_1720);
or U1731 (N_1731,N_1669,N_1674);
nor U1732 (N_1732,N_1710,N_1711);
nor U1733 (N_1733,N_1706,N_1650);
nor U1734 (N_1734,N_1707,N_1662);
or U1735 (N_1735,N_1698,N_1708);
nor U1736 (N_1736,N_1714,N_1681);
or U1737 (N_1737,N_1696,N_1694);
and U1738 (N_1738,N_1709,N_1667);
or U1739 (N_1739,N_1705,N_1657);
or U1740 (N_1740,N_1689,N_1723);
or U1741 (N_1741,N_1703,N_1686);
or U1742 (N_1742,N_1716,N_1688);
nor U1743 (N_1743,N_1704,N_1685);
and U1744 (N_1744,N_1680,N_1695);
nor U1745 (N_1745,N_1713,N_1721);
nor U1746 (N_1746,N_1668,N_1665);
nor U1747 (N_1747,N_1679,N_1715);
nor U1748 (N_1748,N_1699,N_1670);
nor U1749 (N_1749,N_1683,N_1724);
nand U1750 (N_1750,N_1671,N_1700);
or U1751 (N_1751,N_1664,N_1655);
or U1752 (N_1752,N_1717,N_1654);
nand U1753 (N_1753,N_1690,N_1712);
and U1754 (N_1754,N_1673,N_1675);
nor U1755 (N_1755,N_1659,N_1684);
or U1756 (N_1756,N_1672,N_1722);
nor U1757 (N_1757,N_1697,N_1718);
or U1758 (N_1758,N_1682,N_1678);
and U1759 (N_1759,N_1653,N_1692);
nand U1760 (N_1760,N_1701,N_1687);
or U1761 (N_1761,N_1666,N_1719);
nor U1762 (N_1762,N_1660,N_1675);
or U1763 (N_1763,N_1669,N_1695);
or U1764 (N_1764,N_1684,N_1694);
xor U1765 (N_1765,N_1696,N_1705);
and U1766 (N_1766,N_1712,N_1675);
or U1767 (N_1767,N_1707,N_1705);
nand U1768 (N_1768,N_1724,N_1710);
or U1769 (N_1769,N_1706,N_1703);
nand U1770 (N_1770,N_1676,N_1654);
nand U1771 (N_1771,N_1694,N_1682);
or U1772 (N_1772,N_1656,N_1699);
nand U1773 (N_1773,N_1721,N_1653);
nand U1774 (N_1774,N_1672,N_1666);
nand U1775 (N_1775,N_1678,N_1721);
nor U1776 (N_1776,N_1693,N_1656);
nand U1777 (N_1777,N_1651,N_1672);
or U1778 (N_1778,N_1672,N_1705);
nand U1779 (N_1779,N_1705,N_1708);
nand U1780 (N_1780,N_1711,N_1686);
or U1781 (N_1781,N_1702,N_1682);
or U1782 (N_1782,N_1665,N_1702);
and U1783 (N_1783,N_1672,N_1709);
nand U1784 (N_1784,N_1670,N_1708);
nand U1785 (N_1785,N_1651,N_1655);
nor U1786 (N_1786,N_1709,N_1722);
nor U1787 (N_1787,N_1653,N_1709);
nand U1788 (N_1788,N_1688,N_1664);
nand U1789 (N_1789,N_1675,N_1705);
or U1790 (N_1790,N_1651,N_1702);
or U1791 (N_1791,N_1678,N_1651);
nand U1792 (N_1792,N_1676,N_1691);
nand U1793 (N_1793,N_1706,N_1724);
nor U1794 (N_1794,N_1675,N_1710);
nand U1795 (N_1795,N_1701,N_1681);
and U1796 (N_1796,N_1679,N_1656);
nand U1797 (N_1797,N_1691,N_1671);
and U1798 (N_1798,N_1709,N_1658);
xor U1799 (N_1799,N_1705,N_1693);
nand U1800 (N_1800,N_1761,N_1793);
nor U1801 (N_1801,N_1792,N_1777);
nor U1802 (N_1802,N_1752,N_1795);
nor U1803 (N_1803,N_1775,N_1783);
or U1804 (N_1804,N_1726,N_1727);
and U1805 (N_1805,N_1754,N_1759);
or U1806 (N_1806,N_1763,N_1756);
and U1807 (N_1807,N_1766,N_1768);
nand U1808 (N_1808,N_1773,N_1739);
nand U1809 (N_1809,N_1779,N_1797);
nor U1810 (N_1810,N_1769,N_1755);
nand U1811 (N_1811,N_1796,N_1741);
or U1812 (N_1812,N_1767,N_1798);
nand U1813 (N_1813,N_1765,N_1745);
and U1814 (N_1814,N_1758,N_1753);
nor U1815 (N_1815,N_1736,N_1788);
nor U1816 (N_1816,N_1780,N_1762);
nand U1817 (N_1817,N_1731,N_1787);
and U1818 (N_1818,N_1750,N_1742);
and U1819 (N_1819,N_1785,N_1737);
xor U1820 (N_1820,N_1751,N_1778);
nor U1821 (N_1821,N_1784,N_1738);
or U1822 (N_1822,N_1729,N_1786);
nor U1823 (N_1823,N_1794,N_1747);
and U1824 (N_1824,N_1733,N_1764);
nand U1825 (N_1825,N_1749,N_1776);
xor U1826 (N_1826,N_1757,N_1791);
nor U1827 (N_1827,N_1782,N_1740);
nor U1828 (N_1828,N_1746,N_1748);
and U1829 (N_1829,N_1789,N_1735);
nor U1830 (N_1830,N_1730,N_1772);
and U1831 (N_1831,N_1744,N_1743);
nand U1832 (N_1832,N_1734,N_1728);
or U1833 (N_1833,N_1781,N_1799);
nand U1834 (N_1834,N_1774,N_1732);
nand U1835 (N_1835,N_1725,N_1790);
and U1836 (N_1836,N_1771,N_1760);
nor U1837 (N_1837,N_1770,N_1753);
and U1838 (N_1838,N_1734,N_1776);
and U1839 (N_1839,N_1732,N_1755);
nor U1840 (N_1840,N_1746,N_1758);
nor U1841 (N_1841,N_1740,N_1771);
nor U1842 (N_1842,N_1781,N_1756);
and U1843 (N_1843,N_1765,N_1783);
nand U1844 (N_1844,N_1742,N_1744);
or U1845 (N_1845,N_1751,N_1795);
and U1846 (N_1846,N_1761,N_1785);
nor U1847 (N_1847,N_1736,N_1763);
or U1848 (N_1848,N_1776,N_1726);
and U1849 (N_1849,N_1797,N_1759);
or U1850 (N_1850,N_1769,N_1736);
and U1851 (N_1851,N_1785,N_1730);
nand U1852 (N_1852,N_1765,N_1755);
nand U1853 (N_1853,N_1740,N_1739);
or U1854 (N_1854,N_1764,N_1730);
nor U1855 (N_1855,N_1743,N_1771);
and U1856 (N_1856,N_1799,N_1794);
nand U1857 (N_1857,N_1733,N_1753);
nand U1858 (N_1858,N_1790,N_1743);
or U1859 (N_1859,N_1775,N_1731);
and U1860 (N_1860,N_1786,N_1757);
nand U1861 (N_1861,N_1797,N_1785);
or U1862 (N_1862,N_1786,N_1775);
nor U1863 (N_1863,N_1734,N_1742);
xor U1864 (N_1864,N_1785,N_1751);
nor U1865 (N_1865,N_1765,N_1751);
and U1866 (N_1866,N_1796,N_1797);
nor U1867 (N_1867,N_1774,N_1771);
nand U1868 (N_1868,N_1738,N_1765);
nor U1869 (N_1869,N_1769,N_1775);
nor U1870 (N_1870,N_1734,N_1788);
nand U1871 (N_1871,N_1765,N_1733);
nor U1872 (N_1872,N_1747,N_1771);
or U1873 (N_1873,N_1732,N_1782);
xnor U1874 (N_1874,N_1769,N_1772);
or U1875 (N_1875,N_1869,N_1858);
and U1876 (N_1876,N_1811,N_1828);
nor U1877 (N_1877,N_1842,N_1856);
and U1878 (N_1878,N_1848,N_1865);
nand U1879 (N_1879,N_1800,N_1806);
nor U1880 (N_1880,N_1833,N_1810);
nor U1881 (N_1881,N_1863,N_1812);
nand U1882 (N_1882,N_1830,N_1866);
nor U1883 (N_1883,N_1809,N_1831);
and U1884 (N_1884,N_1836,N_1844);
or U1885 (N_1885,N_1843,N_1813);
nand U1886 (N_1886,N_1807,N_1814);
nand U1887 (N_1887,N_1846,N_1847);
and U1888 (N_1888,N_1839,N_1864);
nor U1889 (N_1889,N_1822,N_1835);
and U1890 (N_1890,N_1829,N_1816);
or U1891 (N_1891,N_1818,N_1853);
nand U1892 (N_1892,N_1852,N_1862);
nor U1893 (N_1893,N_1801,N_1855);
nor U1894 (N_1894,N_1802,N_1815);
and U1895 (N_1895,N_1803,N_1808);
or U1896 (N_1896,N_1851,N_1817);
or U1897 (N_1897,N_1823,N_1873);
nand U1898 (N_1898,N_1838,N_1832);
or U1899 (N_1899,N_1854,N_1870);
and U1900 (N_1900,N_1819,N_1867);
nand U1901 (N_1901,N_1861,N_1824);
or U1902 (N_1902,N_1849,N_1868);
and U1903 (N_1903,N_1872,N_1821);
nand U1904 (N_1904,N_1841,N_1860);
nor U1905 (N_1905,N_1805,N_1820);
nand U1906 (N_1906,N_1845,N_1826);
xnor U1907 (N_1907,N_1840,N_1834);
nor U1908 (N_1908,N_1857,N_1825);
and U1909 (N_1909,N_1837,N_1850);
nand U1910 (N_1910,N_1874,N_1827);
nand U1911 (N_1911,N_1804,N_1871);
nor U1912 (N_1912,N_1859,N_1807);
and U1913 (N_1913,N_1825,N_1824);
nand U1914 (N_1914,N_1854,N_1847);
and U1915 (N_1915,N_1847,N_1858);
xor U1916 (N_1916,N_1863,N_1811);
and U1917 (N_1917,N_1836,N_1857);
and U1918 (N_1918,N_1828,N_1814);
and U1919 (N_1919,N_1836,N_1872);
nor U1920 (N_1920,N_1835,N_1843);
nor U1921 (N_1921,N_1842,N_1840);
or U1922 (N_1922,N_1873,N_1868);
and U1923 (N_1923,N_1856,N_1836);
or U1924 (N_1924,N_1867,N_1817);
and U1925 (N_1925,N_1815,N_1803);
or U1926 (N_1926,N_1861,N_1847);
nor U1927 (N_1927,N_1822,N_1818);
or U1928 (N_1928,N_1847,N_1874);
nor U1929 (N_1929,N_1807,N_1819);
or U1930 (N_1930,N_1849,N_1821);
nor U1931 (N_1931,N_1850,N_1821);
or U1932 (N_1932,N_1863,N_1843);
nand U1933 (N_1933,N_1853,N_1825);
xnor U1934 (N_1934,N_1846,N_1801);
nor U1935 (N_1935,N_1868,N_1816);
and U1936 (N_1936,N_1800,N_1822);
nand U1937 (N_1937,N_1826,N_1865);
and U1938 (N_1938,N_1812,N_1873);
and U1939 (N_1939,N_1842,N_1862);
or U1940 (N_1940,N_1825,N_1846);
xnor U1941 (N_1941,N_1836,N_1833);
or U1942 (N_1942,N_1812,N_1826);
nand U1943 (N_1943,N_1848,N_1818);
or U1944 (N_1944,N_1818,N_1854);
nand U1945 (N_1945,N_1835,N_1874);
or U1946 (N_1946,N_1800,N_1818);
and U1947 (N_1947,N_1851,N_1805);
nand U1948 (N_1948,N_1818,N_1836);
nand U1949 (N_1949,N_1843,N_1873);
nand U1950 (N_1950,N_1899,N_1911);
nand U1951 (N_1951,N_1924,N_1931);
nor U1952 (N_1952,N_1879,N_1878);
nand U1953 (N_1953,N_1944,N_1929);
nor U1954 (N_1954,N_1937,N_1908);
nor U1955 (N_1955,N_1925,N_1886);
or U1956 (N_1956,N_1928,N_1885);
nand U1957 (N_1957,N_1915,N_1912);
or U1958 (N_1958,N_1946,N_1910);
nor U1959 (N_1959,N_1895,N_1906);
or U1960 (N_1960,N_1893,N_1947);
and U1961 (N_1961,N_1898,N_1940);
xnor U1962 (N_1962,N_1941,N_1881);
nor U1963 (N_1963,N_1923,N_1875);
nor U1964 (N_1964,N_1914,N_1884);
or U1965 (N_1965,N_1945,N_1936);
and U1966 (N_1966,N_1942,N_1943);
or U1967 (N_1967,N_1896,N_1891);
and U1968 (N_1968,N_1883,N_1921);
nand U1969 (N_1969,N_1932,N_1935);
nor U1970 (N_1970,N_1894,N_1949);
nor U1971 (N_1971,N_1922,N_1927);
nand U1972 (N_1972,N_1938,N_1917);
or U1973 (N_1973,N_1948,N_1926);
and U1974 (N_1974,N_1905,N_1890);
xor U1975 (N_1975,N_1877,N_1916);
nand U1976 (N_1976,N_1913,N_1887);
nand U1977 (N_1977,N_1882,N_1880);
nor U1978 (N_1978,N_1901,N_1933);
or U1979 (N_1979,N_1889,N_1902);
xor U1980 (N_1980,N_1876,N_1907);
nand U1981 (N_1981,N_1918,N_1888);
nor U1982 (N_1982,N_1904,N_1903);
or U1983 (N_1983,N_1897,N_1909);
and U1984 (N_1984,N_1900,N_1934);
xor U1985 (N_1985,N_1930,N_1920);
and U1986 (N_1986,N_1892,N_1919);
or U1987 (N_1987,N_1939,N_1893);
nor U1988 (N_1988,N_1905,N_1923);
xnor U1989 (N_1989,N_1876,N_1945);
and U1990 (N_1990,N_1901,N_1899);
or U1991 (N_1991,N_1876,N_1926);
nand U1992 (N_1992,N_1884,N_1934);
nand U1993 (N_1993,N_1914,N_1924);
or U1994 (N_1994,N_1913,N_1945);
and U1995 (N_1995,N_1877,N_1900);
or U1996 (N_1996,N_1913,N_1875);
nor U1997 (N_1997,N_1917,N_1943);
nor U1998 (N_1998,N_1901,N_1942);
nor U1999 (N_1999,N_1876,N_1941);
xor U2000 (N_2000,N_1907,N_1940);
nor U2001 (N_2001,N_1880,N_1915);
and U2002 (N_2002,N_1914,N_1921);
nand U2003 (N_2003,N_1894,N_1895);
nor U2004 (N_2004,N_1939,N_1923);
or U2005 (N_2005,N_1900,N_1917);
and U2006 (N_2006,N_1921,N_1916);
and U2007 (N_2007,N_1937,N_1930);
or U2008 (N_2008,N_1913,N_1896);
and U2009 (N_2009,N_1939,N_1901);
or U2010 (N_2010,N_1928,N_1948);
and U2011 (N_2011,N_1930,N_1902);
nor U2012 (N_2012,N_1903,N_1938);
and U2013 (N_2013,N_1880,N_1944);
or U2014 (N_2014,N_1921,N_1902);
nand U2015 (N_2015,N_1909,N_1919);
nor U2016 (N_2016,N_1941,N_1935);
nand U2017 (N_2017,N_1904,N_1875);
nand U2018 (N_2018,N_1935,N_1947);
and U2019 (N_2019,N_1928,N_1921);
nand U2020 (N_2020,N_1892,N_1893);
nand U2021 (N_2021,N_1903,N_1925);
or U2022 (N_2022,N_1890,N_1941);
nand U2023 (N_2023,N_1919,N_1877);
nand U2024 (N_2024,N_1930,N_1929);
nor U2025 (N_2025,N_2016,N_1974);
nand U2026 (N_2026,N_2013,N_2022);
nand U2027 (N_2027,N_1966,N_2011);
or U2028 (N_2028,N_1985,N_1986);
and U2029 (N_2029,N_1968,N_2020);
nand U2030 (N_2030,N_1980,N_1999);
and U2031 (N_2031,N_1958,N_1953);
and U2032 (N_2032,N_2017,N_1975);
nand U2033 (N_2033,N_1990,N_2018);
or U2034 (N_2034,N_2008,N_1962);
and U2035 (N_2035,N_1998,N_2001);
nor U2036 (N_2036,N_1981,N_1954);
and U2037 (N_2037,N_2015,N_1959);
and U2038 (N_2038,N_1950,N_1952);
xor U2039 (N_2039,N_1960,N_2005);
or U2040 (N_2040,N_1967,N_1991);
nor U2041 (N_2041,N_2006,N_2012);
or U2042 (N_2042,N_1971,N_2019);
and U2043 (N_2043,N_1973,N_2007);
nor U2044 (N_2044,N_1988,N_2021);
and U2045 (N_2045,N_2023,N_1951);
and U2046 (N_2046,N_1977,N_2024);
or U2047 (N_2047,N_1992,N_2000);
nand U2048 (N_2048,N_1961,N_1978);
or U2049 (N_2049,N_2003,N_1969);
nor U2050 (N_2050,N_1965,N_2014);
nand U2051 (N_2051,N_1997,N_2002);
and U2052 (N_2052,N_2010,N_1982);
or U2053 (N_2053,N_1972,N_1989);
nor U2054 (N_2054,N_1963,N_1964);
and U2055 (N_2055,N_1993,N_1984);
nor U2056 (N_2056,N_1995,N_1956);
nand U2057 (N_2057,N_1957,N_1979);
nor U2058 (N_2058,N_1970,N_1994);
or U2059 (N_2059,N_2009,N_1976);
or U2060 (N_2060,N_2004,N_1987);
nor U2061 (N_2061,N_1996,N_1983);
and U2062 (N_2062,N_1955,N_1951);
nand U2063 (N_2063,N_1969,N_1962);
nor U2064 (N_2064,N_1983,N_2019);
nand U2065 (N_2065,N_1989,N_1957);
nand U2066 (N_2066,N_1957,N_1956);
or U2067 (N_2067,N_1978,N_1997);
and U2068 (N_2068,N_1967,N_2021);
and U2069 (N_2069,N_1963,N_1974);
or U2070 (N_2070,N_2011,N_1956);
and U2071 (N_2071,N_1975,N_2004);
nand U2072 (N_2072,N_2006,N_1991);
nand U2073 (N_2073,N_1978,N_2010);
or U2074 (N_2074,N_2006,N_1977);
and U2075 (N_2075,N_2000,N_1983);
and U2076 (N_2076,N_2021,N_1970);
or U2077 (N_2077,N_2014,N_1988);
nor U2078 (N_2078,N_1990,N_2005);
nand U2079 (N_2079,N_2023,N_1980);
nor U2080 (N_2080,N_1957,N_2021);
nand U2081 (N_2081,N_1976,N_1993);
or U2082 (N_2082,N_2016,N_1983);
nand U2083 (N_2083,N_2014,N_1961);
and U2084 (N_2084,N_2004,N_1991);
or U2085 (N_2085,N_1990,N_2016);
nor U2086 (N_2086,N_1958,N_1954);
nand U2087 (N_2087,N_1976,N_1992);
or U2088 (N_2088,N_2013,N_1965);
nand U2089 (N_2089,N_2019,N_1991);
and U2090 (N_2090,N_1963,N_1961);
or U2091 (N_2091,N_1984,N_2019);
nand U2092 (N_2092,N_1952,N_1974);
or U2093 (N_2093,N_1953,N_1967);
nand U2094 (N_2094,N_1957,N_1958);
and U2095 (N_2095,N_1987,N_1986);
nor U2096 (N_2096,N_1962,N_1973);
nor U2097 (N_2097,N_1966,N_2008);
and U2098 (N_2098,N_1971,N_2009);
nand U2099 (N_2099,N_1986,N_1966);
nand U2100 (N_2100,N_2034,N_2039);
nand U2101 (N_2101,N_2061,N_2095);
or U2102 (N_2102,N_2045,N_2062);
and U2103 (N_2103,N_2099,N_2040);
and U2104 (N_2104,N_2051,N_2079);
and U2105 (N_2105,N_2028,N_2078);
nor U2106 (N_2106,N_2090,N_2033);
and U2107 (N_2107,N_2031,N_2067);
or U2108 (N_2108,N_2037,N_2074);
and U2109 (N_2109,N_2057,N_2089);
or U2110 (N_2110,N_2064,N_2027);
or U2111 (N_2111,N_2093,N_2068);
or U2112 (N_2112,N_2055,N_2035);
and U2113 (N_2113,N_2050,N_2056);
or U2114 (N_2114,N_2094,N_2059);
or U2115 (N_2115,N_2081,N_2065);
nor U2116 (N_2116,N_2046,N_2098);
or U2117 (N_2117,N_2075,N_2087);
and U2118 (N_2118,N_2092,N_2077);
and U2119 (N_2119,N_2026,N_2080);
nand U2120 (N_2120,N_2030,N_2041);
and U2121 (N_2121,N_2083,N_2047);
nor U2122 (N_2122,N_2060,N_2032);
or U2123 (N_2123,N_2052,N_2085);
and U2124 (N_2124,N_2063,N_2088);
nand U2125 (N_2125,N_2082,N_2069);
nand U2126 (N_2126,N_2029,N_2025);
nand U2127 (N_2127,N_2070,N_2048);
nand U2128 (N_2128,N_2053,N_2072);
or U2129 (N_2129,N_2091,N_2044);
or U2130 (N_2130,N_2076,N_2038);
and U2131 (N_2131,N_2043,N_2071);
nand U2132 (N_2132,N_2073,N_2058);
or U2133 (N_2133,N_2084,N_2049);
and U2134 (N_2134,N_2054,N_2096);
nand U2135 (N_2135,N_2097,N_2036);
or U2136 (N_2136,N_2042,N_2086);
or U2137 (N_2137,N_2066,N_2058);
nor U2138 (N_2138,N_2055,N_2074);
nor U2139 (N_2139,N_2085,N_2094);
nor U2140 (N_2140,N_2025,N_2049);
nand U2141 (N_2141,N_2041,N_2066);
or U2142 (N_2142,N_2035,N_2086);
or U2143 (N_2143,N_2073,N_2099);
and U2144 (N_2144,N_2052,N_2029);
and U2145 (N_2145,N_2087,N_2053);
nand U2146 (N_2146,N_2073,N_2094);
nor U2147 (N_2147,N_2081,N_2058);
nor U2148 (N_2148,N_2086,N_2039);
nand U2149 (N_2149,N_2048,N_2072);
nand U2150 (N_2150,N_2034,N_2086);
nor U2151 (N_2151,N_2052,N_2086);
or U2152 (N_2152,N_2041,N_2065);
nand U2153 (N_2153,N_2079,N_2072);
and U2154 (N_2154,N_2039,N_2070);
and U2155 (N_2155,N_2091,N_2060);
or U2156 (N_2156,N_2091,N_2063);
nand U2157 (N_2157,N_2052,N_2047);
nor U2158 (N_2158,N_2046,N_2076);
nand U2159 (N_2159,N_2060,N_2049);
or U2160 (N_2160,N_2031,N_2095);
or U2161 (N_2161,N_2093,N_2063);
or U2162 (N_2162,N_2040,N_2042);
nor U2163 (N_2163,N_2060,N_2025);
and U2164 (N_2164,N_2077,N_2093);
nand U2165 (N_2165,N_2046,N_2062);
or U2166 (N_2166,N_2057,N_2064);
or U2167 (N_2167,N_2052,N_2044);
or U2168 (N_2168,N_2028,N_2072);
nand U2169 (N_2169,N_2040,N_2057);
and U2170 (N_2170,N_2090,N_2044);
or U2171 (N_2171,N_2027,N_2041);
and U2172 (N_2172,N_2054,N_2070);
and U2173 (N_2173,N_2083,N_2051);
or U2174 (N_2174,N_2083,N_2062);
nand U2175 (N_2175,N_2126,N_2136);
or U2176 (N_2176,N_2132,N_2160);
nor U2177 (N_2177,N_2137,N_2114);
nor U2178 (N_2178,N_2139,N_2104);
and U2179 (N_2179,N_2169,N_2105);
nor U2180 (N_2180,N_2148,N_2128);
or U2181 (N_2181,N_2101,N_2144);
nor U2182 (N_2182,N_2173,N_2110);
nor U2183 (N_2183,N_2133,N_2174);
or U2184 (N_2184,N_2131,N_2166);
nand U2185 (N_2185,N_2167,N_2122);
nand U2186 (N_2186,N_2141,N_2117);
nand U2187 (N_2187,N_2162,N_2172);
and U2188 (N_2188,N_2112,N_2147);
or U2189 (N_2189,N_2140,N_2130);
nand U2190 (N_2190,N_2124,N_2164);
or U2191 (N_2191,N_2157,N_2150);
and U2192 (N_2192,N_2106,N_2111);
nor U2193 (N_2193,N_2100,N_2155);
nand U2194 (N_2194,N_2121,N_2171);
and U2195 (N_2195,N_2123,N_2107);
nand U2196 (N_2196,N_2127,N_2153);
and U2197 (N_2197,N_2135,N_2103);
nor U2198 (N_2198,N_2142,N_2145);
or U2199 (N_2199,N_2168,N_2151);
nor U2200 (N_2200,N_2146,N_2158);
or U2201 (N_2201,N_2118,N_2109);
and U2202 (N_2202,N_2154,N_2165);
and U2203 (N_2203,N_2113,N_2134);
nand U2204 (N_2204,N_2138,N_2120);
nor U2205 (N_2205,N_2102,N_2129);
and U2206 (N_2206,N_2159,N_2152);
or U2207 (N_2207,N_2143,N_2170);
nor U2208 (N_2208,N_2125,N_2156);
nor U2209 (N_2209,N_2115,N_2163);
nor U2210 (N_2210,N_2108,N_2119);
nor U2211 (N_2211,N_2116,N_2161);
and U2212 (N_2212,N_2149,N_2123);
xor U2213 (N_2213,N_2153,N_2150);
nor U2214 (N_2214,N_2171,N_2158);
and U2215 (N_2215,N_2128,N_2136);
nor U2216 (N_2216,N_2122,N_2157);
or U2217 (N_2217,N_2174,N_2146);
xnor U2218 (N_2218,N_2111,N_2159);
or U2219 (N_2219,N_2111,N_2171);
or U2220 (N_2220,N_2138,N_2125);
nand U2221 (N_2221,N_2164,N_2152);
and U2222 (N_2222,N_2139,N_2118);
or U2223 (N_2223,N_2174,N_2106);
or U2224 (N_2224,N_2127,N_2140);
and U2225 (N_2225,N_2139,N_2173);
nor U2226 (N_2226,N_2139,N_2150);
nand U2227 (N_2227,N_2159,N_2156);
and U2228 (N_2228,N_2141,N_2165);
or U2229 (N_2229,N_2150,N_2126);
xnor U2230 (N_2230,N_2154,N_2150);
and U2231 (N_2231,N_2104,N_2152);
nor U2232 (N_2232,N_2169,N_2127);
or U2233 (N_2233,N_2129,N_2115);
and U2234 (N_2234,N_2127,N_2135);
nor U2235 (N_2235,N_2128,N_2165);
or U2236 (N_2236,N_2156,N_2149);
nand U2237 (N_2237,N_2174,N_2111);
nand U2238 (N_2238,N_2108,N_2148);
and U2239 (N_2239,N_2130,N_2160);
and U2240 (N_2240,N_2173,N_2141);
xor U2241 (N_2241,N_2142,N_2117);
or U2242 (N_2242,N_2106,N_2164);
nor U2243 (N_2243,N_2108,N_2174);
or U2244 (N_2244,N_2131,N_2152);
and U2245 (N_2245,N_2114,N_2117);
nand U2246 (N_2246,N_2162,N_2157);
or U2247 (N_2247,N_2137,N_2155);
nand U2248 (N_2248,N_2166,N_2114);
and U2249 (N_2249,N_2136,N_2110);
or U2250 (N_2250,N_2232,N_2234);
nor U2251 (N_2251,N_2189,N_2243);
nor U2252 (N_2252,N_2240,N_2213);
nor U2253 (N_2253,N_2238,N_2228);
xnor U2254 (N_2254,N_2193,N_2236);
nand U2255 (N_2255,N_2239,N_2184);
nand U2256 (N_2256,N_2186,N_2199);
nand U2257 (N_2257,N_2177,N_2245);
and U2258 (N_2258,N_2179,N_2202);
nand U2259 (N_2259,N_2246,N_2201);
and U2260 (N_2260,N_2235,N_2211);
or U2261 (N_2261,N_2200,N_2203);
and U2262 (N_2262,N_2181,N_2204);
nor U2263 (N_2263,N_2225,N_2230);
and U2264 (N_2264,N_2242,N_2194);
nand U2265 (N_2265,N_2206,N_2198);
nor U2266 (N_2266,N_2229,N_2247);
nor U2267 (N_2267,N_2188,N_2209);
nand U2268 (N_2268,N_2185,N_2233);
nand U2269 (N_2269,N_2210,N_2248);
xnor U2270 (N_2270,N_2218,N_2208);
nand U2271 (N_2271,N_2217,N_2220);
and U2272 (N_2272,N_2226,N_2231);
xor U2273 (N_2273,N_2222,N_2215);
nor U2274 (N_2274,N_2187,N_2195);
nand U2275 (N_2275,N_2244,N_2176);
xor U2276 (N_2276,N_2227,N_2214);
and U2277 (N_2277,N_2196,N_2207);
nand U2278 (N_2278,N_2175,N_2223);
nor U2279 (N_2279,N_2205,N_2212);
nor U2280 (N_2280,N_2180,N_2192);
nand U2281 (N_2281,N_2178,N_2221);
nor U2282 (N_2282,N_2216,N_2191);
nor U2283 (N_2283,N_2197,N_2224);
nand U2284 (N_2284,N_2249,N_2183);
nand U2285 (N_2285,N_2237,N_2219);
or U2286 (N_2286,N_2182,N_2241);
and U2287 (N_2287,N_2190,N_2241);
and U2288 (N_2288,N_2185,N_2243);
or U2289 (N_2289,N_2197,N_2194);
nor U2290 (N_2290,N_2236,N_2227);
nand U2291 (N_2291,N_2198,N_2177);
or U2292 (N_2292,N_2236,N_2244);
xor U2293 (N_2293,N_2214,N_2212);
nand U2294 (N_2294,N_2230,N_2246);
or U2295 (N_2295,N_2233,N_2235);
or U2296 (N_2296,N_2209,N_2198);
or U2297 (N_2297,N_2200,N_2196);
nand U2298 (N_2298,N_2228,N_2231);
nand U2299 (N_2299,N_2219,N_2195);
nand U2300 (N_2300,N_2182,N_2236);
and U2301 (N_2301,N_2176,N_2228);
nand U2302 (N_2302,N_2207,N_2191);
and U2303 (N_2303,N_2194,N_2240);
nand U2304 (N_2304,N_2183,N_2209);
or U2305 (N_2305,N_2210,N_2207);
nor U2306 (N_2306,N_2228,N_2213);
nand U2307 (N_2307,N_2185,N_2198);
nand U2308 (N_2308,N_2182,N_2178);
and U2309 (N_2309,N_2183,N_2218);
nor U2310 (N_2310,N_2223,N_2219);
nand U2311 (N_2311,N_2180,N_2219);
or U2312 (N_2312,N_2214,N_2229);
or U2313 (N_2313,N_2197,N_2177);
nand U2314 (N_2314,N_2234,N_2194);
nand U2315 (N_2315,N_2217,N_2192);
nand U2316 (N_2316,N_2205,N_2203);
and U2317 (N_2317,N_2211,N_2214);
or U2318 (N_2318,N_2247,N_2201);
xnor U2319 (N_2319,N_2179,N_2194);
nand U2320 (N_2320,N_2186,N_2209);
nor U2321 (N_2321,N_2225,N_2191);
xnor U2322 (N_2322,N_2186,N_2192);
and U2323 (N_2323,N_2245,N_2203);
and U2324 (N_2324,N_2230,N_2177);
nand U2325 (N_2325,N_2255,N_2260);
nand U2326 (N_2326,N_2322,N_2293);
or U2327 (N_2327,N_2299,N_2267);
or U2328 (N_2328,N_2253,N_2315);
nand U2329 (N_2329,N_2309,N_2281);
and U2330 (N_2330,N_2282,N_2317);
nor U2331 (N_2331,N_2308,N_2270);
and U2332 (N_2332,N_2291,N_2321);
and U2333 (N_2333,N_2261,N_2287);
or U2334 (N_2334,N_2285,N_2278);
nand U2335 (N_2335,N_2264,N_2320);
or U2336 (N_2336,N_2279,N_2314);
and U2337 (N_2337,N_2306,N_2259);
and U2338 (N_2338,N_2250,N_2272);
nor U2339 (N_2339,N_2316,N_2286);
and U2340 (N_2340,N_2280,N_2273);
nor U2341 (N_2341,N_2265,N_2269);
nor U2342 (N_2342,N_2294,N_2266);
and U2343 (N_2343,N_2258,N_2263);
or U2344 (N_2344,N_2283,N_2284);
or U2345 (N_2345,N_2311,N_2303);
or U2346 (N_2346,N_2289,N_2288);
nor U2347 (N_2347,N_2310,N_2262);
and U2348 (N_2348,N_2256,N_2300);
and U2349 (N_2349,N_2274,N_2323);
nor U2350 (N_2350,N_2301,N_2277);
nor U2351 (N_2351,N_2276,N_2307);
or U2352 (N_2352,N_2312,N_2318);
or U2353 (N_2353,N_2324,N_2275);
nand U2354 (N_2354,N_2268,N_2292);
nor U2355 (N_2355,N_2305,N_2271);
xnor U2356 (N_2356,N_2298,N_2304);
and U2357 (N_2357,N_2295,N_2302);
and U2358 (N_2358,N_2319,N_2290);
nor U2359 (N_2359,N_2251,N_2313);
nor U2360 (N_2360,N_2257,N_2296);
xor U2361 (N_2361,N_2254,N_2252);
nor U2362 (N_2362,N_2297,N_2310);
xor U2363 (N_2363,N_2282,N_2310);
nor U2364 (N_2364,N_2317,N_2269);
nand U2365 (N_2365,N_2321,N_2257);
nor U2366 (N_2366,N_2267,N_2270);
nor U2367 (N_2367,N_2322,N_2295);
nor U2368 (N_2368,N_2319,N_2282);
or U2369 (N_2369,N_2276,N_2313);
nor U2370 (N_2370,N_2279,N_2315);
nor U2371 (N_2371,N_2296,N_2319);
nand U2372 (N_2372,N_2311,N_2310);
nor U2373 (N_2373,N_2297,N_2315);
nor U2374 (N_2374,N_2266,N_2279);
nor U2375 (N_2375,N_2277,N_2263);
nand U2376 (N_2376,N_2255,N_2304);
nor U2377 (N_2377,N_2263,N_2296);
xor U2378 (N_2378,N_2268,N_2265);
or U2379 (N_2379,N_2258,N_2262);
or U2380 (N_2380,N_2299,N_2296);
xnor U2381 (N_2381,N_2262,N_2251);
or U2382 (N_2382,N_2250,N_2269);
nor U2383 (N_2383,N_2264,N_2322);
and U2384 (N_2384,N_2304,N_2266);
nor U2385 (N_2385,N_2285,N_2288);
nor U2386 (N_2386,N_2251,N_2299);
nand U2387 (N_2387,N_2302,N_2275);
or U2388 (N_2388,N_2279,N_2251);
or U2389 (N_2389,N_2309,N_2290);
nand U2390 (N_2390,N_2297,N_2260);
nor U2391 (N_2391,N_2307,N_2274);
nor U2392 (N_2392,N_2319,N_2318);
nand U2393 (N_2393,N_2266,N_2261);
or U2394 (N_2394,N_2307,N_2267);
and U2395 (N_2395,N_2266,N_2317);
or U2396 (N_2396,N_2313,N_2264);
and U2397 (N_2397,N_2252,N_2301);
or U2398 (N_2398,N_2260,N_2319);
nor U2399 (N_2399,N_2323,N_2292);
nor U2400 (N_2400,N_2351,N_2339);
nand U2401 (N_2401,N_2370,N_2329);
and U2402 (N_2402,N_2385,N_2380);
nand U2403 (N_2403,N_2393,N_2356);
and U2404 (N_2404,N_2359,N_2382);
nand U2405 (N_2405,N_2394,N_2381);
or U2406 (N_2406,N_2379,N_2372);
and U2407 (N_2407,N_2357,N_2353);
nand U2408 (N_2408,N_2389,N_2378);
nor U2409 (N_2409,N_2388,N_2331);
and U2410 (N_2410,N_2342,N_2396);
nand U2411 (N_2411,N_2361,N_2364);
xor U2412 (N_2412,N_2337,N_2358);
and U2413 (N_2413,N_2366,N_2328);
nand U2414 (N_2414,N_2365,N_2330);
nand U2415 (N_2415,N_2354,N_2325);
nor U2416 (N_2416,N_2377,N_2369);
nor U2417 (N_2417,N_2368,N_2363);
nand U2418 (N_2418,N_2336,N_2348);
nand U2419 (N_2419,N_2360,N_2327);
or U2420 (N_2420,N_2375,N_2373);
nor U2421 (N_2421,N_2343,N_2390);
or U2422 (N_2422,N_2335,N_2341);
or U2423 (N_2423,N_2345,N_2367);
or U2424 (N_2424,N_2332,N_2386);
and U2425 (N_2425,N_2384,N_2355);
nor U2426 (N_2426,N_2383,N_2340);
or U2427 (N_2427,N_2376,N_2338);
nor U2428 (N_2428,N_2350,N_2344);
or U2429 (N_2429,N_2362,N_2352);
and U2430 (N_2430,N_2387,N_2347);
nor U2431 (N_2431,N_2391,N_2374);
or U2432 (N_2432,N_2399,N_2397);
and U2433 (N_2433,N_2395,N_2346);
nor U2434 (N_2434,N_2326,N_2334);
nand U2435 (N_2435,N_2371,N_2333);
nand U2436 (N_2436,N_2349,N_2398);
nand U2437 (N_2437,N_2392,N_2336);
and U2438 (N_2438,N_2334,N_2345);
nand U2439 (N_2439,N_2398,N_2355);
and U2440 (N_2440,N_2380,N_2351);
nand U2441 (N_2441,N_2393,N_2351);
and U2442 (N_2442,N_2325,N_2344);
and U2443 (N_2443,N_2341,N_2382);
or U2444 (N_2444,N_2363,N_2360);
nor U2445 (N_2445,N_2343,N_2329);
and U2446 (N_2446,N_2385,N_2338);
nor U2447 (N_2447,N_2395,N_2377);
or U2448 (N_2448,N_2394,N_2374);
or U2449 (N_2449,N_2399,N_2372);
or U2450 (N_2450,N_2391,N_2356);
or U2451 (N_2451,N_2388,N_2379);
or U2452 (N_2452,N_2325,N_2369);
nand U2453 (N_2453,N_2330,N_2379);
nand U2454 (N_2454,N_2329,N_2385);
or U2455 (N_2455,N_2386,N_2346);
and U2456 (N_2456,N_2389,N_2386);
or U2457 (N_2457,N_2330,N_2395);
or U2458 (N_2458,N_2337,N_2381);
xnor U2459 (N_2459,N_2344,N_2381);
and U2460 (N_2460,N_2362,N_2364);
nand U2461 (N_2461,N_2377,N_2373);
and U2462 (N_2462,N_2395,N_2371);
nand U2463 (N_2463,N_2371,N_2392);
and U2464 (N_2464,N_2384,N_2354);
and U2465 (N_2465,N_2367,N_2362);
xor U2466 (N_2466,N_2365,N_2342);
xnor U2467 (N_2467,N_2378,N_2375);
nand U2468 (N_2468,N_2364,N_2383);
xnor U2469 (N_2469,N_2381,N_2339);
or U2470 (N_2470,N_2330,N_2329);
and U2471 (N_2471,N_2372,N_2362);
nor U2472 (N_2472,N_2395,N_2393);
and U2473 (N_2473,N_2338,N_2331);
and U2474 (N_2474,N_2338,N_2383);
xor U2475 (N_2475,N_2465,N_2430);
xnor U2476 (N_2476,N_2453,N_2404);
nor U2477 (N_2477,N_2412,N_2445);
or U2478 (N_2478,N_2459,N_2434);
or U2479 (N_2479,N_2403,N_2426);
and U2480 (N_2480,N_2454,N_2428);
or U2481 (N_2481,N_2448,N_2410);
xor U2482 (N_2482,N_2460,N_2440);
nor U2483 (N_2483,N_2433,N_2463);
and U2484 (N_2484,N_2427,N_2421);
nor U2485 (N_2485,N_2413,N_2467);
nand U2486 (N_2486,N_2456,N_2472);
nand U2487 (N_2487,N_2406,N_2452);
nor U2488 (N_2488,N_2437,N_2446);
or U2489 (N_2489,N_2447,N_2469);
nor U2490 (N_2490,N_2416,N_2400);
or U2491 (N_2491,N_2425,N_2441);
nor U2492 (N_2492,N_2408,N_2466);
and U2493 (N_2493,N_2417,N_2470);
or U2494 (N_2494,N_2415,N_2461);
and U2495 (N_2495,N_2450,N_2401);
and U2496 (N_2496,N_2420,N_2439);
and U2497 (N_2497,N_2402,N_2435);
nand U2498 (N_2498,N_2432,N_2474);
or U2499 (N_2499,N_2449,N_2409);
and U2500 (N_2500,N_2436,N_2443);
nor U2501 (N_2501,N_2438,N_2419);
or U2502 (N_2502,N_2444,N_2464);
and U2503 (N_2503,N_2418,N_2407);
or U2504 (N_2504,N_2473,N_2455);
nor U2505 (N_2505,N_2429,N_2422);
or U2506 (N_2506,N_2442,N_2458);
nand U2507 (N_2507,N_2405,N_2468);
or U2508 (N_2508,N_2471,N_2462);
or U2509 (N_2509,N_2431,N_2424);
nor U2510 (N_2510,N_2457,N_2414);
and U2511 (N_2511,N_2451,N_2411);
and U2512 (N_2512,N_2423,N_2429);
or U2513 (N_2513,N_2427,N_2400);
nor U2514 (N_2514,N_2458,N_2445);
nand U2515 (N_2515,N_2401,N_2465);
nand U2516 (N_2516,N_2408,N_2412);
nand U2517 (N_2517,N_2402,N_2430);
or U2518 (N_2518,N_2445,N_2429);
or U2519 (N_2519,N_2439,N_2419);
nand U2520 (N_2520,N_2438,N_2406);
nand U2521 (N_2521,N_2403,N_2449);
or U2522 (N_2522,N_2419,N_2441);
and U2523 (N_2523,N_2418,N_2434);
nor U2524 (N_2524,N_2438,N_2439);
nand U2525 (N_2525,N_2428,N_2417);
nand U2526 (N_2526,N_2434,N_2437);
nand U2527 (N_2527,N_2459,N_2414);
xnor U2528 (N_2528,N_2420,N_2429);
or U2529 (N_2529,N_2404,N_2461);
nor U2530 (N_2530,N_2449,N_2469);
nor U2531 (N_2531,N_2463,N_2431);
nand U2532 (N_2532,N_2464,N_2408);
or U2533 (N_2533,N_2419,N_2421);
or U2534 (N_2534,N_2412,N_2419);
nand U2535 (N_2535,N_2465,N_2441);
and U2536 (N_2536,N_2433,N_2449);
nand U2537 (N_2537,N_2469,N_2462);
nor U2538 (N_2538,N_2438,N_2408);
xor U2539 (N_2539,N_2413,N_2440);
and U2540 (N_2540,N_2412,N_2430);
and U2541 (N_2541,N_2442,N_2473);
nand U2542 (N_2542,N_2408,N_2416);
or U2543 (N_2543,N_2469,N_2424);
nand U2544 (N_2544,N_2403,N_2460);
or U2545 (N_2545,N_2463,N_2413);
and U2546 (N_2546,N_2457,N_2423);
and U2547 (N_2547,N_2401,N_2453);
xnor U2548 (N_2548,N_2453,N_2438);
nand U2549 (N_2549,N_2463,N_2456);
nor U2550 (N_2550,N_2528,N_2476);
nand U2551 (N_2551,N_2544,N_2542);
and U2552 (N_2552,N_2547,N_2478);
xnor U2553 (N_2553,N_2512,N_2541);
nor U2554 (N_2554,N_2485,N_2515);
and U2555 (N_2555,N_2495,N_2508);
nand U2556 (N_2556,N_2534,N_2537);
or U2557 (N_2557,N_2510,N_2488);
and U2558 (N_2558,N_2536,N_2499);
or U2559 (N_2559,N_2490,N_2525);
or U2560 (N_2560,N_2480,N_2500);
nand U2561 (N_2561,N_2496,N_2477);
and U2562 (N_2562,N_2522,N_2498);
and U2563 (N_2563,N_2501,N_2507);
or U2564 (N_2564,N_2516,N_2513);
or U2565 (N_2565,N_2506,N_2509);
nor U2566 (N_2566,N_2511,N_2484);
nor U2567 (N_2567,N_2491,N_2487);
nand U2568 (N_2568,N_2514,N_2486);
nor U2569 (N_2569,N_2523,N_2531);
nand U2570 (N_2570,N_2504,N_2546);
nor U2571 (N_2571,N_2545,N_2549);
or U2572 (N_2572,N_2540,N_2539);
and U2573 (N_2573,N_2503,N_2521);
nor U2574 (N_2574,N_2526,N_2489);
or U2575 (N_2575,N_2529,N_2492);
and U2576 (N_2576,N_2548,N_2494);
or U2577 (N_2577,N_2538,N_2505);
and U2578 (N_2578,N_2518,N_2520);
nor U2579 (N_2579,N_2533,N_2543);
nor U2580 (N_2580,N_2481,N_2479);
nand U2581 (N_2581,N_2524,N_2493);
or U2582 (N_2582,N_2532,N_2497);
nand U2583 (N_2583,N_2483,N_2502);
nor U2584 (N_2584,N_2535,N_2519);
nor U2585 (N_2585,N_2475,N_2482);
or U2586 (N_2586,N_2530,N_2517);
or U2587 (N_2587,N_2527,N_2531);
nor U2588 (N_2588,N_2488,N_2535);
nor U2589 (N_2589,N_2531,N_2501);
nor U2590 (N_2590,N_2498,N_2476);
or U2591 (N_2591,N_2538,N_2537);
and U2592 (N_2592,N_2478,N_2509);
or U2593 (N_2593,N_2498,N_2519);
nand U2594 (N_2594,N_2497,N_2518);
or U2595 (N_2595,N_2530,N_2516);
and U2596 (N_2596,N_2537,N_2520);
and U2597 (N_2597,N_2504,N_2491);
or U2598 (N_2598,N_2532,N_2527);
nor U2599 (N_2599,N_2506,N_2480);
and U2600 (N_2600,N_2495,N_2522);
and U2601 (N_2601,N_2488,N_2543);
or U2602 (N_2602,N_2481,N_2522);
and U2603 (N_2603,N_2515,N_2524);
or U2604 (N_2604,N_2539,N_2487);
nor U2605 (N_2605,N_2485,N_2536);
or U2606 (N_2606,N_2477,N_2541);
and U2607 (N_2607,N_2530,N_2526);
and U2608 (N_2608,N_2476,N_2536);
and U2609 (N_2609,N_2518,N_2530);
and U2610 (N_2610,N_2510,N_2536);
nor U2611 (N_2611,N_2522,N_2497);
nor U2612 (N_2612,N_2484,N_2525);
or U2613 (N_2613,N_2521,N_2549);
or U2614 (N_2614,N_2504,N_2539);
nand U2615 (N_2615,N_2517,N_2507);
nor U2616 (N_2616,N_2545,N_2541);
or U2617 (N_2617,N_2492,N_2488);
nor U2618 (N_2618,N_2525,N_2546);
nor U2619 (N_2619,N_2545,N_2511);
or U2620 (N_2620,N_2483,N_2485);
nand U2621 (N_2621,N_2535,N_2492);
nor U2622 (N_2622,N_2506,N_2489);
or U2623 (N_2623,N_2506,N_2492);
and U2624 (N_2624,N_2499,N_2505);
and U2625 (N_2625,N_2609,N_2587);
nand U2626 (N_2626,N_2558,N_2556);
and U2627 (N_2627,N_2568,N_2575);
or U2628 (N_2628,N_2617,N_2562);
nor U2629 (N_2629,N_2602,N_2565);
nand U2630 (N_2630,N_2616,N_2576);
nor U2631 (N_2631,N_2560,N_2599);
nor U2632 (N_2632,N_2571,N_2592);
and U2633 (N_2633,N_2583,N_2570);
and U2634 (N_2634,N_2624,N_2574);
and U2635 (N_2635,N_2600,N_2594);
nand U2636 (N_2636,N_2582,N_2577);
or U2637 (N_2637,N_2613,N_2589);
or U2638 (N_2638,N_2607,N_2608);
and U2639 (N_2639,N_2557,N_2623);
or U2640 (N_2640,N_2585,N_2605);
nand U2641 (N_2641,N_2603,N_2578);
nand U2642 (N_2642,N_2566,N_2615);
or U2643 (N_2643,N_2618,N_2590);
nand U2644 (N_2644,N_2606,N_2610);
and U2645 (N_2645,N_2554,N_2550);
nand U2646 (N_2646,N_2569,N_2551);
nor U2647 (N_2647,N_2559,N_2555);
xnor U2648 (N_2648,N_2553,N_2552);
or U2649 (N_2649,N_2595,N_2622);
or U2650 (N_2650,N_2601,N_2580);
or U2651 (N_2651,N_2572,N_2612);
or U2652 (N_2652,N_2564,N_2561);
or U2653 (N_2653,N_2586,N_2593);
and U2654 (N_2654,N_2567,N_2598);
and U2655 (N_2655,N_2604,N_2563);
and U2656 (N_2656,N_2619,N_2579);
nor U2657 (N_2657,N_2596,N_2611);
nand U2658 (N_2658,N_2584,N_2573);
and U2659 (N_2659,N_2581,N_2591);
or U2660 (N_2660,N_2597,N_2620);
or U2661 (N_2661,N_2621,N_2588);
nor U2662 (N_2662,N_2614,N_2559);
and U2663 (N_2663,N_2619,N_2618);
or U2664 (N_2664,N_2571,N_2616);
or U2665 (N_2665,N_2603,N_2616);
or U2666 (N_2666,N_2592,N_2562);
and U2667 (N_2667,N_2594,N_2620);
nand U2668 (N_2668,N_2611,N_2592);
and U2669 (N_2669,N_2574,N_2566);
and U2670 (N_2670,N_2560,N_2592);
or U2671 (N_2671,N_2592,N_2551);
or U2672 (N_2672,N_2566,N_2561);
or U2673 (N_2673,N_2617,N_2564);
nand U2674 (N_2674,N_2588,N_2561);
nand U2675 (N_2675,N_2562,N_2597);
nand U2676 (N_2676,N_2550,N_2589);
nor U2677 (N_2677,N_2587,N_2619);
or U2678 (N_2678,N_2610,N_2605);
nor U2679 (N_2679,N_2558,N_2606);
nor U2680 (N_2680,N_2617,N_2620);
nand U2681 (N_2681,N_2570,N_2590);
and U2682 (N_2682,N_2596,N_2587);
or U2683 (N_2683,N_2598,N_2593);
nor U2684 (N_2684,N_2622,N_2602);
nor U2685 (N_2685,N_2583,N_2601);
nand U2686 (N_2686,N_2610,N_2575);
nor U2687 (N_2687,N_2569,N_2596);
nor U2688 (N_2688,N_2562,N_2624);
nand U2689 (N_2689,N_2585,N_2607);
and U2690 (N_2690,N_2592,N_2584);
or U2691 (N_2691,N_2564,N_2578);
or U2692 (N_2692,N_2555,N_2598);
nand U2693 (N_2693,N_2619,N_2620);
or U2694 (N_2694,N_2556,N_2562);
or U2695 (N_2695,N_2572,N_2607);
and U2696 (N_2696,N_2587,N_2600);
nand U2697 (N_2697,N_2558,N_2596);
nand U2698 (N_2698,N_2571,N_2568);
and U2699 (N_2699,N_2580,N_2572);
nand U2700 (N_2700,N_2637,N_2644);
nand U2701 (N_2701,N_2672,N_2639);
nand U2702 (N_2702,N_2683,N_2675);
nor U2703 (N_2703,N_2665,N_2649);
nor U2704 (N_2704,N_2636,N_2626);
or U2705 (N_2705,N_2692,N_2660);
nand U2706 (N_2706,N_2669,N_2662);
nor U2707 (N_2707,N_2641,N_2635);
nand U2708 (N_2708,N_2699,N_2670);
nand U2709 (N_2709,N_2642,N_2633);
nor U2710 (N_2710,N_2663,N_2659);
and U2711 (N_2711,N_2666,N_2685);
or U2712 (N_2712,N_2679,N_2688);
and U2713 (N_2713,N_2676,N_2627);
and U2714 (N_2714,N_2673,N_2625);
nand U2715 (N_2715,N_2686,N_2678);
nor U2716 (N_2716,N_2650,N_2694);
nand U2717 (N_2717,N_2648,N_2652);
and U2718 (N_2718,N_2645,N_2638);
xor U2719 (N_2719,N_2653,N_2630);
nor U2720 (N_2720,N_2681,N_2646);
nor U2721 (N_2721,N_2680,N_2667);
nor U2722 (N_2722,N_2651,N_2693);
and U2723 (N_2723,N_2643,N_2632);
and U2724 (N_2724,N_2689,N_2664);
nor U2725 (N_2725,N_2684,N_2674);
or U2726 (N_2726,N_2640,N_2687);
or U2727 (N_2727,N_2631,N_2654);
xor U2728 (N_2728,N_2629,N_2657);
nand U2729 (N_2729,N_2668,N_2691);
and U2730 (N_2730,N_2697,N_2634);
or U2731 (N_2731,N_2698,N_2661);
and U2732 (N_2732,N_2695,N_2656);
or U2733 (N_2733,N_2682,N_2655);
nand U2734 (N_2734,N_2647,N_2696);
nor U2735 (N_2735,N_2690,N_2658);
or U2736 (N_2736,N_2677,N_2628);
and U2737 (N_2737,N_2671,N_2674);
nor U2738 (N_2738,N_2643,N_2640);
and U2739 (N_2739,N_2629,N_2655);
or U2740 (N_2740,N_2659,N_2635);
or U2741 (N_2741,N_2679,N_2633);
nand U2742 (N_2742,N_2693,N_2666);
nand U2743 (N_2743,N_2657,N_2627);
xnor U2744 (N_2744,N_2640,N_2683);
or U2745 (N_2745,N_2642,N_2688);
nor U2746 (N_2746,N_2654,N_2666);
nand U2747 (N_2747,N_2677,N_2683);
nor U2748 (N_2748,N_2682,N_2652);
or U2749 (N_2749,N_2655,N_2663);
nand U2750 (N_2750,N_2678,N_2673);
or U2751 (N_2751,N_2665,N_2643);
xnor U2752 (N_2752,N_2654,N_2656);
nor U2753 (N_2753,N_2648,N_2676);
or U2754 (N_2754,N_2668,N_2627);
and U2755 (N_2755,N_2691,N_2643);
nor U2756 (N_2756,N_2629,N_2678);
xnor U2757 (N_2757,N_2631,N_2667);
or U2758 (N_2758,N_2696,N_2677);
nand U2759 (N_2759,N_2674,N_2643);
and U2760 (N_2760,N_2699,N_2676);
and U2761 (N_2761,N_2629,N_2687);
xnor U2762 (N_2762,N_2635,N_2693);
and U2763 (N_2763,N_2635,N_2651);
nor U2764 (N_2764,N_2655,N_2675);
and U2765 (N_2765,N_2654,N_2684);
nor U2766 (N_2766,N_2637,N_2647);
and U2767 (N_2767,N_2671,N_2656);
nor U2768 (N_2768,N_2653,N_2667);
nor U2769 (N_2769,N_2647,N_2635);
and U2770 (N_2770,N_2667,N_2693);
nand U2771 (N_2771,N_2654,N_2696);
nand U2772 (N_2772,N_2692,N_2675);
or U2773 (N_2773,N_2684,N_2659);
or U2774 (N_2774,N_2654,N_2698);
nor U2775 (N_2775,N_2714,N_2762);
or U2776 (N_2776,N_2709,N_2756);
nand U2777 (N_2777,N_2725,N_2771);
nand U2778 (N_2778,N_2740,N_2717);
and U2779 (N_2779,N_2705,N_2750);
or U2780 (N_2780,N_2723,N_2727);
nand U2781 (N_2781,N_2735,N_2721);
nand U2782 (N_2782,N_2764,N_2753);
nor U2783 (N_2783,N_2746,N_2718);
and U2784 (N_2784,N_2736,N_2760);
nor U2785 (N_2785,N_2772,N_2751);
nand U2786 (N_2786,N_2757,N_2761);
nand U2787 (N_2787,N_2742,N_2768);
and U2788 (N_2788,N_2763,N_2766);
nor U2789 (N_2789,N_2707,N_2734);
nand U2790 (N_2790,N_2759,N_2741);
nor U2791 (N_2791,N_2703,N_2758);
nor U2792 (N_2792,N_2732,N_2752);
and U2793 (N_2793,N_2747,N_2755);
or U2794 (N_2794,N_2708,N_2719);
nand U2795 (N_2795,N_2700,N_2743);
or U2796 (N_2796,N_2773,N_2733);
nor U2797 (N_2797,N_2738,N_2730);
and U2798 (N_2798,N_2770,N_2739);
nand U2799 (N_2799,N_2769,N_2710);
or U2800 (N_2800,N_2729,N_2745);
nand U2801 (N_2801,N_2720,N_2765);
or U2802 (N_2802,N_2724,N_2722);
nand U2803 (N_2803,N_2731,N_2749);
or U2804 (N_2804,N_2715,N_2704);
or U2805 (N_2805,N_2702,N_2701);
or U2806 (N_2806,N_2711,N_2754);
nand U2807 (N_2807,N_2716,N_2748);
and U2808 (N_2808,N_2774,N_2706);
and U2809 (N_2809,N_2728,N_2744);
nor U2810 (N_2810,N_2726,N_2712);
and U2811 (N_2811,N_2767,N_2737);
and U2812 (N_2812,N_2713,N_2757);
and U2813 (N_2813,N_2740,N_2723);
and U2814 (N_2814,N_2719,N_2735);
xnor U2815 (N_2815,N_2741,N_2714);
nor U2816 (N_2816,N_2762,N_2718);
and U2817 (N_2817,N_2713,N_2719);
and U2818 (N_2818,N_2747,N_2704);
nor U2819 (N_2819,N_2774,N_2740);
or U2820 (N_2820,N_2763,N_2706);
and U2821 (N_2821,N_2726,N_2711);
nand U2822 (N_2822,N_2731,N_2771);
nand U2823 (N_2823,N_2718,N_2720);
nand U2824 (N_2824,N_2713,N_2726);
or U2825 (N_2825,N_2714,N_2753);
nor U2826 (N_2826,N_2760,N_2767);
and U2827 (N_2827,N_2717,N_2730);
nand U2828 (N_2828,N_2758,N_2764);
nand U2829 (N_2829,N_2764,N_2731);
nor U2830 (N_2830,N_2709,N_2747);
and U2831 (N_2831,N_2751,N_2745);
nand U2832 (N_2832,N_2710,N_2713);
nor U2833 (N_2833,N_2727,N_2702);
and U2834 (N_2834,N_2749,N_2754);
nand U2835 (N_2835,N_2711,N_2712);
xor U2836 (N_2836,N_2738,N_2719);
nand U2837 (N_2837,N_2712,N_2716);
and U2838 (N_2838,N_2722,N_2700);
and U2839 (N_2839,N_2726,N_2755);
and U2840 (N_2840,N_2753,N_2701);
or U2841 (N_2841,N_2747,N_2754);
nor U2842 (N_2842,N_2712,N_2734);
or U2843 (N_2843,N_2735,N_2733);
nor U2844 (N_2844,N_2708,N_2771);
nor U2845 (N_2845,N_2740,N_2716);
or U2846 (N_2846,N_2741,N_2752);
xnor U2847 (N_2847,N_2706,N_2722);
and U2848 (N_2848,N_2765,N_2774);
nand U2849 (N_2849,N_2701,N_2719);
nor U2850 (N_2850,N_2788,N_2818);
or U2851 (N_2851,N_2825,N_2815);
nand U2852 (N_2852,N_2786,N_2841);
and U2853 (N_2853,N_2827,N_2779);
nor U2854 (N_2854,N_2782,N_2811);
or U2855 (N_2855,N_2777,N_2824);
and U2856 (N_2856,N_2833,N_2813);
and U2857 (N_2857,N_2801,N_2822);
or U2858 (N_2858,N_2844,N_2784);
or U2859 (N_2859,N_2778,N_2821);
nand U2860 (N_2860,N_2794,N_2835);
and U2861 (N_2861,N_2843,N_2807);
nand U2862 (N_2862,N_2791,N_2790);
or U2863 (N_2863,N_2849,N_2819);
nor U2864 (N_2864,N_2800,N_2780);
nor U2865 (N_2865,N_2840,N_2805);
or U2866 (N_2866,N_2797,N_2847);
nor U2867 (N_2867,N_2834,N_2814);
and U2868 (N_2868,N_2810,N_2785);
nand U2869 (N_2869,N_2817,N_2842);
or U2870 (N_2870,N_2781,N_2826);
or U2871 (N_2871,N_2812,N_2808);
and U2872 (N_2872,N_2831,N_2793);
or U2873 (N_2873,N_2845,N_2828);
or U2874 (N_2874,N_2795,N_2776);
nand U2875 (N_2875,N_2799,N_2836);
nand U2876 (N_2876,N_2783,N_2809);
or U2877 (N_2877,N_2789,N_2830);
or U2878 (N_2878,N_2804,N_2838);
or U2879 (N_2879,N_2775,N_2823);
nand U2880 (N_2880,N_2802,N_2796);
nand U2881 (N_2881,N_2839,N_2792);
nor U2882 (N_2882,N_2832,N_2829);
nor U2883 (N_2883,N_2837,N_2848);
nor U2884 (N_2884,N_2816,N_2846);
or U2885 (N_2885,N_2820,N_2803);
and U2886 (N_2886,N_2806,N_2787);
or U2887 (N_2887,N_2798,N_2822);
nor U2888 (N_2888,N_2829,N_2828);
or U2889 (N_2889,N_2775,N_2799);
or U2890 (N_2890,N_2775,N_2796);
or U2891 (N_2891,N_2783,N_2800);
or U2892 (N_2892,N_2846,N_2835);
or U2893 (N_2893,N_2817,N_2844);
nor U2894 (N_2894,N_2791,N_2801);
or U2895 (N_2895,N_2786,N_2795);
or U2896 (N_2896,N_2813,N_2834);
and U2897 (N_2897,N_2785,N_2830);
or U2898 (N_2898,N_2841,N_2836);
nand U2899 (N_2899,N_2834,N_2833);
nand U2900 (N_2900,N_2818,N_2815);
nor U2901 (N_2901,N_2779,N_2823);
and U2902 (N_2902,N_2817,N_2836);
nand U2903 (N_2903,N_2780,N_2788);
nand U2904 (N_2904,N_2809,N_2836);
xor U2905 (N_2905,N_2848,N_2819);
nand U2906 (N_2906,N_2842,N_2778);
nand U2907 (N_2907,N_2812,N_2811);
nand U2908 (N_2908,N_2786,N_2791);
nor U2909 (N_2909,N_2809,N_2829);
and U2910 (N_2910,N_2820,N_2810);
and U2911 (N_2911,N_2805,N_2798);
nand U2912 (N_2912,N_2811,N_2795);
nand U2913 (N_2913,N_2775,N_2800);
nand U2914 (N_2914,N_2789,N_2803);
or U2915 (N_2915,N_2780,N_2820);
and U2916 (N_2916,N_2834,N_2844);
and U2917 (N_2917,N_2797,N_2814);
and U2918 (N_2918,N_2792,N_2779);
nor U2919 (N_2919,N_2823,N_2848);
and U2920 (N_2920,N_2839,N_2817);
nand U2921 (N_2921,N_2787,N_2812);
nand U2922 (N_2922,N_2812,N_2778);
and U2923 (N_2923,N_2812,N_2840);
and U2924 (N_2924,N_2847,N_2835);
and U2925 (N_2925,N_2852,N_2874);
and U2926 (N_2926,N_2865,N_2870);
nor U2927 (N_2927,N_2923,N_2913);
nand U2928 (N_2928,N_2875,N_2866);
nor U2929 (N_2929,N_2851,N_2901);
or U2930 (N_2930,N_2919,N_2916);
or U2931 (N_2931,N_2873,N_2859);
nand U2932 (N_2932,N_2882,N_2904);
and U2933 (N_2933,N_2867,N_2921);
nand U2934 (N_2934,N_2890,N_2877);
xor U2935 (N_2935,N_2909,N_2888);
nand U2936 (N_2936,N_2922,N_2906);
nor U2937 (N_2937,N_2915,N_2853);
nand U2938 (N_2938,N_2857,N_2863);
nor U2939 (N_2939,N_2899,N_2918);
nor U2940 (N_2940,N_2881,N_2887);
nor U2941 (N_2941,N_2897,N_2896);
and U2942 (N_2942,N_2902,N_2893);
nand U2943 (N_2943,N_2872,N_2895);
or U2944 (N_2944,N_2910,N_2924);
or U2945 (N_2945,N_2886,N_2889);
and U2946 (N_2946,N_2907,N_2885);
nor U2947 (N_2947,N_2917,N_2880);
and U2948 (N_2948,N_2856,N_2884);
and U2949 (N_2949,N_2860,N_2892);
xor U2950 (N_2950,N_2905,N_2864);
nor U2951 (N_2951,N_2908,N_2854);
and U2952 (N_2952,N_2879,N_2855);
and U2953 (N_2953,N_2903,N_2912);
nand U2954 (N_2954,N_2862,N_2894);
and U2955 (N_2955,N_2891,N_2858);
nor U2956 (N_2956,N_2869,N_2911);
nand U2957 (N_2957,N_2850,N_2878);
nor U2958 (N_2958,N_2876,N_2868);
nand U2959 (N_2959,N_2920,N_2883);
nor U2960 (N_2960,N_2898,N_2900);
nor U2961 (N_2961,N_2861,N_2914);
nor U2962 (N_2962,N_2871,N_2864);
nand U2963 (N_2963,N_2859,N_2901);
and U2964 (N_2964,N_2912,N_2868);
and U2965 (N_2965,N_2879,N_2866);
nand U2966 (N_2966,N_2860,N_2866);
and U2967 (N_2967,N_2886,N_2873);
nor U2968 (N_2968,N_2890,N_2899);
and U2969 (N_2969,N_2897,N_2877);
nand U2970 (N_2970,N_2876,N_2914);
nand U2971 (N_2971,N_2915,N_2860);
nor U2972 (N_2972,N_2883,N_2867);
nand U2973 (N_2973,N_2909,N_2881);
or U2974 (N_2974,N_2919,N_2862);
nand U2975 (N_2975,N_2876,N_2910);
or U2976 (N_2976,N_2890,N_2862);
and U2977 (N_2977,N_2868,N_2865);
and U2978 (N_2978,N_2917,N_2906);
nor U2979 (N_2979,N_2857,N_2924);
or U2980 (N_2980,N_2861,N_2863);
nand U2981 (N_2981,N_2918,N_2857);
nand U2982 (N_2982,N_2889,N_2892);
and U2983 (N_2983,N_2877,N_2850);
nor U2984 (N_2984,N_2899,N_2876);
nand U2985 (N_2985,N_2877,N_2902);
and U2986 (N_2986,N_2903,N_2879);
and U2987 (N_2987,N_2867,N_2922);
and U2988 (N_2988,N_2899,N_2874);
xor U2989 (N_2989,N_2896,N_2910);
and U2990 (N_2990,N_2884,N_2875);
and U2991 (N_2991,N_2877,N_2866);
or U2992 (N_2992,N_2863,N_2877);
nand U2993 (N_2993,N_2875,N_2919);
or U2994 (N_2994,N_2917,N_2877);
nand U2995 (N_2995,N_2898,N_2889);
nor U2996 (N_2996,N_2906,N_2918);
nand U2997 (N_2997,N_2900,N_2893);
nor U2998 (N_2998,N_2860,N_2877);
nor U2999 (N_2999,N_2893,N_2870);
or UO_0 (O_0,N_2995,N_2936);
or UO_1 (O_1,N_2929,N_2949);
nor UO_2 (O_2,N_2977,N_2962);
nand UO_3 (O_3,N_2993,N_2958);
or UO_4 (O_4,N_2986,N_2998);
and UO_5 (O_5,N_2950,N_2952);
nor UO_6 (O_6,N_2956,N_2939);
nor UO_7 (O_7,N_2951,N_2982);
xor UO_8 (O_8,N_2935,N_2969);
nand UO_9 (O_9,N_2944,N_2968);
and UO_10 (O_10,N_2981,N_2974);
or UO_11 (O_11,N_2984,N_2990);
nand UO_12 (O_12,N_2988,N_2925);
or UO_13 (O_13,N_2985,N_2978);
nor UO_14 (O_14,N_2972,N_2964);
nor UO_15 (O_15,N_2961,N_2954);
or UO_16 (O_16,N_2971,N_2963);
and UO_17 (O_17,N_2994,N_2931);
xor UO_18 (O_18,N_2955,N_2975);
and UO_19 (O_19,N_2983,N_2973);
nand UO_20 (O_20,N_2928,N_2941);
nand UO_21 (O_21,N_2937,N_2989);
nor UO_22 (O_22,N_2946,N_2940);
xnor UO_23 (O_23,N_2932,N_2999);
nand UO_24 (O_24,N_2967,N_2948);
nand UO_25 (O_25,N_2959,N_2960);
nor UO_26 (O_26,N_2965,N_2992);
and UO_27 (O_27,N_2927,N_2947);
nand UO_28 (O_28,N_2926,N_2996);
and UO_29 (O_29,N_2970,N_2933);
nand UO_30 (O_30,N_2957,N_2938);
or UO_31 (O_31,N_2979,N_2976);
nor UO_32 (O_32,N_2966,N_2943);
or UO_33 (O_33,N_2934,N_2997);
or UO_34 (O_34,N_2953,N_2942);
or UO_35 (O_35,N_2945,N_2991);
and UO_36 (O_36,N_2930,N_2987);
or UO_37 (O_37,N_2980,N_2965);
or UO_38 (O_38,N_2942,N_2997);
or UO_39 (O_39,N_2947,N_2937);
and UO_40 (O_40,N_2994,N_2963);
or UO_41 (O_41,N_2943,N_2925);
nand UO_42 (O_42,N_2928,N_2948);
xnor UO_43 (O_43,N_2961,N_2935);
nand UO_44 (O_44,N_2949,N_2967);
nand UO_45 (O_45,N_2955,N_2994);
or UO_46 (O_46,N_2946,N_2959);
nor UO_47 (O_47,N_2990,N_2986);
or UO_48 (O_48,N_2956,N_2954);
and UO_49 (O_49,N_2974,N_2953);
nand UO_50 (O_50,N_2966,N_2945);
nor UO_51 (O_51,N_2932,N_2938);
nand UO_52 (O_52,N_2965,N_2949);
nor UO_53 (O_53,N_2999,N_2936);
xnor UO_54 (O_54,N_2946,N_2969);
nand UO_55 (O_55,N_2977,N_2960);
or UO_56 (O_56,N_2967,N_2935);
nand UO_57 (O_57,N_2976,N_2980);
nand UO_58 (O_58,N_2944,N_2940);
or UO_59 (O_59,N_2931,N_2947);
and UO_60 (O_60,N_2944,N_2954);
or UO_61 (O_61,N_2946,N_2984);
nand UO_62 (O_62,N_2989,N_2969);
nor UO_63 (O_63,N_2962,N_2991);
or UO_64 (O_64,N_2954,N_2937);
and UO_65 (O_65,N_2977,N_2944);
nor UO_66 (O_66,N_2937,N_2973);
and UO_67 (O_67,N_2993,N_2976);
and UO_68 (O_68,N_2976,N_2992);
or UO_69 (O_69,N_2995,N_2935);
nor UO_70 (O_70,N_2939,N_2935);
nand UO_71 (O_71,N_2941,N_2958);
or UO_72 (O_72,N_2958,N_2968);
nand UO_73 (O_73,N_2993,N_2981);
nor UO_74 (O_74,N_2985,N_2962);
and UO_75 (O_75,N_2979,N_2997);
nor UO_76 (O_76,N_2972,N_2991);
or UO_77 (O_77,N_2929,N_2948);
nand UO_78 (O_78,N_2998,N_2938);
nor UO_79 (O_79,N_2942,N_2949);
and UO_80 (O_80,N_2955,N_2973);
xnor UO_81 (O_81,N_2993,N_2944);
nand UO_82 (O_82,N_2932,N_2996);
or UO_83 (O_83,N_2967,N_2979);
nor UO_84 (O_84,N_2937,N_2964);
or UO_85 (O_85,N_2935,N_2978);
nand UO_86 (O_86,N_2992,N_2990);
nor UO_87 (O_87,N_2981,N_2991);
nor UO_88 (O_88,N_2979,N_2939);
nand UO_89 (O_89,N_2966,N_2946);
nor UO_90 (O_90,N_2995,N_2989);
or UO_91 (O_91,N_2963,N_2967);
and UO_92 (O_92,N_2945,N_2944);
or UO_93 (O_93,N_2978,N_2987);
or UO_94 (O_94,N_2946,N_2976);
nor UO_95 (O_95,N_2965,N_2929);
or UO_96 (O_96,N_2956,N_2943);
xnor UO_97 (O_97,N_2928,N_2993);
nor UO_98 (O_98,N_2984,N_2989);
nor UO_99 (O_99,N_2963,N_2932);
nor UO_100 (O_100,N_2941,N_2964);
or UO_101 (O_101,N_2963,N_2958);
nand UO_102 (O_102,N_2932,N_2952);
and UO_103 (O_103,N_2998,N_2945);
or UO_104 (O_104,N_2936,N_2948);
nand UO_105 (O_105,N_2930,N_2969);
nor UO_106 (O_106,N_2952,N_2957);
and UO_107 (O_107,N_2968,N_2934);
nand UO_108 (O_108,N_2931,N_2936);
xor UO_109 (O_109,N_2998,N_2978);
nor UO_110 (O_110,N_2984,N_2970);
nand UO_111 (O_111,N_2971,N_2989);
nand UO_112 (O_112,N_2971,N_2975);
or UO_113 (O_113,N_2987,N_2956);
xor UO_114 (O_114,N_2929,N_2926);
nand UO_115 (O_115,N_2927,N_2963);
nor UO_116 (O_116,N_2989,N_2950);
nor UO_117 (O_117,N_2973,N_2977);
nor UO_118 (O_118,N_2980,N_2953);
nand UO_119 (O_119,N_2984,N_2947);
and UO_120 (O_120,N_2976,N_2935);
nor UO_121 (O_121,N_2974,N_2993);
and UO_122 (O_122,N_2952,N_2987);
or UO_123 (O_123,N_2967,N_2969);
nand UO_124 (O_124,N_2950,N_2973);
and UO_125 (O_125,N_2943,N_2978);
or UO_126 (O_126,N_2941,N_2950);
nand UO_127 (O_127,N_2925,N_2989);
or UO_128 (O_128,N_2949,N_2928);
nand UO_129 (O_129,N_2952,N_2986);
nand UO_130 (O_130,N_2932,N_2969);
nor UO_131 (O_131,N_2990,N_2982);
and UO_132 (O_132,N_2947,N_2935);
or UO_133 (O_133,N_2989,N_2980);
or UO_134 (O_134,N_2931,N_2953);
or UO_135 (O_135,N_2961,N_2931);
nand UO_136 (O_136,N_2935,N_2925);
nor UO_137 (O_137,N_2986,N_2940);
xnor UO_138 (O_138,N_2959,N_2984);
nand UO_139 (O_139,N_2980,N_2994);
and UO_140 (O_140,N_2981,N_2938);
nor UO_141 (O_141,N_2996,N_2941);
or UO_142 (O_142,N_2951,N_2948);
and UO_143 (O_143,N_2932,N_2970);
nor UO_144 (O_144,N_2989,N_2972);
and UO_145 (O_145,N_2957,N_2934);
nor UO_146 (O_146,N_2957,N_2999);
and UO_147 (O_147,N_2973,N_2958);
nand UO_148 (O_148,N_2929,N_2956);
nand UO_149 (O_149,N_2994,N_2976);
xnor UO_150 (O_150,N_2941,N_2972);
and UO_151 (O_151,N_2993,N_2989);
and UO_152 (O_152,N_2950,N_2931);
xnor UO_153 (O_153,N_2946,N_2975);
nand UO_154 (O_154,N_2989,N_2942);
or UO_155 (O_155,N_2977,N_2953);
or UO_156 (O_156,N_2976,N_2944);
and UO_157 (O_157,N_2972,N_2926);
or UO_158 (O_158,N_2956,N_2949);
nand UO_159 (O_159,N_2999,N_2993);
nor UO_160 (O_160,N_2965,N_2938);
nand UO_161 (O_161,N_2961,N_2970);
and UO_162 (O_162,N_2951,N_2966);
nand UO_163 (O_163,N_2936,N_2939);
nor UO_164 (O_164,N_2989,N_2994);
nor UO_165 (O_165,N_2934,N_2974);
or UO_166 (O_166,N_2961,N_2937);
and UO_167 (O_167,N_2997,N_2975);
or UO_168 (O_168,N_2958,N_2944);
and UO_169 (O_169,N_2950,N_2960);
nand UO_170 (O_170,N_2928,N_2939);
or UO_171 (O_171,N_2976,N_2972);
xnor UO_172 (O_172,N_2951,N_2983);
nor UO_173 (O_173,N_2982,N_2957);
and UO_174 (O_174,N_2953,N_2985);
and UO_175 (O_175,N_2989,N_2947);
nand UO_176 (O_176,N_2938,N_2970);
xnor UO_177 (O_177,N_2954,N_2980);
or UO_178 (O_178,N_2977,N_2957);
or UO_179 (O_179,N_2974,N_2928);
nor UO_180 (O_180,N_2931,N_2993);
nor UO_181 (O_181,N_2960,N_2983);
or UO_182 (O_182,N_2936,N_2935);
nor UO_183 (O_183,N_2935,N_2937);
and UO_184 (O_184,N_2986,N_2937);
and UO_185 (O_185,N_2971,N_2970);
nand UO_186 (O_186,N_2948,N_2973);
nor UO_187 (O_187,N_2936,N_2945);
or UO_188 (O_188,N_2947,N_2946);
nand UO_189 (O_189,N_2941,N_2974);
and UO_190 (O_190,N_2938,N_2928);
or UO_191 (O_191,N_2941,N_2960);
nand UO_192 (O_192,N_2947,N_2945);
and UO_193 (O_193,N_2928,N_2965);
or UO_194 (O_194,N_2943,N_2990);
nor UO_195 (O_195,N_2947,N_2991);
nor UO_196 (O_196,N_2942,N_2976);
and UO_197 (O_197,N_2943,N_2931);
nand UO_198 (O_198,N_2931,N_2955);
nand UO_199 (O_199,N_2949,N_2934);
and UO_200 (O_200,N_2992,N_2987);
and UO_201 (O_201,N_2981,N_2964);
and UO_202 (O_202,N_2935,N_2996);
or UO_203 (O_203,N_2977,N_2993);
nor UO_204 (O_204,N_2934,N_2961);
and UO_205 (O_205,N_2938,N_2974);
or UO_206 (O_206,N_2964,N_2934);
nor UO_207 (O_207,N_2993,N_2941);
and UO_208 (O_208,N_2990,N_2959);
and UO_209 (O_209,N_2935,N_2981);
and UO_210 (O_210,N_2955,N_2969);
nor UO_211 (O_211,N_2947,N_2976);
or UO_212 (O_212,N_2931,N_2934);
nand UO_213 (O_213,N_2960,N_2969);
nor UO_214 (O_214,N_2946,N_2996);
nor UO_215 (O_215,N_2936,N_2959);
or UO_216 (O_216,N_2991,N_2939);
nor UO_217 (O_217,N_2972,N_2984);
and UO_218 (O_218,N_2964,N_2984);
nand UO_219 (O_219,N_2966,N_2955);
and UO_220 (O_220,N_2994,N_2941);
or UO_221 (O_221,N_2944,N_2959);
nand UO_222 (O_222,N_2985,N_2943);
and UO_223 (O_223,N_2953,N_2959);
nor UO_224 (O_224,N_2962,N_2941);
and UO_225 (O_225,N_2936,N_2973);
and UO_226 (O_226,N_2942,N_2994);
or UO_227 (O_227,N_2955,N_2939);
nand UO_228 (O_228,N_2931,N_2987);
nand UO_229 (O_229,N_2936,N_2996);
or UO_230 (O_230,N_2985,N_2926);
and UO_231 (O_231,N_2965,N_2977);
nor UO_232 (O_232,N_2995,N_2974);
nor UO_233 (O_233,N_2980,N_2947);
and UO_234 (O_234,N_2950,N_2938);
nand UO_235 (O_235,N_2955,N_2985);
and UO_236 (O_236,N_2968,N_2996);
or UO_237 (O_237,N_2990,N_2927);
or UO_238 (O_238,N_2930,N_2958);
xor UO_239 (O_239,N_2997,N_2936);
and UO_240 (O_240,N_2988,N_2927);
and UO_241 (O_241,N_2999,N_2933);
or UO_242 (O_242,N_2949,N_2926);
nand UO_243 (O_243,N_2974,N_2998);
and UO_244 (O_244,N_2993,N_2932);
nand UO_245 (O_245,N_2978,N_2936);
and UO_246 (O_246,N_2927,N_2956);
or UO_247 (O_247,N_2989,N_2927);
and UO_248 (O_248,N_2942,N_2966);
nor UO_249 (O_249,N_2961,N_2930);
nand UO_250 (O_250,N_2978,N_2945);
and UO_251 (O_251,N_2959,N_2928);
or UO_252 (O_252,N_2958,N_2981);
and UO_253 (O_253,N_2987,N_2991);
nand UO_254 (O_254,N_2982,N_2967);
nor UO_255 (O_255,N_2963,N_2962);
xor UO_256 (O_256,N_2981,N_2942);
nand UO_257 (O_257,N_2971,N_2986);
nor UO_258 (O_258,N_2931,N_2940);
nand UO_259 (O_259,N_2986,N_2957);
nand UO_260 (O_260,N_2952,N_2929);
nor UO_261 (O_261,N_2976,N_2939);
nor UO_262 (O_262,N_2996,N_2969);
or UO_263 (O_263,N_2968,N_2985);
nand UO_264 (O_264,N_2972,N_2973);
nor UO_265 (O_265,N_2939,N_2988);
and UO_266 (O_266,N_2975,N_2991);
and UO_267 (O_267,N_2992,N_2961);
and UO_268 (O_268,N_2925,N_2956);
nand UO_269 (O_269,N_2937,N_2962);
or UO_270 (O_270,N_2991,N_2976);
or UO_271 (O_271,N_2940,N_2967);
nand UO_272 (O_272,N_2935,N_2949);
or UO_273 (O_273,N_2981,N_2978);
nor UO_274 (O_274,N_2994,N_2926);
nand UO_275 (O_275,N_2980,N_2938);
or UO_276 (O_276,N_2997,N_2948);
or UO_277 (O_277,N_2943,N_2983);
nor UO_278 (O_278,N_2993,N_2943);
nand UO_279 (O_279,N_2978,N_2955);
nor UO_280 (O_280,N_2967,N_2990);
nand UO_281 (O_281,N_2946,N_2999);
and UO_282 (O_282,N_2992,N_2928);
or UO_283 (O_283,N_2963,N_2951);
or UO_284 (O_284,N_2930,N_2991);
nand UO_285 (O_285,N_2925,N_2953);
nor UO_286 (O_286,N_2974,N_2957);
or UO_287 (O_287,N_2998,N_2939);
and UO_288 (O_288,N_2995,N_2968);
or UO_289 (O_289,N_2948,N_2957);
nor UO_290 (O_290,N_2934,N_2928);
nor UO_291 (O_291,N_2932,N_2931);
nand UO_292 (O_292,N_2987,N_2980);
and UO_293 (O_293,N_2942,N_2963);
xor UO_294 (O_294,N_2969,N_2941);
nand UO_295 (O_295,N_2984,N_2999);
and UO_296 (O_296,N_2981,N_2931);
nor UO_297 (O_297,N_2936,N_2992);
nor UO_298 (O_298,N_2959,N_2952);
nor UO_299 (O_299,N_2977,N_2940);
or UO_300 (O_300,N_2976,N_2930);
or UO_301 (O_301,N_2934,N_2988);
or UO_302 (O_302,N_2957,N_2932);
nor UO_303 (O_303,N_2966,N_2944);
or UO_304 (O_304,N_2968,N_2963);
and UO_305 (O_305,N_2955,N_2926);
nor UO_306 (O_306,N_2974,N_2947);
and UO_307 (O_307,N_2949,N_2970);
xor UO_308 (O_308,N_2993,N_2957);
nand UO_309 (O_309,N_2968,N_2972);
nand UO_310 (O_310,N_2929,N_2988);
and UO_311 (O_311,N_2927,N_2981);
and UO_312 (O_312,N_2935,N_2953);
or UO_313 (O_313,N_2957,N_2926);
or UO_314 (O_314,N_2957,N_2955);
and UO_315 (O_315,N_2958,N_2965);
nand UO_316 (O_316,N_2992,N_2946);
nor UO_317 (O_317,N_2946,N_2995);
nor UO_318 (O_318,N_2965,N_2986);
xor UO_319 (O_319,N_2956,N_2940);
nand UO_320 (O_320,N_2973,N_2978);
nand UO_321 (O_321,N_2955,N_2967);
nor UO_322 (O_322,N_2940,N_2988);
nor UO_323 (O_323,N_2971,N_2995);
nor UO_324 (O_324,N_2980,N_2942);
nand UO_325 (O_325,N_2958,N_2976);
or UO_326 (O_326,N_2954,N_2993);
and UO_327 (O_327,N_2961,N_2955);
or UO_328 (O_328,N_2967,N_2991);
nor UO_329 (O_329,N_2982,N_2977);
nor UO_330 (O_330,N_2987,N_2977);
nor UO_331 (O_331,N_2987,N_2942);
nor UO_332 (O_332,N_2960,N_2995);
nand UO_333 (O_333,N_2935,N_2986);
nor UO_334 (O_334,N_2954,N_2990);
xor UO_335 (O_335,N_2942,N_2932);
nand UO_336 (O_336,N_2970,N_2930);
and UO_337 (O_337,N_2977,N_2929);
or UO_338 (O_338,N_2940,N_2964);
and UO_339 (O_339,N_2925,N_2973);
or UO_340 (O_340,N_2981,N_2939);
or UO_341 (O_341,N_2973,N_2979);
nand UO_342 (O_342,N_2958,N_2984);
nor UO_343 (O_343,N_2973,N_2996);
or UO_344 (O_344,N_2984,N_2949);
nand UO_345 (O_345,N_2945,N_2977);
and UO_346 (O_346,N_2997,N_2976);
or UO_347 (O_347,N_2994,N_2992);
nor UO_348 (O_348,N_2930,N_2980);
nand UO_349 (O_349,N_2981,N_2946);
nor UO_350 (O_350,N_2956,N_2932);
or UO_351 (O_351,N_2939,N_2984);
nand UO_352 (O_352,N_2951,N_2954);
nor UO_353 (O_353,N_2959,N_2995);
or UO_354 (O_354,N_2967,N_2931);
or UO_355 (O_355,N_2973,N_2930);
or UO_356 (O_356,N_2963,N_2933);
and UO_357 (O_357,N_2937,N_2981);
nor UO_358 (O_358,N_2946,N_2926);
nor UO_359 (O_359,N_2943,N_2988);
nor UO_360 (O_360,N_2961,N_2964);
nor UO_361 (O_361,N_2944,N_2951);
or UO_362 (O_362,N_2975,N_2938);
nand UO_363 (O_363,N_2985,N_2933);
nand UO_364 (O_364,N_2930,N_2982);
or UO_365 (O_365,N_2958,N_2926);
nor UO_366 (O_366,N_2933,N_2993);
nand UO_367 (O_367,N_2954,N_2982);
nand UO_368 (O_368,N_2937,N_2975);
or UO_369 (O_369,N_2952,N_2964);
and UO_370 (O_370,N_2948,N_2980);
or UO_371 (O_371,N_2949,N_2937);
xnor UO_372 (O_372,N_2993,N_2959);
or UO_373 (O_373,N_2996,N_2950);
or UO_374 (O_374,N_2982,N_2979);
or UO_375 (O_375,N_2961,N_2971);
nor UO_376 (O_376,N_2998,N_2934);
nand UO_377 (O_377,N_2956,N_2970);
or UO_378 (O_378,N_2999,N_2934);
nand UO_379 (O_379,N_2940,N_2972);
nand UO_380 (O_380,N_2929,N_2958);
or UO_381 (O_381,N_2926,N_2947);
or UO_382 (O_382,N_2930,N_2983);
nand UO_383 (O_383,N_2938,N_2979);
or UO_384 (O_384,N_2962,N_2971);
nand UO_385 (O_385,N_2959,N_2991);
or UO_386 (O_386,N_2988,N_2953);
or UO_387 (O_387,N_2951,N_2946);
and UO_388 (O_388,N_2955,N_2945);
nor UO_389 (O_389,N_2999,N_2967);
nand UO_390 (O_390,N_2971,N_2941);
nor UO_391 (O_391,N_2962,N_2945);
nand UO_392 (O_392,N_2986,N_2964);
xor UO_393 (O_393,N_2998,N_2933);
nor UO_394 (O_394,N_2975,N_2965);
nor UO_395 (O_395,N_2968,N_2962);
nor UO_396 (O_396,N_2948,N_2942);
and UO_397 (O_397,N_2943,N_2967);
or UO_398 (O_398,N_2989,N_2962);
nor UO_399 (O_399,N_2976,N_2963);
nor UO_400 (O_400,N_2991,N_2978);
nand UO_401 (O_401,N_2945,N_2954);
or UO_402 (O_402,N_2971,N_2952);
nor UO_403 (O_403,N_2943,N_2961);
or UO_404 (O_404,N_2953,N_2997);
or UO_405 (O_405,N_2984,N_2986);
or UO_406 (O_406,N_2960,N_2940);
and UO_407 (O_407,N_2971,N_2954);
and UO_408 (O_408,N_2966,N_2936);
and UO_409 (O_409,N_2925,N_2967);
and UO_410 (O_410,N_2970,N_2983);
or UO_411 (O_411,N_2929,N_2954);
or UO_412 (O_412,N_2952,N_2977);
nand UO_413 (O_413,N_2997,N_2970);
and UO_414 (O_414,N_2959,N_2968);
nand UO_415 (O_415,N_2981,N_2999);
and UO_416 (O_416,N_2999,N_2972);
and UO_417 (O_417,N_2989,N_2992);
nor UO_418 (O_418,N_2944,N_2964);
and UO_419 (O_419,N_2997,N_2946);
xnor UO_420 (O_420,N_2995,N_2951);
or UO_421 (O_421,N_2950,N_2977);
nand UO_422 (O_422,N_2946,N_2936);
nand UO_423 (O_423,N_2961,N_2926);
and UO_424 (O_424,N_2928,N_2942);
nor UO_425 (O_425,N_2997,N_2962);
nor UO_426 (O_426,N_2972,N_2966);
nor UO_427 (O_427,N_2952,N_2951);
or UO_428 (O_428,N_2964,N_2943);
and UO_429 (O_429,N_2946,N_2950);
or UO_430 (O_430,N_2939,N_2946);
nand UO_431 (O_431,N_2972,N_2943);
nor UO_432 (O_432,N_2946,N_2985);
nor UO_433 (O_433,N_2934,N_2983);
or UO_434 (O_434,N_2984,N_2942);
or UO_435 (O_435,N_2987,N_2972);
or UO_436 (O_436,N_2934,N_2996);
nand UO_437 (O_437,N_2966,N_2930);
nor UO_438 (O_438,N_2995,N_2987);
or UO_439 (O_439,N_2930,N_2949);
and UO_440 (O_440,N_2973,N_2990);
and UO_441 (O_441,N_2929,N_2934);
nor UO_442 (O_442,N_2987,N_2944);
nor UO_443 (O_443,N_2958,N_2950);
nand UO_444 (O_444,N_2933,N_2960);
and UO_445 (O_445,N_2953,N_2940);
or UO_446 (O_446,N_2989,N_2945);
nand UO_447 (O_447,N_2970,N_2992);
or UO_448 (O_448,N_2941,N_2945);
or UO_449 (O_449,N_2945,N_2969);
nand UO_450 (O_450,N_2954,N_2996);
nor UO_451 (O_451,N_2972,N_2982);
nor UO_452 (O_452,N_2959,N_2940);
or UO_453 (O_453,N_2970,N_2954);
or UO_454 (O_454,N_2996,N_2976);
xnor UO_455 (O_455,N_2950,N_2933);
and UO_456 (O_456,N_2986,N_2953);
and UO_457 (O_457,N_2930,N_2988);
and UO_458 (O_458,N_2938,N_2949);
nand UO_459 (O_459,N_2972,N_2993);
and UO_460 (O_460,N_2927,N_2943);
nand UO_461 (O_461,N_2976,N_2957);
xnor UO_462 (O_462,N_2947,N_2995);
or UO_463 (O_463,N_2962,N_2943);
nor UO_464 (O_464,N_2967,N_2962);
nand UO_465 (O_465,N_2972,N_2929);
nand UO_466 (O_466,N_2986,N_2999);
nor UO_467 (O_467,N_2999,N_2939);
or UO_468 (O_468,N_2969,N_2928);
nor UO_469 (O_469,N_2976,N_2966);
and UO_470 (O_470,N_2989,N_2990);
nand UO_471 (O_471,N_2995,N_2950);
or UO_472 (O_472,N_2925,N_2986);
and UO_473 (O_473,N_2954,N_2946);
and UO_474 (O_474,N_2988,N_2965);
nor UO_475 (O_475,N_2940,N_2949);
xnor UO_476 (O_476,N_2975,N_2953);
nor UO_477 (O_477,N_2947,N_2951);
and UO_478 (O_478,N_2938,N_2963);
nand UO_479 (O_479,N_2981,N_2990);
and UO_480 (O_480,N_2979,N_2993);
xor UO_481 (O_481,N_2926,N_2986);
nand UO_482 (O_482,N_2951,N_2975);
nand UO_483 (O_483,N_2934,N_2975);
nand UO_484 (O_484,N_2956,N_2995);
and UO_485 (O_485,N_2948,N_2938);
or UO_486 (O_486,N_2994,N_2945);
nand UO_487 (O_487,N_2941,N_2957);
and UO_488 (O_488,N_2957,N_2925);
or UO_489 (O_489,N_2966,N_2937);
nand UO_490 (O_490,N_2992,N_2929);
and UO_491 (O_491,N_2986,N_2995);
nor UO_492 (O_492,N_2998,N_2973);
nor UO_493 (O_493,N_2949,N_2953);
or UO_494 (O_494,N_2986,N_2979);
nand UO_495 (O_495,N_2927,N_2976);
or UO_496 (O_496,N_2991,N_2943);
and UO_497 (O_497,N_2974,N_2984);
or UO_498 (O_498,N_2955,N_2962);
and UO_499 (O_499,N_2948,N_2991);
endmodule