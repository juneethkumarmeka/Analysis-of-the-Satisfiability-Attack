module basic_2000_20000_2500_5_levels_10xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
and U0 (N_0,In_1806,In_540);
or U1 (N_1,In_1337,In_171);
xor U2 (N_2,In_309,In_1656);
nand U3 (N_3,In_1930,In_1442);
nor U4 (N_4,In_1854,In_1993);
nand U5 (N_5,In_1435,In_659);
and U6 (N_6,In_429,In_1328);
xnor U7 (N_7,In_924,In_201);
xor U8 (N_8,In_173,In_1549);
xnor U9 (N_9,In_813,In_981);
xor U10 (N_10,In_424,In_1912);
or U11 (N_11,In_392,In_591);
or U12 (N_12,In_1933,In_573);
or U13 (N_13,In_1474,In_1464);
xnor U14 (N_14,In_1770,In_665);
or U15 (N_15,In_1724,In_1762);
and U16 (N_16,In_1106,In_1632);
xor U17 (N_17,In_966,In_1518);
or U18 (N_18,In_1022,In_438);
nand U19 (N_19,In_345,In_1049);
or U20 (N_20,In_751,In_613);
or U21 (N_21,In_1172,In_163);
xnor U22 (N_22,In_445,In_544);
nor U23 (N_23,In_509,In_1669);
or U24 (N_24,In_736,In_1571);
or U25 (N_25,In_449,In_583);
or U26 (N_26,In_6,In_1901);
nand U27 (N_27,In_1784,In_258);
nand U28 (N_28,In_1433,In_1056);
or U29 (N_29,In_1396,In_842);
xor U30 (N_30,In_1871,In_1612);
nand U31 (N_31,In_335,In_437);
xor U32 (N_32,In_655,In_988);
nand U33 (N_33,In_231,In_1849);
and U34 (N_34,In_1230,In_1345);
nor U35 (N_35,In_306,In_1940);
xor U36 (N_36,In_79,In_1629);
or U37 (N_37,In_1832,In_182);
nand U38 (N_38,In_1759,In_1239);
xor U39 (N_39,In_467,In_1187);
nor U40 (N_40,In_77,In_1662);
or U41 (N_41,In_699,In_1405);
nor U42 (N_42,In_564,In_1348);
and U43 (N_43,In_570,In_35);
or U44 (N_44,In_1419,In_1979);
nand U45 (N_45,In_1025,In_1261);
xnor U46 (N_46,In_831,In_688);
and U47 (N_47,In_774,In_280);
or U48 (N_48,In_1986,In_1382);
or U49 (N_49,In_1924,In_1175);
nor U50 (N_50,In_1211,In_958);
xnor U51 (N_51,In_1248,In_1519);
xor U52 (N_52,In_183,In_379);
and U53 (N_53,In_1585,In_1942);
or U54 (N_54,In_1977,In_1387);
or U55 (N_55,In_320,In_17);
or U56 (N_56,In_1263,In_1614);
and U57 (N_57,In_418,In_1658);
and U58 (N_58,In_543,In_1190);
and U59 (N_59,In_610,In_1216);
or U60 (N_60,In_356,In_928);
or U61 (N_61,In_1424,In_542);
or U62 (N_62,In_944,In_1959);
nor U63 (N_63,In_90,In_1031);
and U64 (N_64,In_868,In_760);
xor U65 (N_65,In_1053,In_1683);
xor U66 (N_66,In_649,In_965);
nor U67 (N_67,In_1033,In_128);
xor U68 (N_68,In_210,In_1637);
nand U69 (N_69,In_1293,In_743);
nor U70 (N_70,In_1377,In_1787);
and U71 (N_71,In_553,In_1343);
xor U72 (N_72,In_1452,In_1502);
nand U73 (N_73,In_1587,In_755);
nor U74 (N_74,In_1489,In_1898);
and U75 (N_75,In_219,In_1554);
and U76 (N_76,In_1602,In_1911);
and U77 (N_77,In_839,In_586);
and U78 (N_78,In_880,In_1860);
and U79 (N_79,In_1356,In_1284);
or U80 (N_80,In_908,In_174);
nand U81 (N_81,In_1060,In_945);
and U82 (N_82,In_1527,In_1218);
and U83 (N_83,In_1226,In_1093);
nor U84 (N_84,In_1445,In_888);
or U85 (N_85,In_188,In_702);
nand U86 (N_86,In_1690,In_1529);
nand U87 (N_87,In_1517,In_52);
nand U88 (N_88,In_834,In_512);
nor U89 (N_89,In_1397,In_47);
nor U90 (N_90,In_11,In_346);
and U91 (N_91,In_1707,In_1501);
and U92 (N_92,In_1670,In_1944);
and U93 (N_93,In_1956,In_794);
or U94 (N_94,In_236,In_187);
nor U95 (N_95,In_68,In_176);
nand U96 (N_96,In_1165,In_646);
nor U97 (N_97,In_826,In_1594);
and U98 (N_98,In_377,In_1880);
and U99 (N_99,In_48,In_284);
nor U100 (N_100,In_775,In_262);
and U101 (N_101,In_1753,In_471);
xnor U102 (N_102,In_1668,In_1334);
xnor U103 (N_103,In_724,In_313);
and U104 (N_104,In_1100,In_1644);
nand U105 (N_105,In_216,In_1472);
and U106 (N_106,In_869,In_770);
xor U107 (N_107,In_259,In_1176);
nor U108 (N_108,In_1024,In_264);
and U109 (N_109,In_1941,In_1755);
xor U110 (N_110,In_1819,In_1610);
or U111 (N_111,In_817,In_987);
nor U112 (N_112,In_820,In_1283);
xnor U113 (N_113,In_1758,In_1508);
or U114 (N_114,In_1734,In_582);
or U115 (N_115,In_539,In_365);
nor U116 (N_116,In_239,In_1627);
nor U117 (N_117,In_1116,In_1505);
nor U118 (N_118,In_1254,In_885);
and U119 (N_119,In_864,In_127);
nor U120 (N_120,In_914,In_205);
nand U121 (N_121,In_1423,In_593);
nand U122 (N_122,In_12,In_122);
nand U123 (N_123,In_1847,In_937);
xor U124 (N_124,In_629,In_53);
nor U125 (N_125,In_223,In_490);
nor U126 (N_126,In_685,In_828);
or U127 (N_127,In_631,In_112);
and U128 (N_128,In_177,In_472);
or U129 (N_129,In_1544,In_1076);
nor U130 (N_130,In_461,In_62);
and U131 (N_131,In_920,In_951);
nor U132 (N_132,In_37,In_228);
nor U133 (N_133,In_404,In_768);
and U134 (N_134,In_907,In_1380);
xor U135 (N_135,In_861,In_846);
xor U136 (N_136,In_161,In_1065);
nor U137 (N_137,In_891,In_63);
and U138 (N_138,In_1330,In_138);
and U139 (N_139,In_1524,In_1055);
and U140 (N_140,In_1513,In_1691);
or U141 (N_141,In_633,In_567);
and U142 (N_142,In_957,In_1675);
or U143 (N_143,In_456,In_1272);
or U144 (N_144,In_873,In_855);
nor U145 (N_145,In_1748,In_853);
and U146 (N_146,In_508,In_1362);
nand U147 (N_147,In_1004,In_642);
or U148 (N_148,In_984,In_1915);
and U149 (N_149,In_1546,In_1922);
or U150 (N_150,In_42,In_263);
nand U151 (N_151,In_1998,In_1960);
or U152 (N_152,In_1583,In_1233);
nand U153 (N_153,In_150,In_1968);
xor U154 (N_154,In_65,In_754);
nand U155 (N_155,In_380,In_1002);
nor U156 (N_156,In_1167,In_918);
or U157 (N_157,In_439,In_355);
xor U158 (N_158,In_1342,In_1201);
and U159 (N_159,In_1574,In_144);
nand U160 (N_160,In_712,In_366);
or U161 (N_161,In_511,In_534);
nand U162 (N_162,In_1750,In_874);
xor U163 (N_163,In_190,In_1007);
xnor U164 (N_164,In_501,In_919);
or U165 (N_165,In_316,In_151);
or U166 (N_166,In_103,In_589);
or U167 (N_167,In_268,In_1820);
and U168 (N_168,In_1359,In_1885);
xnor U169 (N_169,In_1962,In_980);
nor U170 (N_170,In_1973,In_369);
or U171 (N_171,In_1028,In_393);
nand U172 (N_172,In_1247,In_1312);
or U173 (N_173,In_506,In_1443);
or U174 (N_174,In_1383,In_332);
or U175 (N_175,In_640,In_178);
or U176 (N_176,In_632,In_1624);
or U177 (N_177,In_795,In_413);
nand U178 (N_178,In_906,In_569);
nand U179 (N_179,In_1034,In_108);
and U180 (N_180,In_91,In_1324);
and U181 (N_181,In_695,In_1005);
or U182 (N_182,In_224,In_1141);
nand U183 (N_183,In_1331,In_1816);
and U184 (N_184,In_1884,In_208);
xnor U185 (N_185,In_1622,In_1696);
nor U186 (N_186,In_478,In_661);
and U187 (N_187,In_587,In_1634);
and U188 (N_188,In_27,In_1064);
or U189 (N_189,In_1238,In_1179);
nand U190 (N_190,In_1109,In_1763);
and U191 (N_191,In_1789,In_1790);
or U192 (N_192,In_1449,In_1409);
nand U193 (N_193,In_1655,In_1894);
and U194 (N_194,In_574,In_1484);
xor U195 (N_195,In_745,In_708);
nand U196 (N_196,In_1754,In_1666);
or U197 (N_197,In_707,In_293);
or U198 (N_198,In_931,In_1514);
and U199 (N_199,In_520,In_358);
nand U200 (N_200,In_1298,In_1794);
xor U201 (N_201,In_865,In_1678);
xnor U202 (N_202,In_590,In_292);
xnor U203 (N_203,In_1204,In_851);
nand U204 (N_204,In_1453,In_962);
xnor U205 (N_205,In_305,In_71);
and U206 (N_206,In_1318,In_247);
and U207 (N_207,In_1999,In_73);
and U208 (N_208,In_222,In_212);
xor U209 (N_209,In_1569,In_1041);
nor U210 (N_210,In_1605,In_694);
or U211 (N_211,In_1378,In_1067);
nor U212 (N_212,In_271,In_1098);
nor U213 (N_213,In_1352,In_1866);
nand U214 (N_214,In_1760,In_1203);
xnor U215 (N_215,In_318,In_39);
and U216 (N_216,In_1843,In_442);
or U217 (N_217,In_1925,In_902);
and U218 (N_218,In_617,In_1596);
or U219 (N_219,In_1835,In_1465);
and U220 (N_220,In_771,In_1647);
and U221 (N_221,In_480,In_1243);
or U222 (N_222,In_1333,In_1083);
nand U223 (N_223,In_1928,In_310);
or U224 (N_224,In_460,In_1711);
nor U225 (N_225,In_719,In_1207);
nand U226 (N_226,In_1000,In_384);
or U227 (N_227,In_1559,In_1557);
or U228 (N_228,In_1572,In_1892);
nand U229 (N_229,In_74,In_1623);
nand U230 (N_230,In_630,In_1972);
nor U231 (N_231,In_110,In_1808);
or U232 (N_232,In_608,In_1511);
nand U233 (N_233,In_457,In_1828);
or U234 (N_234,In_1865,In_535);
and U235 (N_235,In_470,In_936);
and U236 (N_236,In_602,In_515);
nand U237 (N_237,In_961,In_1987);
and U238 (N_238,In_778,In_1277);
or U239 (N_239,In_235,In_1054);
xor U240 (N_240,In_776,In_1607);
or U241 (N_241,In_1209,In_378);
and U242 (N_242,In_1926,In_272);
nor U243 (N_243,In_191,In_837);
nor U244 (N_244,In_514,In_730);
nor U245 (N_245,In_1494,In_725);
nand U246 (N_246,In_25,In_1967);
or U247 (N_247,In_1591,In_1829);
and U248 (N_248,In_376,In_850);
nand U249 (N_249,In_882,In_1151);
or U250 (N_250,In_938,In_519);
or U251 (N_251,In_428,In_815);
nand U252 (N_252,In_166,In_1182);
and U253 (N_253,In_580,In_1032);
nand U254 (N_254,In_890,In_1325);
xnor U255 (N_255,In_1438,In_893);
nand U256 (N_256,In_81,In_1705);
nand U257 (N_257,In_1604,In_1778);
and U258 (N_258,In_1061,In_1785);
xor U259 (N_259,In_18,In_996);
or U260 (N_260,In_835,In_565);
nand U261 (N_261,In_1249,In_1154);
xor U262 (N_262,In_1966,In_1767);
nand U263 (N_263,In_1115,In_1089);
xnor U264 (N_264,In_1456,In_748);
nand U265 (N_265,In_1952,In_1457);
nor U266 (N_266,In_1376,In_13);
nand U267 (N_267,In_967,In_145);
nand U268 (N_268,In_114,In_599);
nand U269 (N_269,In_1162,In_1788);
and U270 (N_270,In_548,In_1772);
nor U271 (N_271,In_1174,In_696);
xor U272 (N_272,In_1426,In_948);
nor U273 (N_273,In_761,In_225);
and U274 (N_274,In_731,In_315);
and U275 (N_275,In_1493,In_611);
or U276 (N_276,In_185,In_1184);
or U277 (N_277,In_1398,In_741);
nor U278 (N_278,In_1598,In_1868);
xor U279 (N_279,In_1907,In_999);
or U280 (N_280,In_381,In_129);
nor U281 (N_281,In_1856,In_1095);
or U282 (N_282,In_1262,In_175);
nor U283 (N_283,In_673,In_648);
and U284 (N_284,In_419,In_1520);
nand U285 (N_285,In_1870,In_406);
and U286 (N_286,In_435,In_1984);
and U287 (N_287,In_949,In_1732);
nor U288 (N_288,In_551,In_1580);
xnor U289 (N_289,In_152,In_1232);
nand U290 (N_290,In_1346,In_275);
nand U291 (N_291,In_141,In_450);
and U292 (N_292,In_1042,In_94);
xor U293 (N_293,In_977,In_1840);
nor U294 (N_294,In_325,In_780);
and U295 (N_295,In_1385,In_1428);
xnor U296 (N_296,In_337,In_1235);
nor U297 (N_297,In_1934,In_1859);
nand U298 (N_298,In_1741,In_1953);
nor U299 (N_299,In_1834,In_1208);
xnor U300 (N_300,In_1735,In_716);
and U301 (N_301,In_1857,In_464);
or U302 (N_302,In_486,In_1475);
xor U303 (N_303,In_1739,In_93);
or U304 (N_304,In_19,In_1918);
and U305 (N_305,In_69,In_604);
or U306 (N_306,In_1771,In_821);
nor U307 (N_307,In_1756,In_405);
nor U308 (N_308,In_703,In_773);
nand U309 (N_309,In_1391,In_1747);
xnor U310 (N_310,In_1228,In_1895);
xor U311 (N_311,In_959,In_441);
nor U312 (N_312,In_623,In_1757);
and U313 (N_313,In_607,In_498);
nand U314 (N_314,In_943,In_915);
and U315 (N_315,In_822,In_1698);
nor U316 (N_316,In_1841,In_522);
and U317 (N_317,In_818,In_1509);
and U318 (N_318,In_339,In_227);
nor U319 (N_319,In_1680,In_85);
xnor U320 (N_320,In_147,In_1412);
nor U321 (N_321,In_287,In_1677);
xor U322 (N_322,In_1321,In_95);
nor U323 (N_323,In_705,In_1581);
nor U324 (N_324,In_283,In_1799);
nor U325 (N_325,In_1145,In_1242);
or U326 (N_326,In_1699,In_321);
or U327 (N_327,In_1467,In_1903);
and U328 (N_328,In_1310,In_1921);
xor U329 (N_329,In_1996,In_83);
xnor U330 (N_330,In_1286,In_1401);
xor U331 (N_331,In_804,In_1477);
and U332 (N_332,In_273,In_679);
nand U333 (N_333,In_326,In_1101);
and U334 (N_334,In_808,In_232);
xnor U335 (N_335,In_1910,In_1439);
or U336 (N_336,In_1703,In_3);
or U337 (N_337,In_711,In_1462);
nand U338 (N_338,In_1480,In_1963);
nor U339 (N_339,In_1710,In_1285);
nor U340 (N_340,In_1969,In_444);
nor U341 (N_341,In_290,In_1006);
nor U342 (N_342,In_603,In_510);
or U343 (N_343,In_80,In_1444);
nand U344 (N_344,In_1315,In_528);
nor U345 (N_345,In_1855,In_389);
nand U346 (N_346,In_394,In_154);
and U347 (N_347,In_911,In_1020);
or U348 (N_348,In_374,In_54);
nor U349 (N_349,In_1679,In_714);
xnor U350 (N_350,In_1384,In_1471);
or U351 (N_351,In_727,In_15);
nand U352 (N_352,In_935,In_1982);
nand U353 (N_353,In_625,In_28);
and U354 (N_354,In_34,In_1210);
and U355 (N_355,In_786,In_664);
or U356 (N_356,In_756,In_485);
and U357 (N_357,In_1863,In_1066);
xor U358 (N_358,In_278,In_1252);
nor U359 (N_359,In_1606,In_1597);
nand U360 (N_360,In_1651,In_340);
nand U361 (N_361,In_217,In_469);
and U362 (N_362,In_518,In_23);
and U363 (N_363,In_1802,In_1815);
xor U364 (N_364,In_677,In_238);
nor U365 (N_365,In_291,In_1316);
or U366 (N_366,In_1305,In_769);
and U367 (N_367,In_1441,In_1500);
nand U368 (N_368,In_1225,In_1879);
and U369 (N_369,In_806,In_876);
or U370 (N_370,In_1023,In_169);
xor U371 (N_371,In_1450,In_706);
and U372 (N_372,In_1399,In_1427);
or U373 (N_373,In_897,In_1811);
xor U374 (N_374,In_1436,In_1395);
and U375 (N_375,In_1186,In_1786);
or U376 (N_376,In_1124,In_483);
and U377 (N_377,In_1831,In_270);
and U378 (N_378,In_1483,In_1869);
xnor U379 (N_379,In_1492,In_1909);
nand U380 (N_380,In_933,In_1957);
nor U381 (N_381,In_1540,In_1833);
nand U382 (N_382,In_871,In_744);
nor U383 (N_383,In_1844,In_494);
or U384 (N_384,In_722,In_1050);
nor U385 (N_385,In_1534,In_1335);
or U386 (N_386,In_1358,In_592);
nand U387 (N_387,In_1288,In_1236);
nand U388 (N_388,In_576,In_803);
nor U389 (N_389,In_811,In_1039);
and U390 (N_390,In_1158,In_165);
nor U391 (N_391,In_1094,In_691);
or U392 (N_392,In_1292,In_1852);
nand U393 (N_393,In_641,In_107);
nor U394 (N_394,In_1686,In_148);
xnor U395 (N_395,In_72,In_1470);
nand U396 (N_396,In_296,In_1777);
and U397 (N_397,In_38,In_372);
or U398 (N_398,In_289,In_809);
xor U399 (N_399,In_1888,In_1241);
or U400 (N_400,In_1481,In_1119);
and U401 (N_401,In_1495,In_1976);
and U402 (N_402,In_1537,In_998);
nor U403 (N_403,In_1914,In_373);
and U404 (N_404,In_67,In_985);
nand U405 (N_405,In_932,In_1370);
nor U406 (N_406,In_1564,In_59);
nand U407 (N_407,In_1231,In_726);
or U408 (N_408,In_1417,In_1814);
xnor U409 (N_409,In_1189,In_1774);
and U410 (N_410,In_982,In_1837);
nor U411 (N_411,In_798,In_492);
or U412 (N_412,In_939,In_357);
nand U413 (N_413,In_1989,In_1223);
and U414 (N_414,In_749,In_1404);
nor U415 (N_415,In_797,In_1040);
nand U416 (N_416,In_180,In_1861);
nand U417 (N_417,In_1127,In_1341);
or U418 (N_418,In_1188,In_913);
and U419 (N_419,In_787,In_1375);
and U420 (N_420,In_1080,In_447);
nand U421 (N_421,In_1932,In_1631);
xor U422 (N_422,In_810,In_361);
nor U423 (N_423,In_1938,In_1582);
xnor U424 (N_424,In_728,In_942);
and U425 (N_425,In_55,In_532);
xor U426 (N_426,In_526,In_1499);
nand U427 (N_427,In_158,In_1074);
nand U428 (N_428,In_1900,In_136);
nor U429 (N_429,In_1311,In_523);
and U430 (N_430,In_1804,In_1864);
nor U431 (N_431,In_563,In_747);
or U432 (N_432,In_343,In_1149);
or U433 (N_433,In_650,In_1515);
xor U434 (N_434,In_253,In_1830);
or U435 (N_435,In_75,In_701);
xnor U436 (N_436,In_1381,In_1221);
nor U437 (N_437,In_1466,In_1729);
nor U438 (N_438,In_934,In_266);
nor U439 (N_439,In_1954,In_1173);
nand U440 (N_440,In_538,In_229);
nand U441 (N_441,In_279,In_683);
or U442 (N_442,In_921,In_1437);
or U443 (N_443,In_1876,In_1652);
xor U444 (N_444,In_1663,In_789);
nand U445 (N_445,In_1649,In_1102);
and U446 (N_446,In_44,In_1166);
xor U447 (N_447,In_622,In_554);
nor U448 (N_448,In_1169,In_1485);
nor U449 (N_449,In_1657,In_1965);
xor U450 (N_450,In_1769,In_1264);
nand U451 (N_451,In_388,In_479);
or U452 (N_452,In_1516,In_105);
and U453 (N_453,In_1827,In_675);
xnor U454 (N_454,In_1560,In_901);
nand U455 (N_455,In_1388,In_1899);
and U456 (N_456,In_1504,In_327);
and U457 (N_457,In_130,In_408);
and U458 (N_458,In_1156,In_1307);
nor U459 (N_459,In_1131,In_896);
nor U460 (N_460,In_595,In_994);
nand U461 (N_461,In_1715,In_417);
and U462 (N_462,In_1822,In_1112);
nor U463 (N_463,In_1974,In_1853);
or U464 (N_464,In_663,In_1037);
or U465 (N_465,In_1733,In_852);
xor U466 (N_466,In_1889,In_1887);
and U467 (N_467,In_1253,In_76);
and U468 (N_468,In_1171,In_654);
nand U469 (N_469,In_1132,In_1881);
or U470 (N_470,In_427,In_1916);
or U471 (N_471,In_1036,In_1927);
or U472 (N_472,In_475,In_240);
or U473 (N_473,In_1995,In_1246);
nand U474 (N_474,In_910,In_1029);
and U475 (N_475,In_858,In_0);
or U476 (N_476,In_160,In_1237);
nand U477 (N_477,In_1320,In_559);
or U478 (N_478,In_1085,In_1543);
and U479 (N_479,In_1146,In_1016);
nor U480 (N_480,In_433,In_1812);
or U481 (N_481,In_342,In_1258);
and U482 (N_482,In_458,In_1270);
nor U483 (N_483,In_1936,In_793);
nor U484 (N_484,In_64,In_1588);
or U485 (N_485,In_740,In_1199);
nand U486 (N_486,In_1882,In_585);
nor U487 (N_487,In_330,In_1458);
or U488 (N_488,In_863,In_1278);
and U489 (N_489,In_681,In_431);
or U490 (N_490,In_892,In_600);
xor U491 (N_491,In_1695,In_57);
or U492 (N_492,In_678,In_1654);
or U493 (N_493,In_1994,In_1374);
and U494 (N_494,In_1648,In_953);
or U495 (N_495,In_277,In_119);
nor U496 (N_496,In_1896,In_98);
and U497 (N_497,In_785,In_434);
xor U498 (N_498,In_1088,In_1009);
and U499 (N_499,In_323,In_643);
and U500 (N_500,In_605,In_370);
nor U501 (N_501,In_1420,In_735);
and U502 (N_502,In_1351,In_1566);
xor U503 (N_503,In_1142,In_347);
nor U504 (N_504,In_671,In_940);
or U505 (N_505,In_1125,In_1287);
xnor U506 (N_506,In_153,In_1958);
or U507 (N_507,In_990,In_1803);
xnor U508 (N_508,In_698,In_1072);
and U509 (N_509,In_213,In_1473);
or U510 (N_510,In_560,In_1206);
nand U511 (N_511,In_7,In_767);
nand U512 (N_512,In_1185,In_849);
nand U513 (N_513,In_1139,In_1177);
nor U514 (N_514,In_146,In_1349);
or U515 (N_515,In_781,In_1545);
nor U516 (N_516,In_1003,In_16);
xor U517 (N_517,In_1422,In_1552);
or U518 (N_518,In_170,In_60);
xor U519 (N_519,In_504,In_1810);
nand U520 (N_520,In_1302,In_1202);
xor U521 (N_521,In_1194,In_1823);
or U522 (N_522,In_672,In_899);
and U523 (N_523,In_973,In_1556);
xor U524 (N_524,In_1180,In_1743);
nor U525 (N_525,In_1908,In_1118);
xor U526 (N_526,In_261,In_903);
nor U527 (N_527,In_979,In_674);
and U528 (N_528,In_328,In_862);
and U529 (N_529,In_21,In_1570);
nand U530 (N_530,In_1394,In_1633);
nor U531 (N_531,In_1975,In_1268);
nand U532 (N_532,In_784,In_215);
xnor U533 (N_533,In_1738,In_1111);
or U534 (N_534,In_1642,In_1027);
nand U535 (N_535,In_1839,In_1608);
xor U536 (N_536,In_1949,In_1801);
nand U537 (N_537,In_156,In_1639);
nand U538 (N_538,In_1048,In_1431);
and U539 (N_539,In_142,In_46);
or U540 (N_540,In_1628,In_624);
or U541 (N_541,In_1558,In_1001);
xnor U542 (N_542,In_584,In_1867);
and U543 (N_543,In_867,In_351);
xor U544 (N_544,In_723,In_964);
nand U545 (N_545,In_1992,In_189);
or U546 (N_546,In_651,In_1086);
and U547 (N_547,In_558,In_14);
nand U548 (N_548,In_399,In_929);
and U549 (N_549,In_308,In_45);
nand U550 (N_550,In_1018,In_513);
nor U551 (N_551,In_86,In_1635);
nor U552 (N_552,In_106,In_923);
nor U553 (N_553,In_1266,In_432);
xor U554 (N_554,In_495,In_1393);
nor U555 (N_555,In_552,In_1719);
nor U556 (N_556,In_8,In_111);
nor U557 (N_557,In_1416,In_887);
nand U558 (N_558,In_1713,In_1138);
and U559 (N_559,In_1297,In_298);
xnor U560 (N_560,In_1990,In_1590);
or U561 (N_561,In_286,In_1660);
xnor U562 (N_562,In_207,In_1157);
nand U563 (N_563,In_1970,In_422);
nand U564 (N_564,In_218,In_267);
xor U565 (N_565,In_58,In_314);
nor U566 (N_566,In_301,In_690);
and U567 (N_567,In_1689,In_423);
nand U568 (N_568,In_1294,In_430);
nor U569 (N_569,In_96,In_1062);
xor U570 (N_570,In_693,In_1836);
xor U571 (N_571,In_1661,In_338);
and U572 (N_572,In_1704,In_26);
nand U573 (N_573,In_1147,In_734);
nand U574 (N_574,In_1213,In_1077);
or U575 (N_575,In_1693,In_415);
xor U576 (N_576,In_1281,In_352);
xor U577 (N_577,In_537,In_1650);
xnor U578 (N_578,In_101,In_615);
and U579 (N_579,In_99,In_1415);
nand U580 (N_580,In_1687,In_1615);
or U581 (N_581,In_1541,In_900);
nor U582 (N_582,In_181,In_516);
nor U583 (N_583,In_1848,In_1536);
nand U584 (N_584,In_89,In_285);
nand U585 (N_585,In_1339,In_995);
and U586 (N_586,In_1671,In_1082);
and U587 (N_587,In_135,In_796);
xor U588 (N_588,In_1653,In_1562);
or U589 (N_589,In_832,In_209);
xor U590 (N_590,In_1198,In_715);
nand U591 (N_591,In_452,In_1796);
nand U592 (N_592,In_952,In_1347);
and U593 (N_593,In_1764,In_549);
nand U594 (N_594,In_1486,In_889);
xor U595 (N_595,In_847,In_1937);
nor U596 (N_596,In_333,In_1800);
nand U597 (N_597,In_1323,In_241);
and U598 (N_598,In_1551,In_524);
xnor U599 (N_599,In_489,In_1776);
nand U600 (N_600,In_386,In_1360);
nand U601 (N_601,In_1134,In_204);
xor U602 (N_602,In_1274,In_1357);
or U603 (N_603,In_878,In_132);
nor U604 (N_604,In_1133,In_297);
xor U605 (N_605,In_667,In_1245);
and U606 (N_606,In_628,In_1573);
and U607 (N_607,In_721,In_668);
and U608 (N_608,In_1267,In_894);
nor U609 (N_609,In_1567,In_1667);
nand U610 (N_610,In_1708,In_1379);
nand U611 (N_611,In_1,In_254);
nand U612 (N_612,In_802,In_319);
and U613 (N_613,In_186,In_709);
and U614 (N_614,In_1659,In_1665);
nor U615 (N_615,In_1120,In_1113);
or U616 (N_616,In_1410,In_1923);
or U617 (N_617,In_1532,In_1081);
nand U618 (N_618,In_1319,In_251);
and U619 (N_619,In_777,In_666);
xor U620 (N_620,In_1256,In_616);
nand U621 (N_621,In_1850,In_1463);
nand U622 (N_622,In_1068,In_684);
nor U623 (N_623,In_1883,In_1069);
xor U624 (N_624,In_1309,In_1366);
and U625 (N_625,In_397,In_505);
or U626 (N_626,In_729,In_436);
and U627 (N_627,In_1161,In_1625);
xnor U628 (N_628,In_653,In_164);
and U629 (N_629,In_1718,In_577);
and U630 (N_630,In_1153,In_1817);
nand U631 (N_631,In_198,In_2);
nor U632 (N_632,In_1681,In_117);
nand U633 (N_633,In_1948,In_1448);
nor U634 (N_634,In_269,In_1550);
nand U635 (N_635,In_476,In_1791);
nand U636 (N_636,In_1364,In_669);
or U637 (N_637,In_477,In_738);
nand U638 (N_638,In_1129,In_1721);
nor U639 (N_639,In_1296,In_1673);
or U640 (N_640,In_499,In_1851);
or U641 (N_641,In_1181,In_636);
xor U642 (N_642,In_997,In_1600);
and U643 (N_643,In_1402,In_1736);
nand U644 (N_644,In_1798,In_805);
and U645 (N_645,In_1122,In_1126);
or U646 (N_646,In_1749,In_1712);
nand U647 (N_647,In_550,In_1136);
xnor U648 (N_648,In_454,In_1961);
nor U649 (N_649,In_1411,In_1353);
nor U650 (N_650,In_1265,In_742);
nor U651 (N_651,In_1105,In_1846);
xor U652 (N_652,In_578,In_1440);
xnor U653 (N_653,In_120,In_1955);
and U654 (N_654,In_838,In_56);
xnor U655 (N_655,In_1140,In_1619);
xor U656 (N_656,In_1107,In_993);
and U657 (N_657,In_704,In_916);
xnor U658 (N_658,In_10,In_24);
or U659 (N_659,In_1079,In_1196);
nor U660 (N_660,In_1217,In_975);
nand U661 (N_661,In_1991,In_1555);
or U662 (N_662,In_410,In_1576);
nor U663 (N_663,In_1392,In_1985);
or U664 (N_664,In_295,In_1700);
or U665 (N_665,In_1616,In_1981);
xnor U666 (N_666,In_234,In_1454);
nor U667 (N_667,In_978,In_1168);
nor U668 (N_668,In_40,In_1640);
nand U669 (N_669,In_1414,In_294);
xnor U670 (N_670,In_588,In_414);
nor U671 (N_671,In_482,In_909);
nor U672 (N_672,In_276,In_1459);
nor U673 (N_673,In_529,In_1931);
or U674 (N_674,In_1858,In_51);
nor U675 (N_675,In_1874,In_1685);
and U676 (N_676,In_502,In_1451);
nor U677 (N_677,In_497,In_1461);
or U678 (N_678,In_1971,In_1701);
and U679 (N_679,In_1664,In_1164);
or U680 (N_680,In_246,In_1222);
or U681 (N_681,In_334,In_1768);
or U682 (N_682,In_1488,In_66);
or U683 (N_683,In_612,In_960);
nand U684 (N_684,In_963,In_1676);
xnor U685 (N_685,In_409,In_403);
nand U686 (N_686,In_1271,In_194);
nor U687 (N_687,In_1694,In_459);
or U688 (N_688,In_686,In_1045);
nor U689 (N_689,In_126,In_886);
or U690 (N_690,In_619,In_1367);
xor U691 (N_691,In_100,In_1313);
and U692 (N_692,In_88,In_1389);
xor U693 (N_693,In_788,In_757);
nor U694 (N_694,In_1244,In_50);
nor U695 (N_695,In_676,In_764);
and U696 (N_696,In_1586,In_1821);
nand U697 (N_697,In_1720,In_249);
or U698 (N_698,In_1725,In_1589);
or U699 (N_699,In_1363,In_1418);
nand U700 (N_700,In_883,In_1008);
nor U701 (N_701,In_488,In_1528);
nor U702 (N_702,In_635,In_1148);
nor U703 (N_703,In_718,In_82);
xor U704 (N_704,In_856,In_779);
xor U705 (N_705,In_1618,In_601);
nor U706 (N_706,In_22,In_398);
or U707 (N_707,In_947,In_1530);
nand U708 (N_708,In_954,In_1943);
nand U709 (N_709,In_1183,In_131);
and U710 (N_710,In_1726,In_1630);
xnor U711 (N_711,In_840,In_1531);
and U712 (N_712,In_300,In_1429);
and U713 (N_713,In_1779,In_1043);
xnor U714 (N_714,In_844,In_884);
nand U715 (N_715,In_870,In_1075);
and U716 (N_716,In_800,In_1727);
xor U717 (N_717,In_739,In_1078);
and U718 (N_718,In_41,In_1684);
or U719 (N_719,In_1476,In_970);
and U720 (N_720,In_1432,In_557);
and U721 (N_721,In_1613,In_1092);
and U722 (N_722,In_115,In_594);
nor U723 (N_723,In_1408,In_1121);
xor U724 (N_724,In_533,In_134);
xnor U725 (N_725,In_481,In_1496);
nor U726 (N_726,In_446,In_1674);
xor U727 (N_727,In_1561,In_1096);
and U728 (N_728,In_989,In_1322);
nand U729 (N_729,In_1250,In_759);
or U730 (N_730,In_303,In_925);
or U731 (N_731,In_1877,In_1893);
nor U732 (N_732,In_1338,In_1063);
nand U733 (N_733,In_956,In_1682);
nand U734 (N_734,In_1214,In_237);
xor U735 (N_735,In_329,In_70);
nor U736 (N_736,In_1455,In_1577);
nor U737 (N_737,In_991,In_1917);
nand U738 (N_738,In_1403,In_579);
xnor U739 (N_739,In_302,In_496);
nand U740 (N_740,In_1872,In_84);
or U741 (N_741,In_1716,In_1523);
and U742 (N_742,In_1824,In_517);
nor U743 (N_743,In_1692,In_572);
nor U744 (N_744,In_1260,In_983);
xor U745 (N_745,In_976,In_912);
and U746 (N_746,In_1752,In_1469);
and U747 (N_747,In_872,In_799);
nand U748 (N_748,In_30,In_1728);
nand U749 (N_749,In_732,In_792);
and U750 (N_750,In_1215,In_1939);
xor U751 (N_751,In_348,In_531);
xor U752 (N_752,In_1220,In_525);
nand U753 (N_753,In_1355,In_1103);
and U754 (N_754,In_1765,In_383);
nand U755 (N_755,In_124,In_1178);
nor U756 (N_756,In_546,In_689);
nor U757 (N_757,In_1117,In_950);
nand U758 (N_758,In_1058,In_1807);
or U759 (N_759,In_658,In_243);
nand U760 (N_760,In_710,In_1688);
or U761 (N_761,In_645,In_791);
xor U762 (N_762,In_697,In_621);
xor U763 (N_763,In_1913,In_626);
nand U764 (N_764,In_1714,In_1782);
nor U765 (N_765,In_1152,In_1781);
and U766 (N_766,In_1170,In_203);
xnor U767 (N_767,In_1084,In_1945);
xnor U768 (N_768,In_1282,In_1601);
nor U769 (N_769,In_1929,In_1336);
and U770 (N_770,In_1978,In_149);
and U771 (N_771,In_443,In_1526);
xor U772 (N_772,In_1902,In_1308);
nand U773 (N_773,In_656,In_200);
or U774 (N_774,In_362,In_197);
xor U775 (N_775,In_1638,In_647);
nand U776 (N_776,In_1091,In_324);
and U777 (N_777,In_487,In_133);
nor U778 (N_778,In_609,In_527);
nor U779 (N_779,In_1737,In_387);
nand U780 (N_780,In_1730,In_1522);
xnor U781 (N_781,In_971,In_1159);
nand U782 (N_782,In_1603,In_260);
and U783 (N_783,In_116,In_829);
nor U784 (N_784,In_1123,In_568);
or U785 (N_785,In_503,In_1110);
xnor U786 (N_786,In_440,In_1950);
or U787 (N_787,In_1160,In_1617);
and U788 (N_788,In_1044,In_536);
nor U789 (N_789,In_1197,In_1035);
and U790 (N_790,In_363,In_922);
or U791 (N_791,In_121,In_1087);
and U792 (N_792,In_78,In_879);
or U793 (N_793,In_462,In_1344);
nand U794 (N_794,In_49,In_118);
nand U795 (N_795,In_1295,In_167);
or U796 (N_796,In_304,In_33);
nor U797 (N_797,In_1626,In_758);
xnor U798 (N_798,In_1406,In_860);
xnor U799 (N_799,In_1951,In_123);
nor U800 (N_800,In_541,In_1997);
xnor U801 (N_801,In_252,In_155);
and U802 (N_802,In_1234,In_843);
nor U803 (N_803,In_825,In_455);
xnor U804 (N_804,In_206,In_1742);
and U805 (N_805,In_1507,In_1538);
or U806 (N_806,In_827,In_733);
nor U807 (N_807,In_1873,In_833);
nand U808 (N_808,In_737,In_1371);
xnor U809 (N_809,In_484,In_113);
and U810 (N_810,In_507,In_1372);
nor U811 (N_811,In_1073,In_812);
nor U812 (N_812,In_1251,In_1609);
nor U813 (N_813,In_1030,In_1090);
or U814 (N_814,In_1135,In_720);
or U815 (N_815,In_257,In_670);
nor U816 (N_816,In_1368,In_1425);
nand U817 (N_817,In_941,In_627);
or U818 (N_818,In_1795,In_1011);
nor U819 (N_819,In_1842,In_875);
and U820 (N_820,In_1047,In_1224);
nor U821 (N_821,In_1497,In_1227);
nand U822 (N_822,In_1611,In_1361);
and U823 (N_823,In_561,In_765);
and U824 (N_824,In_162,In_299);
nand U825 (N_825,In_226,In_1620);
xor U826 (N_826,In_1059,In_946);
nor U827 (N_827,In_1052,In_562);
xor U828 (N_828,In_202,In_391);
nor U829 (N_829,In_1697,In_814);
nand U830 (N_830,In_713,In_1533);
or U831 (N_831,In_193,In_220);
nor U832 (N_832,In_1717,In_214);
xor U833 (N_833,In_1430,In_1304);
or U834 (N_834,In_637,In_104);
and U835 (N_835,In_265,In_349);
or U836 (N_836,In_493,In_545);
nor U837 (N_837,In_1751,In_782);
and U838 (N_838,In_322,In_168);
nand U839 (N_839,In_614,In_1906);
and U840 (N_840,In_1553,In_1192);
nand U841 (N_841,In_426,In_61);
nor U842 (N_842,In_1988,In_468);
xor U843 (N_843,In_184,In_137);
xnor U844 (N_844,In_1332,In_453);
or U845 (N_845,In_1303,In_331);
xor U846 (N_846,In_1130,In_1482);
and U847 (N_847,In_1575,In_762);
and U848 (N_848,In_371,In_596);
or U849 (N_849,In_1809,In_1015);
and U850 (N_850,In_1592,In_157);
or U851 (N_851,In_1521,In_521);
xnor U852 (N_852,In_29,In_1273);
or U853 (N_853,In_930,In_680);
xor U854 (N_854,In_575,In_5);
nand U855 (N_855,In_1300,In_1240);
nand U856 (N_856,In_140,In_783);
nor U857 (N_857,In_555,In_1643);
and U858 (N_858,In_274,In_354);
nor U859 (N_859,In_491,In_350);
xnor U860 (N_860,In_1793,In_692);
nand U861 (N_861,In_657,In_281);
or U862 (N_862,In_192,In_1326);
xor U863 (N_863,In_1070,In_1805);
nand U864 (N_864,In_1599,In_109);
nand U865 (N_865,In_606,In_221);
nor U866 (N_866,In_859,In_1280);
or U867 (N_867,In_1434,In_1539);
xnor U868 (N_868,In_466,In_639);
nor U869 (N_869,In_1446,In_1329);
xor U870 (N_870,In_1723,In_866);
nor U871 (N_871,In_1219,In_801);
or U872 (N_872,In_1792,In_1490);
and U873 (N_873,In_556,In_766);
xnor U874 (N_874,In_1542,In_652);
nand U875 (N_875,In_1299,In_1897);
or U876 (N_876,In_1421,In_644);
nor U877 (N_877,In_700,In_1327);
and U878 (N_878,In_233,In_1890);
nor U879 (N_879,In_1479,In_1875);
xor U880 (N_880,In_43,In_1935);
or U881 (N_881,In_195,In_1818);
xnor U882 (N_882,In_9,In_87);
nor U883 (N_883,In_1825,In_1983);
nor U884 (N_884,In_881,In_230);
nand U885 (N_885,In_36,In_1255);
nor U886 (N_886,In_819,In_1636);
nor U887 (N_887,In_1275,In_1775);
nand U888 (N_888,In_1407,In_848);
nor U889 (N_889,In_530,In_682);
xnor U890 (N_890,In_1862,In_1021);
or U891 (N_891,In_955,In_1340);
nor U892 (N_892,In_1491,In_31);
xor U893 (N_893,In_1826,In_1314);
xnor U894 (N_894,In_196,In_199);
xor U895 (N_895,In_1276,In_311);
nand U896 (N_896,In_1365,In_1019);
nand U897 (N_897,In_255,In_97);
or U898 (N_898,In_1071,In_92);
and U899 (N_899,In_1026,In_1350);
nor U900 (N_900,In_597,In_823);
nor U901 (N_901,In_250,In_772);
or U902 (N_902,In_1097,In_1205);
or U903 (N_903,In_1563,In_746);
and U904 (N_904,In_125,In_1195);
and U905 (N_905,In_927,In_1229);
nor U906 (N_906,In_1354,In_1878);
nand U907 (N_907,In_1904,In_836);
nand U908 (N_908,In_1946,In_634);
nor U909 (N_909,In_1525,In_638);
nand U910 (N_910,In_857,In_1212);
xnor U911 (N_911,In_1200,In_1104);
nand U912 (N_912,In_1744,In_102);
and U913 (N_913,In_1740,In_248);
nor U914 (N_914,In_1289,In_32);
nor U915 (N_915,In_1290,In_1369);
or U916 (N_916,In_1291,In_571);
xnor U917 (N_917,In_904,In_763);
xnor U918 (N_918,In_1114,In_367);
nor U919 (N_919,In_662,In_1163);
and U920 (N_920,In_1057,In_1306);
or U921 (N_921,In_1891,In_845);
nor U922 (N_922,In_1783,In_1099);
or U923 (N_923,In_1773,In_753);
nand U924 (N_924,In_1568,In_359);
or U925 (N_925,In_1731,In_968);
nand U926 (N_926,In_1046,In_282);
and U927 (N_927,In_877,In_905);
and U928 (N_928,In_1746,In_1547);
and U929 (N_929,In_566,In_1498);
and U930 (N_930,In_992,In_1672);
nand U931 (N_931,In_20,In_1645);
xnor U932 (N_932,In_1702,In_1012);
xnor U933 (N_933,In_463,In_1813);
or U934 (N_934,In_620,In_211);
and U935 (N_935,In_717,In_360);
nor U936 (N_936,In_1128,In_1706);
and U937 (N_937,In_390,In_312);
or U938 (N_938,In_1919,In_926);
and U939 (N_939,In_179,In_143);
nand U940 (N_940,In_412,In_1578);
and U941 (N_941,In_687,In_244);
or U942 (N_942,In_1373,In_1279);
and U943 (N_943,In_1646,In_1797);
nor U944 (N_944,In_1980,In_1038);
nor U945 (N_945,In_1641,In_382);
or U946 (N_946,In_395,In_159);
nand U947 (N_947,In_1780,In_824);
or U948 (N_948,In_411,In_986);
nor U949 (N_949,In_1155,In_256);
and U950 (N_950,In_307,In_375);
nand U951 (N_951,In_1413,In_1761);
or U952 (N_952,In_421,In_1051);
nor U953 (N_953,In_425,In_1905);
nand U954 (N_954,In_245,In_1014);
xor U955 (N_955,In_420,In_1010);
xnor U956 (N_956,In_618,In_1460);
and U957 (N_957,In_500,In_1838);
nand U958 (N_958,In_402,In_400);
nor U959 (N_959,In_1845,In_364);
nor U960 (N_960,In_401,In_242);
or U961 (N_961,In_473,In_407);
and U962 (N_962,In_969,In_1579);
and U963 (N_963,In_336,In_917);
nor U964 (N_964,In_1548,In_854);
and U965 (N_965,In_974,In_317);
and U966 (N_966,In_581,In_547);
and U967 (N_967,In_1512,In_660);
nor U968 (N_968,In_139,In_1400);
or U969 (N_969,In_368,In_1137);
nor U970 (N_970,In_448,In_1487);
nand U971 (N_971,In_451,In_1447);
and U972 (N_972,In_1013,In_288);
nor U973 (N_973,In_1766,In_1144);
nor U974 (N_974,In_752,In_1920);
nand U975 (N_975,In_1593,In_816);
nor U976 (N_976,In_598,In_841);
nand U977 (N_977,In_898,In_750);
or U978 (N_978,In_1503,In_1017);
nor U979 (N_979,In_1964,In_1193);
nand U980 (N_980,In_1317,In_1257);
nand U981 (N_981,In_172,In_1584);
xnor U982 (N_982,In_1947,In_1510);
or U983 (N_983,In_1191,In_1595);
nand U984 (N_984,In_1143,In_353);
or U985 (N_985,In_1709,In_1506);
nor U986 (N_986,In_1886,In_341);
nand U987 (N_987,In_1478,In_396);
nor U988 (N_988,In_1269,In_1108);
nand U989 (N_989,In_790,In_1386);
xnor U990 (N_990,In_416,In_972);
nor U991 (N_991,In_1259,In_1722);
xor U992 (N_992,In_830,In_1150);
or U993 (N_993,In_1535,In_474);
or U994 (N_994,In_4,In_1390);
or U995 (N_995,In_895,In_807);
and U996 (N_996,In_465,In_1621);
xor U997 (N_997,In_385,In_344);
nand U998 (N_998,In_1301,In_1468);
nand U999 (N_999,In_1565,In_1745);
or U1000 (N_1000,In_1884,In_1787);
and U1001 (N_1001,In_1086,In_699);
xnor U1002 (N_1002,In_662,In_767);
nor U1003 (N_1003,In_200,In_1073);
nand U1004 (N_1004,In_1957,In_1792);
or U1005 (N_1005,In_1648,In_1460);
nor U1006 (N_1006,In_962,In_934);
xnor U1007 (N_1007,In_901,In_1448);
nand U1008 (N_1008,In_903,In_1878);
nand U1009 (N_1009,In_206,In_1325);
xor U1010 (N_1010,In_151,In_1517);
and U1011 (N_1011,In_226,In_737);
and U1012 (N_1012,In_1024,In_1717);
nand U1013 (N_1013,In_1164,In_892);
or U1014 (N_1014,In_860,In_1578);
nand U1015 (N_1015,In_644,In_319);
nor U1016 (N_1016,In_1924,In_1025);
nand U1017 (N_1017,In_1705,In_1145);
and U1018 (N_1018,In_1179,In_590);
or U1019 (N_1019,In_94,In_139);
nand U1020 (N_1020,In_874,In_1669);
or U1021 (N_1021,In_356,In_637);
and U1022 (N_1022,In_1697,In_419);
or U1023 (N_1023,In_1339,In_458);
or U1024 (N_1024,In_1721,In_1958);
nor U1025 (N_1025,In_1193,In_913);
xnor U1026 (N_1026,In_1621,In_1116);
and U1027 (N_1027,In_663,In_269);
and U1028 (N_1028,In_852,In_939);
and U1029 (N_1029,In_1894,In_543);
and U1030 (N_1030,In_1156,In_1934);
nor U1031 (N_1031,In_166,In_1237);
nor U1032 (N_1032,In_1575,In_1597);
nand U1033 (N_1033,In_1874,In_696);
xnor U1034 (N_1034,In_1996,In_885);
nand U1035 (N_1035,In_1659,In_1958);
xor U1036 (N_1036,In_711,In_272);
nand U1037 (N_1037,In_1725,In_1782);
and U1038 (N_1038,In_1131,In_482);
nor U1039 (N_1039,In_1909,In_200);
xnor U1040 (N_1040,In_648,In_1553);
nand U1041 (N_1041,In_584,In_384);
and U1042 (N_1042,In_1506,In_1548);
and U1043 (N_1043,In_1110,In_446);
and U1044 (N_1044,In_1199,In_1776);
nor U1045 (N_1045,In_260,In_701);
and U1046 (N_1046,In_657,In_56);
xor U1047 (N_1047,In_633,In_1900);
and U1048 (N_1048,In_348,In_1535);
nand U1049 (N_1049,In_1170,In_1520);
or U1050 (N_1050,In_1122,In_152);
xnor U1051 (N_1051,In_719,In_773);
xnor U1052 (N_1052,In_158,In_668);
nand U1053 (N_1053,In_1312,In_832);
nand U1054 (N_1054,In_549,In_537);
and U1055 (N_1055,In_734,In_1747);
nor U1056 (N_1056,In_579,In_1340);
nor U1057 (N_1057,In_1513,In_1312);
nor U1058 (N_1058,In_908,In_942);
and U1059 (N_1059,In_1691,In_1382);
nor U1060 (N_1060,In_26,In_1428);
and U1061 (N_1061,In_720,In_672);
and U1062 (N_1062,In_1538,In_88);
and U1063 (N_1063,In_1204,In_900);
and U1064 (N_1064,In_962,In_1812);
xnor U1065 (N_1065,In_1522,In_1638);
and U1066 (N_1066,In_1968,In_439);
nand U1067 (N_1067,In_69,In_613);
nor U1068 (N_1068,In_814,In_395);
and U1069 (N_1069,In_1292,In_945);
or U1070 (N_1070,In_1769,In_895);
nor U1071 (N_1071,In_1949,In_776);
nand U1072 (N_1072,In_396,In_1275);
nand U1073 (N_1073,In_1792,In_835);
or U1074 (N_1074,In_553,In_910);
nor U1075 (N_1075,In_586,In_243);
and U1076 (N_1076,In_279,In_1116);
and U1077 (N_1077,In_937,In_745);
nand U1078 (N_1078,In_212,In_1262);
or U1079 (N_1079,In_1070,In_1086);
and U1080 (N_1080,In_330,In_1766);
nand U1081 (N_1081,In_1396,In_703);
or U1082 (N_1082,In_1381,In_884);
xor U1083 (N_1083,In_264,In_1157);
nand U1084 (N_1084,In_457,In_1178);
xnor U1085 (N_1085,In_1145,In_377);
and U1086 (N_1086,In_1006,In_1971);
xor U1087 (N_1087,In_415,In_264);
nor U1088 (N_1088,In_1349,In_1837);
or U1089 (N_1089,In_326,In_1656);
or U1090 (N_1090,In_901,In_1386);
nor U1091 (N_1091,In_833,In_292);
nand U1092 (N_1092,In_1932,In_1900);
nor U1093 (N_1093,In_1687,In_195);
and U1094 (N_1094,In_915,In_216);
or U1095 (N_1095,In_1652,In_1340);
or U1096 (N_1096,In_1980,In_82);
nand U1097 (N_1097,In_1195,In_543);
or U1098 (N_1098,In_368,In_374);
xnor U1099 (N_1099,In_711,In_657);
nand U1100 (N_1100,In_1464,In_1899);
and U1101 (N_1101,In_476,In_373);
nand U1102 (N_1102,In_254,In_1598);
xor U1103 (N_1103,In_281,In_1674);
nor U1104 (N_1104,In_1210,In_354);
and U1105 (N_1105,In_1157,In_61);
nand U1106 (N_1106,In_1497,In_734);
and U1107 (N_1107,In_1078,In_63);
nor U1108 (N_1108,In_107,In_1346);
and U1109 (N_1109,In_1218,In_1306);
nand U1110 (N_1110,In_805,In_309);
nand U1111 (N_1111,In_1936,In_326);
xor U1112 (N_1112,In_905,In_1221);
nand U1113 (N_1113,In_1513,In_1078);
xor U1114 (N_1114,In_152,In_188);
nand U1115 (N_1115,In_1210,In_1932);
nand U1116 (N_1116,In_807,In_1890);
nand U1117 (N_1117,In_14,In_1454);
xor U1118 (N_1118,In_1390,In_1030);
xnor U1119 (N_1119,In_1793,In_816);
nor U1120 (N_1120,In_1979,In_204);
and U1121 (N_1121,In_134,In_641);
and U1122 (N_1122,In_511,In_634);
nand U1123 (N_1123,In_1021,In_93);
xor U1124 (N_1124,In_1996,In_840);
or U1125 (N_1125,In_352,In_722);
xnor U1126 (N_1126,In_597,In_178);
or U1127 (N_1127,In_877,In_1326);
nor U1128 (N_1128,In_237,In_515);
and U1129 (N_1129,In_986,In_1093);
nand U1130 (N_1130,In_814,In_410);
nand U1131 (N_1131,In_956,In_1109);
nor U1132 (N_1132,In_823,In_1559);
nor U1133 (N_1133,In_1577,In_1274);
and U1134 (N_1134,In_1856,In_246);
xor U1135 (N_1135,In_1464,In_501);
nand U1136 (N_1136,In_1698,In_986);
nand U1137 (N_1137,In_786,In_936);
xnor U1138 (N_1138,In_1981,In_517);
xnor U1139 (N_1139,In_534,In_208);
xor U1140 (N_1140,In_91,In_142);
nand U1141 (N_1141,In_1247,In_376);
xnor U1142 (N_1142,In_1672,In_681);
nor U1143 (N_1143,In_193,In_209);
nor U1144 (N_1144,In_1041,In_789);
and U1145 (N_1145,In_1522,In_1727);
nand U1146 (N_1146,In_1928,In_969);
and U1147 (N_1147,In_1934,In_764);
and U1148 (N_1148,In_587,In_1907);
xnor U1149 (N_1149,In_1032,In_1948);
nor U1150 (N_1150,In_1444,In_300);
and U1151 (N_1151,In_1034,In_470);
nor U1152 (N_1152,In_344,In_1913);
and U1153 (N_1153,In_327,In_162);
nand U1154 (N_1154,In_1457,In_954);
or U1155 (N_1155,In_244,In_1347);
xnor U1156 (N_1156,In_853,In_1528);
or U1157 (N_1157,In_1479,In_186);
nor U1158 (N_1158,In_1942,In_1435);
and U1159 (N_1159,In_367,In_521);
or U1160 (N_1160,In_1841,In_1627);
nand U1161 (N_1161,In_149,In_1289);
and U1162 (N_1162,In_372,In_791);
and U1163 (N_1163,In_1256,In_1743);
or U1164 (N_1164,In_852,In_981);
and U1165 (N_1165,In_1431,In_1);
nand U1166 (N_1166,In_1147,In_1889);
nor U1167 (N_1167,In_1323,In_1959);
nor U1168 (N_1168,In_606,In_576);
or U1169 (N_1169,In_1002,In_1488);
xor U1170 (N_1170,In_153,In_1213);
xnor U1171 (N_1171,In_36,In_1165);
and U1172 (N_1172,In_747,In_200);
or U1173 (N_1173,In_752,In_1151);
nand U1174 (N_1174,In_1535,In_583);
or U1175 (N_1175,In_1620,In_1748);
or U1176 (N_1176,In_1597,In_1825);
xnor U1177 (N_1177,In_43,In_1588);
xnor U1178 (N_1178,In_82,In_1164);
xor U1179 (N_1179,In_1547,In_220);
nor U1180 (N_1180,In_1191,In_1135);
nand U1181 (N_1181,In_375,In_1704);
nand U1182 (N_1182,In_430,In_1332);
nor U1183 (N_1183,In_589,In_1631);
nor U1184 (N_1184,In_226,In_646);
nand U1185 (N_1185,In_1905,In_1484);
nand U1186 (N_1186,In_1659,In_1359);
or U1187 (N_1187,In_557,In_117);
xnor U1188 (N_1188,In_1709,In_1456);
xor U1189 (N_1189,In_1954,In_41);
or U1190 (N_1190,In_54,In_916);
xor U1191 (N_1191,In_1764,In_203);
nand U1192 (N_1192,In_832,In_1455);
or U1193 (N_1193,In_445,In_1633);
or U1194 (N_1194,In_1817,In_893);
nor U1195 (N_1195,In_1238,In_1377);
nor U1196 (N_1196,In_227,In_956);
xor U1197 (N_1197,In_771,In_1762);
nor U1198 (N_1198,In_1282,In_1332);
xor U1199 (N_1199,In_1786,In_1954);
or U1200 (N_1200,In_1529,In_1745);
nor U1201 (N_1201,In_591,In_918);
and U1202 (N_1202,In_117,In_69);
and U1203 (N_1203,In_1589,In_557);
nand U1204 (N_1204,In_746,In_98);
or U1205 (N_1205,In_1605,In_1441);
nor U1206 (N_1206,In_1698,In_561);
and U1207 (N_1207,In_1130,In_667);
and U1208 (N_1208,In_424,In_1849);
xnor U1209 (N_1209,In_1915,In_295);
and U1210 (N_1210,In_46,In_271);
nand U1211 (N_1211,In_1242,In_514);
and U1212 (N_1212,In_488,In_934);
xnor U1213 (N_1213,In_815,In_1804);
xnor U1214 (N_1214,In_522,In_1529);
xor U1215 (N_1215,In_1791,In_292);
or U1216 (N_1216,In_1138,In_89);
xnor U1217 (N_1217,In_1137,In_962);
xor U1218 (N_1218,In_134,In_1023);
nor U1219 (N_1219,In_1776,In_925);
nor U1220 (N_1220,In_888,In_234);
xor U1221 (N_1221,In_1242,In_1985);
or U1222 (N_1222,In_988,In_35);
nor U1223 (N_1223,In_1109,In_11);
nor U1224 (N_1224,In_467,In_1595);
and U1225 (N_1225,In_1190,In_1583);
or U1226 (N_1226,In_1556,In_1024);
nand U1227 (N_1227,In_1452,In_633);
xor U1228 (N_1228,In_226,In_867);
nand U1229 (N_1229,In_19,In_1760);
nor U1230 (N_1230,In_823,In_1003);
xnor U1231 (N_1231,In_1851,In_975);
nand U1232 (N_1232,In_426,In_1992);
nand U1233 (N_1233,In_486,In_156);
xnor U1234 (N_1234,In_807,In_1281);
xnor U1235 (N_1235,In_1817,In_1964);
xnor U1236 (N_1236,In_846,In_991);
xnor U1237 (N_1237,In_1208,In_792);
or U1238 (N_1238,In_571,In_472);
xnor U1239 (N_1239,In_1608,In_1901);
xnor U1240 (N_1240,In_486,In_1611);
xor U1241 (N_1241,In_209,In_1578);
and U1242 (N_1242,In_703,In_373);
nand U1243 (N_1243,In_1012,In_532);
and U1244 (N_1244,In_489,In_79);
and U1245 (N_1245,In_804,In_202);
nor U1246 (N_1246,In_116,In_407);
nor U1247 (N_1247,In_1929,In_483);
nand U1248 (N_1248,In_1953,In_1734);
or U1249 (N_1249,In_959,In_1713);
nor U1250 (N_1250,In_852,In_1219);
nand U1251 (N_1251,In_1671,In_1759);
or U1252 (N_1252,In_257,In_1571);
nand U1253 (N_1253,In_1718,In_905);
nor U1254 (N_1254,In_1271,In_1988);
xnor U1255 (N_1255,In_1259,In_795);
xor U1256 (N_1256,In_1677,In_1451);
nor U1257 (N_1257,In_826,In_664);
nand U1258 (N_1258,In_1193,In_1564);
nand U1259 (N_1259,In_1133,In_672);
xor U1260 (N_1260,In_1039,In_587);
and U1261 (N_1261,In_1987,In_579);
and U1262 (N_1262,In_144,In_1412);
xnor U1263 (N_1263,In_1927,In_267);
xnor U1264 (N_1264,In_24,In_441);
nand U1265 (N_1265,In_1102,In_19);
xnor U1266 (N_1266,In_1769,In_830);
nor U1267 (N_1267,In_1423,In_1624);
nor U1268 (N_1268,In_330,In_284);
nor U1269 (N_1269,In_1740,In_1784);
and U1270 (N_1270,In_1198,In_1670);
xor U1271 (N_1271,In_855,In_68);
and U1272 (N_1272,In_1384,In_1310);
xor U1273 (N_1273,In_1589,In_1492);
or U1274 (N_1274,In_538,In_1967);
nand U1275 (N_1275,In_903,In_413);
nor U1276 (N_1276,In_897,In_1948);
nand U1277 (N_1277,In_908,In_1652);
and U1278 (N_1278,In_1483,In_1021);
xnor U1279 (N_1279,In_1492,In_724);
xnor U1280 (N_1280,In_1836,In_33);
or U1281 (N_1281,In_1701,In_1108);
nand U1282 (N_1282,In_1903,In_1094);
or U1283 (N_1283,In_1616,In_968);
or U1284 (N_1284,In_681,In_403);
or U1285 (N_1285,In_1899,In_1280);
nand U1286 (N_1286,In_363,In_1608);
nand U1287 (N_1287,In_1767,In_796);
and U1288 (N_1288,In_958,In_1541);
xnor U1289 (N_1289,In_643,In_1517);
nor U1290 (N_1290,In_1995,In_489);
or U1291 (N_1291,In_1142,In_343);
or U1292 (N_1292,In_1258,In_1653);
xor U1293 (N_1293,In_1678,In_1918);
nand U1294 (N_1294,In_1219,In_1621);
or U1295 (N_1295,In_790,In_223);
nor U1296 (N_1296,In_1239,In_1154);
and U1297 (N_1297,In_1776,In_985);
nor U1298 (N_1298,In_1368,In_1937);
and U1299 (N_1299,In_1659,In_908);
nor U1300 (N_1300,In_1947,In_392);
or U1301 (N_1301,In_680,In_1642);
xor U1302 (N_1302,In_1349,In_1744);
nor U1303 (N_1303,In_1227,In_1382);
or U1304 (N_1304,In_591,In_1036);
and U1305 (N_1305,In_1032,In_1287);
or U1306 (N_1306,In_560,In_1170);
and U1307 (N_1307,In_1043,In_379);
nand U1308 (N_1308,In_1043,In_1554);
and U1309 (N_1309,In_1763,In_1180);
and U1310 (N_1310,In_59,In_1036);
xnor U1311 (N_1311,In_964,In_1183);
or U1312 (N_1312,In_460,In_293);
nand U1313 (N_1313,In_1553,In_1166);
or U1314 (N_1314,In_30,In_601);
nand U1315 (N_1315,In_407,In_139);
and U1316 (N_1316,In_414,In_679);
nor U1317 (N_1317,In_1914,In_1996);
or U1318 (N_1318,In_888,In_1025);
or U1319 (N_1319,In_1638,In_1758);
nor U1320 (N_1320,In_233,In_426);
and U1321 (N_1321,In_1039,In_95);
or U1322 (N_1322,In_1770,In_786);
xor U1323 (N_1323,In_1323,In_1657);
nor U1324 (N_1324,In_369,In_1830);
and U1325 (N_1325,In_67,In_1633);
xnor U1326 (N_1326,In_561,In_1230);
nor U1327 (N_1327,In_1535,In_45);
or U1328 (N_1328,In_856,In_1342);
or U1329 (N_1329,In_489,In_1684);
nor U1330 (N_1330,In_525,In_1866);
nor U1331 (N_1331,In_96,In_989);
and U1332 (N_1332,In_1346,In_391);
and U1333 (N_1333,In_1378,In_1522);
xnor U1334 (N_1334,In_1703,In_26);
nand U1335 (N_1335,In_179,In_1205);
nor U1336 (N_1336,In_1279,In_886);
or U1337 (N_1337,In_1983,In_997);
xnor U1338 (N_1338,In_535,In_1772);
or U1339 (N_1339,In_1615,In_1792);
nor U1340 (N_1340,In_720,In_1590);
nand U1341 (N_1341,In_881,In_336);
or U1342 (N_1342,In_1267,In_1835);
nand U1343 (N_1343,In_525,In_1416);
and U1344 (N_1344,In_1823,In_1904);
or U1345 (N_1345,In_1285,In_1542);
nor U1346 (N_1346,In_665,In_1795);
nand U1347 (N_1347,In_1723,In_1194);
xnor U1348 (N_1348,In_1007,In_1773);
or U1349 (N_1349,In_476,In_643);
xnor U1350 (N_1350,In_833,In_752);
and U1351 (N_1351,In_720,In_1766);
nor U1352 (N_1352,In_1426,In_1807);
nor U1353 (N_1353,In_1457,In_480);
or U1354 (N_1354,In_1696,In_723);
or U1355 (N_1355,In_52,In_1831);
xor U1356 (N_1356,In_1822,In_1777);
and U1357 (N_1357,In_561,In_905);
nor U1358 (N_1358,In_1197,In_1348);
nor U1359 (N_1359,In_355,In_217);
xor U1360 (N_1360,In_205,In_1687);
xnor U1361 (N_1361,In_138,In_559);
xor U1362 (N_1362,In_1997,In_1663);
or U1363 (N_1363,In_364,In_19);
or U1364 (N_1364,In_95,In_737);
nand U1365 (N_1365,In_1581,In_1062);
nand U1366 (N_1366,In_1094,In_676);
xnor U1367 (N_1367,In_602,In_1053);
xor U1368 (N_1368,In_90,In_921);
nor U1369 (N_1369,In_1906,In_763);
and U1370 (N_1370,In_223,In_893);
or U1371 (N_1371,In_1928,In_887);
or U1372 (N_1372,In_1337,In_584);
and U1373 (N_1373,In_1869,In_1448);
nand U1374 (N_1374,In_182,In_588);
and U1375 (N_1375,In_150,In_775);
or U1376 (N_1376,In_520,In_1475);
xor U1377 (N_1377,In_1080,In_292);
nand U1378 (N_1378,In_783,In_1457);
xnor U1379 (N_1379,In_1494,In_404);
xor U1380 (N_1380,In_1273,In_1980);
nor U1381 (N_1381,In_1568,In_1510);
nor U1382 (N_1382,In_1083,In_1569);
nand U1383 (N_1383,In_479,In_42);
nor U1384 (N_1384,In_1242,In_597);
or U1385 (N_1385,In_1309,In_1883);
nand U1386 (N_1386,In_1170,In_1821);
and U1387 (N_1387,In_10,In_530);
nor U1388 (N_1388,In_1047,In_225);
and U1389 (N_1389,In_680,In_1155);
and U1390 (N_1390,In_1687,In_1157);
nand U1391 (N_1391,In_641,In_752);
nor U1392 (N_1392,In_1711,In_130);
nand U1393 (N_1393,In_1808,In_1848);
and U1394 (N_1394,In_1203,In_960);
or U1395 (N_1395,In_1432,In_1429);
or U1396 (N_1396,In_1757,In_1684);
xnor U1397 (N_1397,In_1877,In_848);
and U1398 (N_1398,In_874,In_73);
nand U1399 (N_1399,In_1464,In_170);
or U1400 (N_1400,In_552,In_562);
and U1401 (N_1401,In_944,In_1235);
or U1402 (N_1402,In_738,In_1907);
nand U1403 (N_1403,In_51,In_991);
and U1404 (N_1404,In_1569,In_1480);
nor U1405 (N_1405,In_1706,In_1508);
nand U1406 (N_1406,In_1493,In_1790);
nor U1407 (N_1407,In_653,In_1789);
nand U1408 (N_1408,In_1592,In_738);
nand U1409 (N_1409,In_1176,In_1582);
or U1410 (N_1410,In_830,In_1196);
xor U1411 (N_1411,In_109,In_539);
or U1412 (N_1412,In_302,In_800);
nand U1413 (N_1413,In_589,In_1923);
and U1414 (N_1414,In_727,In_1166);
nor U1415 (N_1415,In_1201,In_1857);
and U1416 (N_1416,In_1503,In_1112);
nor U1417 (N_1417,In_1282,In_198);
nand U1418 (N_1418,In_326,In_1587);
nor U1419 (N_1419,In_943,In_1928);
nor U1420 (N_1420,In_77,In_1003);
or U1421 (N_1421,In_418,In_767);
and U1422 (N_1422,In_664,In_4);
nand U1423 (N_1423,In_803,In_60);
or U1424 (N_1424,In_1496,In_1859);
and U1425 (N_1425,In_1616,In_1684);
xnor U1426 (N_1426,In_506,In_1970);
and U1427 (N_1427,In_426,In_693);
nor U1428 (N_1428,In_676,In_625);
xor U1429 (N_1429,In_100,In_717);
nand U1430 (N_1430,In_1077,In_417);
and U1431 (N_1431,In_1073,In_1251);
and U1432 (N_1432,In_1491,In_144);
xnor U1433 (N_1433,In_232,In_588);
or U1434 (N_1434,In_522,In_1333);
nand U1435 (N_1435,In_1609,In_862);
nand U1436 (N_1436,In_1720,In_1999);
xnor U1437 (N_1437,In_1242,In_947);
xor U1438 (N_1438,In_315,In_1649);
nand U1439 (N_1439,In_1753,In_218);
and U1440 (N_1440,In_87,In_955);
and U1441 (N_1441,In_50,In_165);
nand U1442 (N_1442,In_1038,In_167);
or U1443 (N_1443,In_313,In_441);
xor U1444 (N_1444,In_1481,In_630);
and U1445 (N_1445,In_1285,In_1157);
nand U1446 (N_1446,In_704,In_668);
xor U1447 (N_1447,In_755,In_915);
xor U1448 (N_1448,In_1601,In_1754);
or U1449 (N_1449,In_930,In_314);
and U1450 (N_1450,In_1315,In_737);
nand U1451 (N_1451,In_1175,In_108);
nand U1452 (N_1452,In_1278,In_1331);
nor U1453 (N_1453,In_1657,In_864);
nor U1454 (N_1454,In_272,In_298);
and U1455 (N_1455,In_526,In_190);
and U1456 (N_1456,In_346,In_1815);
nand U1457 (N_1457,In_1435,In_1460);
nand U1458 (N_1458,In_1045,In_997);
or U1459 (N_1459,In_639,In_264);
and U1460 (N_1460,In_967,In_1643);
xor U1461 (N_1461,In_1868,In_1753);
nor U1462 (N_1462,In_909,In_1211);
and U1463 (N_1463,In_306,In_172);
nand U1464 (N_1464,In_1226,In_192);
and U1465 (N_1465,In_730,In_700);
nor U1466 (N_1466,In_900,In_957);
nor U1467 (N_1467,In_1014,In_1546);
nor U1468 (N_1468,In_77,In_586);
xor U1469 (N_1469,In_1886,In_1169);
nand U1470 (N_1470,In_1373,In_266);
nand U1471 (N_1471,In_405,In_1878);
xnor U1472 (N_1472,In_3,In_1570);
xor U1473 (N_1473,In_987,In_367);
xnor U1474 (N_1474,In_886,In_1341);
xnor U1475 (N_1475,In_1279,In_1755);
nor U1476 (N_1476,In_177,In_1782);
nor U1477 (N_1477,In_1090,In_769);
nor U1478 (N_1478,In_151,In_1945);
nand U1479 (N_1479,In_699,In_1010);
or U1480 (N_1480,In_930,In_1812);
nor U1481 (N_1481,In_517,In_276);
nor U1482 (N_1482,In_623,In_819);
or U1483 (N_1483,In_830,In_316);
nor U1484 (N_1484,In_515,In_336);
or U1485 (N_1485,In_1038,In_846);
and U1486 (N_1486,In_1460,In_904);
nor U1487 (N_1487,In_627,In_1289);
xnor U1488 (N_1488,In_652,In_1586);
xor U1489 (N_1489,In_1887,In_823);
xnor U1490 (N_1490,In_465,In_149);
or U1491 (N_1491,In_460,In_687);
nand U1492 (N_1492,In_904,In_1082);
or U1493 (N_1493,In_1775,In_753);
xor U1494 (N_1494,In_1982,In_653);
xor U1495 (N_1495,In_1738,In_1630);
or U1496 (N_1496,In_116,In_1670);
and U1497 (N_1497,In_1082,In_1137);
nand U1498 (N_1498,In_1377,In_1996);
or U1499 (N_1499,In_1748,In_463);
and U1500 (N_1500,In_1019,In_1403);
nor U1501 (N_1501,In_1176,In_1844);
nand U1502 (N_1502,In_1789,In_1437);
and U1503 (N_1503,In_639,In_1492);
and U1504 (N_1504,In_759,In_1077);
xnor U1505 (N_1505,In_1286,In_1334);
xor U1506 (N_1506,In_1549,In_877);
nor U1507 (N_1507,In_124,In_319);
nor U1508 (N_1508,In_1433,In_1219);
nand U1509 (N_1509,In_1229,In_1034);
and U1510 (N_1510,In_164,In_1797);
nor U1511 (N_1511,In_182,In_1717);
xor U1512 (N_1512,In_903,In_1729);
nor U1513 (N_1513,In_1033,In_185);
or U1514 (N_1514,In_243,In_525);
nand U1515 (N_1515,In_1601,In_40);
nor U1516 (N_1516,In_792,In_776);
xor U1517 (N_1517,In_798,In_82);
nor U1518 (N_1518,In_1099,In_1204);
xnor U1519 (N_1519,In_338,In_1687);
xnor U1520 (N_1520,In_1652,In_284);
xnor U1521 (N_1521,In_1056,In_387);
xnor U1522 (N_1522,In_25,In_559);
or U1523 (N_1523,In_555,In_1772);
nand U1524 (N_1524,In_1503,In_1765);
xnor U1525 (N_1525,In_150,In_1258);
xnor U1526 (N_1526,In_68,In_1986);
or U1527 (N_1527,In_1594,In_1679);
or U1528 (N_1528,In_400,In_1794);
xnor U1529 (N_1529,In_52,In_407);
nand U1530 (N_1530,In_1614,In_202);
nand U1531 (N_1531,In_481,In_1461);
nand U1532 (N_1532,In_207,In_660);
nand U1533 (N_1533,In_561,In_603);
nor U1534 (N_1534,In_535,In_198);
nor U1535 (N_1535,In_1148,In_478);
or U1536 (N_1536,In_29,In_749);
nor U1537 (N_1537,In_119,In_348);
nand U1538 (N_1538,In_601,In_770);
or U1539 (N_1539,In_1065,In_314);
and U1540 (N_1540,In_500,In_1183);
xnor U1541 (N_1541,In_867,In_9);
and U1542 (N_1542,In_791,In_1892);
or U1543 (N_1543,In_1950,In_872);
nor U1544 (N_1544,In_1284,In_1406);
and U1545 (N_1545,In_678,In_1569);
xor U1546 (N_1546,In_1699,In_65);
nand U1547 (N_1547,In_1913,In_1693);
or U1548 (N_1548,In_1124,In_1670);
or U1549 (N_1549,In_1008,In_925);
or U1550 (N_1550,In_1752,In_633);
xor U1551 (N_1551,In_1902,In_389);
xnor U1552 (N_1552,In_213,In_1846);
nor U1553 (N_1553,In_931,In_1409);
or U1554 (N_1554,In_659,In_60);
nor U1555 (N_1555,In_442,In_1755);
and U1556 (N_1556,In_163,In_888);
xor U1557 (N_1557,In_309,In_898);
xnor U1558 (N_1558,In_900,In_1509);
or U1559 (N_1559,In_1426,In_1845);
nor U1560 (N_1560,In_935,In_1097);
xnor U1561 (N_1561,In_280,In_1063);
nor U1562 (N_1562,In_987,In_1151);
or U1563 (N_1563,In_1692,In_89);
and U1564 (N_1564,In_1064,In_992);
nand U1565 (N_1565,In_276,In_1932);
or U1566 (N_1566,In_387,In_1519);
nand U1567 (N_1567,In_66,In_1907);
nand U1568 (N_1568,In_1607,In_1489);
nor U1569 (N_1569,In_1886,In_976);
and U1570 (N_1570,In_1289,In_1598);
nor U1571 (N_1571,In_1932,In_342);
and U1572 (N_1572,In_759,In_1497);
nor U1573 (N_1573,In_1755,In_1533);
and U1574 (N_1574,In_538,In_1962);
or U1575 (N_1575,In_1341,In_1504);
or U1576 (N_1576,In_149,In_225);
nand U1577 (N_1577,In_275,In_335);
or U1578 (N_1578,In_259,In_1403);
nand U1579 (N_1579,In_1945,In_810);
and U1580 (N_1580,In_1035,In_36);
nor U1581 (N_1581,In_676,In_1288);
or U1582 (N_1582,In_1039,In_511);
or U1583 (N_1583,In_321,In_279);
nor U1584 (N_1584,In_639,In_1933);
xor U1585 (N_1585,In_1385,In_341);
xor U1586 (N_1586,In_114,In_943);
or U1587 (N_1587,In_672,In_500);
or U1588 (N_1588,In_1817,In_377);
xor U1589 (N_1589,In_649,In_337);
xnor U1590 (N_1590,In_886,In_1131);
nor U1591 (N_1591,In_1729,In_569);
nand U1592 (N_1592,In_439,In_1900);
or U1593 (N_1593,In_1190,In_164);
and U1594 (N_1594,In_1401,In_1510);
xnor U1595 (N_1595,In_1165,In_500);
and U1596 (N_1596,In_1958,In_1277);
xor U1597 (N_1597,In_1749,In_85);
or U1598 (N_1598,In_943,In_374);
nor U1599 (N_1599,In_1159,In_1278);
xnor U1600 (N_1600,In_343,In_1863);
nand U1601 (N_1601,In_1798,In_1994);
nand U1602 (N_1602,In_1888,In_696);
nor U1603 (N_1603,In_534,In_372);
nor U1604 (N_1604,In_809,In_1135);
and U1605 (N_1605,In_1811,In_119);
nand U1606 (N_1606,In_929,In_150);
and U1607 (N_1607,In_849,In_1791);
and U1608 (N_1608,In_323,In_1119);
xor U1609 (N_1609,In_1366,In_802);
xnor U1610 (N_1610,In_1896,In_850);
nand U1611 (N_1611,In_902,In_1740);
nand U1612 (N_1612,In_1280,In_977);
nand U1613 (N_1613,In_722,In_203);
nor U1614 (N_1614,In_1047,In_1276);
and U1615 (N_1615,In_1574,In_1914);
xnor U1616 (N_1616,In_346,In_1356);
nand U1617 (N_1617,In_1484,In_492);
nor U1618 (N_1618,In_202,In_969);
or U1619 (N_1619,In_510,In_196);
xnor U1620 (N_1620,In_1352,In_1178);
nor U1621 (N_1621,In_1792,In_1928);
or U1622 (N_1622,In_738,In_76);
nand U1623 (N_1623,In_1825,In_1534);
and U1624 (N_1624,In_787,In_1408);
nor U1625 (N_1625,In_1285,In_1963);
nand U1626 (N_1626,In_1991,In_1446);
or U1627 (N_1627,In_222,In_1290);
xnor U1628 (N_1628,In_627,In_1926);
nand U1629 (N_1629,In_1221,In_1459);
nand U1630 (N_1630,In_41,In_148);
and U1631 (N_1631,In_1937,In_1500);
nor U1632 (N_1632,In_843,In_1033);
and U1633 (N_1633,In_1367,In_833);
nand U1634 (N_1634,In_851,In_572);
and U1635 (N_1635,In_526,In_1811);
and U1636 (N_1636,In_1954,In_1368);
and U1637 (N_1637,In_1793,In_1086);
nand U1638 (N_1638,In_934,In_15);
or U1639 (N_1639,In_1890,In_1986);
xnor U1640 (N_1640,In_903,In_478);
nand U1641 (N_1641,In_1771,In_283);
or U1642 (N_1642,In_1546,In_366);
xnor U1643 (N_1643,In_854,In_33);
nand U1644 (N_1644,In_1228,In_833);
xor U1645 (N_1645,In_1727,In_98);
or U1646 (N_1646,In_1787,In_1401);
and U1647 (N_1647,In_97,In_452);
or U1648 (N_1648,In_434,In_52);
xor U1649 (N_1649,In_1035,In_73);
xnor U1650 (N_1650,In_999,In_844);
xor U1651 (N_1651,In_1217,In_612);
nand U1652 (N_1652,In_631,In_1194);
nor U1653 (N_1653,In_71,In_770);
xnor U1654 (N_1654,In_1412,In_330);
nand U1655 (N_1655,In_1237,In_1371);
nor U1656 (N_1656,In_1057,In_213);
and U1657 (N_1657,In_826,In_309);
nor U1658 (N_1658,In_1852,In_1959);
nor U1659 (N_1659,In_597,In_1879);
xnor U1660 (N_1660,In_1173,In_1267);
nand U1661 (N_1661,In_309,In_21);
and U1662 (N_1662,In_1245,In_1354);
nand U1663 (N_1663,In_1668,In_1165);
or U1664 (N_1664,In_1645,In_1658);
xnor U1665 (N_1665,In_500,In_255);
xnor U1666 (N_1666,In_656,In_1700);
or U1667 (N_1667,In_1977,In_558);
or U1668 (N_1668,In_1038,In_267);
and U1669 (N_1669,In_1068,In_1000);
nor U1670 (N_1670,In_132,In_359);
nor U1671 (N_1671,In_880,In_387);
or U1672 (N_1672,In_96,In_66);
xnor U1673 (N_1673,In_1323,In_1450);
nand U1674 (N_1674,In_1064,In_1357);
and U1675 (N_1675,In_1174,In_488);
or U1676 (N_1676,In_1696,In_1985);
and U1677 (N_1677,In_696,In_1230);
and U1678 (N_1678,In_816,In_558);
xnor U1679 (N_1679,In_1921,In_1307);
nand U1680 (N_1680,In_1111,In_1676);
nor U1681 (N_1681,In_1474,In_814);
xnor U1682 (N_1682,In_1466,In_590);
xnor U1683 (N_1683,In_245,In_502);
and U1684 (N_1684,In_580,In_1044);
xnor U1685 (N_1685,In_1625,In_442);
and U1686 (N_1686,In_294,In_844);
and U1687 (N_1687,In_904,In_1919);
nor U1688 (N_1688,In_162,In_1399);
nor U1689 (N_1689,In_1118,In_891);
and U1690 (N_1690,In_1713,In_1819);
and U1691 (N_1691,In_290,In_816);
xnor U1692 (N_1692,In_192,In_444);
xnor U1693 (N_1693,In_394,In_425);
and U1694 (N_1694,In_688,In_542);
or U1695 (N_1695,In_1044,In_1620);
nor U1696 (N_1696,In_991,In_820);
nor U1697 (N_1697,In_1748,In_1839);
and U1698 (N_1698,In_571,In_780);
xnor U1699 (N_1699,In_1991,In_1183);
nand U1700 (N_1700,In_671,In_1812);
or U1701 (N_1701,In_1399,In_569);
xor U1702 (N_1702,In_460,In_944);
nor U1703 (N_1703,In_559,In_339);
nor U1704 (N_1704,In_270,In_358);
xnor U1705 (N_1705,In_1211,In_1499);
or U1706 (N_1706,In_55,In_1841);
nand U1707 (N_1707,In_1883,In_1668);
and U1708 (N_1708,In_304,In_1698);
xor U1709 (N_1709,In_162,In_613);
nand U1710 (N_1710,In_21,In_98);
and U1711 (N_1711,In_809,In_1186);
and U1712 (N_1712,In_381,In_461);
nor U1713 (N_1713,In_666,In_97);
xnor U1714 (N_1714,In_1906,In_1333);
and U1715 (N_1715,In_1369,In_323);
or U1716 (N_1716,In_1238,In_665);
and U1717 (N_1717,In_1298,In_1827);
and U1718 (N_1718,In_274,In_1075);
and U1719 (N_1719,In_1300,In_1895);
or U1720 (N_1720,In_1021,In_1851);
xnor U1721 (N_1721,In_1284,In_1401);
xor U1722 (N_1722,In_118,In_112);
nand U1723 (N_1723,In_149,In_1979);
nand U1724 (N_1724,In_1885,In_577);
xnor U1725 (N_1725,In_497,In_1649);
xnor U1726 (N_1726,In_819,In_393);
nor U1727 (N_1727,In_1732,In_1639);
and U1728 (N_1728,In_1420,In_1786);
nor U1729 (N_1729,In_1625,In_513);
and U1730 (N_1730,In_1068,In_395);
xor U1731 (N_1731,In_541,In_1473);
nor U1732 (N_1732,In_1501,In_1057);
nor U1733 (N_1733,In_1499,In_1483);
nor U1734 (N_1734,In_1428,In_213);
or U1735 (N_1735,In_525,In_1880);
and U1736 (N_1736,In_543,In_885);
and U1737 (N_1737,In_843,In_228);
nand U1738 (N_1738,In_1088,In_1004);
and U1739 (N_1739,In_603,In_554);
xor U1740 (N_1740,In_1577,In_673);
nor U1741 (N_1741,In_574,In_912);
nor U1742 (N_1742,In_1862,In_1008);
xnor U1743 (N_1743,In_821,In_91);
xnor U1744 (N_1744,In_260,In_1594);
nand U1745 (N_1745,In_509,In_1243);
or U1746 (N_1746,In_338,In_1516);
nand U1747 (N_1747,In_708,In_1742);
xnor U1748 (N_1748,In_1962,In_1613);
nor U1749 (N_1749,In_720,In_670);
nand U1750 (N_1750,In_1341,In_1424);
xnor U1751 (N_1751,In_1997,In_528);
nand U1752 (N_1752,In_429,In_445);
and U1753 (N_1753,In_1406,In_305);
and U1754 (N_1754,In_726,In_411);
or U1755 (N_1755,In_1765,In_329);
nor U1756 (N_1756,In_59,In_511);
nand U1757 (N_1757,In_1381,In_507);
xnor U1758 (N_1758,In_216,In_1985);
xor U1759 (N_1759,In_265,In_1610);
or U1760 (N_1760,In_583,In_1309);
xor U1761 (N_1761,In_1848,In_409);
nand U1762 (N_1762,In_1014,In_1837);
nor U1763 (N_1763,In_1583,In_1034);
or U1764 (N_1764,In_920,In_1002);
nor U1765 (N_1765,In_1288,In_525);
and U1766 (N_1766,In_247,In_785);
or U1767 (N_1767,In_1370,In_651);
and U1768 (N_1768,In_1795,In_325);
xor U1769 (N_1769,In_1374,In_1691);
or U1770 (N_1770,In_1039,In_1720);
xnor U1771 (N_1771,In_573,In_830);
nor U1772 (N_1772,In_825,In_1471);
xor U1773 (N_1773,In_1477,In_369);
and U1774 (N_1774,In_624,In_1374);
and U1775 (N_1775,In_1054,In_1804);
or U1776 (N_1776,In_1905,In_1371);
or U1777 (N_1777,In_1275,In_1081);
or U1778 (N_1778,In_1094,In_878);
and U1779 (N_1779,In_402,In_408);
nand U1780 (N_1780,In_934,In_1619);
and U1781 (N_1781,In_958,In_120);
and U1782 (N_1782,In_1117,In_1840);
nor U1783 (N_1783,In_373,In_559);
and U1784 (N_1784,In_1847,In_806);
nor U1785 (N_1785,In_1047,In_750);
xor U1786 (N_1786,In_960,In_1044);
or U1787 (N_1787,In_897,In_1164);
and U1788 (N_1788,In_690,In_157);
and U1789 (N_1789,In_967,In_529);
or U1790 (N_1790,In_208,In_1394);
and U1791 (N_1791,In_155,In_123);
xnor U1792 (N_1792,In_1545,In_1696);
nand U1793 (N_1793,In_702,In_103);
nor U1794 (N_1794,In_1899,In_1130);
nor U1795 (N_1795,In_123,In_467);
and U1796 (N_1796,In_603,In_1575);
nand U1797 (N_1797,In_782,In_1339);
or U1798 (N_1798,In_1766,In_1082);
nor U1799 (N_1799,In_153,In_1406);
nand U1800 (N_1800,In_396,In_469);
xor U1801 (N_1801,In_926,In_349);
and U1802 (N_1802,In_1028,In_1448);
nor U1803 (N_1803,In_1733,In_646);
xor U1804 (N_1804,In_854,In_1676);
nor U1805 (N_1805,In_917,In_1922);
and U1806 (N_1806,In_1204,In_1631);
nor U1807 (N_1807,In_400,In_160);
xor U1808 (N_1808,In_931,In_293);
nand U1809 (N_1809,In_1756,In_1432);
nand U1810 (N_1810,In_600,In_1312);
xnor U1811 (N_1811,In_794,In_1876);
or U1812 (N_1812,In_228,In_842);
or U1813 (N_1813,In_581,In_759);
nor U1814 (N_1814,In_1075,In_1773);
xnor U1815 (N_1815,In_392,In_1515);
nand U1816 (N_1816,In_716,In_1020);
and U1817 (N_1817,In_314,In_21);
nand U1818 (N_1818,In_403,In_1468);
nor U1819 (N_1819,In_345,In_1070);
or U1820 (N_1820,In_1835,In_776);
nor U1821 (N_1821,In_564,In_1998);
nor U1822 (N_1822,In_1814,In_981);
xor U1823 (N_1823,In_367,In_1201);
and U1824 (N_1824,In_983,In_614);
nand U1825 (N_1825,In_1466,In_1256);
nor U1826 (N_1826,In_443,In_1697);
nor U1827 (N_1827,In_1868,In_898);
or U1828 (N_1828,In_630,In_1179);
and U1829 (N_1829,In_609,In_1241);
xor U1830 (N_1830,In_433,In_511);
nor U1831 (N_1831,In_1786,In_163);
or U1832 (N_1832,In_275,In_410);
xnor U1833 (N_1833,In_325,In_211);
xnor U1834 (N_1834,In_917,In_422);
nor U1835 (N_1835,In_1257,In_891);
xnor U1836 (N_1836,In_1780,In_1691);
nand U1837 (N_1837,In_1625,In_648);
nor U1838 (N_1838,In_1614,In_363);
and U1839 (N_1839,In_1497,In_751);
nand U1840 (N_1840,In_117,In_674);
and U1841 (N_1841,In_1512,In_1189);
and U1842 (N_1842,In_404,In_3);
nand U1843 (N_1843,In_1004,In_906);
nand U1844 (N_1844,In_785,In_39);
and U1845 (N_1845,In_1919,In_1055);
xor U1846 (N_1846,In_1926,In_588);
xor U1847 (N_1847,In_349,In_809);
and U1848 (N_1848,In_1387,In_1970);
and U1849 (N_1849,In_1230,In_399);
or U1850 (N_1850,In_1411,In_1678);
and U1851 (N_1851,In_638,In_1750);
or U1852 (N_1852,In_1514,In_1366);
nor U1853 (N_1853,In_1550,In_353);
nor U1854 (N_1854,In_358,In_796);
xnor U1855 (N_1855,In_854,In_1869);
or U1856 (N_1856,In_113,In_1874);
nand U1857 (N_1857,In_1871,In_1298);
xnor U1858 (N_1858,In_1402,In_655);
xnor U1859 (N_1859,In_1335,In_1722);
nand U1860 (N_1860,In_1727,In_1890);
xor U1861 (N_1861,In_628,In_1458);
nand U1862 (N_1862,In_425,In_1156);
or U1863 (N_1863,In_982,In_1777);
or U1864 (N_1864,In_1701,In_1679);
xnor U1865 (N_1865,In_614,In_1668);
or U1866 (N_1866,In_1155,In_1983);
or U1867 (N_1867,In_727,In_1735);
or U1868 (N_1868,In_353,In_1396);
nand U1869 (N_1869,In_1603,In_1733);
nor U1870 (N_1870,In_822,In_1867);
xnor U1871 (N_1871,In_1959,In_1811);
nand U1872 (N_1872,In_1669,In_1272);
nand U1873 (N_1873,In_1981,In_1017);
and U1874 (N_1874,In_1452,In_190);
or U1875 (N_1875,In_1688,In_1191);
nand U1876 (N_1876,In_712,In_312);
nand U1877 (N_1877,In_642,In_1331);
or U1878 (N_1878,In_1650,In_1543);
nor U1879 (N_1879,In_220,In_1963);
xnor U1880 (N_1880,In_971,In_1183);
xnor U1881 (N_1881,In_71,In_700);
or U1882 (N_1882,In_1999,In_406);
xor U1883 (N_1883,In_1556,In_1941);
nand U1884 (N_1884,In_275,In_1149);
or U1885 (N_1885,In_925,In_349);
xnor U1886 (N_1886,In_645,In_136);
xnor U1887 (N_1887,In_617,In_250);
nor U1888 (N_1888,In_1272,In_1912);
xnor U1889 (N_1889,In_319,In_82);
xor U1890 (N_1890,In_1092,In_1367);
nand U1891 (N_1891,In_376,In_985);
nand U1892 (N_1892,In_615,In_1150);
nor U1893 (N_1893,In_1671,In_285);
nand U1894 (N_1894,In_272,In_555);
nor U1895 (N_1895,In_1046,In_1965);
nand U1896 (N_1896,In_282,In_1794);
or U1897 (N_1897,In_1917,In_91);
and U1898 (N_1898,In_57,In_261);
and U1899 (N_1899,In_1873,In_1947);
or U1900 (N_1900,In_1239,In_1360);
nor U1901 (N_1901,In_250,In_1585);
or U1902 (N_1902,In_165,In_567);
xnor U1903 (N_1903,In_1814,In_1331);
nor U1904 (N_1904,In_1982,In_266);
nand U1905 (N_1905,In_482,In_415);
nor U1906 (N_1906,In_1851,In_1408);
or U1907 (N_1907,In_452,In_258);
nand U1908 (N_1908,In_1069,In_276);
xnor U1909 (N_1909,In_182,In_1906);
and U1910 (N_1910,In_926,In_1822);
and U1911 (N_1911,In_814,In_1270);
and U1912 (N_1912,In_1988,In_1574);
nand U1913 (N_1913,In_187,In_1480);
xnor U1914 (N_1914,In_264,In_1663);
or U1915 (N_1915,In_452,In_404);
or U1916 (N_1916,In_592,In_1429);
nand U1917 (N_1917,In_1960,In_1816);
nor U1918 (N_1918,In_1055,In_337);
and U1919 (N_1919,In_615,In_458);
or U1920 (N_1920,In_161,In_1378);
nand U1921 (N_1921,In_1727,In_86);
and U1922 (N_1922,In_1214,In_1119);
and U1923 (N_1923,In_860,In_995);
xor U1924 (N_1924,In_1917,In_1093);
and U1925 (N_1925,In_1518,In_1387);
xnor U1926 (N_1926,In_1342,In_556);
nand U1927 (N_1927,In_1462,In_428);
xor U1928 (N_1928,In_133,In_1804);
nor U1929 (N_1929,In_969,In_1795);
nor U1930 (N_1930,In_970,In_1225);
nand U1931 (N_1931,In_1168,In_1166);
nor U1932 (N_1932,In_309,In_1102);
nor U1933 (N_1933,In_537,In_1755);
nand U1934 (N_1934,In_1891,In_850);
nor U1935 (N_1935,In_1145,In_118);
xnor U1936 (N_1936,In_222,In_166);
xnor U1937 (N_1937,In_52,In_1186);
and U1938 (N_1938,In_112,In_82);
nor U1939 (N_1939,In_1153,In_989);
nor U1940 (N_1940,In_1639,In_1337);
and U1941 (N_1941,In_175,In_1007);
or U1942 (N_1942,In_152,In_361);
nand U1943 (N_1943,In_1753,In_1194);
or U1944 (N_1944,In_29,In_800);
and U1945 (N_1945,In_422,In_1093);
xor U1946 (N_1946,In_632,In_1689);
xnor U1947 (N_1947,In_1653,In_942);
xor U1948 (N_1948,In_1486,In_1331);
nand U1949 (N_1949,In_213,In_579);
nor U1950 (N_1950,In_376,In_341);
or U1951 (N_1951,In_1394,In_1452);
nand U1952 (N_1952,In_276,In_1499);
and U1953 (N_1953,In_316,In_1547);
xnor U1954 (N_1954,In_628,In_1227);
and U1955 (N_1955,In_1982,In_892);
nor U1956 (N_1956,In_653,In_519);
nand U1957 (N_1957,In_815,In_1822);
or U1958 (N_1958,In_1587,In_940);
xnor U1959 (N_1959,In_688,In_1014);
nor U1960 (N_1960,In_857,In_843);
or U1961 (N_1961,In_1340,In_1470);
and U1962 (N_1962,In_389,In_61);
xor U1963 (N_1963,In_434,In_422);
and U1964 (N_1964,In_505,In_417);
xor U1965 (N_1965,In_41,In_1351);
nand U1966 (N_1966,In_1113,In_1321);
or U1967 (N_1967,In_584,In_956);
xor U1968 (N_1968,In_437,In_474);
nand U1969 (N_1969,In_259,In_1891);
xor U1970 (N_1970,In_1101,In_487);
nand U1971 (N_1971,In_1438,In_1130);
or U1972 (N_1972,In_280,In_166);
or U1973 (N_1973,In_524,In_208);
and U1974 (N_1974,In_974,In_1267);
xor U1975 (N_1975,In_726,In_578);
xnor U1976 (N_1976,In_449,In_457);
and U1977 (N_1977,In_146,In_551);
nand U1978 (N_1978,In_704,In_1421);
and U1979 (N_1979,In_1186,In_1432);
xnor U1980 (N_1980,In_920,In_861);
or U1981 (N_1981,In_1304,In_751);
xor U1982 (N_1982,In_156,In_311);
xnor U1983 (N_1983,In_1865,In_647);
nand U1984 (N_1984,In_268,In_515);
or U1985 (N_1985,In_1204,In_136);
nor U1986 (N_1986,In_829,In_1002);
nand U1987 (N_1987,In_241,In_1736);
nor U1988 (N_1988,In_1025,In_1413);
or U1989 (N_1989,In_1504,In_1337);
and U1990 (N_1990,In_912,In_1061);
and U1991 (N_1991,In_1714,In_1672);
nor U1992 (N_1992,In_1944,In_697);
nand U1993 (N_1993,In_538,In_1458);
or U1994 (N_1994,In_732,In_1994);
xor U1995 (N_1995,In_409,In_1939);
nor U1996 (N_1996,In_1122,In_1163);
xor U1997 (N_1997,In_1697,In_1673);
and U1998 (N_1998,In_1718,In_521);
nand U1999 (N_1999,In_368,In_1092);
and U2000 (N_2000,In_425,In_869);
or U2001 (N_2001,In_1937,In_520);
and U2002 (N_2002,In_346,In_1394);
xor U2003 (N_2003,In_1277,In_74);
nor U2004 (N_2004,In_1980,In_1428);
and U2005 (N_2005,In_96,In_456);
or U2006 (N_2006,In_264,In_1521);
or U2007 (N_2007,In_1430,In_1285);
xnor U2008 (N_2008,In_1720,In_1892);
xnor U2009 (N_2009,In_1802,In_1034);
and U2010 (N_2010,In_1726,In_393);
and U2011 (N_2011,In_1247,In_667);
or U2012 (N_2012,In_1300,In_1047);
and U2013 (N_2013,In_1062,In_1610);
xor U2014 (N_2014,In_1546,In_1114);
and U2015 (N_2015,In_655,In_1489);
and U2016 (N_2016,In_1616,In_1448);
xnor U2017 (N_2017,In_379,In_59);
nor U2018 (N_2018,In_425,In_658);
nand U2019 (N_2019,In_1071,In_489);
nor U2020 (N_2020,In_388,In_949);
nor U2021 (N_2021,In_571,In_1565);
xnor U2022 (N_2022,In_1361,In_841);
or U2023 (N_2023,In_99,In_1870);
nand U2024 (N_2024,In_482,In_1563);
or U2025 (N_2025,In_725,In_553);
nand U2026 (N_2026,In_1021,In_246);
xor U2027 (N_2027,In_747,In_1509);
and U2028 (N_2028,In_1725,In_1501);
nand U2029 (N_2029,In_1637,In_615);
nand U2030 (N_2030,In_1329,In_705);
nor U2031 (N_2031,In_317,In_988);
and U2032 (N_2032,In_1256,In_139);
nor U2033 (N_2033,In_1511,In_419);
or U2034 (N_2034,In_1055,In_588);
nor U2035 (N_2035,In_1877,In_725);
nor U2036 (N_2036,In_497,In_103);
nor U2037 (N_2037,In_235,In_902);
and U2038 (N_2038,In_1471,In_1323);
and U2039 (N_2039,In_137,In_1046);
xor U2040 (N_2040,In_737,In_843);
and U2041 (N_2041,In_1934,In_226);
nor U2042 (N_2042,In_429,In_212);
nor U2043 (N_2043,In_38,In_224);
xor U2044 (N_2044,In_452,In_1424);
or U2045 (N_2045,In_1265,In_1499);
nand U2046 (N_2046,In_676,In_1165);
xor U2047 (N_2047,In_1564,In_497);
and U2048 (N_2048,In_1237,In_485);
nor U2049 (N_2049,In_746,In_1461);
and U2050 (N_2050,In_780,In_1370);
or U2051 (N_2051,In_533,In_1760);
and U2052 (N_2052,In_1294,In_1470);
nand U2053 (N_2053,In_1233,In_74);
and U2054 (N_2054,In_751,In_664);
xor U2055 (N_2055,In_548,In_1025);
or U2056 (N_2056,In_218,In_473);
or U2057 (N_2057,In_828,In_1637);
xor U2058 (N_2058,In_1980,In_902);
xnor U2059 (N_2059,In_281,In_11);
nor U2060 (N_2060,In_115,In_1941);
nor U2061 (N_2061,In_86,In_856);
nand U2062 (N_2062,In_278,In_114);
or U2063 (N_2063,In_1140,In_1856);
or U2064 (N_2064,In_717,In_74);
xor U2065 (N_2065,In_243,In_486);
xor U2066 (N_2066,In_1032,In_1415);
and U2067 (N_2067,In_144,In_702);
xnor U2068 (N_2068,In_1948,In_976);
xnor U2069 (N_2069,In_1955,In_1924);
and U2070 (N_2070,In_228,In_631);
nand U2071 (N_2071,In_1137,In_1136);
xor U2072 (N_2072,In_40,In_1079);
and U2073 (N_2073,In_1507,In_921);
and U2074 (N_2074,In_920,In_152);
and U2075 (N_2075,In_280,In_1767);
xnor U2076 (N_2076,In_621,In_841);
and U2077 (N_2077,In_375,In_688);
or U2078 (N_2078,In_1015,In_164);
or U2079 (N_2079,In_850,In_916);
nand U2080 (N_2080,In_360,In_1735);
nor U2081 (N_2081,In_1333,In_1026);
and U2082 (N_2082,In_1141,In_410);
xnor U2083 (N_2083,In_660,In_568);
and U2084 (N_2084,In_430,In_1195);
nor U2085 (N_2085,In_1340,In_1549);
and U2086 (N_2086,In_963,In_1573);
or U2087 (N_2087,In_347,In_517);
xnor U2088 (N_2088,In_1403,In_1556);
or U2089 (N_2089,In_221,In_1723);
nand U2090 (N_2090,In_1387,In_319);
and U2091 (N_2091,In_965,In_80);
nor U2092 (N_2092,In_1246,In_1499);
and U2093 (N_2093,In_1596,In_1023);
or U2094 (N_2094,In_1935,In_610);
xnor U2095 (N_2095,In_1302,In_1788);
nor U2096 (N_2096,In_241,In_1044);
or U2097 (N_2097,In_1980,In_1829);
and U2098 (N_2098,In_1479,In_474);
nor U2099 (N_2099,In_1018,In_1816);
nor U2100 (N_2100,In_274,In_1135);
or U2101 (N_2101,In_99,In_1316);
or U2102 (N_2102,In_1870,In_494);
and U2103 (N_2103,In_1894,In_137);
nor U2104 (N_2104,In_1663,In_491);
xnor U2105 (N_2105,In_234,In_1220);
and U2106 (N_2106,In_1270,In_1725);
and U2107 (N_2107,In_95,In_378);
or U2108 (N_2108,In_1847,In_1602);
or U2109 (N_2109,In_1054,In_591);
nor U2110 (N_2110,In_1020,In_721);
nor U2111 (N_2111,In_94,In_1298);
and U2112 (N_2112,In_1002,In_938);
xor U2113 (N_2113,In_613,In_1382);
and U2114 (N_2114,In_1887,In_1198);
xnor U2115 (N_2115,In_169,In_1806);
nand U2116 (N_2116,In_307,In_1994);
nand U2117 (N_2117,In_1331,In_641);
xnor U2118 (N_2118,In_693,In_1603);
nor U2119 (N_2119,In_801,In_857);
or U2120 (N_2120,In_1715,In_1918);
nand U2121 (N_2121,In_211,In_663);
xnor U2122 (N_2122,In_1404,In_385);
nor U2123 (N_2123,In_1796,In_1354);
or U2124 (N_2124,In_878,In_545);
and U2125 (N_2125,In_1336,In_1915);
xor U2126 (N_2126,In_50,In_856);
nand U2127 (N_2127,In_699,In_503);
or U2128 (N_2128,In_370,In_430);
xor U2129 (N_2129,In_515,In_1621);
or U2130 (N_2130,In_1836,In_1878);
or U2131 (N_2131,In_640,In_1420);
or U2132 (N_2132,In_313,In_154);
or U2133 (N_2133,In_996,In_512);
xor U2134 (N_2134,In_1990,In_452);
nand U2135 (N_2135,In_455,In_1519);
nand U2136 (N_2136,In_804,In_1979);
or U2137 (N_2137,In_623,In_1940);
or U2138 (N_2138,In_1864,In_912);
and U2139 (N_2139,In_1048,In_977);
nor U2140 (N_2140,In_964,In_760);
nand U2141 (N_2141,In_1736,In_850);
xor U2142 (N_2142,In_1869,In_507);
or U2143 (N_2143,In_4,In_325);
nor U2144 (N_2144,In_1533,In_1511);
xnor U2145 (N_2145,In_1301,In_937);
nand U2146 (N_2146,In_394,In_1140);
or U2147 (N_2147,In_1189,In_1127);
or U2148 (N_2148,In_800,In_231);
xnor U2149 (N_2149,In_995,In_703);
xor U2150 (N_2150,In_1159,In_234);
xnor U2151 (N_2151,In_254,In_1755);
nor U2152 (N_2152,In_890,In_125);
xor U2153 (N_2153,In_622,In_797);
or U2154 (N_2154,In_355,In_1445);
or U2155 (N_2155,In_1633,In_759);
xnor U2156 (N_2156,In_671,In_1822);
xor U2157 (N_2157,In_1346,In_810);
or U2158 (N_2158,In_49,In_153);
nor U2159 (N_2159,In_1031,In_369);
and U2160 (N_2160,In_993,In_1081);
nand U2161 (N_2161,In_952,In_950);
and U2162 (N_2162,In_454,In_929);
or U2163 (N_2163,In_1105,In_778);
xnor U2164 (N_2164,In_1948,In_894);
and U2165 (N_2165,In_797,In_1002);
xor U2166 (N_2166,In_1243,In_125);
or U2167 (N_2167,In_450,In_990);
nor U2168 (N_2168,In_118,In_16);
and U2169 (N_2169,In_76,In_1608);
nor U2170 (N_2170,In_1343,In_811);
xor U2171 (N_2171,In_480,In_753);
nand U2172 (N_2172,In_1076,In_1767);
nand U2173 (N_2173,In_1757,In_372);
nor U2174 (N_2174,In_150,In_1661);
nand U2175 (N_2175,In_170,In_649);
or U2176 (N_2176,In_181,In_347);
or U2177 (N_2177,In_1746,In_469);
nor U2178 (N_2178,In_267,In_1699);
nand U2179 (N_2179,In_479,In_751);
or U2180 (N_2180,In_708,In_1645);
nor U2181 (N_2181,In_255,In_432);
xor U2182 (N_2182,In_730,In_968);
or U2183 (N_2183,In_1579,In_243);
or U2184 (N_2184,In_655,In_1205);
nand U2185 (N_2185,In_1776,In_217);
or U2186 (N_2186,In_1639,In_1504);
nand U2187 (N_2187,In_275,In_1993);
and U2188 (N_2188,In_501,In_1375);
and U2189 (N_2189,In_1972,In_977);
nor U2190 (N_2190,In_401,In_906);
nor U2191 (N_2191,In_518,In_1136);
nand U2192 (N_2192,In_1386,In_403);
nand U2193 (N_2193,In_602,In_166);
nand U2194 (N_2194,In_1027,In_571);
or U2195 (N_2195,In_647,In_516);
or U2196 (N_2196,In_1510,In_422);
xnor U2197 (N_2197,In_1288,In_996);
nor U2198 (N_2198,In_1117,In_28);
xor U2199 (N_2199,In_1250,In_763);
and U2200 (N_2200,In_1002,In_1157);
xnor U2201 (N_2201,In_685,In_1560);
xor U2202 (N_2202,In_237,In_1051);
nand U2203 (N_2203,In_616,In_1626);
xnor U2204 (N_2204,In_6,In_1179);
nand U2205 (N_2205,In_118,In_1732);
nor U2206 (N_2206,In_518,In_981);
nand U2207 (N_2207,In_1692,In_141);
nand U2208 (N_2208,In_1179,In_101);
and U2209 (N_2209,In_810,In_1234);
or U2210 (N_2210,In_1841,In_311);
or U2211 (N_2211,In_147,In_180);
or U2212 (N_2212,In_874,In_799);
xor U2213 (N_2213,In_1720,In_1687);
and U2214 (N_2214,In_1267,In_825);
nand U2215 (N_2215,In_1342,In_310);
nand U2216 (N_2216,In_1868,In_316);
or U2217 (N_2217,In_1906,In_1841);
and U2218 (N_2218,In_545,In_1671);
xor U2219 (N_2219,In_1449,In_477);
or U2220 (N_2220,In_494,In_984);
nand U2221 (N_2221,In_50,In_1512);
xor U2222 (N_2222,In_938,In_190);
and U2223 (N_2223,In_1,In_1282);
nand U2224 (N_2224,In_866,In_444);
nor U2225 (N_2225,In_189,In_244);
nor U2226 (N_2226,In_1893,In_1036);
or U2227 (N_2227,In_366,In_880);
nor U2228 (N_2228,In_1980,In_1272);
nand U2229 (N_2229,In_72,In_1241);
nor U2230 (N_2230,In_1602,In_787);
nor U2231 (N_2231,In_1630,In_865);
nand U2232 (N_2232,In_1352,In_1335);
and U2233 (N_2233,In_1997,In_487);
nor U2234 (N_2234,In_48,In_335);
nand U2235 (N_2235,In_260,In_1397);
nand U2236 (N_2236,In_1037,In_1986);
or U2237 (N_2237,In_1533,In_335);
and U2238 (N_2238,In_1157,In_1528);
or U2239 (N_2239,In_1006,In_654);
or U2240 (N_2240,In_1799,In_20);
or U2241 (N_2241,In_70,In_1840);
nor U2242 (N_2242,In_962,In_984);
or U2243 (N_2243,In_1524,In_770);
and U2244 (N_2244,In_12,In_1110);
nand U2245 (N_2245,In_1492,In_1030);
or U2246 (N_2246,In_1724,In_343);
xnor U2247 (N_2247,In_1449,In_1475);
and U2248 (N_2248,In_257,In_1269);
nand U2249 (N_2249,In_1232,In_306);
xor U2250 (N_2250,In_1112,In_319);
or U2251 (N_2251,In_356,In_1762);
or U2252 (N_2252,In_680,In_1898);
nand U2253 (N_2253,In_1616,In_1568);
nand U2254 (N_2254,In_1212,In_1252);
xor U2255 (N_2255,In_51,In_1136);
and U2256 (N_2256,In_380,In_1397);
or U2257 (N_2257,In_1023,In_1150);
or U2258 (N_2258,In_1277,In_1605);
xnor U2259 (N_2259,In_49,In_1108);
and U2260 (N_2260,In_1844,In_943);
or U2261 (N_2261,In_102,In_1818);
and U2262 (N_2262,In_210,In_461);
xor U2263 (N_2263,In_440,In_1489);
xnor U2264 (N_2264,In_123,In_1746);
xor U2265 (N_2265,In_1637,In_1660);
nand U2266 (N_2266,In_488,In_387);
nor U2267 (N_2267,In_218,In_139);
or U2268 (N_2268,In_1002,In_688);
nand U2269 (N_2269,In_1311,In_1167);
xnor U2270 (N_2270,In_1671,In_1847);
nand U2271 (N_2271,In_1414,In_754);
nor U2272 (N_2272,In_1847,In_1626);
and U2273 (N_2273,In_47,In_306);
or U2274 (N_2274,In_1056,In_1114);
xor U2275 (N_2275,In_1197,In_1543);
nor U2276 (N_2276,In_477,In_954);
nor U2277 (N_2277,In_424,In_576);
xnor U2278 (N_2278,In_528,In_1647);
or U2279 (N_2279,In_720,In_1672);
nor U2280 (N_2280,In_401,In_67);
xor U2281 (N_2281,In_98,In_437);
and U2282 (N_2282,In_1407,In_88);
nor U2283 (N_2283,In_1972,In_1893);
nor U2284 (N_2284,In_841,In_1460);
and U2285 (N_2285,In_676,In_1680);
nand U2286 (N_2286,In_548,In_1533);
nor U2287 (N_2287,In_1639,In_331);
or U2288 (N_2288,In_611,In_92);
nor U2289 (N_2289,In_1339,In_159);
and U2290 (N_2290,In_648,In_184);
xnor U2291 (N_2291,In_1758,In_433);
xor U2292 (N_2292,In_1350,In_1785);
and U2293 (N_2293,In_1878,In_242);
nor U2294 (N_2294,In_1668,In_1699);
or U2295 (N_2295,In_1901,In_7);
xor U2296 (N_2296,In_185,In_868);
nor U2297 (N_2297,In_1472,In_586);
nor U2298 (N_2298,In_1838,In_1721);
xor U2299 (N_2299,In_761,In_1232);
nand U2300 (N_2300,In_710,In_1392);
nor U2301 (N_2301,In_1401,In_1976);
nand U2302 (N_2302,In_1576,In_1172);
nand U2303 (N_2303,In_1448,In_1833);
xor U2304 (N_2304,In_1147,In_1765);
xor U2305 (N_2305,In_125,In_112);
nand U2306 (N_2306,In_1335,In_321);
nand U2307 (N_2307,In_1231,In_50);
nand U2308 (N_2308,In_437,In_1981);
nor U2309 (N_2309,In_824,In_255);
xor U2310 (N_2310,In_348,In_1528);
or U2311 (N_2311,In_1763,In_79);
nor U2312 (N_2312,In_1319,In_1823);
nor U2313 (N_2313,In_787,In_1216);
nor U2314 (N_2314,In_970,In_1257);
or U2315 (N_2315,In_1173,In_1218);
nor U2316 (N_2316,In_228,In_1328);
or U2317 (N_2317,In_426,In_870);
and U2318 (N_2318,In_268,In_1437);
nor U2319 (N_2319,In_662,In_1965);
or U2320 (N_2320,In_1062,In_791);
nand U2321 (N_2321,In_1257,In_1339);
or U2322 (N_2322,In_877,In_1647);
xor U2323 (N_2323,In_221,In_416);
and U2324 (N_2324,In_528,In_877);
and U2325 (N_2325,In_780,In_797);
nand U2326 (N_2326,In_1958,In_1042);
xnor U2327 (N_2327,In_1003,In_733);
or U2328 (N_2328,In_501,In_11);
and U2329 (N_2329,In_1350,In_1491);
xnor U2330 (N_2330,In_1135,In_1776);
nor U2331 (N_2331,In_798,In_1042);
xnor U2332 (N_2332,In_746,In_957);
xor U2333 (N_2333,In_1873,In_1453);
nor U2334 (N_2334,In_1442,In_21);
or U2335 (N_2335,In_1796,In_1738);
nand U2336 (N_2336,In_1784,In_945);
or U2337 (N_2337,In_1589,In_653);
nor U2338 (N_2338,In_1085,In_1821);
xor U2339 (N_2339,In_1657,In_1574);
and U2340 (N_2340,In_1316,In_287);
nand U2341 (N_2341,In_1758,In_1567);
or U2342 (N_2342,In_1059,In_672);
xnor U2343 (N_2343,In_630,In_523);
and U2344 (N_2344,In_1491,In_304);
and U2345 (N_2345,In_114,In_463);
xor U2346 (N_2346,In_684,In_1819);
or U2347 (N_2347,In_391,In_939);
or U2348 (N_2348,In_918,In_1916);
xor U2349 (N_2349,In_415,In_1279);
xnor U2350 (N_2350,In_674,In_1017);
or U2351 (N_2351,In_466,In_587);
nor U2352 (N_2352,In_1624,In_1650);
nand U2353 (N_2353,In_158,In_813);
nor U2354 (N_2354,In_1498,In_172);
or U2355 (N_2355,In_1479,In_888);
nand U2356 (N_2356,In_602,In_1375);
xor U2357 (N_2357,In_180,In_327);
nor U2358 (N_2358,In_199,In_1304);
nand U2359 (N_2359,In_1281,In_321);
nand U2360 (N_2360,In_877,In_783);
nor U2361 (N_2361,In_1658,In_555);
nand U2362 (N_2362,In_1393,In_1272);
and U2363 (N_2363,In_484,In_249);
nand U2364 (N_2364,In_606,In_290);
nand U2365 (N_2365,In_559,In_1185);
or U2366 (N_2366,In_537,In_57);
nor U2367 (N_2367,In_568,In_783);
or U2368 (N_2368,In_378,In_1905);
xor U2369 (N_2369,In_256,In_1364);
and U2370 (N_2370,In_1704,In_1033);
or U2371 (N_2371,In_712,In_105);
nor U2372 (N_2372,In_1265,In_1933);
and U2373 (N_2373,In_1392,In_887);
or U2374 (N_2374,In_1283,In_1378);
nand U2375 (N_2375,In_795,In_959);
xor U2376 (N_2376,In_1321,In_1387);
and U2377 (N_2377,In_95,In_1308);
nor U2378 (N_2378,In_1242,In_1518);
and U2379 (N_2379,In_439,In_707);
or U2380 (N_2380,In_1025,In_675);
xnor U2381 (N_2381,In_1212,In_1778);
nor U2382 (N_2382,In_1339,In_1506);
and U2383 (N_2383,In_214,In_1887);
or U2384 (N_2384,In_0,In_457);
or U2385 (N_2385,In_1369,In_1382);
xor U2386 (N_2386,In_367,In_1524);
nand U2387 (N_2387,In_1755,In_932);
and U2388 (N_2388,In_117,In_434);
and U2389 (N_2389,In_1795,In_1014);
or U2390 (N_2390,In_781,In_1454);
and U2391 (N_2391,In_538,In_1279);
or U2392 (N_2392,In_60,In_879);
xnor U2393 (N_2393,In_491,In_269);
nor U2394 (N_2394,In_189,In_1131);
nor U2395 (N_2395,In_869,In_1318);
nand U2396 (N_2396,In_1482,In_767);
or U2397 (N_2397,In_1517,In_245);
xor U2398 (N_2398,In_577,In_124);
nor U2399 (N_2399,In_1046,In_623);
xnor U2400 (N_2400,In_548,In_1243);
xnor U2401 (N_2401,In_1030,In_1847);
nand U2402 (N_2402,In_1350,In_656);
or U2403 (N_2403,In_240,In_545);
and U2404 (N_2404,In_1567,In_220);
xor U2405 (N_2405,In_1934,In_824);
and U2406 (N_2406,In_1267,In_58);
or U2407 (N_2407,In_919,In_239);
and U2408 (N_2408,In_1440,In_294);
nand U2409 (N_2409,In_1391,In_1305);
nand U2410 (N_2410,In_1129,In_778);
nand U2411 (N_2411,In_575,In_91);
nor U2412 (N_2412,In_1740,In_1707);
nand U2413 (N_2413,In_952,In_1611);
or U2414 (N_2414,In_1633,In_712);
nand U2415 (N_2415,In_129,In_365);
and U2416 (N_2416,In_266,In_1500);
nand U2417 (N_2417,In_1573,In_351);
and U2418 (N_2418,In_249,In_717);
xnor U2419 (N_2419,In_1971,In_1910);
nor U2420 (N_2420,In_1204,In_1608);
xor U2421 (N_2421,In_1572,In_864);
nor U2422 (N_2422,In_1208,In_1440);
nor U2423 (N_2423,In_1644,In_452);
nor U2424 (N_2424,In_452,In_1634);
xor U2425 (N_2425,In_265,In_705);
xnor U2426 (N_2426,In_1427,In_456);
xor U2427 (N_2427,In_881,In_911);
nor U2428 (N_2428,In_1828,In_364);
nor U2429 (N_2429,In_837,In_291);
and U2430 (N_2430,In_1465,In_1984);
nand U2431 (N_2431,In_27,In_1241);
and U2432 (N_2432,In_1190,In_184);
and U2433 (N_2433,In_1672,In_1993);
or U2434 (N_2434,In_1627,In_441);
and U2435 (N_2435,In_838,In_778);
or U2436 (N_2436,In_1915,In_717);
nor U2437 (N_2437,In_923,In_1480);
xnor U2438 (N_2438,In_1191,In_700);
or U2439 (N_2439,In_1957,In_1492);
or U2440 (N_2440,In_1631,In_1928);
nor U2441 (N_2441,In_1951,In_1007);
nand U2442 (N_2442,In_1701,In_464);
or U2443 (N_2443,In_1883,In_1639);
and U2444 (N_2444,In_1770,In_554);
nor U2445 (N_2445,In_555,In_1227);
xor U2446 (N_2446,In_1093,In_1679);
xnor U2447 (N_2447,In_1430,In_351);
xnor U2448 (N_2448,In_1598,In_1438);
or U2449 (N_2449,In_503,In_1153);
and U2450 (N_2450,In_1307,In_145);
and U2451 (N_2451,In_590,In_910);
and U2452 (N_2452,In_514,In_701);
xnor U2453 (N_2453,In_585,In_1908);
nor U2454 (N_2454,In_1223,In_1409);
or U2455 (N_2455,In_1692,In_1029);
or U2456 (N_2456,In_788,In_1724);
and U2457 (N_2457,In_1795,In_1501);
nand U2458 (N_2458,In_1974,In_1602);
nor U2459 (N_2459,In_312,In_561);
and U2460 (N_2460,In_1120,In_1599);
nand U2461 (N_2461,In_1152,In_1632);
nor U2462 (N_2462,In_113,In_536);
xnor U2463 (N_2463,In_1544,In_1332);
or U2464 (N_2464,In_1623,In_928);
xor U2465 (N_2465,In_489,In_900);
nor U2466 (N_2466,In_1678,In_1480);
xor U2467 (N_2467,In_449,In_1268);
and U2468 (N_2468,In_1564,In_785);
nor U2469 (N_2469,In_1656,In_1264);
nor U2470 (N_2470,In_254,In_1629);
or U2471 (N_2471,In_697,In_1401);
or U2472 (N_2472,In_1439,In_724);
nor U2473 (N_2473,In_254,In_1187);
xor U2474 (N_2474,In_1323,In_641);
and U2475 (N_2475,In_372,In_816);
or U2476 (N_2476,In_1681,In_92);
and U2477 (N_2477,In_1601,In_1396);
xor U2478 (N_2478,In_662,In_1723);
nand U2479 (N_2479,In_1654,In_805);
nand U2480 (N_2480,In_682,In_1036);
or U2481 (N_2481,In_1163,In_1272);
xor U2482 (N_2482,In_1301,In_567);
nand U2483 (N_2483,In_1181,In_1848);
nand U2484 (N_2484,In_186,In_413);
and U2485 (N_2485,In_135,In_1732);
nand U2486 (N_2486,In_508,In_813);
nand U2487 (N_2487,In_1889,In_310);
or U2488 (N_2488,In_1428,In_1757);
nand U2489 (N_2489,In_562,In_1745);
nand U2490 (N_2490,In_737,In_86);
and U2491 (N_2491,In_591,In_1470);
nand U2492 (N_2492,In_1439,In_1016);
nand U2493 (N_2493,In_103,In_1269);
nor U2494 (N_2494,In_444,In_477);
or U2495 (N_2495,In_1290,In_1640);
nor U2496 (N_2496,In_162,In_449);
nand U2497 (N_2497,In_457,In_1409);
or U2498 (N_2498,In_934,In_1239);
nor U2499 (N_2499,In_6,In_1174);
nor U2500 (N_2500,In_1491,In_1462);
and U2501 (N_2501,In_366,In_1995);
xnor U2502 (N_2502,In_1036,In_972);
xnor U2503 (N_2503,In_13,In_1190);
nor U2504 (N_2504,In_827,In_1913);
and U2505 (N_2505,In_771,In_235);
nand U2506 (N_2506,In_946,In_1743);
xor U2507 (N_2507,In_1041,In_627);
nor U2508 (N_2508,In_1531,In_753);
and U2509 (N_2509,In_374,In_1215);
xnor U2510 (N_2510,In_932,In_913);
xor U2511 (N_2511,In_1411,In_487);
xor U2512 (N_2512,In_367,In_1075);
nor U2513 (N_2513,In_1297,In_297);
or U2514 (N_2514,In_29,In_883);
or U2515 (N_2515,In_1109,In_979);
nand U2516 (N_2516,In_1209,In_1283);
and U2517 (N_2517,In_1968,In_1718);
xnor U2518 (N_2518,In_57,In_1880);
or U2519 (N_2519,In_1760,In_655);
or U2520 (N_2520,In_865,In_924);
and U2521 (N_2521,In_669,In_1170);
xor U2522 (N_2522,In_735,In_796);
and U2523 (N_2523,In_631,In_554);
and U2524 (N_2524,In_737,In_682);
and U2525 (N_2525,In_612,In_343);
xnor U2526 (N_2526,In_1034,In_1353);
nor U2527 (N_2527,In_171,In_1843);
and U2528 (N_2528,In_116,In_999);
xor U2529 (N_2529,In_1274,In_929);
or U2530 (N_2530,In_234,In_974);
or U2531 (N_2531,In_1855,In_1291);
xor U2532 (N_2532,In_790,In_863);
nor U2533 (N_2533,In_969,In_1080);
and U2534 (N_2534,In_1367,In_274);
nand U2535 (N_2535,In_1983,In_811);
or U2536 (N_2536,In_483,In_1098);
and U2537 (N_2537,In_310,In_1210);
and U2538 (N_2538,In_1984,In_1420);
nor U2539 (N_2539,In_1662,In_670);
and U2540 (N_2540,In_675,In_193);
xnor U2541 (N_2541,In_864,In_1464);
nand U2542 (N_2542,In_1973,In_1235);
xnor U2543 (N_2543,In_381,In_202);
nand U2544 (N_2544,In_1813,In_635);
xor U2545 (N_2545,In_1000,In_1099);
xnor U2546 (N_2546,In_1581,In_883);
xor U2547 (N_2547,In_405,In_298);
and U2548 (N_2548,In_1165,In_711);
nand U2549 (N_2549,In_1353,In_1009);
nand U2550 (N_2550,In_535,In_97);
or U2551 (N_2551,In_321,In_1104);
or U2552 (N_2552,In_941,In_150);
nor U2553 (N_2553,In_1997,In_468);
nand U2554 (N_2554,In_835,In_1740);
nand U2555 (N_2555,In_194,In_307);
and U2556 (N_2556,In_1430,In_206);
or U2557 (N_2557,In_1077,In_916);
nor U2558 (N_2558,In_58,In_638);
or U2559 (N_2559,In_626,In_1724);
nor U2560 (N_2560,In_524,In_1549);
xnor U2561 (N_2561,In_227,In_483);
xnor U2562 (N_2562,In_242,In_1035);
or U2563 (N_2563,In_1780,In_311);
and U2564 (N_2564,In_1555,In_1526);
nand U2565 (N_2565,In_790,In_1716);
xnor U2566 (N_2566,In_776,In_602);
or U2567 (N_2567,In_203,In_700);
or U2568 (N_2568,In_1626,In_1019);
nand U2569 (N_2569,In_1143,In_829);
and U2570 (N_2570,In_1030,In_306);
and U2571 (N_2571,In_1016,In_101);
xnor U2572 (N_2572,In_349,In_598);
nand U2573 (N_2573,In_1741,In_1883);
nor U2574 (N_2574,In_423,In_1390);
or U2575 (N_2575,In_1549,In_492);
xnor U2576 (N_2576,In_610,In_1036);
nor U2577 (N_2577,In_1515,In_683);
or U2578 (N_2578,In_461,In_167);
nand U2579 (N_2579,In_189,In_1866);
or U2580 (N_2580,In_916,In_1978);
nand U2581 (N_2581,In_47,In_322);
or U2582 (N_2582,In_981,In_1242);
and U2583 (N_2583,In_1143,In_599);
xor U2584 (N_2584,In_578,In_1324);
nor U2585 (N_2585,In_1616,In_666);
nor U2586 (N_2586,In_1338,In_1237);
nor U2587 (N_2587,In_1627,In_514);
nor U2588 (N_2588,In_67,In_994);
nor U2589 (N_2589,In_1540,In_829);
xnor U2590 (N_2590,In_1882,In_1614);
nor U2591 (N_2591,In_1412,In_966);
or U2592 (N_2592,In_1224,In_1187);
nand U2593 (N_2593,In_1981,In_287);
or U2594 (N_2594,In_1842,In_94);
or U2595 (N_2595,In_365,In_1280);
xnor U2596 (N_2596,In_1105,In_370);
xnor U2597 (N_2597,In_897,In_86);
nand U2598 (N_2598,In_1547,In_1517);
and U2599 (N_2599,In_1846,In_821);
nand U2600 (N_2600,In_1262,In_944);
or U2601 (N_2601,In_1359,In_263);
nor U2602 (N_2602,In_695,In_47);
or U2603 (N_2603,In_285,In_1641);
and U2604 (N_2604,In_162,In_1327);
and U2605 (N_2605,In_353,In_710);
nand U2606 (N_2606,In_196,In_1687);
nor U2607 (N_2607,In_673,In_483);
and U2608 (N_2608,In_597,In_412);
nor U2609 (N_2609,In_1599,In_1404);
or U2610 (N_2610,In_224,In_1633);
or U2611 (N_2611,In_346,In_741);
or U2612 (N_2612,In_1473,In_823);
or U2613 (N_2613,In_1229,In_264);
xnor U2614 (N_2614,In_1009,In_1475);
xor U2615 (N_2615,In_1818,In_1791);
or U2616 (N_2616,In_1015,In_81);
or U2617 (N_2617,In_1882,In_1188);
nor U2618 (N_2618,In_984,In_1321);
nor U2619 (N_2619,In_1180,In_585);
and U2620 (N_2620,In_1083,In_1283);
nand U2621 (N_2621,In_1232,In_1697);
xnor U2622 (N_2622,In_1036,In_1442);
xor U2623 (N_2623,In_1924,In_694);
nand U2624 (N_2624,In_1235,In_144);
nor U2625 (N_2625,In_873,In_907);
nor U2626 (N_2626,In_423,In_1103);
nor U2627 (N_2627,In_180,In_540);
and U2628 (N_2628,In_369,In_1613);
or U2629 (N_2629,In_688,In_1359);
xnor U2630 (N_2630,In_1008,In_1747);
nand U2631 (N_2631,In_1686,In_1766);
xnor U2632 (N_2632,In_263,In_1267);
nor U2633 (N_2633,In_609,In_541);
nor U2634 (N_2634,In_652,In_1447);
or U2635 (N_2635,In_993,In_791);
and U2636 (N_2636,In_1917,In_1315);
nor U2637 (N_2637,In_984,In_1828);
xnor U2638 (N_2638,In_1033,In_1899);
or U2639 (N_2639,In_142,In_652);
and U2640 (N_2640,In_605,In_240);
and U2641 (N_2641,In_1201,In_401);
or U2642 (N_2642,In_1646,In_170);
nand U2643 (N_2643,In_386,In_334);
and U2644 (N_2644,In_168,In_1964);
nor U2645 (N_2645,In_1320,In_1753);
and U2646 (N_2646,In_181,In_1056);
or U2647 (N_2647,In_1300,In_218);
and U2648 (N_2648,In_677,In_1980);
xor U2649 (N_2649,In_1436,In_971);
or U2650 (N_2650,In_1356,In_1600);
xnor U2651 (N_2651,In_822,In_475);
or U2652 (N_2652,In_1993,In_516);
xnor U2653 (N_2653,In_1286,In_1526);
xor U2654 (N_2654,In_1991,In_1691);
or U2655 (N_2655,In_1040,In_1253);
or U2656 (N_2656,In_1432,In_1835);
nor U2657 (N_2657,In_46,In_444);
or U2658 (N_2658,In_1449,In_486);
or U2659 (N_2659,In_485,In_145);
nand U2660 (N_2660,In_1199,In_1403);
nand U2661 (N_2661,In_1740,In_6);
or U2662 (N_2662,In_895,In_582);
nand U2663 (N_2663,In_500,In_553);
and U2664 (N_2664,In_1684,In_427);
xor U2665 (N_2665,In_1214,In_1300);
or U2666 (N_2666,In_447,In_1833);
xnor U2667 (N_2667,In_1599,In_1297);
nor U2668 (N_2668,In_259,In_413);
xnor U2669 (N_2669,In_1189,In_1952);
nor U2670 (N_2670,In_753,In_1664);
xor U2671 (N_2671,In_1914,In_1043);
nor U2672 (N_2672,In_270,In_963);
or U2673 (N_2673,In_1277,In_1557);
or U2674 (N_2674,In_95,In_794);
nand U2675 (N_2675,In_891,In_1613);
nor U2676 (N_2676,In_867,In_1287);
nand U2677 (N_2677,In_1071,In_637);
nor U2678 (N_2678,In_699,In_1246);
and U2679 (N_2679,In_1683,In_1429);
and U2680 (N_2680,In_1306,In_865);
xor U2681 (N_2681,In_890,In_532);
or U2682 (N_2682,In_1196,In_1949);
xor U2683 (N_2683,In_1214,In_1308);
xnor U2684 (N_2684,In_845,In_799);
nand U2685 (N_2685,In_1390,In_836);
nand U2686 (N_2686,In_1384,In_1638);
and U2687 (N_2687,In_929,In_561);
xnor U2688 (N_2688,In_422,In_1374);
and U2689 (N_2689,In_1192,In_1711);
nor U2690 (N_2690,In_186,In_1557);
xor U2691 (N_2691,In_79,In_244);
nor U2692 (N_2692,In_961,In_418);
nor U2693 (N_2693,In_1817,In_411);
xnor U2694 (N_2694,In_859,In_1513);
and U2695 (N_2695,In_1771,In_818);
nand U2696 (N_2696,In_981,In_503);
xnor U2697 (N_2697,In_1005,In_339);
or U2698 (N_2698,In_1768,In_1453);
and U2699 (N_2699,In_780,In_1845);
nand U2700 (N_2700,In_1032,In_551);
xnor U2701 (N_2701,In_767,In_819);
nand U2702 (N_2702,In_994,In_493);
nand U2703 (N_2703,In_1078,In_1447);
or U2704 (N_2704,In_1,In_906);
xor U2705 (N_2705,In_1643,In_1291);
and U2706 (N_2706,In_1827,In_1143);
and U2707 (N_2707,In_363,In_1898);
nor U2708 (N_2708,In_1397,In_1631);
nor U2709 (N_2709,In_1700,In_232);
or U2710 (N_2710,In_630,In_124);
or U2711 (N_2711,In_1241,In_1528);
xor U2712 (N_2712,In_1614,In_451);
xor U2713 (N_2713,In_509,In_658);
nor U2714 (N_2714,In_1060,In_1314);
xnor U2715 (N_2715,In_1652,In_748);
xor U2716 (N_2716,In_1067,In_1830);
or U2717 (N_2717,In_421,In_996);
and U2718 (N_2718,In_1410,In_335);
nor U2719 (N_2719,In_366,In_916);
or U2720 (N_2720,In_1536,In_783);
xnor U2721 (N_2721,In_1056,In_1235);
and U2722 (N_2722,In_1452,In_1791);
nand U2723 (N_2723,In_558,In_514);
nor U2724 (N_2724,In_1402,In_288);
nor U2725 (N_2725,In_1947,In_1856);
and U2726 (N_2726,In_1518,In_1707);
nor U2727 (N_2727,In_1343,In_1599);
xnor U2728 (N_2728,In_1959,In_1647);
nand U2729 (N_2729,In_517,In_162);
xnor U2730 (N_2730,In_281,In_1451);
nor U2731 (N_2731,In_241,In_52);
and U2732 (N_2732,In_1382,In_633);
and U2733 (N_2733,In_914,In_1276);
and U2734 (N_2734,In_140,In_662);
nand U2735 (N_2735,In_1607,In_603);
nand U2736 (N_2736,In_1689,In_283);
and U2737 (N_2737,In_696,In_603);
xnor U2738 (N_2738,In_1172,In_1167);
nor U2739 (N_2739,In_844,In_462);
nand U2740 (N_2740,In_979,In_1725);
nor U2741 (N_2741,In_1048,In_1448);
or U2742 (N_2742,In_1925,In_1973);
xnor U2743 (N_2743,In_1910,In_1793);
nand U2744 (N_2744,In_825,In_1235);
xor U2745 (N_2745,In_1331,In_1826);
nor U2746 (N_2746,In_262,In_448);
nand U2747 (N_2747,In_1555,In_310);
nand U2748 (N_2748,In_1288,In_379);
and U2749 (N_2749,In_106,In_370);
nand U2750 (N_2750,In_883,In_1937);
xnor U2751 (N_2751,In_446,In_10);
and U2752 (N_2752,In_1523,In_1930);
nand U2753 (N_2753,In_1669,In_1623);
and U2754 (N_2754,In_551,In_1446);
nand U2755 (N_2755,In_584,In_24);
or U2756 (N_2756,In_314,In_87);
nand U2757 (N_2757,In_1017,In_657);
or U2758 (N_2758,In_1189,In_643);
and U2759 (N_2759,In_648,In_1928);
nor U2760 (N_2760,In_420,In_1424);
nand U2761 (N_2761,In_1980,In_68);
or U2762 (N_2762,In_1283,In_1008);
and U2763 (N_2763,In_1123,In_292);
xor U2764 (N_2764,In_1450,In_1476);
nand U2765 (N_2765,In_41,In_597);
nor U2766 (N_2766,In_1628,In_1824);
xnor U2767 (N_2767,In_91,In_491);
xor U2768 (N_2768,In_1086,In_1825);
nand U2769 (N_2769,In_1653,In_64);
and U2770 (N_2770,In_43,In_1075);
nor U2771 (N_2771,In_305,In_1490);
nor U2772 (N_2772,In_1135,In_1761);
or U2773 (N_2773,In_1566,In_821);
xor U2774 (N_2774,In_1232,In_718);
xnor U2775 (N_2775,In_769,In_1761);
xnor U2776 (N_2776,In_605,In_197);
or U2777 (N_2777,In_1116,In_1579);
or U2778 (N_2778,In_1951,In_802);
xor U2779 (N_2779,In_919,In_17);
nand U2780 (N_2780,In_1684,In_520);
or U2781 (N_2781,In_1383,In_607);
nor U2782 (N_2782,In_1536,In_1574);
or U2783 (N_2783,In_1125,In_1094);
and U2784 (N_2784,In_7,In_1878);
or U2785 (N_2785,In_1876,In_1478);
nand U2786 (N_2786,In_1392,In_1149);
or U2787 (N_2787,In_816,In_1452);
xnor U2788 (N_2788,In_970,In_588);
nor U2789 (N_2789,In_194,In_1951);
xor U2790 (N_2790,In_1250,In_1114);
xnor U2791 (N_2791,In_1746,In_677);
and U2792 (N_2792,In_1175,In_1668);
and U2793 (N_2793,In_1053,In_1530);
nand U2794 (N_2794,In_1495,In_48);
or U2795 (N_2795,In_1593,In_1570);
or U2796 (N_2796,In_1824,In_1788);
xnor U2797 (N_2797,In_15,In_992);
nor U2798 (N_2798,In_1000,In_477);
and U2799 (N_2799,In_686,In_891);
nand U2800 (N_2800,In_1577,In_1071);
xor U2801 (N_2801,In_354,In_0);
and U2802 (N_2802,In_1268,In_1683);
nor U2803 (N_2803,In_1777,In_320);
and U2804 (N_2804,In_1624,In_1766);
xnor U2805 (N_2805,In_223,In_960);
or U2806 (N_2806,In_802,In_1852);
nand U2807 (N_2807,In_1737,In_528);
or U2808 (N_2808,In_828,In_1249);
nand U2809 (N_2809,In_1142,In_1149);
nor U2810 (N_2810,In_678,In_1804);
and U2811 (N_2811,In_844,In_1400);
xnor U2812 (N_2812,In_653,In_101);
nor U2813 (N_2813,In_1879,In_212);
or U2814 (N_2814,In_1656,In_274);
nand U2815 (N_2815,In_513,In_734);
and U2816 (N_2816,In_661,In_1350);
and U2817 (N_2817,In_1707,In_754);
nor U2818 (N_2818,In_179,In_903);
xnor U2819 (N_2819,In_492,In_1785);
nand U2820 (N_2820,In_637,In_1030);
nand U2821 (N_2821,In_139,In_1287);
nor U2822 (N_2822,In_1544,In_281);
nor U2823 (N_2823,In_607,In_1779);
xnor U2824 (N_2824,In_1332,In_1467);
and U2825 (N_2825,In_1569,In_421);
xnor U2826 (N_2826,In_651,In_133);
nor U2827 (N_2827,In_779,In_1312);
and U2828 (N_2828,In_1674,In_1696);
and U2829 (N_2829,In_260,In_941);
nand U2830 (N_2830,In_291,In_1860);
and U2831 (N_2831,In_48,In_985);
or U2832 (N_2832,In_1307,In_1328);
nor U2833 (N_2833,In_419,In_1222);
nor U2834 (N_2834,In_1725,In_1231);
xor U2835 (N_2835,In_761,In_760);
and U2836 (N_2836,In_832,In_1590);
and U2837 (N_2837,In_96,In_1901);
nand U2838 (N_2838,In_628,In_1330);
or U2839 (N_2839,In_92,In_1187);
xor U2840 (N_2840,In_345,In_1725);
nand U2841 (N_2841,In_993,In_542);
and U2842 (N_2842,In_1733,In_105);
xnor U2843 (N_2843,In_1609,In_1379);
nor U2844 (N_2844,In_1708,In_1474);
nor U2845 (N_2845,In_1128,In_39);
nand U2846 (N_2846,In_1944,In_194);
or U2847 (N_2847,In_49,In_967);
nand U2848 (N_2848,In_1404,In_1293);
nor U2849 (N_2849,In_1668,In_865);
and U2850 (N_2850,In_1239,In_384);
nor U2851 (N_2851,In_1521,In_1108);
and U2852 (N_2852,In_924,In_1150);
and U2853 (N_2853,In_920,In_921);
or U2854 (N_2854,In_15,In_1153);
or U2855 (N_2855,In_1036,In_1588);
nand U2856 (N_2856,In_1181,In_1633);
nand U2857 (N_2857,In_1564,In_1625);
nand U2858 (N_2858,In_1455,In_688);
and U2859 (N_2859,In_1350,In_471);
nor U2860 (N_2860,In_771,In_1305);
and U2861 (N_2861,In_1965,In_335);
xnor U2862 (N_2862,In_69,In_145);
and U2863 (N_2863,In_649,In_1601);
xnor U2864 (N_2864,In_841,In_999);
or U2865 (N_2865,In_411,In_1745);
or U2866 (N_2866,In_1321,In_1112);
xor U2867 (N_2867,In_1742,In_1700);
or U2868 (N_2868,In_1377,In_1401);
or U2869 (N_2869,In_1570,In_1949);
nand U2870 (N_2870,In_644,In_161);
nor U2871 (N_2871,In_634,In_284);
xnor U2872 (N_2872,In_247,In_768);
xnor U2873 (N_2873,In_1431,In_407);
xnor U2874 (N_2874,In_1494,In_1337);
and U2875 (N_2875,In_958,In_966);
nor U2876 (N_2876,In_593,In_764);
nand U2877 (N_2877,In_381,In_1175);
and U2878 (N_2878,In_1849,In_293);
nor U2879 (N_2879,In_44,In_1212);
nand U2880 (N_2880,In_1820,In_565);
nand U2881 (N_2881,In_1199,In_40);
or U2882 (N_2882,In_1846,In_147);
and U2883 (N_2883,In_1927,In_1779);
nand U2884 (N_2884,In_1350,In_1355);
nor U2885 (N_2885,In_1547,In_1881);
and U2886 (N_2886,In_493,In_1327);
and U2887 (N_2887,In_182,In_653);
nor U2888 (N_2888,In_1730,In_962);
xnor U2889 (N_2889,In_1390,In_793);
nand U2890 (N_2890,In_1798,In_441);
or U2891 (N_2891,In_1544,In_610);
or U2892 (N_2892,In_1062,In_464);
nor U2893 (N_2893,In_757,In_1304);
nand U2894 (N_2894,In_400,In_644);
and U2895 (N_2895,In_194,In_1205);
and U2896 (N_2896,In_441,In_828);
nand U2897 (N_2897,In_201,In_525);
or U2898 (N_2898,In_1424,In_372);
and U2899 (N_2899,In_1749,In_1423);
and U2900 (N_2900,In_1556,In_1324);
nand U2901 (N_2901,In_40,In_381);
or U2902 (N_2902,In_923,In_184);
or U2903 (N_2903,In_1141,In_23);
and U2904 (N_2904,In_672,In_481);
nor U2905 (N_2905,In_482,In_917);
and U2906 (N_2906,In_1414,In_10);
nor U2907 (N_2907,In_1250,In_307);
or U2908 (N_2908,In_182,In_1156);
nor U2909 (N_2909,In_1677,In_52);
xnor U2910 (N_2910,In_1827,In_848);
xor U2911 (N_2911,In_383,In_873);
and U2912 (N_2912,In_156,In_1100);
or U2913 (N_2913,In_1764,In_958);
nand U2914 (N_2914,In_802,In_721);
or U2915 (N_2915,In_827,In_1071);
and U2916 (N_2916,In_1249,In_1150);
xnor U2917 (N_2917,In_1229,In_1198);
or U2918 (N_2918,In_460,In_150);
nor U2919 (N_2919,In_960,In_45);
and U2920 (N_2920,In_819,In_963);
and U2921 (N_2921,In_29,In_1649);
or U2922 (N_2922,In_1501,In_30);
nand U2923 (N_2923,In_747,In_822);
nand U2924 (N_2924,In_1250,In_1989);
nand U2925 (N_2925,In_1496,In_1503);
and U2926 (N_2926,In_210,In_708);
nor U2927 (N_2927,In_348,In_1773);
or U2928 (N_2928,In_528,In_1072);
or U2929 (N_2929,In_1662,In_9);
xor U2930 (N_2930,In_525,In_1864);
or U2931 (N_2931,In_1096,In_110);
xnor U2932 (N_2932,In_270,In_1164);
or U2933 (N_2933,In_692,In_339);
or U2934 (N_2934,In_1801,In_1775);
nand U2935 (N_2935,In_518,In_746);
nand U2936 (N_2936,In_1883,In_1653);
nor U2937 (N_2937,In_25,In_1051);
and U2938 (N_2938,In_1738,In_713);
and U2939 (N_2939,In_1898,In_1878);
xnor U2940 (N_2940,In_1156,In_355);
or U2941 (N_2941,In_1983,In_79);
nand U2942 (N_2942,In_222,In_1555);
nand U2943 (N_2943,In_1693,In_279);
and U2944 (N_2944,In_1038,In_1578);
nor U2945 (N_2945,In_1833,In_1703);
nand U2946 (N_2946,In_1608,In_211);
nor U2947 (N_2947,In_988,In_1959);
nor U2948 (N_2948,In_1871,In_654);
xor U2949 (N_2949,In_1943,In_298);
nor U2950 (N_2950,In_1794,In_1336);
nand U2951 (N_2951,In_1979,In_1167);
or U2952 (N_2952,In_1151,In_367);
nor U2953 (N_2953,In_1318,In_1901);
or U2954 (N_2954,In_114,In_240);
and U2955 (N_2955,In_995,In_1108);
xor U2956 (N_2956,In_1983,In_1520);
or U2957 (N_2957,In_1576,In_944);
xor U2958 (N_2958,In_1336,In_1438);
nor U2959 (N_2959,In_308,In_1715);
or U2960 (N_2960,In_167,In_1650);
or U2961 (N_2961,In_813,In_950);
or U2962 (N_2962,In_521,In_675);
or U2963 (N_2963,In_464,In_870);
nor U2964 (N_2964,In_237,In_1731);
nand U2965 (N_2965,In_1455,In_1345);
or U2966 (N_2966,In_814,In_407);
and U2967 (N_2967,In_335,In_1911);
and U2968 (N_2968,In_766,In_1545);
or U2969 (N_2969,In_1252,In_1197);
and U2970 (N_2970,In_620,In_1357);
xnor U2971 (N_2971,In_1683,In_1998);
nor U2972 (N_2972,In_24,In_402);
and U2973 (N_2973,In_1857,In_340);
or U2974 (N_2974,In_1026,In_332);
nor U2975 (N_2975,In_1406,In_261);
and U2976 (N_2976,In_1325,In_1860);
nor U2977 (N_2977,In_890,In_705);
nand U2978 (N_2978,In_1730,In_1463);
nor U2979 (N_2979,In_950,In_185);
nor U2980 (N_2980,In_1202,In_82);
or U2981 (N_2981,In_1960,In_530);
nand U2982 (N_2982,In_1712,In_939);
xnor U2983 (N_2983,In_1577,In_1671);
and U2984 (N_2984,In_367,In_471);
or U2985 (N_2985,In_1109,In_1314);
and U2986 (N_2986,In_1463,In_613);
xor U2987 (N_2987,In_422,In_406);
or U2988 (N_2988,In_1529,In_29);
nor U2989 (N_2989,In_822,In_1115);
nor U2990 (N_2990,In_798,In_1128);
nor U2991 (N_2991,In_1810,In_1441);
and U2992 (N_2992,In_361,In_426);
and U2993 (N_2993,In_170,In_293);
and U2994 (N_2994,In_329,In_1754);
nand U2995 (N_2995,In_13,In_1579);
or U2996 (N_2996,In_871,In_662);
or U2997 (N_2997,In_786,In_276);
or U2998 (N_2998,In_203,In_1086);
and U2999 (N_2999,In_1709,In_1694);
nor U3000 (N_3000,In_1273,In_1660);
or U3001 (N_3001,In_1154,In_671);
xnor U3002 (N_3002,In_1972,In_1841);
or U3003 (N_3003,In_195,In_1931);
xnor U3004 (N_3004,In_778,In_1225);
nand U3005 (N_3005,In_1070,In_1434);
and U3006 (N_3006,In_1273,In_1008);
nor U3007 (N_3007,In_668,In_1752);
nand U3008 (N_3008,In_203,In_1893);
nor U3009 (N_3009,In_1516,In_261);
or U3010 (N_3010,In_196,In_268);
xnor U3011 (N_3011,In_351,In_1464);
or U3012 (N_3012,In_325,In_1675);
nor U3013 (N_3013,In_1827,In_1081);
and U3014 (N_3014,In_377,In_637);
or U3015 (N_3015,In_1087,In_1674);
or U3016 (N_3016,In_1804,In_403);
nor U3017 (N_3017,In_1247,In_252);
xnor U3018 (N_3018,In_1408,In_512);
nand U3019 (N_3019,In_74,In_1722);
or U3020 (N_3020,In_20,In_113);
nor U3021 (N_3021,In_33,In_861);
xnor U3022 (N_3022,In_252,In_16);
nor U3023 (N_3023,In_1759,In_1958);
or U3024 (N_3024,In_1343,In_1663);
xnor U3025 (N_3025,In_958,In_272);
nor U3026 (N_3026,In_1730,In_161);
and U3027 (N_3027,In_1834,In_1404);
nand U3028 (N_3028,In_1017,In_917);
or U3029 (N_3029,In_1460,In_1498);
nand U3030 (N_3030,In_830,In_548);
or U3031 (N_3031,In_1457,In_1598);
or U3032 (N_3032,In_31,In_200);
and U3033 (N_3033,In_1891,In_905);
and U3034 (N_3034,In_284,In_1799);
nor U3035 (N_3035,In_566,In_1241);
and U3036 (N_3036,In_1478,In_681);
xnor U3037 (N_3037,In_1458,In_7);
nor U3038 (N_3038,In_1026,In_109);
or U3039 (N_3039,In_1351,In_722);
nor U3040 (N_3040,In_1250,In_703);
or U3041 (N_3041,In_210,In_68);
or U3042 (N_3042,In_26,In_1375);
or U3043 (N_3043,In_975,In_1313);
and U3044 (N_3044,In_1218,In_1127);
nor U3045 (N_3045,In_714,In_582);
nor U3046 (N_3046,In_1125,In_1231);
nor U3047 (N_3047,In_410,In_1959);
xnor U3048 (N_3048,In_1502,In_137);
and U3049 (N_3049,In_1021,In_1738);
nand U3050 (N_3050,In_215,In_515);
or U3051 (N_3051,In_568,In_1013);
nor U3052 (N_3052,In_755,In_1703);
and U3053 (N_3053,In_1010,In_226);
xor U3054 (N_3054,In_1211,In_1186);
and U3055 (N_3055,In_1714,In_580);
xnor U3056 (N_3056,In_1178,In_1263);
and U3057 (N_3057,In_1887,In_860);
and U3058 (N_3058,In_750,In_842);
and U3059 (N_3059,In_906,In_504);
nand U3060 (N_3060,In_1120,In_1377);
nand U3061 (N_3061,In_252,In_1870);
xnor U3062 (N_3062,In_569,In_1372);
or U3063 (N_3063,In_1048,In_252);
xnor U3064 (N_3064,In_346,In_1575);
and U3065 (N_3065,In_1679,In_686);
xor U3066 (N_3066,In_291,In_956);
nor U3067 (N_3067,In_294,In_575);
and U3068 (N_3068,In_1823,In_854);
or U3069 (N_3069,In_1816,In_647);
and U3070 (N_3070,In_1065,In_381);
or U3071 (N_3071,In_1414,In_29);
nand U3072 (N_3072,In_1949,In_681);
nand U3073 (N_3073,In_15,In_833);
and U3074 (N_3074,In_228,In_1215);
nand U3075 (N_3075,In_1842,In_862);
nand U3076 (N_3076,In_350,In_178);
and U3077 (N_3077,In_1443,In_847);
xor U3078 (N_3078,In_1824,In_263);
nor U3079 (N_3079,In_1406,In_524);
nand U3080 (N_3080,In_1478,In_1235);
nor U3081 (N_3081,In_832,In_912);
and U3082 (N_3082,In_334,In_1147);
or U3083 (N_3083,In_1432,In_59);
nor U3084 (N_3084,In_247,In_92);
and U3085 (N_3085,In_1679,In_15);
or U3086 (N_3086,In_48,In_1060);
and U3087 (N_3087,In_1459,In_1810);
nand U3088 (N_3088,In_1661,In_858);
or U3089 (N_3089,In_617,In_1258);
or U3090 (N_3090,In_1406,In_1287);
nand U3091 (N_3091,In_1456,In_1522);
or U3092 (N_3092,In_1519,In_1395);
nor U3093 (N_3093,In_24,In_690);
or U3094 (N_3094,In_1352,In_1461);
nor U3095 (N_3095,In_1351,In_718);
and U3096 (N_3096,In_749,In_1145);
xnor U3097 (N_3097,In_1752,In_206);
xnor U3098 (N_3098,In_1716,In_615);
xnor U3099 (N_3099,In_1166,In_1812);
or U3100 (N_3100,In_1295,In_468);
and U3101 (N_3101,In_1701,In_1370);
nand U3102 (N_3102,In_1053,In_1174);
or U3103 (N_3103,In_301,In_616);
nand U3104 (N_3104,In_633,In_684);
nor U3105 (N_3105,In_1706,In_701);
xor U3106 (N_3106,In_946,In_832);
nand U3107 (N_3107,In_279,In_1295);
nand U3108 (N_3108,In_654,In_1858);
and U3109 (N_3109,In_1944,In_163);
nor U3110 (N_3110,In_1623,In_518);
and U3111 (N_3111,In_1500,In_602);
and U3112 (N_3112,In_1339,In_1155);
nand U3113 (N_3113,In_1865,In_117);
nand U3114 (N_3114,In_180,In_1509);
and U3115 (N_3115,In_961,In_1844);
and U3116 (N_3116,In_89,In_1064);
nand U3117 (N_3117,In_1432,In_1377);
nand U3118 (N_3118,In_1159,In_948);
or U3119 (N_3119,In_846,In_1923);
xor U3120 (N_3120,In_132,In_503);
or U3121 (N_3121,In_753,In_433);
or U3122 (N_3122,In_1699,In_603);
nand U3123 (N_3123,In_240,In_306);
nor U3124 (N_3124,In_1416,In_1621);
and U3125 (N_3125,In_999,In_471);
nor U3126 (N_3126,In_1954,In_1582);
xor U3127 (N_3127,In_1103,In_1095);
nand U3128 (N_3128,In_561,In_840);
and U3129 (N_3129,In_588,In_1057);
xnor U3130 (N_3130,In_212,In_958);
and U3131 (N_3131,In_1280,In_1070);
and U3132 (N_3132,In_1591,In_820);
nand U3133 (N_3133,In_211,In_1990);
and U3134 (N_3134,In_1619,In_38);
nand U3135 (N_3135,In_1860,In_245);
or U3136 (N_3136,In_773,In_1956);
nand U3137 (N_3137,In_1099,In_1848);
nand U3138 (N_3138,In_586,In_1477);
and U3139 (N_3139,In_384,In_881);
nand U3140 (N_3140,In_939,In_558);
or U3141 (N_3141,In_567,In_1076);
xor U3142 (N_3142,In_1867,In_1241);
nor U3143 (N_3143,In_1752,In_1227);
nor U3144 (N_3144,In_355,In_1313);
and U3145 (N_3145,In_1402,In_1126);
nor U3146 (N_3146,In_1620,In_855);
or U3147 (N_3147,In_1635,In_569);
and U3148 (N_3148,In_461,In_1978);
xnor U3149 (N_3149,In_547,In_1205);
nand U3150 (N_3150,In_733,In_770);
nand U3151 (N_3151,In_120,In_184);
nor U3152 (N_3152,In_981,In_1083);
nor U3153 (N_3153,In_707,In_566);
nor U3154 (N_3154,In_206,In_678);
nand U3155 (N_3155,In_1985,In_1275);
nand U3156 (N_3156,In_87,In_1969);
xor U3157 (N_3157,In_1366,In_499);
and U3158 (N_3158,In_1117,In_910);
nand U3159 (N_3159,In_625,In_1763);
xor U3160 (N_3160,In_23,In_622);
or U3161 (N_3161,In_775,In_900);
and U3162 (N_3162,In_708,In_1658);
xor U3163 (N_3163,In_945,In_1622);
and U3164 (N_3164,In_1895,In_717);
or U3165 (N_3165,In_1974,In_1078);
nor U3166 (N_3166,In_25,In_1788);
nor U3167 (N_3167,In_346,In_612);
xnor U3168 (N_3168,In_393,In_1250);
xnor U3169 (N_3169,In_130,In_1691);
or U3170 (N_3170,In_760,In_1554);
or U3171 (N_3171,In_20,In_1399);
or U3172 (N_3172,In_45,In_1740);
xor U3173 (N_3173,In_1645,In_60);
nand U3174 (N_3174,In_622,In_1597);
nand U3175 (N_3175,In_565,In_1494);
and U3176 (N_3176,In_1640,In_872);
xor U3177 (N_3177,In_1788,In_1517);
and U3178 (N_3178,In_501,In_1388);
or U3179 (N_3179,In_575,In_462);
nand U3180 (N_3180,In_1905,In_212);
and U3181 (N_3181,In_1271,In_316);
nand U3182 (N_3182,In_175,In_243);
nand U3183 (N_3183,In_854,In_1667);
nor U3184 (N_3184,In_1139,In_978);
or U3185 (N_3185,In_827,In_1068);
nor U3186 (N_3186,In_1608,In_1859);
or U3187 (N_3187,In_682,In_1925);
xnor U3188 (N_3188,In_1729,In_1644);
nand U3189 (N_3189,In_1998,In_881);
and U3190 (N_3190,In_1685,In_629);
or U3191 (N_3191,In_1155,In_1248);
nor U3192 (N_3192,In_1238,In_1158);
nand U3193 (N_3193,In_1875,In_1696);
nor U3194 (N_3194,In_874,In_4);
or U3195 (N_3195,In_347,In_1409);
and U3196 (N_3196,In_130,In_994);
xnor U3197 (N_3197,In_620,In_626);
nor U3198 (N_3198,In_1749,In_1834);
or U3199 (N_3199,In_1937,In_1443);
xor U3200 (N_3200,In_1527,In_1924);
xnor U3201 (N_3201,In_1379,In_893);
and U3202 (N_3202,In_1565,In_366);
xnor U3203 (N_3203,In_650,In_150);
nand U3204 (N_3204,In_1901,In_1416);
xnor U3205 (N_3205,In_1525,In_1951);
xnor U3206 (N_3206,In_1614,In_964);
nand U3207 (N_3207,In_1058,In_386);
nor U3208 (N_3208,In_371,In_1119);
xor U3209 (N_3209,In_613,In_1181);
nor U3210 (N_3210,In_205,In_1684);
or U3211 (N_3211,In_774,In_1557);
nand U3212 (N_3212,In_401,In_253);
xnor U3213 (N_3213,In_1747,In_517);
or U3214 (N_3214,In_356,In_1016);
nand U3215 (N_3215,In_1052,In_1410);
xnor U3216 (N_3216,In_1524,In_1785);
nor U3217 (N_3217,In_1811,In_1354);
or U3218 (N_3218,In_1737,In_1634);
and U3219 (N_3219,In_61,In_1211);
nor U3220 (N_3220,In_1856,In_1233);
nand U3221 (N_3221,In_683,In_708);
or U3222 (N_3222,In_1956,In_1292);
nand U3223 (N_3223,In_1558,In_755);
nand U3224 (N_3224,In_1944,In_1470);
nor U3225 (N_3225,In_90,In_546);
or U3226 (N_3226,In_568,In_1147);
nand U3227 (N_3227,In_1436,In_745);
or U3228 (N_3228,In_981,In_1320);
or U3229 (N_3229,In_1652,In_836);
nor U3230 (N_3230,In_705,In_1189);
and U3231 (N_3231,In_1448,In_1146);
and U3232 (N_3232,In_924,In_1614);
nand U3233 (N_3233,In_899,In_78);
and U3234 (N_3234,In_1535,In_1935);
xor U3235 (N_3235,In_1738,In_1391);
xnor U3236 (N_3236,In_995,In_1728);
nor U3237 (N_3237,In_752,In_1030);
or U3238 (N_3238,In_1147,In_202);
nor U3239 (N_3239,In_567,In_464);
or U3240 (N_3240,In_349,In_137);
nand U3241 (N_3241,In_376,In_1242);
nor U3242 (N_3242,In_1099,In_157);
xnor U3243 (N_3243,In_207,In_843);
xor U3244 (N_3244,In_408,In_632);
nand U3245 (N_3245,In_1615,In_1793);
nand U3246 (N_3246,In_1895,In_1677);
and U3247 (N_3247,In_642,In_1859);
xnor U3248 (N_3248,In_774,In_281);
nor U3249 (N_3249,In_1889,In_817);
nor U3250 (N_3250,In_1250,In_351);
and U3251 (N_3251,In_1795,In_958);
and U3252 (N_3252,In_349,In_148);
nand U3253 (N_3253,In_1697,In_133);
and U3254 (N_3254,In_11,In_447);
nor U3255 (N_3255,In_1477,In_1848);
nor U3256 (N_3256,In_1196,In_670);
nor U3257 (N_3257,In_1710,In_219);
or U3258 (N_3258,In_492,In_1983);
nor U3259 (N_3259,In_775,In_797);
or U3260 (N_3260,In_1562,In_1930);
nand U3261 (N_3261,In_1274,In_1697);
xnor U3262 (N_3262,In_1401,In_1898);
and U3263 (N_3263,In_868,In_902);
or U3264 (N_3264,In_1141,In_1382);
nor U3265 (N_3265,In_1059,In_1337);
nor U3266 (N_3266,In_1536,In_1771);
nor U3267 (N_3267,In_759,In_1801);
nand U3268 (N_3268,In_1169,In_617);
nor U3269 (N_3269,In_1021,In_1858);
nand U3270 (N_3270,In_1782,In_497);
nor U3271 (N_3271,In_1822,In_867);
nor U3272 (N_3272,In_187,In_1402);
xnor U3273 (N_3273,In_1123,In_6);
nor U3274 (N_3274,In_264,In_1156);
or U3275 (N_3275,In_1446,In_373);
nor U3276 (N_3276,In_1048,In_450);
nand U3277 (N_3277,In_391,In_354);
or U3278 (N_3278,In_784,In_1172);
nand U3279 (N_3279,In_1021,In_1463);
or U3280 (N_3280,In_1669,In_261);
and U3281 (N_3281,In_264,In_336);
nand U3282 (N_3282,In_70,In_43);
or U3283 (N_3283,In_914,In_1523);
or U3284 (N_3284,In_1662,In_1574);
xnor U3285 (N_3285,In_338,In_773);
xnor U3286 (N_3286,In_627,In_1530);
nand U3287 (N_3287,In_1156,In_640);
and U3288 (N_3288,In_1077,In_1416);
nand U3289 (N_3289,In_527,In_448);
nor U3290 (N_3290,In_240,In_713);
nand U3291 (N_3291,In_1411,In_254);
or U3292 (N_3292,In_898,In_1126);
nor U3293 (N_3293,In_1220,In_1621);
xnor U3294 (N_3294,In_1143,In_1692);
nor U3295 (N_3295,In_1663,In_511);
or U3296 (N_3296,In_775,In_1315);
nor U3297 (N_3297,In_1369,In_1833);
nand U3298 (N_3298,In_1710,In_695);
nand U3299 (N_3299,In_184,In_1495);
xor U3300 (N_3300,In_858,In_1636);
nor U3301 (N_3301,In_630,In_1177);
and U3302 (N_3302,In_588,In_1995);
nand U3303 (N_3303,In_1148,In_1205);
and U3304 (N_3304,In_709,In_1925);
nand U3305 (N_3305,In_872,In_585);
nand U3306 (N_3306,In_310,In_1158);
xor U3307 (N_3307,In_217,In_386);
and U3308 (N_3308,In_1994,In_1414);
xnor U3309 (N_3309,In_1583,In_1110);
and U3310 (N_3310,In_103,In_577);
nor U3311 (N_3311,In_1822,In_1955);
xnor U3312 (N_3312,In_1369,In_1953);
nor U3313 (N_3313,In_1346,In_1049);
xnor U3314 (N_3314,In_1487,In_545);
and U3315 (N_3315,In_1334,In_1819);
xnor U3316 (N_3316,In_317,In_17);
and U3317 (N_3317,In_1339,In_67);
nand U3318 (N_3318,In_1321,In_36);
or U3319 (N_3319,In_1607,In_1723);
nand U3320 (N_3320,In_1084,In_167);
xor U3321 (N_3321,In_1578,In_1235);
nand U3322 (N_3322,In_780,In_843);
or U3323 (N_3323,In_512,In_1571);
or U3324 (N_3324,In_5,In_1287);
nand U3325 (N_3325,In_1072,In_1293);
and U3326 (N_3326,In_592,In_1490);
nor U3327 (N_3327,In_334,In_1179);
or U3328 (N_3328,In_1056,In_410);
and U3329 (N_3329,In_1368,In_50);
or U3330 (N_3330,In_203,In_746);
xor U3331 (N_3331,In_1910,In_1451);
nor U3332 (N_3332,In_1127,In_623);
and U3333 (N_3333,In_1803,In_168);
xor U3334 (N_3334,In_343,In_710);
nand U3335 (N_3335,In_1565,In_1607);
nor U3336 (N_3336,In_357,In_690);
nor U3337 (N_3337,In_1448,In_92);
xor U3338 (N_3338,In_833,In_189);
nand U3339 (N_3339,In_354,In_1254);
nor U3340 (N_3340,In_505,In_113);
xnor U3341 (N_3341,In_1246,In_329);
or U3342 (N_3342,In_567,In_1726);
or U3343 (N_3343,In_1444,In_1502);
xor U3344 (N_3344,In_874,In_278);
nand U3345 (N_3345,In_412,In_172);
nor U3346 (N_3346,In_924,In_1397);
and U3347 (N_3347,In_1176,In_1781);
or U3348 (N_3348,In_1175,In_1941);
xnor U3349 (N_3349,In_1180,In_1957);
and U3350 (N_3350,In_1192,In_377);
and U3351 (N_3351,In_857,In_201);
or U3352 (N_3352,In_589,In_146);
xor U3353 (N_3353,In_1667,In_547);
and U3354 (N_3354,In_142,In_741);
or U3355 (N_3355,In_1538,In_1632);
and U3356 (N_3356,In_277,In_1541);
nand U3357 (N_3357,In_339,In_916);
nor U3358 (N_3358,In_805,In_455);
or U3359 (N_3359,In_610,In_370);
xnor U3360 (N_3360,In_197,In_193);
and U3361 (N_3361,In_8,In_970);
and U3362 (N_3362,In_1853,In_956);
nor U3363 (N_3363,In_459,In_782);
nor U3364 (N_3364,In_14,In_1511);
nor U3365 (N_3365,In_90,In_230);
nor U3366 (N_3366,In_1441,In_171);
nand U3367 (N_3367,In_164,In_169);
nand U3368 (N_3368,In_1476,In_1202);
and U3369 (N_3369,In_1077,In_1303);
xnor U3370 (N_3370,In_827,In_316);
nor U3371 (N_3371,In_1867,In_199);
xnor U3372 (N_3372,In_1771,In_1465);
or U3373 (N_3373,In_590,In_510);
nand U3374 (N_3374,In_1807,In_863);
and U3375 (N_3375,In_1797,In_194);
xor U3376 (N_3376,In_292,In_1971);
nor U3377 (N_3377,In_1478,In_685);
nor U3378 (N_3378,In_1931,In_25);
nor U3379 (N_3379,In_78,In_1469);
xor U3380 (N_3380,In_1259,In_1336);
or U3381 (N_3381,In_1758,In_1257);
nor U3382 (N_3382,In_835,In_92);
nor U3383 (N_3383,In_241,In_666);
or U3384 (N_3384,In_887,In_1964);
nand U3385 (N_3385,In_1393,In_151);
nand U3386 (N_3386,In_1123,In_140);
xnor U3387 (N_3387,In_1399,In_938);
and U3388 (N_3388,In_261,In_1028);
xnor U3389 (N_3389,In_1887,In_335);
xnor U3390 (N_3390,In_472,In_907);
nor U3391 (N_3391,In_688,In_412);
and U3392 (N_3392,In_1450,In_1565);
or U3393 (N_3393,In_26,In_1558);
nand U3394 (N_3394,In_1273,In_1450);
and U3395 (N_3395,In_1656,In_585);
xnor U3396 (N_3396,In_1804,In_1435);
or U3397 (N_3397,In_928,In_546);
nor U3398 (N_3398,In_972,In_794);
nor U3399 (N_3399,In_1197,In_866);
xnor U3400 (N_3400,In_156,In_35);
and U3401 (N_3401,In_628,In_1365);
xor U3402 (N_3402,In_1835,In_249);
or U3403 (N_3403,In_1971,In_765);
nand U3404 (N_3404,In_815,In_1597);
or U3405 (N_3405,In_517,In_1418);
nor U3406 (N_3406,In_1611,In_1260);
xor U3407 (N_3407,In_254,In_110);
and U3408 (N_3408,In_6,In_889);
xor U3409 (N_3409,In_1275,In_954);
nor U3410 (N_3410,In_535,In_912);
nand U3411 (N_3411,In_514,In_1959);
nand U3412 (N_3412,In_104,In_1819);
xnor U3413 (N_3413,In_466,In_1719);
nor U3414 (N_3414,In_1126,In_1210);
nor U3415 (N_3415,In_1943,In_1330);
or U3416 (N_3416,In_1267,In_88);
and U3417 (N_3417,In_1360,In_943);
or U3418 (N_3418,In_1101,In_141);
or U3419 (N_3419,In_1505,In_1902);
and U3420 (N_3420,In_127,In_1067);
or U3421 (N_3421,In_4,In_346);
or U3422 (N_3422,In_1787,In_866);
nand U3423 (N_3423,In_1987,In_24);
and U3424 (N_3424,In_604,In_1678);
xor U3425 (N_3425,In_1019,In_70);
xor U3426 (N_3426,In_197,In_1309);
nor U3427 (N_3427,In_1738,In_1804);
nand U3428 (N_3428,In_286,In_805);
nand U3429 (N_3429,In_923,In_727);
or U3430 (N_3430,In_71,In_1882);
nand U3431 (N_3431,In_963,In_478);
nand U3432 (N_3432,In_598,In_520);
xnor U3433 (N_3433,In_262,In_1001);
xnor U3434 (N_3434,In_609,In_432);
or U3435 (N_3435,In_349,In_378);
nand U3436 (N_3436,In_509,In_811);
and U3437 (N_3437,In_1594,In_1454);
nand U3438 (N_3438,In_49,In_526);
and U3439 (N_3439,In_759,In_1358);
nand U3440 (N_3440,In_1208,In_431);
nor U3441 (N_3441,In_890,In_1467);
nand U3442 (N_3442,In_513,In_449);
xor U3443 (N_3443,In_1750,In_1873);
nor U3444 (N_3444,In_1698,In_612);
nand U3445 (N_3445,In_683,In_194);
nand U3446 (N_3446,In_1670,In_1882);
nand U3447 (N_3447,In_1191,In_1467);
or U3448 (N_3448,In_129,In_1126);
and U3449 (N_3449,In_1557,In_582);
and U3450 (N_3450,In_1773,In_107);
nor U3451 (N_3451,In_1755,In_1017);
and U3452 (N_3452,In_1238,In_1150);
and U3453 (N_3453,In_1301,In_587);
or U3454 (N_3454,In_1282,In_399);
or U3455 (N_3455,In_393,In_95);
nand U3456 (N_3456,In_54,In_1679);
nor U3457 (N_3457,In_1545,In_1453);
nor U3458 (N_3458,In_1036,In_1147);
nand U3459 (N_3459,In_254,In_1336);
nand U3460 (N_3460,In_396,In_477);
nor U3461 (N_3461,In_1741,In_510);
nand U3462 (N_3462,In_1462,In_83);
nor U3463 (N_3463,In_606,In_455);
or U3464 (N_3464,In_1964,In_1627);
nand U3465 (N_3465,In_1409,In_711);
or U3466 (N_3466,In_1392,In_73);
xor U3467 (N_3467,In_585,In_831);
or U3468 (N_3468,In_359,In_1592);
and U3469 (N_3469,In_1183,In_1928);
xor U3470 (N_3470,In_1772,In_446);
nand U3471 (N_3471,In_1616,In_82);
nand U3472 (N_3472,In_1877,In_1191);
xor U3473 (N_3473,In_1339,In_1675);
nor U3474 (N_3474,In_330,In_1268);
or U3475 (N_3475,In_470,In_848);
nor U3476 (N_3476,In_898,In_512);
or U3477 (N_3477,In_1207,In_1002);
or U3478 (N_3478,In_634,In_1511);
and U3479 (N_3479,In_230,In_162);
and U3480 (N_3480,In_1161,In_1145);
or U3481 (N_3481,In_1494,In_1918);
xnor U3482 (N_3482,In_66,In_1323);
or U3483 (N_3483,In_356,In_1498);
nand U3484 (N_3484,In_1916,In_1357);
xnor U3485 (N_3485,In_1846,In_1205);
or U3486 (N_3486,In_617,In_65);
or U3487 (N_3487,In_1787,In_842);
nand U3488 (N_3488,In_1773,In_1054);
nand U3489 (N_3489,In_965,In_599);
and U3490 (N_3490,In_444,In_1759);
or U3491 (N_3491,In_1168,In_1865);
xor U3492 (N_3492,In_794,In_1025);
or U3493 (N_3493,In_1897,In_791);
xor U3494 (N_3494,In_1500,In_1224);
nand U3495 (N_3495,In_1953,In_982);
xnor U3496 (N_3496,In_1441,In_1786);
nand U3497 (N_3497,In_788,In_34);
nand U3498 (N_3498,In_764,In_369);
xnor U3499 (N_3499,In_1480,In_723);
and U3500 (N_3500,In_1104,In_1299);
nand U3501 (N_3501,In_1066,In_1318);
nor U3502 (N_3502,In_518,In_1730);
nor U3503 (N_3503,In_1554,In_40);
xnor U3504 (N_3504,In_1011,In_350);
and U3505 (N_3505,In_728,In_1947);
or U3506 (N_3506,In_1941,In_1136);
xor U3507 (N_3507,In_527,In_1379);
or U3508 (N_3508,In_817,In_1640);
and U3509 (N_3509,In_1901,In_54);
and U3510 (N_3510,In_1400,In_485);
nor U3511 (N_3511,In_1614,In_1424);
nor U3512 (N_3512,In_415,In_887);
nand U3513 (N_3513,In_1902,In_1771);
nand U3514 (N_3514,In_1665,In_550);
xor U3515 (N_3515,In_49,In_1638);
or U3516 (N_3516,In_1097,In_1718);
nor U3517 (N_3517,In_672,In_455);
or U3518 (N_3518,In_1338,In_636);
or U3519 (N_3519,In_592,In_1163);
nand U3520 (N_3520,In_1240,In_21);
xor U3521 (N_3521,In_1149,In_1331);
or U3522 (N_3522,In_1034,In_1986);
nor U3523 (N_3523,In_1538,In_63);
nor U3524 (N_3524,In_442,In_1893);
nand U3525 (N_3525,In_621,In_791);
xnor U3526 (N_3526,In_1911,In_392);
xnor U3527 (N_3527,In_1200,In_997);
or U3528 (N_3528,In_649,In_1989);
or U3529 (N_3529,In_697,In_1748);
xnor U3530 (N_3530,In_1043,In_561);
nand U3531 (N_3531,In_1677,In_948);
nand U3532 (N_3532,In_1013,In_830);
and U3533 (N_3533,In_413,In_1862);
and U3534 (N_3534,In_333,In_446);
and U3535 (N_3535,In_344,In_1307);
nand U3536 (N_3536,In_1265,In_963);
or U3537 (N_3537,In_1606,In_46);
xnor U3538 (N_3538,In_1280,In_1872);
xnor U3539 (N_3539,In_679,In_1656);
nand U3540 (N_3540,In_13,In_266);
or U3541 (N_3541,In_96,In_395);
or U3542 (N_3542,In_1843,In_1727);
nor U3543 (N_3543,In_903,In_1664);
nand U3544 (N_3544,In_493,In_1143);
and U3545 (N_3545,In_1158,In_482);
and U3546 (N_3546,In_1876,In_518);
and U3547 (N_3547,In_634,In_1043);
nor U3548 (N_3548,In_990,In_1795);
xor U3549 (N_3549,In_1543,In_1702);
and U3550 (N_3550,In_927,In_339);
nand U3551 (N_3551,In_1533,In_1530);
or U3552 (N_3552,In_1280,In_1389);
xnor U3553 (N_3553,In_1218,In_688);
and U3554 (N_3554,In_157,In_1869);
and U3555 (N_3555,In_1149,In_359);
nor U3556 (N_3556,In_1565,In_271);
nand U3557 (N_3557,In_898,In_1340);
nor U3558 (N_3558,In_827,In_1579);
or U3559 (N_3559,In_558,In_46);
nand U3560 (N_3560,In_251,In_413);
or U3561 (N_3561,In_1331,In_1259);
nor U3562 (N_3562,In_1590,In_1926);
nor U3563 (N_3563,In_1149,In_1232);
or U3564 (N_3564,In_1664,In_737);
and U3565 (N_3565,In_956,In_1847);
and U3566 (N_3566,In_809,In_350);
or U3567 (N_3567,In_35,In_1981);
nand U3568 (N_3568,In_626,In_387);
and U3569 (N_3569,In_123,In_1341);
or U3570 (N_3570,In_714,In_215);
xnor U3571 (N_3571,In_1145,In_122);
or U3572 (N_3572,In_481,In_1611);
and U3573 (N_3573,In_1183,In_1833);
nor U3574 (N_3574,In_1897,In_1812);
nand U3575 (N_3575,In_497,In_1629);
and U3576 (N_3576,In_1175,In_1876);
or U3577 (N_3577,In_141,In_170);
xnor U3578 (N_3578,In_1192,In_1741);
xnor U3579 (N_3579,In_310,In_1333);
and U3580 (N_3580,In_1539,In_1050);
nand U3581 (N_3581,In_1377,In_1326);
and U3582 (N_3582,In_1296,In_470);
nor U3583 (N_3583,In_1835,In_749);
nand U3584 (N_3584,In_1178,In_836);
nand U3585 (N_3585,In_900,In_315);
nand U3586 (N_3586,In_1288,In_1176);
nand U3587 (N_3587,In_1137,In_187);
nor U3588 (N_3588,In_1300,In_1971);
xnor U3589 (N_3589,In_270,In_1289);
nor U3590 (N_3590,In_32,In_489);
or U3591 (N_3591,In_1499,In_280);
or U3592 (N_3592,In_1734,In_67);
nand U3593 (N_3593,In_592,In_1763);
nand U3594 (N_3594,In_1625,In_216);
nand U3595 (N_3595,In_17,In_1581);
and U3596 (N_3596,In_1587,In_1518);
and U3597 (N_3597,In_777,In_1536);
nor U3598 (N_3598,In_51,In_1551);
nor U3599 (N_3599,In_1605,In_347);
nor U3600 (N_3600,In_1564,In_273);
nand U3601 (N_3601,In_1255,In_611);
xnor U3602 (N_3602,In_1263,In_1908);
or U3603 (N_3603,In_984,In_1801);
xnor U3604 (N_3604,In_147,In_1622);
and U3605 (N_3605,In_1130,In_1736);
or U3606 (N_3606,In_588,In_1263);
nor U3607 (N_3607,In_1376,In_1508);
nand U3608 (N_3608,In_1847,In_1074);
xor U3609 (N_3609,In_483,In_1761);
xnor U3610 (N_3610,In_1493,In_1132);
or U3611 (N_3611,In_636,In_709);
and U3612 (N_3612,In_518,In_1757);
and U3613 (N_3613,In_1731,In_1950);
nand U3614 (N_3614,In_1773,In_1102);
or U3615 (N_3615,In_1495,In_987);
nor U3616 (N_3616,In_823,In_1034);
nor U3617 (N_3617,In_773,In_361);
nand U3618 (N_3618,In_601,In_1712);
or U3619 (N_3619,In_123,In_1213);
or U3620 (N_3620,In_1528,In_834);
or U3621 (N_3621,In_151,In_890);
xnor U3622 (N_3622,In_382,In_798);
or U3623 (N_3623,In_1456,In_346);
nor U3624 (N_3624,In_190,In_1991);
nand U3625 (N_3625,In_1261,In_732);
or U3626 (N_3626,In_1692,In_1100);
xor U3627 (N_3627,In_640,In_365);
and U3628 (N_3628,In_1962,In_632);
nand U3629 (N_3629,In_1359,In_1451);
or U3630 (N_3630,In_129,In_512);
nor U3631 (N_3631,In_772,In_1894);
nand U3632 (N_3632,In_1339,In_821);
and U3633 (N_3633,In_900,In_948);
and U3634 (N_3634,In_532,In_672);
or U3635 (N_3635,In_1071,In_529);
nor U3636 (N_3636,In_1902,In_1170);
nor U3637 (N_3637,In_1947,In_1924);
nor U3638 (N_3638,In_132,In_1089);
xnor U3639 (N_3639,In_893,In_1895);
and U3640 (N_3640,In_853,In_488);
nor U3641 (N_3641,In_369,In_457);
nand U3642 (N_3642,In_1498,In_1976);
nand U3643 (N_3643,In_103,In_1999);
nor U3644 (N_3644,In_702,In_1470);
and U3645 (N_3645,In_362,In_634);
nor U3646 (N_3646,In_263,In_688);
and U3647 (N_3647,In_738,In_908);
xor U3648 (N_3648,In_1008,In_1656);
nand U3649 (N_3649,In_760,In_1520);
nor U3650 (N_3650,In_1530,In_1601);
xnor U3651 (N_3651,In_1882,In_1604);
xor U3652 (N_3652,In_1072,In_872);
or U3653 (N_3653,In_1968,In_1575);
or U3654 (N_3654,In_1839,In_304);
nand U3655 (N_3655,In_872,In_1645);
nor U3656 (N_3656,In_1279,In_1611);
nand U3657 (N_3657,In_689,In_941);
or U3658 (N_3658,In_1252,In_1951);
xnor U3659 (N_3659,In_1150,In_1320);
or U3660 (N_3660,In_624,In_1441);
xnor U3661 (N_3661,In_116,In_611);
xor U3662 (N_3662,In_310,In_1071);
or U3663 (N_3663,In_553,In_1361);
nand U3664 (N_3664,In_1158,In_1749);
nor U3665 (N_3665,In_1198,In_1261);
nor U3666 (N_3666,In_298,In_197);
nand U3667 (N_3667,In_1208,In_1560);
and U3668 (N_3668,In_1414,In_649);
or U3669 (N_3669,In_1399,In_1847);
xnor U3670 (N_3670,In_1367,In_755);
nor U3671 (N_3671,In_432,In_1598);
nand U3672 (N_3672,In_1555,In_75);
xnor U3673 (N_3673,In_754,In_69);
and U3674 (N_3674,In_780,In_1867);
and U3675 (N_3675,In_579,In_1404);
and U3676 (N_3676,In_35,In_1138);
or U3677 (N_3677,In_1167,In_13);
and U3678 (N_3678,In_1530,In_1558);
nand U3679 (N_3679,In_605,In_1434);
nor U3680 (N_3680,In_291,In_589);
nand U3681 (N_3681,In_458,In_1273);
nor U3682 (N_3682,In_80,In_1964);
or U3683 (N_3683,In_1266,In_112);
nand U3684 (N_3684,In_191,In_1738);
nor U3685 (N_3685,In_449,In_778);
and U3686 (N_3686,In_661,In_1769);
nand U3687 (N_3687,In_84,In_147);
or U3688 (N_3688,In_67,In_901);
nand U3689 (N_3689,In_1519,In_1646);
nor U3690 (N_3690,In_749,In_218);
xnor U3691 (N_3691,In_1149,In_1140);
nor U3692 (N_3692,In_427,In_1845);
nand U3693 (N_3693,In_1189,In_627);
and U3694 (N_3694,In_532,In_1921);
and U3695 (N_3695,In_1071,In_1910);
or U3696 (N_3696,In_873,In_604);
or U3697 (N_3697,In_918,In_791);
nor U3698 (N_3698,In_1029,In_749);
xor U3699 (N_3699,In_1894,In_1001);
xnor U3700 (N_3700,In_1979,In_893);
and U3701 (N_3701,In_81,In_1505);
nand U3702 (N_3702,In_1858,In_1399);
and U3703 (N_3703,In_1654,In_657);
and U3704 (N_3704,In_1668,In_1127);
xor U3705 (N_3705,In_460,In_1968);
nand U3706 (N_3706,In_87,In_36);
xor U3707 (N_3707,In_878,In_1202);
nor U3708 (N_3708,In_1741,In_513);
nor U3709 (N_3709,In_1290,In_929);
or U3710 (N_3710,In_842,In_811);
or U3711 (N_3711,In_1712,In_1558);
and U3712 (N_3712,In_1435,In_1551);
nand U3713 (N_3713,In_1781,In_722);
nand U3714 (N_3714,In_1352,In_872);
and U3715 (N_3715,In_1548,In_757);
xor U3716 (N_3716,In_1840,In_819);
or U3717 (N_3717,In_289,In_1458);
and U3718 (N_3718,In_279,In_737);
nor U3719 (N_3719,In_1541,In_1323);
nand U3720 (N_3720,In_753,In_842);
or U3721 (N_3721,In_1980,In_712);
xor U3722 (N_3722,In_1379,In_1097);
or U3723 (N_3723,In_419,In_1855);
nand U3724 (N_3724,In_938,In_1553);
or U3725 (N_3725,In_759,In_1414);
nor U3726 (N_3726,In_1334,In_340);
and U3727 (N_3727,In_300,In_945);
nor U3728 (N_3728,In_1975,In_542);
xnor U3729 (N_3729,In_1189,In_485);
nand U3730 (N_3730,In_1707,In_441);
nor U3731 (N_3731,In_1509,In_1590);
xor U3732 (N_3732,In_1197,In_708);
nor U3733 (N_3733,In_1806,In_342);
nand U3734 (N_3734,In_1079,In_1796);
and U3735 (N_3735,In_604,In_1692);
or U3736 (N_3736,In_210,In_1128);
and U3737 (N_3737,In_1153,In_1764);
and U3738 (N_3738,In_43,In_196);
xor U3739 (N_3739,In_750,In_382);
or U3740 (N_3740,In_1413,In_1283);
xnor U3741 (N_3741,In_1706,In_1257);
xnor U3742 (N_3742,In_792,In_207);
nand U3743 (N_3743,In_218,In_345);
nand U3744 (N_3744,In_1577,In_1398);
nand U3745 (N_3745,In_843,In_252);
xor U3746 (N_3746,In_1539,In_1140);
nor U3747 (N_3747,In_590,In_975);
or U3748 (N_3748,In_763,In_714);
xnor U3749 (N_3749,In_1879,In_343);
or U3750 (N_3750,In_528,In_489);
or U3751 (N_3751,In_883,In_1587);
nand U3752 (N_3752,In_985,In_719);
and U3753 (N_3753,In_21,In_1025);
xor U3754 (N_3754,In_817,In_1940);
nor U3755 (N_3755,In_113,In_1690);
or U3756 (N_3756,In_1046,In_602);
xor U3757 (N_3757,In_1532,In_1037);
nor U3758 (N_3758,In_1932,In_53);
xnor U3759 (N_3759,In_1096,In_1805);
xor U3760 (N_3760,In_185,In_1340);
or U3761 (N_3761,In_835,In_601);
and U3762 (N_3762,In_1176,In_4);
nor U3763 (N_3763,In_1921,In_1827);
xor U3764 (N_3764,In_643,In_1623);
xor U3765 (N_3765,In_716,In_1698);
xor U3766 (N_3766,In_132,In_464);
and U3767 (N_3767,In_61,In_1210);
and U3768 (N_3768,In_1906,In_1895);
and U3769 (N_3769,In_1989,In_1409);
nand U3770 (N_3770,In_530,In_212);
nor U3771 (N_3771,In_33,In_761);
nor U3772 (N_3772,In_1805,In_256);
xnor U3773 (N_3773,In_1116,In_764);
xnor U3774 (N_3774,In_1046,In_549);
xor U3775 (N_3775,In_155,In_1268);
nand U3776 (N_3776,In_351,In_1470);
and U3777 (N_3777,In_1472,In_106);
xnor U3778 (N_3778,In_1913,In_137);
nor U3779 (N_3779,In_350,In_816);
nand U3780 (N_3780,In_1501,In_1056);
nor U3781 (N_3781,In_1053,In_1316);
xnor U3782 (N_3782,In_625,In_884);
nor U3783 (N_3783,In_1032,In_475);
nand U3784 (N_3784,In_813,In_1337);
nor U3785 (N_3785,In_1315,In_696);
nand U3786 (N_3786,In_313,In_1000);
nor U3787 (N_3787,In_1932,In_1347);
nand U3788 (N_3788,In_273,In_1040);
and U3789 (N_3789,In_127,In_1024);
and U3790 (N_3790,In_1132,In_1386);
and U3791 (N_3791,In_818,In_1278);
or U3792 (N_3792,In_1506,In_1685);
or U3793 (N_3793,In_1967,In_1920);
or U3794 (N_3794,In_1718,In_725);
or U3795 (N_3795,In_1895,In_1430);
xor U3796 (N_3796,In_1369,In_956);
and U3797 (N_3797,In_485,In_429);
nand U3798 (N_3798,In_488,In_18);
nand U3799 (N_3799,In_434,In_1682);
xor U3800 (N_3800,In_27,In_349);
and U3801 (N_3801,In_323,In_303);
nand U3802 (N_3802,In_836,In_59);
nor U3803 (N_3803,In_260,In_712);
and U3804 (N_3804,In_1785,In_230);
nor U3805 (N_3805,In_1620,In_1235);
nor U3806 (N_3806,In_605,In_579);
nand U3807 (N_3807,In_854,In_365);
nand U3808 (N_3808,In_318,In_177);
xnor U3809 (N_3809,In_349,In_1356);
or U3810 (N_3810,In_757,In_278);
nand U3811 (N_3811,In_247,In_43);
nand U3812 (N_3812,In_1829,In_1818);
nand U3813 (N_3813,In_778,In_1757);
nor U3814 (N_3814,In_76,In_1939);
nand U3815 (N_3815,In_1690,In_630);
xor U3816 (N_3816,In_289,In_281);
and U3817 (N_3817,In_1276,In_738);
xnor U3818 (N_3818,In_1292,In_1742);
xor U3819 (N_3819,In_513,In_1946);
and U3820 (N_3820,In_1056,In_618);
xnor U3821 (N_3821,In_1070,In_1111);
or U3822 (N_3822,In_1222,In_1848);
or U3823 (N_3823,In_510,In_1256);
nand U3824 (N_3824,In_1537,In_1708);
and U3825 (N_3825,In_1339,In_189);
nor U3826 (N_3826,In_417,In_75);
xor U3827 (N_3827,In_1239,In_1629);
nor U3828 (N_3828,In_1252,In_1453);
and U3829 (N_3829,In_11,In_1422);
or U3830 (N_3830,In_1261,In_993);
nand U3831 (N_3831,In_445,In_1982);
nand U3832 (N_3832,In_1346,In_322);
nand U3833 (N_3833,In_392,In_425);
or U3834 (N_3834,In_1758,In_1274);
nor U3835 (N_3835,In_321,In_1211);
nor U3836 (N_3836,In_856,In_900);
or U3837 (N_3837,In_1044,In_1950);
nand U3838 (N_3838,In_1416,In_738);
and U3839 (N_3839,In_1633,In_1033);
and U3840 (N_3840,In_1378,In_737);
or U3841 (N_3841,In_787,In_303);
xor U3842 (N_3842,In_1088,In_765);
nand U3843 (N_3843,In_434,In_1923);
xor U3844 (N_3844,In_1656,In_134);
and U3845 (N_3845,In_1300,In_816);
and U3846 (N_3846,In_188,In_1192);
and U3847 (N_3847,In_552,In_720);
xor U3848 (N_3848,In_1346,In_1545);
nor U3849 (N_3849,In_1967,In_990);
and U3850 (N_3850,In_1575,In_1646);
nor U3851 (N_3851,In_1174,In_382);
nor U3852 (N_3852,In_1274,In_293);
nor U3853 (N_3853,In_1620,In_1350);
nor U3854 (N_3854,In_1023,In_1366);
xnor U3855 (N_3855,In_1031,In_1885);
xnor U3856 (N_3856,In_1689,In_829);
or U3857 (N_3857,In_579,In_632);
nor U3858 (N_3858,In_1571,In_1635);
and U3859 (N_3859,In_1528,In_1326);
xor U3860 (N_3860,In_390,In_1069);
nor U3861 (N_3861,In_1650,In_590);
and U3862 (N_3862,In_927,In_1404);
and U3863 (N_3863,In_589,In_79);
nand U3864 (N_3864,In_65,In_690);
nor U3865 (N_3865,In_547,In_1748);
xnor U3866 (N_3866,In_1328,In_632);
xnor U3867 (N_3867,In_386,In_744);
and U3868 (N_3868,In_1024,In_633);
nor U3869 (N_3869,In_158,In_1681);
nor U3870 (N_3870,In_500,In_511);
and U3871 (N_3871,In_1632,In_988);
and U3872 (N_3872,In_394,In_750);
xnor U3873 (N_3873,In_1207,In_1671);
and U3874 (N_3874,In_849,In_337);
nand U3875 (N_3875,In_1244,In_389);
xnor U3876 (N_3876,In_37,In_1581);
and U3877 (N_3877,In_1514,In_1307);
or U3878 (N_3878,In_1893,In_426);
nor U3879 (N_3879,In_1782,In_881);
xnor U3880 (N_3880,In_1291,In_1558);
and U3881 (N_3881,In_1960,In_1782);
nor U3882 (N_3882,In_526,In_77);
and U3883 (N_3883,In_1492,In_1821);
nand U3884 (N_3884,In_698,In_1236);
and U3885 (N_3885,In_1414,In_1154);
and U3886 (N_3886,In_804,In_561);
xor U3887 (N_3887,In_847,In_351);
nand U3888 (N_3888,In_1082,In_982);
or U3889 (N_3889,In_276,In_1091);
or U3890 (N_3890,In_1250,In_478);
nor U3891 (N_3891,In_142,In_562);
nor U3892 (N_3892,In_1245,In_410);
nand U3893 (N_3893,In_1279,In_1430);
nand U3894 (N_3894,In_1712,In_1821);
xnor U3895 (N_3895,In_1758,In_979);
xnor U3896 (N_3896,In_487,In_834);
or U3897 (N_3897,In_1076,In_645);
xor U3898 (N_3898,In_1482,In_1637);
and U3899 (N_3899,In_494,In_797);
and U3900 (N_3900,In_592,In_1632);
xnor U3901 (N_3901,In_1347,In_301);
nor U3902 (N_3902,In_418,In_236);
and U3903 (N_3903,In_1487,In_1321);
and U3904 (N_3904,In_454,In_435);
or U3905 (N_3905,In_183,In_1140);
nor U3906 (N_3906,In_1323,In_1737);
nor U3907 (N_3907,In_385,In_960);
and U3908 (N_3908,In_1017,In_288);
or U3909 (N_3909,In_1525,In_486);
and U3910 (N_3910,In_932,In_694);
or U3911 (N_3911,In_1299,In_1737);
and U3912 (N_3912,In_1589,In_1185);
and U3913 (N_3913,In_1823,In_1205);
nor U3914 (N_3914,In_1306,In_1812);
xnor U3915 (N_3915,In_1198,In_1202);
and U3916 (N_3916,In_713,In_642);
nor U3917 (N_3917,In_1874,In_1752);
xor U3918 (N_3918,In_166,In_862);
or U3919 (N_3919,In_890,In_1796);
and U3920 (N_3920,In_67,In_1638);
nand U3921 (N_3921,In_33,In_135);
or U3922 (N_3922,In_1092,In_1879);
xor U3923 (N_3923,In_424,In_1974);
nand U3924 (N_3924,In_977,In_915);
or U3925 (N_3925,In_1210,In_853);
or U3926 (N_3926,In_845,In_511);
nor U3927 (N_3927,In_1889,In_1241);
or U3928 (N_3928,In_1267,In_1330);
or U3929 (N_3929,In_1138,In_803);
and U3930 (N_3930,In_572,In_4);
and U3931 (N_3931,In_54,In_463);
nor U3932 (N_3932,In_210,In_1336);
nand U3933 (N_3933,In_910,In_1631);
xnor U3934 (N_3934,In_1609,In_1973);
or U3935 (N_3935,In_1895,In_1206);
xnor U3936 (N_3936,In_1345,In_1156);
nand U3937 (N_3937,In_1489,In_247);
nor U3938 (N_3938,In_466,In_260);
or U3939 (N_3939,In_1742,In_1630);
nor U3940 (N_3940,In_1553,In_1481);
nand U3941 (N_3941,In_465,In_1461);
nand U3942 (N_3942,In_1146,In_282);
nor U3943 (N_3943,In_928,In_1765);
and U3944 (N_3944,In_303,In_1746);
and U3945 (N_3945,In_74,In_1813);
or U3946 (N_3946,In_602,In_887);
xor U3947 (N_3947,In_1716,In_385);
xnor U3948 (N_3948,In_1826,In_1175);
and U3949 (N_3949,In_1544,In_592);
and U3950 (N_3950,In_1923,In_1319);
nand U3951 (N_3951,In_1664,In_1313);
and U3952 (N_3952,In_265,In_1116);
or U3953 (N_3953,In_1854,In_316);
nor U3954 (N_3954,In_471,In_1033);
nand U3955 (N_3955,In_1137,In_534);
nor U3956 (N_3956,In_1237,In_176);
or U3957 (N_3957,In_1838,In_1661);
or U3958 (N_3958,In_1286,In_1181);
or U3959 (N_3959,In_1990,In_1639);
and U3960 (N_3960,In_248,In_152);
and U3961 (N_3961,In_21,In_360);
nor U3962 (N_3962,In_427,In_666);
and U3963 (N_3963,In_1526,In_944);
nand U3964 (N_3964,In_1800,In_32);
or U3965 (N_3965,In_1015,In_1013);
nand U3966 (N_3966,In_1766,In_847);
nor U3967 (N_3967,In_228,In_776);
xor U3968 (N_3968,In_1419,In_1394);
xnor U3969 (N_3969,In_1556,In_157);
nand U3970 (N_3970,In_675,In_825);
nand U3971 (N_3971,In_1277,In_376);
or U3972 (N_3972,In_1107,In_99);
nand U3973 (N_3973,In_109,In_789);
xnor U3974 (N_3974,In_1780,In_672);
nand U3975 (N_3975,In_251,In_509);
xor U3976 (N_3976,In_181,In_865);
and U3977 (N_3977,In_192,In_1809);
nor U3978 (N_3978,In_215,In_1445);
nor U3979 (N_3979,In_933,In_219);
nor U3980 (N_3980,In_1595,In_1435);
xor U3981 (N_3981,In_593,In_1587);
nor U3982 (N_3982,In_169,In_1055);
nor U3983 (N_3983,In_1919,In_496);
nor U3984 (N_3984,In_377,In_217);
xnor U3985 (N_3985,In_851,In_1955);
nor U3986 (N_3986,In_1909,In_376);
and U3987 (N_3987,In_1575,In_1785);
or U3988 (N_3988,In_978,In_1099);
or U3989 (N_3989,In_1210,In_1517);
or U3990 (N_3990,In_648,In_1204);
or U3991 (N_3991,In_1715,In_822);
xnor U3992 (N_3992,In_93,In_906);
nand U3993 (N_3993,In_1451,In_1134);
or U3994 (N_3994,In_291,In_820);
or U3995 (N_3995,In_1269,In_1061);
and U3996 (N_3996,In_579,In_1082);
or U3997 (N_3997,In_792,In_897);
nor U3998 (N_3998,In_1817,In_1563);
xnor U3999 (N_3999,In_1531,In_181);
nor U4000 (N_4000,N_1258,N_774);
nor U4001 (N_4001,N_3667,N_3778);
nand U4002 (N_4002,N_502,N_3565);
nor U4003 (N_4003,N_33,N_3216);
nand U4004 (N_4004,N_410,N_472);
nor U4005 (N_4005,N_1814,N_1278);
xor U4006 (N_4006,N_1544,N_3397);
and U4007 (N_4007,N_3969,N_3493);
nor U4008 (N_4008,N_2051,N_955);
and U4009 (N_4009,N_2631,N_3205);
or U4010 (N_4010,N_708,N_1408);
nand U4011 (N_4011,N_2556,N_1533);
xor U4012 (N_4012,N_125,N_1262);
or U4013 (N_4013,N_1692,N_2934);
or U4014 (N_4014,N_1894,N_1630);
or U4015 (N_4015,N_1434,N_2365);
or U4016 (N_4016,N_1261,N_55);
or U4017 (N_4017,N_2148,N_3617);
or U4018 (N_4018,N_2877,N_625);
or U4019 (N_4019,N_1327,N_133);
and U4020 (N_4020,N_3152,N_1609);
or U4021 (N_4021,N_3217,N_747);
nand U4022 (N_4022,N_3151,N_2084);
xnor U4023 (N_4023,N_2081,N_2545);
xor U4024 (N_4024,N_2318,N_617);
or U4025 (N_4025,N_3320,N_1226);
and U4026 (N_4026,N_1682,N_3324);
xor U4027 (N_4027,N_2668,N_2305);
nand U4028 (N_4028,N_1077,N_819);
and U4029 (N_4029,N_2672,N_933);
nor U4030 (N_4030,N_1458,N_2978);
or U4031 (N_4031,N_1191,N_1966);
nor U4032 (N_4032,N_3743,N_233);
and U4033 (N_4033,N_2749,N_3211);
xor U4034 (N_4034,N_1013,N_1748);
xnor U4035 (N_4035,N_3361,N_911);
or U4036 (N_4036,N_1413,N_69);
and U4037 (N_4037,N_1490,N_1018);
or U4038 (N_4038,N_1197,N_3458);
and U4039 (N_4039,N_3715,N_3940);
or U4040 (N_4040,N_1494,N_446);
xnor U4041 (N_4041,N_2239,N_1691);
nor U4042 (N_4042,N_3212,N_3654);
and U4043 (N_4043,N_3054,N_1329);
nand U4044 (N_4044,N_2953,N_2753);
nand U4045 (N_4045,N_3418,N_3358);
and U4046 (N_4046,N_1569,N_977);
or U4047 (N_4047,N_2751,N_1834);
nor U4048 (N_4048,N_713,N_3670);
and U4049 (N_4049,N_374,N_902);
nor U4050 (N_4050,N_2984,N_2251);
nor U4051 (N_4051,N_2093,N_1319);
nor U4052 (N_4052,N_354,N_2769);
and U4053 (N_4053,N_2873,N_1650);
xnor U4054 (N_4054,N_3228,N_208);
and U4055 (N_4055,N_3231,N_797);
nor U4056 (N_4056,N_1656,N_287);
and U4057 (N_4057,N_3428,N_2530);
xor U4058 (N_4058,N_1613,N_1629);
nand U4059 (N_4059,N_2023,N_3705);
and U4060 (N_4060,N_1657,N_905);
and U4061 (N_4061,N_3184,N_749);
xnor U4062 (N_4062,N_147,N_3120);
xnor U4063 (N_4063,N_3407,N_2967);
and U4064 (N_4064,N_82,N_3198);
xor U4065 (N_4065,N_79,N_3197);
nor U4066 (N_4066,N_2332,N_1167);
xnor U4067 (N_4067,N_3094,N_3836);
nor U4068 (N_4068,N_2796,N_2308);
and U4069 (N_4069,N_3804,N_1549);
or U4070 (N_4070,N_2888,N_2536);
nor U4071 (N_4071,N_1610,N_1139);
xor U4072 (N_4072,N_3948,N_1688);
nor U4073 (N_4073,N_1133,N_919);
xor U4074 (N_4074,N_1140,N_3663);
or U4075 (N_4075,N_1425,N_2193);
and U4076 (N_4076,N_2882,N_135);
nand U4077 (N_4077,N_1819,N_636);
nand U4078 (N_4078,N_1782,N_1791);
and U4079 (N_4079,N_1285,N_2198);
xnor U4080 (N_4080,N_1833,N_2259);
nor U4081 (N_4081,N_3404,N_2386);
nand U4082 (N_4082,N_3411,N_2552);
and U4083 (N_4083,N_1385,N_1045);
xnor U4084 (N_4084,N_3134,N_63);
xor U4085 (N_4085,N_3262,N_2976);
or U4086 (N_4086,N_3208,N_2541);
or U4087 (N_4087,N_3082,N_2376);
and U4088 (N_4088,N_859,N_1753);
or U4089 (N_4089,N_3636,N_3895);
or U4090 (N_4090,N_3625,N_1824);
xor U4091 (N_4091,N_1546,N_1811);
nor U4092 (N_4092,N_165,N_1070);
and U4093 (N_4093,N_3306,N_671);
and U4094 (N_4094,N_1214,N_3430);
nor U4095 (N_4095,N_2435,N_1918);
or U4096 (N_4096,N_530,N_1469);
nand U4097 (N_4097,N_909,N_3131);
nor U4098 (N_4098,N_3371,N_2200);
xor U4099 (N_4099,N_1525,N_112);
nand U4100 (N_4100,N_3629,N_763);
xor U4101 (N_4101,N_3766,N_1476);
or U4102 (N_4102,N_2917,N_3147);
nand U4103 (N_4103,N_3317,N_200);
and U4104 (N_4104,N_1574,N_696);
or U4105 (N_4105,N_101,N_3427);
or U4106 (N_4106,N_1522,N_2633);
or U4107 (N_4107,N_407,N_2923);
nor U4108 (N_4108,N_3750,N_3027);
and U4109 (N_4109,N_3635,N_1155);
nand U4110 (N_4110,N_898,N_2272);
nor U4111 (N_4111,N_3410,N_3020);
and U4112 (N_4112,N_510,N_2744);
and U4113 (N_4113,N_3513,N_3392);
nand U4114 (N_4114,N_1798,N_3535);
xor U4115 (N_4115,N_3708,N_303);
or U4116 (N_4116,N_1230,N_2273);
and U4117 (N_4117,N_356,N_1851);
nor U4118 (N_4118,N_2288,N_2129);
xnor U4119 (N_4119,N_958,N_3713);
or U4120 (N_4120,N_362,N_3100);
nor U4121 (N_4121,N_2210,N_569);
and U4122 (N_4122,N_3751,N_3843);
nand U4123 (N_4123,N_1963,N_3105);
nand U4124 (N_4124,N_2643,N_1412);
nor U4125 (N_4125,N_1830,N_2723);
nand U4126 (N_4126,N_1154,N_2721);
xor U4127 (N_4127,N_3898,N_851);
and U4128 (N_4128,N_1930,N_3716);
nor U4129 (N_4129,N_1721,N_499);
nand U4130 (N_4130,N_3383,N_2014);
xnor U4131 (N_4131,N_2295,N_3239);
nand U4132 (N_4132,N_3913,N_2845);
xnor U4133 (N_4133,N_2403,N_2596);
nand U4134 (N_4134,N_2207,N_450);
and U4135 (N_4135,N_2508,N_3987);
nor U4136 (N_4136,N_326,N_2848);
nand U4137 (N_4137,N_325,N_3732);
nor U4138 (N_4138,N_3167,N_2422);
xnor U4139 (N_4139,N_686,N_3219);
nor U4140 (N_4140,N_2881,N_3788);
or U4141 (N_4141,N_1209,N_3976);
or U4142 (N_4142,N_2825,N_1663);
nand U4143 (N_4143,N_3112,N_2851);
nor U4144 (N_4144,N_940,N_2670);
nor U4145 (N_4145,N_3059,N_1792);
and U4146 (N_4146,N_244,N_2526);
and U4147 (N_4147,N_3592,N_1173);
nand U4148 (N_4148,N_1111,N_2886);
nor U4149 (N_4149,N_3735,N_1503);
xor U4150 (N_4150,N_861,N_2082);
and U4151 (N_4151,N_2745,N_787);
and U4152 (N_4152,N_280,N_2489);
xnor U4153 (N_4153,N_1388,N_3793);
and U4154 (N_4154,N_2045,N_3921);
or U4155 (N_4155,N_1607,N_163);
and U4156 (N_4156,N_2918,N_1293);
nor U4157 (N_4157,N_1994,N_3050);
or U4158 (N_4158,N_3539,N_2528);
or U4159 (N_4159,N_2019,N_2074);
nor U4160 (N_4160,N_845,N_1407);
or U4161 (N_4161,N_1182,N_2035);
and U4162 (N_4162,N_1562,N_3156);
and U4163 (N_4163,N_2806,N_2163);
nor U4164 (N_4164,N_990,N_2216);
and U4165 (N_4165,N_3482,N_17);
xnor U4166 (N_4166,N_888,N_3305);
xnor U4167 (N_4167,N_559,N_735);
nor U4168 (N_4168,N_150,N_552);
or U4169 (N_4169,N_1499,N_2680);
nor U4170 (N_4170,N_2218,N_2725);
and U4171 (N_4171,N_1882,N_2361);
xor U4172 (N_4172,N_1436,N_3259);
xnor U4173 (N_4173,N_1342,N_2159);
xnor U4174 (N_4174,N_3160,N_1703);
nand U4175 (N_4175,N_3808,N_842);
xnor U4176 (N_4176,N_341,N_1829);
nand U4177 (N_4177,N_1428,N_433);
and U4178 (N_4178,N_2805,N_2482);
and U4179 (N_4179,N_995,N_3419);
nand U4180 (N_4180,N_1177,N_261);
nor U4181 (N_4181,N_1821,N_0);
nand U4182 (N_4182,N_1697,N_3164);
nand U4183 (N_4183,N_1588,N_1987);
xor U4184 (N_4184,N_1892,N_3562);
or U4185 (N_4185,N_3273,N_75);
nand U4186 (N_4186,N_3462,N_871);
and U4187 (N_4187,N_781,N_1598);
xor U4188 (N_4188,N_914,N_2326);
and U4189 (N_4189,N_3318,N_1913);
nand U4190 (N_4190,N_247,N_179);
and U4191 (N_4191,N_1492,N_1374);
nor U4192 (N_4192,N_3333,N_85);
and U4193 (N_4193,N_299,N_1570);
nand U4194 (N_4194,N_1799,N_1803);
nand U4195 (N_4195,N_293,N_1314);
xnor U4196 (N_4196,N_3832,N_2590);
xor U4197 (N_4197,N_1034,N_382);
or U4198 (N_4198,N_3201,N_1776);
nor U4199 (N_4199,N_1861,N_2184);
or U4200 (N_4200,N_2775,N_635);
and U4201 (N_4201,N_3353,N_1279);
xor U4202 (N_4202,N_1487,N_2060);
nand U4203 (N_4203,N_1781,N_3543);
nand U4204 (N_4204,N_3580,N_1253);
and U4205 (N_4205,N_656,N_222);
and U4206 (N_4206,N_2158,N_1090);
xor U4207 (N_4207,N_191,N_1482);
or U4208 (N_4208,N_2327,N_3557);
or U4209 (N_4209,N_1135,N_1180);
or U4210 (N_4210,N_334,N_2230);
or U4211 (N_4211,N_3450,N_2108);
nand U4212 (N_4212,N_1466,N_3017);
nand U4213 (N_4213,N_3331,N_223);
nand U4214 (N_4214,N_512,N_1835);
or U4215 (N_4215,N_3719,N_1175);
or U4216 (N_4216,N_77,N_115);
xnor U4217 (N_4217,N_3608,N_623);
or U4218 (N_4218,N_295,N_3727);
nor U4219 (N_4219,N_1687,N_1176);
nand U4220 (N_4220,N_306,N_887);
and U4221 (N_4221,N_3413,N_1681);
or U4222 (N_4222,N_3678,N_639);
nor U4223 (N_4223,N_3246,N_1865);
nor U4224 (N_4224,N_3780,N_1827);
nor U4225 (N_4225,N_3453,N_1631);
nor U4226 (N_4226,N_2889,N_22);
or U4227 (N_4227,N_132,N_2286);
and U4228 (N_4228,N_2064,N_363);
xnor U4229 (N_4229,N_1386,N_1148);
nand U4230 (N_4230,N_732,N_941);
nand U4231 (N_4231,N_3126,N_3623);
xnor U4232 (N_4232,N_2503,N_2062);
and U4233 (N_4233,N_2756,N_691);
xor U4234 (N_4234,N_2462,N_2302);
nand U4235 (N_4235,N_335,N_3146);
nor U4236 (N_4236,N_3871,N_43);
and U4237 (N_4237,N_1675,N_3309);
or U4238 (N_4238,N_2950,N_3800);
xor U4239 (N_4239,N_169,N_1920);
nor U4240 (N_4240,N_3174,N_2419);
xnor U4241 (N_4241,N_858,N_1505);
nor U4242 (N_4242,N_3267,N_3589);
nor U4243 (N_4243,N_1537,N_2257);
and U4244 (N_4244,N_2557,N_2479);
and U4245 (N_4245,N_644,N_3442);
nor U4246 (N_4246,N_56,N_3758);
nor U4247 (N_4247,N_3892,N_726);
or U4248 (N_4248,N_3887,N_586);
nor U4249 (N_4249,N_3400,N_1601);
and U4250 (N_4250,N_2319,N_29);
and U4251 (N_4251,N_1310,N_3631);
or U4252 (N_4252,N_28,N_3188);
nor U4253 (N_4253,N_2565,N_2496);
and U4254 (N_4254,N_767,N_2592);
nand U4255 (N_4255,N_3953,N_2451);
or U4256 (N_4256,N_2122,N_703);
nand U4257 (N_4257,N_2088,N_4);
xnor U4258 (N_4258,N_3022,N_641);
or U4259 (N_4259,N_2339,N_2870);
nand U4260 (N_4260,N_2766,N_2442);
and U4261 (N_4261,N_1216,N_1766);
xor U4262 (N_4262,N_3823,N_1001);
xnor U4263 (N_4263,N_1379,N_2811);
nand U4264 (N_4264,N_777,N_1985);
or U4265 (N_4265,N_631,N_1308);
or U4266 (N_4266,N_2788,N_203);
xor U4267 (N_4267,N_113,N_252);
xor U4268 (N_4268,N_3690,N_322);
nand U4269 (N_4269,N_2363,N_606);
and U4270 (N_4270,N_579,N_1528);
or U4271 (N_4271,N_1041,N_221);
and U4272 (N_4272,N_2394,N_406);
or U4273 (N_4273,N_1283,N_849);
and U4274 (N_4274,N_2875,N_1671);
xor U4275 (N_4275,N_1694,N_1243);
nand U4276 (N_4276,N_177,N_156);
xor U4277 (N_4277,N_725,N_2591);
nor U4278 (N_4278,N_2585,N_378);
or U4279 (N_4279,N_3393,N_2812);
and U4280 (N_4280,N_294,N_3399);
and U4281 (N_4281,N_3686,N_2097);
xor U4282 (N_4282,N_1473,N_336);
nor U4283 (N_4283,N_3384,N_3776);
or U4284 (N_4284,N_1967,N_1934);
nand U4285 (N_4285,N_2733,N_3257);
and U4286 (N_4286,N_2347,N_3103);
and U4287 (N_4287,N_3660,N_3598);
and U4288 (N_4288,N_1897,N_442);
xor U4289 (N_4289,N_3834,N_1089);
xor U4290 (N_4290,N_3956,N_3840);
or U4291 (N_4291,N_2427,N_1107);
or U4292 (N_4292,N_2258,N_557);
and U4293 (N_4293,N_2157,N_1165);
and U4294 (N_4294,N_3612,N_2913);
xor U4295 (N_4295,N_218,N_1925);
xnor U4296 (N_4296,N_2377,N_2550);
nand U4297 (N_4297,N_690,N_575);
nor U4298 (N_4298,N_1625,N_2119);
nor U4299 (N_4299,N_3471,N_833);
nor U4300 (N_4300,N_11,N_722);
nor U4301 (N_4301,N_21,N_276);
nand U4302 (N_4302,N_1936,N_1659);
nand U4303 (N_4303,N_360,N_188);
and U4304 (N_4304,N_3559,N_1204);
and U4305 (N_4305,N_1411,N_3073);
or U4306 (N_4306,N_823,N_471);
xor U4307 (N_4307,N_3518,N_1893);
nor U4308 (N_4308,N_122,N_3172);
xnor U4309 (N_4309,N_2666,N_267);
or U4310 (N_4310,N_2385,N_2003);
and U4311 (N_4311,N_1995,N_2411);
nand U4312 (N_4312,N_1723,N_3772);
nor U4313 (N_4313,N_2563,N_669);
nor U4314 (N_4314,N_2267,N_1354);
nand U4315 (N_4315,N_467,N_61);
or U4316 (N_4316,N_1905,N_137);
or U4317 (N_4317,N_707,N_2801);
xor U4318 (N_4318,N_2675,N_1756);
or U4319 (N_4319,N_3611,N_146);
xnor U4320 (N_4320,N_681,N_2697);
xor U4321 (N_4321,N_3524,N_3817);
xnor U4322 (N_4322,N_2543,N_2215);
xnor U4323 (N_4323,N_364,N_680);
or U4324 (N_4324,N_3724,N_477);
nor U4325 (N_4325,N_3304,N_1514);
or U4326 (N_4326,N_3468,N_2842);
nand U4327 (N_4327,N_424,N_2414);
or U4328 (N_4328,N_3764,N_1326);
nand U4329 (N_4329,N_899,N_3047);
or U4330 (N_4330,N_498,N_3374);
nor U4331 (N_4331,N_128,N_2860);
or U4332 (N_4332,N_1933,N_3498);
xnor U4333 (N_4333,N_2219,N_3214);
nor U4334 (N_4334,N_331,N_1431);
nor U4335 (N_4335,N_1576,N_3820);
xnor U4336 (N_4336,N_1768,N_1836);
nand U4337 (N_4337,N_2857,N_1758);
xor U4338 (N_4338,N_3517,N_744);
or U4339 (N_4339,N_3421,N_1347);
xnor U4340 (N_4340,N_1406,N_102);
or U4341 (N_4341,N_1304,N_996);
nand U4342 (N_4342,N_2914,N_952);
or U4343 (N_4343,N_185,N_3789);
or U4344 (N_4344,N_2507,N_1120);
or U4345 (N_4345,N_1048,N_49);
xnor U4346 (N_4346,N_574,N_2061);
or U4347 (N_4347,N_3546,N_870);
xnor U4348 (N_4348,N_1516,N_2448);
and U4349 (N_4349,N_2588,N_3600);
nor U4350 (N_4350,N_922,N_3522);
xnor U4351 (N_4351,N_1668,N_3978);
xor U4352 (N_4352,N_2819,N_1126);
xor U4353 (N_4353,N_1738,N_422);
xor U4354 (N_4354,N_3263,N_313);
or U4355 (N_4355,N_1188,N_2167);
nor U4356 (N_4356,N_1886,N_1825);
or U4357 (N_4357,N_1160,N_3396);
nand U4358 (N_4358,N_2620,N_3348);
and U4359 (N_4359,N_1251,N_2348);
and U4360 (N_4360,N_3191,N_609);
nor U4361 (N_4361,N_3124,N_1423);
nand U4362 (N_4362,N_1853,N_3098);
or U4363 (N_4363,N_1566,N_994);
nor U4364 (N_4364,N_1166,N_2364);
nor U4365 (N_4365,N_219,N_3655);
xnor U4366 (N_4366,N_2760,N_220);
nor U4367 (N_4367,N_1193,N_1683);
or U4368 (N_4368,N_3158,N_3253);
and U4369 (N_4369,N_3376,N_2335);
xor U4370 (N_4370,N_1497,N_1854);
xor U4371 (N_4371,N_1426,N_2637);
nand U4372 (N_4372,N_3283,N_3484);
nor U4373 (N_4373,N_2855,N_2206);
nand U4374 (N_4374,N_3143,N_1396);
nor U4375 (N_4375,N_2424,N_3473);
nor U4376 (N_4376,N_2279,N_1750);
and U4377 (N_4377,N_3029,N_3541);
nand U4378 (N_4378,N_1672,N_799);
nand U4379 (N_4379,N_663,N_2576);
or U4380 (N_4380,N_436,N_1389);
nand U4381 (N_4381,N_2384,N_3662);
or U4382 (N_4382,N_2520,N_330);
or U4383 (N_4383,N_2228,N_1270);
or U4384 (N_4384,N_1628,N_3351);
and U4385 (N_4385,N_1937,N_1390);
or U4386 (N_4386,N_3986,N_2433);
xnor U4387 (N_4387,N_3960,N_1344);
and U4388 (N_4388,N_1444,N_20);
xnor U4389 (N_4389,N_1660,N_3099);
nor U4390 (N_4390,N_3431,N_655);
and U4391 (N_4391,N_2030,N_80);
xor U4392 (N_4392,N_2781,N_1580);
nor U4393 (N_4393,N_3704,N_684);
xnor U4394 (N_4394,N_494,N_2765);
xnor U4395 (N_4395,N_3274,N_3053);
or U4396 (N_4396,N_1540,N_2774);
and U4397 (N_4397,N_1375,N_1059);
nand U4398 (N_4398,N_3616,N_2583);
and U4399 (N_4399,N_1478,N_1759);
xnor U4400 (N_4400,N_965,N_2907);
or U4401 (N_4401,N_2401,N_1032);
nand U4402 (N_4402,N_1929,N_534);
and U4403 (N_4403,N_1075,N_26);
or U4404 (N_4404,N_3774,N_2007);
nor U4405 (N_4405,N_2623,N_3312);
xor U4406 (N_4406,N_803,N_3512);
nand U4407 (N_4407,N_3994,N_3563);
xor U4408 (N_4408,N_2366,N_235);
nand U4409 (N_4409,N_1552,N_1597);
and U4410 (N_4410,N_3307,N_412);
xnor U4411 (N_4411,N_2768,N_3862);
and U4412 (N_4412,N_1856,N_3596);
nand U4413 (N_4413,N_1938,N_3824);
nand U4414 (N_4414,N_2574,N_699);
and U4415 (N_4415,N_496,N_760);
xor U4416 (N_4416,N_2821,N_3116);
nand U4417 (N_4417,N_1713,N_1662);
or U4418 (N_4418,N_2771,N_1736);
and U4419 (N_4419,N_2400,N_558);
or U4420 (N_4420,N_2573,N_3092);
nor U4421 (N_4421,N_988,N_66);
and U4422 (N_4422,N_1764,N_3388);
and U4423 (N_4423,N_2911,N_1394);
nor U4424 (N_4424,N_3221,N_1037);
or U4425 (N_4425,N_956,N_2936);
xnor U4426 (N_4426,N_3526,N_3671);
xnor U4427 (N_4427,N_2296,N_2440);
and U4428 (N_4428,N_525,N_91);
nand U4429 (N_4429,N_3437,N_1169);
and U4430 (N_4430,N_1108,N_3051);
or U4431 (N_4431,N_1383,N_2455);
xor U4432 (N_4432,N_3163,N_2659);
xor U4433 (N_4433,N_2264,N_2430);
or U4434 (N_4434,N_3213,N_184);
or U4435 (N_4435,N_2040,N_194);
and U4436 (N_4436,N_1666,N_342);
xor U4437 (N_4437,N_3108,N_3919);
and U4438 (N_4438,N_1067,N_167);
xnor U4439 (N_4439,N_2867,N_2201);
and U4440 (N_4440,N_127,N_3298);
or U4441 (N_4441,N_3679,N_2194);
xor U4442 (N_4442,N_1454,N_1368);
and U4443 (N_4443,N_1363,N_1415);
or U4444 (N_4444,N_3155,N_2195);
nand U4445 (N_4445,N_2260,N_482);
or U4446 (N_4446,N_1890,N_1735);
nor U4447 (N_4447,N_843,N_1612);
nand U4448 (N_4448,N_3545,N_480);
xor U4449 (N_4449,N_3270,N_2982);
nor U4450 (N_4450,N_3326,N_3902);
nand U4451 (N_4451,N_3136,N_3503);
and U4452 (N_4452,N_1286,N_1360);
nand U4453 (N_4453,N_1266,N_3576);
and U4454 (N_4454,N_3752,N_1062);
xor U4455 (N_4455,N_2485,N_2208);
nand U4456 (N_4456,N_1130,N_1677);
xnor U4457 (N_4457,N_3756,N_401);
xnor U4458 (N_4458,N_1332,N_1084);
or U4459 (N_4459,N_1639,N_3779);
nor U4460 (N_4460,N_969,N_1026);
and U4461 (N_4461,N_2963,N_1489);
nand U4462 (N_4462,N_1584,N_90);
nor U4463 (N_4463,N_462,N_3390);
xnor U4464 (N_4464,N_3579,N_2977);
nand U4465 (N_4465,N_1378,N_3327);
or U4466 (N_4466,N_3173,N_1875);
xor U4467 (N_4467,N_216,N_1618);
xnor U4468 (N_4468,N_1437,N_1777);
nand U4469 (N_4469,N_1008,N_739);
xor U4470 (N_4470,N_3033,N_798);
and U4471 (N_4471,N_415,N_2981);
xnor U4472 (N_4472,N_2933,N_1634);
nand U4473 (N_4473,N_2057,N_3803);
or U4474 (N_4474,N_1299,N_978);
and U4475 (N_4475,N_3060,N_3982);
or U4476 (N_4476,N_1156,N_3499);
nand U4477 (N_4477,N_3179,N_3865);
xor U4478 (N_4478,N_1288,N_1241);
or U4479 (N_4479,N_1734,N_474);
nand U4480 (N_4480,N_923,N_3313);
xnor U4481 (N_4481,N_2992,N_1031);
or U4482 (N_4482,N_1195,N_2227);
or U4483 (N_4483,N_2307,N_371);
and U4484 (N_4484,N_2010,N_879);
nand U4485 (N_4485,N_913,N_2458);
nor U4486 (N_4486,N_3918,N_3627);
or U4487 (N_4487,N_3609,N_2669);
nand U4488 (N_4488,N_2090,N_1701);
xor U4489 (N_4489,N_1158,N_1029);
or U4490 (N_4490,N_2454,N_592);
or U4491 (N_4491,N_867,N_3115);
nor U4492 (N_4492,N_2738,N_2237);
nor U4493 (N_4493,N_3577,N_1947);
nand U4494 (N_4494,N_761,N_1187);
or U4495 (N_4495,N_1124,N_1442);
nand U4496 (N_4496,N_1542,N_2399);
or U4497 (N_4497,N_3220,N_3012);
xnor U4498 (N_4498,N_1318,N_3614);
xnor U4499 (N_4499,N_2612,N_2252);
nand U4500 (N_4500,N_1265,N_3755);
or U4501 (N_4501,N_3447,N_3242);
or U4502 (N_4502,N_2416,N_142);
xnor U4503 (N_4503,N_1112,N_1100);
and U4504 (N_4504,N_328,N_3692);
and U4505 (N_4505,N_3202,N_1742);
xor U4506 (N_4506,N_3300,N_2656);
or U4507 (N_4507,N_893,N_3729);
xor U4508 (N_4508,N_1577,N_672);
nand U4509 (N_4509,N_591,N_1560);
and U4510 (N_4510,N_14,N_506);
or U4511 (N_4511,N_1506,N_2816);
or U4512 (N_4512,N_2047,N_966);
or U4513 (N_4513,N_2728,N_2789);
nor U4514 (N_4514,N_2429,N_3068);
and U4515 (N_4515,N_2406,N_3833);
and U4516 (N_4516,N_1706,N_1194);
or U4517 (N_4517,N_3276,N_775);
or U4518 (N_4518,N_3859,N_1427);
and U4519 (N_4519,N_2931,N_3448);
nor U4520 (N_4520,N_685,N_434);
xor U4521 (N_4521,N_944,N_1535);
xor U4522 (N_4522,N_370,N_2648);
xnor U4523 (N_4523,N_417,N_36);
and U4524 (N_4524,N_349,N_3434);
and U4525 (N_4525,N_2268,N_963);
nand U4526 (N_4526,N_2453,N_1356);
nand U4527 (N_4527,N_613,N_1903);
nand U4528 (N_4528,N_2034,N_3903);
nor U4529 (N_4529,N_2872,N_857);
nand U4530 (N_4530,N_62,N_1794);
and U4531 (N_4531,N_957,N_2730);
xnor U4532 (N_4532,N_1030,N_3868);
and U4533 (N_4533,N_3839,N_2256);
xor U4534 (N_4534,N_430,N_2959);
nand U4535 (N_4535,N_527,N_2311);
nor U4536 (N_4536,N_153,N_201);
or U4537 (N_4537,N_3784,N_126);
nand U4538 (N_4538,N_3284,N_2436);
and U4539 (N_4539,N_1039,N_862);
or U4540 (N_4540,N_2048,N_1295);
xnor U4541 (N_4541,N_637,N_1003);
xor U4542 (N_4542,N_1445,N_2473);
nand U4543 (N_4543,N_2055,N_3821);
xnor U4544 (N_4544,N_243,N_664);
or U4545 (N_4545,N_3561,N_246);
xnor U4546 (N_4546,N_1954,N_3402);
nor U4547 (N_4547,N_910,N_3794);
nor U4548 (N_4548,N_3177,N_3159);
and U4549 (N_4549,N_3486,N_756);
and U4550 (N_4550,N_3377,N_2679);
and U4551 (N_4551,N_388,N_514);
nand U4552 (N_4552,N_2076,N_3718);
nand U4553 (N_4553,N_1483,N_2741);
nor U4554 (N_4554,N_174,N_2874);
nor U4555 (N_4555,N_1060,N_1838);
or U4556 (N_4556,N_214,N_738);
and U4557 (N_4557,N_3538,N_1885);
and U4558 (N_4558,N_423,N_1449);
nor U4559 (N_4559,N_3429,N_3079);
or U4560 (N_4560,N_3008,N_3016);
and U4561 (N_4561,N_3980,N_2232);
nand U4562 (N_4562,N_3785,N_2940);
nand U4563 (N_4563,N_3153,N_694);
nand U4564 (N_4564,N_3796,N_2951);
or U4565 (N_4565,N_2569,N_493);
and U4566 (N_4566,N_3165,N_1719);
nor U4567 (N_4567,N_1145,N_1218);
or U4568 (N_4568,N_3961,N_1098);
nand U4569 (N_4569,N_524,N_392);
xnor U4570 (N_4570,N_2336,N_1136);
xor U4571 (N_4571,N_1769,N_2235);
and U4572 (N_4572,N_673,N_773);
nand U4573 (N_4573,N_307,N_3409);
or U4574 (N_4574,N_542,N_3255);
or U4575 (N_4575,N_1235,N_724);
nor U4576 (N_4576,N_2126,N_2486);
and U4577 (N_4577,N_2107,N_2478);
or U4578 (N_4578,N_1440,N_1648);
and U4579 (N_4579,N_3771,N_297);
or U4580 (N_4580,N_1009,N_3911);
nand U4581 (N_4581,N_2001,N_3040);
and U4582 (N_4582,N_2375,N_1446);
and U4583 (N_4583,N_587,N_2171);
nand U4584 (N_4584,N_543,N_266);
or U4585 (N_4585,N_379,N_743);
nor U4586 (N_4586,N_3835,N_1786);
xnor U4587 (N_4587,N_3977,N_961);
nand U4588 (N_4588,N_640,N_2147);
nand U4589 (N_4589,N_3292,N_1460);
nor U4590 (N_4590,N_1870,N_1614);
and U4591 (N_4591,N_523,N_40);
xor U4592 (N_4592,N_2098,N_894);
and U4593 (N_4593,N_2645,N_2542);
nand U4594 (N_4594,N_2009,N_2640);
and U4595 (N_4595,N_3028,N_187);
or U4596 (N_4596,N_350,N_13);
or U4597 (N_4597,N_316,N_3367);
or U4598 (N_4598,N_1887,N_864);
or U4599 (N_4599,N_1232,N_1474);
nand U4600 (N_4600,N_3841,N_305);
nor U4601 (N_4601,N_239,N_2905);
xor U4602 (N_4602,N_3368,N_3454);
xor U4603 (N_4603,N_352,N_3031);
and U4604 (N_4604,N_1267,N_3746);
and U4605 (N_4605,N_2233,N_869);
and U4606 (N_4606,N_3922,N_2915);
or U4607 (N_4607,N_3652,N_1365);
xnor U4608 (N_4608,N_3350,N_1116);
nand U4609 (N_4609,N_400,N_1101);
xor U4610 (N_4610,N_2011,N_3701);
nor U4611 (N_4611,N_3186,N_947);
and U4612 (N_4612,N_432,N_3056);
or U4613 (N_4613,N_3920,N_3215);
nand U4614 (N_4614,N_854,N_2166);
and U4615 (N_4615,N_65,N_3346);
and U4616 (N_4616,N_2937,N_583);
and U4617 (N_4617,N_2029,N_2960);
and U4618 (N_4618,N_2460,N_2020);
or U4619 (N_4619,N_2885,N_826);
xor U4620 (N_4620,N_3334,N_949);
nand U4621 (N_4621,N_1578,N_2008);
xor U4622 (N_4622,N_1038,N_1707);
or U4623 (N_4623,N_1728,N_2161);
xnor U4624 (N_4624,N_2548,N_2580);
xnor U4625 (N_4625,N_3129,N_230);
nor U4626 (N_4626,N_3574,N_1749);
or U4627 (N_4627,N_3003,N_209);
nand U4628 (N_4628,N_3193,N_1575);
or U4629 (N_4629,N_155,N_76);
nor U4630 (N_4630,N_3065,N_615);
nand U4631 (N_4631,N_2617,N_1548);
nor U4632 (N_4632,N_662,N_402);
nand U4633 (N_4633,N_653,N_2176);
nor U4634 (N_4634,N_3537,N_705);
and U4635 (N_4635,N_384,N_1841);
nand U4636 (N_4636,N_1349,N_2177);
xor U4637 (N_4637,N_1447,N_1088);
xnor U4638 (N_4638,N_3848,N_2673);
and U4639 (N_4639,N_1521,N_3684);
and U4640 (N_4640,N_630,N_1225);
nor U4641 (N_4641,N_1023,N_3519);
or U4642 (N_4642,N_3781,N_2112);
xnor U4643 (N_4643,N_915,N_1901);
and U4644 (N_4644,N_1073,N_1110);
nand U4645 (N_4645,N_3878,N_320);
nand U4646 (N_4646,N_930,N_2804);
xnor U4647 (N_4647,N_1608,N_2006);
nand U4648 (N_4648,N_1464,N_2649);
xor U4649 (N_4649,N_1213,N_580);
or U4650 (N_4650,N_2445,N_3711);
nor U4651 (N_4651,N_251,N_248);
xnor U4652 (N_4652,N_3957,N_1307);
nor U4653 (N_4653,N_1891,N_275);
xnor U4654 (N_4654,N_2152,N_3908);
nor U4655 (N_4655,N_3241,N_2243);
xor U4656 (N_4656,N_2868,N_2566);
and U4657 (N_4657,N_196,N_1545);
and U4658 (N_4658,N_3984,N_87);
xnor U4659 (N_4659,N_504,N_138);
xor U4660 (N_4660,N_1348,N_2891);
or U4661 (N_4661,N_1305,N_39);
nand U4662 (N_4662,N_3849,N_2878);
xnor U4663 (N_4663,N_3698,N_3072);
nor U4664 (N_4664,N_3819,N_1572);
nor U4665 (N_4665,N_1774,N_2609);
xor U4666 (N_4666,N_3485,N_1260);
and U4667 (N_4667,N_1239,N_3013);
or U4668 (N_4668,N_3603,N_3182);
or U4669 (N_4669,N_2983,N_3816);
and U4670 (N_4670,N_3500,N_385);
xor U4671 (N_4671,N_1906,N_2831);
or U4672 (N_4672,N_3904,N_2402);
and U4673 (N_4673,N_2072,N_439);
and U4674 (N_4674,N_1909,N_3110);
and U4675 (N_4675,N_2997,N_2826);
nand U4676 (N_4676,N_1960,N_96);
or U4677 (N_4677,N_2846,N_2901);
and U4678 (N_4678,N_3595,N_2752);
xnor U4679 (N_4679,N_2814,N_714);
nand U4680 (N_4680,N_469,N_616);
or U4681 (N_4681,N_3302,N_367);
xnor U4682 (N_4682,N_3886,N_2145);
xor U4683 (N_4683,N_3693,N_217);
nor U4684 (N_4684,N_1670,N_1652);
or U4685 (N_4685,N_945,N_1465);
nand U4686 (N_4686,N_3247,N_2379);
nor U4687 (N_4687,N_3689,N_245);
nand U4688 (N_4688,N_1939,N_1689);
xnor U4689 (N_4689,N_1941,N_3741);
nand U4690 (N_4690,N_2438,N_814);
nand U4691 (N_4691,N_2892,N_3476);
xor U4692 (N_4692,N_2964,N_2249);
xor U4693 (N_4693,N_1876,N_490);
and U4694 (N_4694,N_2075,N_567);
nor U4695 (N_4695,N_647,N_440);
or U4696 (N_4696,N_1565,N_2452);
or U4697 (N_4697,N_2080,N_3465);
and U4698 (N_4698,N_2972,N_1185);
or U4699 (N_4699,N_1357,N_759);
xor U4700 (N_4700,N_121,N_628);
and U4701 (N_4701,N_1808,N_2408);
nor U4702 (N_4702,N_1724,N_110);
and U4703 (N_4703,N_3695,N_234);
or U4704 (N_4704,N_1884,N_2667);
nor U4705 (N_4705,N_1069,N_3093);
or U4706 (N_4706,N_3507,N_3584);
and U4707 (N_4707,N_985,N_2839);
nand U4708 (N_4708,N_3869,N_3606);
nor U4709 (N_4709,N_912,N_2944);
nor U4710 (N_4710,N_2903,N_397);
and U4711 (N_4711,N_1944,N_540);
and U4712 (N_4712,N_2527,N_1526);
or U4713 (N_4713,N_3728,N_3858);
nand U4714 (N_4714,N_1534,N_537);
and U4715 (N_4715,N_1956,N_3408);
nor U4716 (N_4716,N_2919,N_1531);
xor U4717 (N_4717,N_2568,N_972);
nor U4718 (N_4718,N_116,N_2511);
xnor U4719 (N_4719,N_1704,N_2115);
nor U4720 (N_4720,N_1813,N_199);
nor U4721 (N_4721,N_3000,N_1731);
or U4722 (N_4722,N_2884,N_2660);
xnor U4723 (N_4723,N_1164,N_2736);
xnor U4724 (N_4724,N_2534,N_3268);
or U4725 (N_4725,N_1914,N_2263);
or U4726 (N_4726,N_3899,N_1298);
nor U4727 (N_4727,N_2705,N_2734);
and U4728 (N_4728,N_2676,N_2614);
nand U4729 (N_4729,N_1498,N_3573);
or U4730 (N_4730,N_3385,N_2920);
xor U4731 (N_4731,N_2797,N_820);
or U4732 (N_4732,N_497,N_329);
xor U4733 (N_4733,N_1717,N_929);
nor U4734 (N_4734,N_2975,N_2290);
xor U4735 (N_4735,N_2431,N_2012);
or U4736 (N_4736,N_2740,N_853);
or U4737 (N_4737,N_3387,N_3472);
nand U4738 (N_4738,N_3638,N_2532);
or U4739 (N_4739,N_2642,N_3861);
xnor U4740 (N_4740,N_2085,N_2360);
nand U4741 (N_4741,N_614,N_2099);
or U4742 (N_4742,N_802,N_3145);
or U4743 (N_4743,N_3210,N_338);
and U4744 (N_4744,N_1452,N_339);
and U4745 (N_4745,N_2417,N_1292);
or U4746 (N_4746,N_2750,N_346);
nor U4747 (N_4747,N_932,N_2735);
nor U4748 (N_4748,N_1333,N_931);
nand U4749 (N_4749,N_2102,N_1405);
or U4750 (N_4750,N_3002,N_3974);
xnor U4751 (N_4751,N_2456,N_2196);
and U4752 (N_4752,N_2632,N_678);
or U4753 (N_4753,N_302,N_836);
xnor U4754 (N_4754,N_3882,N_1561);
and U4755 (N_4755,N_3915,N_1796);
nand U4756 (N_4756,N_256,N_1);
nor U4757 (N_4757,N_300,N_2372);
xnor U4758 (N_4758,N_3506,N_2475);
nor U4759 (N_4759,N_1541,N_1081);
or U4760 (N_4760,N_1144,N_3332);
and U4761 (N_4761,N_3618,N_3291);
nand U4762 (N_4762,N_37,N_429);
and U4763 (N_4763,N_2261,N_3032);
and U4764 (N_4764,N_3720,N_2017);
xnor U4765 (N_4765,N_1712,N_3687);
nor U4766 (N_4766,N_3280,N_2764);
or U4767 (N_4767,N_3810,N_3176);
nor U4768 (N_4768,N_403,N_1178);
or U4769 (N_4769,N_231,N_2989);
nand U4770 (N_4770,N_3489,N_3425);
and U4771 (N_4771,N_1096,N_3795);
xor U4772 (N_4772,N_3649,N_3085);
xor U4773 (N_4773,N_856,N_1282);
nand U4774 (N_4774,N_193,N_311);
nor U4775 (N_4775,N_210,N_1690);
nor U4776 (N_4776,N_315,N_517);
xnor U4777 (N_4777,N_1276,N_951);
nor U4778 (N_4778,N_1429,N_413);
nand U4779 (N_4779,N_262,N_148);
xor U4780 (N_4780,N_3586,N_1700);
or U4781 (N_4781,N_3492,N_813);
or U4782 (N_4782,N_2276,N_3285);
and U4783 (N_4783,N_3502,N_438);
xnor U4784 (N_4784,N_737,N_1019);
and U4785 (N_4785,N_1393,N_3637);
nand U4786 (N_4786,N_1309,N_427);
xor U4787 (N_4787,N_2840,N_2844);
xnor U4788 (N_4788,N_3850,N_1847);
xor U4789 (N_4789,N_3157,N_3301);
xor U4790 (N_4790,N_1515,N_2236);
xnor U4791 (N_4791,N_3224,N_3490);
nand U4792 (N_4792,N_2646,N_2658);
nor U4793 (N_4793,N_3791,N_2459);
nand U4794 (N_4794,N_3733,N_987);
and U4795 (N_4795,N_619,N_1094);
xnor U4796 (N_4796,N_989,N_1477);
and U4797 (N_4797,N_2564,N_563);
xnor U4798 (N_4798,N_3161,N_638);
nor U4799 (N_4799,N_3916,N_1711);
or U4800 (N_4800,N_1364,N_3964);
and U4801 (N_4801,N_3130,N_1510);
nand U4802 (N_4802,N_288,N_355);
or U4803 (N_4803,N_3078,N_1227);
or U4804 (N_4804,N_1083,N_1346);
and U4805 (N_4805,N_10,N_828);
and U4806 (N_4806,N_908,N_528);
or U4807 (N_4807,N_182,N_2495);
nand U4808 (N_4808,N_794,N_242);
nand U4809 (N_4809,N_3703,N_2310);
or U4810 (N_4810,N_2762,N_1767);
nor U4811 (N_4811,N_380,N_3846);
nand U4812 (N_4812,N_2850,N_3232);
xnor U4813 (N_4813,N_3426,N_2359);
xor U4814 (N_4814,N_2150,N_3494);
or U4815 (N_4815,N_2794,N_154);
or U4816 (N_4816,N_2540,N_1118);
nor U4817 (N_4817,N_1432,N_3757);
nor U4818 (N_4818,N_1486,N_2362);
xnor U4819 (N_4819,N_1222,N_2837);
and U4820 (N_4820,N_610,N_3917);
and U4821 (N_4821,N_1698,N_2686);
nor U4822 (N_4822,N_3782,N_298);
nand U4823 (N_4823,N_3610,N_1667);
nor U4824 (N_4824,N_134,N_3805);
xnor U4825 (N_4825,N_1990,N_3714);
or U4826 (N_4826,N_414,N_3240);
and U4827 (N_4827,N_3590,N_1973);
nor U4828 (N_4828,N_2859,N_2197);
nor U4829 (N_4829,N_1035,N_974);
nand U4830 (N_4830,N_3281,N_437);
and U4831 (N_4831,N_3761,N_3483);
or U4832 (N_4832,N_3905,N_3166);
and U4833 (N_4833,N_645,N_1849);
xnor U4834 (N_4834,N_3699,N_3934);
and U4835 (N_4835,N_3725,N_576);
and U4836 (N_4836,N_1518,N_1801);
nand U4837 (N_4837,N_2823,N_3287);
xor U4838 (N_4838,N_1959,N_249);
nor U4839 (N_4839,N_2785,N_3370);
xnor U4840 (N_4840,N_3991,N_3516);
nor U4841 (N_4841,N_9,N_2863);
and U4842 (N_4842,N_3090,N_100);
xor U4843 (N_4843,N_2560,N_2289);
xnor U4844 (N_4844,N_2961,N_3323);
or U4845 (N_4845,N_1046,N_2613);
xor U4846 (N_4846,N_3286,N_2866);
and U4847 (N_4847,N_2293,N_3009);
nor U4848 (N_4848,N_1845,N_1201);
nor U4849 (N_4849,N_3531,N_601);
or U4850 (N_4850,N_822,N_3933);
nor U4851 (N_4851,N_1969,N_1828);
nor U4852 (N_4852,N_2357,N_582);
xor U4853 (N_4853,N_1867,N_1085);
and U4854 (N_4854,N_2059,N_3569);
and U4855 (N_4855,N_1932,N_1616);
xor U4856 (N_4856,N_3477,N_855);
nor U4857 (N_4857,N_3925,N_229);
nand U4858 (N_4858,N_3842,N_3007);
nor U4859 (N_4859,N_3673,N_3455);
nand U4860 (N_4860,N_1183,N_2712);
and U4861 (N_4861,N_2134,N_1842);
xor U4862 (N_4862,N_3550,N_1422);
nand U4863 (N_4863,N_2052,N_1086);
nor U4864 (N_4864,N_1674,N_1313);
nor U4865 (N_4865,N_741,N_3653);
xor U4866 (N_4866,N_3544,N_2284);
nand U4867 (N_4867,N_3011,N_2449);
nand U4868 (N_4868,N_3487,N_2229);
nand U4869 (N_4869,N_2342,N_1788);
nor U4870 (N_4870,N_3289,N_2423);
and U4871 (N_4871,N_2634,N_500);
or U4872 (N_4872,N_1047,N_3706);
xnor U4873 (N_4873,N_1633,N_327);
xor U4874 (N_4874,N_1150,N_1301);
xnor U4875 (N_4875,N_3983,N_2847);
and U4876 (N_4876,N_1807,N_283);
xor U4877 (N_4877,N_1512,N_3787);
xor U4878 (N_4878,N_3456,N_1718);
nand U4879 (N_4879,N_889,N_883);
nor U4880 (N_4880,N_3417,N_1461);
or U4881 (N_4881,N_2494,N_2465);
and U4882 (N_4882,N_1564,N_3547);
nor U4883 (N_4883,N_1806,N_2329);
and U4884 (N_4884,N_3150,N_3504);
xnor U4885 (N_4885,N_281,N_720);
nand U4886 (N_4886,N_3081,N_3549);
nor U4887 (N_4887,N_3314,N_2469);
xor U4888 (N_4888,N_1269,N_2586);
and U4889 (N_4889,N_259,N_3329);
or U4890 (N_4890,N_2682,N_2350);
or U4891 (N_4891,N_2803,N_2502);
and U4892 (N_4892,N_1589,N_704);
or U4893 (N_4893,N_2116,N_1832);
nor U4894 (N_4894,N_3480,N_2572);
xnor U4895 (N_4895,N_573,N_3035);
xnor U4896 (N_4896,N_550,N_599);
xor U4897 (N_4897,N_1057,N_1547);
xor U4898 (N_4898,N_3192,N_1238);
nor U4899 (N_4899,N_3685,N_2641);
and U4900 (N_4900,N_730,N_3578);
or U4901 (N_4901,N_309,N_2558);
xnor U4902 (N_4902,N_1507,N_620);
xor U4903 (N_4903,N_2678,N_3135);
xnor U4904 (N_4904,N_2708,N_3356);
and U4905 (N_4905,N_3950,N_1179);
xor U4906 (N_4906,N_2044,N_3668);
and U4907 (N_4907,N_865,N_565);
or U4908 (N_4908,N_1273,N_3797);
nand U4909 (N_4909,N_1463,N_1014);
or U4910 (N_4910,N_529,N_1850);
and U4911 (N_4911,N_3885,N_398);
and U4912 (N_4912,N_748,N_805);
xnor U4913 (N_4913,N_593,N_3770);
or U4914 (N_4914,N_2024,N_1091);
and U4915 (N_4915,N_2209,N_3602);
nand U4916 (N_4916,N_1189,N_1462);
and U4917 (N_4917,N_2117,N_3343);
nand U4918 (N_4918,N_3227,N_2958);
nand U4919 (N_4919,N_1645,N_3658);
nor U4920 (N_4920,N_736,N_3405);
and U4921 (N_4921,N_1161,N_2644);
and U4922 (N_4922,N_1641,N_3495);
xnor U4923 (N_4923,N_2555,N_2079);
or U4924 (N_4924,N_1186,N_1055);
nand U4925 (N_4925,N_745,N_332);
xnor U4926 (N_4926,N_2488,N_2204);
or U4927 (N_4927,N_2538,N_3931);
xnor U4928 (N_4928,N_224,N_2761);
or U4929 (N_4929,N_793,N_2087);
xor U4930 (N_4930,N_2337,N_661);
nor U4931 (N_4931,N_1392,N_2038);
or U4932 (N_4932,N_2818,N_2058);
or U4933 (N_4933,N_2720,N_3867);
xnor U4934 (N_4934,N_939,N_52);
xnor U4935 (N_4935,N_1664,N_578);
nor U4936 (N_4936,N_3521,N_2518);
nand U4937 (N_4937,N_1250,N_1131);
xor U4938 (N_4938,N_1146,N_83);
xor U4939 (N_4939,N_1200,N_3245);
and U4940 (N_4940,N_1002,N_2225);
nor U4941 (N_4941,N_3266,N_1555);
or U4942 (N_4942,N_698,N_3624);
nand U4943 (N_4943,N_2820,N_1479);
nor U4944 (N_4944,N_431,N_1311);
xnor U4945 (N_4945,N_1284,N_2281);
xnor U4946 (N_4946,N_2248,N_1603);
xor U4947 (N_4947,N_3070,N_2164);
and U4948 (N_4948,N_588,N_3463);
nor U4949 (N_4949,N_758,N_2807);
or U4950 (N_4950,N_795,N_2094);
nor U4951 (N_4951,N_589,N_2601);
nor U4952 (N_4952,N_3501,N_1468);
nand U4953 (N_4953,N_1583,N_1852);
xor U4954 (N_4954,N_2835,N_1999);
nand U4955 (N_4955,N_3644,N_3949);
nor U4956 (N_4956,N_2579,N_882);
or U4957 (N_4957,N_2013,N_375);
or U4958 (N_4958,N_381,N_762);
nor U4959 (N_4959,N_2303,N_1143);
nand U4960 (N_4960,N_852,N_3069);
or U4961 (N_4961,N_2322,N_709);
nand U4962 (N_4962,N_1398,N_3347);
nand U4963 (N_4963,N_1079,N_3847);
xor U4964 (N_4964,N_2477,N_2822);
or U4965 (N_4965,N_3464,N_1430);
and U4966 (N_4966,N_2898,N_683);
nor U4967 (N_4967,N_372,N_2121);
xnor U4968 (N_4968,N_3939,N_804);
nor U4969 (N_4969,N_3375,N_786);
nand U4970 (N_4970,N_1900,N_3540);
and U4971 (N_4971,N_3140,N_572);
nor U4972 (N_4972,N_3822,N_1170);
or U4973 (N_4973,N_785,N_3515);
and U4974 (N_4974,N_2856,N_1095);
nand U4975 (N_4975,N_522,N_2381);
nand U4976 (N_4976,N_2226,N_257);
nand U4977 (N_4977,N_2409,N_3005);
and U4978 (N_4978,N_3250,N_3024);
nor U4979 (N_4979,N_3989,N_1303);
or U4980 (N_4980,N_396,N_2629);
or U4981 (N_4981,N_484,N_348);
xor U4982 (N_4982,N_106,N_585);
xnor U4983 (N_4983,N_2214,N_3132);
and U4984 (N_4984,N_752,N_161);
nand U4985 (N_4985,N_1401,N_3747);
and U4986 (N_4986,N_2597,N_1132);
nand U4987 (N_4987,N_2246,N_1644);
nor U4988 (N_4988,N_195,N_1586);
nand U4989 (N_4989,N_466,N_612);
nand U4990 (N_4990,N_1658,N_1527);
or U4991 (N_4991,N_1289,N_1623);
or U4992 (N_4992,N_3813,N_3591);
or U4993 (N_4993,N_361,N_3406);
or U4994 (N_4994,N_1831,N_3675);
nand U4995 (N_4995,N_2993,N_3536);
nand U4996 (N_4996,N_3038,N_1377);
and U4997 (N_4997,N_1256,N_2146);
or U4998 (N_4998,N_1244,N_1922);
and U4999 (N_4999,N_943,N_3765);
or U5000 (N_5000,N_1746,N_3801);
and U5001 (N_5001,N_2777,N_1071);
or U5002 (N_5002,N_1236,N_1988);
or U5003 (N_5003,N_353,N_1991);
nor U5004 (N_5004,N_2428,N_860);
nand U5005 (N_5005,N_2033,N_1050);
xor U5006 (N_5006,N_3736,N_1414);
or U5007 (N_5007,N_273,N_2779);
or U5008 (N_5008,N_3555,N_1117);
and U5009 (N_5009,N_136,N_1382);
or U5010 (N_5010,N_3890,N_3587);
and U5011 (N_5011,N_1653,N_1402);
nor U5012 (N_5012,N_391,N_2651);
nor U5013 (N_5013,N_78,N_1676);
nand U5014 (N_5014,N_3626,N_2387);
and U5015 (N_5015,N_1595,N_130);
nor U5016 (N_5016,N_3479,N_2037);
or U5017 (N_5017,N_1336,N_2299);
and U5018 (N_5018,N_2965,N_3196);
and U5019 (N_5019,N_3365,N_3330);
nand U5020 (N_5020,N_3643,N_2748);
nand U5021 (N_5021,N_411,N_3064);
or U5022 (N_5022,N_3738,N_3533);
xor U5023 (N_5023,N_2142,N_3941);
nor U5024 (N_5024,N_3648,N_18);
and U5025 (N_5025,N_3601,N_2900);
and U5026 (N_5026,N_1306,N_2426);
and U5027 (N_5027,N_757,N_755);
nor U5028 (N_5028,N_1017,N_3460);
xor U5029 (N_5029,N_3440,N_2471);
xor U5030 (N_5030,N_2962,N_677);
or U5031 (N_5031,N_3530,N_2285);
nor U5032 (N_5032,N_175,N_2832);
xnor U5033 (N_5033,N_2397,N_2661);
nand U5034 (N_5034,N_825,N_3061);
nand U5035 (N_5035,N_3873,N_1877);
and U5036 (N_5036,N_688,N_2611);
and U5037 (N_5037,N_2988,N_1350);
or U5038 (N_5038,N_3230,N_2833);
nand U5039 (N_5039,N_2089,N_3628);
and U5040 (N_5040,N_416,N_2066);
xor U5041 (N_5041,N_1435,N_1992);
nor U5042 (N_5042,N_834,N_734);
xnor U5043 (N_5043,N_1280,N_2185);
xnor U5044 (N_5044,N_531,N_3491);
or U5045 (N_5045,N_817,N_2787);
xnor U5046 (N_5046,N_3646,N_2340);
and U5047 (N_5047,N_2879,N_228);
nand U5048 (N_5048,N_168,N_3171);
xnor U5049 (N_5049,N_776,N_873);
and U5050 (N_5050,N_3768,N_84);
nor U5051 (N_5051,N_1322,N_841);
nor U5052 (N_5052,N_1076,N_511);
nand U5053 (N_5053,N_3594,N_3420);
or U5054 (N_5054,N_553,N_3074);
nor U5055 (N_5055,N_2179,N_1470);
and U5056 (N_5056,N_2188,N_2512);
and U5057 (N_5057,N_2523,N_1958);
or U5058 (N_5058,N_3802,N_3677);
or U5059 (N_5059,N_2584,N_1190);
or U5060 (N_5060,N_1297,N_2809);
and U5061 (N_5061,N_921,N_750);
or U5062 (N_5062,N_1387,N_1579);
nor U5063 (N_5063,N_2280,N_3807);
or U5064 (N_5064,N_3086,N_2786);
nor U5065 (N_5065,N_3030,N_213);
nand U5066 (N_5066,N_3508,N_1028);
or U5067 (N_5067,N_1312,N_368);
nand U5068 (N_5068,N_1800,N_304);
nand U5069 (N_5069,N_284,N_1904);
nand U5070 (N_5070,N_973,N_568);
nor U5071 (N_5071,N_3702,N_687);
or U5072 (N_5072,N_1404,N_3233);
or U5073 (N_5073,N_3062,N_1484);
nand U5074 (N_5074,N_1582,N_2217);
or U5075 (N_5075,N_2966,N_308);
and U5076 (N_5076,N_2368,N_1626);
and U5077 (N_5077,N_1259,N_1787);
and U5078 (N_5078,N_2447,N_3855);
and U5079 (N_5079,N_2439,N_1457);
nor U5080 (N_5080,N_212,N_3700);
xnor U5081 (N_5081,N_265,N_2306);
and U5082 (N_5082,N_1553,N_2767);
or U5083 (N_5083,N_674,N_1661);
nand U5084 (N_5084,N_1593,N_1338);
nand U5085 (N_5085,N_3605,N_2684);
nor U5086 (N_5086,N_321,N_2491);
and U5087 (N_5087,N_3910,N_2902);
xor U5088 (N_5088,N_408,N_1495);
and U5089 (N_5089,N_541,N_3900);
nor U5090 (N_5090,N_157,N_1433);
or U5091 (N_5091,N_2355,N_1121);
or U5092 (N_5092,N_3527,N_2896);
nor U5093 (N_5093,N_2068,N_3010);
or U5094 (N_5094,N_3023,N_241);
xnor U5095 (N_5095,N_2425,N_3352);
and U5096 (N_5096,N_626,N_285);
nor U5097 (N_5097,N_2954,N_204);
nand U5098 (N_5098,N_1320,N_926);
or U5099 (N_5099,N_2405,N_460);
xor U5100 (N_5100,N_1924,N_98);
or U5101 (N_5101,N_1729,N_2912);
and U5102 (N_5102,N_1196,N_1056);
nor U5103 (N_5103,N_2894,N_23);
nor U5104 (N_5104,N_3044,N_840);
or U5105 (N_5105,N_3520,N_2378);
or U5106 (N_5106,N_2404,N_2986);
nor U5107 (N_5107,N_733,N_3872);
xor U5108 (N_5108,N_897,N_3278);
nor U5109 (N_5109,N_3809,N_2343);
xnor U5110 (N_5110,N_3866,N_2713);
nand U5111 (N_5111,N_3478,N_1805);
nor U5112 (N_5112,N_1337,N_2412);
and U5113 (N_5113,N_1551,N_2698);
xnor U5114 (N_5114,N_3339,N_3988);
xor U5115 (N_5115,N_1997,N_1705);
nand U5116 (N_5116,N_3026,N_962);
nand U5117 (N_5117,N_3433,N_2493);
and U5118 (N_5118,N_279,N_1594);
or U5119 (N_5119,N_2810,N_1785);
xnor U5120 (N_5120,N_3095,N_2042);
nor U5121 (N_5121,N_3597,N_1974);
nor U5122 (N_5122,N_1760,N_340);
and U5123 (N_5123,N_2685,N_1783);
nand U5124 (N_5124,N_1419,N_464);
xor U5125 (N_5125,N_2109,N_1568);
or U5126 (N_5126,N_1157,N_1501);
and U5127 (N_5127,N_1208,N_3058);
nor U5128 (N_5128,N_3942,N_3914);
and U5129 (N_5129,N_310,N_453);
or U5130 (N_5130,N_1684,N_2970);
or U5131 (N_5131,N_3357,N_3321);
nand U5132 (N_5132,N_3615,N_1080);
and U5133 (N_5133,N_1456,N_3993);
and U5134 (N_5134,N_1485,N_3057);
nor U5135 (N_5135,N_2509,N_712);
or U5136 (N_5136,N_358,N_850);
and U5137 (N_5137,N_492,N_2205);
or U5138 (N_5138,N_1860,N_2525);
or U5139 (N_5139,N_1373,N_2689);
xnor U5140 (N_5140,N_2792,N_3683);
xnor U5141 (N_5141,N_425,N_3944);
or U5142 (N_5142,N_2671,N_1268);
xor U5143 (N_5143,N_968,N_679);
nor U5144 (N_5144,N_3566,N_2865);
xnor U5145 (N_5145,N_667,N_3360);
or U5146 (N_5146,N_1007,N_2895);
nor U5147 (N_5147,N_3509,N_659);
nor U5148 (N_5148,N_907,N_1837);
or U5149 (N_5149,N_2211,N_2784);
nand U5150 (N_5150,N_3379,N_3181);
nand U5151 (N_5151,N_1020,N_2654);
xnor U5152 (N_5152,N_3234,N_3097);
and U5153 (N_5153,N_409,N_1946);
nand U5154 (N_5154,N_809,N_1989);
and U5155 (N_5155,N_1931,N_2716);
nor U5156 (N_5156,N_2711,N_1714);
nor U5157 (N_5157,N_2598,N_2928);
or U5158 (N_5158,N_171,N_2421);
nand U5159 (N_5159,N_2991,N_2559);
nand U5160 (N_5160,N_1151,N_2985);
nand U5161 (N_5161,N_3879,N_2553);
or U5162 (N_5162,N_878,N_3310);
or U5163 (N_5163,N_682,N_2253);
nor U5164 (N_5164,N_481,N_3682);
nor U5165 (N_5165,N_2500,N_2655);
xor U5166 (N_5166,N_675,N_1036);
xnor U5167 (N_5167,N_1006,N_1669);
nor U5168 (N_5168,N_1955,N_1982);
xor U5169 (N_5169,N_3992,N_2467);
xnor U5170 (N_5170,N_532,N_1646);
and U5171 (N_5171,N_2824,N_390);
nand U5172 (N_5172,N_1596,N_3830);
or U5173 (N_5173,N_884,N_2772);
and U5174 (N_5174,N_1859,N_1696);
or U5175 (N_5175,N_3632,N_1708);
nor U5176 (N_5176,N_928,N_751);
xor U5177 (N_5177,N_3523,N_3014);
or U5178 (N_5178,N_721,N_47);
nor U5179 (N_5179,N_143,N_2808);
xor U5180 (N_5180,N_3588,N_3923);
xor U5181 (N_5181,N_3349,N_1863);
nor U5182 (N_5182,N_727,N_1115);
nand U5183 (N_5183,N_1271,N_3665);
nor U5184 (N_5184,N_2636,N_2665);
nor U5185 (N_5185,N_2155,N_2770);
and U5186 (N_5186,N_1355,N_2275);
nand U5187 (N_5187,N_70,N_1453);
or U5188 (N_5188,N_723,N_2924);
xor U5189 (N_5189,N_1246,N_1902);
nand U5190 (N_5190,N_2746,N_1043);
and U5191 (N_5191,N_3336,N_1252);
nand U5192 (N_5192,N_2544,N_2893);
and U5193 (N_5193,N_1908,N_1249);
xor U5194 (N_5194,N_535,N_1104);
and U5195 (N_5195,N_149,N_1439);
and U5196 (N_5196,N_333,N_486);
or U5197 (N_5197,N_3386,N_3083);
xnor U5198 (N_5198,N_3812,N_728);
or U5199 (N_5199,N_2739,N_2942);
xor U5200 (N_5200,N_2829,N_1840);
and U5201 (N_5201,N_3851,N_95);
nor U5202 (N_5202,N_964,N_3581);
or U5203 (N_5203,N_632,N_1951);
xnor U5204 (N_5204,N_526,N_2737);
nor U5205 (N_5205,N_3113,N_2571);
or U5206 (N_5206,N_2071,N_1000);
nor U5207 (N_5207,N_3883,N_519);
xor U5208 (N_5208,N_2298,N_198);
nor U5209 (N_5209,N_3651,N_986);
nor U5210 (N_5210,N_3,N_3141);
nor U5211 (N_5211,N_3138,N_1438);
nor U5212 (N_5212,N_1567,N_3676);
xor U5213 (N_5213,N_1105,N_2053);
nor U5214 (N_5214,N_448,N_1651);
or U5215 (N_5215,N_598,N_3190);
nand U5216 (N_5216,N_515,N_3998);
and U5217 (N_5217,N_520,N_51);
or U5218 (N_5218,N_1957,N_3554);
and U5219 (N_5219,N_821,N_633);
xnor U5220 (N_5220,N_2266,N_3340);
or U5221 (N_5221,N_2170,N_838);
or U5222 (N_5222,N_876,N_546);
xnor U5223 (N_5223,N_3189,N_3947);
nand U5224 (N_5224,N_1732,N_979);
nor U5225 (N_5225,N_1330,N_1381);
nor U5226 (N_5226,N_2100,N_158);
nor U5227 (N_5227,N_2349,N_2095);
nor U5228 (N_5228,N_2105,N_657);
nand U5229 (N_5229,N_689,N_3183);
and U5230 (N_5230,N_1720,N_2638);
nor U5231 (N_5231,N_1093,N_2172);
and U5232 (N_5232,N_2065,N_1275);
nand U5233 (N_5233,N_999,N_3880);
xnor U5234 (N_5234,N_2876,N_3681);
and U5235 (N_5235,N_3264,N_2309);
nand U5236 (N_5236,N_3344,N_1942);
xnor U5237 (N_5237,N_981,N_2313);
xor U5238 (N_5238,N_3640,N_2304);
and U5239 (N_5239,N_1370,N_2320);
or U5240 (N_5240,N_1638,N_1215);
nand U5241 (N_5241,N_935,N_2791);
nor U5242 (N_5242,N_717,N_2930);
nand U5243 (N_5243,N_1380,N_3532);
nor U5244 (N_5244,N_1410,N_3045);
xnor U5245 (N_5245,N_3474,N_772);
or U5246 (N_5246,N_3080,N_435);
xor U5247 (N_5247,N_2754,N_2463);
or U5248 (N_5248,N_937,N_954);
nand U5249 (N_5249,N_1128,N_2470);
or U5250 (N_5250,N_2519,N_1358);
xor U5251 (N_5251,N_3203,N_2706);
nand U5252 (N_5252,N_3717,N_2254);
or U5253 (N_5253,N_796,N_2952);
nand U5254 (N_5254,N_377,N_3548);
nor U5255 (N_5255,N_1919,N_2747);
xnor U5256 (N_5256,N_181,N_2815);
nor U5257 (N_5257,N_2717,N_2139);
nand U5258 (N_5258,N_1125,N_2546);
nor U5259 (N_5259,N_452,N_1519);
nand U5260 (N_5260,N_3525,N_959);
or U5261 (N_5261,N_2278,N_2935);
nand U5262 (N_5262,N_1581,N_3006);
nand U5263 (N_5263,N_554,N_1403);
and U5264 (N_5264,N_34,N_192);
nand U5265 (N_5265,N_3043,N_3709);
and U5266 (N_5266,N_2481,N_1986);
or U5267 (N_5267,N_1102,N_607);
and U5268 (N_5268,N_2124,N_114);
xor U5269 (N_5269,N_1025,N_1754);
or U5270 (N_5270,N_2474,N_3067);
or U5271 (N_5271,N_1743,N_1780);
and U5272 (N_5272,N_3423,N_503);
nand U5273 (N_5273,N_71,N_3558);
nor U5274 (N_5274,N_792,N_197);
xnor U5275 (N_5275,N_3019,N_445);
nand U5276 (N_5276,N_2492,N_788);
and U5277 (N_5277,N_1636,N_1127);
and U5278 (N_5278,N_2,N_1895);
or U5279 (N_5279,N_754,N_815);
and U5280 (N_5280,N_1968,N_1976);
xnor U5281 (N_5281,N_31,N_746);
nor U5282 (N_5282,N_2270,N_1097);
and U5283 (N_5283,N_1878,N_2140);
xor U5284 (N_5284,N_2990,N_2973);
xor U5285 (N_5285,N_3424,N_3398);
and U5286 (N_5286,N_560,N_3279);
or U5287 (N_5287,N_1420,N_2245);
xor U5288 (N_5288,N_983,N_837);
nor U5289 (N_5289,N_2688,N_2929);
xor U5290 (N_5290,N_1202,N_2247);
nand U5291 (N_5291,N_2778,N_301);
xnor U5292 (N_5292,N_2974,N_1763);
nor U5293 (N_5293,N_2370,N_2487);
nand U5294 (N_5294,N_507,N_2262);
and U5295 (N_5295,N_2581,N_1334);
xnor U5296 (N_5296,N_2595,N_3382);
and U5297 (N_5297,N_1740,N_501);
xor U5298 (N_5298,N_1417,N_1072);
or U5299 (N_5299,N_621,N_1087);
xnor U5300 (N_5300,N_3337,N_1467);
or U5301 (N_5301,N_19,N_3952);
nand U5302 (N_5302,N_904,N_2653);
and U5303 (N_5303,N_3127,N_139);
and U5304 (N_5304,N_2004,N_1680);
nor U5305 (N_5305,N_3666,N_890);
nand U5306 (N_5306,N_3445,N_1443);
nor U5307 (N_5307,N_2939,N_1281);
nor U5308 (N_5308,N_2224,N_564);
or U5309 (N_5309,N_141,N_2858);
nor U5310 (N_5310,N_123,N_895);
or U5311 (N_5311,N_3710,N_2466);
nand U5312 (N_5312,N_2798,N_900);
nor U5313 (N_5313,N_1248,N_896);
xnor U5314 (N_5314,N_3979,N_2398);
or U5315 (N_5315,N_2628,N_2341);
nor U5316 (N_5316,N_2524,N_1012);
xor U5317 (N_5317,N_3897,N_3244);
nand U5318 (N_5318,N_1491,N_2691);
and U5319 (N_5319,N_533,N_359);
nor U5320 (N_5320,N_3137,N_2650);
nand U5321 (N_5321,N_1761,N_344);
or U5322 (N_5322,N_3180,N_2323);
and U5323 (N_5323,N_151,N_1068);
or U5324 (N_5324,N_2154,N_3363);
xnor U5325 (N_5325,N_1826,N_769);
nor U5326 (N_5326,N_3265,N_629);
nand U5327 (N_5327,N_780,N_459);
or U5328 (N_5328,N_3935,N_3488);
and U5329 (N_5329,N_652,N_3926);
or U5330 (N_5330,N_2639,N_1061);
or U5331 (N_5331,N_2619,N_885);
xor U5332 (N_5332,N_2432,N_715);
and U5333 (N_5333,N_1302,N_2561);
nor U5334 (N_5334,N_2143,N_2325);
xor U5335 (N_5335,N_3207,N_1231);
nor U5336 (N_5336,N_991,N_3252);
xor U5337 (N_5337,N_1011,N_1779);
xor U5338 (N_5338,N_1784,N_1866);
nand U5339 (N_5339,N_3439,N_190);
xor U5340 (N_5340,N_3260,N_2608);
and U5341 (N_5341,N_597,N_3786);
or U5342 (N_5342,N_3860,N_312);
and U5343 (N_5343,N_1082,N_3696);
or U5344 (N_5344,N_1171,N_648);
xnor U5345 (N_5345,N_3272,N_255);
or U5346 (N_5346,N_1843,N_2916);
nor U5347 (N_5347,N_975,N_2328);
and U5348 (N_5348,N_108,N_3707);
xnor U5349 (N_5349,N_3745,N_2562);
or U5350 (N_5350,N_2625,N_2718);
xnor U5351 (N_5351,N_646,N_1635);
and U5352 (N_5352,N_1765,N_1015);
or U5353 (N_5353,N_2605,N_3107);
xor U5354 (N_5354,N_2593,N_274);
xor U5355 (N_5355,N_2710,N_3894);
nor U5356 (N_5356,N_1790,N_3844);
nor U5357 (N_5357,N_3657,N_2758);
and U5358 (N_5358,N_697,N_8);
nand U5359 (N_5359,N_1054,N_3037);
xor U5360 (N_5360,N_2022,N_1153);
nor U5361 (N_5361,N_1977,N_289);
nor U5362 (N_5362,N_2120,N_2358);
nor U5363 (N_5363,N_3018,N_1868);
or U5364 (N_5364,N_2817,N_1678);
and U5365 (N_5365,N_2703,N_3856);
or U5366 (N_5366,N_2241,N_2316);
nand U5367 (N_5367,N_848,N_1817);
nor U5368 (N_5368,N_189,N_830);
nand U5369 (N_5369,N_2707,N_2173);
and U5370 (N_5370,N_863,N_2443);
nand U5371 (N_5371,N_1109,N_1727);
xnor U5372 (N_5372,N_54,N_1324);
nor U5373 (N_5373,N_2418,N_2664);
or U5374 (N_5374,N_3364,N_3066);
and U5375 (N_5375,N_2927,N_2000);
or U5376 (N_5376,N_2925,N_1472);
nand U5377 (N_5377,N_2137,N_3827);
nand U5378 (N_5378,N_2692,N_1395);
or U5379 (N_5379,N_3990,N_3731);
xor U5380 (N_5380,N_2681,N_455);
or U5381 (N_5381,N_3106,N_2514);
nor U5382 (N_5382,N_918,N_3634);
or U5383 (N_5383,N_3854,N_3089);
nor U5384 (N_5384,N_2002,N_3102);
xnor U5385 (N_5385,N_1053,N_2111);
xnor U5386 (N_5386,N_2283,N_3888);
xnor U5387 (N_5387,N_1710,N_1590);
and U5388 (N_5388,N_3659,N_3443);
xor U5389 (N_5389,N_1606,N_891);
and U5390 (N_5390,N_2222,N_2624);
or U5391 (N_5391,N_1184,N_88);
xnor U5392 (N_5392,N_731,N_164);
nor U5393 (N_5393,N_1113,N_1198);
nand U5394 (N_5394,N_3389,N_2719);
and U5395 (N_5395,N_3958,N_3620);
and U5396 (N_5396,N_2828,N_548);
xor U5397 (N_5397,N_2016,N_2932);
nand U5398 (N_5398,N_1063,N_544);
nand U5399 (N_5399,N_1571,N_3052);
and U5400 (N_5400,N_145,N_701);
and U5401 (N_5401,N_654,N_2338);
or U5402 (N_5402,N_3222,N_1733);
or U5403 (N_5403,N_1673,N_282);
nand U5404 (N_5404,N_2971,N_536);
xnor U5405 (N_5405,N_716,N_3362);
and U5406 (N_5406,N_1245,N_72);
or U5407 (N_5407,N_545,N_2136);
and U5408 (N_5408,N_710,N_2906);
nor U5409 (N_5409,N_3104,N_2181);
or U5410 (N_5410,N_1772,N_2420);
nor U5411 (N_5411,N_1159,N_993);
and U5412 (N_5412,N_1953,N_2162);
xor U5413 (N_5413,N_386,N_2615);
nor U5414 (N_5414,N_1615,N_3818);
or U5415 (N_5415,N_3096,N_2616);
xor U5416 (N_5416,N_3889,N_2314);
and U5417 (N_5417,N_1078,N_650);
nand U5418 (N_5418,N_1820,N_2183);
xnor U5419 (N_5419,N_1910,N_451);
and U5420 (N_5420,N_3560,N_2575);
and U5421 (N_5421,N_1873,N_3972);
or U5422 (N_5422,N_1795,N_1889);
or U5423 (N_5423,N_3744,N_3630);
and U5424 (N_5424,N_3261,N_92);
nand U5425 (N_5425,N_1872,N_476);
nor U5426 (N_5426,N_3583,N_2407);
or U5427 (N_5427,N_516,N_3907);
xor U5428 (N_5428,N_104,N_3282);
and U5429 (N_5429,N_2199,N_1459);
nor U5430 (N_5430,N_1257,N_948);
or U5431 (N_5431,N_3664,N_2582);
and U5432 (N_5432,N_3621,N_2943);
and U5433 (N_5433,N_1316,N_2599);
or U5434 (N_5434,N_2255,N_3401);
or U5435 (N_5435,N_3162,N_693);
or U5436 (N_5436,N_206,N_1632);
nor U5437 (N_5437,N_604,N_1092);
or U5438 (N_5438,N_1010,N_602);
xnor U5439 (N_5439,N_3929,N_3943);
and U5440 (N_5440,N_1351,N_3354);
nand U5441 (N_5441,N_1051,N_2630);
xor U5442 (N_5442,N_2269,N_665);
and U5443 (N_5443,N_3996,N_1722);
nand U5444 (N_5444,N_998,N_3295);
nor U5445 (N_5445,N_3924,N_1793);
or U5446 (N_5446,N_2499,N_551);
xor U5447 (N_5447,N_3529,N_3380);
or U5448 (N_5448,N_1587,N_2356);
xnor U5449 (N_5449,N_99,N_1163);
nand U5450 (N_5450,N_159,N_207);
or U5451 (N_5451,N_24,N_3223);
nand U5452 (N_5452,N_2321,N_1296);
nand U5453 (N_5453,N_925,N_68);
or U5454 (N_5454,N_1418,N_2941);
or U5455 (N_5455,N_3109,N_1620);
and U5456 (N_5456,N_2212,N_1778);
nand U5457 (N_5457,N_2369,N_2464);
or U5458 (N_5458,N_1052,N_668);
or U5459 (N_5459,N_3981,N_25);
and U5460 (N_5460,N_3722,N_118);
or U5461 (N_5461,N_3457,N_3893);
nor U5462 (N_5462,N_2125,N_421);
or U5463 (N_5463,N_2333,N_3852);
nand U5464 (N_5464,N_1539,N_1424);
and U5465 (N_5465,N_2504,N_3826);
xor U5466 (N_5466,N_1563,N_3084);
and U5467 (N_5467,N_343,N_1049);
and U5468 (N_5468,N_1898,N_2203);
or U5469 (N_5469,N_3119,N_622);
and U5470 (N_5470,N_590,N_3642);
xor U5471 (N_5471,N_1450,N_2151);
xnor U5472 (N_5472,N_982,N_2086);
or U5473 (N_5473,N_3760,N_800);
nand U5474 (N_5474,N_2497,N_3034);
xor U5475 (N_5475,N_2521,N_2135);
nand U5476 (N_5476,N_1816,N_1855);
or U5477 (N_5477,N_1172,N_1205);
nor U5478 (N_5478,N_2683,N_324);
and U5479 (N_5479,N_976,N_278);
or U5480 (N_5480,N_3748,N_2345);
or U5481 (N_5481,N_357,N_1294);
or U5482 (N_5482,N_1004,N_1916);
nor U5483 (N_5483,N_3088,N_566);
nand U5484 (N_5484,N_2175,N_3936);
nor U5485 (N_5485,N_1726,N_847);
or U5486 (N_5486,N_2551,N_3039);
or U5487 (N_5487,N_3328,N_226);
nand U5488 (N_5488,N_605,N_323);
and U5489 (N_5489,N_3694,N_1971);
nor U5490 (N_5490,N_1685,N_3271);
or U5491 (N_5491,N_1804,N_1331);
and U5492 (N_5492,N_1812,N_917);
or U5493 (N_5493,N_3514,N_1040);
nor U5494 (N_5494,N_508,N_1556);
xnor U5495 (N_5495,N_1899,N_1600);
nand U5496 (N_5496,N_2780,N_2996);
nand U5497 (N_5497,N_3414,N_3619);
nand U5498 (N_5498,N_3258,N_3783);
xor U5499 (N_5499,N_227,N_1640);
nand U5500 (N_5500,N_3049,N_44);
xnor U5501 (N_5501,N_3995,N_906);
nand U5502 (N_5502,N_2662,N_3829);
xor U5503 (N_5503,N_2897,N_1359);
nor U5504 (N_5504,N_2652,N_2354);
nand U5505 (N_5505,N_3542,N_1504);
xor U5506 (N_5506,N_1233,N_465);
xnor U5507 (N_5507,N_2979,N_3004);
nand U5508 (N_5508,N_2618,N_3599);
xor U5509 (N_5509,N_3730,N_1362);
xor U5510 (N_5510,N_3048,N_967);
nor U5511 (N_5511,N_1880,N_3534);
xnor U5512 (N_5512,N_1119,N_1964);
xnor U5513 (N_5513,N_3825,N_2647);
or U5514 (N_5514,N_766,N_2128);
nand U5515 (N_5515,N_1686,N_1224);
and U5516 (N_5516,N_2312,N_3200);
nor U5517 (N_5517,N_2391,N_2265);
nor U5518 (N_5518,N_2510,N_831);
and U5519 (N_5519,N_2202,N_1591);
xor U5520 (N_5520,N_38,N_264);
nor U5521 (N_5521,N_2517,N_1042);
nand U5522 (N_5522,N_2063,N_3142);
nor U5523 (N_5523,N_3149,N_317);
nand U5524 (N_5524,N_2096,N_35);
or U5525 (N_5525,N_2554,N_1605);
xor U5526 (N_5526,N_1945,N_1550);
nand U5527 (N_5527,N_1416,N_2073);
xnor U5528 (N_5528,N_3199,N_2505);
nand U5529 (N_5529,N_1229,N_1181);
xor U5530 (N_5530,N_1122,N_3297);
and U5531 (N_5531,N_1979,N_984);
nor U5532 (N_5532,N_2790,N_2904);
nand U5533 (N_5533,N_1520,N_232);
xnor U5534 (N_5534,N_58,N_2015);
xnor U5535 (N_5535,N_505,N_131);
nand U5536 (N_5536,N_2827,N_394);
and U5537 (N_5537,N_292,N_2549);
and U5538 (N_5538,N_649,N_3243);
nand U5539 (N_5539,N_2687,N_3906);
nor U5540 (N_5540,N_237,N_3754);
nand U5541 (N_5541,N_3645,N_1844);
nand U5542 (N_5542,N_719,N_2300);
nor U5543 (N_5543,N_2191,N_1005);
xnor U5544 (N_5544,N_1602,N_3999);
and U5545 (N_5545,N_827,N_2244);
and U5546 (N_5546,N_1896,N_489);
nor U5547 (N_5547,N_2287,N_1192);
xnor U5548 (N_5548,N_383,N_3639);
or U5549 (N_5549,N_2980,N_3496);
nor U5550 (N_5550,N_3381,N_124);
or U5551 (N_5551,N_3467,N_1621);
nand U5552 (N_5552,N_1234,N_449);
nand U5553 (N_5553,N_1341,N_2395);
nand U5554 (N_5554,N_2987,N_2674);
nand U5555 (N_5555,N_1228,N_1372);
and U5556 (N_5556,N_3122,N_2577);
nor U5557 (N_5557,N_3395,N_880);
and U5558 (N_5558,N_2297,N_2317);
or U5559 (N_5559,N_240,N_180);
nor U5560 (N_5560,N_2373,N_2776);
or U5561 (N_5561,N_2250,N_3585);
xnor U5562 (N_5562,N_3721,N_2709);
xnor U5563 (N_5563,N_2330,N_3814);
and U5564 (N_5564,N_2131,N_1255);
or U5565 (N_5565,N_600,N_3481);
and U5566 (N_5566,N_874,N_183);
and U5567 (N_5567,N_2871,N_3691);
and U5568 (N_5568,N_3853,N_458);
or U5569 (N_5569,N_2437,N_46);
nand U5570 (N_5570,N_2955,N_1409);
or U5571 (N_5571,N_3773,N_2602);
xnor U5572 (N_5572,N_3299,N_980);
and U5573 (N_5573,N_3604,N_2367);
or U5574 (N_5574,N_3087,N_3740);
xnor U5575 (N_5575,N_570,N_1361);
and U5576 (N_5576,N_2025,N_934);
xnor U5577 (N_5577,N_2132,N_2374);
nor U5578 (N_5578,N_1219,N_1815);
nor U5579 (N_5579,N_3769,N_832);
xor U5580 (N_5580,N_2998,N_1274);
or U5581 (N_5581,N_811,N_3742);
nor U5582 (N_5582,N_1961,N_3967);
nand U5583 (N_5583,N_3311,N_3945);
or U5584 (N_5584,N_577,N_2506);
nor U5585 (N_5585,N_2600,N_3403);
and U5586 (N_5586,N_2133,N_801);
nand U5587 (N_5587,N_1371,N_211);
nand U5588 (N_5588,N_892,N_1883);
or U5589 (N_5589,N_81,N_2947);
nand U5590 (N_5590,N_561,N_2783);
and U5591 (N_5591,N_509,N_290);
xnor U5592 (N_5592,N_3975,N_816);
or U5593 (N_5593,N_778,N_1725);
and U5594 (N_5594,N_1074,N_3435);
nor U5595 (N_5595,N_1142,N_618);
nand U5596 (N_5596,N_426,N_3139);
nand U5597 (N_5597,N_2083,N_936);
xnor U5598 (N_5598,N_3378,N_971);
or U5599 (N_5599,N_3169,N_810);
and U5600 (N_5600,N_27,N_806);
or U5601 (N_5601,N_1471,N_1210);
and U5602 (N_5602,N_89,N_2714);
or U5603 (N_5603,N_205,N_3238);
or U5604 (N_5604,N_93,N_3734);
nand U5605 (N_5605,N_2192,N_2383);
nand U5606 (N_5606,N_107,N_2849);
or U5607 (N_5607,N_1524,N_2149);
and U5608 (N_5608,N_753,N_2570);
xnor U5609 (N_5609,N_2036,N_1475);
nor U5610 (N_5610,N_3342,N_3475);
nor U5611 (N_5611,N_2726,N_1716);
and U5612 (N_5612,N_3930,N_2021);
or U5613 (N_5613,N_634,N_627);
xnor U5614 (N_5614,N_3901,N_73);
nor U5615 (N_5615,N_2627,N_1978);
xor U5616 (N_5616,N_1789,N_1532);
xnor U5617 (N_5617,N_3248,N_1762);
nor U5618 (N_5618,N_3674,N_1523);
xor U5619 (N_5619,N_2324,N_581);
xor U5620 (N_5620,N_1321,N_3575);
nor U5621 (N_5621,N_521,N_2104);
and U5622 (N_5622,N_103,N_1715);
nand U5623 (N_5623,N_658,N_2843);
nand U5624 (N_5624,N_3359,N_1223);
xor U5625 (N_5625,N_457,N_1496);
xor U5626 (N_5626,N_3951,N_594);
or U5627 (N_5627,N_1242,N_3876);
nand U5628 (N_5628,N_463,N_3712);
and U5629 (N_5629,N_1926,N_1024);
or U5630 (N_5630,N_97,N_2515);
and U5631 (N_5631,N_2315,N_1771);
and U5632 (N_5632,N_3254,N_202);
nor U5633 (N_5633,N_3891,N_2589);
nand U5634 (N_5634,N_2834,N_1822);
xnor U5635 (N_5635,N_447,N_3938);
and U5636 (N_5636,N_3622,N_2731);
nor U5637 (N_5637,N_2138,N_176);
xor U5638 (N_5638,N_2231,N_2945);
nor U5639 (N_5639,N_718,N_2186);
nor U5640 (N_5640,N_1611,N_3118);
and U5641 (N_5641,N_3593,N_5);
nor U5642 (N_5642,N_2704,N_1907);
nor U5643 (N_5643,N_3237,N_129);
and U5644 (N_5644,N_475,N_2331);
and U5645 (N_5645,N_1654,N_2622);
nand U5646 (N_5646,N_487,N_1665);
or U5647 (N_5647,N_3775,N_1206);
and U5648 (N_5648,N_3269,N_3296);
nand U5649 (N_5649,N_347,N_789);
nor U5650 (N_5650,N_3505,N_1911);
xnor U5651 (N_5651,N_3111,N_270);
nand U5652 (N_5652,N_160,N_2160);
nor U5653 (N_5653,N_443,N_59);
nor U5654 (N_5654,N_3194,N_562);
nand U5655 (N_5655,N_3680,N_140);
and U5656 (N_5656,N_2050,N_2852);
xnor U5657 (N_5657,N_2444,N_1928);
nor U5658 (N_5658,N_2539,N_3451);
nand U5659 (N_5659,N_405,N_3799);
and U5660 (N_5660,N_1655,N_2690);
xnor U5661 (N_5661,N_399,N_2793);
nor U5662 (N_5662,N_3568,N_1530);
xnor U5663 (N_5663,N_3209,N_700);
nor U5664 (N_5664,N_1912,N_2156);
or U5665 (N_5665,N_2663,N_2141);
nor U5666 (N_5666,N_2031,N_109);
and U5667 (N_5667,N_1695,N_3875);
nand U5668 (N_5668,N_2103,N_3218);
nand U5669 (N_5669,N_1679,N_868);
or U5670 (N_5670,N_2334,N_3669);
or U5671 (N_5671,N_1809,N_596);
xnor U5672 (N_5672,N_1343,N_404);
and U5673 (N_5673,N_2567,N_549);
and U5674 (N_5674,N_3178,N_706);
xnor U5675 (N_5675,N_373,N_3510);
or U5676 (N_5676,N_1797,N_152);
and U5677 (N_5677,N_571,N_2657);
xor U5678 (N_5678,N_2292,N_387);
xor U5679 (N_5679,N_2018,N_3055);
nand U5680 (N_5680,N_2110,N_2271);
nand U5681 (N_5681,N_253,N_473);
xor U5682 (N_5682,N_3962,N_2180);
nor U5683 (N_5683,N_86,N_418);
xor U5684 (N_5684,N_60,N_2956);
or U5685 (N_5685,N_3341,N_120);
xnor U5686 (N_5686,N_2168,N_2606);
nand U5687 (N_5687,N_1975,N_1367);
and U5688 (N_5688,N_2635,N_2291);
nor U5689 (N_5689,N_94,N_2861);
or U5690 (N_5690,N_1340,N_2946);
nand U5691 (N_5691,N_2389,N_2393);
or U5692 (N_5692,N_444,N_1984);
nor U5693 (N_5693,N_178,N_1287);
nand U5694 (N_5694,N_3963,N_366);
nand U5695 (N_5695,N_1016,N_3206);
or U5696 (N_5696,N_3912,N_3927);
nand U5697 (N_5697,N_1864,N_3461);
xor U5698 (N_5698,N_3128,N_2056);
and U5699 (N_5699,N_3968,N_3415);
and U5700 (N_5700,N_877,N_2484);
nand U5701 (N_5701,N_1557,N_3966);
nor U5702 (N_5702,N_1300,N_2301);
nor U5703 (N_5703,N_119,N_818);
xnor U5704 (N_5704,N_2165,N_2130);
nor U5705 (N_5705,N_1451,N_483);
and U5706 (N_5706,N_3965,N_924);
or U5707 (N_5707,N_319,N_337);
nand U5708 (N_5708,N_3556,N_2380);
and U5709 (N_5709,N_269,N_2213);
and U5710 (N_5710,N_3932,N_651);
nand U5711 (N_5711,N_1846,N_584);
or U5712 (N_5712,N_3641,N_3185);
or U5713 (N_5713,N_3777,N_3438);
nand U5714 (N_5714,N_835,N_277);
nor U5715 (N_5715,N_1325,N_3650);
or U5716 (N_5716,N_2724,N_782);
nand U5717 (N_5717,N_2026,N_3369);
or U5718 (N_5718,N_3225,N_2067);
or U5719 (N_5719,N_1637,N_960);
nor U5720 (N_5720,N_3441,N_1915);
and U5721 (N_5721,N_3338,N_846);
nor U5722 (N_5722,N_824,N_1573);
or U5723 (N_5723,N_3572,N_173);
nand U5724 (N_5724,N_2223,N_2938);
nor U5725 (N_5725,N_45,N_3446);
or U5726 (N_5726,N_3121,N_3168);
nor U5727 (N_5727,N_2533,N_296);
xor U5728 (N_5728,N_1058,N_2743);
nor U5729 (N_5729,N_3204,N_1559);
nand U5730 (N_5730,N_2799,N_970);
and U5731 (N_5731,N_2468,N_2480);
nand U5732 (N_5732,N_791,N_3997);
xnor U5733 (N_5733,N_1923,N_3607);
nand U5734 (N_5734,N_1277,N_1599);
xnor U5735 (N_5735,N_1839,N_2450);
nand U5736 (N_5736,N_2910,N_1757);
nand U5737 (N_5737,N_2144,N_1345);
or U5738 (N_5738,N_3970,N_2594);
or U5739 (N_5739,N_1481,N_603);
nor U5740 (N_5740,N_2106,N_3792);
nor U5741 (N_5741,N_547,N_3831);
and U5742 (N_5742,N_1751,N_389);
and U5743 (N_5743,N_2294,N_2277);
or U5744 (N_5744,N_3075,N_2621);
xor U5745 (N_5745,N_3688,N_454);
xor U5746 (N_5746,N_2382,N_1400);
xnor U5747 (N_5747,N_1493,N_2169);
or U5748 (N_5748,N_3937,N_997);
or U5749 (N_5749,N_16,N_2949);
and U5750 (N_5750,N_1996,N_1099);
or U5751 (N_5751,N_1737,N_186);
xor U5752 (N_5752,N_1366,N_1962);
nor U5753 (N_5753,N_2696,N_2054);
xnor U5754 (N_5754,N_263,N_2802);
xor U5755 (N_5755,N_946,N_1702);
or U5756 (N_5756,N_2841,N_15);
xnor U5757 (N_5757,N_3837,N_495);
and U5758 (N_5758,N_3001,N_768);
and U5759 (N_5759,N_3798,N_1543);
nand U5760 (N_5760,N_215,N_1323);
and U5761 (N_5761,N_3647,N_1254);
nand U5762 (N_5762,N_42,N_3256);
or U5763 (N_5763,N_2396,N_1965);
xnor U5764 (N_5764,N_2078,N_513);
and U5765 (N_5765,N_901,N_3759);
nand U5766 (N_5766,N_3582,N_3955);
xor U5767 (N_5767,N_2887,N_1770);
xor U5768 (N_5768,N_3811,N_2813);
and U5769 (N_5769,N_3863,N_2242);
and U5770 (N_5770,N_3170,N_2742);
or U5771 (N_5771,N_488,N_3444);
nand U5772 (N_5772,N_2862,N_2123);
or U5773 (N_5773,N_3954,N_2729);
nor U5774 (N_5774,N_3726,N_2501);
and U5775 (N_5775,N_643,N_3973);
or U5776 (N_5776,N_3739,N_1203);
nor U5777 (N_5777,N_1917,N_1810);
xor U5778 (N_5778,N_2221,N_1391);
nor U5779 (N_5779,N_1106,N_7);
nor U5780 (N_5780,N_268,N_1818);
xnor U5781 (N_5781,N_872,N_53);
or U5782 (N_5782,N_2101,N_3470);
nor U5783 (N_5783,N_3763,N_1949);
nor U5784 (N_5784,N_1174,N_1970);
nand U5785 (N_5785,N_2153,N_3091);
or U5786 (N_5786,N_1739,N_1509);
nand U5787 (N_5787,N_2410,N_2607);
or U5788 (N_5788,N_1272,N_2344);
or U5789 (N_5789,N_2603,N_3672);
nor U5790 (N_5790,N_2476,N_1290);
nor U5791 (N_5791,N_1538,N_3845);
and U5792 (N_5792,N_624,N_1149);
xor U5793 (N_5793,N_1848,N_2388);
nand U5794 (N_5794,N_1857,N_172);
and U5795 (N_5795,N_1624,N_30);
and U5796 (N_5796,N_3432,N_992);
xnor U5797 (N_5797,N_2457,N_3046);
xor U5798 (N_5798,N_2854,N_3762);
nor U5799 (N_5799,N_2968,N_3790);
xor U5800 (N_5800,N_2763,N_2039);
and U5801 (N_5801,N_1352,N_345);
or U5802 (N_5802,N_3749,N_3697);
or U5803 (N_5803,N_236,N_3251);
or U5804 (N_5804,N_770,N_225);
and U5805 (N_5805,N_3391,N_3567);
xnor U5806 (N_5806,N_676,N_702);
or U5807 (N_5807,N_1217,N_3896);
nor U5808 (N_5808,N_286,N_1129);
and U5809 (N_5809,N_3325,N_162);
and U5810 (N_5810,N_2694,N_1858);
xor U5811 (N_5811,N_3767,N_2190);
or U5812 (N_5812,N_3373,N_1871);
xnor U5813 (N_5813,N_2715,N_2921);
or U5814 (N_5814,N_170,N_1480);
nand U5815 (N_5815,N_470,N_2529);
nor U5816 (N_5816,N_938,N_3101);
nand U5817 (N_5817,N_1529,N_2032);
nor U5818 (N_5818,N_875,N_1747);
nor U5819 (N_5819,N_2041,N_3319);
xor U5820 (N_5820,N_2352,N_3815);
and U5821 (N_5821,N_2999,N_556);
nand U5822 (N_5822,N_369,N_478);
xor U5823 (N_5823,N_642,N_1943);
or U5824 (N_5824,N_2604,N_844);
xor U5825 (N_5825,N_1168,N_3071);
nor U5826 (N_5826,N_1881,N_3946);
xnor U5827 (N_5827,N_441,N_318);
nor U5828 (N_5828,N_1536,N_1137);
or U5829 (N_5829,N_3315,N_670);
and U5830 (N_5830,N_3322,N_2127);
and U5831 (N_5831,N_260,N_2702);
and U5832 (N_5832,N_608,N_1141);
and U5833 (N_5833,N_1240,N_2371);
or U5834 (N_5834,N_1064,N_3290);
or U5835 (N_5835,N_1317,N_1237);
and U5836 (N_5836,N_807,N_1619);
nand U5837 (N_5837,N_3466,N_3661);
nor U5838 (N_5838,N_3959,N_3042);
nand U5839 (N_5839,N_2220,N_3806);
or U5840 (N_5840,N_3277,N_2883);
or U5841 (N_5841,N_1207,N_2043);
and U5842 (N_5842,N_3497,N_3076);
xor U5843 (N_5843,N_942,N_1823);
xor U5844 (N_5844,N_479,N_2699);
or U5845 (N_5845,N_1397,N_2490);
nor U5846 (N_5846,N_3117,N_2864);
xnor U5847 (N_5847,N_1033,N_1021);
nand U5848 (N_5848,N_2908,N_3633);
xnor U5849 (N_5849,N_3025,N_866);
or U5850 (N_5850,N_2701,N_1399);
nor U5851 (N_5851,N_2274,N_105);
xor U5852 (N_5852,N_3656,N_2522);
nor U5853 (N_5853,N_485,N_2483);
xnor U5854 (N_5854,N_1940,N_419);
xnor U5855 (N_5855,N_2836,N_1869);
or U5856 (N_5856,N_1741,N_1755);
xnor U5857 (N_5857,N_764,N_1643);
and U5858 (N_5858,N_314,N_3838);
xor U5859 (N_5859,N_2234,N_2782);
nor U5860 (N_5860,N_67,N_2413);
nand U5861 (N_5861,N_254,N_376);
xor U5862 (N_5862,N_1554,N_886);
nand U5863 (N_5863,N_3552,N_518);
or U5864 (N_5864,N_538,N_1315);
and U5865 (N_5865,N_1730,N_3366);
and U5866 (N_5866,N_1993,N_3394);
nand U5867 (N_5867,N_1199,N_272);
or U5868 (N_5868,N_3303,N_1123);
xor U5869 (N_5869,N_1585,N_2415);
or U5870 (N_5870,N_3928,N_3123);
or U5871 (N_5871,N_2531,N_3436);
or U5872 (N_5872,N_1627,N_1022);
xor U5873 (N_5873,N_1212,N_2027);
or U5874 (N_5874,N_3195,N_3570);
nor U5875 (N_5875,N_3316,N_779);
nor U5876 (N_5876,N_1369,N_3528);
nand U5877 (N_5877,N_1513,N_166);
xnor U5878 (N_5878,N_2346,N_1065);
and U5879 (N_5879,N_2869,N_2995);
and U5880 (N_5880,N_729,N_611);
or U5881 (N_5881,N_3422,N_1879);
xnor U5882 (N_5882,N_2899,N_1642);
nand U5883 (N_5883,N_790,N_3449);
nor U5884 (N_5884,N_2677,N_3857);
or U5885 (N_5885,N_2838,N_3564);
or U5886 (N_5886,N_1114,N_2434);
nand U5887 (N_5887,N_1134,N_2446);
xor U5888 (N_5888,N_2092,N_1211);
xnor U5889 (N_5889,N_2351,N_666);
xnor U5890 (N_5890,N_2049,N_1972);
xor U5891 (N_5891,N_1649,N_3753);
and U5892 (N_5892,N_271,N_3372);
or U5893 (N_5893,N_1647,N_3154);
nand U5894 (N_5894,N_2282,N_2722);
nor U5895 (N_5895,N_2113,N_6);
and U5896 (N_5896,N_2693,N_3864);
nor U5897 (N_5897,N_2178,N_291);
nor U5898 (N_5898,N_2795,N_3235);
and U5899 (N_5899,N_2626,N_3148);
or U5900 (N_5900,N_3877,N_839);
nor U5901 (N_5901,N_1264,N_3870);
or U5902 (N_5902,N_2441,N_3828);
xor U5903 (N_5903,N_1699,N_2922);
xnor U5904 (N_5904,N_1980,N_660);
or U5905 (N_5905,N_953,N_50);
and U5906 (N_5906,N_1500,N_3459);
or U5907 (N_5907,N_1138,N_2028);
or U5908 (N_5908,N_117,N_1511);
or U5909 (N_5909,N_1328,N_1147);
and U5910 (N_5910,N_2187,N_1488);
nor U5911 (N_5911,N_1066,N_3553);
nand U5912 (N_5912,N_1935,N_3511);
xnor U5913 (N_5913,N_1802,N_2880);
nor U5914 (N_5914,N_784,N_1263);
xnor U5915 (N_5915,N_1622,N_1888);
xnor U5916 (N_5916,N_2969,N_3114);
nand U5917 (N_5917,N_3985,N_1502);
nand U5918 (N_5918,N_2700,N_1441);
or U5919 (N_5919,N_2114,N_393);
xnor U5920 (N_5920,N_1744,N_3293);
nand U5921 (N_5921,N_1950,N_57);
nand U5922 (N_5922,N_2070,N_2461);
xor U5923 (N_5923,N_1455,N_1152);
or U5924 (N_5924,N_539,N_2005);
or U5925 (N_5925,N_1421,N_927);
nor U5926 (N_5926,N_2240,N_1376);
nor U5927 (N_5927,N_2537,N_250);
or U5928 (N_5928,N_3308,N_3613);
or U5929 (N_5929,N_1448,N_903);
nand U5930 (N_5930,N_3236,N_2909);
nor U5931 (N_5931,N_742,N_2238);
and U5932 (N_5932,N_48,N_3294);
and U5933 (N_5933,N_2773,N_1247);
and U5934 (N_5934,N_1558,N_2853);
nand U5935 (N_5935,N_2535,N_2610);
nand U5936 (N_5936,N_3884,N_1775);
nor U5937 (N_5937,N_2174,N_3345);
nor U5938 (N_5938,N_3288,N_3881);
nor U5939 (N_5939,N_3469,N_1693);
or U5940 (N_5940,N_2695,N_3571);
nand U5941 (N_5941,N_3229,N_771);
xor U5942 (N_5942,N_3015,N_2077);
xnor U5943 (N_5943,N_2353,N_258);
nor U5944 (N_5944,N_2118,N_920);
or U5945 (N_5945,N_2800,N_2182);
and U5946 (N_5946,N_2759,N_1103);
or U5947 (N_5947,N_2755,N_1709);
xor U5948 (N_5948,N_1617,N_3187);
or U5949 (N_5949,N_2732,N_2390);
or U5950 (N_5950,N_395,N_1044);
xnor U5951 (N_5951,N_1353,N_2727);
nand U5952 (N_5952,N_12,N_1592);
and U5953 (N_5953,N_711,N_468);
or U5954 (N_5954,N_3133,N_950);
or U5955 (N_5955,N_812,N_1773);
or U5956 (N_5956,N_3551,N_783);
xnor U5957 (N_5957,N_2994,N_2547);
xnor U5958 (N_5958,N_420,N_595);
and U5959 (N_5959,N_740,N_555);
or U5960 (N_5960,N_2757,N_2069);
nor U5961 (N_5961,N_365,N_2046);
nor U5962 (N_5962,N_238,N_1335);
or U5963 (N_5963,N_2189,N_64);
nor U5964 (N_5964,N_2830,N_3021);
and U5965 (N_5965,N_1948,N_2472);
or U5966 (N_5966,N_3874,N_1291);
or U5967 (N_5967,N_3737,N_428);
and U5968 (N_5968,N_881,N_461);
and U5969 (N_5969,N_692,N_1752);
xnor U5970 (N_5970,N_1998,N_1508);
xnor U5971 (N_5971,N_3125,N_2578);
nor U5972 (N_5972,N_144,N_2091);
and U5973 (N_5973,N_491,N_32);
and U5974 (N_5974,N_351,N_3275);
nand U5975 (N_5975,N_3077,N_1162);
nor U5976 (N_5976,N_1221,N_3723);
and U5977 (N_5977,N_2587,N_829);
xnor U5978 (N_5978,N_765,N_2957);
or U5979 (N_5979,N_3036,N_3226);
and U5980 (N_5980,N_1604,N_2948);
xnor U5981 (N_5981,N_3063,N_916);
and U5982 (N_5982,N_3416,N_111);
nor U5983 (N_5983,N_1220,N_1981);
nand U5984 (N_5984,N_1927,N_2890);
and U5985 (N_5985,N_1517,N_2926);
nor U5986 (N_5986,N_3355,N_2516);
nor U5987 (N_5987,N_1745,N_41);
nor U5988 (N_5988,N_3909,N_695);
or U5989 (N_5989,N_3971,N_1027);
nand U5990 (N_5990,N_2498,N_1339);
nand U5991 (N_5991,N_3412,N_1874);
or U5992 (N_5992,N_3249,N_2392);
or U5993 (N_5993,N_1952,N_1983);
nor U5994 (N_5994,N_456,N_3144);
nor U5995 (N_5995,N_1921,N_3335);
and U5996 (N_5996,N_2513,N_1862);
or U5997 (N_5997,N_3452,N_808);
and U5998 (N_5998,N_3175,N_1384);
nor U5999 (N_5999,N_74,N_3041);
xor U6000 (N_6000,N_3432,N_3807);
or U6001 (N_6001,N_692,N_3140);
and U6002 (N_6002,N_2356,N_386);
xor U6003 (N_6003,N_93,N_2650);
nor U6004 (N_6004,N_712,N_3604);
nor U6005 (N_6005,N_2304,N_3144);
xor U6006 (N_6006,N_3059,N_3440);
xor U6007 (N_6007,N_3844,N_3689);
xor U6008 (N_6008,N_1821,N_3687);
and U6009 (N_6009,N_722,N_2959);
nor U6010 (N_6010,N_2870,N_2636);
nor U6011 (N_6011,N_1764,N_1787);
nand U6012 (N_6012,N_1319,N_1956);
nor U6013 (N_6013,N_1157,N_2603);
or U6014 (N_6014,N_355,N_2167);
xnor U6015 (N_6015,N_7,N_1980);
and U6016 (N_6016,N_1616,N_1885);
and U6017 (N_6017,N_2832,N_1537);
nand U6018 (N_6018,N_1586,N_575);
or U6019 (N_6019,N_1436,N_3490);
or U6020 (N_6020,N_1494,N_3622);
and U6021 (N_6021,N_2206,N_382);
nor U6022 (N_6022,N_600,N_2335);
nor U6023 (N_6023,N_2151,N_257);
nor U6024 (N_6024,N_1807,N_3117);
nand U6025 (N_6025,N_211,N_2808);
or U6026 (N_6026,N_3109,N_3357);
or U6027 (N_6027,N_319,N_1117);
nand U6028 (N_6028,N_2752,N_789);
xor U6029 (N_6029,N_237,N_2514);
nor U6030 (N_6030,N_3726,N_2879);
nand U6031 (N_6031,N_2968,N_3166);
or U6032 (N_6032,N_1072,N_3148);
nor U6033 (N_6033,N_1852,N_1055);
or U6034 (N_6034,N_310,N_1721);
nor U6035 (N_6035,N_83,N_1184);
nor U6036 (N_6036,N_1869,N_839);
xnor U6037 (N_6037,N_2964,N_496);
nor U6038 (N_6038,N_2104,N_3102);
xnor U6039 (N_6039,N_469,N_1837);
nand U6040 (N_6040,N_1186,N_62);
xnor U6041 (N_6041,N_2155,N_3196);
xor U6042 (N_6042,N_373,N_2083);
xor U6043 (N_6043,N_2358,N_2934);
xor U6044 (N_6044,N_325,N_109);
or U6045 (N_6045,N_2633,N_847);
or U6046 (N_6046,N_2913,N_25);
nor U6047 (N_6047,N_220,N_2883);
nand U6048 (N_6048,N_2946,N_1819);
and U6049 (N_6049,N_1588,N_3583);
and U6050 (N_6050,N_487,N_3293);
or U6051 (N_6051,N_3135,N_2886);
nand U6052 (N_6052,N_278,N_3235);
or U6053 (N_6053,N_3683,N_1502);
xnor U6054 (N_6054,N_3099,N_910);
xor U6055 (N_6055,N_2954,N_2682);
or U6056 (N_6056,N_2140,N_2271);
nand U6057 (N_6057,N_2057,N_3094);
nand U6058 (N_6058,N_312,N_102);
nand U6059 (N_6059,N_1726,N_2491);
and U6060 (N_6060,N_1599,N_3985);
xnor U6061 (N_6061,N_3338,N_278);
or U6062 (N_6062,N_1387,N_1838);
or U6063 (N_6063,N_3684,N_3424);
or U6064 (N_6064,N_773,N_2045);
and U6065 (N_6065,N_599,N_2513);
nor U6066 (N_6066,N_2751,N_1043);
xor U6067 (N_6067,N_1,N_1173);
nor U6068 (N_6068,N_2466,N_602);
and U6069 (N_6069,N_412,N_1005);
xnor U6070 (N_6070,N_3135,N_3861);
and U6071 (N_6071,N_735,N_3900);
and U6072 (N_6072,N_3331,N_2068);
xor U6073 (N_6073,N_2039,N_459);
nor U6074 (N_6074,N_2384,N_1080);
and U6075 (N_6075,N_1347,N_543);
or U6076 (N_6076,N_1749,N_3917);
and U6077 (N_6077,N_2127,N_1442);
and U6078 (N_6078,N_2238,N_3792);
xor U6079 (N_6079,N_1948,N_3988);
nor U6080 (N_6080,N_3716,N_1055);
nor U6081 (N_6081,N_1588,N_414);
nor U6082 (N_6082,N_1096,N_3463);
nand U6083 (N_6083,N_3814,N_785);
nand U6084 (N_6084,N_1260,N_2283);
nor U6085 (N_6085,N_182,N_215);
or U6086 (N_6086,N_193,N_928);
xnor U6087 (N_6087,N_2035,N_2238);
xnor U6088 (N_6088,N_2964,N_1904);
and U6089 (N_6089,N_469,N_3741);
and U6090 (N_6090,N_1943,N_1462);
xor U6091 (N_6091,N_3544,N_1387);
and U6092 (N_6092,N_1530,N_822);
or U6093 (N_6093,N_1812,N_843);
and U6094 (N_6094,N_963,N_3626);
nor U6095 (N_6095,N_887,N_579);
nor U6096 (N_6096,N_3685,N_1792);
nor U6097 (N_6097,N_1762,N_2570);
nand U6098 (N_6098,N_1163,N_1112);
or U6099 (N_6099,N_3466,N_1965);
xnor U6100 (N_6100,N_3462,N_2143);
nand U6101 (N_6101,N_1757,N_1440);
or U6102 (N_6102,N_2413,N_3923);
or U6103 (N_6103,N_3694,N_566);
nor U6104 (N_6104,N_3420,N_2894);
xnor U6105 (N_6105,N_2024,N_1312);
nor U6106 (N_6106,N_1704,N_3763);
or U6107 (N_6107,N_3585,N_3550);
or U6108 (N_6108,N_2286,N_119);
nor U6109 (N_6109,N_1116,N_3171);
or U6110 (N_6110,N_2166,N_1244);
and U6111 (N_6111,N_3545,N_3808);
and U6112 (N_6112,N_3945,N_3441);
nor U6113 (N_6113,N_1546,N_3370);
or U6114 (N_6114,N_541,N_3421);
and U6115 (N_6115,N_1344,N_3697);
and U6116 (N_6116,N_2822,N_2300);
xnor U6117 (N_6117,N_2309,N_318);
nor U6118 (N_6118,N_3804,N_3127);
nand U6119 (N_6119,N_1625,N_1609);
xnor U6120 (N_6120,N_931,N_538);
nand U6121 (N_6121,N_297,N_2821);
or U6122 (N_6122,N_1949,N_1199);
and U6123 (N_6123,N_105,N_3787);
xor U6124 (N_6124,N_2403,N_3988);
nand U6125 (N_6125,N_3335,N_1872);
or U6126 (N_6126,N_1468,N_3130);
nand U6127 (N_6127,N_3052,N_1400);
and U6128 (N_6128,N_3314,N_2253);
xor U6129 (N_6129,N_3962,N_2364);
and U6130 (N_6130,N_2233,N_1031);
nor U6131 (N_6131,N_970,N_3402);
xnor U6132 (N_6132,N_604,N_298);
nand U6133 (N_6133,N_1823,N_943);
and U6134 (N_6134,N_2575,N_3727);
and U6135 (N_6135,N_336,N_2852);
nand U6136 (N_6136,N_942,N_574);
nor U6137 (N_6137,N_1222,N_456);
nor U6138 (N_6138,N_509,N_3397);
or U6139 (N_6139,N_1211,N_90);
or U6140 (N_6140,N_3139,N_741);
and U6141 (N_6141,N_3379,N_52);
nand U6142 (N_6142,N_774,N_2052);
nand U6143 (N_6143,N_1450,N_1400);
xnor U6144 (N_6144,N_2985,N_2063);
or U6145 (N_6145,N_3653,N_3279);
or U6146 (N_6146,N_754,N_922);
and U6147 (N_6147,N_1111,N_395);
and U6148 (N_6148,N_1381,N_1948);
or U6149 (N_6149,N_1101,N_2916);
and U6150 (N_6150,N_2847,N_233);
or U6151 (N_6151,N_2259,N_2345);
nor U6152 (N_6152,N_390,N_2073);
and U6153 (N_6153,N_1246,N_3940);
nor U6154 (N_6154,N_2606,N_1045);
nor U6155 (N_6155,N_584,N_1163);
or U6156 (N_6156,N_3962,N_206);
nand U6157 (N_6157,N_2610,N_3748);
or U6158 (N_6158,N_376,N_3589);
nor U6159 (N_6159,N_3434,N_1583);
or U6160 (N_6160,N_1078,N_1192);
nor U6161 (N_6161,N_1811,N_178);
xor U6162 (N_6162,N_494,N_1891);
nor U6163 (N_6163,N_556,N_3300);
nand U6164 (N_6164,N_1012,N_1480);
xnor U6165 (N_6165,N_2610,N_955);
nand U6166 (N_6166,N_1320,N_436);
nand U6167 (N_6167,N_1440,N_1108);
or U6168 (N_6168,N_1814,N_1640);
or U6169 (N_6169,N_600,N_472);
nor U6170 (N_6170,N_2187,N_2411);
nand U6171 (N_6171,N_75,N_3101);
or U6172 (N_6172,N_1167,N_2451);
xor U6173 (N_6173,N_1579,N_1375);
nor U6174 (N_6174,N_126,N_661);
nor U6175 (N_6175,N_2719,N_599);
xor U6176 (N_6176,N_2249,N_3118);
nor U6177 (N_6177,N_1702,N_1652);
nand U6178 (N_6178,N_3621,N_340);
nor U6179 (N_6179,N_602,N_3441);
or U6180 (N_6180,N_3884,N_644);
xnor U6181 (N_6181,N_3008,N_1037);
xnor U6182 (N_6182,N_2645,N_2945);
and U6183 (N_6183,N_2812,N_2180);
nor U6184 (N_6184,N_292,N_1941);
nor U6185 (N_6185,N_3213,N_1652);
nand U6186 (N_6186,N_1819,N_2569);
nand U6187 (N_6187,N_3149,N_3992);
or U6188 (N_6188,N_2396,N_2930);
xor U6189 (N_6189,N_3721,N_1608);
nand U6190 (N_6190,N_1144,N_1417);
and U6191 (N_6191,N_1318,N_816);
xor U6192 (N_6192,N_2714,N_1555);
and U6193 (N_6193,N_2719,N_2536);
and U6194 (N_6194,N_1730,N_1234);
xnor U6195 (N_6195,N_159,N_757);
nor U6196 (N_6196,N_2631,N_2394);
or U6197 (N_6197,N_2001,N_648);
xor U6198 (N_6198,N_3452,N_2791);
nand U6199 (N_6199,N_3489,N_1172);
xnor U6200 (N_6200,N_2224,N_1658);
or U6201 (N_6201,N_2731,N_1870);
nor U6202 (N_6202,N_808,N_2697);
or U6203 (N_6203,N_1008,N_3043);
or U6204 (N_6204,N_2655,N_2097);
and U6205 (N_6205,N_1279,N_1296);
xor U6206 (N_6206,N_2512,N_617);
xnor U6207 (N_6207,N_3162,N_3585);
xor U6208 (N_6208,N_927,N_471);
and U6209 (N_6209,N_1755,N_401);
and U6210 (N_6210,N_507,N_3640);
xor U6211 (N_6211,N_1,N_1378);
or U6212 (N_6212,N_3805,N_1142);
nor U6213 (N_6213,N_1520,N_704);
xor U6214 (N_6214,N_1802,N_268);
or U6215 (N_6215,N_3729,N_2956);
nor U6216 (N_6216,N_370,N_3479);
and U6217 (N_6217,N_3714,N_162);
xor U6218 (N_6218,N_3423,N_1232);
nor U6219 (N_6219,N_451,N_2078);
nand U6220 (N_6220,N_2649,N_1213);
nand U6221 (N_6221,N_1269,N_762);
nand U6222 (N_6222,N_2183,N_3621);
xnor U6223 (N_6223,N_2444,N_627);
or U6224 (N_6224,N_3681,N_1162);
xnor U6225 (N_6225,N_785,N_3403);
xnor U6226 (N_6226,N_1598,N_2900);
nor U6227 (N_6227,N_2913,N_1593);
nor U6228 (N_6228,N_3465,N_3517);
and U6229 (N_6229,N_1764,N_476);
nand U6230 (N_6230,N_399,N_3062);
xnor U6231 (N_6231,N_3006,N_5);
nor U6232 (N_6232,N_2029,N_3029);
nor U6233 (N_6233,N_289,N_583);
nand U6234 (N_6234,N_3096,N_3459);
or U6235 (N_6235,N_20,N_1266);
xnor U6236 (N_6236,N_3260,N_3344);
nand U6237 (N_6237,N_793,N_900);
nand U6238 (N_6238,N_517,N_841);
xnor U6239 (N_6239,N_2382,N_2311);
and U6240 (N_6240,N_144,N_2331);
and U6241 (N_6241,N_3489,N_2214);
xnor U6242 (N_6242,N_2836,N_3122);
nand U6243 (N_6243,N_3092,N_1654);
nor U6244 (N_6244,N_3476,N_2420);
or U6245 (N_6245,N_2039,N_1842);
nor U6246 (N_6246,N_187,N_2715);
nand U6247 (N_6247,N_943,N_2808);
or U6248 (N_6248,N_697,N_1366);
and U6249 (N_6249,N_1068,N_2571);
and U6250 (N_6250,N_710,N_954);
nand U6251 (N_6251,N_991,N_2770);
nor U6252 (N_6252,N_2087,N_630);
nand U6253 (N_6253,N_11,N_1159);
nor U6254 (N_6254,N_708,N_686);
nor U6255 (N_6255,N_64,N_3988);
and U6256 (N_6256,N_1160,N_2037);
and U6257 (N_6257,N_601,N_1962);
or U6258 (N_6258,N_2236,N_3434);
xor U6259 (N_6259,N_3268,N_1158);
nor U6260 (N_6260,N_3165,N_300);
xor U6261 (N_6261,N_2747,N_1895);
nor U6262 (N_6262,N_28,N_3834);
nand U6263 (N_6263,N_1512,N_3398);
nor U6264 (N_6264,N_3327,N_3896);
xnor U6265 (N_6265,N_3549,N_1556);
nand U6266 (N_6266,N_2730,N_182);
nand U6267 (N_6267,N_83,N_57);
nor U6268 (N_6268,N_301,N_1114);
nor U6269 (N_6269,N_1199,N_1021);
or U6270 (N_6270,N_985,N_2186);
and U6271 (N_6271,N_3775,N_563);
and U6272 (N_6272,N_90,N_2323);
nor U6273 (N_6273,N_1997,N_572);
nor U6274 (N_6274,N_1842,N_3644);
xor U6275 (N_6275,N_1807,N_1031);
nand U6276 (N_6276,N_1457,N_719);
nor U6277 (N_6277,N_3038,N_3648);
nor U6278 (N_6278,N_1923,N_3440);
or U6279 (N_6279,N_440,N_181);
nor U6280 (N_6280,N_2798,N_2499);
or U6281 (N_6281,N_3697,N_3834);
and U6282 (N_6282,N_1663,N_3693);
and U6283 (N_6283,N_1544,N_3136);
nand U6284 (N_6284,N_2062,N_2912);
and U6285 (N_6285,N_1745,N_3455);
nor U6286 (N_6286,N_3674,N_1139);
and U6287 (N_6287,N_678,N_939);
and U6288 (N_6288,N_3948,N_359);
xnor U6289 (N_6289,N_3664,N_389);
nor U6290 (N_6290,N_3887,N_3865);
nor U6291 (N_6291,N_3490,N_1621);
nor U6292 (N_6292,N_3475,N_246);
or U6293 (N_6293,N_1776,N_1246);
nand U6294 (N_6294,N_347,N_1305);
or U6295 (N_6295,N_400,N_2485);
nand U6296 (N_6296,N_2624,N_210);
xor U6297 (N_6297,N_1911,N_3276);
xor U6298 (N_6298,N_3029,N_1009);
or U6299 (N_6299,N_1740,N_2910);
and U6300 (N_6300,N_3052,N_1880);
xnor U6301 (N_6301,N_903,N_1504);
nand U6302 (N_6302,N_1536,N_240);
nor U6303 (N_6303,N_29,N_1894);
xor U6304 (N_6304,N_1885,N_1076);
or U6305 (N_6305,N_1807,N_528);
and U6306 (N_6306,N_1661,N_3581);
and U6307 (N_6307,N_1694,N_3632);
xnor U6308 (N_6308,N_3515,N_1531);
nand U6309 (N_6309,N_420,N_3310);
nor U6310 (N_6310,N_2648,N_2359);
or U6311 (N_6311,N_3926,N_3067);
nor U6312 (N_6312,N_490,N_2077);
and U6313 (N_6313,N_3488,N_1766);
nand U6314 (N_6314,N_529,N_1463);
or U6315 (N_6315,N_1731,N_1080);
xnor U6316 (N_6316,N_2905,N_3764);
xnor U6317 (N_6317,N_1541,N_73);
or U6318 (N_6318,N_1987,N_2238);
and U6319 (N_6319,N_698,N_3356);
or U6320 (N_6320,N_3721,N_21);
nand U6321 (N_6321,N_2859,N_3549);
xor U6322 (N_6322,N_3661,N_1259);
nor U6323 (N_6323,N_1114,N_2374);
xnor U6324 (N_6324,N_535,N_3089);
nand U6325 (N_6325,N_2162,N_2849);
or U6326 (N_6326,N_2563,N_1960);
xnor U6327 (N_6327,N_2290,N_3369);
or U6328 (N_6328,N_1350,N_904);
nand U6329 (N_6329,N_2675,N_643);
or U6330 (N_6330,N_3014,N_1340);
nand U6331 (N_6331,N_3920,N_2594);
nor U6332 (N_6332,N_1296,N_2323);
xor U6333 (N_6333,N_2030,N_1581);
or U6334 (N_6334,N_284,N_2899);
xnor U6335 (N_6335,N_361,N_752);
xor U6336 (N_6336,N_2754,N_3428);
nand U6337 (N_6337,N_1878,N_266);
nor U6338 (N_6338,N_2212,N_2127);
and U6339 (N_6339,N_887,N_2481);
or U6340 (N_6340,N_3263,N_1860);
or U6341 (N_6341,N_2277,N_1970);
nand U6342 (N_6342,N_1926,N_872);
or U6343 (N_6343,N_1093,N_3419);
nor U6344 (N_6344,N_3231,N_3398);
nand U6345 (N_6345,N_2426,N_1812);
and U6346 (N_6346,N_539,N_3921);
and U6347 (N_6347,N_3405,N_2624);
nand U6348 (N_6348,N_1487,N_243);
nand U6349 (N_6349,N_3292,N_2068);
nand U6350 (N_6350,N_718,N_3018);
xnor U6351 (N_6351,N_64,N_1807);
and U6352 (N_6352,N_1118,N_643);
nor U6353 (N_6353,N_2922,N_2573);
and U6354 (N_6354,N_3567,N_1758);
xnor U6355 (N_6355,N_544,N_611);
nand U6356 (N_6356,N_775,N_1608);
xnor U6357 (N_6357,N_634,N_224);
or U6358 (N_6358,N_3354,N_2607);
nand U6359 (N_6359,N_1064,N_1371);
or U6360 (N_6360,N_1537,N_2297);
nor U6361 (N_6361,N_2514,N_3007);
and U6362 (N_6362,N_3076,N_3255);
xor U6363 (N_6363,N_2593,N_388);
and U6364 (N_6364,N_2836,N_3401);
xor U6365 (N_6365,N_564,N_597);
nand U6366 (N_6366,N_1766,N_574);
nand U6367 (N_6367,N_3339,N_2623);
or U6368 (N_6368,N_914,N_3667);
nand U6369 (N_6369,N_1893,N_1809);
nand U6370 (N_6370,N_854,N_3519);
nor U6371 (N_6371,N_1637,N_2883);
or U6372 (N_6372,N_997,N_1174);
nand U6373 (N_6373,N_3575,N_3649);
xor U6374 (N_6374,N_3446,N_528);
or U6375 (N_6375,N_169,N_1369);
or U6376 (N_6376,N_1231,N_2327);
and U6377 (N_6377,N_3134,N_3309);
or U6378 (N_6378,N_1854,N_420);
nand U6379 (N_6379,N_1857,N_484);
and U6380 (N_6380,N_3478,N_3990);
or U6381 (N_6381,N_3608,N_1915);
xnor U6382 (N_6382,N_2533,N_837);
xor U6383 (N_6383,N_896,N_2029);
or U6384 (N_6384,N_1607,N_3012);
and U6385 (N_6385,N_3817,N_2495);
nor U6386 (N_6386,N_110,N_314);
and U6387 (N_6387,N_2211,N_3441);
and U6388 (N_6388,N_1092,N_3097);
nor U6389 (N_6389,N_11,N_2202);
or U6390 (N_6390,N_1706,N_2169);
nand U6391 (N_6391,N_1337,N_597);
xnor U6392 (N_6392,N_3402,N_559);
nand U6393 (N_6393,N_3769,N_2325);
and U6394 (N_6394,N_3718,N_3583);
and U6395 (N_6395,N_2885,N_336);
nand U6396 (N_6396,N_1047,N_3707);
nor U6397 (N_6397,N_2932,N_1015);
nand U6398 (N_6398,N_1392,N_2453);
nor U6399 (N_6399,N_1975,N_162);
or U6400 (N_6400,N_2481,N_5);
or U6401 (N_6401,N_2325,N_874);
xnor U6402 (N_6402,N_3637,N_3359);
or U6403 (N_6403,N_1133,N_2770);
nor U6404 (N_6404,N_2038,N_782);
nand U6405 (N_6405,N_1003,N_1084);
or U6406 (N_6406,N_247,N_1006);
and U6407 (N_6407,N_2049,N_3860);
or U6408 (N_6408,N_698,N_2471);
xor U6409 (N_6409,N_3023,N_1253);
or U6410 (N_6410,N_1518,N_3995);
and U6411 (N_6411,N_931,N_2086);
nor U6412 (N_6412,N_1598,N_950);
nand U6413 (N_6413,N_2490,N_999);
nor U6414 (N_6414,N_3280,N_3691);
xor U6415 (N_6415,N_2957,N_3074);
or U6416 (N_6416,N_811,N_3510);
xnor U6417 (N_6417,N_2714,N_2243);
or U6418 (N_6418,N_3147,N_545);
and U6419 (N_6419,N_2898,N_2805);
nor U6420 (N_6420,N_3533,N_2254);
xor U6421 (N_6421,N_2718,N_3294);
or U6422 (N_6422,N_800,N_859);
xor U6423 (N_6423,N_3062,N_821);
xor U6424 (N_6424,N_593,N_2651);
xor U6425 (N_6425,N_3117,N_3433);
and U6426 (N_6426,N_2116,N_3671);
and U6427 (N_6427,N_1812,N_1760);
or U6428 (N_6428,N_351,N_3334);
and U6429 (N_6429,N_936,N_1900);
nand U6430 (N_6430,N_1690,N_219);
nor U6431 (N_6431,N_93,N_231);
nor U6432 (N_6432,N_2658,N_2293);
or U6433 (N_6433,N_2436,N_656);
xnor U6434 (N_6434,N_1004,N_823);
nor U6435 (N_6435,N_2051,N_2663);
nor U6436 (N_6436,N_3722,N_3805);
and U6437 (N_6437,N_3382,N_845);
nor U6438 (N_6438,N_93,N_2730);
xor U6439 (N_6439,N_247,N_950);
nand U6440 (N_6440,N_266,N_1103);
nor U6441 (N_6441,N_330,N_1881);
xnor U6442 (N_6442,N_1542,N_1124);
or U6443 (N_6443,N_474,N_399);
and U6444 (N_6444,N_1675,N_2559);
xnor U6445 (N_6445,N_1885,N_474);
nand U6446 (N_6446,N_679,N_1566);
xnor U6447 (N_6447,N_1995,N_918);
nor U6448 (N_6448,N_3920,N_3086);
or U6449 (N_6449,N_3078,N_1122);
and U6450 (N_6450,N_1898,N_1324);
nand U6451 (N_6451,N_3070,N_2096);
and U6452 (N_6452,N_2069,N_2904);
xnor U6453 (N_6453,N_3461,N_417);
nand U6454 (N_6454,N_3047,N_96);
and U6455 (N_6455,N_533,N_3251);
and U6456 (N_6456,N_1528,N_3781);
nor U6457 (N_6457,N_446,N_2913);
xor U6458 (N_6458,N_1752,N_138);
nor U6459 (N_6459,N_3943,N_373);
nor U6460 (N_6460,N_2339,N_790);
nand U6461 (N_6461,N_3785,N_1781);
nor U6462 (N_6462,N_3136,N_587);
or U6463 (N_6463,N_1215,N_1406);
xnor U6464 (N_6464,N_3859,N_2204);
or U6465 (N_6465,N_3547,N_566);
xnor U6466 (N_6466,N_1973,N_2544);
nor U6467 (N_6467,N_1698,N_1460);
or U6468 (N_6468,N_163,N_3925);
nor U6469 (N_6469,N_3792,N_3912);
xnor U6470 (N_6470,N_3392,N_3478);
nand U6471 (N_6471,N_994,N_569);
nor U6472 (N_6472,N_2846,N_3112);
and U6473 (N_6473,N_2169,N_1158);
or U6474 (N_6474,N_480,N_2243);
nand U6475 (N_6475,N_835,N_571);
or U6476 (N_6476,N_215,N_1524);
xnor U6477 (N_6477,N_2835,N_2932);
and U6478 (N_6478,N_612,N_3193);
and U6479 (N_6479,N_2879,N_896);
and U6480 (N_6480,N_3321,N_1551);
and U6481 (N_6481,N_3762,N_3851);
and U6482 (N_6482,N_615,N_2120);
nor U6483 (N_6483,N_3843,N_822);
and U6484 (N_6484,N_33,N_2457);
or U6485 (N_6485,N_2615,N_3521);
and U6486 (N_6486,N_2828,N_828);
and U6487 (N_6487,N_1234,N_3692);
or U6488 (N_6488,N_2847,N_2540);
nor U6489 (N_6489,N_2071,N_360);
nand U6490 (N_6490,N_512,N_1226);
or U6491 (N_6491,N_2884,N_1233);
nand U6492 (N_6492,N_1738,N_1588);
or U6493 (N_6493,N_1578,N_954);
nand U6494 (N_6494,N_2386,N_2243);
nand U6495 (N_6495,N_64,N_2874);
or U6496 (N_6496,N_632,N_634);
nand U6497 (N_6497,N_2970,N_3374);
xor U6498 (N_6498,N_1159,N_937);
nand U6499 (N_6499,N_2550,N_2861);
and U6500 (N_6500,N_2448,N_1677);
xnor U6501 (N_6501,N_812,N_177);
and U6502 (N_6502,N_3154,N_1419);
and U6503 (N_6503,N_897,N_2048);
nand U6504 (N_6504,N_370,N_2011);
and U6505 (N_6505,N_1008,N_971);
or U6506 (N_6506,N_1435,N_2236);
and U6507 (N_6507,N_2409,N_139);
nand U6508 (N_6508,N_2684,N_2498);
and U6509 (N_6509,N_2246,N_1710);
and U6510 (N_6510,N_750,N_3249);
and U6511 (N_6511,N_2893,N_1850);
nor U6512 (N_6512,N_1720,N_3888);
or U6513 (N_6513,N_524,N_3853);
nor U6514 (N_6514,N_3111,N_453);
xor U6515 (N_6515,N_546,N_1932);
nor U6516 (N_6516,N_1214,N_1386);
and U6517 (N_6517,N_168,N_946);
xor U6518 (N_6518,N_771,N_3869);
nand U6519 (N_6519,N_1746,N_1720);
nand U6520 (N_6520,N_1745,N_375);
and U6521 (N_6521,N_2958,N_1614);
xnor U6522 (N_6522,N_1477,N_2437);
and U6523 (N_6523,N_3928,N_2596);
nor U6524 (N_6524,N_2287,N_2207);
xor U6525 (N_6525,N_2343,N_3119);
nor U6526 (N_6526,N_1534,N_1948);
xor U6527 (N_6527,N_1563,N_3955);
nor U6528 (N_6528,N_3275,N_745);
xnor U6529 (N_6529,N_279,N_1691);
or U6530 (N_6530,N_450,N_793);
and U6531 (N_6531,N_3970,N_3199);
xor U6532 (N_6532,N_2299,N_2394);
and U6533 (N_6533,N_325,N_99);
or U6534 (N_6534,N_2432,N_2128);
or U6535 (N_6535,N_2084,N_1327);
or U6536 (N_6536,N_3435,N_465);
xnor U6537 (N_6537,N_1629,N_730);
and U6538 (N_6538,N_1519,N_3355);
nor U6539 (N_6539,N_2425,N_3689);
xor U6540 (N_6540,N_2636,N_2345);
nor U6541 (N_6541,N_1872,N_422);
nand U6542 (N_6542,N_3017,N_3105);
or U6543 (N_6543,N_1786,N_2326);
and U6544 (N_6544,N_1890,N_2583);
or U6545 (N_6545,N_2694,N_634);
or U6546 (N_6546,N_2840,N_1816);
nand U6547 (N_6547,N_1074,N_3633);
nor U6548 (N_6548,N_2665,N_1798);
and U6549 (N_6549,N_3859,N_1148);
nor U6550 (N_6550,N_2520,N_3863);
and U6551 (N_6551,N_1314,N_970);
nand U6552 (N_6552,N_530,N_810);
nand U6553 (N_6553,N_1822,N_2056);
nand U6554 (N_6554,N_2349,N_2299);
and U6555 (N_6555,N_2529,N_1062);
nor U6556 (N_6556,N_3451,N_3371);
nor U6557 (N_6557,N_2826,N_1964);
nor U6558 (N_6558,N_3164,N_958);
nor U6559 (N_6559,N_1874,N_1509);
nand U6560 (N_6560,N_216,N_3046);
nor U6561 (N_6561,N_1612,N_3696);
or U6562 (N_6562,N_1695,N_3993);
xor U6563 (N_6563,N_3852,N_3364);
and U6564 (N_6564,N_149,N_3896);
nor U6565 (N_6565,N_132,N_3084);
or U6566 (N_6566,N_2243,N_723);
nor U6567 (N_6567,N_678,N_3955);
nand U6568 (N_6568,N_3419,N_2553);
xnor U6569 (N_6569,N_2613,N_3420);
nor U6570 (N_6570,N_1182,N_1876);
xor U6571 (N_6571,N_3944,N_3338);
or U6572 (N_6572,N_1190,N_1283);
nand U6573 (N_6573,N_2692,N_3585);
and U6574 (N_6574,N_766,N_3878);
nand U6575 (N_6575,N_2936,N_2986);
xor U6576 (N_6576,N_1239,N_3529);
and U6577 (N_6577,N_1439,N_125);
nand U6578 (N_6578,N_2179,N_1346);
or U6579 (N_6579,N_2679,N_1921);
or U6580 (N_6580,N_3684,N_3807);
nor U6581 (N_6581,N_3712,N_286);
xnor U6582 (N_6582,N_3446,N_784);
and U6583 (N_6583,N_3115,N_1531);
nand U6584 (N_6584,N_1506,N_688);
or U6585 (N_6585,N_1348,N_2988);
and U6586 (N_6586,N_1153,N_1273);
xor U6587 (N_6587,N_2610,N_3705);
xnor U6588 (N_6588,N_277,N_416);
and U6589 (N_6589,N_2881,N_8);
nand U6590 (N_6590,N_1187,N_236);
xnor U6591 (N_6591,N_1880,N_1850);
xnor U6592 (N_6592,N_3295,N_3561);
nand U6593 (N_6593,N_2783,N_1721);
and U6594 (N_6594,N_1520,N_2339);
and U6595 (N_6595,N_2443,N_1432);
nor U6596 (N_6596,N_1421,N_2252);
and U6597 (N_6597,N_1216,N_2974);
and U6598 (N_6598,N_2284,N_3965);
xnor U6599 (N_6599,N_1540,N_3387);
and U6600 (N_6600,N_3024,N_3041);
and U6601 (N_6601,N_3363,N_495);
or U6602 (N_6602,N_2760,N_3273);
or U6603 (N_6603,N_1289,N_736);
nand U6604 (N_6604,N_2023,N_1736);
nor U6605 (N_6605,N_888,N_1917);
and U6606 (N_6606,N_3683,N_2348);
and U6607 (N_6607,N_3391,N_1358);
nand U6608 (N_6608,N_2152,N_56);
nand U6609 (N_6609,N_2040,N_1361);
or U6610 (N_6610,N_2497,N_123);
xnor U6611 (N_6611,N_378,N_2450);
nor U6612 (N_6612,N_2754,N_157);
and U6613 (N_6613,N_3861,N_3082);
or U6614 (N_6614,N_324,N_2921);
or U6615 (N_6615,N_3374,N_3126);
or U6616 (N_6616,N_508,N_2063);
nand U6617 (N_6617,N_3561,N_1791);
nand U6618 (N_6618,N_2962,N_253);
nor U6619 (N_6619,N_1416,N_1701);
xor U6620 (N_6620,N_3460,N_2119);
nor U6621 (N_6621,N_3471,N_2398);
xnor U6622 (N_6622,N_2079,N_173);
or U6623 (N_6623,N_3322,N_2060);
or U6624 (N_6624,N_1111,N_1441);
or U6625 (N_6625,N_2377,N_1737);
nor U6626 (N_6626,N_3103,N_2571);
nand U6627 (N_6627,N_3796,N_93);
nand U6628 (N_6628,N_507,N_401);
nor U6629 (N_6629,N_25,N_201);
and U6630 (N_6630,N_2442,N_835);
xor U6631 (N_6631,N_869,N_1455);
nand U6632 (N_6632,N_3416,N_818);
and U6633 (N_6633,N_984,N_221);
xnor U6634 (N_6634,N_1776,N_1445);
and U6635 (N_6635,N_3664,N_2364);
nand U6636 (N_6636,N_1276,N_1280);
nand U6637 (N_6637,N_754,N_1488);
or U6638 (N_6638,N_1012,N_1573);
nor U6639 (N_6639,N_2846,N_3658);
nor U6640 (N_6640,N_1019,N_2820);
and U6641 (N_6641,N_144,N_1847);
xor U6642 (N_6642,N_2803,N_3457);
xnor U6643 (N_6643,N_1223,N_3256);
nor U6644 (N_6644,N_1590,N_1227);
or U6645 (N_6645,N_1754,N_2824);
nand U6646 (N_6646,N_3740,N_3447);
nor U6647 (N_6647,N_3999,N_2090);
nand U6648 (N_6648,N_1834,N_1124);
nor U6649 (N_6649,N_3368,N_743);
nor U6650 (N_6650,N_735,N_2204);
and U6651 (N_6651,N_3909,N_2524);
or U6652 (N_6652,N_2750,N_2240);
nor U6653 (N_6653,N_935,N_1242);
nand U6654 (N_6654,N_617,N_782);
xor U6655 (N_6655,N_1228,N_2915);
nor U6656 (N_6656,N_2263,N_3240);
nor U6657 (N_6657,N_1746,N_3520);
or U6658 (N_6658,N_2682,N_3113);
nor U6659 (N_6659,N_3019,N_3710);
and U6660 (N_6660,N_2510,N_1516);
or U6661 (N_6661,N_2676,N_110);
or U6662 (N_6662,N_1494,N_339);
xor U6663 (N_6663,N_2180,N_2664);
or U6664 (N_6664,N_3276,N_273);
nor U6665 (N_6665,N_1582,N_911);
nand U6666 (N_6666,N_624,N_325);
nand U6667 (N_6667,N_3283,N_3432);
xor U6668 (N_6668,N_715,N_2162);
nand U6669 (N_6669,N_465,N_2199);
xnor U6670 (N_6670,N_1912,N_2408);
or U6671 (N_6671,N_2230,N_339);
and U6672 (N_6672,N_2712,N_3391);
xnor U6673 (N_6673,N_658,N_680);
nor U6674 (N_6674,N_3844,N_3920);
and U6675 (N_6675,N_2799,N_1477);
and U6676 (N_6676,N_3270,N_3349);
or U6677 (N_6677,N_392,N_2901);
and U6678 (N_6678,N_2613,N_3814);
or U6679 (N_6679,N_1457,N_2846);
xor U6680 (N_6680,N_2718,N_2427);
nand U6681 (N_6681,N_1704,N_2722);
nor U6682 (N_6682,N_299,N_396);
and U6683 (N_6683,N_2318,N_1655);
nor U6684 (N_6684,N_2021,N_1586);
and U6685 (N_6685,N_3277,N_2992);
nand U6686 (N_6686,N_3529,N_1949);
and U6687 (N_6687,N_1219,N_2769);
or U6688 (N_6688,N_385,N_1122);
and U6689 (N_6689,N_3360,N_3916);
nor U6690 (N_6690,N_984,N_630);
or U6691 (N_6691,N_3949,N_2915);
nand U6692 (N_6692,N_2703,N_1863);
xor U6693 (N_6693,N_1631,N_3676);
or U6694 (N_6694,N_3776,N_1003);
nor U6695 (N_6695,N_38,N_2129);
and U6696 (N_6696,N_1749,N_198);
nor U6697 (N_6697,N_288,N_1408);
or U6698 (N_6698,N_3770,N_3809);
xor U6699 (N_6699,N_1463,N_1843);
xnor U6700 (N_6700,N_3847,N_393);
nor U6701 (N_6701,N_2372,N_1);
nor U6702 (N_6702,N_3927,N_2649);
xor U6703 (N_6703,N_476,N_175);
xor U6704 (N_6704,N_474,N_3427);
nand U6705 (N_6705,N_2992,N_1162);
and U6706 (N_6706,N_209,N_3043);
and U6707 (N_6707,N_941,N_1207);
and U6708 (N_6708,N_1834,N_1319);
xor U6709 (N_6709,N_1903,N_2361);
and U6710 (N_6710,N_344,N_1137);
nand U6711 (N_6711,N_1108,N_1552);
xor U6712 (N_6712,N_1647,N_656);
and U6713 (N_6713,N_3938,N_1849);
and U6714 (N_6714,N_2238,N_3931);
or U6715 (N_6715,N_1601,N_3367);
nand U6716 (N_6716,N_1123,N_3804);
nor U6717 (N_6717,N_868,N_815);
nand U6718 (N_6718,N_2391,N_1737);
and U6719 (N_6719,N_1992,N_1326);
and U6720 (N_6720,N_395,N_641);
and U6721 (N_6721,N_104,N_3977);
or U6722 (N_6722,N_778,N_2846);
xor U6723 (N_6723,N_1190,N_2173);
nor U6724 (N_6724,N_941,N_10);
and U6725 (N_6725,N_561,N_1110);
nand U6726 (N_6726,N_3001,N_2192);
and U6727 (N_6727,N_1686,N_2166);
or U6728 (N_6728,N_2254,N_1196);
or U6729 (N_6729,N_3226,N_2295);
nand U6730 (N_6730,N_1489,N_1028);
nand U6731 (N_6731,N_1738,N_953);
nor U6732 (N_6732,N_236,N_2956);
nor U6733 (N_6733,N_1248,N_1268);
nor U6734 (N_6734,N_599,N_112);
nor U6735 (N_6735,N_3406,N_55);
xnor U6736 (N_6736,N_2498,N_3425);
xnor U6737 (N_6737,N_272,N_617);
nor U6738 (N_6738,N_152,N_206);
nand U6739 (N_6739,N_1113,N_141);
and U6740 (N_6740,N_2396,N_2313);
or U6741 (N_6741,N_541,N_615);
and U6742 (N_6742,N_2645,N_2404);
nor U6743 (N_6743,N_1662,N_2190);
nand U6744 (N_6744,N_2199,N_3267);
nor U6745 (N_6745,N_1613,N_91);
and U6746 (N_6746,N_1567,N_1334);
or U6747 (N_6747,N_3238,N_1924);
nor U6748 (N_6748,N_1015,N_568);
nor U6749 (N_6749,N_3319,N_766);
xnor U6750 (N_6750,N_2683,N_1577);
or U6751 (N_6751,N_1724,N_2822);
and U6752 (N_6752,N_1434,N_2156);
nand U6753 (N_6753,N_887,N_1954);
and U6754 (N_6754,N_3977,N_3004);
nor U6755 (N_6755,N_2555,N_77);
and U6756 (N_6756,N_2332,N_2535);
xor U6757 (N_6757,N_1656,N_3435);
nand U6758 (N_6758,N_3433,N_452);
xor U6759 (N_6759,N_1290,N_2072);
or U6760 (N_6760,N_3359,N_3154);
or U6761 (N_6761,N_3227,N_3808);
or U6762 (N_6762,N_377,N_3134);
nand U6763 (N_6763,N_2816,N_1686);
and U6764 (N_6764,N_234,N_394);
nand U6765 (N_6765,N_1533,N_3991);
nor U6766 (N_6766,N_735,N_675);
or U6767 (N_6767,N_3542,N_1323);
nand U6768 (N_6768,N_1649,N_751);
xor U6769 (N_6769,N_2934,N_341);
xor U6770 (N_6770,N_3624,N_80);
or U6771 (N_6771,N_1612,N_1948);
or U6772 (N_6772,N_3657,N_3888);
and U6773 (N_6773,N_1715,N_1444);
and U6774 (N_6774,N_313,N_1795);
xnor U6775 (N_6775,N_3246,N_2865);
and U6776 (N_6776,N_2535,N_3462);
or U6777 (N_6777,N_462,N_4);
and U6778 (N_6778,N_652,N_1392);
nand U6779 (N_6779,N_2427,N_1806);
and U6780 (N_6780,N_716,N_2755);
or U6781 (N_6781,N_88,N_711);
and U6782 (N_6782,N_3833,N_2000);
xnor U6783 (N_6783,N_1750,N_3315);
and U6784 (N_6784,N_2508,N_1155);
or U6785 (N_6785,N_3934,N_1836);
xor U6786 (N_6786,N_3431,N_2867);
or U6787 (N_6787,N_1265,N_1070);
xnor U6788 (N_6788,N_2005,N_1490);
nor U6789 (N_6789,N_866,N_1190);
nand U6790 (N_6790,N_730,N_920);
nor U6791 (N_6791,N_3061,N_1929);
xnor U6792 (N_6792,N_1649,N_3107);
xnor U6793 (N_6793,N_919,N_2590);
xnor U6794 (N_6794,N_3617,N_3216);
nor U6795 (N_6795,N_3184,N_2008);
and U6796 (N_6796,N_28,N_1732);
xor U6797 (N_6797,N_271,N_1938);
xor U6798 (N_6798,N_562,N_883);
and U6799 (N_6799,N_2067,N_828);
nor U6800 (N_6800,N_1842,N_1432);
and U6801 (N_6801,N_3481,N_747);
or U6802 (N_6802,N_5,N_522);
or U6803 (N_6803,N_2587,N_2037);
xnor U6804 (N_6804,N_3591,N_3030);
nor U6805 (N_6805,N_901,N_1323);
or U6806 (N_6806,N_2868,N_852);
nor U6807 (N_6807,N_3223,N_3421);
and U6808 (N_6808,N_1350,N_1896);
nor U6809 (N_6809,N_1244,N_3929);
nand U6810 (N_6810,N_3076,N_3893);
nand U6811 (N_6811,N_709,N_2117);
and U6812 (N_6812,N_261,N_3973);
or U6813 (N_6813,N_3819,N_242);
nor U6814 (N_6814,N_3703,N_8);
nand U6815 (N_6815,N_3248,N_765);
xor U6816 (N_6816,N_1926,N_875);
nand U6817 (N_6817,N_447,N_442);
or U6818 (N_6818,N_2122,N_43);
xor U6819 (N_6819,N_1959,N_3626);
nand U6820 (N_6820,N_1926,N_2456);
nor U6821 (N_6821,N_3270,N_1016);
xor U6822 (N_6822,N_3768,N_461);
nor U6823 (N_6823,N_2622,N_1233);
nand U6824 (N_6824,N_578,N_1677);
xor U6825 (N_6825,N_957,N_688);
xor U6826 (N_6826,N_2461,N_654);
xor U6827 (N_6827,N_1287,N_988);
and U6828 (N_6828,N_2400,N_3591);
xor U6829 (N_6829,N_1874,N_1294);
nor U6830 (N_6830,N_148,N_1088);
nor U6831 (N_6831,N_3733,N_1684);
nor U6832 (N_6832,N_2343,N_1809);
nor U6833 (N_6833,N_374,N_1504);
nand U6834 (N_6834,N_2249,N_2090);
xnor U6835 (N_6835,N_3390,N_2492);
and U6836 (N_6836,N_2836,N_1799);
nand U6837 (N_6837,N_1668,N_3417);
xor U6838 (N_6838,N_381,N_2692);
nor U6839 (N_6839,N_1943,N_3602);
nor U6840 (N_6840,N_2249,N_3123);
nor U6841 (N_6841,N_2961,N_1500);
and U6842 (N_6842,N_2087,N_1579);
and U6843 (N_6843,N_1182,N_2257);
nor U6844 (N_6844,N_355,N_2331);
xnor U6845 (N_6845,N_3482,N_860);
xor U6846 (N_6846,N_1759,N_2083);
nor U6847 (N_6847,N_3671,N_1928);
nand U6848 (N_6848,N_370,N_1162);
nor U6849 (N_6849,N_1067,N_1726);
and U6850 (N_6850,N_3376,N_369);
or U6851 (N_6851,N_674,N_1794);
nand U6852 (N_6852,N_3665,N_314);
nand U6853 (N_6853,N_3369,N_2091);
nor U6854 (N_6854,N_3110,N_3038);
xor U6855 (N_6855,N_2372,N_1909);
nor U6856 (N_6856,N_736,N_37);
xnor U6857 (N_6857,N_3822,N_2010);
xor U6858 (N_6858,N_3877,N_3273);
xnor U6859 (N_6859,N_2632,N_597);
xnor U6860 (N_6860,N_2192,N_467);
and U6861 (N_6861,N_2264,N_371);
nor U6862 (N_6862,N_2489,N_2605);
nor U6863 (N_6863,N_2602,N_3435);
or U6864 (N_6864,N_394,N_686);
nor U6865 (N_6865,N_2627,N_3813);
xor U6866 (N_6866,N_3765,N_2939);
and U6867 (N_6867,N_1722,N_55);
xor U6868 (N_6868,N_421,N_249);
nand U6869 (N_6869,N_2477,N_428);
nand U6870 (N_6870,N_3524,N_538);
nor U6871 (N_6871,N_1937,N_2281);
nor U6872 (N_6872,N_643,N_2758);
nor U6873 (N_6873,N_2947,N_3863);
nand U6874 (N_6874,N_1387,N_2802);
and U6875 (N_6875,N_1274,N_2164);
nand U6876 (N_6876,N_129,N_322);
or U6877 (N_6877,N_2479,N_2187);
and U6878 (N_6878,N_398,N_1052);
nor U6879 (N_6879,N_276,N_3380);
nor U6880 (N_6880,N_3241,N_3803);
nand U6881 (N_6881,N_1464,N_2485);
xor U6882 (N_6882,N_3739,N_2326);
xor U6883 (N_6883,N_900,N_2701);
and U6884 (N_6884,N_2699,N_1492);
and U6885 (N_6885,N_923,N_2003);
nand U6886 (N_6886,N_2775,N_2813);
and U6887 (N_6887,N_1538,N_2404);
nand U6888 (N_6888,N_1534,N_1860);
xor U6889 (N_6889,N_1025,N_3939);
or U6890 (N_6890,N_2015,N_1513);
nand U6891 (N_6891,N_257,N_1201);
or U6892 (N_6892,N_2912,N_1899);
nor U6893 (N_6893,N_26,N_3575);
and U6894 (N_6894,N_2681,N_3155);
and U6895 (N_6895,N_66,N_1728);
xor U6896 (N_6896,N_2734,N_911);
nor U6897 (N_6897,N_3296,N_2225);
or U6898 (N_6898,N_2582,N_127);
nand U6899 (N_6899,N_1237,N_60);
and U6900 (N_6900,N_3367,N_1139);
nand U6901 (N_6901,N_2958,N_613);
nand U6902 (N_6902,N_2862,N_1423);
nand U6903 (N_6903,N_1829,N_1952);
nor U6904 (N_6904,N_2590,N_3679);
nor U6905 (N_6905,N_859,N_2810);
nand U6906 (N_6906,N_149,N_3499);
or U6907 (N_6907,N_1751,N_1326);
and U6908 (N_6908,N_712,N_529);
and U6909 (N_6909,N_2955,N_1490);
nor U6910 (N_6910,N_1295,N_166);
or U6911 (N_6911,N_2044,N_2116);
xnor U6912 (N_6912,N_2199,N_1346);
nor U6913 (N_6913,N_921,N_3005);
or U6914 (N_6914,N_3806,N_2456);
or U6915 (N_6915,N_1940,N_1044);
or U6916 (N_6916,N_2718,N_3889);
nand U6917 (N_6917,N_2001,N_3588);
xor U6918 (N_6918,N_3706,N_3581);
and U6919 (N_6919,N_1238,N_2320);
nand U6920 (N_6920,N_2643,N_2178);
xor U6921 (N_6921,N_1645,N_1278);
xnor U6922 (N_6922,N_2845,N_3461);
and U6923 (N_6923,N_3905,N_2274);
and U6924 (N_6924,N_1948,N_1179);
nor U6925 (N_6925,N_615,N_3021);
or U6926 (N_6926,N_1412,N_3503);
nand U6927 (N_6927,N_1717,N_1382);
xnor U6928 (N_6928,N_522,N_2016);
xor U6929 (N_6929,N_968,N_977);
xor U6930 (N_6930,N_2971,N_1877);
nor U6931 (N_6931,N_855,N_3728);
and U6932 (N_6932,N_975,N_138);
nor U6933 (N_6933,N_224,N_3379);
nor U6934 (N_6934,N_2602,N_1652);
and U6935 (N_6935,N_420,N_797);
xor U6936 (N_6936,N_251,N_2022);
or U6937 (N_6937,N_2456,N_1500);
nor U6938 (N_6938,N_2706,N_3180);
or U6939 (N_6939,N_792,N_2997);
nand U6940 (N_6940,N_2719,N_3462);
or U6941 (N_6941,N_594,N_3285);
or U6942 (N_6942,N_3886,N_479);
and U6943 (N_6943,N_1240,N_242);
or U6944 (N_6944,N_3660,N_1678);
nand U6945 (N_6945,N_2175,N_3572);
nor U6946 (N_6946,N_1411,N_3192);
nor U6947 (N_6947,N_754,N_2425);
xnor U6948 (N_6948,N_3752,N_3093);
nand U6949 (N_6949,N_2315,N_1566);
and U6950 (N_6950,N_2977,N_1295);
xnor U6951 (N_6951,N_3980,N_846);
or U6952 (N_6952,N_2856,N_1931);
or U6953 (N_6953,N_3065,N_2930);
nor U6954 (N_6954,N_1596,N_1649);
nand U6955 (N_6955,N_3175,N_2741);
nand U6956 (N_6956,N_3180,N_709);
and U6957 (N_6957,N_2688,N_1411);
xor U6958 (N_6958,N_1575,N_2219);
and U6959 (N_6959,N_2100,N_946);
and U6960 (N_6960,N_796,N_2794);
and U6961 (N_6961,N_118,N_3413);
and U6962 (N_6962,N_211,N_2299);
nor U6963 (N_6963,N_3242,N_2333);
or U6964 (N_6964,N_508,N_3966);
xnor U6965 (N_6965,N_625,N_2449);
nor U6966 (N_6966,N_1232,N_1208);
nor U6967 (N_6967,N_3628,N_814);
or U6968 (N_6968,N_1056,N_481);
and U6969 (N_6969,N_31,N_2513);
or U6970 (N_6970,N_2798,N_1986);
nand U6971 (N_6971,N_2276,N_1539);
and U6972 (N_6972,N_3560,N_3333);
nor U6973 (N_6973,N_838,N_2337);
nand U6974 (N_6974,N_3501,N_112);
xnor U6975 (N_6975,N_3164,N_2151);
nand U6976 (N_6976,N_2955,N_3298);
nand U6977 (N_6977,N_3006,N_2184);
or U6978 (N_6978,N_3975,N_895);
nand U6979 (N_6979,N_2205,N_3346);
and U6980 (N_6980,N_2614,N_394);
nand U6981 (N_6981,N_3760,N_2260);
nor U6982 (N_6982,N_2176,N_2107);
or U6983 (N_6983,N_1196,N_3533);
xor U6984 (N_6984,N_3559,N_3934);
xor U6985 (N_6985,N_178,N_2806);
and U6986 (N_6986,N_3907,N_1132);
nand U6987 (N_6987,N_3299,N_562);
xor U6988 (N_6988,N_1170,N_1883);
nand U6989 (N_6989,N_2840,N_3940);
xnor U6990 (N_6990,N_3346,N_855);
and U6991 (N_6991,N_632,N_1665);
or U6992 (N_6992,N_3901,N_3250);
or U6993 (N_6993,N_1373,N_834);
and U6994 (N_6994,N_2200,N_2380);
nor U6995 (N_6995,N_1072,N_14);
or U6996 (N_6996,N_2419,N_2540);
nand U6997 (N_6997,N_1972,N_3648);
and U6998 (N_6998,N_3692,N_1032);
nor U6999 (N_6999,N_3242,N_1845);
nand U7000 (N_7000,N_78,N_3782);
and U7001 (N_7001,N_3981,N_1523);
or U7002 (N_7002,N_3014,N_3184);
or U7003 (N_7003,N_317,N_3278);
and U7004 (N_7004,N_2280,N_1338);
nand U7005 (N_7005,N_2585,N_2614);
or U7006 (N_7006,N_477,N_2765);
nor U7007 (N_7007,N_994,N_1452);
nand U7008 (N_7008,N_3609,N_2452);
or U7009 (N_7009,N_665,N_1661);
and U7010 (N_7010,N_3920,N_1890);
xor U7011 (N_7011,N_3409,N_2579);
or U7012 (N_7012,N_105,N_146);
xor U7013 (N_7013,N_2384,N_627);
nor U7014 (N_7014,N_2647,N_421);
nor U7015 (N_7015,N_2002,N_2841);
nand U7016 (N_7016,N_1136,N_2060);
and U7017 (N_7017,N_3640,N_153);
or U7018 (N_7018,N_456,N_795);
and U7019 (N_7019,N_1301,N_1888);
nor U7020 (N_7020,N_55,N_1301);
nand U7021 (N_7021,N_2157,N_2090);
nor U7022 (N_7022,N_2724,N_1124);
nand U7023 (N_7023,N_1475,N_2288);
xnor U7024 (N_7024,N_476,N_216);
nand U7025 (N_7025,N_3012,N_1180);
nand U7026 (N_7026,N_821,N_3808);
and U7027 (N_7027,N_2027,N_364);
nor U7028 (N_7028,N_1547,N_1724);
nand U7029 (N_7029,N_2187,N_1397);
or U7030 (N_7030,N_3703,N_3679);
and U7031 (N_7031,N_2783,N_999);
nand U7032 (N_7032,N_2192,N_1833);
or U7033 (N_7033,N_1025,N_861);
or U7034 (N_7034,N_1699,N_1824);
xnor U7035 (N_7035,N_1189,N_3079);
nand U7036 (N_7036,N_1193,N_3420);
or U7037 (N_7037,N_3616,N_899);
and U7038 (N_7038,N_2423,N_3753);
xnor U7039 (N_7039,N_193,N_2168);
nor U7040 (N_7040,N_2957,N_2839);
nand U7041 (N_7041,N_3679,N_865);
and U7042 (N_7042,N_3728,N_112);
xnor U7043 (N_7043,N_495,N_2889);
nor U7044 (N_7044,N_1613,N_1561);
or U7045 (N_7045,N_3650,N_1164);
and U7046 (N_7046,N_2953,N_521);
or U7047 (N_7047,N_3856,N_119);
or U7048 (N_7048,N_2310,N_310);
and U7049 (N_7049,N_3777,N_2120);
nand U7050 (N_7050,N_703,N_1109);
nand U7051 (N_7051,N_2799,N_2513);
nand U7052 (N_7052,N_1503,N_1743);
and U7053 (N_7053,N_83,N_3809);
xor U7054 (N_7054,N_1497,N_313);
nand U7055 (N_7055,N_296,N_1803);
xnor U7056 (N_7056,N_717,N_2497);
nor U7057 (N_7057,N_1012,N_2985);
or U7058 (N_7058,N_1629,N_2330);
and U7059 (N_7059,N_2871,N_743);
nor U7060 (N_7060,N_3347,N_202);
nand U7061 (N_7061,N_2364,N_689);
and U7062 (N_7062,N_1613,N_3099);
xor U7063 (N_7063,N_1021,N_279);
nand U7064 (N_7064,N_3745,N_2022);
or U7065 (N_7065,N_1318,N_1440);
xnor U7066 (N_7066,N_2209,N_3254);
nand U7067 (N_7067,N_87,N_1580);
nor U7068 (N_7068,N_3885,N_3229);
xor U7069 (N_7069,N_2826,N_438);
nor U7070 (N_7070,N_308,N_1188);
nand U7071 (N_7071,N_1813,N_2077);
nor U7072 (N_7072,N_3634,N_3476);
or U7073 (N_7073,N_1876,N_579);
xnor U7074 (N_7074,N_199,N_2048);
nor U7075 (N_7075,N_3693,N_2628);
nand U7076 (N_7076,N_2361,N_2688);
xnor U7077 (N_7077,N_368,N_837);
nand U7078 (N_7078,N_1143,N_96);
xor U7079 (N_7079,N_815,N_823);
xnor U7080 (N_7080,N_1569,N_2581);
or U7081 (N_7081,N_3696,N_1518);
and U7082 (N_7082,N_987,N_2355);
nor U7083 (N_7083,N_3789,N_3677);
or U7084 (N_7084,N_663,N_3737);
nor U7085 (N_7085,N_1434,N_20);
nand U7086 (N_7086,N_2799,N_564);
xor U7087 (N_7087,N_2386,N_2039);
nand U7088 (N_7088,N_3214,N_3037);
xor U7089 (N_7089,N_2193,N_114);
xnor U7090 (N_7090,N_1699,N_667);
nand U7091 (N_7091,N_1796,N_202);
nor U7092 (N_7092,N_1152,N_3246);
nand U7093 (N_7093,N_3980,N_1597);
nor U7094 (N_7094,N_3262,N_2792);
or U7095 (N_7095,N_936,N_831);
xor U7096 (N_7096,N_659,N_3654);
and U7097 (N_7097,N_924,N_2347);
and U7098 (N_7098,N_289,N_1395);
xor U7099 (N_7099,N_180,N_884);
nor U7100 (N_7100,N_2508,N_3794);
xor U7101 (N_7101,N_1003,N_2890);
and U7102 (N_7102,N_1999,N_573);
nand U7103 (N_7103,N_1680,N_3727);
and U7104 (N_7104,N_3195,N_271);
or U7105 (N_7105,N_1707,N_2606);
nand U7106 (N_7106,N_1282,N_3342);
nor U7107 (N_7107,N_1747,N_764);
nor U7108 (N_7108,N_742,N_2268);
nand U7109 (N_7109,N_796,N_2522);
nor U7110 (N_7110,N_1671,N_2853);
or U7111 (N_7111,N_3212,N_246);
xnor U7112 (N_7112,N_60,N_1142);
or U7113 (N_7113,N_2712,N_2319);
and U7114 (N_7114,N_545,N_2975);
nand U7115 (N_7115,N_3688,N_207);
nor U7116 (N_7116,N_2534,N_25);
nor U7117 (N_7117,N_502,N_3461);
xor U7118 (N_7118,N_1653,N_815);
xnor U7119 (N_7119,N_2538,N_304);
nand U7120 (N_7120,N_3497,N_3534);
or U7121 (N_7121,N_524,N_2682);
nor U7122 (N_7122,N_219,N_1782);
and U7123 (N_7123,N_446,N_2302);
xor U7124 (N_7124,N_768,N_2935);
or U7125 (N_7125,N_3263,N_2983);
xnor U7126 (N_7126,N_1715,N_1437);
xor U7127 (N_7127,N_2962,N_3213);
nor U7128 (N_7128,N_1513,N_707);
xnor U7129 (N_7129,N_1264,N_1041);
and U7130 (N_7130,N_588,N_2039);
nand U7131 (N_7131,N_891,N_2270);
nor U7132 (N_7132,N_3433,N_1683);
nor U7133 (N_7133,N_1624,N_1173);
nor U7134 (N_7134,N_1441,N_851);
nand U7135 (N_7135,N_159,N_3609);
nand U7136 (N_7136,N_115,N_492);
xor U7137 (N_7137,N_1401,N_3822);
xor U7138 (N_7138,N_2963,N_3703);
xor U7139 (N_7139,N_1025,N_1172);
xor U7140 (N_7140,N_2999,N_1897);
and U7141 (N_7141,N_1362,N_3656);
nor U7142 (N_7142,N_3446,N_2081);
nand U7143 (N_7143,N_891,N_2461);
and U7144 (N_7144,N_55,N_722);
or U7145 (N_7145,N_3914,N_2543);
and U7146 (N_7146,N_2751,N_1162);
nor U7147 (N_7147,N_3056,N_3624);
or U7148 (N_7148,N_1600,N_2616);
nor U7149 (N_7149,N_503,N_197);
and U7150 (N_7150,N_3876,N_1460);
or U7151 (N_7151,N_1400,N_3506);
and U7152 (N_7152,N_2637,N_2885);
nor U7153 (N_7153,N_1092,N_1639);
or U7154 (N_7154,N_359,N_1063);
nor U7155 (N_7155,N_1935,N_3267);
xor U7156 (N_7156,N_3672,N_1286);
nor U7157 (N_7157,N_1129,N_2815);
and U7158 (N_7158,N_342,N_3426);
and U7159 (N_7159,N_2675,N_3283);
xnor U7160 (N_7160,N_3531,N_1436);
nand U7161 (N_7161,N_3294,N_824);
xnor U7162 (N_7162,N_3583,N_2968);
nand U7163 (N_7163,N_117,N_2121);
and U7164 (N_7164,N_1233,N_1545);
xor U7165 (N_7165,N_2873,N_1422);
and U7166 (N_7166,N_471,N_2681);
xor U7167 (N_7167,N_1396,N_3648);
xor U7168 (N_7168,N_3563,N_1233);
xnor U7169 (N_7169,N_2279,N_2491);
xnor U7170 (N_7170,N_811,N_3202);
xor U7171 (N_7171,N_3201,N_2152);
xor U7172 (N_7172,N_2972,N_3399);
xnor U7173 (N_7173,N_3800,N_2143);
and U7174 (N_7174,N_3633,N_1126);
nand U7175 (N_7175,N_197,N_3559);
xnor U7176 (N_7176,N_2793,N_975);
and U7177 (N_7177,N_3332,N_1130);
nor U7178 (N_7178,N_3168,N_1447);
or U7179 (N_7179,N_508,N_1184);
or U7180 (N_7180,N_1020,N_1412);
or U7181 (N_7181,N_698,N_1612);
and U7182 (N_7182,N_3840,N_1516);
nor U7183 (N_7183,N_591,N_1688);
xor U7184 (N_7184,N_3325,N_2382);
and U7185 (N_7185,N_2384,N_2574);
xor U7186 (N_7186,N_2495,N_2058);
xor U7187 (N_7187,N_1740,N_2257);
xnor U7188 (N_7188,N_263,N_154);
or U7189 (N_7189,N_3849,N_2737);
nor U7190 (N_7190,N_1157,N_3032);
and U7191 (N_7191,N_2947,N_2988);
xor U7192 (N_7192,N_1424,N_982);
xnor U7193 (N_7193,N_1379,N_3113);
nand U7194 (N_7194,N_2134,N_2429);
and U7195 (N_7195,N_3447,N_1591);
or U7196 (N_7196,N_2145,N_3949);
nand U7197 (N_7197,N_3,N_888);
nand U7198 (N_7198,N_2494,N_207);
xnor U7199 (N_7199,N_1040,N_2698);
xnor U7200 (N_7200,N_3310,N_3342);
xnor U7201 (N_7201,N_3429,N_2334);
xor U7202 (N_7202,N_623,N_415);
xor U7203 (N_7203,N_2511,N_1403);
and U7204 (N_7204,N_2133,N_3717);
and U7205 (N_7205,N_744,N_1334);
nor U7206 (N_7206,N_192,N_929);
or U7207 (N_7207,N_2128,N_3503);
xor U7208 (N_7208,N_1782,N_696);
and U7209 (N_7209,N_1843,N_1126);
nor U7210 (N_7210,N_3731,N_370);
nand U7211 (N_7211,N_2900,N_220);
nor U7212 (N_7212,N_3841,N_3366);
and U7213 (N_7213,N_3630,N_1054);
and U7214 (N_7214,N_3980,N_2146);
nand U7215 (N_7215,N_2488,N_91);
or U7216 (N_7216,N_3519,N_2012);
or U7217 (N_7217,N_2796,N_2703);
and U7218 (N_7218,N_1481,N_769);
nand U7219 (N_7219,N_231,N_3156);
nand U7220 (N_7220,N_517,N_148);
xor U7221 (N_7221,N_3292,N_1115);
nor U7222 (N_7222,N_132,N_947);
nor U7223 (N_7223,N_1258,N_3289);
nand U7224 (N_7224,N_468,N_190);
nand U7225 (N_7225,N_3514,N_334);
xor U7226 (N_7226,N_3055,N_3036);
and U7227 (N_7227,N_2696,N_3312);
nand U7228 (N_7228,N_1750,N_2563);
nand U7229 (N_7229,N_545,N_1095);
xor U7230 (N_7230,N_653,N_3394);
or U7231 (N_7231,N_1186,N_654);
and U7232 (N_7232,N_1315,N_1803);
nor U7233 (N_7233,N_363,N_1926);
or U7234 (N_7234,N_3022,N_62);
nand U7235 (N_7235,N_2561,N_731);
xor U7236 (N_7236,N_3751,N_1447);
and U7237 (N_7237,N_1945,N_1161);
or U7238 (N_7238,N_3040,N_547);
and U7239 (N_7239,N_3183,N_2715);
xor U7240 (N_7240,N_2322,N_839);
nand U7241 (N_7241,N_3049,N_1136);
and U7242 (N_7242,N_87,N_948);
and U7243 (N_7243,N_2278,N_1683);
xor U7244 (N_7244,N_3212,N_477);
nor U7245 (N_7245,N_1170,N_1496);
xnor U7246 (N_7246,N_2631,N_1886);
nand U7247 (N_7247,N_927,N_664);
or U7248 (N_7248,N_2558,N_3165);
xnor U7249 (N_7249,N_3895,N_1075);
xor U7250 (N_7250,N_2618,N_97);
nand U7251 (N_7251,N_3097,N_3739);
xnor U7252 (N_7252,N_2259,N_2973);
nand U7253 (N_7253,N_810,N_2738);
nor U7254 (N_7254,N_1417,N_1701);
and U7255 (N_7255,N_3840,N_1001);
or U7256 (N_7256,N_2293,N_764);
nor U7257 (N_7257,N_2717,N_1361);
or U7258 (N_7258,N_2214,N_868);
or U7259 (N_7259,N_3632,N_559);
xor U7260 (N_7260,N_1509,N_2761);
and U7261 (N_7261,N_3295,N_3615);
nand U7262 (N_7262,N_2433,N_2393);
nor U7263 (N_7263,N_190,N_1344);
nor U7264 (N_7264,N_1178,N_1535);
xor U7265 (N_7265,N_540,N_732);
or U7266 (N_7266,N_2742,N_3160);
nand U7267 (N_7267,N_325,N_3511);
nand U7268 (N_7268,N_3403,N_2853);
nor U7269 (N_7269,N_468,N_1144);
xnor U7270 (N_7270,N_820,N_1262);
xor U7271 (N_7271,N_3945,N_818);
or U7272 (N_7272,N_1624,N_609);
nor U7273 (N_7273,N_105,N_3232);
nor U7274 (N_7274,N_3185,N_1185);
xor U7275 (N_7275,N_3711,N_3782);
nor U7276 (N_7276,N_443,N_1696);
nor U7277 (N_7277,N_2295,N_1242);
or U7278 (N_7278,N_2749,N_2750);
nor U7279 (N_7279,N_2184,N_338);
nor U7280 (N_7280,N_200,N_2700);
and U7281 (N_7281,N_2964,N_3224);
or U7282 (N_7282,N_1876,N_3620);
nand U7283 (N_7283,N_3883,N_3216);
nand U7284 (N_7284,N_3079,N_2314);
nand U7285 (N_7285,N_642,N_1056);
xor U7286 (N_7286,N_1616,N_1444);
nor U7287 (N_7287,N_2058,N_877);
xor U7288 (N_7288,N_1582,N_3596);
nor U7289 (N_7289,N_742,N_2822);
and U7290 (N_7290,N_3304,N_2632);
and U7291 (N_7291,N_1957,N_2205);
or U7292 (N_7292,N_3879,N_654);
nand U7293 (N_7293,N_362,N_3227);
xnor U7294 (N_7294,N_3763,N_473);
nand U7295 (N_7295,N_214,N_1381);
or U7296 (N_7296,N_733,N_293);
nor U7297 (N_7297,N_2695,N_766);
or U7298 (N_7298,N_2856,N_3803);
nor U7299 (N_7299,N_2205,N_690);
nand U7300 (N_7300,N_108,N_1606);
nand U7301 (N_7301,N_2020,N_29);
nand U7302 (N_7302,N_755,N_209);
nand U7303 (N_7303,N_197,N_1503);
xnor U7304 (N_7304,N_3006,N_1585);
xnor U7305 (N_7305,N_1986,N_3668);
nor U7306 (N_7306,N_229,N_3875);
nor U7307 (N_7307,N_3787,N_2185);
or U7308 (N_7308,N_250,N_2504);
nand U7309 (N_7309,N_564,N_292);
xor U7310 (N_7310,N_3487,N_1465);
xnor U7311 (N_7311,N_1147,N_1513);
or U7312 (N_7312,N_2096,N_831);
xnor U7313 (N_7313,N_180,N_2530);
xnor U7314 (N_7314,N_574,N_1983);
and U7315 (N_7315,N_2354,N_3586);
nor U7316 (N_7316,N_2018,N_2135);
and U7317 (N_7317,N_150,N_1719);
xnor U7318 (N_7318,N_2858,N_3791);
xnor U7319 (N_7319,N_1401,N_2340);
or U7320 (N_7320,N_865,N_2282);
and U7321 (N_7321,N_1857,N_802);
nor U7322 (N_7322,N_2402,N_3788);
nor U7323 (N_7323,N_3576,N_3130);
xor U7324 (N_7324,N_2930,N_2070);
nor U7325 (N_7325,N_2215,N_2218);
nand U7326 (N_7326,N_2032,N_2189);
nand U7327 (N_7327,N_2214,N_610);
or U7328 (N_7328,N_2841,N_1900);
nor U7329 (N_7329,N_3284,N_1474);
and U7330 (N_7330,N_3911,N_2996);
xor U7331 (N_7331,N_3049,N_1147);
or U7332 (N_7332,N_2201,N_2408);
nor U7333 (N_7333,N_1784,N_782);
nand U7334 (N_7334,N_3119,N_3234);
nand U7335 (N_7335,N_1036,N_2472);
nand U7336 (N_7336,N_1214,N_3781);
and U7337 (N_7337,N_2033,N_1994);
nor U7338 (N_7338,N_2304,N_3670);
and U7339 (N_7339,N_2580,N_869);
nor U7340 (N_7340,N_988,N_3317);
nand U7341 (N_7341,N_2526,N_1213);
or U7342 (N_7342,N_1749,N_204);
or U7343 (N_7343,N_619,N_2606);
or U7344 (N_7344,N_2587,N_2310);
xnor U7345 (N_7345,N_3149,N_2737);
xnor U7346 (N_7346,N_2650,N_3931);
xor U7347 (N_7347,N_1916,N_2877);
or U7348 (N_7348,N_3914,N_1882);
or U7349 (N_7349,N_1648,N_3326);
and U7350 (N_7350,N_1345,N_3539);
nand U7351 (N_7351,N_9,N_2713);
nand U7352 (N_7352,N_2114,N_3879);
nor U7353 (N_7353,N_2627,N_543);
nand U7354 (N_7354,N_984,N_2710);
nand U7355 (N_7355,N_2512,N_3109);
xnor U7356 (N_7356,N_1670,N_2023);
or U7357 (N_7357,N_1623,N_3354);
and U7358 (N_7358,N_3393,N_3645);
nand U7359 (N_7359,N_24,N_1978);
and U7360 (N_7360,N_1950,N_1964);
nand U7361 (N_7361,N_1661,N_3804);
nand U7362 (N_7362,N_3692,N_724);
nor U7363 (N_7363,N_3889,N_2559);
or U7364 (N_7364,N_2763,N_3337);
and U7365 (N_7365,N_591,N_1566);
nor U7366 (N_7366,N_3838,N_3778);
nand U7367 (N_7367,N_3709,N_2715);
or U7368 (N_7368,N_3452,N_3225);
or U7369 (N_7369,N_3755,N_3234);
xor U7370 (N_7370,N_3155,N_2262);
and U7371 (N_7371,N_471,N_500);
nor U7372 (N_7372,N_2577,N_3759);
or U7373 (N_7373,N_736,N_151);
nand U7374 (N_7374,N_3502,N_3944);
nand U7375 (N_7375,N_1665,N_134);
nand U7376 (N_7376,N_3032,N_2778);
nand U7377 (N_7377,N_635,N_1073);
nand U7378 (N_7378,N_412,N_2630);
and U7379 (N_7379,N_3999,N_3346);
nand U7380 (N_7380,N_1789,N_3022);
xnor U7381 (N_7381,N_2772,N_3629);
or U7382 (N_7382,N_3104,N_1744);
nand U7383 (N_7383,N_3891,N_3444);
nand U7384 (N_7384,N_366,N_3573);
xnor U7385 (N_7385,N_958,N_2506);
nand U7386 (N_7386,N_1138,N_953);
and U7387 (N_7387,N_2222,N_2155);
nand U7388 (N_7388,N_1444,N_3707);
nor U7389 (N_7389,N_3851,N_3777);
and U7390 (N_7390,N_2393,N_1228);
or U7391 (N_7391,N_702,N_3474);
nor U7392 (N_7392,N_2244,N_3956);
nor U7393 (N_7393,N_1,N_453);
and U7394 (N_7394,N_119,N_1970);
xor U7395 (N_7395,N_469,N_787);
nand U7396 (N_7396,N_1561,N_15);
or U7397 (N_7397,N_1841,N_3112);
and U7398 (N_7398,N_936,N_1317);
xnor U7399 (N_7399,N_179,N_2891);
xor U7400 (N_7400,N_2095,N_1648);
nor U7401 (N_7401,N_14,N_1713);
and U7402 (N_7402,N_1847,N_2038);
nand U7403 (N_7403,N_1491,N_450);
and U7404 (N_7404,N_2199,N_1153);
or U7405 (N_7405,N_2309,N_1466);
nor U7406 (N_7406,N_1756,N_2330);
nor U7407 (N_7407,N_107,N_3716);
xnor U7408 (N_7408,N_3077,N_145);
or U7409 (N_7409,N_2350,N_3122);
nand U7410 (N_7410,N_2699,N_2212);
nor U7411 (N_7411,N_1885,N_2255);
nor U7412 (N_7412,N_2715,N_1338);
xor U7413 (N_7413,N_2188,N_2870);
nand U7414 (N_7414,N_1890,N_1233);
nor U7415 (N_7415,N_1460,N_2469);
xnor U7416 (N_7416,N_1110,N_3893);
nor U7417 (N_7417,N_3013,N_2554);
xnor U7418 (N_7418,N_1896,N_1831);
nor U7419 (N_7419,N_856,N_1707);
and U7420 (N_7420,N_1074,N_1331);
nor U7421 (N_7421,N_189,N_1554);
or U7422 (N_7422,N_1041,N_1407);
nor U7423 (N_7423,N_944,N_498);
nor U7424 (N_7424,N_900,N_3403);
and U7425 (N_7425,N_1492,N_2127);
nand U7426 (N_7426,N_3841,N_3276);
and U7427 (N_7427,N_194,N_2586);
or U7428 (N_7428,N_2708,N_1001);
nand U7429 (N_7429,N_2788,N_2239);
xnor U7430 (N_7430,N_825,N_3645);
nor U7431 (N_7431,N_2994,N_3658);
or U7432 (N_7432,N_1185,N_1329);
nor U7433 (N_7433,N_2206,N_1280);
xnor U7434 (N_7434,N_3659,N_3771);
nor U7435 (N_7435,N_3027,N_770);
xor U7436 (N_7436,N_592,N_3020);
or U7437 (N_7437,N_1244,N_642);
or U7438 (N_7438,N_2567,N_3137);
or U7439 (N_7439,N_3473,N_2264);
and U7440 (N_7440,N_3610,N_3152);
nor U7441 (N_7441,N_230,N_458);
or U7442 (N_7442,N_875,N_2951);
or U7443 (N_7443,N_376,N_1821);
xnor U7444 (N_7444,N_2670,N_1088);
or U7445 (N_7445,N_2361,N_1190);
xnor U7446 (N_7446,N_271,N_740);
and U7447 (N_7447,N_915,N_355);
xnor U7448 (N_7448,N_442,N_741);
and U7449 (N_7449,N_1974,N_277);
or U7450 (N_7450,N_2718,N_2903);
or U7451 (N_7451,N_3817,N_3185);
nor U7452 (N_7452,N_1098,N_3386);
nor U7453 (N_7453,N_2218,N_1444);
nor U7454 (N_7454,N_2501,N_1263);
nor U7455 (N_7455,N_3660,N_1547);
xor U7456 (N_7456,N_3436,N_2426);
or U7457 (N_7457,N_1219,N_2985);
or U7458 (N_7458,N_684,N_1529);
xor U7459 (N_7459,N_687,N_2782);
or U7460 (N_7460,N_3299,N_3460);
and U7461 (N_7461,N_3798,N_924);
xnor U7462 (N_7462,N_3940,N_705);
and U7463 (N_7463,N_1468,N_3717);
and U7464 (N_7464,N_270,N_3928);
nor U7465 (N_7465,N_152,N_1687);
and U7466 (N_7466,N_3835,N_3063);
nand U7467 (N_7467,N_3099,N_3320);
xor U7468 (N_7468,N_1705,N_323);
or U7469 (N_7469,N_419,N_3029);
or U7470 (N_7470,N_2949,N_2739);
and U7471 (N_7471,N_195,N_244);
nor U7472 (N_7472,N_2283,N_434);
xnor U7473 (N_7473,N_2398,N_3890);
and U7474 (N_7474,N_2289,N_2551);
and U7475 (N_7475,N_1405,N_2317);
or U7476 (N_7476,N_2355,N_3793);
nor U7477 (N_7477,N_2121,N_2022);
and U7478 (N_7478,N_603,N_3051);
xor U7479 (N_7479,N_3519,N_2630);
xor U7480 (N_7480,N_1129,N_3408);
xnor U7481 (N_7481,N_2910,N_3182);
xor U7482 (N_7482,N_3759,N_1206);
nand U7483 (N_7483,N_92,N_2092);
xnor U7484 (N_7484,N_297,N_65);
and U7485 (N_7485,N_185,N_1292);
or U7486 (N_7486,N_2913,N_3723);
xnor U7487 (N_7487,N_140,N_3163);
or U7488 (N_7488,N_183,N_2121);
xor U7489 (N_7489,N_344,N_2999);
nand U7490 (N_7490,N_3414,N_810);
xnor U7491 (N_7491,N_148,N_1919);
xnor U7492 (N_7492,N_2197,N_3983);
xnor U7493 (N_7493,N_3466,N_2467);
or U7494 (N_7494,N_222,N_2652);
nand U7495 (N_7495,N_1216,N_3713);
xnor U7496 (N_7496,N_1911,N_1590);
nor U7497 (N_7497,N_3638,N_2272);
or U7498 (N_7498,N_3774,N_1740);
or U7499 (N_7499,N_3423,N_2066);
xnor U7500 (N_7500,N_17,N_968);
nor U7501 (N_7501,N_2708,N_2722);
and U7502 (N_7502,N_435,N_3843);
xnor U7503 (N_7503,N_3376,N_648);
and U7504 (N_7504,N_639,N_948);
xnor U7505 (N_7505,N_1172,N_2707);
nor U7506 (N_7506,N_2006,N_2338);
nand U7507 (N_7507,N_291,N_1761);
nor U7508 (N_7508,N_3574,N_2457);
and U7509 (N_7509,N_661,N_3316);
xor U7510 (N_7510,N_2734,N_1914);
nand U7511 (N_7511,N_1824,N_6);
or U7512 (N_7512,N_513,N_938);
nor U7513 (N_7513,N_3482,N_2069);
xnor U7514 (N_7514,N_3226,N_3039);
nor U7515 (N_7515,N_2663,N_20);
nor U7516 (N_7516,N_3995,N_401);
nand U7517 (N_7517,N_1852,N_308);
nand U7518 (N_7518,N_613,N_3236);
and U7519 (N_7519,N_2616,N_1187);
nor U7520 (N_7520,N_2049,N_836);
nand U7521 (N_7521,N_1861,N_3741);
xor U7522 (N_7522,N_1562,N_1328);
nor U7523 (N_7523,N_2173,N_3289);
nand U7524 (N_7524,N_1153,N_3824);
xor U7525 (N_7525,N_1016,N_998);
xor U7526 (N_7526,N_499,N_378);
nand U7527 (N_7527,N_3225,N_2181);
and U7528 (N_7528,N_196,N_543);
nand U7529 (N_7529,N_920,N_3423);
nor U7530 (N_7530,N_2604,N_3673);
or U7531 (N_7531,N_3337,N_1636);
and U7532 (N_7532,N_2151,N_1858);
nand U7533 (N_7533,N_661,N_367);
xnor U7534 (N_7534,N_1418,N_3262);
nand U7535 (N_7535,N_3479,N_2563);
nand U7536 (N_7536,N_610,N_3437);
nand U7537 (N_7537,N_1528,N_2159);
and U7538 (N_7538,N_2178,N_582);
xnor U7539 (N_7539,N_3430,N_2617);
nand U7540 (N_7540,N_3846,N_1239);
or U7541 (N_7541,N_276,N_2382);
or U7542 (N_7542,N_3558,N_48);
or U7543 (N_7543,N_162,N_904);
nor U7544 (N_7544,N_1109,N_3052);
or U7545 (N_7545,N_3972,N_967);
nand U7546 (N_7546,N_2098,N_1355);
or U7547 (N_7547,N_357,N_3084);
nor U7548 (N_7548,N_1552,N_3586);
and U7549 (N_7549,N_1629,N_2859);
or U7550 (N_7550,N_3983,N_3825);
xor U7551 (N_7551,N_3284,N_700);
nand U7552 (N_7552,N_2297,N_3498);
or U7553 (N_7553,N_3488,N_825);
or U7554 (N_7554,N_156,N_2061);
nand U7555 (N_7555,N_3661,N_2507);
nor U7556 (N_7556,N_2203,N_1576);
and U7557 (N_7557,N_773,N_438);
or U7558 (N_7558,N_1277,N_3020);
nor U7559 (N_7559,N_2864,N_698);
xor U7560 (N_7560,N_3981,N_2951);
xnor U7561 (N_7561,N_3108,N_686);
nor U7562 (N_7562,N_319,N_276);
nor U7563 (N_7563,N_3864,N_2405);
nor U7564 (N_7564,N_1762,N_2596);
nor U7565 (N_7565,N_3205,N_678);
and U7566 (N_7566,N_967,N_2415);
or U7567 (N_7567,N_3286,N_1474);
or U7568 (N_7568,N_2857,N_1898);
and U7569 (N_7569,N_1244,N_3958);
nand U7570 (N_7570,N_2194,N_3265);
nor U7571 (N_7571,N_716,N_991);
nand U7572 (N_7572,N_2075,N_3785);
or U7573 (N_7573,N_3440,N_1221);
xnor U7574 (N_7574,N_733,N_402);
nand U7575 (N_7575,N_2369,N_1396);
nand U7576 (N_7576,N_1215,N_2306);
xor U7577 (N_7577,N_3638,N_885);
nor U7578 (N_7578,N_2100,N_2712);
nor U7579 (N_7579,N_3335,N_3872);
nand U7580 (N_7580,N_1308,N_905);
and U7581 (N_7581,N_3614,N_2067);
and U7582 (N_7582,N_2942,N_2866);
nand U7583 (N_7583,N_3441,N_1865);
or U7584 (N_7584,N_190,N_820);
or U7585 (N_7585,N_1197,N_3276);
xnor U7586 (N_7586,N_1033,N_1686);
xnor U7587 (N_7587,N_1620,N_2163);
nor U7588 (N_7588,N_1046,N_3737);
nand U7589 (N_7589,N_57,N_3980);
nand U7590 (N_7590,N_2701,N_3651);
and U7591 (N_7591,N_2377,N_3948);
nand U7592 (N_7592,N_3507,N_3907);
or U7593 (N_7593,N_3867,N_3441);
xor U7594 (N_7594,N_1651,N_2175);
or U7595 (N_7595,N_2074,N_3424);
xor U7596 (N_7596,N_1445,N_1340);
or U7597 (N_7597,N_1985,N_164);
xnor U7598 (N_7598,N_1279,N_1157);
and U7599 (N_7599,N_864,N_625);
nor U7600 (N_7600,N_3565,N_1816);
or U7601 (N_7601,N_3959,N_1651);
nor U7602 (N_7602,N_1225,N_1105);
nor U7603 (N_7603,N_2446,N_303);
nand U7604 (N_7604,N_1785,N_1796);
or U7605 (N_7605,N_762,N_3623);
or U7606 (N_7606,N_3550,N_25);
and U7607 (N_7607,N_2693,N_3440);
or U7608 (N_7608,N_817,N_2781);
or U7609 (N_7609,N_825,N_3387);
nand U7610 (N_7610,N_64,N_1432);
and U7611 (N_7611,N_87,N_765);
nand U7612 (N_7612,N_2780,N_2799);
and U7613 (N_7613,N_3570,N_2670);
nand U7614 (N_7614,N_1656,N_2719);
xor U7615 (N_7615,N_883,N_2070);
or U7616 (N_7616,N_1385,N_736);
or U7617 (N_7617,N_1632,N_3255);
nand U7618 (N_7618,N_3705,N_1130);
and U7619 (N_7619,N_3421,N_2684);
and U7620 (N_7620,N_1882,N_1989);
nand U7621 (N_7621,N_3135,N_1328);
nor U7622 (N_7622,N_3276,N_2915);
xnor U7623 (N_7623,N_1508,N_246);
xor U7624 (N_7624,N_19,N_1874);
nor U7625 (N_7625,N_2171,N_3961);
xnor U7626 (N_7626,N_1779,N_3877);
nand U7627 (N_7627,N_3745,N_1648);
xnor U7628 (N_7628,N_1495,N_768);
and U7629 (N_7629,N_343,N_3982);
nor U7630 (N_7630,N_3577,N_227);
xnor U7631 (N_7631,N_3149,N_2577);
nand U7632 (N_7632,N_3707,N_3828);
and U7633 (N_7633,N_1787,N_3609);
and U7634 (N_7634,N_3310,N_1616);
or U7635 (N_7635,N_1245,N_2239);
or U7636 (N_7636,N_413,N_30);
xor U7637 (N_7637,N_545,N_3199);
nor U7638 (N_7638,N_3169,N_135);
xnor U7639 (N_7639,N_784,N_2213);
and U7640 (N_7640,N_280,N_1015);
xnor U7641 (N_7641,N_1987,N_3655);
and U7642 (N_7642,N_1337,N_3544);
nand U7643 (N_7643,N_3999,N_1136);
and U7644 (N_7644,N_2344,N_3165);
nor U7645 (N_7645,N_2431,N_2643);
xnor U7646 (N_7646,N_1605,N_2163);
nand U7647 (N_7647,N_222,N_1918);
or U7648 (N_7648,N_2197,N_3303);
xor U7649 (N_7649,N_2999,N_2877);
xnor U7650 (N_7650,N_3099,N_2202);
nor U7651 (N_7651,N_1671,N_2610);
nor U7652 (N_7652,N_3322,N_1593);
nor U7653 (N_7653,N_3336,N_3497);
or U7654 (N_7654,N_723,N_3177);
or U7655 (N_7655,N_1331,N_3296);
nand U7656 (N_7656,N_3178,N_3831);
and U7657 (N_7657,N_795,N_2057);
nor U7658 (N_7658,N_695,N_1592);
or U7659 (N_7659,N_3079,N_2904);
nand U7660 (N_7660,N_1930,N_1909);
nand U7661 (N_7661,N_2582,N_1007);
or U7662 (N_7662,N_664,N_1416);
xor U7663 (N_7663,N_707,N_3075);
nor U7664 (N_7664,N_320,N_3510);
nand U7665 (N_7665,N_2451,N_42);
or U7666 (N_7666,N_2206,N_3139);
nand U7667 (N_7667,N_368,N_3671);
xnor U7668 (N_7668,N_411,N_2478);
nor U7669 (N_7669,N_3451,N_377);
and U7670 (N_7670,N_1399,N_1621);
xnor U7671 (N_7671,N_775,N_600);
and U7672 (N_7672,N_2431,N_1469);
xnor U7673 (N_7673,N_465,N_2855);
or U7674 (N_7674,N_3316,N_441);
xor U7675 (N_7675,N_91,N_3732);
xnor U7676 (N_7676,N_1001,N_933);
xor U7677 (N_7677,N_3494,N_2740);
nand U7678 (N_7678,N_1483,N_3112);
or U7679 (N_7679,N_1966,N_3638);
xnor U7680 (N_7680,N_3594,N_665);
nand U7681 (N_7681,N_3448,N_2057);
nand U7682 (N_7682,N_2578,N_1773);
or U7683 (N_7683,N_660,N_2159);
nor U7684 (N_7684,N_1609,N_3051);
xor U7685 (N_7685,N_942,N_937);
nand U7686 (N_7686,N_223,N_2542);
nand U7687 (N_7687,N_184,N_1247);
and U7688 (N_7688,N_3027,N_3151);
and U7689 (N_7689,N_2265,N_1568);
nor U7690 (N_7690,N_2654,N_1292);
xnor U7691 (N_7691,N_1440,N_596);
xor U7692 (N_7692,N_2014,N_1545);
xnor U7693 (N_7693,N_3778,N_3240);
nor U7694 (N_7694,N_2112,N_840);
or U7695 (N_7695,N_3655,N_2052);
and U7696 (N_7696,N_17,N_1743);
or U7697 (N_7697,N_1837,N_1068);
xnor U7698 (N_7698,N_957,N_1345);
nor U7699 (N_7699,N_1769,N_2873);
and U7700 (N_7700,N_980,N_3057);
and U7701 (N_7701,N_165,N_3036);
nor U7702 (N_7702,N_272,N_1797);
or U7703 (N_7703,N_1081,N_2546);
xor U7704 (N_7704,N_1792,N_2468);
nand U7705 (N_7705,N_2466,N_1235);
xnor U7706 (N_7706,N_1566,N_2704);
and U7707 (N_7707,N_107,N_1545);
nor U7708 (N_7708,N_3348,N_2601);
xnor U7709 (N_7709,N_1105,N_1953);
and U7710 (N_7710,N_2832,N_1432);
and U7711 (N_7711,N_3643,N_426);
nor U7712 (N_7712,N_1666,N_3571);
xnor U7713 (N_7713,N_2974,N_3389);
xor U7714 (N_7714,N_2712,N_3748);
xor U7715 (N_7715,N_1994,N_456);
nand U7716 (N_7716,N_1081,N_1149);
xnor U7717 (N_7717,N_417,N_3061);
nand U7718 (N_7718,N_2839,N_1020);
xnor U7719 (N_7719,N_85,N_1372);
xnor U7720 (N_7720,N_2813,N_86);
xor U7721 (N_7721,N_1796,N_225);
xor U7722 (N_7722,N_324,N_2828);
xnor U7723 (N_7723,N_1367,N_3362);
and U7724 (N_7724,N_1670,N_951);
xnor U7725 (N_7725,N_2504,N_3287);
nor U7726 (N_7726,N_1618,N_1908);
xor U7727 (N_7727,N_1815,N_3128);
or U7728 (N_7728,N_3313,N_15);
nor U7729 (N_7729,N_1848,N_486);
nand U7730 (N_7730,N_266,N_2821);
or U7731 (N_7731,N_2869,N_2906);
xor U7732 (N_7732,N_3161,N_3421);
or U7733 (N_7733,N_1200,N_3756);
and U7734 (N_7734,N_2312,N_2233);
xor U7735 (N_7735,N_2702,N_1801);
nor U7736 (N_7736,N_3243,N_1481);
or U7737 (N_7737,N_3580,N_2695);
xnor U7738 (N_7738,N_579,N_1301);
or U7739 (N_7739,N_2235,N_3343);
xor U7740 (N_7740,N_2868,N_1297);
nand U7741 (N_7741,N_3009,N_2542);
nor U7742 (N_7742,N_3517,N_1352);
or U7743 (N_7743,N_1984,N_662);
nand U7744 (N_7744,N_2339,N_3324);
xor U7745 (N_7745,N_1093,N_884);
xnor U7746 (N_7746,N_1885,N_3452);
and U7747 (N_7747,N_3005,N_86);
nor U7748 (N_7748,N_2554,N_3883);
xnor U7749 (N_7749,N_2493,N_1282);
xnor U7750 (N_7750,N_3521,N_10);
xnor U7751 (N_7751,N_3943,N_2211);
xnor U7752 (N_7752,N_2143,N_1739);
xnor U7753 (N_7753,N_2561,N_300);
and U7754 (N_7754,N_2095,N_943);
or U7755 (N_7755,N_1342,N_1029);
and U7756 (N_7756,N_3877,N_3010);
nand U7757 (N_7757,N_966,N_3028);
or U7758 (N_7758,N_1612,N_2471);
nand U7759 (N_7759,N_335,N_3652);
nand U7760 (N_7760,N_771,N_3020);
or U7761 (N_7761,N_3945,N_874);
nand U7762 (N_7762,N_144,N_10);
or U7763 (N_7763,N_1735,N_2806);
nor U7764 (N_7764,N_1218,N_1501);
xnor U7765 (N_7765,N_1408,N_2828);
nand U7766 (N_7766,N_3322,N_3754);
and U7767 (N_7767,N_264,N_798);
or U7768 (N_7768,N_1077,N_2724);
and U7769 (N_7769,N_2832,N_1368);
nand U7770 (N_7770,N_3719,N_759);
nand U7771 (N_7771,N_0,N_3175);
or U7772 (N_7772,N_682,N_3350);
xor U7773 (N_7773,N_3274,N_639);
and U7774 (N_7774,N_500,N_2481);
nand U7775 (N_7775,N_2749,N_1186);
or U7776 (N_7776,N_1508,N_816);
and U7777 (N_7777,N_1851,N_3898);
nand U7778 (N_7778,N_2264,N_3498);
or U7779 (N_7779,N_169,N_3036);
nand U7780 (N_7780,N_3839,N_1395);
or U7781 (N_7781,N_1609,N_1343);
and U7782 (N_7782,N_195,N_2475);
nand U7783 (N_7783,N_500,N_1542);
nand U7784 (N_7784,N_1751,N_1666);
or U7785 (N_7785,N_3996,N_751);
nand U7786 (N_7786,N_1525,N_1106);
nor U7787 (N_7787,N_3355,N_1647);
or U7788 (N_7788,N_1925,N_1793);
or U7789 (N_7789,N_3862,N_1642);
nor U7790 (N_7790,N_2380,N_3315);
or U7791 (N_7791,N_249,N_1402);
nor U7792 (N_7792,N_1395,N_3922);
nand U7793 (N_7793,N_3329,N_330);
nand U7794 (N_7794,N_1633,N_314);
nor U7795 (N_7795,N_2335,N_3577);
or U7796 (N_7796,N_902,N_243);
xnor U7797 (N_7797,N_508,N_3254);
or U7798 (N_7798,N_2138,N_1172);
and U7799 (N_7799,N_1255,N_3719);
or U7800 (N_7800,N_1263,N_3708);
nor U7801 (N_7801,N_2020,N_3933);
nand U7802 (N_7802,N_3034,N_3985);
xnor U7803 (N_7803,N_1487,N_519);
nor U7804 (N_7804,N_738,N_963);
and U7805 (N_7805,N_120,N_2324);
and U7806 (N_7806,N_3471,N_2201);
nand U7807 (N_7807,N_3360,N_3166);
nand U7808 (N_7808,N_1863,N_939);
or U7809 (N_7809,N_2652,N_2045);
xor U7810 (N_7810,N_2285,N_3387);
xnor U7811 (N_7811,N_502,N_821);
or U7812 (N_7812,N_650,N_1102);
or U7813 (N_7813,N_3518,N_1483);
nor U7814 (N_7814,N_3596,N_1955);
and U7815 (N_7815,N_2878,N_401);
and U7816 (N_7816,N_1993,N_1093);
and U7817 (N_7817,N_2511,N_3603);
nor U7818 (N_7818,N_3437,N_1992);
and U7819 (N_7819,N_789,N_43);
nand U7820 (N_7820,N_3512,N_2564);
nor U7821 (N_7821,N_2470,N_452);
xnor U7822 (N_7822,N_802,N_2827);
and U7823 (N_7823,N_2332,N_2652);
nand U7824 (N_7824,N_3007,N_3530);
and U7825 (N_7825,N_1546,N_2087);
and U7826 (N_7826,N_666,N_1404);
nor U7827 (N_7827,N_1181,N_1746);
and U7828 (N_7828,N_2111,N_37);
or U7829 (N_7829,N_3027,N_2211);
and U7830 (N_7830,N_1506,N_1513);
and U7831 (N_7831,N_3017,N_3357);
or U7832 (N_7832,N_639,N_431);
nand U7833 (N_7833,N_928,N_2290);
and U7834 (N_7834,N_1031,N_1214);
xor U7835 (N_7835,N_46,N_2774);
xnor U7836 (N_7836,N_132,N_2399);
and U7837 (N_7837,N_1926,N_142);
nor U7838 (N_7838,N_1025,N_3423);
nand U7839 (N_7839,N_25,N_108);
or U7840 (N_7840,N_1553,N_2202);
or U7841 (N_7841,N_714,N_3944);
nand U7842 (N_7842,N_254,N_441);
nor U7843 (N_7843,N_3901,N_2089);
or U7844 (N_7844,N_1097,N_1724);
or U7845 (N_7845,N_3494,N_21);
nor U7846 (N_7846,N_926,N_258);
xnor U7847 (N_7847,N_2276,N_3835);
and U7848 (N_7848,N_1641,N_2758);
nor U7849 (N_7849,N_3374,N_3980);
and U7850 (N_7850,N_3119,N_3252);
xnor U7851 (N_7851,N_609,N_669);
nand U7852 (N_7852,N_2823,N_2419);
nand U7853 (N_7853,N_1556,N_3168);
nand U7854 (N_7854,N_722,N_1343);
and U7855 (N_7855,N_750,N_3730);
xnor U7856 (N_7856,N_39,N_1015);
nor U7857 (N_7857,N_201,N_3143);
nand U7858 (N_7858,N_3291,N_450);
nor U7859 (N_7859,N_3381,N_2098);
nor U7860 (N_7860,N_2290,N_2784);
nand U7861 (N_7861,N_2390,N_3023);
or U7862 (N_7862,N_1793,N_1734);
nor U7863 (N_7863,N_458,N_1702);
nand U7864 (N_7864,N_1669,N_3050);
and U7865 (N_7865,N_2969,N_2278);
nor U7866 (N_7866,N_2306,N_727);
xnor U7867 (N_7867,N_1859,N_3765);
or U7868 (N_7868,N_1086,N_2725);
nor U7869 (N_7869,N_1237,N_2447);
or U7870 (N_7870,N_598,N_1567);
nor U7871 (N_7871,N_3492,N_3169);
and U7872 (N_7872,N_73,N_1522);
and U7873 (N_7873,N_2864,N_3003);
nor U7874 (N_7874,N_3629,N_527);
xnor U7875 (N_7875,N_2913,N_3555);
and U7876 (N_7876,N_2674,N_967);
and U7877 (N_7877,N_820,N_3619);
nand U7878 (N_7878,N_1624,N_3832);
nor U7879 (N_7879,N_2117,N_1002);
xnor U7880 (N_7880,N_1054,N_2606);
or U7881 (N_7881,N_3083,N_855);
xor U7882 (N_7882,N_2416,N_1444);
xnor U7883 (N_7883,N_2231,N_9);
nand U7884 (N_7884,N_2470,N_3182);
or U7885 (N_7885,N_3590,N_136);
nor U7886 (N_7886,N_2802,N_3741);
or U7887 (N_7887,N_2519,N_2056);
xnor U7888 (N_7888,N_690,N_3338);
and U7889 (N_7889,N_726,N_917);
nand U7890 (N_7890,N_964,N_2948);
and U7891 (N_7891,N_1987,N_1550);
or U7892 (N_7892,N_3766,N_1695);
nand U7893 (N_7893,N_2828,N_1678);
nand U7894 (N_7894,N_3504,N_2074);
and U7895 (N_7895,N_563,N_738);
xor U7896 (N_7896,N_1073,N_1250);
or U7897 (N_7897,N_2497,N_1752);
and U7898 (N_7898,N_1875,N_3182);
nor U7899 (N_7899,N_436,N_2933);
and U7900 (N_7900,N_2503,N_3945);
xor U7901 (N_7901,N_3070,N_3599);
or U7902 (N_7902,N_875,N_1687);
nand U7903 (N_7903,N_1108,N_949);
xor U7904 (N_7904,N_1267,N_3542);
nor U7905 (N_7905,N_1107,N_2500);
nor U7906 (N_7906,N_1074,N_3238);
and U7907 (N_7907,N_2613,N_2799);
nor U7908 (N_7908,N_1602,N_428);
nand U7909 (N_7909,N_2303,N_1265);
nand U7910 (N_7910,N_2877,N_2860);
nor U7911 (N_7911,N_664,N_1032);
nor U7912 (N_7912,N_2999,N_3676);
and U7913 (N_7913,N_1258,N_808);
nand U7914 (N_7914,N_2000,N_2538);
and U7915 (N_7915,N_35,N_3506);
xnor U7916 (N_7916,N_1484,N_546);
nand U7917 (N_7917,N_1805,N_3315);
and U7918 (N_7918,N_1690,N_1100);
nand U7919 (N_7919,N_473,N_501);
or U7920 (N_7920,N_2905,N_2095);
nor U7921 (N_7921,N_1738,N_3224);
or U7922 (N_7922,N_2545,N_1815);
and U7923 (N_7923,N_2964,N_1794);
and U7924 (N_7924,N_2852,N_1872);
nor U7925 (N_7925,N_1314,N_832);
and U7926 (N_7926,N_2965,N_383);
xnor U7927 (N_7927,N_2353,N_2343);
xnor U7928 (N_7928,N_3400,N_799);
and U7929 (N_7929,N_1845,N_2547);
nor U7930 (N_7930,N_1566,N_2606);
nor U7931 (N_7931,N_1337,N_330);
xnor U7932 (N_7932,N_3411,N_1217);
xnor U7933 (N_7933,N_2209,N_3969);
and U7934 (N_7934,N_1924,N_2848);
xor U7935 (N_7935,N_2542,N_3687);
and U7936 (N_7936,N_2915,N_3209);
nand U7937 (N_7937,N_2381,N_2812);
xnor U7938 (N_7938,N_895,N_2569);
xnor U7939 (N_7939,N_3059,N_3228);
nor U7940 (N_7940,N_3031,N_1051);
xnor U7941 (N_7941,N_2519,N_1624);
or U7942 (N_7942,N_3170,N_542);
or U7943 (N_7943,N_2533,N_3893);
or U7944 (N_7944,N_1852,N_1233);
or U7945 (N_7945,N_467,N_1983);
nor U7946 (N_7946,N_1433,N_2222);
nand U7947 (N_7947,N_637,N_3518);
and U7948 (N_7948,N_2584,N_1769);
xor U7949 (N_7949,N_2666,N_2194);
or U7950 (N_7950,N_1223,N_3110);
xor U7951 (N_7951,N_1995,N_2409);
nand U7952 (N_7952,N_3026,N_9);
or U7953 (N_7953,N_531,N_2554);
nor U7954 (N_7954,N_3177,N_3330);
nor U7955 (N_7955,N_1298,N_3330);
and U7956 (N_7956,N_314,N_2758);
nor U7957 (N_7957,N_473,N_2633);
or U7958 (N_7958,N_2380,N_2484);
nand U7959 (N_7959,N_1074,N_2486);
xor U7960 (N_7960,N_215,N_3858);
nand U7961 (N_7961,N_1617,N_448);
and U7962 (N_7962,N_980,N_1841);
nor U7963 (N_7963,N_1193,N_151);
or U7964 (N_7964,N_3658,N_89);
nand U7965 (N_7965,N_2394,N_2416);
or U7966 (N_7966,N_466,N_2673);
or U7967 (N_7967,N_3989,N_286);
nand U7968 (N_7968,N_2998,N_3798);
nand U7969 (N_7969,N_1445,N_3711);
nor U7970 (N_7970,N_277,N_5);
nor U7971 (N_7971,N_3566,N_3391);
or U7972 (N_7972,N_688,N_3311);
or U7973 (N_7973,N_1437,N_653);
nand U7974 (N_7974,N_631,N_3206);
xor U7975 (N_7975,N_1800,N_3667);
nand U7976 (N_7976,N_294,N_3407);
nor U7977 (N_7977,N_2201,N_2327);
xor U7978 (N_7978,N_2250,N_3020);
and U7979 (N_7979,N_1177,N_3829);
nor U7980 (N_7980,N_3297,N_3236);
nand U7981 (N_7981,N_1547,N_611);
nor U7982 (N_7982,N_3999,N_3123);
and U7983 (N_7983,N_802,N_645);
xor U7984 (N_7984,N_3036,N_536);
xor U7985 (N_7985,N_3129,N_2167);
xor U7986 (N_7986,N_597,N_1616);
nand U7987 (N_7987,N_3841,N_1313);
and U7988 (N_7988,N_2345,N_1609);
nand U7989 (N_7989,N_2211,N_3743);
nor U7990 (N_7990,N_3247,N_2262);
nand U7991 (N_7991,N_1713,N_740);
or U7992 (N_7992,N_136,N_2135);
nand U7993 (N_7993,N_1724,N_2580);
or U7994 (N_7994,N_301,N_1679);
nand U7995 (N_7995,N_209,N_2600);
or U7996 (N_7996,N_1881,N_400);
xnor U7997 (N_7997,N_2756,N_2605);
xor U7998 (N_7998,N_2447,N_2307);
xor U7999 (N_7999,N_1276,N_3154);
or U8000 (N_8000,N_5686,N_4536);
nand U8001 (N_8001,N_6435,N_7096);
xnor U8002 (N_8002,N_7976,N_5786);
xnor U8003 (N_8003,N_4670,N_5919);
nor U8004 (N_8004,N_7233,N_6286);
nand U8005 (N_8005,N_5925,N_4209);
nand U8006 (N_8006,N_5666,N_6314);
or U8007 (N_8007,N_6759,N_5589);
xnor U8008 (N_8008,N_4838,N_6019);
and U8009 (N_8009,N_6091,N_4099);
nand U8010 (N_8010,N_5213,N_4085);
nor U8011 (N_8011,N_5565,N_6264);
and U8012 (N_8012,N_7048,N_4003);
xnor U8013 (N_8013,N_5246,N_5875);
xor U8014 (N_8014,N_6026,N_4278);
nand U8015 (N_8015,N_7305,N_5651);
nor U8016 (N_8016,N_5777,N_7139);
or U8017 (N_8017,N_7847,N_7119);
xnor U8018 (N_8018,N_7970,N_6644);
and U8019 (N_8019,N_4100,N_7310);
or U8020 (N_8020,N_5753,N_5042);
or U8021 (N_8021,N_6399,N_6084);
and U8022 (N_8022,N_4873,N_7682);
and U8023 (N_8023,N_4671,N_6082);
xor U8024 (N_8024,N_7498,N_6604);
or U8025 (N_8025,N_6169,N_4999);
and U8026 (N_8026,N_5233,N_4458);
and U8027 (N_8027,N_5820,N_6765);
or U8028 (N_8028,N_5403,N_6320);
and U8029 (N_8029,N_4421,N_7930);
and U8030 (N_8030,N_6700,N_6027);
and U8031 (N_8031,N_4729,N_4684);
xnor U8032 (N_8032,N_6328,N_5255);
nor U8033 (N_8033,N_5383,N_4176);
nor U8034 (N_8034,N_5755,N_6959);
xnor U8035 (N_8035,N_6887,N_6459);
and U8036 (N_8036,N_6311,N_6442);
nor U8037 (N_8037,N_7629,N_7858);
or U8038 (N_8038,N_7422,N_6635);
and U8039 (N_8039,N_5237,N_5927);
nor U8040 (N_8040,N_7525,N_6977);
or U8041 (N_8041,N_7809,N_7217);
and U8042 (N_8042,N_4706,N_5493);
or U8043 (N_8043,N_4925,N_7785);
nand U8044 (N_8044,N_4403,N_4881);
nand U8045 (N_8045,N_6258,N_5293);
and U8046 (N_8046,N_5949,N_7000);
or U8047 (N_8047,N_5936,N_5709);
xor U8048 (N_8048,N_4444,N_7739);
nor U8049 (N_8049,N_5609,N_5327);
xnor U8050 (N_8050,N_5997,N_5215);
and U8051 (N_8051,N_5677,N_7447);
or U8052 (N_8052,N_5521,N_5423);
nor U8053 (N_8053,N_4262,N_4975);
nor U8054 (N_8054,N_6556,N_6770);
nand U8055 (N_8055,N_5156,N_4328);
nand U8056 (N_8056,N_4185,N_5010);
nor U8057 (N_8057,N_6901,N_4463);
or U8058 (N_8058,N_5166,N_7870);
and U8059 (N_8059,N_6637,N_6292);
nor U8060 (N_8060,N_4749,N_6496);
and U8061 (N_8061,N_5445,N_6192);
and U8062 (N_8062,N_5569,N_5228);
xor U8063 (N_8063,N_7397,N_7430);
nand U8064 (N_8064,N_7060,N_6937);
xnor U8065 (N_8065,N_5204,N_6089);
or U8066 (N_8066,N_5514,N_6346);
nor U8067 (N_8067,N_4139,N_5211);
nor U8068 (N_8068,N_5703,N_4007);
nand U8069 (N_8069,N_5003,N_4534);
xnor U8070 (N_8070,N_5803,N_5561);
nand U8071 (N_8071,N_6131,N_7802);
or U8072 (N_8072,N_7883,N_7330);
xor U8073 (N_8073,N_6003,N_7579);
xnor U8074 (N_8074,N_7088,N_6821);
and U8075 (N_8075,N_4108,N_5274);
xor U8076 (N_8076,N_7190,N_6795);
xor U8077 (N_8077,N_5314,N_4736);
nand U8078 (N_8078,N_4618,N_6119);
and U8079 (N_8079,N_6491,N_4906);
and U8080 (N_8080,N_4845,N_6042);
nand U8081 (N_8081,N_5349,N_6515);
and U8082 (N_8082,N_7024,N_5184);
nor U8083 (N_8083,N_7596,N_4627);
nand U8084 (N_8084,N_5548,N_4713);
or U8085 (N_8085,N_4979,N_4771);
or U8086 (N_8086,N_7303,N_5095);
xnor U8087 (N_8087,N_6362,N_5100);
xor U8088 (N_8088,N_7507,N_7594);
xor U8089 (N_8089,N_4383,N_4254);
nand U8090 (N_8090,N_6088,N_5976);
or U8091 (N_8091,N_6625,N_7894);
nor U8092 (N_8092,N_7974,N_6798);
and U8093 (N_8093,N_4918,N_7972);
nor U8094 (N_8094,N_4561,N_5394);
nor U8095 (N_8095,N_5887,N_6121);
or U8096 (N_8096,N_4879,N_5012);
or U8097 (N_8097,N_7202,N_6882);
and U8098 (N_8098,N_4700,N_4689);
xnor U8099 (N_8099,N_7353,N_7228);
or U8100 (N_8100,N_6032,N_4158);
xor U8101 (N_8101,N_4018,N_5279);
and U8102 (N_8102,N_4593,N_7725);
nor U8103 (N_8103,N_7775,N_6253);
and U8104 (N_8104,N_6841,N_5115);
nand U8105 (N_8105,N_4981,N_7319);
nor U8106 (N_8106,N_7999,N_5412);
or U8107 (N_8107,N_7003,N_7044);
or U8108 (N_8108,N_6373,N_5417);
nand U8109 (N_8109,N_4516,N_7564);
or U8110 (N_8110,N_4560,N_7335);
nand U8111 (N_8111,N_5057,N_5190);
nand U8112 (N_8112,N_4799,N_5853);
or U8113 (N_8113,N_6024,N_4142);
xor U8114 (N_8114,N_4371,N_7278);
xnor U8115 (N_8115,N_7997,N_4160);
or U8116 (N_8116,N_7328,N_4407);
nand U8117 (N_8117,N_6233,N_6554);
xnor U8118 (N_8118,N_4600,N_6403);
or U8119 (N_8119,N_4079,N_7144);
nor U8120 (N_8120,N_5076,N_7573);
nor U8121 (N_8121,N_7534,N_6610);
nor U8122 (N_8122,N_6230,N_7929);
nand U8123 (N_8123,N_4204,N_5982);
xor U8124 (N_8124,N_6334,N_7206);
and U8125 (N_8125,N_6071,N_4166);
or U8126 (N_8126,N_7711,N_6506);
xnor U8127 (N_8127,N_7820,N_6653);
nand U8128 (N_8128,N_5835,N_4459);
nor U8129 (N_8129,N_7313,N_4575);
xor U8130 (N_8130,N_7674,N_4569);
nor U8131 (N_8131,N_7668,N_4573);
nor U8132 (N_8132,N_7673,N_4062);
nor U8133 (N_8133,N_4287,N_5747);
nor U8134 (N_8134,N_5942,N_6492);
or U8135 (N_8135,N_4603,N_7936);
and U8136 (N_8136,N_5087,N_6113);
and U8137 (N_8137,N_7355,N_7829);
nor U8138 (N_8138,N_5231,N_5890);
nor U8139 (N_8139,N_5765,N_4572);
and U8140 (N_8140,N_7720,N_6702);
nand U8141 (N_8141,N_7680,N_7971);
or U8142 (N_8142,N_6087,N_5583);
nor U8143 (N_8143,N_5490,N_6828);
xnor U8144 (N_8144,N_5483,N_4563);
nand U8145 (N_8145,N_7757,N_4261);
nor U8146 (N_8146,N_5200,N_5431);
xnor U8147 (N_8147,N_5654,N_4368);
nor U8148 (N_8148,N_6561,N_6249);
or U8149 (N_8149,N_4414,N_7798);
and U8150 (N_8150,N_5433,N_4239);
nand U8151 (N_8151,N_4241,N_6200);
xor U8152 (N_8152,N_5921,N_7194);
and U8153 (N_8153,N_6667,N_7158);
nor U8154 (N_8154,N_4882,N_5612);
xnor U8155 (N_8155,N_6085,N_6592);
and U8156 (N_8156,N_7318,N_4682);
or U8157 (N_8157,N_5261,N_5014);
nand U8158 (N_8158,N_6699,N_5754);
xor U8159 (N_8159,N_6966,N_4098);
nor U8160 (N_8160,N_6464,N_7253);
or U8161 (N_8161,N_5733,N_5234);
nor U8162 (N_8162,N_6234,N_6438);
and U8163 (N_8163,N_5044,N_7382);
or U8164 (N_8164,N_6248,N_6886);
or U8165 (N_8165,N_5800,N_5779);
or U8166 (N_8166,N_4372,N_4657);
and U8167 (N_8167,N_5103,N_6444);
nor U8168 (N_8168,N_4978,N_4112);
or U8169 (N_8169,N_5716,N_7499);
nor U8170 (N_8170,N_7376,N_4402);
or U8171 (N_8171,N_6753,N_5556);
and U8172 (N_8172,N_5099,N_4299);
and U8173 (N_8173,N_4964,N_4221);
or U8174 (N_8174,N_4253,N_4486);
or U8175 (N_8175,N_6266,N_6204);
nand U8176 (N_8176,N_5298,N_5283);
or U8177 (N_8177,N_4794,N_5790);
nand U8178 (N_8178,N_7654,N_7022);
or U8179 (N_8179,N_5524,N_7331);
nand U8180 (N_8180,N_4584,N_6251);
nand U8181 (N_8181,N_6460,N_7272);
nand U8182 (N_8182,N_6244,N_4776);
nor U8183 (N_8183,N_6914,N_5460);
or U8184 (N_8184,N_5407,N_5880);
xor U8185 (N_8185,N_7617,N_5276);
nor U8186 (N_8186,N_6895,N_6980);
nor U8187 (N_8187,N_7645,N_4240);
nand U8188 (N_8188,N_5128,N_6735);
nand U8189 (N_8189,N_6861,N_6796);
and U8190 (N_8190,N_4958,N_5983);
or U8191 (N_8191,N_6158,N_4592);
and U8192 (N_8192,N_7098,N_7954);
xor U8193 (N_8193,N_7411,N_6767);
nand U8194 (N_8194,N_5140,N_4988);
and U8195 (N_8195,N_7333,N_5110);
and U8196 (N_8196,N_5148,N_5415);
xor U8197 (N_8197,N_6427,N_5097);
nand U8198 (N_8198,N_4417,N_6504);
xor U8199 (N_8199,N_7016,N_5635);
nor U8200 (N_8200,N_5137,N_6799);
nand U8201 (N_8201,N_5046,N_5817);
nor U8202 (N_8202,N_4331,N_4909);
nand U8203 (N_8203,N_6407,N_5322);
xnor U8204 (N_8204,N_4191,N_7759);
nor U8205 (N_8205,N_4440,N_6546);
or U8206 (N_8206,N_5304,N_7213);
or U8207 (N_8207,N_7203,N_6331);
and U8208 (N_8208,N_7643,N_7708);
xor U8209 (N_8209,N_6065,N_4704);
or U8210 (N_8210,N_6171,N_7616);
xor U8211 (N_8211,N_7961,N_5068);
nor U8212 (N_8212,N_6811,N_6381);
or U8213 (N_8213,N_7084,N_5009);
xor U8214 (N_8214,N_6899,N_4103);
xor U8215 (N_8215,N_7501,N_7293);
and U8216 (N_8216,N_6461,N_5756);
xor U8217 (N_8217,N_7298,N_5264);
or U8218 (N_8218,N_7769,N_7689);
or U8219 (N_8219,N_7188,N_5638);
nor U8220 (N_8220,N_4753,N_6724);
xor U8221 (N_8221,N_7345,N_7101);
xor U8222 (N_8222,N_7666,N_7089);
and U8223 (N_8223,N_5713,N_4597);
xnor U8224 (N_8224,N_7286,N_7464);
nand U8225 (N_8225,N_7237,N_4654);
nor U8226 (N_8226,N_6415,N_4567);
nor U8227 (N_8227,N_5792,N_6788);
nor U8228 (N_8228,N_4957,N_4798);
and U8229 (N_8229,N_5449,N_4778);
xor U8230 (N_8230,N_7749,N_7209);
or U8231 (N_8231,N_4376,N_7923);
nand U8232 (N_8232,N_4849,N_7690);
xor U8233 (N_8233,N_5888,N_5426);
or U8234 (N_8234,N_7231,N_6284);
nand U8235 (N_8235,N_6099,N_7037);
or U8236 (N_8236,N_7518,N_7425);
nand U8237 (N_8237,N_4012,N_5176);
xnor U8238 (N_8238,N_6695,N_6650);
xnor U8239 (N_8239,N_4820,N_4456);
or U8240 (N_8240,N_5785,N_5039);
nand U8241 (N_8241,N_5051,N_6478);
nor U8242 (N_8242,N_4038,N_6487);
xnor U8243 (N_8243,N_7861,N_6547);
nand U8244 (N_8244,N_5249,N_5650);
and U8245 (N_8245,N_6618,N_4770);
nor U8246 (N_8246,N_7812,N_5189);
xor U8247 (N_8247,N_5430,N_7186);
nor U8248 (N_8248,N_5389,N_5992);
xnor U8249 (N_8249,N_7788,N_6866);
and U8250 (N_8250,N_7106,N_6536);
nand U8251 (N_8251,N_7919,N_4015);
nand U8252 (N_8252,N_6455,N_5463);
nand U8253 (N_8253,N_4467,N_4468);
nor U8254 (N_8254,N_6100,N_4984);
xor U8255 (N_8255,N_7362,N_7289);
nand U8256 (N_8256,N_5109,N_6458);
nand U8257 (N_8257,N_4844,N_5610);
nor U8258 (N_8258,N_7255,N_4392);
xnor U8259 (N_8259,N_6350,N_4303);
nand U8260 (N_8260,N_7762,N_4867);
or U8261 (N_8261,N_7364,N_6275);
or U8262 (N_8262,N_4009,N_6053);
nor U8263 (N_8263,N_7577,N_7783);
nor U8264 (N_8264,N_6832,N_7124);
nor U8265 (N_8265,N_4452,N_6462);
nor U8266 (N_8266,N_7572,N_5341);
or U8267 (N_8267,N_7181,N_4435);
or U8268 (N_8268,N_7995,N_6897);
and U8269 (N_8269,N_4117,N_7230);
nand U8270 (N_8270,N_4310,N_6179);
and U8271 (N_8271,N_4132,N_5542);
and U8272 (N_8272,N_6921,N_6274);
and U8273 (N_8273,N_6007,N_6578);
nand U8274 (N_8274,N_6909,N_6060);
and U8275 (N_8275,N_6668,N_4217);
nand U8276 (N_8276,N_5294,N_6593);
and U8277 (N_8277,N_6675,N_4939);
xnor U8278 (N_8278,N_5823,N_7996);
nand U8279 (N_8279,N_6202,N_5476);
nand U8280 (N_8280,N_6992,N_4199);
or U8281 (N_8281,N_6135,N_7859);
nor U8282 (N_8282,N_7457,N_4974);
xor U8283 (N_8283,N_6540,N_4248);
nand U8284 (N_8284,N_5985,N_4041);
nand U8285 (N_8285,N_7872,N_5523);
or U8286 (N_8286,N_6919,N_4963);
nand U8287 (N_8287,N_6271,N_5954);
and U8288 (N_8288,N_5735,N_6645);
and U8289 (N_8289,N_7151,N_4751);
nand U8290 (N_8290,N_5029,N_6490);
xnor U8291 (N_8291,N_6047,N_7803);
nor U8292 (N_8292,N_5065,N_4748);
xor U8293 (N_8293,N_6391,N_7655);
nor U8294 (N_8294,N_5136,N_4045);
nand U8295 (N_8295,N_5059,N_5938);
nand U8296 (N_8296,N_5512,N_6541);
and U8297 (N_8297,N_7201,N_4238);
nand U8298 (N_8298,N_4551,N_5002);
xnor U8299 (N_8299,N_6107,N_6104);
nor U8300 (N_8300,N_6693,N_6711);
nand U8301 (N_8301,N_7307,N_7160);
nand U8302 (N_8302,N_6090,N_7465);
nand U8303 (N_8303,N_7412,N_7477);
or U8304 (N_8304,N_5229,N_5152);
or U8305 (N_8305,N_5006,N_6378);
nand U8306 (N_8306,N_7892,N_7746);
xor U8307 (N_8307,N_6539,N_6446);
nand U8308 (N_8308,N_7012,N_5209);
and U8309 (N_8309,N_7570,N_6452);
nor U8310 (N_8310,N_4789,N_5257);
and U8311 (N_8311,N_7831,N_5480);
and U8312 (N_8312,N_7890,N_5477);
xnor U8313 (N_8313,N_6359,N_6660);
or U8314 (N_8314,N_7463,N_5054);
xor U8315 (N_8315,N_5282,N_7434);
nor U8316 (N_8316,N_6126,N_5337);
xnor U8317 (N_8317,N_5865,N_7911);
and U8318 (N_8318,N_6370,N_6228);
and U8319 (N_8319,N_7446,N_4497);
nand U8320 (N_8320,N_4752,N_6960);
and U8321 (N_8321,N_6677,N_5132);
or U8322 (N_8322,N_4201,N_5309);
or U8323 (N_8323,N_6979,N_6039);
xor U8324 (N_8324,N_5434,N_4650);
or U8325 (N_8325,N_5290,N_7719);
nand U8326 (N_8326,N_6077,N_7659);
nor U8327 (N_8327,N_7386,N_4431);
nor U8328 (N_8328,N_5035,N_5766);
nand U8329 (N_8329,N_7508,N_7854);
nor U8330 (N_8330,N_6873,N_7410);
or U8331 (N_8331,N_6754,N_7952);
and U8332 (N_8332,N_4227,N_4330);
and U8333 (N_8333,N_6422,N_6136);
xor U8334 (N_8334,N_7295,N_6776);
nand U8335 (N_8335,N_5296,N_6568);
nor U8336 (N_8336,N_6844,N_6591);
or U8337 (N_8337,N_7753,N_7462);
xor U8338 (N_8338,N_5826,N_5939);
nand U8339 (N_8339,N_5535,N_6252);
nand U8340 (N_8340,N_7852,N_4797);
nand U8341 (N_8341,N_6752,N_5909);
nand U8342 (N_8342,N_5188,N_5926);
or U8343 (N_8343,N_6820,N_7834);
or U8344 (N_8344,N_6726,N_6269);
xnor U8345 (N_8345,N_6563,N_7069);
or U8346 (N_8346,N_5288,N_7320);
xor U8347 (N_8347,N_5578,N_4149);
or U8348 (N_8348,N_7322,N_4134);
or U8349 (N_8349,N_5157,N_6582);
and U8350 (N_8350,N_5697,N_5683);
nor U8351 (N_8351,N_4515,N_4430);
and U8352 (N_8352,N_7943,N_4523);
and U8353 (N_8353,N_5558,N_7724);
nand U8354 (N_8354,N_6656,N_6041);
nand U8355 (N_8355,N_7049,N_6925);
nor U8356 (N_8356,N_6709,N_5810);
nor U8357 (N_8357,N_4295,N_7374);
nor U8358 (N_8358,N_4314,N_5883);
and U8359 (N_8359,N_4510,N_7728);
or U8360 (N_8360,N_7704,N_5172);
nor U8361 (N_8361,N_5278,N_6146);
nor U8362 (N_8362,N_7560,N_5267);
nand U8363 (N_8363,N_7765,N_4664);
or U8364 (N_8364,N_5685,N_6559);
nor U8365 (N_8365,N_4047,N_5427);
xor U8366 (N_8366,N_5915,N_7758);
and U8367 (N_8367,N_4023,N_7801);
and U8368 (N_8368,N_6936,N_4812);
or U8369 (N_8369,N_5838,N_5967);
nor U8370 (N_8370,N_7350,N_4090);
and U8371 (N_8371,N_5284,N_6383);
or U8372 (N_8372,N_6166,N_4089);
nand U8373 (N_8373,N_6846,N_5272);
xnor U8374 (N_8374,N_5472,N_7405);
nand U8375 (N_8375,N_5382,N_7169);
and U8376 (N_8376,N_4623,N_5644);
or U8377 (N_8377,N_5575,N_5637);
and U8378 (N_8378,N_6658,N_7061);
or U8379 (N_8379,N_4271,N_6893);
nor U8380 (N_8380,N_7977,N_5707);
xnor U8381 (N_8381,N_7848,N_6574);
nor U8382 (N_8382,N_7926,N_4503);
xnor U8383 (N_8383,N_6967,N_7326);
or U8384 (N_8384,N_4629,N_4070);
or U8385 (N_8385,N_5491,N_5311);
nor U8386 (N_8386,N_7085,N_7232);
nor U8387 (N_8387,N_4276,N_4605);
xor U8388 (N_8388,N_7933,N_5958);
nor U8389 (N_8389,N_6222,N_5884);
and U8390 (N_8390,N_5050,N_7161);
or U8391 (N_8391,N_6527,N_5834);
or U8392 (N_8392,N_6564,N_6508);
nand U8393 (N_8393,N_4533,N_6819);
xor U8394 (N_8394,N_5413,N_5180);
nand U8395 (N_8395,N_7850,N_6175);
nand U8396 (N_8396,N_4487,N_7437);
or U8397 (N_8397,N_7723,N_4300);
or U8398 (N_8398,N_6984,N_4116);
nand U8399 (N_8399,N_7262,N_6127);
nor U8400 (N_8400,N_6953,N_4692);
and U8401 (N_8401,N_6868,N_5398);
or U8402 (N_8402,N_4839,N_4231);
and U8403 (N_8403,N_4842,N_4944);
or U8404 (N_8404,N_4399,N_7945);
xnor U8405 (N_8405,N_6017,N_6774);
nand U8406 (N_8406,N_5776,N_7214);
and U8407 (N_8407,N_5253,N_4270);
or U8408 (N_8408,N_7165,N_4352);
and U8409 (N_8409,N_6607,N_4756);
nor U8410 (N_8410,N_4324,N_6137);
nand U8411 (N_8411,N_5139,N_6079);
or U8412 (N_8412,N_6758,N_6766);
nor U8413 (N_8413,N_7433,N_6229);
and U8414 (N_8414,N_7524,N_6296);
or U8415 (N_8415,N_7302,N_7367);
nor U8416 (N_8416,N_6588,N_5328);
nor U8417 (N_8417,N_5673,N_6646);
nand U8418 (N_8418,N_7291,N_5443);
and U8419 (N_8419,N_7274,N_4308);
and U8420 (N_8420,N_4024,N_5592);
and U8421 (N_8421,N_5120,N_6297);
or U8422 (N_8422,N_6513,N_4790);
nand U8423 (N_8423,N_5235,N_5814);
or U8424 (N_8424,N_5966,N_6521);
xor U8425 (N_8425,N_4195,N_7445);
nand U8426 (N_8426,N_6096,N_4102);
nor U8427 (N_8427,N_5342,N_7480);
nor U8428 (N_8428,N_5153,N_7806);
xnor U8429 (N_8429,N_6876,N_6694);
xor U8430 (N_8430,N_4601,N_7729);
nor U8431 (N_8431,N_7369,N_5581);
nor U8432 (N_8432,N_4211,N_4907);
nand U8433 (N_8433,N_7460,N_7162);
nand U8434 (N_8434,N_7876,N_6425);
or U8435 (N_8435,N_4883,N_6982);
or U8436 (N_8436,N_7251,N_7222);
nor U8437 (N_8437,N_4937,N_6302);
or U8438 (N_8438,N_6057,N_7844);
and U8439 (N_8439,N_5981,N_4189);
and U8440 (N_8440,N_5669,N_7799);
nor U8441 (N_8441,N_4923,N_5271);
nand U8442 (N_8442,N_6343,N_5321);
and U8443 (N_8443,N_7939,N_4080);
and U8444 (N_8444,N_7384,N_5998);
nand U8445 (N_8445,N_5496,N_5961);
nor U8446 (N_8446,N_4942,N_6920);
and U8447 (N_8447,N_4986,N_4680);
xor U8448 (N_8448,N_7562,N_4316);
or U8449 (N_8449,N_5912,N_5841);
and U8450 (N_8450,N_4955,N_6998);
xnor U8451 (N_8451,N_4767,N_4181);
nand U8452 (N_8452,N_4606,N_7709);
xnor U8453 (N_8453,N_4707,N_5344);
and U8454 (N_8454,N_7816,N_6288);
nor U8455 (N_8455,N_7781,N_4448);
or U8456 (N_8456,N_5175,N_5993);
nor U8457 (N_8457,N_5316,N_5080);
nor U8458 (N_8458,N_7034,N_7440);
nor U8459 (N_8459,N_6836,N_7587);
or U8460 (N_8460,N_5366,N_6737);
xor U8461 (N_8461,N_6631,N_4759);
xnor U8462 (N_8462,N_7697,N_7389);
nor U8463 (N_8463,N_4810,N_7567);
nand U8464 (N_8464,N_6584,N_4594);
and U8465 (N_8465,N_4137,N_5027);
nand U8466 (N_8466,N_5079,N_7884);
nor U8467 (N_8467,N_7893,N_4246);
nand U8468 (N_8468,N_5395,N_7885);
nor U8469 (N_8469,N_6214,N_4951);
or U8470 (N_8470,N_6557,N_4162);
nand U8471 (N_8471,N_7716,N_6197);
xnor U8472 (N_8472,N_6898,N_6958);
and U8473 (N_8473,N_4768,N_5595);
nor U8474 (N_8474,N_7613,N_7955);
xnor U8475 (N_8475,N_5808,N_5658);
nand U8476 (N_8476,N_4866,N_7946);
nand U8477 (N_8477,N_7082,N_7441);
nand U8478 (N_8478,N_4972,N_4422);
nand U8479 (N_8479,N_7978,N_4390);
or U8480 (N_8480,N_7862,N_7123);
xnor U8481 (N_8481,N_5141,N_5094);
nor U8482 (N_8482,N_4348,N_5931);
xor U8483 (N_8483,N_6125,N_5601);
and U8484 (N_8484,N_5183,N_5024);
nor U8485 (N_8485,N_4291,N_4110);
and U8486 (N_8486,N_7150,N_7640);
nor U8487 (N_8487,N_6410,N_5177);
xor U8488 (N_8488,N_6738,N_7621);
xnor U8489 (N_8489,N_7242,N_4095);
nor U8490 (N_8490,N_5971,N_4679);
nand U8491 (N_8491,N_6560,N_6883);
nor U8492 (N_8492,N_5361,N_5886);
nor U8493 (N_8493,N_5317,N_5406);
nand U8494 (N_8494,N_4658,N_4107);
and U8495 (N_8495,N_7630,N_7368);
nand U8496 (N_8496,N_5292,N_4474);
nand U8497 (N_8497,N_4847,N_5326);
xor U8498 (N_8498,N_6161,N_6713);
nor U8499 (N_8499,N_6888,N_4581);
nand U8500 (N_8500,N_4512,N_6045);
nor U8501 (N_8501,N_7281,N_6122);
or U8502 (N_8502,N_7273,N_4609);
nand U8503 (N_8503,N_7647,N_7207);
nand U8504 (N_8504,N_7731,N_6388);
nor U8505 (N_8505,N_5354,N_4053);
xor U8506 (N_8506,N_5332,N_7268);
and U8507 (N_8507,N_4354,N_4877);
nor U8508 (N_8508,N_6316,N_6479);
nor U8509 (N_8509,N_7135,N_7735);
and U8510 (N_8510,N_6358,N_5421);
nor U8511 (N_8511,N_5362,N_7490);
or U8512 (N_8512,N_6312,N_4932);
or U8513 (N_8513,N_5989,N_7512);
and U8514 (N_8514,N_6186,N_7905);
and U8515 (N_8515,N_5026,N_7133);
xor U8516 (N_8516,N_6589,N_6360);
or U8517 (N_8517,N_7159,N_6243);
nand U8518 (N_8518,N_4173,N_4690);
nand U8519 (N_8519,N_6185,N_5481);
and U8520 (N_8520,N_6948,N_4744);
and U8521 (N_8521,N_5519,N_5378);
nand U8522 (N_8522,N_4373,N_6285);
and U8523 (N_8523,N_4441,N_5479);
or U8524 (N_8524,N_4578,N_5988);
xor U8525 (N_8525,N_4857,N_4801);
xor U8526 (N_8526,N_5259,N_7467);
xor U8527 (N_8527,N_4129,N_4338);
nor U8528 (N_8528,N_5442,N_7359);
nand U8529 (N_8529,N_7042,N_4822);
nand U8530 (N_8530,N_6237,N_4547);
xor U8531 (N_8531,N_7975,N_4213);
nor U8532 (N_8532,N_7418,N_5784);
nand U8533 (N_8533,N_4126,N_5910);
nand U8534 (N_8534,N_4072,N_4656);
nand U8535 (N_8535,N_5247,N_6154);
or U8536 (N_8536,N_7537,N_5446);
nand U8537 (N_8537,N_4335,N_5108);
nand U8538 (N_8538,N_6986,N_7553);
xor U8539 (N_8539,N_6613,N_5082);
nor U8540 (N_8540,N_5130,N_7900);
xnor U8541 (N_8541,N_6333,N_7492);
nor U8542 (N_8542,N_7707,N_7436);
nor U8543 (N_8543,N_6142,N_7592);
or U8544 (N_8544,N_7244,N_4966);
nand U8545 (N_8545,N_5216,N_7611);
xnor U8546 (N_8546,N_7452,N_7265);
xor U8547 (N_8547,N_5487,N_4983);
nand U8548 (N_8548,N_4445,N_4428);
nand U8549 (N_8549,N_6217,N_5263);
and U8550 (N_8550,N_5867,N_5225);
or U8551 (N_8551,N_7473,N_6354);
and U8552 (N_8552,N_6031,N_7196);
nor U8553 (N_8553,N_5798,N_6174);
nand U8554 (N_8554,N_5088,N_7113);
and U8555 (N_8555,N_7683,N_4566);
and U8556 (N_8556,N_5844,N_5439);
and U8557 (N_8557,N_7316,N_5310);
nor U8558 (N_8558,N_5258,N_6398);
and U8559 (N_8559,N_5762,N_4283);
nand U8560 (N_8560,N_4384,N_4637);
nor U8561 (N_8561,N_5159,N_6262);
nor U8562 (N_8562,N_5662,N_4073);
and U8563 (N_8563,N_7973,N_6235);
nor U8564 (N_8564,N_6128,N_5757);
or U8565 (N_8565,N_7821,N_6250);
and U8566 (N_8566,N_5384,N_7083);
or U8567 (N_8567,N_4040,N_7672);
xnor U8568 (N_8568,N_7363,N_4343);
nand U8569 (N_8569,N_5725,N_7426);
nand U8570 (N_8570,N_4900,N_4553);
xor U8571 (N_8571,N_7609,N_4723);
xor U8572 (N_8572,N_7815,N_5151);
or U8573 (N_8573,N_6981,N_7148);
nor U8574 (N_8574,N_5657,N_5907);
and U8575 (N_8575,N_4028,N_7845);
nor U8576 (N_8576,N_6669,N_5582);
and U8577 (N_8577,N_6859,N_7784);
xor U8578 (N_8578,N_6801,N_4168);
xor U8579 (N_8579,N_4323,N_6015);
nand U8580 (N_8580,N_7050,N_4935);
or U8581 (N_8581,N_5952,N_4538);
nand U8582 (N_8582,N_5829,N_6005);
nor U8583 (N_8583,N_6657,N_7636);
nor U8584 (N_8584,N_5659,N_7324);
or U8585 (N_8585,N_5913,N_7880);
or U8586 (N_8586,N_6777,N_7379);
or U8587 (N_8587,N_4022,N_7669);
or U8588 (N_8588,N_4010,N_6627);
or U8589 (N_8589,N_4885,N_5179);
nor U8590 (N_8590,N_4780,N_7472);
nand U8591 (N_8591,N_6188,N_5369);
nand U8592 (N_8592,N_7075,N_7782);
and U8593 (N_8593,N_5598,N_5849);
xor U8594 (N_8594,N_5078,N_5739);
nor U8595 (N_8595,N_5458,N_6511);
nand U8596 (N_8596,N_4161,N_4333);
or U8597 (N_8597,N_7878,N_5603);
nand U8598 (N_8598,N_7469,N_5870);
xnor U8599 (N_8599,N_7078,N_5712);
or U8600 (N_8600,N_6830,N_5904);
xor U8601 (N_8601,N_4406,N_6226);
or U8602 (N_8602,N_4720,N_7432);
xor U8603 (N_8603,N_6787,N_6678);
and U8604 (N_8604,N_4361,N_5593);
and U8605 (N_8605,N_4889,N_7226);
nor U8606 (N_8606,N_4504,N_4825);
or U8607 (N_8607,N_7420,N_6392);
nand U8608 (N_8608,N_5862,N_4642);
and U8609 (N_8609,N_7413,N_7391);
and U8610 (N_8610,N_4380,N_4728);
nand U8611 (N_8611,N_6522,N_7011);
nand U8612 (N_8612,N_4284,N_5429);
and U8613 (N_8613,N_6189,N_7521);
nor U8614 (N_8614,N_6950,N_4363);
nand U8615 (N_8615,N_6434,N_4321);
or U8616 (N_8616,N_4194,N_4598);
xor U8617 (N_8617,N_6149,N_4815);
or U8618 (N_8618,N_7631,N_5011);
and U8619 (N_8619,N_4084,N_6323);
nand U8620 (N_8620,N_7375,N_5286);
nand U8621 (N_8621,N_7252,N_4763);
nor U8622 (N_8622,N_6183,N_5693);
or U8623 (N_8623,N_6703,N_6000);
nor U8624 (N_8624,N_4643,N_5680);
or U8625 (N_8625,N_4919,N_5016);
and U8626 (N_8626,N_7476,N_4470);
nand U8627 (N_8627,N_6151,N_5195);
and U8628 (N_8628,N_7021,N_5874);
and U8629 (N_8629,N_6771,N_7195);
and U8630 (N_8630,N_4389,N_4946);
and U8631 (N_8631,N_5365,N_4187);
or U8632 (N_8632,N_6433,N_6355);
nand U8633 (N_8633,N_4904,N_5484);
or U8634 (N_8634,N_4218,N_7824);
nor U8635 (N_8635,N_7510,N_4386);
xor U8636 (N_8636,N_4197,N_4150);
xnor U8637 (N_8637,N_5062,N_4841);
xor U8638 (N_8638,N_4762,N_4396);
nand U8639 (N_8639,N_5104,N_5056);
or U8640 (N_8640,N_6353,N_7239);
and U8641 (N_8641,N_5174,N_4631);
nand U8642 (N_8642,N_5782,N_6672);
nand U8643 (N_8643,N_7461,N_5113);
nand U8644 (N_8644,N_6587,N_5007);
and U8645 (N_8645,N_7957,N_4147);
nor U8646 (N_8646,N_5379,N_7540);
nand U8647 (N_8647,N_7653,N_4897);
and U8648 (N_8648,N_5118,N_6431);
or U8649 (N_8649,N_6651,N_7365);
nor U8650 (N_8650,N_4659,N_7138);
nor U8651 (N_8651,N_5559,N_4346);
and U8652 (N_8652,N_5866,N_4302);
xor U8653 (N_8653,N_4863,N_7344);
xnor U8654 (N_8654,N_6822,N_6684);
xor U8655 (N_8655,N_6319,N_7056);
or U8656 (N_8656,N_5048,N_4113);
nor U8657 (N_8657,N_4228,N_7535);
nand U8658 (N_8658,N_6530,N_7401);
or U8659 (N_8659,N_5498,N_7141);
xnor U8660 (N_8660,N_6416,N_5015);
xor U8661 (N_8661,N_7068,N_6803);
xnor U8662 (N_8662,N_7532,N_5710);
nor U8663 (N_8663,N_6313,N_6855);
nand U8664 (N_8664,N_4269,N_6437);
nand U8665 (N_8665,N_4524,N_7311);
xor U8666 (N_8666,N_5456,N_7726);
nand U8667 (N_8667,N_4258,N_4587);
nand U8668 (N_8668,N_4229,N_4876);
nand U8669 (N_8669,N_7429,N_7804);
nor U8670 (N_8670,N_7453,N_7904);
xor U8671 (N_8671,N_4721,N_5796);
or U8672 (N_8672,N_7882,N_4491);
or U8673 (N_8673,N_6309,N_7392);
or U8674 (N_8674,N_7651,N_5055);
xnor U8675 (N_8675,N_4483,N_5937);
and U8676 (N_8676,N_4400,N_6781);
or U8677 (N_8677,N_7602,N_6238);
and U8678 (N_8678,N_7623,N_4992);
xor U8679 (N_8679,N_4086,N_7964);
xnor U8680 (N_8680,N_6916,N_6413);
or U8681 (N_8681,N_7591,N_7204);
and U8682 (N_8682,N_6002,N_7015);
or U8683 (N_8683,N_7205,N_4465);
nor U8684 (N_8684,N_5318,N_7646);
nor U8685 (N_8685,N_4954,N_4950);
nand U8686 (N_8686,N_7544,N_7179);
xor U8687 (N_8687,N_7571,N_6011);
and U8688 (N_8688,N_6147,N_6351);
and U8689 (N_8689,N_7170,N_4641);
xor U8690 (N_8690,N_6681,N_4370);
nand U8691 (N_8691,N_7633,N_7055);
and U8692 (N_8692,N_6810,N_4968);
or U8693 (N_8693,N_5974,N_4469);
or U8694 (N_8694,N_7583,N_7542);
and U8695 (N_8695,N_6385,N_6797);
nor U8696 (N_8696,N_5688,N_4987);
nor U8697 (N_8697,N_6199,N_6549);
nor U8698 (N_8698,N_6764,N_5117);
nor U8699 (N_8699,N_5005,N_7092);
xor U8700 (N_8700,N_5457,N_4746);
and U8701 (N_8701,N_6064,N_7514);
xor U8702 (N_8702,N_7776,N_5464);
or U8703 (N_8703,N_6469,N_6762);
xnor U8704 (N_8704,N_4029,N_7360);
or U8705 (N_8705,N_4930,N_4552);
xor U8706 (N_8706,N_7054,N_6187);
nor U8707 (N_8707,N_6662,N_7466);
or U8708 (N_8708,N_4297,N_7875);
nand U8709 (N_8709,N_5729,N_7180);
nand U8710 (N_8710,N_4829,N_4438);
nand U8711 (N_8711,N_7131,N_5528);
xnor U8712 (N_8712,N_7387,N_6182);
and U8713 (N_8713,N_6287,N_6903);
nor U8714 (N_8714,N_7593,N_5122);
nor U8715 (N_8715,N_5678,N_5114);
or U8716 (N_8716,N_4779,N_4455);
nand U8717 (N_8717,N_4008,N_5550);
nand U8718 (N_8718,N_6594,N_7155);
nand U8719 (N_8719,N_5679,N_6159);
or U8720 (N_8720,N_7734,N_4424);
nand U8721 (N_8721,N_6364,N_7342);
xor U8722 (N_8722,N_6931,N_6736);
and U8723 (N_8723,N_5526,N_7114);
nor U8724 (N_8724,N_7404,N_6585);
and U8725 (N_8725,N_5008,N_6938);
or U8726 (N_8726,N_6679,N_7221);
or U8727 (N_8727,N_7912,N_4724);
or U8728 (N_8728,N_5663,N_6834);
or U8729 (N_8729,N_7910,N_4959);
xnor U8730 (N_8730,N_7863,N_5649);
or U8731 (N_8731,N_4017,N_5553);
or U8732 (N_8732,N_5614,N_7241);
and U8733 (N_8733,N_4317,N_7366);
nor U8734 (N_8734,N_5277,N_4661);
and U8735 (N_8735,N_5631,N_5715);
or U8736 (N_8736,N_7126,N_5897);
or U8737 (N_8737,N_4105,N_4385);
nor U8738 (N_8738,N_6342,N_7143);
or U8739 (N_8739,N_6377,N_4039);
nor U8740 (N_8740,N_4479,N_4886);
nand U8741 (N_8741,N_5617,N_7608);
and U8742 (N_8742,N_4188,N_6940);
nand U8743 (N_8743,N_7035,N_7699);
xor U8744 (N_8744,N_6232,N_6441);
xnor U8745 (N_8745,N_6659,N_6671);
or U8746 (N_8746,N_7770,N_5232);
nand U8747 (N_8747,N_7773,N_4929);
nand U8748 (N_8748,N_7721,N_5218);
xnor U8749 (N_8749,N_7787,N_6831);
nor U8750 (N_8750,N_7810,N_5990);
and U8751 (N_8751,N_7886,N_7898);
or U8752 (N_8752,N_6691,N_6756);
xnor U8753 (N_8753,N_4887,N_7377);
nand U8754 (N_8754,N_7455,N_7130);
or U8755 (N_8755,N_4945,N_7030);
or U8756 (N_8756,N_5422,N_6507);
nand U8757 (N_8757,N_6384,N_6509);
or U8758 (N_8758,N_7182,N_5783);
and U8759 (N_8759,N_6372,N_7442);
or U8760 (N_8760,N_4170,N_6545);
xnor U8761 (N_8761,N_5914,N_6664);
xnor U8762 (N_8762,N_5742,N_7308);
xor U8763 (N_8763,N_5242,N_6265);
nand U8764 (N_8764,N_7010,N_7153);
and U8765 (N_8765,N_7520,N_5576);
nor U8766 (N_8766,N_6375,N_5948);
nand U8767 (N_8767,N_5124,N_5373);
xor U8768 (N_8768,N_4216,N_7023);
or U8769 (N_8769,N_5469,N_5695);
or U8770 (N_8770,N_4802,N_5248);
and U8771 (N_8771,N_4823,N_5254);
nor U8772 (N_8772,N_5780,N_7164);
nand U8773 (N_8773,N_7070,N_4274);
or U8774 (N_8774,N_4537,N_4914);
and U8775 (N_8775,N_7963,N_5339);
or U8776 (N_8776,N_7417,N_5227);
xnor U8777 (N_8777,N_4306,N_4702);
nor U8778 (N_8778,N_5185,N_7622);
or U8779 (N_8779,N_6902,N_6544);
nand U8780 (N_8780,N_5643,N_6745);
and U8781 (N_8781,N_6923,N_6790);
or U8782 (N_8782,N_7513,N_4948);
nor U8783 (N_8783,N_6917,N_6387);
or U8784 (N_8784,N_6957,N_6338);
and U8785 (N_8785,N_7671,N_6386);
nor U8786 (N_8786,N_7825,N_4043);
and U8787 (N_8787,N_4232,N_5545);
nor U8788 (N_8788,N_4737,N_5889);
xor U8789 (N_8789,N_4522,N_4519);
xor U8790 (N_8790,N_6643,N_4687);
xor U8791 (N_8791,N_7229,N_4837);
or U8792 (N_8792,N_6946,N_4869);
xnor U8793 (N_8793,N_5205,N_5830);
nand U8794 (N_8794,N_7053,N_6519);
nor U8795 (N_8795,N_7396,N_4377);
xnor U8796 (N_8796,N_6874,N_5831);
nand U8797 (N_8797,N_4715,N_5187);
xor U8798 (N_8798,N_7751,N_4579);
or U8799 (N_8799,N_4157,N_7352);
nor U8800 (N_8800,N_4521,N_7888);
nand U8801 (N_8801,N_5538,N_5420);
and U8802 (N_8802,N_4275,N_5455);
and U8803 (N_8803,N_5475,N_6969);
or U8804 (N_8804,N_4111,N_4875);
or U8805 (N_8805,N_7941,N_4016);
or U8806 (N_8806,N_7650,N_4153);
nand U8807 (N_8807,N_5034,N_6043);
xor U8808 (N_8808,N_5291,N_4071);
nor U8809 (N_8809,N_7712,N_6303);
and U8810 (N_8810,N_7865,N_6623);
xor U8811 (N_8811,N_5208,N_6739);
and U8812 (N_8812,N_7771,N_5217);
nand U8813 (N_8813,N_6029,N_5127);
nand U8814 (N_8814,N_4864,N_7599);
xnor U8815 (N_8815,N_4446,N_5674);
and U8816 (N_8816,N_7927,N_6349);
nor U8817 (N_8817,N_7294,N_7832);
xnor U8818 (N_8818,N_5932,N_6922);
xor U8819 (N_8819,N_4076,N_4545);
nand U8820 (N_8820,N_4068,N_7129);
or U8821 (N_8821,N_4374,N_4234);
xnor U8822 (N_8822,N_5758,N_5408);
nor U8823 (N_8823,N_5922,N_4808);
and U8824 (N_8824,N_4683,N_4742);
and U8825 (N_8825,N_6722,N_6617);
or U8826 (N_8826,N_6473,N_7547);
and U8827 (N_8827,N_7754,N_6133);
nand U8828 (N_8828,N_4644,N_4765);
xor U8829 (N_8829,N_5623,N_5251);
xor U8830 (N_8830,N_6255,N_6573);
or U8831 (N_8831,N_6366,N_5386);
xor U8832 (N_8832,N_7236,N_5173);
xor U8833 (N_8833,N_6880,N_7415);
nor U8834 (N_8834,N_7626,N_6470);
nand U8835 (N_8835,N_5397,N_5864);
xor U8836 (N_8836,N_6389,N_6793);
xor U8837 (N_8837,N_5905,N_6030);
or U8838 (N_8838,N_5627,N_5499);
nand U8839 (N_8839,N_5517,N_7531);
nand U8840 (N_8840,N_4439,N_4685);
and U8841 (N_8841,N_5143,N_4910);
and U8842 (N_8842,N_6432,N_4473);
nor U8843 (N_8843,N_7965,N_7595);
nand U8844 (N_8844,N_6395,N_4764);
and U8845 (N_8845,N_4260,N_6773);
nor U8846 (N_8846,N_4998,N_5855);
nand U8847 (N_8847,N_7225,N_6523);
or U8848 (N_8848,N_7555,N_7256);
nor U8849 (N_8849,N_5199,N_6294);
nor U8850 (N_8850,N_7706,N_6991);
xnor U8851 (N_8851,N_7189,N_5178);
or U8852 (N_8852,N_4582,N_6181);
and U8853 (N_8853,N_5060,N_7047);
nand U8854 (N_8854,N_6911,N_6418);
xor U8855 (N_8855,N_5773,N_7134);
and U8856 (N_8856,N_5676,N_5312);
nor U8857 (N_8857,N_6254,N_5353);
and U8858 (N_8858,N_7488,N_4013);
xor U8859 (N_8859,N_6004,N_6097);
and U8860 (N_8860,N_6697,N_5873);
xor U8861 (N_8861,N_4596,N_6581);
or U8862 (N_8862,N_7315,N_5852);
or U8863 (N_8863,N_6048,N_5878);
nor U8864 (N_8864,N_4645,N_4961);
or U8865 (N_8865,N_4394,N_6116);
or U8866 (N_8866,N_4758,N_4714);
nand U8867 (N_8867,N_7086,N_4436);
xor U8868 (N_8868,N_6369,N_5877);
nand U8869 (N_8869,N_7791,N_5037);
nand U8870 (N_8870,N_6676,N_4250);
nor U8871 (N_8871,N_5706,N_6839);
and U8872 (N_8872,N_7400,N_7925);
and U8873 (N_8873,N_6712,N_6805);
and U8874 (N_8874,N_5791,N_7074);
or U8875 (N_8875,N_5381,N_6598);
nand U8876 (N_8876,N_5764,N_5568);
and U8877 (N_8877,N_5020,N_4688);
and U8878 (N_8878,N_7924,N_6497);
xnor U8879 (N_8879,N_4546,N_7001);
and U8880 (N_8880,N_5105,N_4011);
and U8881 (N_8881,N_5471,N_7740);
or U8882 (N_8882,N_4878,N_7842);
xnor U8883 (N_8883,N_4655,N_4437);
or U8884 (N_8884,N_4064,N_4871);
or U8885 (N_8885,N_6411,N_6538);
nand U8886 (N_8886,N_4353,N_5198);
nand U8887 (N_8887,N_5690,N_7747);
or U8888 (N_8888,N_7115,N_4663);
nor U8889 (N_8889,N_6954,N_6477);
xor U8890 (N_8890,N_4119,N_4451);
or U8891 (N_8891,N_7979,N_7568);
nand U8892 (N_8892,N_4027,N_6069);
and U8893 (N_8893,N_5720,N_4529);
xnor U8894 (N_8894,N_4318,N_5859);
and U8895 (N_8895,N_7097,N_6216);
xnor U8896 (N_8896,N_6575,N_4607);
xor U8897 (N_8897,N_6412,N_6476);
nor U8898 (N_8898,N_4457,N_7981);
or U8899 (N_8899,N_4941,N_4156);
or U8900 (N_8900,N_5269,N_7867);
and U8901 (N_8901,N_7336,N_6583);
and U8902 (N_8902,N_7701,N_7212);
nand U8903 (N_8903,N_4398,N_5847);
or U8904 (N_8904,N_4855,N_5653);
and U8905 (N_8905,N_5280,N_5169);
and U8906 (N_8906,N_6246,N_5401);
and U8907 (N_8907,N_7687,N_4577);
nand U8908 (N_8908,N_7664,N_6962);
nand U8909 (N_8909,N_5734,N_7306);
nor U8910 (N_8910,N_6336,N_6223);
nor U8911 (N_8911,N_5513,N_6965);
and U8912 (N_8912,N_5694,N_4492);
xor U8913 (N_8913,N_6791,N_6239);
nand U8914 (N_8914,N_4936,N_4182);
nand U8915 (N_8915,N_5134,N_7424);
or U8916 (N_8916,N_5634,N_5750);
nand U8917 (N_8917,N_6865,N_7676);
xnor U8918 (N_8918,N_4336,N_6315);
xnor U8919 (N_8919,N_7009,N_7279);
xnor U8920 (N_8920,N_7087,N_4674);
nor U8921 (N_8921,N_4681,N_6371);
nand U8922 (N_8922,N_7146,N_7730);
nand U8923 (N_8923,N_4286,N_4613);
nor U8924 (N_8924,N_6500,N_5146);
and U8925 (N_8925,N_7471,N_6356);
and U8926 (N_8926,N_4419,N_4520);
nor U8927 (N_8927,N_6059,N_6908);
or U8928 (N_8928,N_7323,N_7122);
or U8929 (N_8929,N_6225,N_5885);
nand U8930 (N_8930,N_6802,N_7779);
nor U8931 (N_8931,N_7271,N_4583);
xor U8932 (N_8932,N_6929,N_5655);
nor U8933 (N_8933,N_6361,N_4462);
nor U8934 (N_8934,N_4741,N_5052);
or U8935 (N_8935,N_4273,N_4827);
xor U8936 (N_8936,N_7777,N_6760);
nand U8937 (N_8937,N_7175,N_5736);
nor U8938 (N_8938,N_5943,N_4840);
xnor U8939 (N_8939,N_4292,N_6118);
or U8940 (N_8940,N_7649,N_7830);
nand U8941 (N_8941,N_7632,N_5980);
or U8942 (N_8942,N_5996,N_7267);
or U8943 (N_8943,N_6963,N_6382);
or U8944 (N_8944,N_4888,N_7358);
nor U8945 (N_8945,N_5801,N_4811);
nor U8946 (N_8946,N_6022,N_5671);
nor U8947 (N_8947,N_5301,N_5168);
and U8948 (N_8948,N_5092,N_7566);
nand U8949 (N_8949,N_4634,N_5017);
and U8950 (N_8950,N_7710,N_5769);
nor U8951 (N_8951,N_7907,N_7556);
nand U8952 (N_8952,N_7625,N_5768);
or U8953 (N_8953,N_5539,N_5911);
nand U8954 (N_8954,N_7887,N_7227);
and U8955 (N_8955,N_7045,N_7479);
or U8956 (N_8956,N_6930,N_4078);
and U8957 (N_8957,N_7183,N_6488);
nand U8958 (N_8958,N_7624,N_4101);
nor U8959 (N_8959,N_5516,N_4391);
and U8960 (N_8960,N_4481,N_6330);
xor U8961 (N_8961,N_7772,N_4025);
nor U8962 (N_8962,N_4397,N_7263);
xor U8963 (N_8963,N_7660,N_4953);
nand U8964 (N_8964,N_6636,N_7057);
and U8965 (N_8965,N_6178,N_4511);
nor U8966 (N_8966,N_5624,N_7216);
or U8967 (N_8967,N_7814,N_4740);
nand U8968 (N_8968,N_5566,N_6579);
nand U8969 (N_8969,N_6468,N_7679);
xnor U8970 (N_8970,N_6537,N_5836);
and U8971 (N_8971,N_7818,N_4559);
nand U8972 (N_8972,N_7491,N_5672);
and U8973 (N_8973,N_5700,N_7557);
nor U8974 (N_8974,N_5454,N_5632);
and U8975 (N_8975,N_4912,N_4146);
xor U8976 (N_8976,N_5302,N_6755);
or U8977 (N_8977,N_4621,N_6439);
nor U8978 (N_8978,N_5567,N_6453);
nand U8979 (N_8979,N_5957,N_6157);
and U8980 (N_8980,N_7127,N_4805);
nand U8981 (N_8981,N_4539,N_6654);
nor U8982 (N_8982,N_6293,N_7109);
xnor U8983 (N_8983,N_7634,N_5774);
nand U8984 (N_8984,N_4356,N_7678);
or U8985 (N_8985,N_7018,N_5876);
xor U8986 (N_8986,N_5075,N_7685);
xor U8987 (N_8987,N_6020,N_4920);
nand U8988 (N_8988,N_7639,N_7243);
xnor U8989 (N_8989,N_4750,N_6164);
nand U8990 (N_8990,N_4136,N_6608);
or U8991 (N_8991,N_5868,N_4891);
nand U8992 (N_8992,N_4813,N_5719);
xnor U8993 (N_8993,N_4703,N_7506);
or U8994 (N_8994,N_4528,N_5018);
nor U8995 (N_8995,N_6817,N_5947);
or U8996 (N_8996,N_5067,N_7703);
nand U8997 (N_8997,N_4622,N_7110);
nand U8998 (N_8998,N_7220,N_4179);
xnor U8999 (N_8999,N_7896,N_6555);
xnor U9000 (N_9000,N_7484,N_6707);
nor U9001 (N_9001,N_6879,N_5319);
or U9002 (N_9002,N_4235,N_5206);
and U9003 (N_9003,N_5850,N_6054);
nand U9004 (N_9004,N_4207,N_6421);
xor U9005 (N_9005,N_7667,N_4934);
or U9006 (N_9006,N_5991,N_5424);
nor U9007 (N_9007,N_6337,N_6008);
or U9008 (N_9008,N_6494,N_6501);
nor U9009 (N_9009,N_4364,N_6430);
or U9010 (N_9010,N_5138,N_4517);
nor U9011 (N_9011,N_4393,N_7421);
xnor U9012 (N_9012,N_7147,N_5028);
or U9013 (N_9013,N_6357,N_4970);
or U9014 (N_9014,N_7527,N_6106);
nand U9015 (N_9015,N_5203,N_7969);
and U9016 (N_9016,N_7822,N_5409);
nand U9017 (N_9017,N_5116,N_5502);
nand U9018 (N_9018,N_6590,N_7198);
nor U9019 (N_9019,N_6290,N_4382);
or U9020 (N_9020,N_6108,N_5622);
xnor U9021 (N_9021,N_5001,N_7373);
xor U9022 (N_9022,N_6721,N_7913);
and U9023 (N_9023,N_6449,N_5459);
xnor U9024 (N_9024,N_6851,N_4557);
or U9025 (N_9025,N_6601,N_6904);
nand U9026 (N_9026,N_7841,N_4787);
nor U9027 (N_9027,N_6816,N_6600);
and U9028 (N_9028,N_6552,N_7760);
or U9029 (N_9029,N_6926,N_6665);
or U9030 (N_9030,N_4461,N_5031);
nor U9031 (N_9031,N_7727,N_6747);
and U9032 (N_9032,N_4044,N_5273);
nor U9033 (N_9033,N_7090,N_5995);
nand U9034 (N_9034,N_6864,N_7584);
xnor U9035 (N_9035,N_7511,N_5440);
xor U9036 (N_9036,N_5647,N_6208);
xor U9037 (N_9037,N_6376,N_5058);
and U9038 (N_9038,N_4610,N_6471);
and U9039 (N_9039,N_5970,N_5920);
nand U9040 (N_9040,N_5391,N_7116);
or U9041 (N_9041,N_7992,N_6823);
and U9042 (N_9042,N_7300,N_6704);
nor U9043 (N_9043,N_6040,N_7827);
nand U9044 (N_9044,N_5812,N_6768);
nand U9045 (N_9045,N_4667,N_7732);
or U9046 (N_9046,N_6055,N_4174);
or U9047 (N_9047,N_5737,N_7607);
xnor U9048 (N_9048,N_5793,N_6051);
nor U9049 (N_9049,N_5816,N_4997);
or U9050 (N_9050,N_6804,N_6997);
nand U9051 (N_9051,N_6450,N_5586);
xnor U9052 (N_9052,N_6109,N_5738);
nand U9053 (N_9053,N_7052,N_4733);
or U9054 (N_9054,N_4858,N_6145);
nand U9055 (N_9055,N_5805,N_6184);
xor U9056 (N_9056,N_6889,N_5744);
nor U9057 (N_9057,N_7065,N_7062);
and U9058 (N_9058,N_5040,N_4947);
nand U9059 (N_9059,N_7517,N_5360);
or U9060 (N_9060,N_4296,N_4048);
nand U9061 (N_9061,N_6326,N_5376);
nand U9062 (N_9062,N_4896,N_4619);
xnor U9063 (N_9063,N_7990,N_5144);
nand U9064 (N_9064,N_7597,N_7276);
nand U9065 (N_9065,N_4718,N_4666);
nor U9066 (N_9066,N_6729,N_4927);
and U9067 (N_9067,N_7167,N_7794);
nor U9068 (N_9068,N_6078,N_5554);
xnor U9069 (N_9069,N_4036,N_6193);
or U9070 (N_9070,N_4075,N_5220);
xor U9071 (N_9071,N_7656,N_5219);
nand U9072 (N_9072,N_5473,N_5093);
or U9073 (N_9073,N_5534,N_6769);
nand U9074 (N_9074,N_4880,N_4226);
xnor U9075 (N_9075,N_5681,N_5063);
nand U9076 (N_9076,N_5101,N_5438);
xnor U9077 (N_9077,N_5824,N_4052);
or U9078 (N_9078,N_6036,N_7028);
xor U9079 (N_9079,N_5846,N_5606);
nor U9080 (N_9080,N_7828,N_5845);
nor U9081 (N_9081,N_6942,N_5084);
nand U9082 (N_9082,N_6101,N_7007);
xnor U9083 (N_9083,N_5732,N_7817);
nor U9084 (N_9084,N_4525,N_4285);
nor U9085 (N_9085,N_4874,N_6247);
xnor U9086 (N_9086,N_6571,N_5308);
nand U9087 (N_9087,N_5551,N_5832);
nor U9088 (N_9088,N_7986,N_4388);
and U9089 (N_9089,N_6451,N_6632);
nand U9090 (N_9090,N_6327,N_4245);
nand U9091 (N_9091,N_4507,N_4359);
nand U9092 (N_9092,N_7394,N_4775);
xor U9093 (N_9093,N_6445,N_5323);
nor U9094 (N_9094,N_4660,N_6972);
nand U9095 (N_9095,N_5201,N_5945);
and U9096 (N_9096,N_6633,N_6010);
nand U9097 (N_9097,N_7582,N_5306);
nor U9098 (N_9098,N_7917,N_6038);
nor U9099 (N_9099,N_6021,N_5214);
xnor U9100 (N_9100,N_5049,N_5879);
nor U9101 (N_9101,N_7002,N_4135);
and U9102 (N_9102,N_5973,N_7013);
and U9103 (N_9103,N_5025,N_7836);
and U9104 (N_9104,N_6550,N_7259);
and U9105 (N_9105,N_4589,N_5083);
nand U9106 (N_9106,N_4466,N_7357);
and U9107 (N_9107,N_4649,N_7786);
and U9108 (N_9108,N_7877,N_7390);
or U9109 (N_9109,N_6289,N_7528);
xnor U9110 (N_9110,N_7208,N_6614);
nor U9111 (N_9111,N_7610,N_4322);
xor U9112 (N_9112,N_7843,N_7670);
or U9113 (N_9113,N_6784,N_6975);
xnor U9114 (N_9114,N_4651,N_4784);
or U9115 (N_9115,N_6503,N_4063);
nor U9116 (N_9116,N_6117,N_5416);
nor U9117 (N_9117,N_4732,N_6144);
nand U9118 (N_9118,N_4434,N_4279);
nor U9119 (N_9119,N_5555,N_7743);
xor U9120 (N_9120,N_7459,N_6153);
nand U9121 (N_9121,N_4087,N_6849);
nand U9122 (N_9122,N_6429,N_6927);
xor U9123 (N_9123,N_5165,N_5540);
nor U9124 (N_9124,N_5226,N_5435);
or U9125 (N_9125,N_5488,N_4646);
nand U9126 (N_9126,N_4115,N_6340);
nor U9127 (N_9127,N_7789,N_5789);
xor U9128 (N_9128,N_7014,N_5243);
nand U9129 (N_9129,N_4378,N_6687);
or U9130 (N_9130,N_6562,N_5392);
xor U9131 (N_9131,N_5728,N_7156);
xnor U9132 (N_9132,N_5858,N_4976);
nand U9133 (N_9133,N_5642,N_4532);
or U9134 (N_9134,N_6134,N_5781);
xnor U9135 (N_9135,N_4337,N_6565);
and U9136 (N_9136,N_6138,N_6443);
nand U9137 (N_9137,N_5667,N_5045);
xnor U9138 (N_9138,N_6641,N_5452);
xor U9139 (N_9139,N_7652,N_7099);
xor U9140 (N_9140,N_4818,N_6304);
nor U9141 (N_9141,N_5533,N_4614);
and U9142 (N_9142,N_5066,N_7619);
and U9143 (N_9143,N_4320,N_7889);
xnor U9144 (N_9144,N_6746,N_4004);
and U9145 (N_9145,N_4484,N_6763);
and U9146 (N_9146,N_5358,N_4200);
xor U9147 (N_9147,N_6428,N_7304);
and U9148 (N_9148,N_6025,N_7448);
or U9149 (N_9149,N_4716,N_4037);
nor U9150 (N_9150,N_5161,N_4791);
and U9151 (N_9151,N_4427,N_5794);
xor U9152 (N_9152,N_7589,N_7895);
or U9153 (N_9153,N_4639,N_4611);
or U9154 (N_9154,N_5000,N_4982);
nand U9155 (N_9155,N_5448,N_4243);
nor U9156 (N_9156,N_6012,N_4861);
nor U9157 (N_9157,N_4006,N_4046);
nand U9158 (N_9158,N_6692,N_6698);
xnor U9159 (N_9159,N_7588,N_7288);
and U9160 (N_9160,N_7046,N_5708);
xnor U9161 (N_9161,N_7258,N_6306);
nor U9162 (N_9162,N_7605,N_5543);
nor U9163 (N_9163,N_4514,N_5466);
or U9164 (N_9164,N_5916,N_5574);
xor U9165 (N_9165,N_4588,N_6070);
xnor U9166 (N_9166,N_5380,N_6505);
nand U9167 (N_9167,N_4809,N_7980);
xor U9168 (N_9168,N_6824,N_4148);
and U9169 (N_9169,N_5387,N_4362);
nand U9170 (N_9170,N_4313,N_6273);
xnor U9171 (N_9171,N_6259,N_4186);
xnor U9172 (N_9172,N_5385,N_6172);
xnor U9173 (N_9173,N_5158,N_4726);
nand U9174 (N_9174,N_5425,N_4083);
xor U9175 (N_9175,N_4705,N_7966);
and U9176 (N_9176,N_6525,N_6985);
or U9177 (N_9177,N_7958,N_6609);
or U9178 (N_9178,N_6493,N_4432);
xnor U9179 (N_9179,N_4502,N_6531);
and U9180 (N_9180,N_4120,N_4711);
or U9181 (N_9181,N_6673,N_7103);
and U9182 (N_9182,N_4505,N_4496);
or U9183 (N_9183,N_6295,N_7292);
nor U9184 (N_9184,N_6955,N_5745);
and U9185 (N_9185,N_4178,N_4734);
and U9186 (N_9186,N_5133,N_4995);
or U9187 (N_9187,N_4903,N_4266);
xnor U9188 (N_9188,N_7173,N_5241);
or U9189 (N_9189,N_5740,N_6177);
or U9190 (N_9190,N_5450,N_6063);
xor U9191 (N_9191,N_5515,N_6792);
xnor U9192 (N_9192,N_4082,N_5021);
nor U9193 (N_9193,N_4648,N_5297);
nor U9194 (N_9194,N_7698,N_4977);
xnor U9195 (N_9195,N_4282,N_5331);
nand U9196 (N_9196,N_7247,N_5461);
or U9197 (N_9197,N_4558,N_5091);
or U9198 (N_9198,N_4803,N_7994);
or U9199 (N_9199,N_7509,N_4617);
and U9200 (N_9200,N_7839,N_7043);
and U9201 (N_9201,N_6961,N_5470);
or U9202 (N_9202,N_5303,N_7197);
nor U9203 (N_9203,N_4745,N_4014);
nor U9204 (N_9204,N_6885,N_5608);
or U9205 (N_9205,N_5402,N_4738);
or U9206 (N_9206,N_4916,N_4856);
or U9207 (N_9207,N_6716,N_5577);
nand U9208 (N_9208,N_4127,N_6683);
nor U9209 (N_9209,N_4405,N_4251);
nor U9210 (N_9210,N_6329,N_5089);
nand U9211 (N_9211,N_6674,N_4743);
xor U9212 (N_9212,N_6414,N_7416);
nor U9213 (N_9213,N_6814,N_7541);
or U9214 (N_9214,N_4404,N_5518);
and U9215 (N_9215,N_7503,N_4220);
nand U9216 (N_9216,N_4668,N_4628);
xnor U9217 (N_9217,N_5307,N_4210);
xnor U9218 (N_9218,N_4425,N_5934);
or U9219 (N_9219,N_6454,N_5537);
nand U9220 (N_9220,N_5660,N_5315);
and U9221 (N_9221,N_4054,N_6173);
and U9222 (N_9222,N_5908,N_7266);
nor U9223 (N_9223,N_6730,N_4247);
xor U9224 (N_9224,N_5351,N_4712);
xnor U9225 (N_9225,N_4379,N_4118);
nand U9226 (N_9226,N_4094,N_7700);
or U9227 (N_9227,N_6682,N_7427);
nand U9228 (N_9228,N_6068,N_7805);
nor U9229 (N_9229,N_4485,N_5571);
and U9230 (N_9230,N_5717,N_7618);
nor U9231 (N_9231,N_7193,N_7111);
nand U9232 (N_9232,N_7581,N_6964);
nor U9233 (N_9233,N_5953,N_5895);
xnor U9234 (N_9234,N_5839,N_6083);
and U9235 (N_9235,N_4125,N_5616);
or U9236 (N_9236,N_6152,N_5125);
nand U9237 (N_9237,N_4760,N_6332);
xnor U9238 (N_9238,N_6837,N_6520);
and U9239 (N_9239,N_5987,N_5019);
xnor U9240 (N_9240,N_5504,N_7128);
xor U9241 (N_9241,N_6409,N_4691);
nand U9242 (N_9242,N_4230,N_6789);
nand U9243 (N_9243,N_5325,N_5702);
nor U9244 (N_9244,N_7879,N_4002);
nor U9245 (N_9245,N_4350,N_6815);
nor U9246 (N_9246,N_4786,N_7800);
xnor U9247 (N_9247,N_6016,N_5192);
or U9248 (N_9248,N_6436,N_7297);
xor U9249 (N_9249,N_6474,N_7178);
or U9250 (N_9250,N_6742,N_6028);
xnor U9251 (N_9251,N_4568,N_7172);
nand U9252 (N_9252,N_7403,N_7257);
or U9253 (N_9253,N_6843,N_4673);
nand U9254 (N_9254,N_5154,N_7019);
and U9255 (N_9255,N_6586,N_5486);
nor U9256 (N_9256,N_7552,N_5840);
or U9257 (N_9257,N_7768,N_4991);
xor U9258 (N_9258,N_4277,N_5506);
or U9259 (N_9259,N_4632,N_5636);
nand U9260 (N_9260,N_6597,N_6924);
and U9261 (N_9261,N_7029,N_6858);
nand U9262 (N_9262,N_7321,N_5726);
and U9263 (N_9263,N_4928,N_7792);
nand U9264 (N_9264,N_4612,N_5500);
and U9265 (N_9265,N_5906,N_4365);
nand U9266 (N_9266,N_7550,N_4727);
nand U9267 (N_9267,N_4021,N_6896);
nor U9268 (N_9268,N_4556,N_7406);
xor U9269 (N_9269,N_6240,N_5604);
nand U9270 (N_9270,N_4267,N_7285);
or U9271 (N_9271,N_6209,N_6532);
nor U9272 (N_9272,N_6321,N_5333);
or U9273 (N_9273,N_7250,N_6176);
nor U9274 (N_9274,N_6510,N_7505);
nor U9275 (N_9275,N_5536,N_5964);
or U9276 (N_9276,N_5935,N_7811);
nor U9277 (N_9277,N_6498,N_6605);
nand U9278 (N_9278,N_6480,N_6221);
nor U9279 (N_9279,N_6404,N_4693);
nor U9280 (N_9280,N_4349,N_5334);
or U9281 (N_9281,N_4905,N_7025);
xnor U9282 (N_9282,N_4624,N_7184);
xor U9283 (N_9283,N_5552,N_7960);
or U9284 (N_9284,N_4931,N_7516);
xor U9285 (N_9285,N_6853,N_4675);
nand U9286 (N_9286,N_4513,N_7117);
or U9287 (N_9287,N_7987,N_4949);
nor U9288 (N_9288,N_4574,N_5721);
or U9289 (N_9289,N_4926,N_4854);
xnor U9290 (N_9290,N_4325,N_7371);
or U9291 (N_9291,N_6484,N_5107);
xor U9292 (N_9292,N_6475,N_5645);
xor U9293 (N_9293,N_4548,N_6518);
nand U9294 (N_9294,N_5718,N_6649);
nor U9295 (N_9295,N_6092,N_4475);
and U9296 (N_9296,N_5857,N_4924);
nor U9297 (N_9297,N_6270,N_4184);
nand U9298 (N_9298,N_4183,N_7058);
nor U9299 (N_9299,N_5492,N_4785);
xor U9300 (N_9300,N_4154,N_5494);
or U9301 (N_9301,N_4595,N_6877);
xnor U9302 (N_9302,N_7334,N_7211);
xnor U9303 (N_9303,N_7327,N_7808);
xnor U9304 (N_9304,N_6339,N_7813);
nor U9305 (N_9305,N_7493,N_4527);
or U9306 (N_9306,N_6867,N_4761);
nand U9307 (N_9307,N_7027,N_7388);
nand U9308 (N_9308,N_7989,N_4489);
nor U9309 (N_9309,N_6772,N_5861);
nor U9310 (N_9310,N_4301,N_4477);
or U9311 (N_9311,N_5444,N_6095);
or U9312 (N_9312,N_7314,N_4549);
or U9313 (N_9313,N_4993,N_6102);
and U9314 (N_9314,N_7356,N_7094);
and U9315 (N_9315,N_5530,N_6751);
xor U9316 (N_9316,N_4755,N_4423);
or U9317 (N_9317,N_4409,N_5013);
nand U9318 (N_9318,N_6213,N_5788);
nor U9319 (N_9319,N_5162,N_5123);
and U9320 (N_9320,N_5182,N_5268);
xnor U9321 (N_9321,N_4033,N_4387);
xnor U9322 (N_9322,N_7280,N_4943);
nor U9323 (N_9323,N_5639,N_6034);
or U9324 (N_9324,N_6932,N_5797);
xnor U9325 (N_9325,N_4635,N_6093);
xnor U9326 (N_9326,N_4215,N_6130);
xor U9327 (N_9327,N_4019,N_7688);
xnor U9328 (N_9328,N_4665,N_7983);
xor U9329 (N_9329,N_7860,N_5320);
nor U9330 (N_9330,N_7601,N_4351);
or U9331 (N_9331,N_4591,N_4772);
nand U9332 (N_9332,N_6263,N_4899);
nand U9333 (N_9333,N_4782,N_4807);
xor U9334 (N_9334,N_4032,N_5340);
xnor U9335 (N_9335,N_5224,N_5748);
nor U9336 (N_9336,N_5474,N_6818);
xor U9337 (N_9337,N_7104,N_7269);
nand U9338 (N_9338,N_7475,N_5096);
nand U9339 (N_9339,N_6272,N_6363);
and U9340 (N_9340,N_6978,N_6934);
nor U9341 (N_9341,N_7934,N_4777);
nor U9342 (N_9342,N_4034,N_5363);
and U9343 (N_9343,N_6622,N_5965);
and U9344 (N_9344,N_6685,N_6307);
nor U9345 (N_9345,N_5656,N_5629);
nand U9346 (N_9346,N_4307,N_4312);
or U9347 (N_9347,N_4294,N_6949);
or U9348 (N_9348,N_5564,N_7408);
or U9349 (N_9349,N_7486,N_4447);
xor U9350 (N_9350,N_5081,N_5752);
nand U9351 (N_9351,N_4788,N_6688);
and U9352 (N_9352,N_4401,N_6080);
or U9353 (N_9353,N_5372,N_4535);
nand U9354 (N_9354,N_4342,N_4848);
or U9355 (N_9355,N_7764,N_4795);
and U9356 (N_9356,N_7565,N_7657);
and U9357 (N_9357,N_5896,N_6783);
nor U9358 (N_9358,N_4824,N_7745);
or U9359 (N_9359,N_7684,N_6928);
nor U9360 (N_9360,N_5465,N_5324);
and U9361 (N_9361,N_7340,N_7439);
or U9362 (N_9362,N_6139,N_5607);
xor U9363 (N_9363,N_4699,N_7443);
nand U9364 (N_9364,N_4850,N_7152);
and U9365 (N_9365,N_5563,N_5682);
or U9366 (N_9366,N_4985,N_4290);
nor U9367 (N_9367,N_6809,N_5085);
nand U9368 (N_9368,N_6367,N_5347);
xnor U9369 (N_9369,N_5428,N_5170);
or U9370 (N_9370,N_5202,N_6014);
xor U9371 (N_9371,N_5004,N_6611);
or U9372 (N_9372,N_6267,N_6569);
or U9373 (N_9373,N_7489,N_5352);
nand U9374 (N_9374,N_4662,N_4792);
xor U9375 (N_9375,N_4526,N_6405);
nand U9376 (N_9376,N_4630,N_6467);
xor U9377 (N_9377,N_4092,N_5410);
nand U9378 (N_9378,N_5611,N_5437);
xor U9379 (N_9379,N_4429,N_6690);
nand U9380 (N_9380,N_4530,N_7284);
nand U9381 (N_9381,N_5511,N_4159);
nand U9382 (N_9382,N_7642,N_5270);
or U9383 (N_9383,N_4580,N_5600);
or U9384 (N_9384,N_6835,N_4177);
xor U9385 (N_9385,N_7337,N_4205);
xnor U9386 (N_9386,N_5591,N_7899);
nand U9387 (N_9387,N_6180,N_7105);
or U9388 (N_9388,N_4093,N_6165);
nand U9389 (N_9389,N_6778,N_5106);
nand U9390 (N_9390,N_6913,N_6242);
nand U9391 (N_9391,N_6241,N_6277);
nor U9392 (N_9392,N_7264,N_5390);
nand U9393 (N_9393,N_7663,N_5368);
and U9394 (N_9394,N_5684,N_6170);
or U9395 (N_9395,N_5262,N_6140);
xnor U9396 (N_9396,N_6894,N_7032);
or U9397 (N_9397,N_7095,N_6308);
nor U9398 (N_9398,N_6124,N_5405);
nor U9399 (N_9399,N_6743,N_4846);
nand U9400 (N_9400,N_6725,N_4001);
and U9401 (N_9401,N_7067,N_5357);
nor U9402 (N_9402,N_5570,N_7951);
nor U9403 (N_9403,N_7851,N_5854);
xor U9404 (N_9404,N_7793,N_5984);
or U9405 (N_9405,N_7662,N_6871);
nor U9406 (N_9406,N_4175,N_6160);
nand U9407 (N_9407,N_4367,N_5236);
xor U9408 (N_9408,N_5374,N_7691);
xor U9409 (N_9409,N_5585,N_6995);
and U9410 (N_9410,N_5287,N_7920);
xnor U9411 (N_9411,N_5223,N_5881);
and U9412 (N_9412,N_7748,N_5275);
and U9413 (N_9413,N_6906,N_6542);
and U9414 (N_9414,N_7628,N_6741);
nor U9415 (N_9415,N_7347,N_5557);
and U9416 (N_9416,N_6419,N_6129);
or U9417 (N_9417,N_5207,N_7778);
and U9418 (N_9418,N_7399,N_7533);
nand U9419 (N_9419,N_5393,N_7423);
xnor U9420 (N_9420,N_4698,N_5281);
or U9421 (N_9421,N_7240,N_6621);
and U9422 (N_9422,N_5579,N_6076);
nand U9423 (N_9423,N_4493,N_5580);
xnor U9424 (N_9424,N_6167,N_7031);
nand U9425 (N_9425,N_6447,N_7395);
nand U9426 (N_9426,N_7638,N_4834);
and U9427 (N_9427,N_7495,N_4754);
or U9428 (N_9428,N_5061,N_4042);
xor U9429 (N_9429,N_4066,N_4242);
or U9430 (N_9430,N_6833,N_4898);
nor U9431 (N_9431,N_7487,N_4859);
nor U9432 (N_9432,N_4051,N_6325);
and U9433 (N_9433,N_4626,N_6067);
xor U9434 (N_9434,N_7837,N_5602);
nor U9435 (N_9435,N_5648,N_4506);
or U9436 (N_9436,N_7857,N_4570);
xor U9437 (N_9437,N_7774,N_5171);
nor U9438 (N_9438,N_6800,N_7346);
xnor U9439 (N_9439,N_5086,N_5619);
xor U9440 (N_9440,N_7932,N_7361);
xor U9441 (N_9441,N_7339,N_6220);
nor U9442 (N_9442,N_5451,N_7414);
xnor U9443 (N_9443,N_4225,N_4500);
or U9444 (N_9444,N_5547,N_5111);
nand U9445 (N_9445,N_5069,N_5147);
or U9446 (N_9446,N_5359,N_7718);
or U9447 (N_9447,N_5819,N_7051);
xor U9448 (N_9448,N_5900,N_6892);
nor U9449 (N_9449,N_4233,N_5572);
nor U9450 (N_9450,N_6860,N_4171);
nor U9451 (N_9451,N_7504,N_7040);
xnor U9452 (N_9452,N_6884,N_6424);
nand U9453 (N_9453,N_5265,N_7341);
and U9454 (N_9454,N_5871,N_7496);
and U9455 (N_9455,N_7329,N_5497);
and U9456 (N_9456,N_6870,N_6749);
nor U9457 (N_9457,N_6120,N_4357);
and U9458 (N_9458,N_5149,N_6499);
or U9459 (N_9459,N_7036,N_6335);
nand U9460 (N_9460,N_6483,N_4793);
nor U9461 (N_9461,N_6224,N_4005);
nand U9462 (N_9462,N_6379,N_4138);
nand U9463 (N_9463,N_6155,N_5345);
and U9464 (N_9464,N_4341,N_4480);
xor U9465 (N_9465,N_6941,N_6299);
nand U9466 (N_9466,N_4636,N_4190);
nor U9467 (N_9467,N_6744,N_6465);
xor U9468 (N_9468,N_4917,N_5842);
or U9469 (N_9469,N_6023,N_5256);
or U9470 (N_9470,N_6996,N_6486);
nor U9471 (N_9471,N_5771,N_6638);
or U9472 (N_9472,N_4224,N_6448);
xor U9473 (N_9473,N_4460,N_4114);
and U9474 (N_9474,N_6533,N_4843);
and U9475 (N_9475,N_6718,N_6875);
xor U9476 (N_9476,N_5828,N_5955);
and U9477 (N_9477,N_5799,N_4332);
and U9478 (N_9478,N_7819,N_5724);
and U9479 (N_9479,N_5917,N_5620);
or U9480 (N_9480,N_4155,N_6580);
xnor U9481 (N_9481,N_7988,N_6190);
and U9482 (N_9482,N_7695,N_4952);
nand U9483 (N_9483,N_5240,N_4124);
nand U9484 (N_9484,N_5630,N_6062);
nand U9485 (N_9485,N_6516,N_5238);
and U9486 (N_9486,N_5767,N_7080);
xor U9487 (N_9487,N_7833,N_5388);
or U9488 (N_9488,N_7906,N_7738);
xor U9489 (N_9489,N_5963,N_7538);
or U9490 (N_9490,N_7661,N_6786);
xnor U9491 (N_9491,N_6374,N_6740);
nor U9492 (N_9492,N_6061,N_6105);
xor U9493 (N_9493,N_7354,N_4722);
xnor U9494 (N_9494,N_4830,N_6988);
or U9495 (N_9495,N_6918,N_4638);
nand U9496 (N_9496,N_4747,N_7163);
or U9497 (N_9497,N_6282,N_4531);
xnor U9498 (N_9498,N_5522,N_6599);
and U9499 (N_9499,N_6115,N_4550);
nor U9500 (N_9500,N_4061,N_5640);
and U9501 (N_9501,N_7752,N_5503);
xnor U9502 (N_9502,N_4585,N_5163);
nand U9503 (N_9503,N_4731,N_7299);
xnor U9504 (N_9504,N_5260,N_6380);
xnor U9505 (N_9505,N_7187,N_4298);
or U9506 (N_9506,N_4956,N_5300);
xor U9507 (N_9507,N_7967,N_7693);
nor U9508 (N_9508,N_6619,N_7948);
or U9509 (N_9509,N_6857,N_7838);
nor U9510 (N_9510,N_4049,N_6686);
nand U9511 (N_9511,N_6485,N_7283);
and U9512 (N_9512,N_7615,N_5541);
nor U9513 (N_9513,N_7468,N_7270);
xnor U9514 (N_9514,N_4565,N_7549);
nor U9515 (N_9515,N_7066,N_5155);
or U9516 (N_9516,N_4814,N_4164);
nor U9517 (N_9517,N_7702,N_4677);
nor U9518 (N_9518,N_6779,N_5441);
or U9519 (N_9519,N_6281,N_6974);
and U9520 (N_9520,N_5419,N_7071);
nand U9521 (N_9521,N_7301,N_4442);
or U9522 (N_9522,N_7260,N_5596);
nand U9523 (N_9523,N_5833,N_5962);
xor U9524 (N_9524,N_7548,N_5944);
and U9525 (N_9525,N_6035,N_5239);
and U9526 (N_9526,N_5743,N_7871);
xnor U9527 (N_9527,N_6013,N_7530);
and U9528 (N_9528,N_5336,N_7755);
nand U9529 (N_9529,N_5489,N_4272);
or U9530 (N_9530,N_6968,N_6710);
or U9531 (N_9531,N_4562,N_6775);
nor U9532 (N_9532,N_4625,N_7174);
nor U9533 (N_9533,N_6970,N_4031);
or U9534 (N_9534,N_6211,N_7254);
or U9535 (N_9535,N_7575,N_4835);
nand U9536 (N_9536,N_5064,N_4109);
nor U9537 (N_9537,N_6987,N_7215);
xnor U9538 (N_9538,N_4449,N_6098);
nand U9539 (N_9539,N_5705,N_4326);
and U9540 (N_9540,N_4223,N_6037);
and U9541 (N_9541,N_4259,N_6976);
nor U9542 (N_9542,N_6808,N_4647);
or U9543 (N_9543,N_4488,N_7559);
xnor U9544 (N_9544,N_5355,N_5856);
nor U9545 (N_9545,N_6195,N_6842);
nor U9546 (N_9546,N_7984,N_6215);
and U9547 (N_9547,N_5121,N_6847);
and U9548 (N_9548,N_7210,N_6734);
and U9549 (N_9549,N_7790,N_4151);
nor U9550 (N_9550,N_5946,N_5338);
nand U9551 (N_9551,N_5562,N_5821);
and U9552 (N_9552,N_7017,N_7381);
nand U9553 (N_9553,N_4214,N_5675);
xor U9554 (N_9554,N_6347,N_5749);
xor U9555 (N_9555,N_4980,N_4544);
or U9556 (N_9556,N_4416,N_5102);
nor U9557 (N_9557,N_6680,N_6905);
xor U9558 (N_9558,N_4056,N_7908);
or U9559 (N_9559,N_4327,N_7223);
or U9560 (N_9560,N_7962,N_4345);
nor U9561 (N_9561,N_6075,N_7635);
and U9562 (N_9562,N_6206,N_6207);
xnor U9563 (N_9563,N_6123,N_4540);
or U9564 (N_9564,N_6390,N_5704);
or U9565 (N_9565,N_4412,N_7332);
nand U9566 (N_9566,N_6322,N_7959);
or U9567 (N_9567,N_7949,N_6856);
nand U9568 (N_9568,N_4686,N_7004);
and U9569 (N_9569,N_6191,N_4757);
or U9570 (N_9570,N_6634,N_6629);
xnor U9571 (N_9571,N_7079,N_4735);
xnor U9572 (N_9572,N_6344,N_4450);
nand U9573 (N_9573,N_5723,N_6648);
nor U9574 (N_9574,N_4911,N_7677);
nor U9575 (N_9575,N_4020,N_4088);
nor U9576 (N_9576,N_5923,N_7554);
and U9577 (N_9577,N_7586,N_6852);
or U9578 (N_9578,N_7235,N_4311);
nand U9579 (N_9579,N_4832,N_5689);
nor U9580 (N_9580,N_6990,N_4141);
nor U9581 (N_9581,N_4140,N_7072);
and U9582 (N_9582,N_4960,N_7166);
xor U9583 (N_9583,N_5892,N_4265);
nand U9584 (N_9584,N_6642,N_6661);
nand U9585 (N_9585,N_4709,N_4347);
nor U9586 (N_9586,N_4901,N_4862);
or U9587 (N_9587,N_7612,N_6891);
xnor U9588 (N_9588,N_5860,N_7985);
xor U9589 (N_9589,N_5509,N_5244);
or U9590 (N_9590,N_6081,N_4494);
nor U9591 (N_9591,N_6394,N_7737);
or U9592 (N_9592,N_5289,N_4908);
nand U9593 (N_9593,N_7402,N_6576);
xnor U9594 (N_9594,N_5775,N_7909);
nand U9595 (N_9595,N_7914,N_5560);
nand U9596 (N_9596,N_7020,N_5722);
nand U9597 (N_9597,N_7199,N_4800);
and U9598 (N_9598,N_4608,N_4555);
nor U9599 (N_9599,N_4133,N_7091);
and U9600 (N_9600,N_5901,N_7766);
xnor U9601 (N_9601,N_6201,N_5119);
xor U9602 (N_9602,N_5986,N_6044);
or U9603 (N_9603,N_4599,N_5071);
and U9604 (N_9604,N_7419,N_6163);
and U9605 (N_9605,N_6009,N_6268);
and U9606 (N_9606,N_4143,N_4395);
nand U9607 (N_9607,N_6050,N_5587);
nor U9608 (N_9608,N_6993,N_4264);
nor U9609 (N_9609,N_6049,N_5145);
nand U9610 (N_9610,N_4355,N_7840);
and U9611 (N_9611,N_7574,N_5770);
nor U9612 (N_9612,N_4454,N_5924);
and U9613 (N_9613,N_7918,N_5778);
or U9614 (N_9614,N_7742,N_4055);
xnor U9615 (N_9615,N_7275,N_7185);
or U9616 (N_9616,N_6862,N_5940);
or U9617 (N_9617,N_5371,N_4067);
and U9618 (N_9618,N_7717,N_6994);
nand U9619 (N_9619,N_5584,N_6141);
nand U9620 (N_9620,N_4694,N_5837);
nand U9621 (N_9621,N_7246,N_5597);
nand U9622 (N_9622,N_5532,N_7081);
or U9623 (N_9623,N_7500,N_7551);
or U9624 (N_9624,N_4678,N_4131);
or U9625 (N_9625,N_6577,N_7100);
xor U9626 (N_9626,N_4192,N_5941);
or U9627 (N_9627,N_4464,N_6733);
xnor U9628 (N_9628,N_6933,N_6983);
or U9629 (N_9629,N_7937,N_6567);
nand U9630 (N_9630,N_4030,N_5787);
nor U9631 (N_9631,N_4212,N_7325);
or U9632 (N_9632,N_5482,N_6463);
xnor U9633 (N_9633,N_7756,N_7519);
and U9634 (N_9634,N_7590,N_7132);
nor U9635 (N_9635,N_5621,N_6348);
or U9636 (N_9636,N_5348,N_6352);
nor U9637 (N_9637,N_5313,N_6052);
or U9638 (N_9638,N_5827,N_5030);
and U9639 (N_9639,N_7993,N_4816);
and U9640 (N_9640,N_7526,N_7797);
nand U9641 (N_9641,N_4410,N_4334);
nand U9642 (N_9642,N_6553,N_4701);
nor U9643 (N_9643,N_4969,N_5299);
nor U9644 (N_9644,N_5252,N_5822);
xor U9645 (N_9645,N_4571,N_4167);
xnor U9646 (N_9646,N_4193,N_6761);
xor U9647 (N_9647,N_4938,N_5618);
nor U9648 (N_9648,N_6812,N_7176);
nor U9649 (N_9649,N_6417,N_6219);
xnor U9650 (N_9650,N_4994,N_7780);
nand U9651 (N_9651,N_4222,N_6456);
and U9652 (N_9652,N_5544,N_5751);
and U9653 (N_9653,N_5994,N_4990);
nor U9654 (N_9654,N_7428,N_5520);
or U9655 (N_9655,N_5795,N_6001);
nand U9656 (N_9656,N_6212,N_7177);
nor U9657 (N_9657,N_4249,N_6850);
nor U9658 (N_9658,N_6956,N_5959);
nor U9659 (N_9659,N_4208,N_4708);
nor U9660 (N_9660,N_6717,N_5032);
nor U9661 (N_9661,N_7968,N_5929);
nand U9662 (N_9662,N_7378,N_6732);
nor U9663 (N_9663,N_4620,N_6514);
nor U9664 (N_9664,N_7902,N_5305);
xor U9665 (N_9665,N_7916,N_4590);
nand U9666 (N_9666,N_5763,N_6402);
or U9667 (N_9667,N_5670,N_4498);
or U9668 (N_9668,N_4872,N_6345);
or U9669 (N_9669,N_7849,N_5933);
and U9670 (N_9670,N_7370,N_4305);
or U9671 (N_9671,N_4828,N_6046);
or U9672 (N_9672,N_4554,N_6543);
xor U9673 (N_9673,N_5696,N_4163);
nor U9674 (N_9674,N_5730,N_7648);
or U9675 (N_9675,N_7807,N_5350);
and U9676 (N_9676,N_5164,N_4719);
and U9677 (N_9677,N_4868,N_6782);
nand U9678 (N_9678,N_7482,N_4196);
xnor U9679 (N_9679,N_5181,N_6757);
xor U9680 (N_9680,N_5977,N_5098);
or U9681 (N_9681,N_7942,N_4739);
nor U9682 (N_9682,N_7991,N_5573);
nor U9683 (N_9683,N_7407,N_4518);
xor U9684 (N_9684,N_6612,N_4490);
nand U9685 (N_9685,N_5230,N_6785);
xor U9686 (N_9686,N_6094,N_6630);
and U9687 (N_9687,N_4057,N_5400);
nor U9688 (N_9688,N_5731,N_4915);
or U9689 (N_9689,N_4989,N_5701);
nand U9690 (N_9690,N_5129,N_5664);
and U9691 (N_9691,N_6566,N_5266);
nor U9692 (N_9692,N_7502,N_4833);
or U9693 (N_9693,N_6033,N_6620);
xor U9694 (N_9694,N_4281,N_4826);
nand U9695 (N_9695,N_7604,N_6073);
or U9696 (N_9696,N_7953,N_5818);
or U9697 (N_9697,N_5999,N_6420);
and U9698 (N_9698,N_7855,N_6526);
nand U9699 (N_9699,N_5191,N_5646);
nor U9700 (N_9700,N_4172,N_7380);
nand U9701 (N_9701,N_7722,N_6548);
and U9702 (N_9702,N_6715,N_6162);
and U9703 (N_9703,N_4509,N_5212);
nand U9704 (N_9704,N_4697,N_5804);
nand U9705 (N_9705,N_7287,N_6652);
or U9706 (N_9706,N_6595,N_6301);
xnor U9707 (N_9707,N_7470,N_4769);
and U9708 (N_9708,N_5468,N_6952);
or U9709 (N_9709,N_5447,N_7846);
nand U9710 (N_9710,N_5978,N_5928);
xor U9711 (N_9711,N_5869,N_6205);
xnor U9712 (N_9712,N_4268,N_4344);
nor U9713 (N_9713,N_6481,N_6132);
xor U9714 (N_9714,N_7112,N_6489);
xnor U9715 (N_9715,N_4640,N_4050);
nor U9716 (N_9716,N_7956,N_5507);
or U9717 (N_9717,N_5432,N_4852);
or U9718 (N_9718,N_7869,N_5197);
and U9719 (N_9719,N_6058,N_7705);
nor U9720 (N_9720,N_4602,N_6148);
nand U9721 (N_9721,N_7224,N_4288);
xor U9722 (N_9722,N_7826,N_7835);
or U9723 (N_9723,N_5142,N_5531);
nand U9724 (N_9724,N_4074,N_4819);
nor U9725 (N_9725,N_7120,N_7750);
and U9726 (N_9726,N_6845,N_5692);
or U9727 (N_9727,N_6647,N_7317);
nor U9728 (N_9728,N_6103,N_5968);
or U9729 (N_9729,N_4870,N_4059);
nand U9730 (N_9730,N_4892,N_7149);
or U9731 (N_9731,N_5074,N_4501);
xor U9732 (N_9732,N_5038,N_6529);
nor U9733 (N_9733,N_4077,N_5053);
or U9734 (N_9734,N_6502,N_6944);
nor U9735 (N_9735,N_6524,N_7349);
nand U9736 (N_9736,N_7873,N_7931);
nor U9737 (N_9737,N_7481,N_5160);
xnor U9738 (N_9738,N_7715,N_4413);
xor U9739 (N_9739,N_4152,N_5641);
xnor U9740 (N_9740,N_7343,N_5467);
nand U9741 (N_9741,N_7008,N_6110);
xnor U9742 (N_9742,N_7154,N_6551);
xor U9743 (N_9743,N_6472,N_7219);
nand U9744 (N_9744,N_5525,N_7903);
nand U9745 (N_9745,N_5546,N_6397);
nand U9746 (N_9746,N_7763,N_7383);
or U9747 (N_9747,N_4304,N_4358);
xor U9748 (N_9748,N_7494,N_7897);
xnor U9749 (N_9749,N_6056,N_7121);
and U9750 (N_9750,N_5903,N_5367);
or U9751 (N_9751,N_7454,N_5126);
nor U9752 (N_9752,N_7950,N_5370);
nand U9753 (N_9753,N_4106,N_5411);
and U9754 (N_9754,N_6440,N_7658);
nor U9755 (N_9755,N_7823,N_6257);
nand U9756 (N_9756,N_7077,N_4000);
nand U9757 (N_9757,N_4730,N_4123);
nor U9758 (N_9758,N_7351,N_6558);
and U9759 (N_9759,N_5399,N_5112);
xor U9760 (N_9760,N_6018,N_7191);
nand U9761 (N_9761,N_5759,N_7665);
nand U9762 (N_9762,N_4256,N_7982);
nor U9763 (N_9763,N_5529,N_4576);
nor U9764 (N_9764,N_6150,N_4895);
nor U9765 (N_9765,N_5414,N_4478);
nor U9766 (N_9766,N_6827,N_4145);
and U9767 (N_9767,N_4366,N_4426);
and U9768 (N_9768,N_6196,N_5041);
or U9769 (N_9769,N_6806,N_6066);
nor U9770 (N_9770,N_5043,N_6624);
nor U9771 (N_9771,N_7546,N_4339);
nor U9772 (N_9772,N_4962,N_6719);
xnor U9773 (N_9773,N_6198,N_7076);
or U9774 (N_9774,N_6260,N_5806);
or U9775 (N_9775,N_7641,N_7245);
or U9776 (N_9776,N_6278,N_7497);
nor U9777 (N_9777,N_4375,N_4418);
xnor U9778 (N_9778,N_6528,N_6006);
xnor U9779 (N_9779,N_7947,N_7059);
nand U9780 (N_9780,N_7543,N_7928);
nor U9781 (N_9781,N_7529,N_4289);
xnor U9782 (N_9782,N_5898,N_7450);
or U9783 (N_9783,N_6236,N_5221);
nor U9784 (N_9784,N_5613,N_6943);
and U9785 (N_9785,N_7545,N_4360);
or U9786 (N_9786,N_6280,N_7696);
nand U9787 (N_9787,N_7438,N_7039);
xnor U9788 (N_9788,N_4860,N_6794);
xnor U9789 (N_9789,N_7580,N_6143);
and U9790 (N_9790,N_6807,N_4122);
nor U9791 (N_9791,N_7171,N_5809);
nand U9792 (N_9792,N_4902,N_5073);
xnor U9793 (N_9793,N_5918,N_6112);
and U9794 (N_9794,N_7736,N_6393);
or U9795 (N_9795,N_7338,N_6596);
xnor U9796 (N_9796,N_4633,N_4471);
xnor U9797 (N_9797,N_7102,N_7603);
nand U9798 (N_9798,N_4696,N_4263);
xnor U9799 (N_9799,N_7714,N_7692);
or U9800 (N_9800,N_6276,N_7409);
and U9801 (N_9801,N_6291,N_4408);
nor U9802 (N_9802,N_7868,N_4203);
nand U9803 (N_9803,N_7157,N_4165);
nand U9804 (N_9804,N_6723,N_4971);
nand U9805 (N_9805,N_4766,N_4616);
nor U9806 (N_9806,N_4415,N_6535);
nor U9807 (N_9807,N_4219,N_7290);
and U9808 (N_9808,N_4104,N_7485);
nand U9809 (N_9809,N_5960,N_5746);
nor U9810 (N_9810,N_5843,N_5902);
xnor U9811 (N_9811,N_6408,N_5687);
or U9812 (N_9812,N_7644,N_7282);
xor U9813 (N_9813,N_5699,N_6720);
nor U9814 (N_9814,N_6111,N_7600);
or U9815 (N_9815,N_7938,N_4026);
and U9816 (N_9816,N_5501,N_5033);
or U9817 (N_9817,N_6457,N_6951);
and U9818 (N_9818,N_7922,N_6748);
nor U9819 (N_9819,N_5330,N_4081);
and U9820 (N_9820,N_5979,N_5807);
nand U9821 (N_9821,N_5364,N_5899);
xor U9822 (N_9822,N_4420,N_5802);
and U9823 (N_9823,N_5741,N_7107);
and U9824 (N_9824,N_7598,N_5711);
or U9825 (N_9825,N_4781,N_4060);
xnor U9826 (N_9826,N_4315,N_6245);
or U9827 (N_9827,N_5485,N_6825);
nand U9828 (N_9828,N_4796,N_5418);
nor U9829 (N_9829,N_5625,N_4725);
nor U9830 (N_9830,N_5356,N_7041);
and U9831 (N_9831,N_6826,N_7536);
or U9832 (N_9832,N_6708,N_6878);
or U9833 (N_9833,N_4309,N_6670);
xnor U9834 (N_9834,N_5022,N_6863);
nor U9835 (N_9835,N_4604,N_7026);
and U9836 (N_9836,N_6999,N_5285);
xnor U9837 (N_9837,N_7713,N_5527);
nand U9838 (N_9838,N_4236,N_6973);
nand U9839 (N_9839,N_4508,N_4443);
and U9840 (N_9840,N_4851,N_6168);
and U9841 (N_9841,N_4967,N_7478);
nor U9842 (N_9842,N_6655,N_7145);
or U9843 (N_9843,N_4653,N_5714);
or U9844 (N_9844,N_5335,N_6256);
nor U9845 (N_9845,N_5510,N_6283);
nor U9846 (N_9846,N_7108,N_4921);
nand U9847 (N_9847,N_7944,N_5894);
nand U9848 (N_9848,N_5863,N_6666);
xor U9849 (N_9849,N_4821,N_4202);
or U9850 (N_9850,N_6156,N_6663);
or U9851 (N_9851,N_6300,N_5872);
and U9852 (N_9852,N_5661,N_5760);
nand U9853 (N_9853,N_7585,N_6365);
nand U9854 (N_9854,N_5375,N_5131);
or U9855 (N_9855,N_6072,N_5950);
nand U9856 (N_9856,N_4097,N_4280);
nand U9857 (N_9857,N_5135,N_5626);
nand U9858 (N_9858,N_5194,N_6939);
nand U9859 (N_9859,N_5167,N_4586);
nor U9860 (N_9860,N_5590,N_7238);
nand U9861 (N_9861,N_5588,N_4672);
nand U9862 (N_9862,N_6114,N_5462);
nor U9863 (N_9863,N_4996,N_6231);
or U9864 (N_9864,N_6696,N_7093);
and U9865 (N_9865,N_7614,N_6971);
xor U9866 (N_9866,N_7767,N_4894);
xor U9867 (N_9867,N_7309,N_4433);
and U9868 (N_9868,N_5956,N_6606);
nor U9869 (N_9869,N_7578,N_6910);
and U9870 (N_9870,N_6512,N_6086);
nor U9871 (N_9871,N_4940,N_4206);
nand U9872 (N_9872,N_4252,N_5186);
nor U9873 (N_9873,N_7681,N_5549);
nor U9874 (N_9874,N_6570,N_5691);
xor U9875 (N_9875,N_5505,N_6881);
nand U9876 (N_9876,N_7733,N_7312);
nor U9877 (N_9877,N_6401,N_6626);
nand U9878 (N_9878,N_5848,N_7063);
and U9879 (N_9879,N_4257,N_4853);
nor U9880 (N_9880,N_5196,N_5150);
nor U9881 (N_9881,N_4542,N_5975);
and U9882 (N_9882,N_7393,N_4669);
nor U9883 (N_9883,N_5070,N_4913);
or U9884 (N_9884,N_6194,N_6872);
or U9885 (N_9885,N_6848,N_7118);
and U9886 (N_9886,N_4244,N_4128);
nor U9887 (N_9887,N_7033,N_7874);
or U9888 (N_9888,N_5772,N_7561);
xnor U9889 (N_9889,N_7866,N_6368);
nor U9890 (N_9890,N_7856,N_4476);
and U9891 (N_9891,N_4319,N_6639);
or U9892 (N_9892,N_5665,N_5969);
nor U9893 (N_9893,N_6210,N_7142);
and U9894 (N_9894,N_4065,N_5250);
nand U9895 (N_9895,N_5893,N_7795);
and U9896 (N_9896,N_4965,N_6305);
nand U9897 (N_9897,N_4255,N_7277);
and U9898 (N_9898,N_7372,N_6572);
xor U9899 (N_9899,N_4096,N_6615);
or U9900 (N_9900,N_6706,N_7921);
or U9901 (N_9901,N_4130,N_4543);
nor U9902 (N_9902,N_7348,N_6750);
nor U9903 (N_9903,N_7451,N_4831);
nor U9904 (N_9904,N_7125,N_7006);
xnor U9905 (N_9905,N_6495,N_6341);
nor U9906 (N_9906,N_7005,N_6890);
nand U9907 (N_9907,N_6406,N_5495);
or U9908 (N_9908,N_4237,N_7741);
and U9909 (N_9909,N_7435,N_7444);
and U9910 (N_9910,N_4717,N_4773);
nand U9911 (N_9911,N_6318,N_6705);
or U9912 (N_9912,N_5508,N_7515);
nand U9913 (N_9913,N_7398,N_4499);
nor U9914 (N_9914,N_5346,N_6915);
or U9915 (N_9915,N_7576,N_5951);
xnor U9916 (N_9916,N_5815,N_7456);
and U9917 (N_9917,N_5090,N_5077);
and U9918 (N_9918,N_5891,N_5404);
or U9919 (N_9919,N_6838,N_6840);
nor U9920 (N_9920,N_5047,N_6701);
nand U9921 (N_9921,N_6640,N_4121);
xnor U9922 (N_9922,N_5668,N_4058);
or U9923 (N_9923,N_7038,N_6074);
or U9924 (N_9924,N_7915,N_7523);
nand U9925 (N_9925,N_6602,N_7796);
or U9926 (N_9926,N_6912,N_6400);
nor U9927 (N_9927,N_4340,N_5072);
nand U9928 (N_9928,N_7539,N_5930);
nand U9929 (N_9929,N_7563,N_4973);
or U9930 (N_9930,N_5727,N_7483);
nand U9931 (N_9931,N_7458,N_5594);
xor U9932 (N_9932,N_6534,N_6780);
or U9933 (N_9933,N_7449,N_6714);
or U9934 (N_9934,N_5811,N_6227);
xor U9935 (N_9935,N_7569,N_5245);
xor U9936 (N_9936,N_4495,N_5343);
or U9937 (N_9937,N_5329,N_4381);
or U9938 (N_9938,N_6829,N_5851);
nand U9939 (N_9939,N_6947,N_5436);
nand U9940 (N_9940,N_7474,N_7140);
xnor U9941 (N_9941,N_7168,N_4482);
xnor U9942 (N_9942,N_5222,N_7558);
or U9943 (N_9943,N_7686,N_7136);
nand U9944 (N_9944,N_6396,N_6900);
nand U9945 (N_9945,N_4783,N_5193);
nor U9946 (N_9946,N_6935,N_4884);
nand U9947 (N_9947,N_6854,N_7073);
or U9948 (N_9948,N_4817,N_4804);
or U9949 (N_9949,N_6218,N_4472);
xor U9950 (N_9950,N_4035,N_7675);
xnor U9951 (N_9951,N_7261,N_7192);
nand U9952 (N_9952,N_6869,N_4652);
nand U9953 (N_9953,N_7627,N_5210);
nand U9954 (N_9954,N_7522,N_6279);
xor U9955 (N_9955,N_4169,N_4806);
nand U9956 (N_9956,N_6989,N_6482);
and U9957 (N_9957,N_4710,N_5036);
xnor U9958 (N_9958,N_7761,N_4922);
or U9959 (N_9959,N_4615,N_6813);
and U9960 (N_9960,N_4329,N_4836);
or U9961 (N_9961,N_4774,N_4933);
nand U9962 (N_9962,N_6907,N_7064);
or U9963 (N_9963,N_7901,N_6603);
nor U9964 (N_9964,N_5972,N_6203);
and U9965 (N_9965,N_4091,N_4069);
nor U9966 (N_9966,N_7248,N_6423);
and U9967 (N_9967,N_7431,N_7218);
xor U9968 (N_9968,N_4144,N_5698);
xor U9969 (N_9969,N_4411,N_6317);
nor U9970 (N_9970,N_4369,N_7385);
xnor U9971 (N_9971,N_6298,N_6426);
xor U9972 (N_9972,N_5023,N_7694);
xnor U9973 (N_9973,N_6324,N_6261);
or U9974 (N_9974,N_4293,N_7620);
and U9975 (N_9975,N_5478,N_6616);
nand U9976 (N_9976,N_7744,N_4893);
nand U9977 (N_9977,N_5825,N_4541);
nor U9978 (N_9978,N_7935,N_7864);
nor U9979 (N_9979,N_4676,N_4180);
nor U9980 (N_9980,N_7998,N_5761);
nand U9981 (N_9981,N_7137,N_7940);
nor U9982 (N_9982,N_6727,N_5652);
nor U9983 (N_9983,N_5377,N_5882);
nor U9984 (N_9984,N_4890,N_5295);
nor U9985 (N_9985,N_7234,N_5396);
xnor U9986 (N_9986,N_7881,N_5605);
and U9987 (N_9987,N_7296,N_6689);
nand U9988 (N_9988,N_6628,N_7249);
xor U9989 (N_9989,N_5628,N_4564);
and U9990 (N_9990,N_7637,N_4198);
nor U9991 (N_9991,N_6517,N_7200);
nand U9992 (N_9992,N_6728,N_5599);
xnor U9993 (N_9993,N_6945,N_7853);
or U9994 (N_9994,N_4453,N_6466);
nand U9995 (N_9995,N_4865,N_5615);
nand U9996 (N_9996,N_6310,N_7606);
or U9997 (N_9997,N_6731,N_5633);
nor U9998 (N_9998,N_5453,N_5813);
xnor U9999 (N_9999,N_4695,N_7891);
and U10000 (N_10000,N_7881,N_5883);
nand U10001 (N_10001,N_4846,N_4388);
xnor U10002 (N_10002,N_7980,N_6575);
nand U10003 (N_10003,N_7367,N_4277);
and U10004 (N_10004,N_4618,N_6131);
nand U10005 (N_10005,N_4202,N_6481);
or U10006 (N_10006,N_5843,N_4640);
nand U10007 (N_10007,N_4347,N_7932);
or U10008 (N_10008,N_4834,N_5159);
nor U10009 (N_10009,N_7611,N_6942);
or U10010 (N_10010,N_5806,N_4824);
nor U10011 (N_10011,N_6141,N_4820);
xor U10012 (N_10012,N_4572,N_5209);
and U10013 (N_10013,N_7493,N_6503);
nor U10014 (N_10014,N_7784,N_7749);
and U10015 (N_10015,N_5111,N_5487);
xor U10016 (N_10016,N_4909,N_4963);
nand U10017 (N_10017,N_6148,N_4435);
and U10018 (N_10018,N_7846,N_6393);
or U10019 (N_10019,N_5555,N_5789);
nand U10020 (N_10020,N_6704,N_4562);
or U10021 (N_10021,N_7023,N_4038);
and U10022 (N_10022,N_6934,N_6332);
or U10023 (N_10023,N_7777,N_5831);
or U10024 (N_10024,N_4168,N_7387);
nor U10025 (N_10025,N_5966,N_5524);
and U10026 (N_10026,N_7267,N_7564);
nand U10027 (N_10027,N_5431,N_5922);
nand U10028 (N_10028,N_4338,N_6476);
nand U10029 (N_10029,N_5014,N_4000);
or U10030 (N_10030,N_5559,N_6566);
and U10031 (N_10031,N_5847,N_4645);
or U10032 (N_10032,N_5927,N_4142);
nand U10033 (N_10033,N_7225,N_6743);
nor U10034 (N_10034,N_6128,N_7652);
or U10035 (N_10035,N_4888,N_6295);
and U10036 (N_10036,N_4952,N_6648);
xnor U10037 (N_10037,N_4484,N_6365);
or U10038 (N_10038,N_4815,N_5528);
nor U10039 (N_10039,N_5465,N_6040);
or U10040 (N_10040,N_5831,N_5663);
nor U10041 (N_10041,N_5583,N_4003);
nand U10042 (N_10042,N_6287,N_6105);
and U10043 (N_10043,N_6532,N_4048);
nor U10044 (N_10044,N_7644,N_7972);
nand U10045 (N_10045,N_4005,N_7938);
xnor U10046 (N_10046,N_4935,N_6478);
nand U10047 (N_10047,N_4298,N_5350);
nor U10048 (N_10048,N_4662,N_5428);
and U10049 (N_10049,N_7603,N_7859);
xor U10050 (N_10050,N_6239,N_5631);
nor U10051 (N_10051,N_6351,N_4129);
xnor U10052 (N_10052,N_5570,N_4834);
xor U10053 (N_10053,N_6182,N_7231);
nor U10054 (N_10054,N_5027,N_4203);
xnor U10055 (N_10055,N_5908,N_5964);
or U10056 (N_10056,N_4015,N_5240);
and U10057 (N_10057,N_7127,N_7754);
xor U10058 (N_10058,N_6267,N_5144);
xor U10059 (N_10059,N_5676,N_4194);
nand U10060 (N_10060,N_6947,N_5633);
nand U10061 (N_10061,N_7063,N_5958);
nand U10062 (N_10062,N_5472,N_4479);
nor U10063 (N_10063,N_6952,N_4764);
xnor U10064 (N_10064,N_4090,N_5813);
or U10065 (N_10065,N_7867,N_6175);
nand U10066 (N_10066,N_7509,N_5690);
xor U10067 (N_10067,N_5306,N_6886);
xor U10068 (N_10068,N_6820,N_6028);
nand U10069 (N_10069,N_4172,N_5531);
and U10070 (N_10070,N_5385,N_6780);
nand U10071 (N_10071,N_4401,N_7272);
nand U10072 (N_10072,N_7730,N_5688);
and U10073 (N_10073,N_5945,N_6649);
or U10074 (N_10074,N_4192,N_4322);
nor U10075 (N_10075,N_4937,N_7994);
or U10076 (N_10076,N_5730,N_7045);
nand U10077 (N_10077,N_6858,N_4995);
and U10078 (N_10078,N_4383,N_5437);
nand U10079 (N_10079,N_7753,N_6607);
xor U10080 (N_10080,N_4055,N_6756);
or U10081 (N_10081,N_5379,N_4446);
nand U10082 (N_10082,N_6406,N_6540);
nand U10083 (N_10083,N_7829,N_7392);
xor U10084 (N_10084,N_5237,N_4184);
nand U10085 (N_10085,N_5280,N_7666);
nor U10086 (N_10086,N_6332,N_5551);
or U10087 (N_10087,N_6111,N_4270);
xnor U10088 (N_10088,N_4582,N_6071);
xor U10089 (N_10089,N_6725,N_5957);
or U10090 (N_10090,N_5431,N_4889);
xnor U10091 (N_10091,N_4782,N_7115);
and U10092 (N_10092,N_7973,N_4775);
or U10093 (N_10093,N_5529,N_5333);
and U10094 (N_10094,N_7611,N_4020);
nand U10095 (N_10095,N_5951,N_7409);
xnor U10096 (N_10096,N_6032,N_4442);
xor U10097 (N_10097,N_5086,N_6789);
nor U10098 (N_10098,N_6716,N_7413);
and U10099 (N_10099,N_7072,N_7849);
nand U10100 (N_10100,N_7521,N_7388);
nand U10101 (N_10101,N_7012,N_5832);
xnor U10102 (N_10102,N_5233,N_7764);
and U10103 (N_10103,N_4131,N_6989);
nor U10104 (N_10104,N_7405,N_7479);
nor U10105 (N_10105,N_4336,N_4964);
xor U10106 (N_10106,N_5981,N_7555);
or U10107 (N_10107,N_4054,N_5636);
or U10108 (N_10108,N_7036,N_6836);
and U10109 (N_10109,N_4024,N_7743);
xnor U10110 (N_10110,N_5601,N_6399);
and U10111 (N_10111,N_5700,N_4978);
nand U10112 (N_10112,N_5820,N_6266);
nand U10113 (N_10113,N_5045,N_4856);
nand U10114 (N_10114,N_4924,N_6867);
and U10115 (N_10115,N_6898,N_6825);
or U10116 (N_10116,N_4117,N_7792);
and U10117 (N_10117,N_5643,N_6843);
xnor U10118 (N_10118,N_5152,N_6415);
nor U10119 (N_10119,N_4900,N_4456);
and U10120 (N_10120,N_5065,N_5278);
or U10121 (N_10121,N_6134,N_7401);
nand U10122 (N_10122,N_4381,N_6321);
nand U10123 (N_10123,N_4323,N_4147);
xor U10124 (N_10124,N_4710,N_5872);
or U10125 (N_10125,N_7050,N_6229);
and U10126 (N_10126,N_5677,N_6184);
or U10127 (N_10127,N_5574,N_7852);
and U10128 (N_10128,N_5708,N_5238);
or U10129 (N_10129,N_7633,N_4575);
nand U10130 (N_10130,N_7069,N_7537);
nand U10131 (N_10131,N_4940,N_4885);
and U10132 (N_10132,N_7215,N_5396);
nor U10133 (N_10133,N_4231,N_6015);
and U10134 (N_10134,N_5630,N_7540);
or U10135 (N_10135,N_4863,N_7658);
nor U10136 (N_10136,N_6260,N_4583);
xor U10137 (N_10137,N_4073,N_4993);
and U10138 (N_10138,N_4431,N_4734);
nor U10139 (N_10139,N_4005,N_6987);
or U10140 (N_10140,N_5281,N_4257);
or U10141 (N_10141,N_4282,N_6200);
or U10142 (N_10142,N_4162,N_5729);
or U10143 (N_10143,N_4762,N_5846);
and U10144 (N_10144,N_5268,N_6586);
or U10145 (N_10145,N_7788,N_5542);
nor U10146 (N_10146,N_6471,N_5384);
nor U10147 (N_10147,N_7289,N_4777);
and U10148 (N_10148,N_6904,N_7945);
or U10149 (N_10149,N_5489,N_6368);
nand U10150 (N_10150,N_7515,N_7699);
nor U10151 (N_10151,N_5620,N_7574);
and U10152 (N_10152,N_7228,N_5978);
nor U10153 (N_10153,N_5129,N_6717);
and U10154 (N_10154,N_5012,N_5347);
or U10155 (N_10155,N_4219,N_5129);
nand U10156 (N_10156,N_5216,N_4319);
and U10157 (N_10157,N_4025,N_7137);
xnor U10158 (N_10158,N_7041,N_7557);
or U10159 (N_10159,N_4359,N_4724);
or U10160 (N_10160,N_4650,N_7205);
and U10161 (N_10161,N_4389,N_4977);
and U10162 (N_10162,N_5237,N_4515);
xor U10163 (N_10163,N_4932,N_7344);
nand U10164 (N_10164,N_7590,N_6786);
nand U10165 (N_10165,N_5620,N_5228);
nand U10166 (N_10166,N_4650,N_7772);
nor U10167 (N_10167,N_4868,N_5400);
or U10168 (N_10168,N_5227,N_7786);
or U10169 (N_10169,N_6410,N_5562);
or U10170 (N_10170,N_4790,N_5790);
or U10171 (N_10171,N_6757,N_5371);
or U10172 (N_10172,N_5800,N_4597);
or U10173 (N_10173,N_7987,N_7686);
or U10174 (N_10174,N_6154,N_4816);
nand U10175 (N_10175,N_4139,N_6171);
nor U10176 (N_10176,N_5364,N_7008);
and U10177 (N_10177,N_5381,N_6704);
nand U10178 (N_10178,N_6832,N_6261);
xor U10179 (N_10179,N_7888,N_7819);
nand U10180 (N_10180,N_4536,N_7884);
nand U10181 (N_10181,N_6276,N_5596);
nor U10182 (N_10182,N_7822,N_5561);
or U10183 (N_10183,N_6456,N_6979);
nor U10184 (N_10184,N_7817,N_6591);
nand U10185 (N_10185,N_4882,N_5209);
nand U10186 (N_10186,N_4635,N_4006);
nand U10187 (N_10187,N_6121,N_6543);
nand U10188 (N_10188,N_7687,N_7725);
nand U10189 (N_10189,N_5339,N_6861);
nand U10190 (N_10190,N_6156,N_5727);
nand U10191 (N_10191,N_7270,N_5810);
nand U10192 (N_10192,N_7796,N_5887);
and U10193 (N_10193,N_6147,N_6932);
nor U10194 (N_10194,N_7150,N_7451);
and U10195 (N_10195,N_5829,N_7406);
or U10196 (N_10196,N_7088,N_4024);
or U10197 (N_10197,N_4842,N_5128);
or U10198 (N_10198,N_7503,N_5192);
nor U10199 (N_10199,N_6357,N_4211);
nor U10200 (N_10200,N_6699,N_4403);
or U10201 (N_10201,N_4478,N_4752);
nand U10202 (N_10202,N_6970,N_4351);
xnor U10203 (N_10203,N_4686,N_7347);
nand U10204 (N_10204,N_5893,N_6531);
xor U10205 (N_10205,N_6401,N_7176);
nand U10206 (N_10206,N_5770,N_6243);
nand U10207 (N_10207,N_7599,N_5268);
nand U10208 (N_10208,N_6306,N_7161);
or U10209 (N_10209,N_7198,N_4062);
or U10210 (N_10210,N_6588,N_7916);
xor U10211 (N_10211,N_5846,N_4796);
or U10212 (N_10212,N_4691,N_5913);
or U10213 (N_10213,N_7858,N_4101);
nor U10214 (N_10214,N_4661,N_6856);
nand U10215 (N_10215,N_4293,N_5020);
nand U10216 (N_10216,N_7970,N_7464);
nor U10217 (N_10217,N_7305,N_5862);
nor U10218 (N_10218,N_6605,N_7758);
nand U10219 (N_10219,N_5362,N_6791);
xnor U10220 (N_10220,N_4315,N_7208);
xor U10221 (N_10221,N_6059,N_4141);
or U10222 (N_10222,N_5252,N_5310);
or U10223 (N_10223,N_5045,N_6456);
xor U10224 (N_10224,N_7373,N_6946);
and U10225 (N_10225,N_7928,N_6529);
and U10226 (N_10226,N_4327,N_5165);
and U10227 (N_10227,N_5494,N_4964);
xor U10228 (N_10228,N_6757,N_6368);
nand U10229 (N_10229,N_6720,N_5859);
and U10230 (N_10230,N_7495,N_6099);
nand U10231 (N_10231,N_6544,N_5127);
xor U10232 (N_10232,N_6870,N_6701);
or U10233 (N_10233,N_5077,N_4878);
or U10234 (N_10234,N_5218,N_5723);
and U10235 (N_10235,N_4290,N_7530);
nand U10236 (N_10236,N_4831,N_7170);
xnor U10237 (N_10237,N_4516,N_4974);
nand U10238 (N_10238,N_5107,N_6149);
or U10239 (N_10239,N_7107,N_4529);
nor U10240 (N_10240,N_5102,N_5925);
xnor U10241 (N_10241,N_6576,N_4343);
or U10242 (N_10242,N_4473,N_4410);
nor U10243 (N_10243,N_6615,N_5071);
or U10244 (N_10244,N_7020,N_7011);
xor U10245 (N_10245,N_4991,N_7770);
xor U10246 (N_10246,N_6291,N_5251);
xor U10247 (N_10247,N_5005,N_5462);
and U10248 (N_10248,N_4109,N_6553);
nor U10249 (N_10249,N_4913,N_4884);
nand U10250 (N_10250,N_4329,N_6008);
nor U10251 (N_10251,N_6064,N_7173);
or U10252 (N_10252,N_5664,N_7904);
nor U10253 (N_10253,N_4558,N_7713);
xnor U10254 (N_10254,N_6103,N_4769);
and U10255 (N_10255,N_4944,N_6273);
and U10256 (N_10256,N_5367,N_5793);
nand U10257 (N_10257,N_5470,N_5905);
nor U10258 (N_10258,N_6673,N_6136);
xor U10259 (N_10259,N_6068,N_5335);
nand U10260 (N_10260,N_6160,N_5229);
xnor U10261 (N_10261,N_7628,N_5545);
nand U10262 (N_10262,N_5496,N_4990);
nand U10263 (N_10263,N_5542,N_6075);
nand U10264 (N_10264,N_5142,N_7405);
nor U10265 (N_10265,N_6643,N_6687);
nand U10266 (N_10266,N_7083,N_7480);
nor U10267 (N_10267,N_5479,N_7648);
or U10268 (N_10268,N_6995,N_7042);
or U10269 (N_10269,N_4691,N_6379);
or U10270 (N_10270,N_7461,N_7434);
and U10271 (N_10271,N_7975,N_5787);
nand U10272 (N_10272,N_4752,N_6890);
nor U10273 (N_10273,N_7658,N_6462);
nand U10274 (N_10274,N_7457,N_7025);
or U10275 (N_10275,N_7108,N_7889);
xor U10276 (N_10276,N_7880,N_5911);
xnor U10277 (N_10277,N_5129,N_6000);
or U10278 (N_10278,N_6530,N_4423);
xor U10279 (N_10279,N_5947,N_6306);
nor U10280 (N_10280,N_6724,N_6729);
nand U10281 (N_10281,N_7484,N_4736);
or U10282 (N_10282,N_6075,N_5534);
nand U10283 (N_10283,N_5311,N_4598);
nor U10284 (N_10284,N_5863,N_5336);
xor U10285 (N_10285,N_5088,N_4261);
nand U10286 (N_10286,N_6184,N_6896);
and U10287 (N_10287,N_4585,N_5445);
xnor U10288 (N_10288,N_7304,N_5904);
nor U10289 (N_10289,N_7888,N_5553);
and U10290 (N_10290,N_6052,N_6227);
and U10291 (N_10291,N_5515,N_7319);
nand U10292 (N_10292,N_6193,N_6319);
xor U10293 (N_10293,N_7539,N_7123);
nand U10294 (N_10294,N_4239,N_7623);
nor U10295 (N_10295,N_6935,N_6704);
and U10296 (N_10296,N_7080,N_6993);
xor U10297 (N_10297,N_7301,N_6488);
nand U10298 (N_10298,N_6423,N_7501);
or U10299 (N_10299,N_5100,N_6885);
nand U10300 (N_10300,N_6145,N_5754);
or U10301 (N_10301,N_5784,N_4264);
nor U10302 (N_10302,N_5534,N_5723);
nor U10303 (N_10303,N_5032,N_7691);
or U10304 (N_10304,N_7801,N_5893);
and U10305 (N_10305,N_5537,N_6412);
nor U10306 (N_10306,N_5433,N_4114);
and U10307 (N_10307,N_7589,N_6734);
nor U10308 (N_10308,N_7786,N_6364);
or U10309 (N_10309,N_4114,N_6886);
nand U10310 (N_10310,N_4256,N_5840);
and U10311 (N_10311,N_6599,N_6600);
nor U10312 (N_10312,N_6128,N_5651);
or U10313 (N_10313,N_5585,N_5256);
nand U10314 (N_10314,N_6086,N_7710);
nor U10315 (N_10315,N_4769,N_5877);
or U10316 (N_10316,N_5065,N_4862);
nand U10317 (N_10317,N_5397,N_4378);
nor U10318 (N_10318,N_6919,N_5822);
or U10319 (N_10319,N_5956,N_5547);
or U10320 (N_10320,N_6715,N_7625);
nand U10321 (N_10321,N_4239,N_4186);
xnor U10322 (N_10322,N_4781,N_6479);
xor U10323 (N_10323,N_5868,N_4253);
nor U10324 (N_10324,N_5201,N_4690);
nand U10325 (N_10325,N_4480,N_6861);
nand U10326 (N_10326,N_6054,N_6874);
xor U10327 (N_10327,N_4646,N_5802);
nor U10328 (N_10328,N_4931,N_6743);
nor U10329 (N_10329,N_4109,N_6092);
or U10330 (N_10330,N_4663,N_5995);
or U10331 (N_10331,N_4141,N_7137);
xor U10332 (N_10332,N_6120,N_6404);
nor U10333 (N_10333,N_5018,N_4367);
or U10334 (N_10334,N_5413,N_6675);
or U10335 (N_10335,N_6807,N_6862);
xnor U10336 (N_10336,N_5137,N_7856);
nand U10337 (N_10337,N_7858,N_5117);
nand U10338 (N_10338,N_4587,N_5887);
xor U10339 (N_10339,N_6748,N_6433);
xor U10340 (N_10340,N_5816,N_7528);
nor U10341 (N_10341,N_4138,N_4698);
nor U10342 (N_10342,N_7001,N_4975);
nand U10343 (N_10343,N_7511,N_5137);
or U10344 (N_10344,N_6093,N_4392);
or U10345 (N_10345,N_7119,N_4323);
and U10346 (N_10346,N_5810,N_6690);
or U10347 (N_10347,N_6504,N_7544);
nor U10348 (N_10348,N_7565,N_4078);
and U10349 (N_10349,N_7721,N_4722);
or U10350 (N_10350,N_5340,N_5867);
or U10351 (N_10351,N_5734,N_4232);
or U10352 (N_10352,N_4367,N_6794);
xor U10353 (N_10353,N_5523,N_6940);
and U10354 (N_10354,N_7161,N_4969);
or U10355 (N_10355,N_5507,N_6531);
and U10356 (N_10356,N_4588,N_7371);
nor U10357 (N_10357,N_5686,N_6685);
xor U10358 (N_10358,N_5597,N_4911);
nand U10359 (N_10359,N_6350,N_5170);
and U10360 (N_10360,N_7709,N_7450);
and U10361 (N_10361,N_7336,N_7333);
or U10362 (N_10362,N_7621,N_6500);
xnor U10363 (N_10363,N_6075,N_6716);
nor U10364 (N_10364,N_6746,N_6829);
and U10365 (N_10365,N_5024,N_5610);
nand U10366 (N_10366,N_7131,N_4570);
or U10367 (N_10367,N_5775,N_4180);
xor U10368 (N_10368,N_6438,N_7130);
nand U10369 (N_10369,N_5590,N_7449);
or U10370 (N_10370,N_6314,N_5108);
nand U10371 (N_10371,N_5596,N_6424);
xor U10372 (N_10372,N_4055,N_5193);
nor U10373 (N_10373,N_5941,N_7507);
xor U10374 (N_10374,N_5827,N_7947);
nor U10375 (N_10375,N_7576,N_7734);
xnor U10376 (N_10376,N_5714,N_7231);
xor U10377 (N_10377,N_4866,N_4262);
nor U10378 (N_10378,N_5008,N_5809);
xnor U10379 (N_10379,N_7369,N_6946);
nand U10380 (N_10380,N_5866,N_4454);
xor U10381 (N_10381,N_4079,N_6859);
nand U10382 (N_10382,N_7978,N_5818);
xnor U10383 (N_10383,N_7770,N_5673);
or U10384 (N_10384,N_6985,N_7344);
or U10385 (N_10385,N_7071,N_4386);
xor U10386 (N_10386,N_7749,N_4118);
nor U10387 (N_10387,N_5392,N_4880);
xnor U10388 (N_10388,N_6735,N_6910);
xnor U10389 (N_10389,N_7874,N_6451);
and U10390 (N_10390,N_7330,N_6970);
or U10391 (N_10391,N_5819,N_4612);
xnor U10392 (N_10392,N_5935,N_5037);
xor U10393 (N_10393,N_6127,N_4720);
xnor U10394 (N_10394,N_4580,N_7156);
xnor U10395 (N_10395,N_6238,N_6849);
xor U10396 (N_10396,N_6026,N_7693);
xnor U10397 (N_10397,N_6513,N_7144);
nor U10398 (N_10398,N_4812,N_5977);
nand U10399 (N_10399,N_5686,N_6993);
nand U10400 (N_10400,N_5258,N_7975);
xnor U10401 (N_10401,N_7237,N_6969);
or U10402 (N_10402,N_7082,N_6326);
xor U10403 (N_10403,N_4646,N_6556);
or U10404 (N_10404,N_5610,N_5553);
and U10405 (N_10405,N_5077,N_5296);
or U10406 (N_10406,N_7476,N_6428);
or U10407 (N_10407,N_7749,N_5122);
and U10408 (N_10408,N_7027,N_5787);
nand U10409 (N_10409,N_6787,N_4444);
nor U10410 (N_10410,N_6456,N_4529);
nor U10411 (N_10411,N_4085,N_5676);
and U10412 (N_10412,N_6366,N_7396);
xor U10413 (N_10413,N_6408,N_5168);
and U10414 (N_10414,N_4109,N_6146);
nor U10415 (N_10415,N_5921,N_4220);
nand U10416 (N_10416,N_4533,N_5179);
or U10417 (N_10417,N_6261,N_7165);
or U10418 (N_10418,N_4669,N_4689);
nand U10419 (N_10419,N_6680,N_4796);
nand U10420 (N_10420,N_6913,N_4671);
and U10421 (N_10421,N_4334,N_6937);
xnor U10422 (N_10422,N_4069,N_6952);
or U10423 (N_10423,N_5696,N_7054);
or U10424 (N_10424,N_4122,N_4524);
and U10425 (N_10425,N_7855,N_6613);
and U10426 (N_10426,N_6744,N_4416);
or U10427 (N_10427,N_4411,N_5524);
nand U10428 (N_10428,N_4295,N_6683);
nand U10429 (N_10429,N_4560,N_4151);
or U10430 (N_10430,N_5214,N_4210);
nor U10431 (N_10431,N_4045,N_6033);
and U10432 (N_10432,N_4700,N_5042);
xnor U10433 (N_10433,N_5755,N_7636);
xor U10434 (N_10434,N_4704,N_7867);
nand U10435 (N_10435,N_7568,N_5071);
nor U10436 (N_10436,N_4593,N_6756);
nor U10437 (N_10437,N_6670,N_6943);
or U10438 (N_10438,N_6072,N_7394);
and U10439 (N_10439,N_5427,N_7772);
nor U10440 (N_10440,N_7995,N_7270);
xor U10441 (N_10441,N_7691,N_6677);
nor U10442 (N_10442,N_4541,N_4686);
and U10443 (N_10443,N_4196,N_7907);
or U10444 (N_10444,N_4138,N_6576);
xnor U10445 (N_10445,N_7452,N_7315);
and U10446 (N_10446,N_6819,N_5300);
nor U10447 (N_10447,N_6085,N_6710);
nor U10448 (N_10448,N_4443,N_6279);
xnor U10449 (N_10449,N_7622,N_6038);
xor U10450 (N_10450,N_7558,N_7608);
xor U10451 (N_10451,N_4225,N_4389);
or U10452 (N_10452,N_4034,N_6945);
xnor U10453 (N_10453,N_6731,N_7855);
nor U10454 (N_10454,N_4319,N_6234);
nor U10455 (N_10455,N_6671,N_6835);
nand U10456 (N_10456,N_7541,N_6050);
nand U10457 (N_10457,N_6276,N_4505);
or U10458 (N_10458,N_5132,N_4689);
and U10459 (N_10459,N_6431,N_6458);
or U10460 (N_10460,N_5732,N_7907);
nor U10461 (N_10461,N_7312,N_5506);
nor U10462 (N_10462,N_5885,N_4644);
or U10463 (N_10463,N_7479,N_7349);
or U10464 (N_10464,N_5061,N_6586);
nor U10465 (N_10465,N_5097,N_5595);
xor U10466 (N_10466,N_5941,N_5886);
nor U10467 (N_10467,N_4428,N_6787);
nor U10468 (N_10468,N_7663,N_5195);
and U10469 (N_10469,N_5557,N_6091);
xor U10470 (N_10470,N_6550,N_5695);
nand U10471 (N_10471,N_6245,N_4884);
nand U10472 (N_10472,N_6479,N_4647);
nand U10473 (N_10473,N_6351,N_7714);
nand U10474 (N_10474,N_4922,N_4601);
nor U10475 (N_10475,N_6777,N_4709);
and U10476 (N_10476,N_7534,N_7735);
or U10477 (N_10477,N_5280,N_6714);
nor U10478 (N_10478,N_6802,N_5304);
xor U10479 (N_10479,N_5243,N_6090);
and U10480 (N_10480,N_4245,N_7532);
xor U10481 (N_10481,N_7323,N_5354);
and U10482 (N_10482,N_4367,N_5889);
and U10483 (N_10483,N_5317,N_4683);
and U10484 (N_10484,N_5002,N_4203);
nor U10485 (N_10485,N_6154,N_5395);
or U10486 (N_10486,N_5125,N_6164);
nor U10487 (N_10487,N_6726,N_4784);
or U10488 (N_10488,N_4475,N_5642);
nor U10489 (N_10489,N_5325,N_6726);
and U10490 (N_10490,N_7552,N_7096);
or U10491 (N_10491,N_5542,N_4202);
nor U10492 (N_10492,N_4286,N_4141);
and U10493 (N_10493,N_6103,N_5145);
or U10494 (N_10494,N_5372,N_6708);
or U10495 (N_10495,N_4011,N_4106);
nand U10496 (N_10496,N_5121,N_4856);
nand U10497 (N_10497,N_6549,N_7589);
or U10498 (N_10498,N_6368,N_4780);
nor U10499 (N_10499,N_5628,N_7067);
or U10500 (N_10500,N_7217,N_6613);
nor U10501 (N_10501,N_4163,N_7819);
or U10502 (N_10502,N_7910,N_7428);
and U10503 (N_10503,N_6481,N_7666);
xor U10504 (N_10504,N_5049,N_5930);
or U10505 (N_10505,N_5678,N_5900);
or U10506 (N_10506,N_6532,N_4086);
and U10507 (N_10507,N_4113,N_7507);
nand U10508 (N_10508,N_5492,N_6067);
nand U10509 (N_10509,N_4834,N_7398);
or U10510 (N_10510,N_7666,N_7750);
xnor U10511 (N_10511,N_7157,N_5371);
or U10512 (N_10512,N_4975,N_4604);
nor U10513 (N_10513,N_5082,N_4715);
or U10514 (N_10514,N_4878,N_4459);
nor U10515 (N_10515,N_4650,N_7350);
xnor U10516 (N_10516,N_4580,N_7952);
or U10517 (N_10517,N_6563,N_7362);
xor U10518 (N_10518,N_4060,N_7354);
nor U10519 (N_10519,N_7579,N_4880);
nor U10520 (N_10520,N_6039,N_5240);
or U10521 (N_10521,N_7549,N_7400);
and U10522 (N_10522,N_7095,N_5351);
nor U10523 (N_10523,N_5186,N_7400);
xnor U10524 (N_10524,N_4260,N_7728);
or U10525 (N_10525,N_7892,N_5701);
nor U10526 (N_10526,N_7970,N_4390);
and U10527 (N_10527,N_5235,N_6045);
nor U10528 (N_10528,N_4285,N_5036);
nand U10529 (N_10529,N_5673,N_4867);
nand U10530 (N_10530,N_5759,N_7266);
nand U10531 (N_10531,N_7486,N_5249);
xnor U10532 (N_10532,N_4389,N_6354);
nor U10533 (N_10533,N_7528,N_4248);
or U10534 (N_10534,N_5429,N_7258);
and U10535 (N_10535,N_5616,N_7189);
xor U10536 (N_10536,N_5495,N_4011);
nand U10537 (N_10537,N_4776,N_6776);
nor U10538 (N_10538,N_7754,N_6154);
xor U10539 (N_10539,N_4618,N_7303);
nand U10540 (N_10540,N_4818,N_4396);
or U10541 (N_10541,N_7583,N_4964);
and U10542 (N_10542,N_4582,N_4228);
xnor U10543 (N_10543,N_5951,N_4958);
nand U10544 (N_10544,N_7432,N_4002);
and U10545 (N_10545,N_7423,N_7250);
xnor U10546 (N_10546,N_7476,N_5693);
xnor U10547 (N_10547,N_6952,N_6994);
nand U10548 (N_10548,N_7036,N_4200);
nand U10549 (N_10549,N_5433,N_4720);
and U10550 (N_10550,N_5548,N_5521);
nand U10551 (N_10551,N_7111,N_7071);
nor U10552 (N_10552,N_5528,N_4496);
or U10553 (N_10553,N_6991,N_7819);
and U10554 (N_10554,N_4701,N_6967);
and U10555 (N_10555,N_6621,N_5955);
xnor U10556 (N_10556,N_7757,N_7675);
nor U10557 (N_10557,N_6663,N_4924);
nor U10558 (N_10558,N_4655,N_4202);
nor U10559 (N_10559,N_5429,N_5601);
nor U10560 (N_10560,N_6193,N_6809);
and U10561 (N_10561,N_6247,N_4455);
nor U10562 (N_10562,N_7507,N_7545);
and U10563 (N_10563,N_6029,N_7002);
nand U10564 (N_10564,N_5146,N_6700);
or U10565 (N_10565,N_4710,N_4286);
or U10566 (N_10566,N_5121,N_4729);
xor U10567 (N_10567,N_7393,N_7106);
or U10568 (N_10568,N_5661,N_4221);
nand U10569 (N_10569,N_7625,N_6280);
and U10570 (N_10570,N_4170,N_6234);
and U10571 (N_10571,N_5515,N_7717);
nand U10572 (N_10572,N_6224,N_7835);
xnor U10573 (N_10573,N_6080,N_7472);
and U10574 (N_10574,N_5053,N_5031);
and U10575 (N_10575,N_6499,N_5297);
nand U10576 (N_10576,N_4934,N_5416);
nor U10577 (N_10577,N_4002,N_5734);
and U10578 (N_10578,N_5951,N_4873);
nor U10579 (N_10579,N_4842,N_4082);
or U10580 (N_10580,N_5660,N_6186);
or U10581 (N_10581,N_4564,N_4307);
and U10582 (N_10582,N_7943,N_5970);
xor U10583 (N_10583,N_7741,N_5779);
nand U10584 (N_10584,N_7153,N_5768);
nand U10585 (N_10585,N_5558,N_7336);
nor U10586 (N_10586,N_6771,N_7754);
nor U10587 (N_10587,N_5719,N_7238);
xnor U10588 (N_10588,N_5548,N_5761);
xnor U10589 (N_10589,N_6157,N_6177);
xnor U10590 (N_10590,N_4896,N_5792);
or U10591 (N_10591,N_7281,N_4550);
nand U10592 (N_10592,N_4012,N_6924);
or U10593 (N_10593,N_5418,N_7365);
xnor U10594 (N_10594,N_4921,N_6978);
and U10595 (N_10595,N_7395,N_4818);
or U10596 (N_10596,N_7611,N_4968);
nor U10597 (N_10597,N_7809,N_5825);
or U10598 (N_10598,N_4110,N_7072);
and U10599 (N_10599,N_7416,N_4805);
nand U10600 (N_10600,N_5572,N_7058);
xnor U10601 (N_10601,N_4083,N_4645);
nor U10602 (N_10602,N_7532,N_5183);
or U10603 (N_10603,N_5995,N_7864);
nor U10604 (N_10604,N_4435,N_5612);
nor U10605 (N_10605,N_4920,N_5344);
nand U10606 (N_10606,N_7695,N_7800);
and U10607 (N_10607,N_5338,N_6079);
nor U10608 (N_10608,N_4119,N_5748);
or U10609 (N_10609,N_6672,N_5524);
nor U10610 (N_10610,N_5576,N_6848);
xor U10611 (N_10611,N_6520,N_5655);
xor U10612 (N_10612,N_5631,N_6608);
or U10613 (N_10613,N_5338,N_7581);
or U10614 (N_10614,N_6118,N_6987);
nand U10615 (N_10615,N_7681,N_5132);
nand U10616 (N_10616,N_6264,N_4124);
or U10617 (N_10617,N_4890,N_6501);
and U10618 (N_10618,N_7745,N_4599);
xor U10619 (N_10619,N_7816,N_6071);
nor U10620 (N_10620,N_5434,N_7533);
or U10621 (N_10621,N_5937,N_7658);
or U10622 (N_10622,N_6288,N_6186);
or U10623 (N_10623,N_7274,N_6675);
xnor U10624 (N_10624,N_4784,N_5553);
or U10625 (N_10625,N_6096,N_6989);
nor U10626 (N_10626,N_6275,N_5553);
nor U10627 (N_10627,N_5067,N_4276);
nor U10628 (N_10628,N_6697,N_5540);
nor U10629 (N_10629,N_7127,N_5792);
nand U10630 (N_10630,N_5280,N_4512);
or U10631 (N_10631,N_6830,N_7113);
and U10632 (N_10632,N_4558,N_7443);
xor U10633 (N_10633,N_6543,N_7775);
or U10634 (N_10634,N_5753,N_4306);
xnor U10635 (N_10635,N_4709,N_7323);
nor U10636 (N_10636,N_6175,N_5937);
xnor U10637 (N_10637,N_6210,N_7027);
nor U10638 (N_10638,N_4877,N_5799);
and U10639 (N_10639,N_6744,N_7981);
and U10640 (N_10640,N_6261,N_7889);
nor U10641 (N_10641,N_4902,N_5301);
and U10642 (N_10642,N_6134,N_5702);
and U10643 (N_10643,N_7026,N_6683);
or U10644 (N_10644,N_7124,N_5553);
and U10645 (N_10645,N_6046,N_4800);
nand U10646 (N_10646,N_6903,N_5017);
or U10647 (N_10647,N_4201,N_6744);
nand U10648 (N_10648,N_7830,N_5641);
nor U10649 (N_10649,N_7674,N_4109);
nand U10650 (N_10650,N_6677,N_6334);
nor U10651 (N_10651,N_6182,N_6966);
xor U10652 (N_10652,N_7884,N_5359);
and U10653 (N_10653,N_5893,N_7453);
nand U10654 (N_10654,N_6647,N_5083);
or U10655 (N_10655,N_5707,N_6265);
nor U10656 (N_10656,N_4484,N_4980);
or U10657 (N_10657,N_5622,N_6732);
xor U10658 (N_10658,N_4746,N_4142);
xor U10659 (N_10659,N_6026,N_7310);
or U10660 (N_10660,N_7823,N_5041);
nand U10661 (N_10661,N_5326,N_5576);
xor U10662 (N_10662,N_4995,N_4587);
nor U10663 (N_10663,N_4545,N_7619);
or U10664 (N_10664,N_4309,N_5392);
nand U10665 (N_10665,N_7063,N_5052);
xnor U10666 (N_10666,N_6828,N_7566);
and U10667 (N_10667,N_5971,N_5558);
xor U10668 (N_10668,N_5694,N_5093);
nor U10669 (N_10669,N_7543,N_4452);
and U10670 (N_10670,N_6886,N_5730);
nand U10671 (N_10671,N_4261,N_4452);
and U10672 (N_10672,N_6745,N_6507);
or U10673 (N_10673,N_4103,N_4106);
nand U10674 (N_10674,N_7466,N_6682);
nor U10675 (N_10675,N_5941,N_7060);
and U10676 (N_10676,N_6021,N_5464);
or U10677 (N_10677,N_6016,N_4270);
xor U10678 (N_10678,N_5360,N_5030);
nand U10679 (N_10679,N_4757,N_6356);
and U10680 (N_10680,N_4619,N_5555);
and U10681 (N_10681,N_7183,N_4159);
nor U10682 (N_10682,N_5060,N_5969);
or U10683 (N_10683,N_5595,N_6094);
nand U10684 (N_10684,N_6293,N_5863);
nor U10685 (N_10685,N_5960,N_6306);
xor U10686 (N_10686,N_4149,N_4760);
xor U10687 (N_10687,N_4741,N_4618);
xnor U10688 (N_10688,N_4676,N_4276);
xor U10689 (N_10689,N_4635,N_7996);
nor U10690 (N_10690,N_4033,N_4060);
or U10691 (N_10691,N_5067,N_5652);
nand U10692 (N_10692,N_6145,N_7823);
nor U10693 (N_10693,N_7133,N_4209);
or U10694 (N_10694,N_5645,N_4747);
nand U10695 (N_10695,N_6094,N_4055);
and U10696 (N_10696,N_4357,N_4811);
and U10697 (N_10697,N_4126,N_5919);
or U10698 (N_10698,N_6205,N_5396);
and U10699 (N_10699,N_7314,N_4513);
or U10700 (N_10700,N_7702,N_5798);
xor U10701 (N_10701,N_6119,N_7146);
xor U10702 (N_10702,N_7798,N_4708);
nor U10703 (N_10703,N_4355,N_6025);
nor U10704 (N_10704,N_6863,N_4631);
xor U10705 (N_10705,N_6550,N_7997);
nor U10706 (N_10706,N_7414,N_7572);
nand U10707 (N_10707,N_5418,N_6852);
and U10708 (N_10708,N_7879,N_6578);
nand U10709 (N_10709,N_7473,N_6458);
nor U10710 (N_10710,N_7229,N_7086);
nor U10711 (N_10711,N_6754,N_4426);
nand U10712 (N_10712,N_7840,N_6782);
nand U10713 (N_10713,N_5695,N_7903);
nor U10714 (N_10714,N_7831,N_5449);
and U10715 (N_10715,N_6354,N_6653);
nand U10716 (N_10716,N_4701,N_7123);
or U10717 (N_10717,N_4828,N_6733);
xor U10718 (N_10718,N_4030,N_7892);
xnor U10719 (N_10719,N_4968,N_7151);
xnor U10720 (N_10720,N_6065,N_7467);
nor U10721 (N_10721,N_6011,N_5857);
xor U10722 (N_10722,N_5710,N_7600);
xor U10723 (N_10723,N_7620,N_5970);
nor U10724 (N_10724,N_6991,N_4676);
and U10725 (N_10725,N_5558,N_4963);
xnor U10726 (N_10726,N_5263,N_4790);
or U10727 (N_10727,N_5607,N_4679);
nand U10728 (N_10728,N_5571,N_6882);
nor U10729 (N_10729,N_7041,N_4606);
nand U10730 (N_10730,N_6506,N_4600);
nand U10731 (N_10731,N_4301,N_7597);
or U10732 (N_10732,N_7231,N_7324);
or U10733 (N_10733,N_7809,N_6137);
xor U10734 (N_10734,N_4536,N_7335);
xnor U10735 (N_10735,N_5578,N_5091);
nand U10736 (N_10736,N_6355,N_6622);
and U10737 (N_10737,N_7137,N_5640);
nand U10738 (N_10738,N_6687,N_4828);
xor U10739 (N_10739,N_4279,N_4183);
nor U10740 (N_10740,N_6600,N_5652);
nand U10741 (N_10741,N_4960,N_5552);
and U10742 (N_10742,N_5505,N_6935);
and U10743 (N_10743,N_7620,N_5429);
and U10744 (N_10744,N_7036,N_6441);
nor U10745 (N_10745,N_4521,N_7520);
xnor U10746 (N_10746,N_4841,N_5255);
xor U10747 (N_10747,N_4542,N_5487);
nor U10748 (N_10748,N_4353,N_5781);
and U10749 (N_10749,N_6378,N_4142);
or U10750 (N_10750,N_4228,N_7854);
or U10751 (N_10751,N_5902,N_5907);
nand U10752 (N_10752,N_4844,N_6100);
nand U10753 (N_10753,N_5297,N_5975);
and U10754 (N_10754,N_7949,N_4579);
nor U10755 (N_10755,N_5142,N_7081);
nor U10756 (N_10756,N_7792,N_6417);
nor U10757 (N_10757,N_5728,N_4299);
and U10758 (N_10758,N_5634,N_6427);
nor U10759 (N_10759,N_4457,N_4895);
and U10760 (N_10760,N_7184,N_6769);
xor U10761 (N_10761,N_6717,N_6366);
nor U10762 (N_10762,N_4107,N_4936);
nor U10763 (N_10763,N_4807,N_4610);
and U10764 (N_10764,N_7554,N_5479);
and U10765 (N_10765,N_7624,N_7634);
nand U10766 (N_10766,N_4298,N_7561);
or U10767 (N_10767,N_6504,N_7615);
nand U10768 (N_10768,N_5664,N_4951);
xor U10769 (N_10769,N_5600,N_5386);
nand U10770 (N_10770,N_5270,N_4219);
or U10771 (N_10771,N_6417,N_6464);
xor U10772 (N_10772,N_4184,N_7988);
nand U10773 (N_10773,N_4180,N_7123);
and U10774 (N_10774,N_6152,N_6574);
xor U10775 (N_10775,N_7371,N_6899);
or U10776 (N_10776,N_4941,N_7699);
nand U10777 (N_10777,N_6817,N_4523);
and U10778 (N_10778,N_7650,N_6950);
and U10779 (N_10779,N_5113,N_7147);
xnor U10780 (N_10780,N_6851,N_4915);
xnor U10781 (N_10781,N_5846,N_6452);
nand U10782 (N_10782,N_5830,N_4357);
or U10783 (N_10783,N_7834,N_6368);
xor U10784 (N_10784,N_7262,N_5062);
xnor U10785 (N_10785,N_6259,N_6866);
nand U10786 (N_10786,N_4266,N_5495);
nand U10787 (N_10787,N_6919,N_6160);
nand U10788 (N_10788,N_4191,N_6725);
nand U10789 (N_10789,N_7425,N_6981);
nand U10790 (N_10790,N_6336,N_5418);
and U10791 (N_10791,N_4279,N_7305);
and U10792 (N_10792,N_5751,N_6219);
and U10793 (N_10793,N_6290,N_7903);
xnor U10794 (N_10794,N_7307,N_5561);
or U10795 (N_10795,N_6675,N_4354);
nor U10796 (N_10796,N_7484,N_7456);
and U10797 (N_10797,N_5638,N_6442);
nand U10798 (N_10798,N_5150,N_5361);
nand U10799 (N_10799,N_5902,N_6857);
nor U10800 (N_10800,N_6197,N_5222);
nor U10801 (N_10801,N_7422,N_7007);
and U10802 (N_10802,N_4929,N_7915);
nor U10803 (N_10803,N_5453,N_7132);
xor U10804 (N_10804,N_7089,N_6881);
xor U10805 (N_10805,N_5143,N_5703);
or U10806 (N_10806,N_4939,N_5017);
nor U10807 (N_10807,N_5595,N_7165);
nor U10808 (N_10808,N_7740,N_5842);
nor U10809 (N_10809,N_6017,N_5049);
or U10810 (N_10810,N_6933,N_5996);
or U10811 (N_10811,N_5094,N_7521);
nand U10812 (N_10812,N_6818,N_7735);
nor U10813 (N_10813,N_7450,N_5548);
xor U10814 (N_10814,N_5044,N_5136);
and U10815 (N_10815,N_6849,N_6099);
or U10816 (N_10816,N_5786,N_6658);
nor U10817 (N_10817,N_7627,N_5912);
or U10818 (N_10818,N_4148,N_5703);
nand U10819 (N_10819,N_6445,N_6965);
nor U10820 (N_10820,N_5429,N_5017);
and U10821 (N_10821,N_4084,N_6517);
and U10822 (N_10822,N_7777,N_7923);
xor U10823 (N_10823,N_4783,N_6327);
nor U10824 (N_10824,N_4945,N_4316);
nand U10825 (N_10825,N_5299,N_7756);
or U10826 (N_10826,N_5977,N_5458);
nor U10827 (N_10827,N_7539,N_4009);
xor U10828 (N_10828,N_6957,N_4965);
or U10829 (N_10829,N_7237,N_5292);
and U10830 (N_10830,N_4811,N_7635);
nor U10831 (N_10831,N_6161,N_6122);
and U10832 (N_10832,N_4818,N_5955);
and U10833 (N_10833,N_7977,N_4134);
or U10834 (N_10834,N_7298,N_6023);
xor U10835 (N_10835,N_4058,N_4577);
xor U10836 (N_10836,N_4962,N_5519);
nand U10837 (N_10837,N_5166,N_6904);
nand U10838 (N_10838,N_7278,N_7817);
or U10839 (N_10839,N_5555,N_7329);
or U10840 (N_10840,N_6695,N_7770);
xor U10841 (N_10841,N_6820,N_4200);
nand U10842 (N_10842,N_5640,N_6357);
nand U10843 (N_10843,N_7873,N_7489);
nor U10844 (N_10844,N_5861,N_5874);
or U10845 (N_10845,N_4124,N_5588);
xor U10846 (N_10846,N_6137,N_6947);
nor U10847 (N_10847,N_4048,N_6902);
xor U10848 (N_10848,N_7378,N_4699);
xnor U10849 (N_10849,N_4704,N_5818);
nand U10850 (N_10850,N_4146,N_7349);
xnor U10851 (N_10851,N_4865,N_5579);
or U10852 (N_10852,N_4749,N_5460);
xnor U10853 (N_10853,N_6559,N_5020);
or U10854 (N_10854,N_6120,N_6036);
nand U10855 (N_10855,N_6617,N_4863);
nand U10856 (N_10856,N_5362,N_6505);
and U10857 (N_10857,N_6661,N_4573);
and U10858 (N_10858,N_7644,N_5890);
or U10859 (N_10859,N_7948,N_7400);
and U10860 (N_10860,N_6711,N_5461);
and U10861 (N_10861,N_4553,N_7131);
xor U10862 (N_10862,N_7112,N_4483);
or U10863 (N_10863,N_5890,N_5356);
nor U10864 (N_10864,N_7931,N_6950);
or U10865 (N_10865,N_4288,N_7679);
nand U10866 (N_10866,N_5464,N_7170);
or U10867 (N_10867,N_6586,N_5665);
xnor U10868 (N_10868,N_6010,N_5412);
and U10869 (N_10869,N_5385,N_5594);
xnor U10870 (N_10870,N_6419,N_4290);
nor U10871 (N_10871,N_6858,N_7642);
nand U10872 (N_10872,N_7254,N_4267);
or U10873 (N_10873,N_6491,N_4357);
nor U10874 (N_10874,N_5713,N_7490);
and U10875 (N_10875,N_5392,N_7554);
xor U10876 (N_10876,N_4138,N_7330);
or U10877 (N_10877,N_4485,N_4205);
or U10878 (N_10878,N_5717,N_7439);
and U10879 (N_10879,N_5696,N_7531);
nor U10880 (N_10880,N_4925,N_7395);
or U10881 (N_10881,N_6729,N_6281);
or U10882 (N_10882,N_5631,N_5465);
nor U10883 (N_10883,N_7521,N_4925);
nand U10884 (N_10884,N_6467,N_4516);
nor U10885 (N_10885,N_6073,N_6667);
nor U10886 (N_10886,N_5960,N_6925);
nor U10887 (N_10887,N_7084,N_4053);
nor U10888 (N_10888,N_6254,N_6363);
nand U10889 (N_10889,N_5518,N_4377);
xor U10890 (N_10890,N_4850,N_7946);
nand U10891 (N_10891,N_5573,N_4102);
nor U10892 (N_10892,N_4654,N_5552);
xor U10893 (N_10893,N_6900,N_4789);
nand U10894 (N_10894,N_4333,N_7263);
and U10895 (N_10895,N_5830,N_4878);
and U10896 (N_10896,N_4398,N_4331);
nand U10897 (N_10897,N_4065,N_5943);
and U10898 (N_10898,N_6440,N_5330);
and U10899 (N_10899,N_7162,N_4610);
and U10900 (N_10900,N_4926,N_5499);
xnor U10901 (N_10901,N_7808,N_7922);
nor U10902 (N_10902,N_7805,N_6752);
and U10903 (N_10903,N_6955,N_5182);
and U10904 (N_10904,N_5222,N_5659);
nand U10905 (N_10905,N_6928,N_5369);
xor U10906 (N_10906,N_5739,N_4645);
xor U10907 (N_10907,N_6290,N_7172);
nand U10908 (N_10908,N_6336,N_6579);
nand U10909 (N_10909,N_6206,N_4965);
or U10910 (N_10910,N_4310,N_4600);
or U10911 (N_10911,N_6118,N_4838);
nand U10912 (N_10912,N_6384,N_5598);
xor U10913 (N_10913,N_5832,N_7289);
or U10914 (N_10914,N_7062,N_7622);
xor U10915 (N_10915,N_4432,N_4169);
and U10916 (N_10916,N_6390,N_5161);
nand U10917 (N_10917,N_6407,N_6395);
nand U10918 (N_10918,N_5557,N_5966);
or U10919 (N_10919,N_7875,N_6771);
xnor U10920 (N_10920,N_4592,N_5525);
nand U10921 (N_10921,N_5368,N_7485);
or U10922 (N_10922,N_4713,N_7050);
or U10923 (N_10923,N_4353,N_7680);
nor U10924 (N_10924,N_5964,N_7356);
or U10925 (N_10925,N_7252,N_7910);
or U10926 (N_10926,N_6287,N_4077);
or U10927 (N_10927,N_7231,N_4709);
xnor U10928 (N_10928,N_6858,N_5112);
nor U10929 (N_10929,N_4882,N_7529);
nor U10930 (N_10930,N_5862,N_4702);
nor U10931 (N_10931,N_4718,N_6253);
or U10932 (N_10932,N_5736,N_4499);
nor U10933 (N_10933,N_5135,N_4898);
nand U10934 (N_10934,N_4437,N_4269);
xor U10935 (N_10935,N_6339,N_6351);
or U10936 (N_10936,N_5162,N_5144);
and U10937 (N_10937,N_5973,N_4854);
xnor U10938 (N_10938,N_4156,N_6580);
nand U10939 (N_10939,N_4616,N_4283);
or U10940 (N_10940,N_7224,N_7840);
or U10941 (N_10941,N_6683,N_5131);
xnor U10942 (N_10942,N_5413,N_7514);
nor U10943 (N_10943,N_4370,N_4056);
or U10944 (N_10944,N_4482,N_5937);
nor U10945 (N_10945,N_7655,N_6908);
or U10946 (N_10946,N_4654,N_4529);
and U10947 (N_10947,N_5946,N_6198);
nand U10948 (N_10948,N_7143,N_6927);
and U10949 (N_10949,N_4055,N_4893);
or U10950 (N_10950,N_5394,N_5535);
nand U10951 (N_10951,N_7775,N_4516);
xor U10952 (N_10952,N_5154,N_6807);
xnor U10953 (N_10953,N_5071,N_5321);
or U10954 (N_10954,N_6730,N_4829);
xnor U10955 (N_10955,N_6833,N_5563);
nand U10956 (N_10956,N_4577,N_5752);
or U10957 (N_10957,N_7135,N_5459);
nand U10958 (N_10958,N_4556,N_5331);
and U10959 (N_10959,N_6148,N_6618);
or U10960 (N_10960,N_6981,N_6306);
and U10961 (N_10961,N_7498,N_6187);
nand U10962 (N_10962,N_7465,N_6580);
nand U10963 (N_10963,N_5335,N_7405);
nor U10964 (N_10964,N_6222,N_7811);
xnor U10965 (N_10965,N_6168,N_5926);
or U10966 (N_10966,N_7509,N_6293);
and U10967 (N_10967,N_5915,N_4870);
or U10968 (N_10968,N_7167,N_4160);
nor U10969 (N_10969,N_4557,N_5861);
or U10970 (N_10970,N_7670,N_6334);
xor U10971 (N_10971,N_6155,N_6862);
nand U10972 (N_10972,N_7182,N_5430);
xnor U10973 (N_10973,N_4120,N_7426);
and U10974 (N_10974,N_7347,N_6427);
or U10975 (N_10975,N_4030,N_7071);
nor U10976 (N_10976,N_7155,N_7857);
and U10977 (N_10977,N_4062,N_7329);
or U10978 (N_10978,N_4224,N_4659);
nand U10979 (N_10979,N_5070,N_4167);
xnor U10980 (N_10980,N_6034,N_7350);
or U10981 (N_10981,N_4411,N_5601);
and U10982 (N_10982,N_6610,N_4071);
or U10983 (N_10983,N_6708,N_5812);
xor U10984 (N_10984,N_6088,N_7501);
and U10985 (N_10985,N_4508,N_7671);
nand U10986 (N_10986,N_5632,N_6752);
or U10987 (N_10987,N_7343,N_6937);
nor U10988 (N_10988,N_5543,N_7268);
nand U10989 (N_10989,N_4550,N_4597);
nor U10990 (N_10990,N_7107,N_5707);
or U10991 (N_10991,N_6138,N_5416);
xnor U10992 (N_10992,N_6402,N_7084);
or U10993 (N_10993,N_6014,N_7687);
and U10994 (N_10994,N_6088,N_6439);
and U10995 (N_10995,N_6364,N_4468);
or U10996 (N_10996,N_6116,N_4504);
xnor U10997 (N_10997,N_7517,N_7180);
xnor U10998 (N_10998,N_6146,N_7732);
nor U10999 (N_10999,N_4573,N_7297);
or U11000 (N_11000,N_6315,N_6009);
nand U11001 (N_11001,N_6994,N_6581);
nor U11002 (N_11002,N_6326,N_7578);
or U11003 (N_11003,N_4145,N_6711);
xor U11004 (N_11004,N_5213,N_4217);
xnor U11005 (N_11005,N_5078,N_7998);
or U11006 (N_11006,N_7298,N_4579);
and U11007 (N_11007,N_5795,N_6052);
and U11008 (N_11008,N_4834,N_4728);
xnor U11009 (N_11009,N_5961,N_4191);
nand U11010 (N_11010,N_5681,N_5608);
or U11011 (N_11011,N_7497,N_6060);
xnor U11012 (N_11012,N_5440,N_6735);
xnor U11013 (N_11013,N_4837,N_7359);
xnor U11014 (N_11014,N_6418,N_5759);
nor U11015 (N_11015,N_4729,N_6743);
xor U11016 (N_11016,N_7552,N_7785);
nor U11017 (N_11017,N_5652,N_7844);
xnor U11018 (N_11018,N_6809,N_6652);
and U11019 (N_11019,N_4211,N_7310);
xnor U11020 (N_11020,N_5752,N_7870);
nor U11021 (N_11021,N_4958,N_4220);
nor U11022 (N_11022,N_4742,N_6215);
and U11023 (N_11023,N_7858,N_4798);
or U11024 (N_11024,N_6605,N_6512);
or U11025 (N_11025,N_4648,N_7890);
nand U11026 (N_11026,N_7490,N_7402);
or U11027 (N_11027,N_7654,N_5676);
and U11028 (N_11028,N_7625,N_4776);
nor U11029 (N_11029,N_5718,N_7248);
and U11030 (N_11030,N_5085,N_5955);
nand U11031 (N_11031,N_7535,N_7086);
and U11032 (N_11032,N_4215,N_5269);
and U11033 (N_11033,N_7017,N_4351);
nor U11034 (N_11034,N_5897,N_4976);
nand U11035 (N_11035,N_4835,N_6117);
nand U11036 (N_11036,N_5584,N_5617);
nand U11037 (N_11037,N_5081,N_7504);
xnor U11038 (N_11038,N_5422,N_6761);
and U11039 (N_11039,N_4857,N_5390);
nor U11040 (N_11040,N_4384,N_4633);
and U11041 (N_11041,N_4763,N_7139);
and U11042 (N_11042,N_6827,N_4485);
nand U11043 (N_11043,N_5587,N_6840);
nor U11044 (N_11044,N_7836,N_5049);
or U11045 (N_11045,N_5416,N_7154);
or U11046 (N_11046,N_6894,N_5555);
or U11047 (N_11047,N_6629,N_6014);
nand U11048 (N_11048,N_4228,N_7061);
nand U11049 (N_11049,N_4032,N_7832);
nand U11050 (N_11050,N_6644,N_4350);
nand U11051 (N_11051,N_7952,N_5999);
and U11052 (N_11052,N_4092,N_6707);
and U11053 (N_11053,N_7968,N_4880);
xnor U11054 (N_11054,N_5360,N_4304);
xor U11055 (N_11055,N_6568,N_6080);
nor U11056 (N_11056,N_6373,N_4830);
and U11057 (N_11057,N_4630,N_4383);
and U11058 (N_11058,N_7883,N_7426);
xnor U11059 (N_11059,N_7790,N_4215);
nand U11060 (N_11060,N_4517,N_5156);
or U11061 (N_11061,N_4722,N_4452);
nor U11062 (N_11062,N_4277,N_4465);
xor U11063 (N_11063,N_5483,N_7952);
and U11064 (N_11064,N_4898,N_5145);
nand U11065 (N_11065,N_6538,N_7745);
or U11066 (N_11066,N_4343,N_4166);
nor U11067 (N_11067,N_4969,N_7909);
nor U11068 (N_11068,N_6276,N_4493);
xnor U11069 (N_11069,N_4847,N_5543);
xnor U11070 (N_11070,N_4919,N_5585);
xnor U11071 (N_11071,N_5791,N_7980);
nor U11072 (N_11072,N_5250,N_5917);
or U11073 (N_11073,N_5693,N_6739);
and U11074 (N_11074,N_6895,N_6241);
or U11075 (N_11075,N_4347,N_5224);
nand U11076 (N_11076,N_7787,N_6859);
and U11077 (N_11077,N_6374,N_7762);
or U11078 (N_11078,N_7627,N_7063);
or U11079 (N_11079,N_6888,N_4408);
nand U11080 (N_11080,N_4065,N_5698);
nand U11081 (N_11081,N_7610,N_5339);
xor U11082 (N_11082,N_5630,N_5648);
and U11083 (N_11083,N_4366,N_6467);
nand U11084 (N_11084,N_7115,N_5786);
xor U11085 (N_11085,N_7955,N_7291);
xnor U11086 (N_11086,N_4039,N_4315);
and U11087 (N_11087,N_4133,N_6170);
nand U11088 (N_11088,N_5391,N_5161);
xnor U11089 (N_11089,N_4712,N_7796);
xnor U11090 (N_11090,N_4837,N_6303);
or U11091 (N_11091,N_6670,N_7674);
and U11092 (N_11092,N_4519,N_4573);
nand U11093 (N_11093,N_4722,N_4123);
nor U11094 (N_11094,N_7622,N_6461);
and U11095 (N_11095,N_4824,N_4560);
xnor U11096 (N_11096,N_7871,N_7283);
xnor U11097 (N_11097,N_7931,N_6700);
and U11098 (N_11098,N_4374,N_6147);
and U11099 (N_11099,N_5129,N_6047);
xnor U11100 (N_11100,N_7081,N_7012);
nor U11101 (N_11101,N_4602,N_5360);
xor U11102 (N_11102,N_5723,N_7751);
or U11103 (N_11103,N_7551,N_5207);
nor U11104 (N_11104,N_7854,N_7641);
or U11105 (N_11105,N_7170,N_7637);
nor U11106 (N_11106,N_4435,N_6464);
or U11107 (N_11107,N_7727,N_4398);
xor U11108 (N_11108,N_6221,N_5359);
nor U11109 (N_11109,N_7137,N_7691);
nand U11110 (N_11110,N_4468,N_6641);
xor U11111 (N_11111,N_5157,N_5451);
nand U11112 (N_11112,N_4620,N_7691);
and U11113 (N_11113,N_6924,N_4973);
nor U11114 (N_11114,N_5275,N_4697);
nor U11115 (N_11115,N_5762,N_6355);
and U11116 (N_11116,N_5672,N_6342);
nor U11117 (N_11117,N_4515,N_6841);
nor U11118 (N_11118,N_6201,N_7083);
xor U11119 (N_11119,N_4659,N_6418);
nor U11120 (N_11120,N_6603,N_4295);
xor U11121 (N_11121,N_4453,N_5916);
or U11122 (N_11122,N_6242,N_7998);
and U11123 (N_11123,N_4167,N_4171);
and U11124 (N_11124,N_6240,N_7401);
xnor U11125 (N_11125,N_5928,N_6506);
nand U11126 (N_11126,N_6841,N_4580);
and U11127 (N_11127,N_7771,N_5275);
nor U11128 (N_11128,N_5012,N_4888);
or U11129 (N_11129,N_4837,N_5470);
and U11130 (N_11130,N_5817,N_5672);
and U11131 (N_11131,N_7992,N_6951);
nor U11132 (N_11132,N_7895,N_4841);
xor U11133 (N_11133,N_7921,N_4444);
nor U11134 (N_11134,N_7693,N_6935);
xnor U11135 (N_11135,N_4892,N_5637);
and U11136 (N_11136,N_5453,N_7122);
nand U11137 (N_11137,N_4824,N_5128);
xor U11138 (N_11138,N_4971,N_4133);
or U11139 (N_11139,N_4086,N_7872);
or U11140 (N_11140,N_6033,N_4353);
nor U11141 (N_11141,N_5926,N_4980);
and U11142 (N_11142,N_7679,N_7400);
nand U11143 (N_11143,N_4014,N_4041);
or U11144 (N_11144,N_7342,N_4064);
xnor U11145 (N_11145,N_4084,N_5872);
or U11146 (N_11146,N_5430,N_6269);
or U11147 (N_11147,N_5919,N_5405);
or U11148 (N_11148,N_7077,N_7420);
nor U11149 (N_11149,N_4217,N_5017);
or U11150 (N_11150,N_5639,N_7375);
xnor U11151 (N_11151,N_6159,N_7380);
nand U11152 (N_11152,N_5006,N_5305);
or U11153 (N_11153,N_7937,N_7510);
xnor U11154 (N_11154,N_7646,N_7962);
and U11155 (N_11155,N_4211,N_5761);
nor U11156 (N_11156,N_5835,N_4744);
xnor U11157 (N_11157,N_7479,N_6692);
xor U11158 (N_11158,N_5930,N_4926);
or U11159 (N_11159,N_4300,N_4328);
and U11160 (N_11160,N_7846,N_4675);
xor U11161 (N_11161,N_5292,N_5782);
or U11162 (N_11162,N_7577,N_7512);
xor U11163 (N_11163,N_6190,N_6687);
or U11164 (N_11164,N_7503,N_6208);
nand U11165 (N_11165,N_5456,N_7810);
xor U11166 (N_11166,N_6105,N_7017);
nor U11167 (N_11167,N_6329,N_6948);
and U11168 (N_11168,N_4792,N_5132);
or U11169 (N_11169,N_7837,N_7523);
nand U11170 (N_11170,N_5358,N_6481);
nand U11171 (N_11171,N_5034,N_6933);
or U11172 (N_11172,N_6171,N_6346);
or U11173 (N_11173,N_5487,N_6744);
nor U11174 (N_11174,N_7499,N_6958);
or U11175 (N_11175,N_7909,N_5021);
or U11176 (N_11176,N_5413,N_6367);
nand U11177 (N_11177,N_4016,N_6310);
nand U11178 (N_11178,N_7323,N_6898);
and U11179 (N_11179,N_4843,N_4575);
xnor U11180 (N_11180,N_4544,N_4068);
nor U11181 (N_11181,N_7530,N_7303);
and U11182 (N_11182,N_5950,N_4550);
nand U11183 (N_11183,N_4066,N_7565);
xor U11184 (N_11184,N_7170,N_4371);
and U11185 (N_11185,N_5269,N_4331);
and U11186 (N_11186,N_6722,N_6003);
or U11187 (N_11187,N_6598,N_5420);
or U11188 (N_11188,N_7249,N_4767);
or U11189 (N_11189,N_4739,N_6496);
xor U11190 (N_11190,N_7386,N_4653);
or U11191 (N_11191,N_5631,N_4704);
nor U11192 (N_11192,N_6049,N_6118);
and U11193 (N_11193,N_6785,N_7086);
nor U11194 (N_11194,N_4688,N_7543);
and U11195 (N_11195,N_4776,N_4219);
nand U11196 (N_11196,N_7101,N_5942);
nand U11197 (N_11197,N_7647,N_6113);
nand U11198 (N_11198,N_4117,N_6075);
and U11199 (N_11199,N_4033,N_7431);
xor U11200 (N_11200,N_6409,N_6264);
and U11201 (N_11201,N_5602,N_7382);
xor U11202 (N_11202,N_5480,N_6736);
and U11203 (N_11203,N_5312,N_4320);
nor U11204 (N_11204,N_4389,N_5361);
and U11205 (N_11205,N_4613,N_6625);
nand U11206 (N_11206,N_5134,N_4840);
xor U11207 (N_11207,N_4197,N_5470);
or U11208 (N_11208,N_4602,N_5316);
or U11209 (N_11209,N_5023,N_4452);
xnor U11210 (N_11210,N_6214,N_4086);
or U11211 (N_11211,N_7650,N_4839);
nor U11212 (N_11212,N_7429,N_5018);
nor U11213 (N_11213,N_7328,N_6002);
nand U11214 (N_11214,N_6089,N_4921);
xor U11215 (N_11215,N_5044,N_7116);
and U11216 (N_11216,N_7252,N_7740);
xor U11217 (N_11217,N_4996,N_5092);
nand U11218 (N_11218,N_6857,N_5334);
and U11219 (N_11219,N_4521,N_7071);
xor U11220 (N_11220,N_5700,N_5549);
nor U11221 (N_11221,N_4177,N_6295);
nand U11222 (N_11222,N_6721,N_4715);
nor U11223 (N_11223,N_7603,N_6832);
and U11224 (N_11224,N_5018,N_7305);
xor U11225 (N_11225,N_5450,N_5377);
xor U11226 (N_11226,N_7846,N_4963);
nor U11227 (N_11227,N_5042,N_6185);
xor U11228 (N_11228,N_6630,N_6710);
nor U11229 (N_11229,N_5890,N_6812);
and U11230 (N_11230,N_4908,N_5345);
or U11231 (N_11231,N_4136,N_7616);
nor U11232 (N_11232,N_7369,N_4670);
nand U11233 (N_11233,N_6813,N_7404);
nor U11234 (N_11234,N_6875,N_7011);
xnor U11235 (N_11235,N_4138,N_6578);
nand U11236 (N_11236,N_7530,N_4607);
nor U11237 (N_11237,N_5594,N_4189);
or U11238 (N_11238,N_7058,N_5100);
nor U11239 (N_11239,N_4523,N_7415);
nand U11240 (N_11240,N_6409,N_6314);
nand U11241 (N_11241,N_4816,N_4282);
nor U11242 (N_11242,N_7028,N_7429);
xnor U11243 (N_11243,N_5949,N_6439);
nand U11244 (N_11244,N_5810,N_5153);
and U11245 (N_11245,N_7746,N_4988);
nor U11246 (N_11246,N_7477,N_5361);
nor U11247 (N_11247,N_4185,N_5135);
and U11248 (N_11248,N_6808,N_7647);
or U11249 (N_11249,N_4818,N_4345);
and U11250 (N_11250,N_5468,N_4778);
and U11251 (N_11251,N_5667,N_6826);
and U11252 (N_11252,N_7172,N_5127);
nand U11253 (N_11253,N_5510,N_7276);
and U11254 (N_11254,N_6335,N_7335);
nor U11255 (N_11255,N_4039,N_7843);
nand U11256 (N_11256,N_4260,N_7489);
or U11257 (N_11257,N_7480,N_6771);
or U11258 (N_11258,N_5995,N_6655);
xnor U11259 (N_11259,N_4825,N_5463);
nor U11260 (N_11260,N_7756,N_6766);
nand U11261 (N_11261,N_5288,N_7641);
nand U11262 (N_11262,N_6966,N_6041);
xnor U11263 (N_11263,N_5975,N_7459);
xnor U11264 (N_11264,N_5714,N_6621);
and U11265 (N_11265,N_4446,N_5078);
and U11266 (N_11266,N_6941,N_7557);
nand U11267 (N_11267,N_4103,N_6097);
nand U11268 (N_11268,N_7818,N_4589);
or U11269 (N_11269,N_4361,N_7887);
nand U11270 (N_11270,N_5235,N_5268);
and U11271 (N_11271,N_7164,N_7687);
xor U11272 (N_11272,N_6965,N_7146);
nand U11273 (N_11273,N_6136,N_5580);
xnor U11274 (N_11274,N_5105,N_4784);
xor U11275 (N_11275,N_5549,N_4554);
or U11276 (N_11276,N_5300,N_7726);
nand U11277 (N_11277,N_7521,N_5640);
nand U11278 (N_11278,N_5293,N_7736);
nand U11279 (N_11279,N_5344,N_4601);
xnor U11280 (N_11280,N_5621,N_5049);
nor U11281 (N_11281,N_4727,N_4517);
nor U11282 (N_11282,N_7142,N_4963);
and U11283 (N_11283,N_4479,N_4975);
xor U11284 (N_11284,N_6595,N_4964);
nand U11285 (N_11285,N_7435,N_4975);
xor U11286 (N_11286,N_6452,N_7587);
or U11287 (N_11287,N_4447,N_4968);
xnor U11288 (N_11288,N_6717,N_7086);
and U11289 (N_11289,N_7206,N_7659);
xor U11290 (N_11290,N_6308,N_6162);
or U11291 (N_11291,N_7797,N_7208);
nor U11292 (N_11292,N_4960,N_5928);
or U11293 (N_11293,N_4887,N_6321);
and U11294 (N_11294,N_6703,N_5041);
nand U11295 (N_11295,N_4481,N_6946);
and U11296 (N_11296,N_4400,N_5390);
or U11297 (N_11297,N_6447,N_6212);
or U11298 (N_11298,N_6168,N_6076);
xnor U11299 (N_11299,N_4474,N_4234);
and U11300 (N_11300,N_5242,N_7772);
nor U11301 (N_11301,N_4756,N_5580);
xor U11302 (N_11302,N_7575,N_7504);
and U11303 (N_11303,N_6985,N_7576);
nor U11304 (N_11304,N_4553,N_6436);
xnor U11305 (N_11305,N_7658,N_5525);
nand U11306 (N_11306,N_7356,N_6164);
or U11307 (N_11307,N_6848,N_7306);
xnor U11308 (N_11308,N_7350,N_5950);
nand U11309 (N_11309,N_7977,N_4077);
or U11310 (N_11310,N_4820,N_4217);
or U11311 (N_11311,N_6981,N_4082);
nand U11312 (N_11312,N_7288,N_5552);
or U11313 (N_11313,N_7474,N_5299);
and U11314 (N_11314,N_5601,N_7605);
xor U11315 (N_11315,N_7017,N_7294);
and U11316 (N_11316,N_6418,N_5887);
nor U11317 (N_11317,N_4966,N_6438);
and U11318 (N_11318,N_5284,N_6141);
xnor U11319 (N_11319,N_5457,N_7888);
xnor U11320 (N_11320,N_7584,N_7219);
nand U11321 (N_11321,N_5542,N_7521);
nor U11322 (N_11322,N_5975,N_4907);
xor U11323 (N_11323,N_7588,N_7107);
nand U11324 (N_11324,N_6282,N_5183);
nand U11325 (N_11325,N_7518,N_6585);
and U11326 (N_11326,N_4473,N_6469);
xnor U11327 (N_11327,N_5399,N_4301);
nand U11328 (N_11328,N_7816,N_7247);
and U11329 (N_11329,N_4644,N_6656);
or U11330 (N_11330,N_6826,N_7246);
nand U11331 (N_11331,N_6045,N_7227);
nand U11332 (N_11332,N_7721,N_7290);
xnor U11333 (N_11333,N_4731,N_7320);
and U11334 (N_11334,N_5690,N_4338);
and U11335 (N_11335,N_4917,N_4574);
and U11336 (N_11336,N_5006,N_6321);
and U11337 (N_11337,N_4105,N_7883);
nand U11338 (N_11338,N_4096,N_6800);
nand U11339 (N_11339,N_4921,N_5478);
xnor U11340 (N_11340,N_7758,N_4491);
and U11341 (N_11341,N_6302,N_5534);
and U11342 (N_11342,N_7715,N_6228);
nor U11343 (N_11343,N_7090,N_5175);
xor U11344 (N_11344,N_7662,N_6081);
xnor U11345 (N_11345,N_7274,N_4943);
nand U11346 (N_11346,N_6270,N_6722);
or U11347 (N_11347,N_4138,N_6579);
and U11348 (N_11348,N_5249,N_7442);
xor U11349 (N_11349,N_4908,N_5937);
nor U11350 (N_11350,N_4523,N_5739);
xnor U11351 (N_11351,N_5230,N_4093);
and U11352 (N_11352,N_4064,N_5625);
nor U11353 (N_11353,N_6960,N_4486);
or U11354 (N_11354,N_6383,N_6277);
nor U11355 (N_11355,N_4570,N_5491);
or U11356 (N_11356,N_5392,N_5503);
nor U11357 (N_11357,N_4716,N_4954);
or U11358 (N_11358,N_5014,N_4455);
nand U11359 (N_11359,N_5649,N_6624);
nor U11360 (N_11360,N_7878,N_5306);
nand U11361 (N_11361,N_5867,N_4530);
and U11362 (N_11362,N_6174,N_4250);
and U11363 (N_11363,N_5466,N_6023);
or U11364 (N_11364,N_5602,N_4241);
xor U11365 (N_11365,N_4751,N_4940);
or U11366 (N_11366,N_4713,N_7235);
nand U11367 (N_11367,N_7019,N_4104);
and U11368 (N_11368,N_5694,N_7739);
and U11369 (N_11369,N_6355,N_6858);
xnor U11370 (N_11370,N_5580,N_4186);
and U11371 (N_11371,N_4435,N_7155);
xor U11372 (N_11372,N_7333,N_5376);
nand U11373 (N_11373,N_5314,N_5109);
and U11374 (N_11374,N_6185,N_5307);
xnor U11375 (N_11375,N_5301,N_4748);
or U11376 (N_11376,N_7638,N_4749);
nand U11377 (N_11377,N_4649,N_5675);
nand U11378 (N_11378,N_6884,N_4258);
nand U11379 (N_11379,N_5529,N_4581);
nand U11380 (N_11380,N_5065,N_4961);
nand U11381 (N_11381,N_6752,N_6529);
or U11382 (N_11382,N_5041,N_5924);
and U11383 (N_11383,N_5408,N_7201);
xor U11384 (N_11384,N_7852,N_6565);
xnor U11385 (N_11385,N_7783,N_4427);
nand U11386 (N_11386,N_5146,N_6069);
nand U11387 (N_11387,N_5632,N_6738);
nor U11388 (N_11388,N_7098,N_7930);
or U11389 (N_11389,N_7756,N_5371);
and U11390 (N_11390,N_6998,N_5733);
or U11391 (N_11391,N_4423,N_5822);
nor U11392 (N_11392,N_4334,N_7021);
xnor U11393 (N_11393,N_6207,N_7977);
and U11394 (N_11394,N_7286,N_6563);
nor U11395 (N_11395,N_6008,N_5459);
or U11396 (N_11396,N_7464,N_6839);
xnor U11397 (N_11397,N_6153,N_4430);
nor U11398 (N_11398,N_4968,N_5796);
nor U11399 (N_11399,N_7194,N_7228);
nor U11400 (N_11400,N_5870,N_6766);
or U11401 (N_11401,N_5443,N_6173);
or U11402 (N_11402,N_5501,N_7385);
and U11403 (N_11403,N_5482,N_4659);
nor U11404 (N_11404,N_6818,N_7325);
nand U11405 (N_11405,N_5371,N_6487);
or U11406 (N_11406,N_6408,N_6316);
nor U11407 (N_11407,N_6587,N_4606);
or U11408 (N_11408,N_5386,N_6253);
or U11409 (N_11409,N_7940,N_5840);
nand U11410 (N_11410,N_4302,N_7398);
or U11411 (N_11411,N_7376,N_4567);
xnor U11412 (N_11412,N_6692,N_4908);
or U11413 (N_11413,N_4211,N_6313);
and U11414 (N_11414,N_7856,N_6941);
and U11415 (N_11415,N_5022,N_5587);
nor U11416 (N_11416,N_6830,N_6463);
and U11417 (N_11417,N_7784,N_6634);
or U11418 (N_11418,N_7774,N_5053);
or U11419 (N_11419,N_6711,N_5217);
nand U11420 (N_11420,N_7856,N_7180);
nor U11421 (N_11421,N_6907,N_6054);
or U11422 (N_11422,N_6650,N_5040);
and U11423 (N_11423,N_6396,N_4320);
xnor U11424 (N_11424,N_4392,N_5705);
and U11425 (N_11425,N_7785,N_7942);
and U11426 (N_11426,N_7419,N_7425);
xor U11427 (N_11427,N_5564,N_5878);
nand U11428 (N_11428,N_6404,N_4559);
and U11429 (N_11429,N_5989,N_5897);
and U11430 (N_11430,N_7290,N_5927);
or U11431 (N_11431,N_6792,N_7273);
and U11432 (N_11432,N_6457,N_5977);
and U11433 (N_11433,N_5508,N_6764);
or U11434 (N_11434,N_7869,N_5893);
or U11435 (N_11435,N_4993,N_7964);
or U11436 (N_11436,N_5169,N_4573);
and U11437 (N_11437,N_5977,N_6510);
and U11438 (N_11438,N_6682,N_6433);
nand U11439 (N_11439,N_6312,N_5157);
nand U11440 (N_11440,N_4524,N_4635);
nand U11441 (N_11441,N_6210,N_7649);
nand U11442 (N_11442,N_4856,N_5355);
xor U11443 (N_11443,N_4289,N_5727);
nor U11444 (N_11444,N_5661,N_5005);
or U11445 (N_11445,N_7558,N_7481);
nand U11446 (N_11446,N_6795,N_6188);
xor U11447 (N_11447,N_7060,N_7016);
and U11448 (N_11448,N_7576,N_6813);
and U11449 (N_11449,N_5842,N_7448);
nor U11450 (N_11450,N_4488,N_5763);
nand U11451 (N_11451,N_6523,N_4343);
and U11452 (N_11452,N_5307,N_7846);
or U11453 (N_11453,N_7421,N_7207);
and U11454 (N_11454,N_5752,N_7169);
nor U11455 (N_11455,N_4511,N_7112);
nand U11456 (N_11456,N_7599,N_7198);
nand U11457 (N_11457,N_5399,N_4350);
nand U11458 (N_11458,N_7984,N_6510);
and U11459 (N_11459,N_6290,N_4996);
xnor U11460 (N_11460,N_5112,N_4194);
and U11461 (N_11461,N_5569,N_7194);
nand U11462 (N_11462,N_6460,N_5892);
xor U11463 (N_11463,N_6278,N_7685);
or U11464 (N_11464,N_7128,N_6099);
nand U11465 (N_11465,N_7513,N_7491);
and U11466 (N_11466,N_4724,N_6369);
or U11467 (N_11467,N_5555,N_7035);
nand U11468 (N_11468,N_7555,N_6647);
nand U11469 (N_11469,N_7022,N_5522);
nand U11470 (N_11470,N_7832,N_7384);
and U11471 (N_11471,N_4750,N_5536);
or U11472 (N_11472,N_4775,N_5236);
xor U11473 (N_11473,N_5594,N_6985);
and U11474 (N_11474,N_7972,N_5001);
nor U11475 (N_11475,N_7346,N_7396);
nor U11476 (N_11476,N_7231,N_7810);
or U11477 (N_11477,N_4147,N_4561);
xnor U11478 (N_11478,N_6106,N_4062);
or U11479 (N_11479,N_6518,N_7550);
xnor U11480 (N_11480,N_7515,N_6040);
and U11481 (N_11481,N_5866,N_4072);
xor U11482 (N_11482,N_7124,N_5143);
nand U11483 (N_11483,N_4775,N_6851);
xor U11484 (N_11484,N_5551,N_6199);
nand U11485 (N_11485,N_7172,N_7310);
and U11486 (N_11486,N_5142,N_7857);
and U11487 (N_11487,N_4359,N_4196);
xnor U11488 (N_11488,N_4992,N_6181);
nor U11489 (N_11489,N_7225,N_7041);
nand U11490 (N_11490,N_7840,N_7266);
and U11491 (N_11491,N_7709,N_7185);
nor U11492 (N_11492,N_4351,N_5098);
and U11493 (N_11493,N_4631,N_6255);
and U11494 (N_11494,N_4927,N_4461);
or U11495 (N_11495,N_5820,N_6506);
xor U11496 (N_11496,N_4020,N_5052);
xnor U11497 (N_11497,N_6195,N_4300);
or U11498 (N_11498,N_6309,N_7493);
or U11499 (N_11499,N_6691,N_7178);
and U11500 (N_11500,N_6660,N_6922);
nand U11501 (N_11501,N_5559,N_7062);
nor U11502 (N_11502,N_7334,N_4443);
xor U11503 (N_11503,N_7808,N_7867);
or U11504 (N_11504,N_6941,N_6690);
nor U11505 (N_11505,N_6634,N_7261);
xnor U11506 (N_11506,N_5092,N_7638);
xor U11507 (N_11507,N_6307,N_5971);
xnor U11508 (N_11508,N_7521,N_7784);
xnor U11509 (N_11509,N_7532,N_6892);
nand U11510 (N_11510,N_7390,N_5853);
nand U11511 (N_11511,N_4050,N_5292);
nand U11512 (N_11512,N_7604,N_5626);
or U11513 (N_11513,N_5982,N_6481);
or U11514 (N_11514,N_5601,N_6792);
nand U11515 (N_11515,N_5471,N_6458);
nor U11516 (N_11516,N_7854,N_7991);
and U11517 (N_11517,N_4129,N_5691);
nor U11518 (N_11518,N_5842,N_4661);
xor U11519 (N_11519,N_4370,N_5165);
xnor U11520 (N_11520,N_4322,N_4406);
or U11521 (N_11521,N_4549,N_6362);
nand U11522 (N_11522,N_7017,N_4187);
nand U11523 (N_11523,N_4782,N_4204);
or U11524 (N_11524,N_6345,N_7789);
and U11525 (N_11525,N_4818,N_6467);
or U11526 (N_11526,N_7336,N_5461);
nand U11527 (N_11527,N_7200,N_5695);
or U11528 (N_11528,N_5699,N_5523);
nor U11529 (N_11529,N_6835,N_7719);
or U11530 (N_11530,N_4014,N_6584);
nor U11531 (N_11531,N_6832,N_6369);
and U11532 (N_11532,N_6965,N_4126);
xnor U11533 (N_11533,N_5591,N_5483);
and U11534 (N_11534,N_4300,N_7664);
nand U11535 (N_11535,N_6919,N_5006);
or U11536 (N_11536,N_5924,N_7928);
xnor U11537 (N_11537,N_4111,N_7524);
nor U11538 (N_11538,N_4138,N_6203);
and U11539 (N_11539,N_4986,N_6211);
nand U11540 (N_11540,N_7526,N_5297);
or U11541 (N_11541,N_6945,N_6367);
or U11542 (N_11542,N_5921,N_4063);
nor U11543 (N_11543,N_4053,N_5632);
xnor U11544 (N_11544,N_5551,N_6715);
nand U11545 (N_11545,N_7987,N_4417);
or U11546 (N_11546,N_6089,N_7998);
xor U11547 (N_11547,N_6085,N_7315);
or U11548 (N_11548,N_7847,N_6054);
and U11549 (N_11549,N_5712,N_7247);
or U11550 (N_11550,N_4397,N_5629);
nor U11551 (N_11551,N_7481,N_7131);
or U11552 (N_11552,N_6912,N_4249);
or U11553 (N_11553,N_6696,N_6099);
xnor U11554 (N_11554,N_5153,N_4740);
and U11555 (N_11555,N_7424,N_4094);
xor U11556 (N_11556,N_4335,N_7788);
nand U11557 (N_11557,N_4059,N_7812);
nand U11558 (N_11558,N_6046,N_4142);
xor U11559 (N_11559,N_7838,N_7837);
nand U11560 (N_11560,N_5790,N_7968);
or U11561 (N_11561,N_7805,N_7076);
nor U11562 (N_11562,N_5320,N_4381);
xor U11563 (N_11563,N_5613,N_7418);
nor U11564 (N_11564,N_5798,N_4464);
nand U11565 (N_11565,N_6264,N_7694);
xor U11566 (N_11566,N_7719,N_6911);
and U11567 (N_11567,N_6304,N_7466);
xnor U11568 (N_11568,N_6997,N_6412);
xnor U11569 (N_11569,N_6722,N_6433);
or U11570 (N_11570,N_7019,N_4737);
and U11571 (N_11571,N_7381,N_7824);
nor U11572 (N_11572,N_6303,N_5210);
xnor U11573 (N_11573,N_6611,N_5327);
nand U11574 (N_11574,N_7992,N_4293);
and U11575 (N_11575,N_4664,N_5513);
or U11576 (N_11576,N_4716,N_4845);
nor U11577 (N_11577,N_7759,N_7060);
nor U11578 (N_11578,N_4703,N_6360);
or U11579 (N_11579,N_7574,N_4180);
and U11580 (N_11580,N_4867,N_4785);
nand U11581 (N_11581,N_5892,N_7728);
or U11582 (N_11582,N_7779,N_4209);
nand U11583 (N_11583,N_7573,N_7574);
xor U11584 (N_11584,N_4181,N_5976);
and U11585 (N_11585,N_4586,N_5808);
xnor U11586 (N_11586,N_5636,N_5857);
nor U11587 (N_11587,N_6930,N_7619);
nand U11588 (N_11588,N_5151,N_4514);
nand U11589 (N_11589,N_7709,N_4169);
xor U11590 (N_11590,N_6300,N_6550);
nor U11591 (N_11591,N_4461,N_6832);
nor U11592 (N_11592,N_7850,N_7397);
xor U11593 (N_11593,N_7713,N_5063);
and U11594 (N_11594,N_4130,N_6599);
nor U11595 (N_11595,N_4282,N_5917);
or U11596 (N_11596,N_4120,N_5899);
or U11597 (N_11597,N_7496,N_6781);
and U11598 (N_11598,N_5451,N_5840);
xnor U11599 (N_11599,N_4720,N_7502);
or U11600 (N_11600,N_7392,N_4092);
xor U11601 (N_11601,N_6498,N_7656);
xnor U11602 (N_11602,N_5888,N_6012);
nand U11603 (N_11603,N_4450,N_7671);
nor U11604 (N_11604,N_7900,N_5233);
xnor U11605 (N_11605,N_4862,N_5888);
or U11606 (N_11606,N_5174,N_5979);
xor U11607 (N_11607,N_6230,N_4413);
nand U11608 (N_11608,N_5328,N_5110);
nor U11609 (N_11609,N_5428,N_4827);
xor U11610 (N_11610,N_6436,N_4550);
nor U11611 (N_11611,N_4109,N_5287);
nand U11612 (N_11612,N_7827,N_7347);
xnor U11613 (N_11613,N_5542,N_6346);
nor U11614 (N_11614,N_7111,N_4993);
and U11615 (N_11615,N_4701,N_6038);
nor U11616 (N_11616,N_4387,N_6497);
and U11617 (N_11617,N_7029,N_5452);
nand U11618 (N_11618,N_7875,N_5251);
xor U11619 (N_11619,N_4465,N_6016);
or U11620 (N_11620,N_4711,N_7008);
xor U11621 (N_11621,N_7106,N_5836);
nand U11622 (N_11622,N_7307,N_5603);
or U11623 (N_11623,N_5217,N_5464);
nand U11624 (N_11624,N_7070,N_7341);
or U11625 (N_11625,N_4323,N_4740);
nor U11626 (N_11626,N_7459,N_7521);
nand U11627 (N_11627,N_6792,N_5046);
or U11628 (N_11628,N_6855,N_7402);
nand U11629 (N_11629,N_6983,N_5475);
nor U11630 (N_11630,N_5369,N_6662);
nand U11631 (N_11631,N_4333,N_4387);
and U11632 (N_11632,N_4068,N_6319);
and U11633 (N_11633,N_7090,N_4113);
nor U11634 (N_11634,N_7435,N_6366);
or U11635 (N_11635,N_4417,N_6866);
nor U11636 (N_11636,N_5539,N_7007);
nand U11637 (N_11637,N_6678,N_5916);
xnor U11638 (N_11638,N_6915,N_4302);
nand U11639 (N_11639,N_7951,N_7666);
or U11640 (N_11640,N_4216,N_4127);
nor U11641 (N_11641,N_5527,N_5874);
and U11642 (N_11642,N_7568,N_5349);
nor U11643 (N_11643,N_6159,N_7173);
or U11644 (N_11644,N_5619,N_5300);
or U11645 (N_11645,N_6195,N_7762);
or U11646 (N_11646,N_7158,N_7864);
nor U11647 (N_11647,N_7173,N_5647);
and U11648 (N_11648,N_6003,N_6126);
xnor U11649 (N_11649,N_6398,N_5127);
xnor U11650 (N_11650,N_5200,N_5540);
nand U11651 (N_11651,N_5156,N_6267);
xnor U11652 (N_11652,N_4711,N_7756);
or U11653 (N_11653,N_6919,N_4037);
xnor U11654 (N_11654,N_5198,N_5111);
nand U11655 (N_11655,N_6413,N_6432);
nor U11656 (N_11656,N_6767,N_4739);
xor U11657 (N_11657,N_5714,N_7542);
nand U11658 (N_11658,N_7347,N_6475);
and U11659 (N_11659,N_6811,N_5113);
or U11660 (N_11660,N_6447,N_6775);
or U11661 (N_11661,N_7593,N_6397);
nand U11662 (N_11662,N_7376,N_7659);
xor U11663 (N_11663,N_5770,N_7435);
or U11664 (N_11664,N_7709,N_6025);
nand U11665 (N_11665,N_6490,N_7577);
nand U11666 (N_11666,N_5348,N_6457);
and U11667 (N_11667,N_4765,N_7670);
nand U11668 (N_11668,N_7338,N_6363);
nor U11669 (N_11669,N_6938,N_6666);
and U11670 (N_11670,N_7538,N_4408);
nand U11671 (N_11671,N_4343,N_4537);
nand U11672 (N_11672,N_5940,N_6110);
nor U11673 (N_11673,N_5886,N_4850);
or U11674 (N_11674,N_4846,N_4791);
or U11675 (N_11675,N_5668,N_4998);
or U11676 (N_11676,N_6339,N_7011);
and U11677 (N_11677,N_7155,N_7289);
or U11678 (N_11678,N_4293,N_7041);
nand U11679 (N_11679,N_6363,N_7059);
or U11680 (N_11680,N_7160,N_6500);
nor U11681 (N_11681,N_7757,N_4923);
xor U11682 (N_11682,N_4398,N_4035);
xnor U11683 (N_11683,N_5052,N_6694);
xnor U11684 (N_11684,N_7936,N_7877);
or U11685 (N_11685,N_6543,N_6096);
or U11686 (N_11686,N_5953,N_6532);
nand U11687 (N_11687,N_4101,N_4150);
xnor U11688 (N_11688,N_7846,N_6974);
nand U11689 (N_11689,N_4344,N_6551);
or U11690 (N_11690,N_6870,N_6630);
nor U11691 (N_11691,N_6264,N_4483);
xnor U11692 (N_11692,N_6756,N_6343);
xor U11693 (N_11693,N_5706,N_5511);
nor U11694 (N_11694,N_7396,N_5883);
nand U11695 (N_11695,N_4300,N_7085);
or U11696 (N_11696,N_4088,N_4684);
and U11697 (N_11697,N_5036,N_6673);
and U11698 (N_11698,N_6409,N_5753);
nand U11699 (N_11699,N_5750,N_4494);
nor U11700 (N_11700,N_6087,N_6875);
or U11701 (N_11701,N_7754,N_6296);
nand U11702 (N_11702,N_7276,N_4038);
xor U11703 (N_11703,N_5261,N_4095);
or U11704 (N_11704,N_7560,N_4034);
nand U11705 (N_11705,N_6357,N_5517);
or U11706 (N_11706,N_5535,N_5227);
nand U11707 (N_11707,N_7169,N_4785);
nor U11708 (N_11708,N_4736,N_5955);
nor U11709 (N_11709,N_5929,N_6041);
or U11710 (N_11710,N_5342,N_6168);
xnor U11711 (N_11711,N_7987,N_6694);
nand U11712 (N_11712,N_4814,N_6741);
and U11713 (N_11713,N_6685,N_4769);
nand U11714 (N_11714,N_5739,N_6135);
nor U11715 (N_11715,N_5320,N_7396);
and U11716 (N_11716,N_6349,N_5601);
xnor U11717 (N_11717,N_6838,N_4417);
nor U11718 (N_11718,N_6896,N_6785);
nor U11719 (N_11719,N_4431,N_7542);
nand U11720 (N_11720,N_5428,N_6818);
nand U11721 (N_11721,N_4178,N_4322);
xor U11722 (N_11722,N_7128,N_5267);
nand U11723 (N_11723,N_6634,N_4302);
and U11724 (N_11724,N_7679,N_5400);
or U11725 (N_11725,N_6266,N_7328);
or U11726 (N_11726,N_6766,N_6294);
nand U11727 (N_11727,N_7170,N_4281);
nand U11728 (N_11728,N_7618,N_6621);
nor U11729 (N_11729,N_6838,N_6905);
nand U11730 (N_11730,N_6621,N_7425);
and U11731 (N_11731,N_5483,N_4604);
and U11732 (N_11732,N_7642,N_5805);
or U11733 (N_11733,N_6760,N_4658);
nand U11734 (N_11734,N_7223,N_5234);
xnor U11735 (N_11735,N_6422,N_6112);
xnor U11736 (N_11736,N_4610,N_5881);
xor U11737 (N_11737,N_6272,N_6405);
nand U11738 (N_11738,N_5594,N_5034);
xnor U11739 (N_11739,N_4520,N_4254);
nor U11740 (N_11740,N_6120,N_5869);
nand U11741 (N_11741,N_5429,N_4518);
xnor U11742 (N_11742,N_6749,N_6325);
or U11743 (N_11743,N_5771,N_5887);
or U11744 (N_11744,N_5256,N_6088);
or U11745 (N_11745,N_4576,N_7469);
and U11746 (N_11746,N_5441,N_7258);
and U11747 (N_11747,N_4619,N_4733);
or U11748 (N_11748,N_6754,N_6614);
and U11749 (N_11749,N_5803,N_7003);
or U11750 (N_11750,N_6011,N_7720);
and U11751 (N_11751,N_6238,N_7241);
nor U11752 (N_11752,N_7660,N_7910);
and U11753 (N_11753,N_4419,N_5400);
nor U11754 (N_11754,N_4598,N_7212);
or U11755 (N_11755,N_4934,N_7425);
xnor U11756 (N_11756,N_5885,N_5789);
and U11757 (N_11757,N_4811,N_7829);
xnor U11758 (N_11758,N_7654,N_4626);
nor U11759 (N_11759,N_4330,N_6642);
nand U11760 (N_11760,N_7424,N_6870);
or U11761 (N_11761,N_6731,N_6436);
and U11762 (N_11762,N_7565,N_6896);
nand U11763 (N_11763,N_6982,N_5030);
nand U11764 (N_11764,N_4775,N_7763);
or U11765 (N_11765,N_6678,N_4037);
xor U11766 (N_11766,N_6496,N_5903);
nor U11767 (N_11767,N_5421,N_4846);
or U11768 (N_11768,N_7426,N_5232);
or U11769 (N_11769,N_5994,N_6005);
nor U11770 (N_11770,N_7823,N_4533);
nor U11771 (N_11771,N_6311,N_5955);
or U11772 (N_11772,N_5752,N_5813);
xor U11773 (N_11773,N_4639,N_4720);
xnor U11774 (N_11774,N_7015,N_7774);
nand U11775 (N_11775,N_5882,N_6440);
nor U11776 (N_11776,N_7026,N_5242);
xor U11777 (N_11777,N_5050,N_5706);
nand U11778 (N_11778,N_5046,N_7291);
xnor U11779 (N_11779,N_7778,N_7034);
or U11780 (N_11780,N_4838,N_7184);
or U11781 (N_11781,N_4174,N_6292);
nor U11782 (N_11782,N_4537,N_5948);
or U11783 (N_11783,N_4694,N_5117);
or U11784 (N_11784,N_6518,N_4785);
xnor U11785 (N_11785,N_6610,N_7642);
or U11786 (N_11786,N_7239,N_7783);
and U11787 (N_11787,N_5114,N_6506);
xor U11788 (N_11788,N_7505,N_5328);
or U11789 (N_11789,N_6070,N_7922);
nand U11790 (N_11790,N_7261,N_5805);
xnor U11791 (N_11791,N_7939,N_7422);
xor U11792 (N_11792,N_4856,N_5901);
xor U11793 (N_11793,N_4082,N_5562);
or U11794 (N_11794,N_7962,N_6393);
nand U11795 (N_11795,N_4008,N_4687);
xnor U11796 (N_11796,N_6334,N_4112);
nand U11797 (N_11797,N_6786,N_5908);
nor U11798 (N_11798,N_5060,N_5944);
and U11799 (N_11799,N_7685,N_7824);
nor U11800 (N_11800,N_4047,N_4685);
and U11801 (N_11801,N_5846,N_5752);
or U11802 (N_11802,N_5491,N_4213);
nor U11803 (N_11803,N_6062,N_5077);
or U11804 (N_11804,N_7506,N_7841);
xnor U11805 (N_11805,N_6906,N_5870);
or U11806 (N_11806,N_7701,N_6739);
or U11807 (N_11807,N_5530,N_6680);
nor U11808 (N_11808,N_4858,N_5561);
or U11809 (N_11809,N_5469,N_7514);
nand U11810 (N_11810,N_7081,N_7529);
nor U11811 (N_11811,N_7946,N_6839);
nor U11812 (N_11812,N_6013,N_6383);
nor U11813 (N_11813,N_7260,N_4681);
or U11814 (N_11814,N_6536,N_4565);
xor U11815 (N_11815,N_7448,N_5063);
nand U11816 (N_11816,N_5113,N_6927);
or U11817 (N_11817,N_6024,N_6542);
nor U11818 (N_11818,N_5062,N_7007);
nand U11819 (N_11819,N_7266,N_6431);
and U11820 (N_11820,N_4430,N_5212);
or U11821 (N_11821,N_6550,N_4894);
xor U11822 (N_11822,N_7072,N_4198);
xnor U11823 (N_11823,N_7141,N_7638);
and U11824 (N_11824,N_5669,N_5278);
and U11825 (N_11825,N_5364,N_4016);
and U11826 (N_11826,N_7478,N_4929);
nor U11827 (N_11827,N_4577,N_5988);
nand U11828 (N_11828,N_5156,N_6600);
xnor U11829 (N_11829,N_7857,N_7527);
nor U11830 (N_11830,N_5234,N_6479);
xnor U11831 (N_11831,N_5997,N_7128);
nor U11832 (N_11832,N_7121,N_5393);
xnor U11833 (N_11833,N_6062,N_4904);
xnor U11834 (N_11834,N_5491,N_4813);
and U11835 (N_11835,N_4050,N_7632);
or U11836 (N_11836,N_4305,N_7530);
nor U11837 (N_11837,N_4929,N_4863);
or U11838 (N_11838,N_5331,N_5522);
nor U11839 (N_11839,N_7912,N_7646);
xor U11840 (N_11840,N_5078,N_4964);
nand U11841 (N_11841,N_6690,N_4742);
and U11842 (N_11842,N_7388,N_4854);
xnor U11843 (N_11843,N_7876,N_5436);
and U11844 (N_11844,N_4146,N_6770);
and U11845 (N_11845,N_4943,N_7290);
nand U11846 (N_11846,N_7874,N_4199);
nand U11847 (N_11847,N_5144,N_5699);
xor U11848 (N_11848,N_5326,N_6080);
and U11849 (N_11849,N_7250,N_7000);
xnor U11850 (N_11850,N_7628,N_6842);
xor U11851 (N_11851,N_5814,N_5576);
xor U11852 (N_11852,N_5744,N_5513);
xnor U11853 (N_11853,N_6521,N_7995);
or U11854 (N_11854,N_5156,N_4361);
and U11855 (N_11855,N_6657,N_7288);
and U11856 (N_11856,N_7871,N_4031);
xnor U11857 (N_11857,N_6187,N_4693);
nand U11858 (N_11858,N_5339,N_7861);
nor U11859 (N_11859,N_6446,N_7256);
nor U11860 (N_11860,N_5343,N_4907);
nand U11861 (N_11861,N_6887,N_7933);
xnor U11862 (N_11862,N_5119,N_4262);
xnor U11863 (N_11863,N_6266,N_7944);
nor U11864 (N_11864,N_7622,N_7993);
nand U11865 (N_11865,N_6612,N_4574);
nor U11866 (N_11866,N_4538,N_4147);
nand U11867 (N_11867,N_4165,N_6799);
and U11868 (N_11868,N_4390,N_6694);
and U11869 (N_11869,N_6323,N_5390);
or U11870 (N_11870,N_6583,N_7048);
nor U11871 (N_11871,N_7876,N_7190);
nor U11872 (N_11872,N_6910,N_7657);
nor U11873 (N_11873,N_4038,N_4569);
nor U11874 (N_11874,N_5965,N_6981);
xnor U11875 (N_11875,N_7211,N_5123);
nor U11876 (N_11876,N_7177,N_6624);
nor U11877 (N_11877,N_6203,N_5905);
or U11878 (N_11878,N_4274,N_7900);
nor U11879 (N_11879,N_6467,N_7574);
nor U11880 (N_11880,N_5372,N_5457);
nand U11881 (N_11881,N_5310,N_6780);
and U11882 (N_11882,N_5746,N_4288);
nor U11883 (N_11883,N_5504,N_5755);
nand U11884 (N_11884,N_6576,N_6957);
and U11885 (N_11885,N_5589,N_4768);
and U11886 (N_11886,N_5762,N_5276);
or U11887 (N_11887,N_5944,N_7021);
or U11888 (N_11888,N_7171,N_4152);
or U11889 (N_11889,N_5873,N_7046);
nor U11890 (N_11890,N_6784,N_6386);
nor U11891 (N_11891,N_7273,N_4284);
xnor U11892 (N_11892,N_7763,N_7135);
nor U11893 (N_11893,N_4628,N_5648);
or U11894 (N_11894,N_4367,N_6462);
and U11895 (N_11895,N_4726,N_4403);
nor U11896 (N_11896,N_6990,N_4258);
nor U11897 (N_11897,N_5325,N_5301);
nor U11898 (N_11898,N_7381,N_7902);
or U11899 (N_11899,N_6137,N_4719);
or U11900 (N_11900,N_7439,N_4283);
nand U11901 (N_11901,N_5210,N_6282);
or U11902 (N_11902,N_6519,N_6966);
or U11903 (N_11903,N_7026,N_7968);
nand U11904 (N_11904,N_4141,N_5161);
xnor U11905 (N_11905,N_4616,N_4472);
and U11906 (N_11906,N_5531,N_7405);
xor U11907 (N_11907,N_7388,N_4167);
or U11908 (N_11908,N_4166,N_7722);
nor U11909 (N_11909,N_6788,N_4984);
and U11910 (N_11910,N_4622,N_7735);
or U11911 (N_11911,N_5107,N_4256);
xnor U11912 (N_11912,N_6968,N_5896);
or U11913 (N_11913,N_5333,N_7402);
nor U11914 (N_11914,N_4705,N_4632);
and U11915 (N_11915,N_6914,N_7641);
xnor U11916 (N_11916,N_4874,N_6522);
nor U11917 (N_11917,N_7214,N_5824);
nand U11918 (N_11918,N_5063,N_4961);
nand U11919 (N_11919,N_6971,N_5498);
nor U11920 (N_11920,N_4866,N_5284);
or U11921 (N_11921,N_5795,N_5418);
xor U11922 (N_11922,N_6075,N_4104);
nor U11923 (N_11923,N_6494,N_5427);
nand U11924 (N_11924,N_4773,N_6218);
and U11925 (N_11925,N_4467,N_4856);
xnor U11926 (N_11926,N_4770,N_5003);
nand U11927 (N_11927,N_6907,N_4566);
nand U11928 (N_11928,N_7972,N_5621);
and U11929 (N_11929,N_7201,N_7948);
and U11930 (N_11930,N_6871,N_4784);
or U11931 (N_11931,N_7071,N_5965);
xnor U11932 (N_11932,N_7046,N_4153);
and U11933 (N_11933,N_5510,N_5960);
or U11934 (N_11934,N_4240,N_6897);
nand U11935 (N_11935,N_4545,N_6789);
xnor U11936 (N_11936,N_6252,N_5568);
nor U11937 (N_11937,N_7156,N_4846);
and U11938 (N_11938,N_5987,N_7623);
nand U11939 (N_11939,N_5049,N_5806);
xor U11940 (N_11940,N_4373,N_6016);
nand U11941 (N_11941,N_4643,N_4454);
and U11942 (N_11942,N_4026,N_5060);
nor U11943 (N_11943,N_6001,N_4920);
nor U11944 (N_11944,N_5096,N_4507);
nor U11945 (N_11945,N_6196,N_7236);
or U11946 (N_11946,N_5511,N_4957);
or U11947 (N_11947,N_6921,N_5795);
xor U11948 (N_11948,N_6353,N_7564);
nand U11949 (N_11949,N_4243,N_6526);
nor U11950 (N_11950,N_6737,N_6465);
nor U11951 (N_11951,N_6354,N_7325);
or U11952 (N_11952,N_4301,N_5401);
xor U11953 (N_11953,N_4018,N_6587);
nor U11954 (N_11954,N_6535,N_4351);
xnor U11955 (N_11955,N_4994,N_7258);
nor U11956 (N_11956,N_6113,N_5062);
or U11957 (N_11957,N_4196,N_7343);
or U11958 (N_11958,N_7026,N_7325);
xor U11959 (N_11959,N_6995,N_6753);
nand U11960 (N_11960,N_5827,N_6921);
nor U11961 (N_11961,N_6530,N_6971);
xnor U11962 (N_11962,N_4201,N_5809);
or U11963 (N_11963,N_7291,N_7180);
or U11964 (N_11964,N_4779,N_4310);
or U11965 (N_11965,N_7580,N_5428);
nor U11966 (N_11966,N_5760,N_5841);
or U11967 (N_11967,N_4919,N_6287);
nor U11968 (N_11968,N_4668,N_4376);
nand U11969 (N_11969,N_4354,N_4031);
nor U11970 (N_11970,N_5952,N_5546);
and U11971 (N_11971,N_4289,N_5473);
xnor U11972 (N_11972,N_6670,N_4888);
or U11973 (N_11973,N_6078,N_5460);
xnor U11974 (N_11974,N_7983,N_5554);
and U11975 (N_11975,N_7915,N_5920);
or U11976 (N_11976,N_7165,N_6973);
and U11977 (N_11977,N_6100,N_4457);
nor U11978 (N_11978,N_4336,N_4636);
nor U11979 (N_11979,N_4089,N_6927);
nand U11980 (N_11980,N_7675,N_6601);
nand U11981 (N_11981,N_6911,N_6733);
nor U11982 (N_11982,N_4521,N_6379);
and U11983 (N_11983,N_7277,N_4465);
or U11984 (N_11984,N_7460,N_5292);
xor U11985 (N_11985,N_7759,N_7327);
xor U11986 (N_11986,N_4480,N_7855);
and U11987 (N_11987,N_5442,N_4054);
xnor U11988 (N_11988,N_4643,N_4234);
xnor U11989 (N_11989,N_6715,N_4674);
nor U11990 (N_11990,N_7160,N_6038);
and U11991 (N_11991,N_5379,N_4438);
nor U11992 (N_11992,N_5610,N_4744);
or U11993 (N_11993,N_7216,N_6844);
xnor U11994 (N_11994,N_6282,N_6841);
and U11995 (N_11995,N_4842,N_7232);
and U11996 (N_11996,N_5482,N_4513);
and U11997 (N_11997,N_5403,N_5934);
xor U11998 (N_11998,N_4752,N_7782);
nor U11999 (N_11999,N_4079,N_6653);
or U12000 (N_12000,N_8801,N_10669);
nand U12001 (N_12001,N_11062,N_11628);
nor U12002 (N_12002,N_9377,N_11927);
nand U12003 (N_12003,N_10554,N_10562);
nand U12004 (N_12004,N_10300,N_11100);
and U12005 (N_12005,N_11633,N_8003);
or U12006 (N_12006,N_9644,N_8942);
or U12007 (N_12007,N_8273,N_11460);
xnor U12008 (N_12008,N_9142,N_8720);
nand U12009 (N_12009,N_8282,N_10072);
or U12010 (N_12010,N_10955,N_11138);
nand U12011 (N_12011,N_10149,N_8344);
nand U12012 (N_12012,N_8024,N_8033);
nor U12013 (N_12013,N_10268,N_9060);
nor U12014 (N_12014,N_9482,N_10534);
nand U12015 (N_12015,N_8687,N_9519);
nand U12016 (N_12016,N_10459,N_8046);
or U12017 (N_12017,N_8343,N_9278);
nor U12018 (N_12018,N_11403,N_9096);
and U12019 (N_12019,N_9488,N_11027);
nor U12020 (N_12020,N_11468,N_9921);
or U12021 (N_12021,N_9343,N_10897);
or U12022 (N_12022,N_8658,N_9266);
nand U12023 (N_12023,N_10789,N_8380);
xor U12024 (N_12024,N_10209,N_10707);
nand U12025 (N_12025,N_8618,N_11083);
or U12026 (N_12026,N_11706,N_8692);
xnor U12027 (N_12027,N_10423,N_8679);
and U12028 (N_12028,N_10478,N_11840);
nand U12029 (N_12029,N_8596,N_8021);
nand U12030 (N_12030,N_10768,N_9734);
or U12031 (N_12031,N_8504,N_8394);
or U12032 (N_12032,N_10041,N_9535);
nor U12033 (N_12033,N_9677,N_8850);
nand U12034 (N_12034,N_8253,N_10689);
or U12035 (N_12035,N_11408,N_11570);
nand U12036 (N_12036,N_10801,N_9688);
xor U12037 (N_12037,N_10227,N_8385);
xor U12038 (N_12038,N_8861,N_8249);
or U12039 (N_12039,N_8075,N_9848);
nor U12040 (N_12040,N_11187,N_9703);
or U12041 (N_12041,N_11447,N_9822);
and U12042 (N_12042,N_9505,N_9107);
and U12043 (N_12043,N_11026,N_9575);
nor U12044 (N_12044,N_11907,N_9083);
nor U12045 (N_12045,N_9379,N_11271);
xor U12046 (N_12046,N_9296,N_9633);
and U12047 (N_12047,N_10463,N_8613);
nand U12048 (N_12048,N_10568,N_8925);
nor U12049 (N_12049,N_8510,N_11631);
and U12050 (N_12050,N_8152,N_11462);
nor U12051 (N_12051,N_10857,N_9075);
xnor U12052 (N_12052,N_8659,N_8677);
nor U12053 (N_12053,N_9156,N_8774);
xor U12054 (N_12054,N_9857,N_10754);
and U12055 (N_12055,N_11801,N_10238);
nand U12056 (N_12056,N_9784,N_10296);
or U12057 (N_12057,N_11317,N_11134);
and U12058 (N_12058,N_11194,N_8970);
and U12059 (N_12059,N_10825,N_10861);
and U12060 (N_12060,N_11803,N_10087);
nand U12061 (N_12061,N_9346,N_10661);
xor U12062 (N_12062,N_10059,N_8633);
xor U12063 (N_12063,N_10682,N_10543);
or U12064 (N_12064,N_11791,N_10582);
nor U12065 (N_12065,N_8845,N_11510);
nand U12066 (N_12066,N_10908,N_11857);
and U12067 (N_12067,N_10623,N_10635);
xor U12068 (N_12068,N_8146,N_10926);
xor U12069 (N_12069,N_10721,N_8975);
xnor U12070 (N_12070,N_10921,N_9972);
and U12071 (N_12071,N_8827,N_11144);
nor U12072 (N_12072,N_11133,N_10678);
and U12073 (N_12073,N_11367,N_10931);
and U12074 (N_12074,N_11389,N_8560);
nor U12075 (N_12075,N_10972,N_10406);
or U12076 (N_12076,N_10605,N_10697);
nand U12077 (N_12077,N_11395,N_11917);
nand U12078 (N_12078,N_10984,N_9390);
and U12079 (N_12079,N_9173,N_11061);
nor U12080 (N_12080,N_11797,N_11856);
xor U12081 (N_12081,N_9255,N_11048);
or U12082 (N_12082,N_9963,N_11418);
nand U12083 (N_12083,N_9120,N_9329);
xor U12084 (N_12084,N_11357,N_9995);
and U12085 (N_12085,N_9757,N_11988);
or U12086 (N_12086,N_11701,N_10276);
and U12087 (N_12087,N_11452,N_9418);
nand U12088 (N_12088,N_11627,N_8668);
nand U12089 (N_12089,N_11214,N_9154);
nand U12090 (N_12090,N_10853,N_11788);
xor U12091 (N_12091,N_8214,N_11198);
nor U12092 (N_12092,N_11255,N_8911);
or U12093 (N_12093,N_11672,N_8290);
and U12094 (N_12094,N_11125,N_9617);
and U12095 (N_12095,N_10080,N_8260);
and U12096 (N_12096,N_11757,N_10540);
nor U12097 (N_12097,N_9686,N_11190);
and U12098 (N_12098,N_11596,N_10819);
xor U12099 (N_12099,N_10654,N_11126);
xor U12100 (N_12100,N_10330,N_11542);
or U12101 (N_12101,N_11912,N_10901);
or U12102 (N_12102,N_9497,N_9594);
xnor U12103 (N_12103,N_11810,N_10672);
and U12104 (N_12104,N_9898,N_9770);
or U12105 (N_12105,N_10085,N_10814);
nand U12106 (N_12106,N_8949,N_10929);
xor U12107 (N_12107,N_11915,N_11305);
and U12108 (N_12108,N_8811,N_9899);
nand U12109 (N_12109,N_9609,N_8795);
nand U12110 (N_12110,N_11943,N_9009);
xnor U12111 (N_12111,N_10128,N_8713);
xor U12112 (N_12112,N_9803,N_8841);
nand U12113 (N_12113,N_11262,N_10660);
xnor U12114 (N_12114,N_8515,N_8370);
nand U12115 (N_12115,N_10992,N_9289);
or U12116 (N_12116,N_9614,N_10140);
and U12117 (N_12117,N_8245,N_11379);
xor U12118 (N_12118,N_9680,N_10407);
nand U12119 (N_12119,N_10860,N_9578);
or U12120 (N_12120,N_11623,N_10737);
nor U12121 (N_12121,N_8113,N_11834);
or U12122 (N_12122,N_8400,N_10551);
and U12123 (N_12123,N_8621,N_8000);
xor U12124 (N_12124,N_8163,N_10420);
nor U12125 (N_12125,N_8413,N_9270);
and U12126 (N_12126,N_11747,N_8788);
nor U12127 (N_12127,N_10442,N_11949);
xnor U12128 (N_12128,N_10160,N_11303);
and U12129 (N_12129,N_11446,N_11240);
nor U12130 (N_12130,N_10448,N_10146);
or U12131 (N_12131,N_11310,N_11783);
xnor U12132 (N_12132,N_8275,N_10791);
xnor U12133 (N_12133,N_8476,N_11975);
and U12134 (N_12134,N_8746,N_9025);
or U12135 (N_12135,N_11899,N_10460);
and U12136 (N_12136,N_9481,N_9068);
nand U12137 (N_12137,N_10638,N_10387);
and U12138 (N_12138,N_8017,N_8660);
nand U12139 (N_12139,N_8092,N_8080);
or U12140 (N_12140,N_9947,N_8629);
xnor U12141 (N_12141,N_9211,N_9542);
and U12142 (N_12142,N_8954,N_10286);
nand U12143 (N_12143,N_9220,N_10105);
or U12144 (N_12144,N_11984,N_11195);
and U12145 (N_12145,N_11977,N_11354);
or U12146 (N_12146,N_9375,N_10077);
xnor U12147 (N_12147,N_9072,N_10915);
nor U12148 (N_12148,N_10251,N_9268);
xor U12149 (N_12149,N_8201,N_8698);
or U12150 (N_12150,N_11171,N_9162);
and U12151 (N_12151,N_11396,N_9619);
and U12152 (N_12152,N_10625,N_9102);
xnor U12153 (N_12153,N_11853,N_8759);
xnor U12154 (N_12154,N_10439,N_9694);
xnor U12155 (N_12155,N_10469,N_11444);
xnor U12156 (N_12156,N_10132,N_10364);
xnor U12157 (N_12157,N_10696,N_9417);
and U12158 (N_12158,N_9664,N_9900);
xnor U12159 (N_12159,N_9217,N_9853);
or U12160 (N_12160,N_8948,N_11843);
xor U12161 (N_12161,N_10928,N_10710);
and U12162 (N_12162,N_11170,N_11934);
xor U12163 (N_12163,N_9565,N_9554);
xnor U12164 (N_12164,N_11050,N_8064);
or U12165 (N_12165,N_8548,N_9082);
or U12166 (N_12166,N_9029,N_11555);
and U12167 (N_12167,N_10662,N_9933);
nand U12168 (N_12168,N_8247,N_10099);
and U12169 (N_12169,N_8611,N_8182);
and U12170 (N_12170,N_11445,N_9378);
and U12171 (N_12171,N_11095,N_11343);
nor U12172 (N_12172,N_8386,N_10020);
and U12173 (N_12173,N_8213,N_9568);
nand U12174 (N_12174,N_10967,N_8234);
and U12175 (N_12175,N_10609,N_8124);
xnor U12176 (N_12176,N_11210,N_8812);
xnor U12177 (N_12177,N_8688,N_8379);
or U12178 (N_12178,N_10254,N_8381);
or U12179 (N_12179,N_10036,N_9733);
nor U12180 (N_12180,N_11252,N_9206);
nor U12181 (N_12181,N_9386,N_10629);
and U12182 (N_12182,N_10771,N_11852);
and U12183 (N_12183,N_8357,N_11192);
or U12184 (N_12184,N_9787,N_8741);
or U12185 (N_12185,N_8019,N_9984);
nand U12186 (N_12186,N_9915,N_11412);
nand U12187 (N_12187,N_9501,N_9732);
xor U12188 (N_12188,N_11495,N_8434);
xor U12189 (N_12189,N_10143,N_8312);
xnor U12190 (N_12190,N_9807,N_9952);
and U12191 (N_12191,N_11093,N_11146);
nor U12192 (N_12192,N_10292,N_8109);
and U12193 (N_12193,N_8155,N_10461);
and U12194 (N_12194,N_9994,N_11320);
and U12195 (N_12195,N_11224,N_8428);
and U12196 (N_12196,N_11835,N_8060);
nand U12197 (N_12197,N_10844,N_11060);
nor U12198 (N_12198,N_9105,N_9618);
or U12199 (N_12199,N_9502,N_10311);
nor U12200 (N_12200,N_9167,N_10436);
or U12201 (N_12201,N_9191,N_9698);
nand U12202 (N_12202,N_11593,N_8545);
or U12203 (N_12203,N_11951,N_9998);
nand U12204 (N_12204,N_8244,N_8221);
or U12205 (N_12205,N_10475,N_9650);
and U12206 (N_12206,N_9786,N_9392);
nand U12207 (N_12207,N_8461,N_10088);
xor U12208 (N_12208,N_10007,N_9610);
xor U12209 (N_12209,N_10224,N_8885);
xnor U12210 (N_12210,N_9456,N_8543);
or U12211 (N_12211,N_9937,N_11941);
or U12212 (N_12212,N_8868,N_9338);
xor U12213 (N_12213,N_11945,N_8009);
xnor U12214 (N_12214,N_8958,N_11331);
and U12215 (N_12215,N_10298,N_8835);
xnor U12216 (N_12216,N_9846,N_9826);
and U12217 (N_12217,N_9422,N_10647);
xnor U12218 (N_12218,N_10148,N_10802);
nand U12219 (N_12219,N_9337,N_9741);
nor U12220 (N_12220,N_8316,N_10904);
and U12221 (N_12221,N_11333,N_10985);
xor U12222 (N_12222,N_9116,N_10242);
xor U12223 (N_12223,N_8297,N_8619);
nand U12224 (N_12224,N_9896,N_9495);
nand U12225 (N_12225,N_10177,N_11417);
nand U12226 (N_12226,N_10025,N_10004);
xnor U12227 (N_12227,N_11457,N_10206);
nor U12228 (N_12228,N_11286,N_9978);
or U12229 (N_12229,N_9226,N_10550);
nor U12230 (N_12230,N_10376,N_9180);
nand U12231 (N_12231,N_9288,N_9553);
nand U12232 (N_12232,N_11487,N_9150);
or U12233 (N_12233,N_11830,N_8578);
and U12234 (N_12234,N_8765,N_8976);
nand U12235 (N_12235,N_11115,N_10966);
and U12236 (N_12236,N_8036,N_11266);
and U12237 (N_12237,N_9945,N_11731);
nand U12238 (N_12238,N_11157,N_8410);
nand U12239 (N_12239,N_10455,N_10161);
nand U12240 (N_12240,N_10103,N_11324);
nand U12241 (N_12241,N_9508,N_8709);
nor U12242 (N_12242,N_9484,N_9074);
nor U12243 (N_12243,N_9325,N_10715);
nand U12244 (N_12244,N_11361,N_10846);
nor U12245 (N_12245,N_10917,N_9717);
nor U12246 (N_12246,N_9696,N_8294);
and U12247 (N_12247,N_9611,N_9547);
nand U12248 (N_12248,N_9756,N_9451);
and U12249 (N_12249,N_8797,N_10441);
nor U12250 (N_12250,N_10450,N_10750);
xnor U12251 (N_12251,N_11568,N_9317);
nand U12252 (N_12252,N_8169,N_11787);
and U12253 (N_12253,N_8206,N_11537);
and U12254 (N_12254,N_10354,N_8541);
nor U12255 (N_12255,N_11557,N_9636);
nor U12256 (N_12256,N_11287,N_11616);
or U12257 (N_12257,N_8291,N_10485);
xor U12258 (N_12258,N_10916,N_9605);
nand U12259 (N_12259,N_9870,N_11072);
xnor U12260 (N_12260,N_10282,N_8646);
or U12261 (N_12261,N_11066,N_9111);
and U12262 (N_12262,N_11229,N_11097);
or U12263 (N_12263,N_11993,N_8027);
nor U12264 (N_12264,N_11328,N_8965);
nand U12265 (N_12265,N_8779,N_11879);
xor U12266 (N_12266,N_9023,N_11275);
and U12267 (N_12267,N_10070,N_11531);
nand U12268 (N_12268,N_10333,N_10365);
nor U12269 (N_12269,N_8023,N_9174);
xnor U12270 (N_12270,N_11521,N_10872);
or U12271 (N_12271,N_10351,N_10604);
or U12272 (N_12272,N_11520,N_8278);
or U12273 (N_12273,N_8893,N_10892);
nor U12274 (N_12274,N_8743,N_9880);
and U12275 (N_12275,N_9960,N_8956);
nor U12276 (N_12276,N_10449,N_9308);
nor U12277 (N_12277,N_11663,N_11442);
nor U12278 (N_12278,N_11349,N_8389);
or U12279 (N_12279,N_11360,N_11903);
nand U12280 (N_12280,N_11878,N_9799);
and U12281 (N_12281,N_8753,N_11792);
nor U12282 (N_12282,N_9719,N_9052);
xnor U12283 (N_12283,N_8849,N_8922);
or U12284 (N_12284,N_8934,N_10862);
nor U12285 (N_12285,N_11505,N_9195);
or U12286 (N_12286,N_10795,N_8286);
nand U12287 (N_12287,N_8558,N_8448);
and U12288 (N_12288,N_8160,N_9510);
or U12289 (N_12289,N_11178,N_9890);
or U12290 (N_12290,N_9975,N_11676);
or U12291 (N_12291,N_9118,N_9967);
and U12292 (N_12292,N_9494,N_11765);
or U12293 (N_12293,N_11599,N_11164);
or U12294 (N_12294,N_9835,N_8396);
nor U12295 (N_12295,N_11067,N_9948);
and U12296 (N_12296,N_8222,N_11109);
xor U12297 (N_12297,N_9672,N_10035);
nand U12298 (N_12298,N_8284,N_11696);
nand U12299 (N_12299,N_11786,N_8772);
nand U12300 (N_12300,N_10272,N_11148);
and U12301 (N_12301,N_10769,N_11808);
xor U12302 (N_12302,N_9475,N_11269);
xnor U12303 (N_12303,N_8997,N_11433);
and U12304 (N_12304,N_11506,N_8905);
or U12305 (N_12305,N_8988,N_9403);
xor U12306 (N_12306,N_9916,N_11486);
nand U12307 (N_12307,N_8355,N_9269);
or U12308 (N_12308,N_11575,N_10338);
and U12309 (N_12309,N_9743,N_9991);
nand U12310 (N_12310,N_8866,N_8580);
nor U12311 (N_12311,N_10889,N_8289);
xnor U12312 (N_12312,N_10782,N_10060);
nand U12313 (N_12313,N_9586,N_8083);
or U12314 (N_12314,N_11390,N_10842);
nor U12315 (N_12315,N_11166,N_11959);
nor U12316 (N_12316,N_8590,N_8963);
nand U12317 (N_12317,N_9716,N_10038);
and U12318 (N_12318,N_10044,N_9398);
xor U12319 (N_12319,N_10001,N_9791);
and U12320 (N_12320,N_9059,N_8823);
xnor U12321 (N_12321,N_10367,N_11260);
or U12322 (N_12322,N_11637,N_11400);
nand U12323 (N_12323,N_10111,N_10528);
or U12324 (N_12324,N_11074,N_10850);
xnor U12325 (N_12325,N_9094,N_11587);
or U12326 (N_12326,N_11176,N_11458);
nand U12327 (N_12327,N_11896,N_9276);
nand U12328 (N_12328,N_11319,N_8681);
or U12329 (N_12329,N_11113,N_11140);
xnor U12330 (N_12330,N_10776,N_8585);
nand U12331 (N_12331,N_11848,N_11244);
and U12332 (N_12332,N_8393,N_10040);
or U12333 (N_12333,N_9530,N_8451);
nand U12334 (N_12334,N_9902,N_8650);
xnor U12335 (N_12335,N_10307,N_10773);
xnor U12336 (N_12336,N_11450,N_9834);
nor U12337 (N_12337,N_8130,N_10095);
nor U12338 (N_12338,N_9368,N_9792);
nand U12339 (N_12339,N_10980,N_11997);
and U12340 (N_12340,N_8272,N_9969);
and U12341 (N_12341,N_9265,N_8601);
xnor U12342 (N_12342,N_10462,N_9907);
nor U12343 (N_12343,N_10948,N_9360);
nor U12344 (N_12344,N_8239,N_10610);
or U12345 (N_12345,N_8862,N_10358);
xor U12346 (N_12346,N_10526,N_11182);
and U12347 (N_12347,N_9958,N_9012);
and U12348 (N_12348,N_8460,N_9005);
nor U12349 (N_12349,N_10233,N_8199);
xnor U12350 (N_12350,N_8492,N_8360);
nor U12351 (N_12351,N_9628,N_8517);
nand U12352 (N_12352,N_11092,N_9333);
nand U12353 (N_12353,N_8856,N_11184);
and U12354 (N_12354,N_8215,N_9942);
xnor U12355 (N_12355,N_10123,N_8656);
nor U12356 (N_12356,N_11010,N_10433);
xnor U12357 (N_12357,N_10626,N_10071);
and U12358 (N_12358,N_9097,N_10440);
nand U12359 (N_12359,N_11529,N_8441);
xnor U12360 (N_12360,N_10685,N_11274);
and U12361 (N_12361,N_10936,N_11035);
nor U12362 (N_12362,N_11130,N_10404);
or U12363 (N_12363,N_10642,N_11985);
and U12364 (N_12364,N_10285,N_9349);
nand U12365 (N_12365,N_8531,N_11567);
and U12366 (N_12366,N_11365,N_9992);
nor U12367 (N_12367,N_9877,N_10775);
nor U12368 (N_12368,N_10848,N_9175);
nor U12369 (N_12369,N_11987,N_9558);
and U12370 (N_12370,N_9491,N_9539);
xnor U12371 (N_12371,N_11090,N_8755);
nand U12372 (N_12372,N_11401,N_9305);
nor U12373 (N_12373,N_9421,N_11370);
or U12374 (N_12374,N_10016,N_10878);
or U12375 (N_12375,N_9122,N_11494);
and U12376 (N_12376,N_10246,N_11105);
nand U12377 (N_12377,N_10067,N_9630);
nand U12378 (N_12378,N_8686,N_10632);
nand U12379 (N_12379,N_10480,N_9626);
nand U12380 (N_12380,N_11006,N_11029);
nor U12381 (N_12381,N_11872,N_9040);
and U12382 (N_12382,N_9085,N_10633);
nand U12383 (N_12383,N_9436,N_8847);
and U12384 (N_12384,N_9706,N_9742);
xor U12385 (N_12385,N_8595,N_9204);
nand U12386 (N_12386,N_9241,N_9013);
nand U12387 (N_12387,N_11267,N_11315);
nand U12388 (N_12388,N_9767,N_11895);
or U12389 (N_12389,N_10882,N_9016);
xor U12390 (N_12390,N_10294,N_11308);
or U12391 (N_12391,N_10415,N_8354);
xor U12392 (N_12392,N_11761,N_10756);
and U12393 (N_12393,N_8600,N_11102);
or U12394 (N_12394,N_8562,N_11758);
nand U12395 (N_12395,N_10097,N_11764);
or U12396 (N_12396,N_11038,N_11524);
xor U12397 (N_12397,N_10466,N_10347);
xnor U12398 (N_12398,N_11772,N_8261);
xor U12399 (N_12399,N_10797,N_8998);
nor U12400 (N_12400,N_10470,N_11992);
and U12401 (N_12401,N_9215,N_11558);
and U12402 (N_12402,N_11366,N_11338);
nor U12403 (N_12403,N_9393,N_11776);
nor U12404 (N_12404,N_8884,N_10708);
nand U12405 (N_12405,N_9882,N_10956);
xnor U12406 (N_12406,N_9312,N_8513);
nor U12407 (N_12407,N_11394,N_8615);
and U12408 (N_12408,N_11173,N_9034);
and U12409 (N_12409,N_10947,N_11629);
and U12410 (N_12410,N_11384,N_11768);
xor U12411 (N_12411,N_11794,N_11953);
nand U12412 (N_12412,N_10890,N_11159);
xnor U12413 (N_12413,N_10836,N_9026);
xor U12414 (N_12414,N_9261,N_8156);
nand U12415 (N_12415,N_8143,N_8346);
and U12416 (N_12416,N_11238,N_9897);
xnor U12417 (N_12417,N_10509,N_8194);
xnor U12418 (N_12418,N_11250,N_9738);
nand U12419 (N_12419,N_11527,N_9090);
xor U12420 (N_12420,N_8511,N_11024);
or U12421 (N_12421,N_8931,N_11737);
and U12422 (N_12422,N_11265,N_9214);
nor U12423 (N_12423,N_9621,N_9997);
nor U12424 (N_12424,N_11534,N_9950);
xor U12425 (N_12425,N_9449,N_9182);
nor U12426 (N_12426,N_9509,N_9582);
and U12427 (N_12427,N_10288,N_8821);
or U12428 (N_12428,N_10187,N_8906);
xnor U12429 (N_12429,N_10614,N_9273);
xnor U12430 (N_12430,N_9177,N_8702);
and U12431 (N_12431,N_8808,N_8056);
and U12432 (N_12432,N_11581,N_11241);
xor U12433 (N_12433,N_8421,N_10377);
or U12434 (N_12434,N_11504,N_8737);
and U12435 (N_12435,N_8736,N_11617);
xor U12436 (N_12436,N_8707,N_8525);
nor U12437 (N_12437,N_8387,N_8154);
nor U12438 (N_12438,N_8010,N_8699);
nor U12439 (N_12439,N_9450,N_10297);
nand U12440 (N_12440,N_10714,N_10817);
or U12441 (N_12441,N_10727,N_10930);
or U12442 (N_12442,N_8121,N_10029);
or U12443 (N_12443,N_11829,N_8719);
and U12444 (N_12444,N_8820,N_10845);
nor U12445 (N_12445,N_10223,N_8614);
nor U12446 (N_12446,N_9710,N_10747);
nor U12447 (N_12447,N_9181,N_8458);
and U12448 (N_12448,N_9341,N_9859);
nor U12449 (N_12449,N_8363,N_8876);
nand U12450 (N_12450,N_9410,N_8890);
xnor U12451 (N_12451,N_8353,N_11604);
nor U12452 (N_12452,N_9336,N_10784);
nand U12453 (N_12453,N_9866,N_11179);
nor U12454 (N_12454,N_10127,N_10217);
or U12455 (N_12455,N_11806,N_9810);
nand U12456 (N_12456,N_8832,N_10028);
nor U12457 (N_12457,N_10345,N_10263);
nor U12458 (N_12458,N_11796,N_9662);
nand U12459 (N_12459,N_10202,N_11422);
or U12460 (N_12460,N_9207,N_9259);
or U12461 (N_12461,N_11656,N_10843);
xnor U12462 (N_12462,N_8077,N_8325);
xor U12463 (N_12463,N_9193,N_8184);
nor U12464 (N_12464,N_9855,N_10849);
nor U12465 (N_12465,N_10113,N_10082);
nand U12466 (N_12466,N_9556,N_11231);
nand U12467 (N_12467,N_10222,N_9458);
or U12468 (N_12468,N_11711,N_11918);
nor U12469 (N_12469,N_9832,N_8824);
and U12470 (N_12470,N_8303,N_9924);
nand U12471 (N_12471,N_11058,N_10116);
xor U12472 (N_12472,N_8809,N_8120);
xor U12473 (N_12473,N_10022,N_11775);
and U12474 (N_12474,N_11847,N_9093);
nand U12475 (N_12475,N_11112,N_11456);
xor U12476 (N_12476,N_10164,N_9223);
nor U12477 (N_12477,N_10675,N_10050);
and U12478 (N_12478,N_10250,N_11259);
nor U12479 (N_12479,N_9399,N_8391);
and U12480 (N_12480,N_9244,N_9697);
or U12481 (N_12481,N_8048,N_11223);
or U12482 (N_12482,N_10018,N_11428);
xnor U12483 (N_12483,N_10374,N_8833);
xor U12484 (N_12484,N_8480,N_11364);
nand U12485 (N_12485,N_8361,N_9340);
nand U12486 (N_12486,N_10884,N_11302);
nand U12487 (N_12487,N_10500,N_11559);
or U12488 (N_12488,N_8414,N_9871);
or U12489 (N_12489,N_9500,N_11968);
xor U12490 (N_12490,N_11948,N_10840);
and U12491 (N_12491,N_10758,N_9764);
or U12492 (N_12492,N_10053,N_9309);
or U12493 (N_12493,N_9382,N_11409);
xor U12494 (N_12494,N_9461,N_8996);
nand U12495 (N_12495,N_8044,N_10738);
nor U12496 (N_12496,N_8701,N_9601);
or U12497 (N_12497,N_8671,N_10361);
nor U12498 (N_12498,N_9641,N_11924);
nand U12499 (N_12499,N_8994,N_10368);
nand U12500 (N_12500,N_9374,N_10946);
xnor U12501 (N_12501,N_8776,N_11831);
or U12502 (N_12502,N_9361,N_11342);
nand U12503 (N_12503,N_11723,N_9161);
nand U12504 (N_12504,N_8170,N_9777);
nand U12505 (N_12505,N_11419,N_11508);
xnor U12506 (N_12506,N_10181,N_11956);
or U12507 (N_12507,N_8445,N_10467);
nor U12508 (N_12508,N_11750,N_11325);
xor U12509 (N_12509,N_8299,N_9649);
and U12510 (N_12510,N_10213,N_8935);
nor U12511 (N_12511,N_8054,N_8773);
xor U12512 (N_12512,N_10389,N_10235);
or U12513 (N_12513,N_9842,N_11769);
xor U12514 (N_12514,N_8235,N_11964);
xor U12515 (N_12515,N_8165,N_8859);
and U12516 (N_12516,N_9858,N_11398);
xnor U12517 (N_12517,N_10665,N_8657);
and U12518 (N_12518,N_10839,N_10229);
or U12519 (N_12519,N_8481,N_11870);
nor U12520 (N_12520,N_10961,N_11128);
nand U12521 (N_12521,N_8676,N_9128);
xnor U12522 (N_12522,N_11222,N_8277);
or U12523 (N_12523,N_8095,N_11785);
and U12524 (N_12524,N_8848,N_11919);
xor U12525 (N_12525,N_11474,N_9811);
nand U12526 (N_12526,N_11978,N_8257);
nor U12527 (N_12527,N_9473,N_10692);
nor U12528 (N_12528,N_8546,N_11429);
and U12529 (N_12529,N_11264,N_10519);
or U12530 (N_12530,N_11018,N_8305);
or U12531 (N_12531,N_8606,N_10011);
nand U12532 (N_12532,N_10739,N_10785);
nor U12533 (N_12533,N_9977,N_10525);
xnor U12534 (N_12534,N_11689,N_8584);
xor U12535 (N_12535,N_9964,N_9380);
nand U12536 (N_12536,N_11290,N_9253);
nand U12537 (N_12537,N_11730,N_8723);
or U12538 (N_12538,N_9454,N_11553);
nor U12539 (N_12539,N_10555,N_10249);
or U12540 (N_12540,N_8536,N_8496);
and U12541 (N_12541,N_11397,N_11845);
and U12542 (N_12542,N_10464,N_8830);
xnor U12543 (N_12543,N_11086,N_10953);
and U12544 (N_12544,N_8384,N_11334);
and U12545 (N_12545,N_11547,N_8961);
nand U12546 (N_12546,N_10107,N_10706);
and U12547 (N_12547,N_8136,N_8116);
or U12548 (N_12548,N_9163,N_10287);
xor U12549 (N_12549,N_10813,N_9247);
or U12550 (N_12550,N_8050,N_10178);
or U12551 (N_12551,N_9236,N_8932);
or U12552 (N_12552,N_9033,N_9302);
nand U12553 (N_12553,N_10987,N_10386);
xnor U12554 (N_12554,N_11432,N_9721);
or U12555 (N_12555,N_8557,N_9304);
nand U12556 (N_12556,N_8509,N_8336);
or U12557 (N_12557,N_10468,N_9541);
or U12558 (N_12558,N_9000,N_10834);
or U12559 (N_12559,N_9047,N_11522);
nand U12560 (N_12560,N_11756,N_10688);
xnor U12561 (N_12561,N_10650,N_8764);
nand U12562 (N_12562,N_9019,N_11549);
nor U12563 (N_12563,N_9754,N_8205);
nor U12564 (N_12564,N_9592,N_11552);
nor U12565 (N_12565,N_11082,N_9965);
and U12566 (N_12566,N_9583,N_9692);
nand U12567 (N_12567,N_9574,N_8452);
and U12568 (N_12568,N_8415,N_8897);
xnor U12569 (N_12569,N_10064,N_9457);
or U12570 (N_12570,N_8258,N_10990);
nor U12571 (N_12571,N_9989,N_11005);
nor U12572 (N_12572,N_9366,N_11002);
nor U12573 (N_12573,N_8020,N_9512);
nand U12574 (N_12574,N_8528,N_10938);
xnor U12575 (N_12575,N_8127,N_11117);
and U12576 (N_12576,N_9318,N_9283);
nand U12577 (N_12577,N_10913,N_8675);
and U12578 (N_12578,N_11132,N_11770);
nand U12579 (N_12579,N_9479,N_8732);
or U12580 (N_12580,N_11634,N_9543);
xor U12581 (N_12581,N_9844,N_8852);
xnor U12582 (N_12582,N_10530,N_11888);
xor U12583 (N_12583,N_10349,N_9232);
and U12584 (N_12584,N_8666,N_10234);
nor U12585 (N_12585,N_11382,N_9735);
nand U12586 (N_12586,N_8062,N_11963);
xnor U12587 (N_12587,N_11391,N_10651);
xor U12588 (N_12588,N_10532,N_8128);
and U12589 (N_12589,N_10106,N_9885);
or U12590 (N_12590,N_11344,N_9426);
and U12591 (N_12591,N_10876,N_8990);
xnor U12592 (N_12592,N_10894,N_10186);
and U12593 (N_12593,N_11213,N_9860);
xnor U12594 (N_12594,N_9936,N_9225);
and U12595 (N_12595,N_10552,N_8899);
xor U12596 (N_12596,N_9091,N_10313);
or U12597 (N_12597,N_10295,N_10541);
or U12598 (N_12598,N_9838,N_8813);
nand U12599 (N_12599,N_9158,N_10165);
nor U12600 (N_12600,N_8814,N_9579);
or U12601 (N_12601,N_10139,N_10870);
and U12602 (N_12602,N_9271,N_11296);
or U12603 (N_12603,N_10763,N_10057);
nand U12604 (N_12604,N_11536,N_10498);
nand U12605 (N_12605,N_9981,N_10606);
and U12606 (N_12606,N_10799,N_9065);
nor U12607 (N_12607,N_11124,N_11864);
xnor U12608 (N_12608,N_9886,N_11261);
nor U12609 (N_12609,N_8800,N_8267);
nor U12610 (N_12610,N_9546,N_9383);
xor U12611 (N_12611,N_11055,N_11332);
xor U12612 (N_12612,N_11154,N_10435);
nand U12613 (N_12613,N_8602,N_9645);
nor U12614 (N_12614,N_8318,N_8315);
xnor U12615 (N_12615,N_10031,N_8691);
and U12616 (N_12616,N_10172,N_9749);
xor U12617 (N_12617,N_9441,N_10950);
nor U12618 (N_12618,N_10400,N_8846);
nor U12619 (N_12619,N_8678,N_9796);
or U12620 (N_12620,N_9808,N_11283);
nand U12621 (N_12621,N_9865,N_11695);
nand U12622 (N_12622,N_11116,N_9058);
or U12623 (N_12623,N_10527,N_11538);
xor U12624 (N_12624,N_10201,N_9196);
nor U12625 (N_12625,N_11920,N_10047);
nand U12626 (N_12626,N_11817,N_8716);
nand U12627 (N_12627,N_9245,N_11185);
or U12628 (N_12628,N_9595,N_9252);
and U12629 (N_12629,N_8901,N_9708);
nor U12630 (N_12630,N_9001,N_9711);
nor U12631 (N_12631,N_11297,N_10410);
or U12632 (N_12632,N_9109,N_10197);
nor U12633 (N_12633,N_11550,N_11322);
and U12634 (N_12634,N_8437,N_10312);
nand U12635 (N_12635,N_9282,N_10228);
nor U12636 (N_12636,N_10275,N_8921);
nor U12637 (N_12637,N_8474,N_9171);
and U12638 (N_12638,N_11571,N_9095);
xor U12639 (N_12639,N_10616,N_10521);
xor U12640 (N_12640,N_8519,N_11685);
xor U12641 (N_12641,N_10216,N_8203);
nor U12642 (N_12642,N_10914,N_8367);
nor U12643 (N_12643,N_10658,N_11386);
and U12644 (N_12644,N_11661,N_11574);
xor U12645 (N_12645,N_11475,N_8626);
nor U12646 (N_12646,N_8424,N_11971);
or U12647 (N_12647,N_9912,N_11209);
or U12648 (N_12648,N_9800,N_9291);
nor U12649 (N_12649,N_10378,N_8376);
xnor U12650 (N_12650,N_9419,N_11602);
or U12651 (N_12651,N_8039,N_11811);
nor U12652 (N_12652,N_8636,N_10594);
or U12653 (N_12653,N_8300,N_11839);
nand U12654 (N_12654,N_8574,N_10879);
nand U12655 (N_12655,N_11678,N_11603);
nor U12656 (N_12656,N_9467,N_9188);
nand U12657 (N_12657,N_11651,N_9227);
nand U12658 (N_12658,N_10155,N_11877);
xnor U12659 (N_12659,N_11659,N_11618);
nor U12660 (N_12660,N_10559,N_8332);
nor U12661 (N_12661,N_8487,N_10253);
nor U12662 (N_12662,N_10900,N_10501);
nand U12663 (N_12663,N_9407,N_10580);
and U12664 (N_12664,N_10393,N_9387);
nand U12665 (N_12665,N_8647,N_10362);
nand U12666 (N_12666,N_9257,N_8964);
nor U12667 (N_12667,N_8125,N_11533);
xnor U12668 (N_12668,N_9514,N_8803);
nand U12669 (N_12669,N_9597,N_8193);
nor U12670 (N_12670,N_8631,N_11782);
and U12671 (N_12671,N_11299,N_8412);
nand U12672 (N_12672,N_10120,N_11608);
and U12673 (N_12673,N_10147,N_10934);
nor U12674 (N_12674,N_8960,N_9761);
or U12675 (N_12675,N_8564,N_11636);
nand U12676 (N_12676,N_9045,N_10200);
and U12677 (N_12677,N_9164,N_11104);
nor U12678 (N_12678,N_10712,N_10150);
and U12679 (N_12679,N_8270,N_10189);
nor U12680 (N_12680,N_9474,N_10002);
nor U12681 (N_12681,N_9608,N_10693);
xnor U12682 (N_12682,N_11193,N_10005);
xnor U12683 (N_12683,N_9246,N_11362);
nor U12684 (N_12684,N_10667,N_8323);
xnor U12685 (N_12685,N_9112,N_8350);
nor U12686 (N_12686,N_9737,N_9203);
nand U12687 (N_12687,N_9311,N_8818);
and U12688 (N_12688,N_11795,N_11045);
or U12689 (N_12689,N_9793,N_9923);
xor U12690 (N_12690,N_10701,N_11800);
nand U12691 (N_12691,N_8750,N_8326);
xnor U12692 (N_12692,N_9993,N_9493);
or U12693 (N_12693,N_11946,N_11515);
nor U12694 (N_12694,N_11858,N_8166);
and U12695 (N_12695,N_10163,N_10680);
and U12696 (N_12696,N_11900,N_9813);
nor U12697 (N_12697,N_11614,N_8628);
and U12698 (N_12698,N_10729,N_11813);
xnor U12699 (N_12699,N_9224,N_8763);
xnor U12700 (N_12700,N_8144,N_9599);
nor U12701 (N_12701,N_10816,N_10649);
or U12702 (N_12702,N_8787,N_9632);
nand U12703 (N_12703,N_11648,N_8188);
nor U12704 (N_12704,N_10355,N_8673);
and U12705 (N_12705,N_8107,N_8034);
xnor U12706 (N_12706,N_8430,N_9462);
nand U12707 (N_12707,N_8173,N_8076);
nor U12708 (N_12708,N_10291,N_10304);
nor U12709 (N_12709,N_11420,N_9205);
or U12710 (N_12710,N_11199,N_10597);
and U12711 (N_12711,N_11610,N_10416);
and U12712 (N_12712,N_11647,N_11497);
and U12713 (N_12713,N_8067,N_8588);
nand U12714 (N_12714,N_9637,N_9080);
nor U12715 (N_12715,N_8609,N_8822);
or U12716 (N_12716,N_10428,N_8926);
xor U12717 (N_12717,N_9759,N_8503);
and U12718 (N_12718,N_11551,N_10671);
xor U12719 (N_12719,N_11556,N_8979);
and U12720 (N_12720,N_10270,N_11991);
nand U12721 (N_12721,N_10166,N_11908);
or U12722 (N_12722,N_10430,N_8212);
nor U12723 (N_12723,N_10537,N_11855);
nor U12724 (N_12724,N_8575,N_11478);
nand U12725 (N_12725,N_11989,N_9179);
and U12726 (N_12726,N_10278,N_10587);
or U12727 (N_12727,N_8223,N_9357);
nor U12728 (N_12728,N_9646,N_10212);
xor U12729 (N_12729,N_9358,N_10506);
xnor U12730 (N_12730,N_8045,N_10944);
and U12731 (N_12731,N_9771,N_9200);
or U12732 (N_12732,N_10772,N_11326);
xnor U12733 (N_12733,N_9856,N_10144);
or U12734 (N_12734,N_8697,N_11799);
or U12735 (N_12735,N_8924,N_9447);
nor U12736 (N_12736,N_8991,N_8655);
nor U12737 (N_12737,N_9388,N_9157);
nor U12738 (N_12738,N_11894,N_11207);
and U12739 (N_12739,N_10989,N_11329);
or U12740 (N_12740,N_9668,N_11339);
nand U12741 (N_12741,N_11047,N_11402);
or U12742 (N_12742,N_8189,N_11854);
xnor U12743 (N_12743,N_8108,N_8532);
xor U12744 (N_12744,N_9593,N_8138);
and U12745 (N_12745,N_11609,N_8368);
xnor U12746 (N_12746,N_8630,N_11704);
or U12747 (N_12747,N_10013,N_10078);
nor U12748 (N_12748,N_8978,N_11205);
or U12749 (N_12749,N_10725,N_9248);
or U12750 (N_12750,N_8047,N_9117);
xor U12751 (N_12751,N_9453,N_10247);
xnor U12752 (N_12752,N_10100,N_10793);
nor U12753 (N_12753,N_11385,N_10949);
nor U12754 (N_12754,N_11824,N_10856);
or U12755 (N_12755,N_10553,N_11675);
nand U12756 (N_12756,N_8274,N_8153);
or U12757 (N_12757,N_10136,N_8625);
and U12758 (N_12758,N_8006,N_8106);
or U12759 (N_12759,N_11172,N_10104);
or U12760 (N_12760,N_11741,N_8190);
nand U12761 (N_12761,N_9854,N_9272);
xor U12762 (N_12762,N_11226,N_10713);
nor U12763 (N_12763,N_9986,N_8623);
nor U12764 (N_12764,N_11720,N_10258);
or U12765 (N_12765,N_8470,N_9103);
or U12766 (N_12766,N_8035,N_9194);
nor U12767 (N_12767,N_11668,N_9141);
nor U12768 (N_12768,N_10910,N_9354);
nand U12769 (N_12769,N_11499,N_8871);
xor U12770 (N_12770,N_8896,N_9166);
and U12771 (N_12771,N_10520,N_9286);
or U12772 (N_12772,N_10348,N_9321);
xor U12773 (N_12773,N_8877,N_8340);
xor U12774 (N_12774,N_9691,N_9262);
xor U12775 (N_12775,N_11073,N_8250);
or U12776 (N_12776,N_8187,N_8456);
nor U12777 (N_12777,N_8420,N_8306);
and U12778 (N_12778,N_9251,N_8241);
nor U12779 (N_12779,N_8292,N_11763);
or U12780 (N_12780,N_11606,N_10684);
and U12781 (N_12781,N_9683,N_11211);
and U12782 (N_12782,N_11077,N_11814);
nand U12783 (N_12783,N_8912,N_9687);
xor U12784 (N_12784,N_11330,N_8112);
nor U12785 (N_12785,N_8887,N_8218);
xor U12786 (N_12786,N_8909,N_11022);
or U12787 (N_12787,N_10852,N_8798);
nor U12788 (N_12788,N_11034,N_10158);
nor U12789 (N_12789,N_11065,N_10267);
nor U12790 (N_12790,N_9218,N_9779);
xnor U12791 (N_12791,N_11930,N_8756);
and U12792 (N_12792,N_9152,N_11191);
nand U12793 (N_12793,N_8168,N_10806);
nand U12794 (N_12794,N_10476,N_11314);
xor U12795 (N_12795,N_11539,N_11511);
nand U12796 (N_12796,N_10301,N_9930);
nor U12797 (N_12797,N_9264,N_10592);
or U12798 (N_12798,N_10741,N_10379);
or U12799 (N_12799,N_9730,N_9805);
xnor U12800 (N_12800,N_11860,N_10248);
and U12801 (N_12801,N_9715,N_11106);
nor U12802 (N_12802,N_11476,N_11519);
and U12803 (N_12803,N_9824,N_8770);
and U12804 (N_12804,N_8603,N_10726);
nand U12805 (N_12805,N_10051,N_11108);
nor U12806 (N_12806,N_10627,N_10920);
or U12807 (N_12807,N_9391,N_11316);
xnor U12808 (N_12808,N_8507,N_10299);
or U12809 (N_12809,N_10655,N_8276);
nor U12810 (N_12810,N_9140,N_9801);
nand U12811 (N_12811,N_9365,N_8141);
nor U12812 (N_12812,N_11425,N_8857);
nor U12813 (N_12813,N_9216,N_8836);
nor U12814 (N_12814,N_11165,N_9699);
or U12815 (N_12815,N_11972,N_8708);
and U12816 (N_12816,N_10743,N_8139);
xnor U12817 (N_12817,N_10119,N_11718);
nand U12818 (N_12818,N_11893,N_9110);
and U12819 (N_12819,N_11023,N_10804);
and U12820 (N_12820,N_8417,N_11158);
nand U12821 (N_12821,N_10831,N_9443);
and U12822 (N_12822,N_10422,N_10774);
xor U12823 (N_12823,N_10975,N_8690);
nand U12824 (N_12824,N_9529,N_8296);
nor U12825 (N_12825,N_9465,N_11111);
nand U12826 (N_12826,N_10512,N_9055);
or U12827 (N_12827,N_10924,N_8936);
nand U12828 (N_12828,N_11649,N_9127);
nand U12829 (N_12829,N_9004,N_10613);
or U12830 (N_12830,N_9100,N_11392);
nor U12831 (N_12831,N_10762,N_8914);
or U12832 (N_12832,N_11143,N_9752);
and U12833 (N_12833,N_10432,N_9788);
and U12834 (N_12834,N_11196,N_9613);
nor U12835 (N_12835,N_11163,N_8374);
nor U12836 (N_12836,N_11300,N_9996);
xor U12837 (N_12837,N_10426,N_10342);
and U12838 (N_12838,N_11020,N_11423);
nor U12839 (N_12839,N_11742,N_8971);
nor U12840 (N_12840,N_10483,N_8771);
nor U12841 (N_12841,N_11543,N_11383);
nand U12842 (N_12842,N_10033,N_10858);
nor U12843 (N_12843,N_11818,N_8878);
xor U12844 (N_12844,N_10009,N_9516);
xnor U12845 (N_12845,N_11019,N_8262);
nor U12846 (N_12846,N_10427,N_11220);
and U12847 (N_12847,N_8640,N_10438);
nand U12848 (N_12848,N_10652,N_9239);
xor U12849 (N_12849,N_10644,N_10000);
xnor U12850 (N_12850,N_10728,N_8538);
or U12851 (N_12851,N_8438,N_8450);
nand U12852 (N_12852,N_8372,N_11561);
xnor U12853 (N_12853,N_9988,N_10830);
and U12854 (N_12854,N_10873,N_11721);
xor U12855 (N_12855,N_9661,N_8442);
and U12856 (N_12856,N_10086,N_9750);
nor U12857 (N_12857,N_8418,N_10593);
or U12858 (N_12858,N_10445,N_11336);
and U12859 (N_12859,N_10765,N_8022);
xnor U12860 (N_12860,N_8320,N_8717);
and U12861 (N_12861,N_10280,N_9620);
nor U12862 (N_12862,N_11639,N_11044);
and U12863 (N_12863,N_8685,N_11348);
and U12864 (N_12864,N_8747,N_9775);
and U12865 (N_12865,N_8745,N_10073);
nor U12866 (N_12866,N_11327,N_8662);
or U12867 (N_12867,N_9657,N_9098);
or U12868 (N_12868,N_9562,N_9929);
nand U12869 (N_12869,N_10335,N_11393);
or U12870 (N_12870,N_9222,N_9159);
or U12871 (N_12871,N_9843,N_11033);
nor U12872 (N_12872,N_9971,N_11625);
xor U12873 (N_12873,N_8680,N_9178);
and U12874 (N_12874,N_11345,N_8117);
nand U12875 (N_12875,N_10939,N_8984);
xnor U12876 (N_12876,N_10927,N_8041);
or U12877 (N_12877,N_11512,N_11355);
and U12878 (N_12878,N_8007,N_11725);
nor U12879 (N_12879,N_9727,N_11523);
or U12880 (N_12880,N_8059,N_10601);
nand U12881 (N_12881,N_10343,N_8775);
and U12882 (N_12882,N_11901,N_9552);
nor U12883 (N_12883,N_8140,N_8683);
xor U12884 (N_12884,N_10244,N_11726);
nor U12885 (N_12885,N_8612,N_8569);
nand U12886 (N_12886,N_10488,N_9201);
xor U12887 (N_12887,N_8865,N_10179);
or U12888 (N_12888,N_9551,N_11217);
xor U12889 (N_12889,N_11576,N_9490);
and U12890 (N_12890,N_8307,N_8159);
and U12891 (N_12891,N_9656,N_9428);
and U12892 (N_12892,N_8178,N_9723);
xor U12893 (N_12893,N_9731,N_9471);
and U12894 (N_12894,N_11640,N_10711);
xor U12895 (N_12895,N_8025,N_10350);
or U12896 (N_12896,N_10999,N_8293);
xnor U12897 (N_12897,N_9638,N_8069);
xor U12898 (N_12898,N_10863,N_11615);
xor U12899 (N_12899,N_9445,N_8648);
nor U12900 (N_12900,N_8335,N_11436);
or U12901 (N_12901,N_8653,N_9518);
or U12902 (N_12902,N_9705,N_11693);
nor U12903 (N_12903,N_9041,N_8134);
nor U12904 (N_12904,N_9381,N_9762);
xor U12905 (N_12905,N_9359,N_9797);
and U12906 (N_12906,N_11754,N_10152);
nand U12907 (N_12907,N_11546,N_10818);
nand U12908 (N_12908,N_8913,N_8313);
and U12909 (N_12909,N_9212,N_10810);
xor U12910 (N_12910,N_8598,N_10993);
nor U12911 (N_12911,N_8843,N_11036);
xnor U12912 (N_12912,N_8181,N_11431);
xnor U12913 (N_12913,N_9024,N_9433);
nor U12914 (N_12914,N_11619,N_11258);
nand U12915 (N_12915,N_8784,N_9483);
nor U12916 (N_12916,N_10369,N_10722);
nand U12917 (N_12917,N_11215,N_8256);
and U12918 (N_12918,N_11740,N_9079);
nor U12919 (N_12919,N_8579,N_10184);
and U12920 (N_12920,N_10066,N_8288);
nor U12921 (N_12921,N_11744,N_11983);
or U12922 (N_12922,N_11218,N_9294);
nor U12923 (N_12923,N_9676,N_9648);
or U12924 (N_12924,N_8957,N_11644);
and U12925 (N_12925,N_10971,N_11174);
nor U12926 (N_12926,N_8339,N_10108);
xor U12927 (N_12927,N_9260,N_9054);
xor U12928 (N_12928,N_8985,N_10363);
and U12929 (N_12929,N_9351,N_9673);
nor U12930 (N_12930,N_11188,N_8542);
xnor U12931 (N_12931,N_8457,N_9463);
or U12932 (N_12932,N_11999,N_8953);
and U12933 (N_12933,N_9307,N_8444);
nand U12934 (N_12934,N_10225,N_9430);
or U12935 (N_12935,N_10643,N_8785);
nor U12936 (N_12936,N_8482,N_8592);
or U12937 (N_12937,N_11586,N_11007);
nand U12938 (N_12938,N_10563,N_9720);
nand U12939 (N_12939,N_8501,N_9913);
nand U12940 (N_12940,N_11986,N_11595);
xnor U12941 (N_12941,N_9536,N_9961);
or U12942 (N_12942,N_8220,N_10912);
nor U12943 (N_12943,N_8137,N_8710);
xnor U12944 (N_12944,N_9424,N_8616);
and U12945 (N_12945,N_10828,N_11594);
or U12946 (N_12946,N_9833,N_8358);
xor U12947 (N_12947,N_8014,N_8087);
nor U12948 (N_12948,N_8524,N_10717);
nor U12949 (N_12949,N_10641,N_8977);
or U12950 (N_12950,N_11844,N_10536);
and U12951 (N_12951,N_10600,N_8583);
or U12952 (N_12952,N_10815,N_11821);
and U12953 (N_12953,N_9342,N_8281);
nand U12954 (N_12954,N_11263,N_10317);
or U12955 (N_12955,N_8469,N_8742);
and U12956 (N_12956,N_8563,N_8030);
and U12957 (N_12957,N_9622,N_11256);
nor U12958 (N_12958,N_8219,N_10231);
xnor U12959 (N_12959,N_11554,N_9598);
xor U12960 (N_12960,N_9078,N_10390);
nor U12961 (N_12961,N_10940,N_11381);
nand U12962 (N_12962,N_10770,N_10023);
nor U12963 (N_12963,N_9520,N_10042);
xor U12964 (N_12964,N_10207,N_9330);
and U12965 (N_12965,N_10723,N_11247);
or U12966 (N_12966,N_11532,N_11954);
nand U12967 (N_12967,N_9088,N_11597);
xnor U12968 (N_12968,N_8094,N_9385);
or U12969 (N_12969,N_8783,N_8903);
or U12970 (N_12970,N_8645,N_11937);
and U12971 (N_12971,N_10173,N_11734);
or U12972 (N_12972,N_11923,N_9751);
nor U12973 (N_12973,N_8390,N_8207);
and U12974 (N_12974,N_8388,N_9790);
nand U12975 (N_12975,N_8377,N_10273);
xnor U12976 (N_12976,N_11642,N_11680);
and U12977 (N_12977,N_9966,N_9922);
or U12978 (N_12978,N_8028,N_10686);
or U12979 (N_12979,N_10193,N_8649);
nor U12980 (N_12980,N_8726,N_8534);
nor U12981 (N_12981,N_8587,N_10063);
nor U12982 (N_12982,N_9533,N_9123);
and U12983 (N_12983,N_8280,N_9957);
and U12984 (N_12984,N_8074,N_11600);
and U12985 (N_12985,N_9667,N_10503);
xnor U12986 (N_12986,N_11098,N_11270);
or U12987 (N_12987,N_8008,N_11114);
or U12988 (N_12988,N_11490,N_11779);
or U12989 (N_12989,N_8466,N_10262);
or U12990 (N_12990,N_9517,N_9655);
or U12991 (N_12991,N_9487,N_10569);
xor U12992 (N_12992,N_11939,N_10510);
xnor U12993 (N_12993,N_8319,N_10308);
xnor U12994 (N_12994,N_8179,N_11588);
or U12995 (N_12995,N_10925,N_9186);
nor U12996 (N_12996,N_9504,N_11753);
nor U12997 (N_12997,N_11724,N_11683);
xor U12998 (N_12998,N_8804,N_10046);
nand U12999 (N_12999,N_11572,N_10677);
nor U13000 (N_13000,N_10578,N_11874);
or U13001 (N_13001,N_8637,N_10375);
or U13002 (N_13002,N_10497,N_10024);
nand U13003 (N_13003,N_11583,N_8927);
nand U13004 (N_13004,N_9316,N_11491);
xnor U13005 (N_13005,N_8635,N_11040);
and U13006 (N_13006,N_11849,N_11237);
or U13007 (N_13007,N_10798,N_8570);
nand U13008 (N_13008,N_9469,N_8266);
nor U13009 (N_13009,N_8485,N_10631);
xor U13010 (N_13010,N_10511,N_11032);
xor U13011 (N_13011,N_11358,N_11046);
or U13012 (N_13012,N_9576,N_8265);
xor U13013 (N_13013,N_11690,N_11996);
nor U13014 (N_13014,N_9658,N_8052);
nor U13015 (N_13015,N_10887,N_11807);
and U13016 (N_13016,N_8467,N_9198);
nand U13017 (N_13017,N_10911,N_10637);
or U13018 (N_13018,N_11716,N_9612);
xor U13019 (N_13019,N_11932,N_9402);
or U13020 (N_13020,N_10360,N_10484);
nand U13021 (N_13021,N_11890,N_9147);
and U13022 (N_13022,N_10006,N_8547);
nor U13023 (N_13023,N_8142,N_9852);
nor U13024 (N_13024,N_11347,N_11043);
and U13025 (N_13025,N_8910,N_11015);
and U13026 (N_13026,N_10102,N_8053);
nand U13027 (N_13027,N_8972,N_9927);
nand U13028 (N_13028,N_8348,N_11921);
nor U13029 (N_13029,N_8255,N_9669);
nand U13030 (N_13030,N_11885,N_9084);
xor U13031 (N_13031,N_11482,N_9039);
and U13032 (N_13032,N_8529,N_8624);
or U13033 (N_13033,N_11748,N_8177);
or U13034 (N_13034,N_9812,N_11103);
xor U13035 (N_13035,N_9460,N_11415);
nor U13036 (N_13036,N_11882,N_10670);
and U13037 (N_13037,N_8695,N_11498);
or U13038 (N_13038,N_8089,N_11202);
nor U13039 (N_13039,N_8566,N_9908);
or U13040 (N_13040,N_10336,N_9567);
nand U13041 (N_13041,N_9132,N_11728);
and U13042 (N_13042,N_10425,N_11732);
and U13043 (N_13043,N_9396,N_8729);
nor U13044 (N_13044,N_9339,N_11825);
nor U13045 (N_13045,N_10185,N_10952);
and U13046 (N_13046,N_8001,N_11012);
nand U13047 (N_13047,N_9032,N_8383);
and U13048 (N_13048,N_10973,N_10564);
xor U13049 (N_13049,N_8351,N_9076);
and U13050 (N_13050,N_8597,N_10402);
xor U13051 (N_13051,N_8475,N_10142);
or U13052 (N_13052,N_11410,N_8724);
or U13053 (N_13053,N_11416,N_10043);
or U13054 (N_13054,N_11502,N_8943);
xor U13055 (N_13055,N_11119,N_11413);
nand U13056 (N_13056,N_8490,N_8392);
nor U13057 (N_13057,N_9679,N_9124);
nand U13058 (N_13058,N_9384,N_8195);
and U13059 (N_13059,N_10443,N_11236);
or U13060 (N_13060,N_11970,N_10603);
or U13061 (N_13061,N_8049,N_9600);
xnor U13062 (N_13062,N_11307,N_11037);
nand U13063 (N_13063,N_9081,N_8228);
or U13064 (N_13064,N_10218,N_11070);
or U13065 (N_13065,N_9755,N_9435);
xnor U13066 (N_13066,N_10780,N_11380);
nand U13067 (N_13067,N_10092,N_8037);
and U13068 (N_13068,N_10465,N_10357);
xor U13069 (N_13069,N_9873,N_9146);
nand U13070 (N_13070,N_11246,N_10724);
xor U13071 (N_13071,N_11933,N_11230);
or U13072 (N_13072,N_8242,N_9663);
nor U13073 (N_13073,N_8617,N_9869);
and U13074 (N_13074,N_11911,N_9439);
or U13075 (N_13075,N_11155,N_8766);
xnor U13076 (N_13076,N_8484,N_9839);
or U13077 (N_13077,N_8860,N_11461);
nand U13078 (N_13078,N_11826,N_9344);
or U13079 (N_13079,N_9753,N_10409);
xor U13080 (N_13080,N_8439,N_9666);
nor U13081 (N_13081,N_8711,N_8012);
nand U13082 (N_13082,N_10869,N_8073);
nor U13083 (N_13083,N_9538,N_11359);
nor U13084 (N_13084,N_10612,N_10683);
or U13085 (N_13085,N_8663,N_10957);
nor U13086 (N_13086,N_8722,N_10145);
nor U13087 (N_13087,N_8435,N_9889);
nor U13088 (N_13088,N_10585,N_11008);
and U13089 (N_13089,N_10787,N_10719);
or U13090 (N_13090,N_9104,N_8641);
or U13091 (N_13091,N_8432,N_8918);
or U13092 (N_13092,N_10052,N_9371);
and U13093 (N_13093,N_11995,N_8553);
xor U13094 (N_13094,N_10691,N_9955);
nor U13095 (N_13095,N_8900,N_8907);
nor U13096 (N_13096,N_10766,N_10502);
nor U13097 (N_13097,N_9370,N_10620);
or U13098 (N_13098,N_10524,N_10855);
nand U13099 (N_13099,N_8454,N_10499);
and U13100 (N_13100,N_8802,N_11674);
xnor U13101 (N_13101,N_8131,N_9279);
nor U13102 (N_13102,N_11094,N_9470);
and U13103 (N_13103,N_10720,N_10960);
nand U13104 (N_13104,N_8639,N_9695);
nand U13105 (N_13105,N_11544,N_10457);
nor U13106 (N_13106,N_9744,N_10491);
and U13107 (N_13107,N_9240,N_9867);
xnor U13108 (N_13108,N_8886,N_9549);
xnor U13109 (N_13109,N_10607,N_8644);
nor U13110 (N_13110,N_11802,N_11545);
nor U13111 (N_13111,N_11735,N_9557);
xnor U13112 (N_13112,N_11011,N_9028);
or U13113 (N_13113,N_9373,N_8967);
or U13114 (N_13114,N_11780,N_9086);
or U13115 (N_13115,N_10114,N_8171);
nor U13116 (N_13116,N_11714,N_9413);
nand U13117 (N_13117,N_9532,N_8705);
and U13118 (N_13118,N_10575,N_11580);
and U13119 (N_13119,N_9176,N_10579);
nand U13120 (N_13120,N_11669,N_8167);
nor U13121 (N_13121,N_8793,N_9724);
nand U13122 (N_13122,N_8593,N_9561);
nand U13123 (N_13123,N_11301,N_8995);
and U13124 (N_13124,N_9021,N_11239);
nand U13125 (N_13125,N_9712,N_9748);
xor U13126 (N_13126,N_10081,N_10583);
nand U13127 (N_13127,N_8149,N_9883);
xor U13128 (N_13128,N_9295,N_10823);
nand U13129 (N_13129,N_8004,N_8883);
nor U13130 (N_13130,N_11657,N_11156);
nand U13131 (N_13131,N_11931,N_10919);
nor U13132 (N_13132,N_10049,N_10690);
xor U13133 (N_13133,N_10545,N_9229);
xnor U13134 (N_13134,N_10126,N_10664);
or U13135 (N_13135,N_8158,N_9414);
or U13136 (N_13136,N_10918,N_8780);
xnor U13137 (N_13137,N_11277,N_8079);
nor U13138 (N_13138,N_9910,N_8129);
and U13139 (N_13139,N_10157,N_9643);
nand U13140 (N_13140,N_8070,N_8086);
and U13141 (N_13141,N_11535,N_8544);
nor U13142 (N_13142,N_11662,N_9604);
nand U13143 (N_13143,N_9531,N_10174);
or U13144 (N_13144,N_10065,N_10056);
xor U13145 (N_13145,N_10284,N_10327);
nor U13146 (N_13146,N_10154,N_9829);
nor U13147 (N_13147,N_10026,N_8940);
nand U13148 (N_13148,N_10833,N_11936);
nor U13149 (N_13149,N_9736,N_11733);
and U13150 (N_13150,N_9943,N_9250);
nand U13151 (N_13151,N_8969,N_9670);
or U13152 (N_13152,N_11405,N_11057);
xnor U13153 (N_13153,N_11118,N_11755);
nor U13154 (N_13154,N_10951,N_9693);
or U13155 (N_13155,N_11208,N_10962);
and U13156 (N_13156,N_8259,N_8211);
or U13157 (N_13157,N_8478,N_10800);
and U13158 (N_13158,N_11658,N_11201);
nand U13159 (N_13159,N_8327,N_9849);
xnor U13160 (N_13160,N_8431,N_11762);
and U13161 (N_13161,N_8522,N_10970);
or U13162 (N_13162,N_8285,N_9409);
and U13163 (N_13163,N_11186,N_10112);
and U13164 (N_13164,N_8917,N_11017);
nand U13165 (N_13165,N_11962,N_10408);
or U13166 (N_13166,N_8817,N_9726);
and U13167 (N_13167,N_9209,N_9878);
nand U13168 (N_13168,N_11664,N_10841);
and U13169 (N_13169,N_9804,N_8436);
or U13170 (N_13170,N_9092,N_11145);
nor U13171 (N_13171,N_9106,N_9763);
or U13172 (N_13172,N_9395,N_10907);
nor U13173 (N_13173,N_8881,N_11592);
or U13174 (N_13174,N_10319,N_11251);
nand U13175 (N_13175,N_10986,N_10230);
nand U13176 (N_13176,N_9234,N_9895);
or U13177 (N_13177,N_9789,N_8301);
or U13178 (N_13178,N_10079,N_9503);
nor U13179 (N_13179,N_11909,N_8689);
xnor U13180 (N_13180,N_8842,N_11980);
or U13181 (N_13181,N_10954,N_9893);
xnor U13182 (N_13182,N_8364,N_9434);
nor U13183 (N_13183,N_8605,N_10820);
nor U13184 (N_13184,N_8892,N_9350);
nor U13185 (N_13185,N_10659,N_11940);
nor U13186 (N_13186,N_9027,N_11085);
and U13187 (N_13187,N_10260,N_8586);
nor U13188 (N_13188,N_9362,N_8864);
or U13189 (N_13189,N_9682,N_8651);
xnor U13190 (N_13190,N_10454,N_10337);
or U13191 (N_13191,N_11692,N_10783);
xnor U13192 (N_13192,N_8568,N_8494);
xor U13193 (N_13193,N_9327,N_8254);
or U13194 (N_13194,N_11850,N_11833);
and U13195 (N_13195,N_9781,N_9782);
and U13196 (N_13196,N_8237,N_8331);
or U13197 (N_13197,N_11150,N_10522);
nand U13198 (N_13198,N_9184,N_10083);
and U13199 (N_13199,N_9652,N_10030);
xor U13200 (N_13200,N_9809,N_9629);
or U13201 (N_13201,N_10544,N_8426);
or U13202 (N_13202,N_10352,N_10208);
nor U13203 (N_13203,N_9326,N_9202);
nand U13204 (N_13204,N_8693,N_8781);
and U13205 (N_13205,N_9903,N_11851);
nand U13206 (N_13206,N_8298,N_9071);
and U13207 (N_13207,N_9564,N_8634);
nor U13208 (N_13208,N_11404,N_10240);
nand U13209 (N_13209,N_10334,N_8499);
or U13210 (N_13210,N_11910,N_11906);
nor U13211 (N_13211,N_11717,N_11873);
and U13212 (N_13212,N_11961,N_9951);
nand U13213 (N_13213,N_8362,N_9440);
nor U13214 (N_13214,N_11960,N_9496);
or U13215 (N_13215,N_11738,N_8162);
xor U13216 (N_13216,N_11059,N_11031);
nand U13217 (N_13217,N_9070,N_8135);
nand U13218 (N_13218,N_11777,N_8739);
or U13219 (N_13219,N_9237,N_10935);
and U13220 (N_13220,N_8758,N_10821);
xnor U13221 (N_13221,N_10125,N_8264);
and U13222 (N_13222,N_8479,N_8760);
nor U13223 (N_13223,N_9647,N_11289);
nor U13224 (N_13224,N_9847,N_8341);
nor U13225 (N_13225,N_9064,N_11411);
nand U13226 (N_13226,N_11189,N_11448);
nor U13227 (N_13227,N_8589,N_10803);
xor U13228 (N_13228,N_11950,N_9363);
xor U13229 (N_13229,N_9372,N_8133);
or U13230 (N_13230,N_11626,N_10996);
nor U13231 (N_13231,N_8981,N_9828);
xnor U13232 (N_13232,N_9256,N_8365);
nor U13233 (N_13233,N_8040,N_9155);
and U13234 (N_13234,N_9573,N_10141);
and U13235 (N_13235,N_11784,N_11175);
nand U13236 (N_13236,N_8898,N_9845);
and U13237 (N_13237,N_10958,N_11484);
and U13238 (N_13238,N_9795,N_9587);
or U13239 (N_13239,N_10391,N_10874);
nor U13240 (N_13240,N_11569,N_8347);
nand U13241 (N_13241,N_10182,N_10109);
nand U13242 (N_13242,N_9115,N_9904);
and U13243 (N_13243,N_8700,N_10264);
and U13244 (N_13244,N_8725,N_8727);
nor U13245 (N_13245,N_10734,N_11123);
xor U13246 (N_13246,N_8071,N_11232);
nor U13247 (N_13247,N_10630,N_10531);
xnor U13248 (N_13248,N_11697,N_10344);
nor U13249 (N_13249,N_11234,N_11467);
or U13250 (N_13250,N_8567,N_9872);
and U13251 (N_13251,N_10191,N_8919);
nor U13252 (N_13252,N_11601,N_8945);
nor U13253 (N_13253,N_9464,N_10539);
or U13254 (N_13254,N_11548,N_8103);
xor U13255 (N_13255,N_11611,N_10090);
nor U13256 (N_13256,N_9420,N_10757);
xnor U13257 (N_13257,N_11707,N_8248);
nand U13258 (N_13258,N_11042,N_10382);
nand U13259 (N_13259,N_9675,N_11025);
nor U13260 (N_13260,N_10405,N_11253);
and U13261 (N_13261,N_9780,N_8356);
xor U13262 (N_13262,N_10493,N_10546);
nand U13263 (N_13263,N_8858,N_9400);
nand U13264 (N_13264,N_8923,N_11994);
xnor U13265 (N_13265,N_9635,N_8721);
nor U13266 (N_13266,N_11180,N_11162);
nand U13267 (N_13267,N_8488,N_10969);
xnor U13268 (N_13268,N_11233,N_8473);
xnor U13269 (N_13269,N_9061,N_9415);
and U13270 (N_13270,N_11667,N_10274);
nor U13271 (N_13271,N_11679,N_9660);
or U13272 (N_13272,N_9659,N_8665);
or U13273 (N_13273,N_9405,N_11793);
nand U13274 (N_13274,N_8072,N_10129);
and U13275 (N_13275,N_9293,N_11276);
or U13276 (N_13276,N_9528,N_9863);
nand U13277 (N_13277,N_9258,N_8622);
nor U13278 (N_13278,N_9003,N_10744);
xor U13279 (N_13279,N_9982,N_11976);
xor U13280 (N_13280,N_9148,N_10674);
xnor U13281 (N_13281,N_9486,N_8096);
or U13282 (N_13282,N_8632,N_10847);
or U13283 (N_13283,N_8761,N_11778);
nor U13284 (N_13284,N_10309,N_9401);
and U13285 (N_13285,N_10322,N_8123);
xnor U13286 (N_13286,N_9973,N_10325);
nand U13287 (N_13287,N_8638,N_9485);
xnor U13288 (N_13288,N_9353,N_10896);
nor U13289 (N_13289,N_10255,N_8302);
nor U13290 (N_13290,N_11699,N_11079);
and U13291 (N_13291,N_10203,N_10622);
nand U13292 (N_13292,N_10668,N_8915);
xor U13293 (N_13293,N_9515,N_11928);
or U13294 (N_13294,N_10981,N_9429);
xnor U13295 (N_13295,N_10507,N_10764);
and U13296 (N_13296,N_11613,N_11285);
nor U13297 (N_13297,N_8459,N_9772);
and U13298 (N_13298,N_11091,N_8403);
nor U13299 (N_13299,N_11279,N_9213);
and U13300 (N_13300,N_10061,N_11488);
xnor U13301 (N_13301,N_10751,N_9591);
nor U13302 (N_13302,N_10796,N_8031);
or U13303 (N_13303,N_8714,N_9654);
or U13304 (N_13304,N_9581,N_11009);
nand U13305 (N_13305,N_8225,N_10266);
or U13306 (N_13306,N_8829,N_10963);
or U13307 (N_13307,N_8754,N_11493);
xnor U13308 (N_13308,N_10964,N_11562);
nand U13309 (N_13309,N_9850,N_9149);
nand U13310 (N_13310,N_10571,N_10054);
xnor U13311 (N_13311,N_10101,N_8198);
nand U13312 (N_13312,N_10210,N_8744);
and U13313 (N_13313,N_10169,N_10281);
xnor U13314 (N_13314,N_11063,N_11832);
nand U13315 (N_13315,N_11715,N_11013);
and U13316 (N_13316,N_10742,N_9037);
xnor U13317 (N_13317,N_9275,N_11049);
nand U13318 (N_13318,N_8229,N_10137);
nand U13319 (N_13319,N_8516,N_10731);
nand U13320 (N_13320,N_10988,N_9815);
xor U13321 (N_13321,N_8643,N_10807);
xnor U13322 (N_13322,N_10385,N_10557);
nor U13323 (N_13323,N_9231,N_9499);
nand U13324 (N_13324,N_10589,N_10434);
and U13325 (N_13325,N_9544,N_9560);
or U13326 (N_13326,N_8078,N_10548);
and U13327 (N_13327,N_11816,N_8068);
xnor U13328 (N_13328,N_9550,N_11078);
nand U13329 (N_13329,N_9187,N_8851);
nor U13330 (N_13330,N_11916,N_10666);
and U13331 (N_13331,N_8704,N_11710);
xor U13332 (N_13332,N_8375,N_10736);
xor U13333 (N_13333,N_11030,N_11935);
nor U13334 (N_13334,N_8093,N_9022);
nand U13335 (N_13335,N_11612,N_9057);
or U13336 (N_13336,N_9489,N_10289);
nand U13337 (N_13337,N_8674,N_11686);
or U13338 (N_13338,N_9616,N_11459);
and U13339 (N_13339,N_11424,N_9210);
and U13340 (N_13340,N_10482,N_9299);
nor U13341 (N_13341,N_8872,N_11660);
or U13342 (N_13342,N_11406,N_11076);
or U13343 (N_13343,N_10381,N_10220);
or U13344 (N_13344,N_9840,N_10321);
or U13345 (N_13345,N_10902,N_10451);
xnor U13346 (N_13346,N_11760,N_10906);
nand U13347 (N_13347,N_9714,N_10192);
or U13348 (N_13348,N_11990,N_10735);
and U13349 (N_13349,N_9876,N_11501);
or U13350 (N_13350,N_11705,N_11621);
nor U13351 (N_13351,N_10805,N_10883);
and U13352 (N_13352,N_10974,N_11228);
or U13353 (N_13353,N_9874,N_11922);
xnor U13354 (N_13354,N_11868,N_10411);
nor U13355 (N_13355,N_11096,N_8512);
or U13356 (N_13356,N_11709,N_10959);
nand U13357 (N_13357,N_9891,N_8952);
nor U13358 (N_13358,N_8102,N_11350);
nor U13359 (N_13359,N_8661,N_11957);
nand U13360 (N_13360,N_8550,N_8051);
xor U13361 (N_13361,N_9263,N_10424);
or U13362 (N_13362,N_11646,N_8422);
nor U13363 (N_13363,N_10794,N_11080);
or U13364 (N_13364,N_10866,N_8837);
and U13365 (N_13365,N_11243,N_11670);
nand U13366 (N_13366,N_8240,N_10891);
or U13367 (N_13367,N_10159,N_10074);
and U13368 (N_13368,N_10346,N_8084);
nor U13369 (N_13369,N_11880,N_9758);
xor U13370 (N_13370,N_8929,N_8894);
or U13371 (N_13371,N_11859,N_11454);
and U13372 (N_13372,N_10331,N_11671);
nand U13373 (N_13373,N_9319,N_9077);
and U13374 (N_13374,N_10138,N_8594);
nand U13375 (N_13375,N_11471,N_10558);
nand U13376 (N_13376,N_8366,N_10700);
nand U13377 (N_13377,N_10535,N_8712);
nand U13378 (N_13378,N_9769,N_8328);
or U13379 (N_13379,N_9932,N_9101);
and U13380 (N_13380,N_10663,N_8715);
nand U13381 (N_13381,N_10968,N_11407);
xnor U13382 (N_13382,N_8013,N_11056);
nor U13383 (N_13383,N_8200,N_9911);
nand U13384 (N_13384,N_11691,N_8853);
and U13385 (N_13385,N_11719,N_11897);
xor U13386 (N_13386,N_11819,N_9423);
nor U13387 (N_13387,N_10514,N_11700);
nand U13388 (N_13388,N_10403,N_10941);
nor U13389 (N_13389,N_10646,N_8669);
and U13390 (N_13390,N_8728,N_8191);
nand U13391 (N_13391,N_11421,N_8933);
nand U13392 (N_13392,N_10694,N_8147);
xor U13393 (N_13393,N_9785,N_10565);
xor U13394 (N_13394,N_8489,N_8309);
xnor U13395 (N_13395,N_8398,N_11598);
nor U13396 (N_13396,N_8989,N_10215);
nand U13397 (N_13397,N_8032,N_11838);
nand U13398 (N_13398,N_11254,N_10115);
nand U13399 (N_13399,N_8164,N_11729);
nor U13400 (N_13400,N_11883,N_10437);
nor U13401 (N_13401,N_8694,N_8767);
nand U13402 (N_13402,N_9477,N_9702);
and U13403 (N_13403,N_10602,N_8446);
and U13404 (N_13404,N_10076,N_11516);
and U13405 (N_13405,N_10808,N_8321);
nor U13406 (N_13406,N_8535,N_11485);
nand U13407 (N_13407,N_11891,N_11281);
and U13408 (N_13408,N_10252,N_11638);
or U13409 (N_13409,N_11469,N_8082);
nand U13410 (N_13410,N_9596,N_8786);
nor U13411 (N_13411,N_8792,N_11451);
nand U13412 (N_13412,N_10318,N_11876);
nor U13413 (N_13413,N_9347,N_8338);
or U13414 (N_13414,N_9394,N_9281);
and U13415 (N_13415,N_10131,N_8399);
nor U13416 (N_13416,N_11958,N_8642);
and U13417 (N_13417,N_11881,N_9397);
nor U13418 (N_13418,N_11135,N_8369);
nor U13419 (N_13419,N_9778,N_9783);
or U13420 (N_13420,N_8055,N_11480);
nand U13421 (N_13421,N_8825,N_9976);
nand U13422 (N_13422,N_11866,N_8029);
nand U13423 (N_13423,N_10965,N_8591);
and U13424 (N_13424,N_11483,N_8405);
nor U13425 (N_13425,N_10414,N_10718);
and U13426 (N_13426,N_8232,N_10885);
nor U13427 (N_13427,N_9129,N_8453);
nand U13428 (N_13428,N_9642,N_8202);
nor U13429 (N_13429,N_9355,N_9219);
xnor U13430 (N_13430,N_9841,N_10673);
nand U13431 (N_13431,N_9480,N_8493);
or U13432 (N_13432,N_8789,N_8349);
nor U13433 (N_13433,N_9653,N_11886);
and U13434 (N_13434,N_11641,N_9238);
xnor U13435 (N_13435,N_8816,N_9233);
or U13436 (N_13436,N_10495,N_9277);
or U13437 (N_13437,N_10134,N_8607);
nand U13438 (N_13438,N_10290,N_10135);
nand U13439 (N_13439,N_10709,N_8283);
nand U13440 (N_13440,N_10922,N_11153);
nand U13441 (N_13441,N_9946,N_11292);
or U13442 (N_13442,N_8874,N_11064);
nor U13443 (N_13443,N_9681,N_11069);
and U13444 (N_13444,N_9718,N_11579);
and U13445 (N_13445,N_11812,N_10617);
or U13446 (N_13446,N_9053,N_11318);
or U13447 (N_13447,N_8805,N_9802);
nand U13448 (N_13448,N_9243,N_8937);
xnor U13449 (N_13449,N_9523,N_8521);
or U13450 (N_13450,N_9934,N_11500);
xnor U13451 (N_13451,N_10581,N_10226);
and U13452 (N_13452,N_8185,N_8941);
nand U13453 (N_13453,N_10293,N_9507);
xor U13454 (N_13454,N_10781,N_10826);
nor U13455 (N_13455,N_8980,N_8224);
xor U13456 (N_13456,N_9114,N_8433);
and U13457 (N_13457,N_8682,N_11248);
xor U13458 (N_13458,N_11666,N_8831);
or U13459 (N_13459,N_9559,N_8738);
xor U13460 (N_13460,N_8419,N_9139);
xor U13461 (N_13461,N_8097,N_11294);
and U13462 (N_13462,N_10778,N_8844);
nor U13463 (N_13463,N_11887,N_9773);
or U13464 (N_13464,N_11311,N_10190);
and U13465 (N_13465,N_10221,N_9949);
or U13466 (N_13466,N_9131,N_11973);
xor U13467 (N_13467,N_10905,N_11759);
and U13468 (N_13468,N_10219,N_8352);
nand U13469 (N_13469,N_9492,N_9938);
xor U13470 (N_13470,N_11000,N_10943);
nor U13471 (N_13471,N_8063,N_10628);
xor U13472 (N_13472,N_8287,N_8506);
or U13473 (N_13473,N_10326,N_8938);
nor U13474 (N_13474,N_11346,N_10384);
and U13475 (N_13475,N_8016,N_8581);
nor U13476 (N_13476,N_11127,N_11071);
nand U13477 (N_13477,N_9980,N_9577);
xor U13478 (N_13478,N_9427,N_11842);
nand U13479 (N_13479,N_9684,N_11712);
or U13480 (N_13480,N_9894,N_8058);
or U13481 (N_13481,N_10595,N_9455);
nand U13482 (N_13482,N_10812,N_10513);
nor U13483 (N_13483,N_8620,N_9452);
nor U13484 (N_13484,N_11650,N_11681);
nor U13485 (N_13485,N_11841,N_10310);
nand U13486 (N_13486,N_11470,N_9728);
xor U13487 (N_13487,N_9603,N_11206);
nand U13488 (N_13488,N_8443,N_11944);
or U13489 (N_13489,N_8498,N_9153);
nor U13490 (N_13490,N_9035,N_10366);
xnor U13491 (N_13491,N_9983,N_9524);
or U13492 (N_13492,N_8928,N_8119);
and U13493 (N_13493,N_10977,N_9130);
or U13494 (N_13494,N_11369,N_11507);
xor U13495 (N_13495,N_8962,N_9700);
xnor U13496 (N_13496,N_9459,N_11242);
xor U13497 (N_13497,N_11273,N_8002);
xor U13498 (N_13498,N_11200,N_10516);
and U13499 (N_13499,N_8533,N_9827);
or U13500 (N_13500,N_10740,N_11727);
xor U13501 (N_13501,N_11304,N_10835);
nor U13502 (N_13502,N_9689,N_9051);
xor U13503 (N_13503,N_9615,N_10639);
nor U13504 (N_13504,N_9280,N_8778);
or U13505 (N_13505,N_10560,N_9031);
and U13506 (N_13506,N_8854,N_9589);
or U13507 (N_13507,N_10302,N_11509);
nor U13508 (N_13508,N_8599,N_10395);
xnor U13509 (N_13509,N_9954,N_11889);
and U13510 (N_13510,N_9138,N_11745);
or U13511 (N_13511,N_10933,N_9739);
nor U13512 (N_13512,N_11167,N_8317);
and U13513 (N_13513,N_10117,N_11645);
or U13514 (N_13514,N_10653,N_10893);
and U13515 (N_13515,N_8819,N_10909);
and U13516 (N_13516,N_9760,N_8150);
nor U13517 (N_13517,N_10167,N_9287);
and U13518 (N_13518,N_8799,N_8888);
and U13519 (N_13519,N_10979,N_11904);
nor U13520 (N_13520,N_10624,N_10444);
xnor U13521 (N_13521,N_11052,N_11414);
nor U13522 (N_13522,N_10392,N_9956);
nor U13523 (N_13523,N_11177,N_9136);
nor U13524 (N_13524,N_9412,N_11028);
nor U13525 (N_13525,N_8706,N_11643);
nor U13526 (N_13526,N_9468,N_8186);
nor U13527 (N_13527,N_8057,N_8081);
nand U13528 (N_13528,N_11773,N_9940);
nor U13529 (N_13529,N_8210,N_10611);
or U13530 (N_13530,N_9297,N_8373);
xnor U13531 (N_13531,N_10490,N_9376);
or U13532 (N_13532,N_8828,N_9119);
xor U13533 (N_13533,N_11129,N_8122);
nand U13534 (N_13534,N_11905,N_8974);
nand U13535 (N_13535,N_9446,N_9563);
and U13536 (N_13536,N_8855,N_9411);
nand U13537 (N_13537,N_9746,N_8172);
nand U13538 (N_13538,N_11688,N_10561);
and U13539 (N_13539,N_9066,N_10452);
and U13540 (N_13540,N_11566,N_8371);
or U13541 (N_13541,N_8703,N_9121);
xor U13542 (N_13542,N_11288,N_10586);
nand U13543 (N_13543,N_9525,N_8610);
xor U13544 (N_13544,N_8889,N_8526);
nor U13545 (N_13545,N_10978,N_8982);
or U13546 (N_13546,N_11525,N_9126);
or U13547 (N_13547,N_9067,N_11298);
nand U13548 (N_13548,N_10786,N_8582);
xor U13549 (N_13549,N_9135,N_8330);
or U13550 (N_13550,N_10590,N_11967);
xor U13551 (N_13551,N_11203,N_9014);
nand U13552 (N_13552,N_10733,N_9511);
or U13553 (N_13553,N_9555,N_11722);
xnor U13554 (N_13554,N_11295,N_11221);
and U13555 (N_13555,N_8115,N_10332);
xor U13556 (N_13556,N_9042,N_11440);
nand U13557 (N_13557,N_10196,N_9006);
nand U13558 (N_13558,N_8670,N_11053);
nand U13559 (N_13559,N_11684,N_9884);
or U13560 (N_13560,N_11152,N_9431);
and U13561 (N_13561,N_10899,N_10383);
and U13562 (N_13562,N_9050,N_9918);
xnor U13563 (N_13563,N_11752,N_11564);
and U13564 (N_13564,N_11438,N_8148);
or U13565 (N_13565,N_8667,N_9925);
or U13566 (N_13566,N_8986,N_8502);
xnor U13567 (N_13567,N_8324,N_9625);
and U13568 (N_13568,N_10767,N_8867);
nand U13569 (N_13569,N_11340,N_11573);
xor U13570 (N_13570,N_9335,N_11227);
or U13571 (N_13571,N_11590,N_9862);
nand U13572 (N_13572,N_9944,N_9313);
nor U13573 (N_13573,N_11655,N_9044);
xnor U13574 (N_13574,N_9624,N_10777);
nor U13575 (N_13575,N_9987,N_10645);
or U13576 (N_13576,N_10489,N_9063);
nor U13577 (N_13577,N_10566,N_8333);
and U13578 (N_13578,N_9472,N_9825);
and U13579 (N_13579,N_11284,N_8066);
nand U13580 (N_13580,N_8483,N_10039);
nand U13581 (N_13581,N_10676,N_8464);
and U13582 (N_13582,N_9919,N_11087);
and U13583 (N_13583,N_11282,N_11149);
and U13584 (N_13584,N_10371,N_10245);
and U13585 (N_13585,N_8768,N_10417);
xor U13586 (N_13586,N_10474,N_10471);
xor U13587 (N_13587,N_9823,N_10871);
nand U13588 (N_13588,N_11075,N_8902);
and U13589 (N_13589,N_9043,N_9073);
nor U13590 (N_13590,N_11160,N_9089);
and U13591 (N_13591,N_9831,N_10323);
nor U13592 (N_13592,N_8101,N_10657);
and U13593 (N_13593,N_8565,N_10256);
and U13594 (N_13594,N_9527,N_8099);
nor U13595 (N_13595,N_11387,N_10122);
nand U13596 (N_13596,N_8577,N_8314);
and U13597 (N_13597,N_10877,N_9953);
nor U13598 (N_13598,N_8110,N_11449);
xor U13599 (N_13599,N_11947,N_8425);
xor U13600 (N_13600,N_10110,N_11473);
nand U13601 (N_13601,N_9018,N_10170);
nor U13602 (N_13602,N_9639,N_11465);
xnor U13603 (N_13603,N_8271,N_11528);
nor U13604 (N_13604,N_9254,N_8161);
and U13605 (N_13605,N_8561,N_9267);
nor U13606 (N_13606,N_8378,N_10472);
and U13607 (N_13607,N_10648,N_10091);
xor U13608 (N_13608,N_11698,N_9183);
and U13609 (N_13609,N_9406,N_11268);
and U13610 (N_13610,N_11966,N_10994);
or U13611 (N_13611,N_11863,N_8608);
and U13612 (N_13612,N_8730,N_8794);
nor U13613 (N_13613,N_9534,N_11142);
or U13614 (N_13614,N_10194,N_10353);
and U13615 (N_13615,N_10412,N_9671);
nand U13616 (N_13616,N_9315,N_10180);
xnor U13617 (N_13617,N_8308,N_10211);
or U13618 (N_13618,N_11181,N_11489);
nor U13619 (N_13619,N_9345,N_9572);
xnor U13620 (N_13620,N_9334,N_8950);
nor U13621 (N_13621,N_9584,N_8449);
and U13622 (N_13622,N_10372,N_11736);
nor U13623 (N_13623,N_9545,N_9151);
nor U13624 (N_13624,N_8559,N_10687);
or U13625 (N_13625,N_9701,N_11430);
and U13626 (N_13626,N_10494,N_9300);
and U13627 (N_13627,N_8838,N_10021);
and U13628 (N_13628,N_8404,N_9962);
or U13629 (N_13629,N_11702,N_10239);
nor U13630 (N_13630,N_11088,N_9928);
nor U13631 (N_13631,N_8005,N_11353);
or U13632 (N_13632,N_10591,N_8329);
nand U13633 (N_13633,N_11313,N_8204);
xnor U13634 (N_13634,N_9169,N_9709);
nand U13635 (N_13635,N_9145,N_11371);
nand U13636 (N_13636,N_11435,N_11653);
nand U13637 (N_13637,N_8916,N_9537);
or U13638 (N_13638,N_11443,N_10995);
and U13639 (N_13639,N_10538,N_11373);
or U13640 (N_13640,N_9048,N_8196);
nor U13641 (N_13641,N_10019,N_9125);
nand U13642 (N_13642,N_9144,N_9134);
nor U13643 (N_13643,N_11925,N_8718);
xor U13644 (N_13644,N_8556,N_9170);
xor U13645 (N_13645,N_9685,N_9369);
and U13646 (N_13646,N_9038,N_11272);
nand U13647 (N_13647,N_9046,N_8520);
nand U13648 (N_13648,N_11257,N_10027);
nor U13649 (N_13649,N_9665,N_11183);
xnor U13650 (N_13650,N_11565,N_8796);
or U13651 (N_13651,N_8895,N_8508);
and U13652 (N_13652,N_9875,N_10130);
xor U13653 (N_13653,N_11427,N_10542);
xor U13654 (N_13654,N_10529,N_10008);
and U13655 (N_13655,N_10824,N_9920);
nor U13656 (N_13656,N_10547,N_11926);
nand U13657 (N_13657,N_10615,N_8752);
xnor U13658 (N_13658,N_8537,N_8268);
and U13659 (N_13659,N_9707,N_9806);
or U13660 (N_13660,N_11492,N_11068);
nor U13661 (N_13661,N_10875,N_10055);
nor U13662 (N_13662,N_8091,N_9794);
nor U13663 (N_13663,N_9230,N_9985);
nand U13664 (N_13664,N_8939,N_11136);
xor U13665 (N_13665,N_9513,N_8100);
nand U13666 (N_13666,N_10168,N_8551);
xor U13667 (N_13667,N_9814,N_8908);
nand U13668 (N_13668,N_10356,N_11374);
or U13669 (N_13669,N_8993,N_8252);
nor U13670 (N_13670,N_10479,N_11439);
nand U13671 (N_13671,N_8790,N_10570);
xnor U13672 (N_13672,N_8279,N_9968);
or U13673 (N_13673,N_11212,N_10084);
xor U13674 (N_13674,N_10431,N_9087);
nand U13675 (N_13675,N_9364,N_10704);
and U13676 (N_13676,N_8038,N_11479);
and U13677 (N_13677,N_8497,N_11426);
xor U13678 (N_13678,N_9010,N_10419);
and U13679 (N_13679,N_8197,N_11084);
nand U13680 (N_13680,N_8782,N_10329);
nor U13681 (N_13681,N_10746,N_8295);
and U13682 (N_13682,N_10271,N_10447);
and U13683 (N_13683,N_10397,N_9506);
and U13684 (N_13684,N_8500,N_11846);
and U13685 (N_13685,N_8408,N_10396);
nor U13686 (N_13686,N_9623,N_9939);
nor U13687 (N_13687,N_10314,N_8251);
nor U13688 (N_13688,N_10518,N_11399);
nor U13689 (N_13689,N_9221,N_10093);
nor U13690 (N_13690,N_8992,N_11875);
and U13691 (N_13691,N_10037,N_8118);
nor U13692 (N_13692,N_10556,N_8227);
and U13693 (N_13693,N_8238,N_11131);
xor U13694 (N_13694,N_11837,N_8955);
xor U13695 (N_13695,N_11577,N_9030);
or U13696 (N_13696,N_11309,N_9974);
or U13697 (N_13697,N_8870,N_9817);
xnor U13698 (N_13698,N_9931,N_8429);
nor U13699 (N_13699,N_10014,N_9776);
nand U13700 (N_13700,N_9909,N_11463);
nor U13701 (N_13701,N_8757,N_8409);
and U13702 (N_13702,N_8875,N_11003);
nand U13703 (N_13703,N_10761,N_10324);
nor U13704 (N_13704,N_10898,N_8652);
or U13705 (N_13705,N_9292,N_11151);
or U13706 (N_13706,N_9056,N_10572);
or U13707 (N_13707,N_11121,N_11477);
xnor U13708 (N_13708,N_10517,N_11694);
xnor U13709 (N_13709,N_9298,N_8879);
nor U13710 (N_13710,N_10373,N_10577);
nor U13711 (N_13711,N_9320,N_11820);
nor U13712 (N_13712,N_9285,N_11168);
xnor U13713 (N_13713,N_8654,N_11466);
nand U13714 (N_13714,N_8104,N_8840);
and U13715 (N_13715,N_11965,N_8105);
xnor U13716 (N_13716,N_10864,N_10283);
nor U13717 (N_13717,N_8192,N_8180);
or U13718 (N_13718,N_9160,N_8174);
nand U13719 (N_13719,N_9008,N_10058);
nor U13720 (N_13720,N_11378,N_9526);
nor U13721 (N_13721,N_11929,N_10748);
xor U13722 (N_13722,N_9999,N_10421);
nand U13723 (N_13723,N_11902,N_9367);
xor U13724 (N_13724,N_8777,N_9332);
nor U13725 (N_13725,N_9906,N_8322);
nand U13726 (N_13726,N_11938,N_11541);
nand U13727 (N_13727,N_10788,N_9168);
nor U13728 (N_13728,N_11204,N_10175);
or U13729 (N_13729,N_9819,N_9015);
and U13730 (N_13730,N_9917,N_10156);
xnor U13731 (N_13731,N_9651,N_10010);
nand U13732 (N_13732,N_10923,N_10305);
or U13733 (N_13733,N_11517,N_8807);
and U13734 (N_13734,N_11815,N_10991);
nand U13735 (N_13735,N_11453,N_9189);
or U13736 (N_13736,N_8217,N_9228);
nand U13737 (N_13737,N_11225,N_9442);
and U13738 (N_13738,N_10976,N_9725);
and U13739 (N_13739,N_9747,N_10303);
xnor U13740 (N_13740,N_11743,N_9331);
or U13741 (N_13741,N_8749,N_10188);
xnor U13742 (N_13742,N_9585,N_11898);
and U13743 (N_13743,N_9498,N_8423);
or U13744 (N_13744,N_10118,N_8337);
xor U13745 (N_13745,N_11766,N_8735);
xor U13746 (N_13746,N_9133,N_11141);
or U13747 (N_13747,N_9069,N_10837);
nor U13748 (N_13748,N_10232,N_9323);
or U13749 (N_13749,N_10399,N_8090);
xnor U13750 (N_13750,N_8733,N_10827);
or U13751 (N_13751,N_9678,N_11952);
nor U13752 (N_13752,N_10012,N_9432);
or U13753 (N_13753,N_9570,N_9356);
nand U13754 (N_13754,N_8216,N_9002);
nor U13755 (N_13755,N_9099,N_9438);
nor U13756 (N_13756,N_9197,N_11751);
xnor U13757 (N_13757,N_11441,N_11805);
nor U13758 (N_13758,N_10176,N_8740);
and U13759 (N_13759,N_11622,N_9892);
or U13760 (N_13760,N_10881,N_9830);
or U13761 (N_13761,N_11620,N_10446);
nor U13762 (N_13762,N_11001,N_10341);
nor U13763 (N_13763,N_10634,N_11455);
nor U13764 (N_13764,N_10997,N_9249);
and U13765 (N_13765,N_11039,N_10133);
and U13766 (N_13766,N_11913,N_8552);
and U13767 (N_13767,N_9017,N_11673);
xnor U13768 (N_13768,N_10533,N_8684);
xor U13769 (N_13769,N_8233,N_8427);
or U13770 (N_13770,N_9979,N_10069);
nand U13771 (N_13771,N_8145,N_11337);
and U13772 (N_13772,N_9816,N_9740);
xor U13773 (N_13773,N_11472,N_9879);
or U13774 (N_13774,N_11278,N_9729);
xor U13775 (N_13775,N_8382,N_11335);
or U13776 (N_13776,N_10151,N_11713);
xnor U13777 (N_13777,N_11605,N_11914);
nand U13778 (N_13778,N_10477,N_8839);
and U13779 (N_13779,N_9766,N_10243);
and U13780 (N_13780,N_9888,N_10549);
nor U13781 (N_13781,N_10204,N_11363);
or U13782 (N_13782,N_9348,N_8269);
and U13783 (N_13783,N_10588,N_8477);
nor U13784 (N_13784,N_10505,N_8230);
xnor U13785 (N_13785,N_8126,N_11739);
nor U13786 (N_13786,N_9274,N_10045);
or U13787 (N_13787,N_9864,N_11865);
or U13788 (N_13788,N_9185,N_8447);
nand U13789 (N_13789,N_10496,N_10886);
nand U13790 (N_13790,N_8696,N_8026);
xor U13791 (N_13791,N_8407,N_11979);
nand U13792 (N_13792,N_9242,N_9352);
nor U13793 (N_13793,N_11377,N_10453);
nor U13794 (N_13794,N_10618,N_9634);
and U13795 (N_13795,N_11585,N_11351);
nand U13796 (N_13796,N_9521,N_10598);
xnor U13797 (N_13797,N_8183,N_10456);
nor U13798 (N_13798,N_10822,N_9607);
nor U13799 (N_13799,N_10573,N_9290);
or U13800 (N_13800,N_8440,N_11607);
nand U13801 (N_13801,N_8465,N_11998);
nor U13802 (N_13802,N_11578,N_9765);
xnor U13803 (N_13803,N_11372,N_9571);
nand U13804 (N_13804,N_8572,N_11513);
and U13805 (N_13805,N_10937,N_9192);
nor U13806 (N_13806,N_8208,N_9328);
nor U13807 (N_13807,N_9444,N_10124);
xnor U13808 (N_13808,N_10903,N_8401);
and U13809 (N_13809,N_9404,N_8462);
nand U13810 (N_13810,N_10205,N_9303);
or U13811 (N_13811,N_11081,N_10982);
or U13812 (N_13812,N_11437,N_8791);
nand U13813 (N_13813,N_8514,N_10094);
and U13814 (N_13814,N_10048,N_8959);
xor U13815 (N_13815,N_8088,N_9722);
nor U13816 (N_13816,N_8157,N_8518);
xnor U13817 (N_13817,N_11589,N_8576);
xor U13818 (N_13818,N_11560,N_8539);
and U13819 (N_13819,N_11514,N_10760);
nor U13820 (N_13820,N_9745,N_10429);
xor U13821 (N_13821,N_11871,N_9324);
nand U13822 (N_13822,N_8209,N_10017);
nor U13823 (N_13823,N_10998,N_9704);
xor U13824 (N_13824,N_11789,N_11481);
nand U13825 (N_13825,N_8627,N_8397);
or U13826 (N_13826,N_9310,N_8304);
nand U13827 (N_13827,N_11969,N_9165);
and U13828 (N_13828,N_8175,N_11434);
or U13829 (N_13829,N_9322,N_8236);
xnor U13830 (N_13830,N_10695,N_10942);
nor U13831 (N_13831,N_11464,N_8151);
or U13832 (N_13832,N_9959,N_11376);
xor U13833 (N_13833,N_9301,N_10867);
nor U13834 (N_13834,N_8455,N_8769);
nor U13835 (N_13835,N_8869,N_11388);
or U13836 (N_13836,N_10306,N_11021);
xor U13837 (N_13837,N_10621,N_11708);
or U13838 (N_13838,N_10656,N_10779);
xnor U13839 (N_13839,N_8486,N_9690);
or U13840 (N_13840,N_8762,N_11051);
and U13841 (N_13841,N_11665,N_9137);
nand U13842 (N_13842,N_8904,N_9580);
nor U13843 (N_13843,N_9284,N_10195);
xnor U13844 (N_13844,N_9314,N_11139);
nor U13845 (N_13845,N_11041,N_11530);
xor U13846 (N_13846,N_9926,N_11746);
and U13847 (N_13847,N_11861,N_11828);
or U13848 (N_13848,N_11016,N_10068);
xnor U13849 (N_13849,N_10486,N_11089);
xor U13850 (N_13850,N_8015,N_8523);
or U13851 (N_13851,N_8863,N_10574);
nand U13852 (N_13852,N_8555,N_11804);
nand U13853 (N_13853,N_8826,N_10859);
nor U13854 (N_13854,N_10851,N_10932);
nor U13855 (N_13855,N_11677,N_9062);
and U13856 (N_13856,N_10732,N_10608);
nand U13857 (N_13857,N_11682,N_9437);
xnor U13858 (N_13858,N_11107,N_9448);
or U13859 (N_13859,N_9020,N_10749);
xor U13860 (N_13860,N_8973,N_9905);
nor U13861 (N_13861,N_10075,N_10596);
and U13862 (N_13862,N_9007,N_8132);
nor U13863 (N_13863,N_10790,N_10269);
nor U13864 (N_13864,N_8751,N_10759);
and U13865 (N_13865,N_10945,N_11632);
xor U13866 (N_13866,N_10829,N_10183);
nor U13867 (N_13867,N_11341,N_8416);
nand U13868 (N_13868,N_9798,N_8085);
nand U13869 (N_13869,N_10983,N_10705);
nand U13870 (N_13870,N_10153,N_11219);
xnor U13871 (N_13871,N_9820,N_8947);
nand U13872 (N_13872,N_9199,N_8176);
or U13873 (N_13873,N_11687,N_11942);
or U13874 (N_13874,N_11749,N_11809);
nor U13875 (N_13875,N_11827,N_10198);
xor U13876 (N_13876,N_9818,N_10340);
or U13877 (N_13877,N_11306,N_10098);
and U13878 (N_13878,N_9836,N_10380);
nand U13879 (N_13879,N_8664,N_8061);
nand U13880 (N_13880,N_10895,N_11147);
nor U13881 (N_13881,N_11375,N_11312);
and U13882 (N_13882,N_10261,N_8554);
or U13883 (N_13883,N_9540,N_11892);
or U13884 (N_13884,N_11099,N_8472);
nand U13885 (N_13885,N_8930,N_11584);
nand U13886 (N_13886,N_8604,N_11368);
nor U13887 (N_13887,N_8920,N_8311);
or U13888 (N_13888,N_10888,N_11955);
nand U13889 (N_13889,N_9478,N_10716);
nor U13890 (N_13890,N_8880,N_10241);
nor U13891 (N_13891,N_11767,N_11004);
nand U13892 (N_13892,N_9640,N_9466);
and U13893 (N_13893,N_8463,N_9881);
or U13894 (N_13894,N_11014,N_8549);
nor U13895 (N_13895,N_10487,N_10681);
or U13896 (N_13896,N_11291,N_10865);
nand U13897 (N_13897,N_10003,N_10394);
or U13898 (N_13898,N_10636,N_8968);
and U13899 (N_13899,N_10838,N_8114);
nand U13900 (N_13900,N_11790,N_11862);
nand U13901 (N_13901,N_10567,N_10640);
nand U13902 (N_13902,N_8491,N_10032);
or U13903 (N_13903,N_11137,N_10619);
nand U13904 (N_13904,N_9011,N_11249);
nand U13905 (N_13905,N_11280,N_9713);
xnor U13906 (N_13906,N_11974,N_8530);
and U13907 (N_13907,N_11216,N_11101);
xnor U13908 (N_13908,N_10315,N_9590);
nor U13909 (N_13909,N_10370,N_11540);
xnor U13910 (N_13910,N_10121,N_11836);
or U13911 (N_13911,N_11110,N_8834);
nor U13912 (N_13912,N_11654,N_10753);
or U13913 (N_13913,N_11169,N_10745);
and U13914 (N_13914,N_9887,N_10576);
nor U13915 (N_13915,N_10755,N_8243);
nand U13916 (N_13916,N_11518,N_11120);
xnor U13917 (N_13917,N_8983,N_11884);
xor U13918 (N_13918,N_8042,N_8672);
nor U13919 (N_13919,N_8966,N_9821);
nor U13920 (N_13920,N_8310,N_8098);
nand U13921 (N_13921,N_11624,N_9851);
xnor U13922 (N_13922,N_8345,N_9941);
nand U13923 (N_13923,N_11293,N_8111);
xor U13924 (N_13924,N_8571,N_9208);
or U13925 (N_13925,N_10199,N_9990);
or U13926 (N_13926,N_10388,N_10698);
xor U13927 (N_13927,N_10171,N_9970);
nand U13928 (N_13928,N_8471,N_10279);
nand U13929 (N_13929,N_9768,N_10316);
nor U13930 (N_13930,N_9914,N_11822);
nand U13931 (N_13931,N_9861,N_10492);
nor U13932 (N_13932,N_9566,N_9935);
nor U13933 (N_13933,N_8540,N_11703);
xnor U13934 (N_13934,N_8527,N_11981);
nand U13935 (N_13935,N_9113,N_9408);
nand U13936 (N_13936,N_10339,N_9416);
and U13937 (N_13937,N_11982,N_8748);
or U13938 (N_13938,N_8043,N_10089);
and U13939 (N_13939,N_9548,N_11356);
nor U13940 (N_13940,N_9674,N_9627);
and U13941 (N_13941,N_11563,N_8734);
xor U13942 (N_13942,N_8882,N_11781);
nor U13943 (N_13943,N_9837,N_9190);
or U13944 (N_13944,N_10015,N_8011);
or U13945 (N_13945,N_11869,N_9049);
nor U13946 (N_13946,N_9143,N_8987);
xor U13947 (N_13947,N_10679,N_9901);
nand U13948 (N_13948,N_8406,N_10034);
nand U13949 (N_13949,N_8263,N_11635);
nand U13950 (N_13950,N_9606,N_10062);
and U13951 (N_13951,N_8944,N_10792);
xor U13952 (N_13952,N_10096,N_8359);
nor U13953 (N_13953,N_10398,N_11321);
and U13954 (N_13954,N_10473,N_8731);
nand U13955 (N_13955,N_8246,N_10702);
nand U13956 (N_13956,N_10259,N_10504);
nand U13957 (N_13957,N_9588,N_11652);
nand U13958 (N_13958,N_8231,N_8999);
nand U13959 (N_13959,N_10811,N_10868);
xnor U13960 (N_13960,N_11582,N_10214);
nor U13961 (N_13961,N_8495,N_8468);
and U13962 (N_13962,N_10832,N_8226);
nor U13963 (N_13963,N_9036,N_11867);
nand U13964 (N_13964,N_9108,N_9774);
or U13965 (N_13965,N_10809,N_8402);
nor U13966 (N_13966,N_9235,N_10481);
xnor U13967 (N_13967,N_9631,N_9602);
xnor U13968 (N_13968,N_10401,N_8951);
nor U13969 (N_13969,N_11823,N_10265);
nand U13970 (N_13970,N_8018,N_10237);
xnor U13971 (N_13971,N_11161,N_9476);
nand U13972 (N_13972,N_9306,N_11235);
xor U13973 (N_13973,N_11774,N_11054);
nor U13974 (N_13974,N_8395,N_8873);
nor U13975 (N_13975,N_10277,N_8806);
xnor U13976 (N_13976,N_8065,N_11197);
and U13977 (N_13977,N_11771,N_10257);
and U13978 (N_13978,N_8334,N_8573);
nand U13979 (N_13979,N_10162,N_10752);
xnor U13980 (N_13980,N_9522,N_8505);
nor U13981 (N_13981,N_11526,N_10508);
nand U13982 (N_13982,N_10703,N_8342);
and U13983 (N_13983,N_11503,N_10236);
nor U13984 (N_13984,N_10458,N_10328);
nor U13985 (N_13985,N_11245,N_10730);
nor U13986 (N_13986,N_10359,N_11496);
and U13987 (N_13987,N_11630,N_8411);
or U13988 (N_13988,N_9425,N_8946);
and U13989 (N_13989,N_10599,N_10515);
nand U13990 (N_13990,N_10523,N_11591);
nor U13991 (N_13991,N_11122,N_10699);
or U13992 (N_13992,N_10413,N_10854);
xor U13993 (N_13993,N_9569,N_11798);
xor U13994 (N_13994,N_10584,N_11352);
or U13995 (N_13995,N_9172,N_10418);
and U13996 (N_13996,N_11323,N_10320);
nor U13997 (N_13997,N_10880,N_9868);
and U13998 (N_13998,N_9389,N_8810);
or U13999 (N_13999,N_8815,N_8891);
and U14000 (N_14000,N_8081,N_9659);
nand U14001 (N_14001,N_8905,N_9932);
and U14002 (N_14002,N_10984,N_11001);
or U14003 (N_14003,N_10139,N_8796);
or U14004 (N_14004,N_9953,N_11582);
xor U14005 (N_14005,N_10499,N_9738);
xor U14006 (N_14006,N_8227,N_9123);
and U14007 (N_14007,N_8603,N_10580);
nor U14008 (N_14008,N_10622,N_11921);
and U14009 (N_14009,N_8122,N_11886);
nand U14010 (N_14010,N_8594,N_11499);
nor U14011 (N_14011,N_8923,N_11379);
and U14012 (N_14012,N_10009,N_9014);
nor U14013 (N_14013,N_10255,N_9124);
xnor U14014 (N_14014,N_8306,N_10217);
xor U14015 (N_14015,N_11647,N_9871);
nor U14016 (N_14016,N_8466,N_9682);
or U14017 (N_14017,N_11864,N_8837);
or U14018 (N_14018,N_10590,N_9261);
nand U14019 (N_14019,N_9612,N_10629);
and U14020 (N_14020,N_10766,N_10476);
and U14021 (N_14021,N_10493,N_8661);
nand U14022 (N_14022,N_10758,N_11682);
or U14023 (N_14023,N_9431,N_8008);
xnor U14024 (N_14024,N_11272,N_10991);
and U14025 (N_14025,N_9129,N_10916);
and U14026 (N_14026,N_10139,N_8605);
xnor U14027 (N_14027,N_10071,N_8957);
xnor U14028 (N_14028,N_9516,N_10116);
nor U14029 (N_14029,N_9697,N_9197);
nor U14030 (N_14030,N_8639,N_11397);
nor U14031 (N_14031,N_10719,N_10819);
or U14032 (N_14032,N_9955,N_8093);
nor U14033 (N_14033,N_11236,N_9756);
nor U14034 (N_14034,N_8523,N_10521);
and U14035 (N_14035,N_11005,N_8498);
and U14036 (N_14036,N_8937,N_10063);
xor U14037 (N_14037,N_9014,N_9473);
nor U14038 (N_14038,N_9356,N_10772);
xor U14039 (N_14039,N_9720,N_10317);
and U14040 (N_14040,N_8251,N_10485);
xnor U14041 (N_14041,N_8810,N_10320);
nand U14042 (N_14042,N_10461,N_9349);
nand U14043 (N_14043,N_8120,N_9038);
and U14044 (N_14044,N_11580,N_11308);
nand U14045 (N_14045,N_9752,N_10181);
or U14046 (N_14046,N_10749,N_11607);
or U14047 (N_14047,N_10874,N_11876);
nand U14048 (N_14048,N_9883,N_8945);
or U14049 (N_14049,N_9386,N_8581);
and U14050 (N_14050,N_9611,N_11863);
xnor U14051 (N_14051,N_10916,N_11479);
nand U14052 (N_14052,N_11686,N_8950);
or U14053 (N_14053,N_8492,N_9197);
and U14054 (N_14054,N_9984,N_11740);
nand U14055 (N_14055,N_11965,N_10174);
xnor U14056 (N_14056,N_8943,N_8611);
and U14057 (N_14057,N_9815,N_11346);
or U14058 (N_14058,N_8775,N_10286);
nand U14059 (N_14059,N_9084,N_11997);
nand U14060 (N_14060,N_9272,N_9684);
and U14061 (N_14061,N_9399,N_10443);
and U14062 (N_14062,N_11190,N_10427);
nor U14063 (N_14063,N_10836,N_9600);
nand U14064 (N_14064,N_11578,N_10215);
xor U14065 (N_14065,N_8904,N_11355);
or U14066 (N_14066,N_9230,N_8237);
nor U14067 (N_14067,N_9209,N_8280);
nand U14068 (N_14068,N_10873,N_10174);
and U14069 (N_14069,N_9706,N_10845);
xor U14070 (N_14070,N_10499,N_10187);
nor U14071 (N_14071,N_9024,N_10880);
or U14072 (N_14072,N_9090,N_10330);
xor U14073 (N_14073,N_10544,N_11353);
xor U14074 (N_14074,N_11834,N_8042);
xnor U14075 (N_14075,N_11435,N_10777);
or U14076 (N_14076,N_11134,N_11544);
or U14077 (N_14077,N_10942,N_8694);
and U14078 (N_14078,N_8268,N_11805);
xnor U14079 (N_14079,N_8636,N_10515);
xnor U14080 (N_14080,N_8016,N_8579);
nor U14081 (N_14081,N_8683,N_8427);
and U14082 (N_14082,N_9244,N_8676);
nor U14083 (N_14083,N_10463,N_10530);
nor U14084 (N_14084,N_10351,N_10283);
nor U14085 (N_14085,N_8791,N_10510);
nor U14086 (N_14086,N_8293,N_10799);
xor U14087 (N_14087,N_10321,N_10750);
xor U14088 (N_14088,N_10904,N_8863);
or U14089 (N_14089,N_9742,N_8058);
nor U14090 (N_14090,N_10510,N_8671);
and U14091 (N_14091,N_8987,N_10888);
and U14092 (N_14092,N_9895,N_8154);
xor U14093 (N_14093,N_11706,N_9055);
or U14094 (N_14094,N_9648,N_11178);
nor U14095 (N_14095,N_9179,N_8838);
nand U14096 (N_14096,N_8279,N_8698);
and U14097 (N_14097,N_8266,N_10643);
xor U14098 (N_14098,N_10449,N_8111);
nand U14099 (N_14099,N_10504,N_9073);
or U14100 (N_14100,N_10924,N_10914);
nor U14101 (N_14101,N_11561,N_8263);
nor U14102 (N_14102,N_10098,N_8417);
xnor U14103 (N_14103,N_9338,N_8036);
nand U14104 (N_14104,N_10548,N_8387);
and U14105 (N_14105,N_9723,N_9186);
xnor U14106 (N_14106,N_11039,N_11897);
nand U14107 (N_14107,N_11122,N_10120);
xnor U14108 (N_14108,N_10812,N_8547);
nor U14109 (N_14109,N_11110,N_9639);
or U14110 (N_14110,N_10636,N_9234);
and U14111 (N_14111,N_8746,N_11439);
nor U14112 (N_14112,N_11052,N_11982);
nor U14113 (N_14113,N_9244,N_10324);
or U14114 (N_14114,N_11743,N_9394);
nor U14115 (N_14115,N_9300,N_11386);
xnor U14116 (N_14116,N_11063,N_10771);
or U14117 (N_14117,N_8350,N_10280);
nand U14118 (N_14118,N_9245,N_8911);
and U14119 (N_14119,N_11763,N_10901);
nand U14120 (N_14120,N_10969,N_8718);
xnor U14121 (N_14121,N_8183,N_9897);
nor U14122 (N_14122,N_10000,N_11394);
xor U14123 (N_14123,N_9454,N_10059);
nor U14124 (N_14124,N_11903,N_9461);
and U14125 (N_14125,N_11072,N_11555);
xor U14126 (N_14126,N_11223,N_8955);
or U14127 (N_14127,N_9940,N_9088);
nor U14128 (N_14128,N_8770,N_9636);
xor U14129 (N_14129,N_10568,N_9973);
and U14130 (N_14130,N_10575,N_11596);
xor U14131 (N_14131,N_9774,N_9959);
xnor U14132 (N_14132,N_11009,N_8207);
nor U14133 (N_14133,N_10560,N_8446);
xnor U14134 (N_14134,N_10930,N_10277);
nand U14135 (N_14135,N_11455,N_9185);
or U14136 (N_14136,N_10829,N_10436);
nor U14137 (N_14137,N_10311,N_10198);
xnor U14138 (N_14138,N_8456,N_11230);
nand U14139 (N_14139,N_10018,N_11304);
or U14140 (N_14140,N_10184,N_10930);
xor U14141 (N_14141,N_9267,N_11784);
or U14142 (N_14142,N_11315,N_9109);
and U14143 (N_14143,N_8741,N_11475);
xnor U14144 (N_14144,N_9611,N_11234);
and U14145 (N_14145,N_11350,N_9749);
or U14146 (N_14146,N_10969,N_11245);
nor U14147 (N_14147,N_8622,N_11194);
xor U14148 (N_14148,N_8729,N_9932);
nor U14149 (N_14149,N_9768,N_10575);
nor U14150 (N_14150,N_10805,N_10465);
nand U14151 (N_14151,N_10035,N_8004);
and U14152 (N_14152,N_11870,N_9910);
nor U14153 (N_14153,N_9949,N_11323);
or U14154 (N_14154,N_8213,N_11726);
xor U14155 (N_14155,N_8221,N_10104);
xnor U14156 (N_14156,N_11176,N_9368);
xnor U14157 (N_14157,N_11783,N_11376);
xor U14158 (N_14158,N_10797,N_11199);
nor U14159 (N_14159,N_11670,N_8470);
and U14160 (N_14160,N_10358,N_8062);
and U14161 (N_14161,N_8148,N_9928);
or U14162 (N_14162,N_11854,N_8141);
xnor U14163 (N_14163,N_8147,N_9732);
xor U14164 (N_14164,N_10201,N_9089);
nor U14165 (N_14165,N_9470,N_8395);
nand U14166 (N_14166,N_11995,N_10933);
xor U14167 (N_14167,N_9889,N_8756);
xnor U14168 (N_14168,N_9011,N_8462);
nor U14169 (N_14169,N_9775,N_11254);
nor U14170 (N_14170,N_11015,N_8483);
nor U14171 (N_14171,N_8037,N_8463);
or U14172 (N_14172,N_10392,N_10988);
xnor U14173 (N_14173,N_9283,N_10482);
nand U14174 (N_14174,N_9544,N_11675);
nand U14175 (N_14175,N_11402,N_10267);
nor U14176 (N_14176,N_9239,N_9755);
or U14177 (N_14177,N_9846,N_8372);
nand U14178 (N_14178,N_8906,N_10603);
nand U14179 (N_14179,N_9080,N_8809);
nor U14180 (N_14180,N_9314,N_8398);
nand U14181 (N_14181,N_9335,N_10269);
or U14182 (N_14182,N_8624,N_8369);
xnor U14183 (N_14183,N_11877,N_10378);
xnor U14184 (N_14184,N_8313,N_11258);
nor U14185 (N_14185,N_8864,N_11391);
xnor U14186 (N_14186,N_8400,N_8062);
xor U14187 (N_14187,N_11253,N_9556);
nor U14188 (N_14188,N_8950,N_8831);
nor U14189 (N_14189,N_10657,N_8348);
nand U14190 (N_14190,N_11250,N_8393);
xor U14191 (N_14191,N_11883,N_11803);
nor U14192 (N_14192,N_10008,N_11837);
nand U14193 (N_14193,N_8021,N_11501);
nor U14194 (N_14194,N_11296,N_11377);
xor U14195 (N_14195,N_9585,N_11114);
xnor U14196 (N_14196,N_8523,N_11822);
xnor U14197 (N_14197,N_10814,N_10227);
and U14198 (N_14198,N_10321,N_9487);
and U14199 (N_14199,N_9792,N_11546);
or U14200 (N_14200,N_9491,N_8684);
or U14201 (N_14201,N_10477,N_11361);
nand U14202 (N_14202,N_10954,N_10596);
xor U14203 (N_14203,N_9649,N_8790);
nand U14204 (N_14204,N_10531,N_9400);
nand U14205 (N_14205,N_11539,N_11016);
or U14206 (N_14206,N_10669,N_9611);
and U14207 (N_14207,N_8619,N_10456);
and U14208 (N_14208,N_9797,N_11162);
or U14209 (N_14209,N_11044,N_10469);
xnor U14210 (N_14210,N_10626,N_9285);
nor U14211 (N_14211,N_9631,N_8195);
nand U14212 (N_14212,N_9090,N_8620);
or U14213 (N_14213,N_10632,N_11492);
nor U14214 (N_14214,N_9319,N_11176);
xor U14215 (N_14215,N_9343,N_8415);
nor U14216 (N_14216,N_10721,N_10877);
or U14217 (N_14217,N_11866,N_9714);
nand U14218 (N_14218,N_10634,N_9764);
xnor U14219 (N_14219,N_9757,N_8811);
and U14220 (N_14220,N_9141,N_9368);
nand U14221 (N_14221,N_10333,N_8508);
or U14222 (N_14222,N_10320,N_9893);
nor U14223 (N_14223,N_11706,N_9062);
or U14224 (N_14224,N_8164,N_9776);
nand U14225 (N_14225,N_8101,N_11398);
xor U14226 (N_14226,N_11518,N_10393);
nor U14227 (N_14227,N_11979,N_8026);
nand U14228 (N_14228,N_8621,N_10079);
xnor U14229 (N_14229,N_10360,N_11464);
nor U14230 (N_14230,N_11321,N_11217);
xor U14231 (N_14231,N_9239,N_9899);
and U14232 (N_14232,N_10585,N_9358);
and U14233 (N_14233,N_9634,N_8424);
nand U14234 (N_14234,N_9457,N_9517);
xnor U14235 (N_14235,N_10555,N_9244);
nor U14236 (N_14236,N_11534,N_10164);
and U14237 (N_14237,N_10257,N_9150);
and U14238 (N_14238,N_9050,N_8658);
nand U14239 (N_14239,N_11167,N_11374);
and U14240 (N_14240,N_8802,N_8465);
xnor U14241 (N_14241,N_9342,N_11636);
nand U14242 (N_14242,N_10484,N_10725);
nand U14243 (N_14243,N_10186,N_11622);
or U14244 (N_14244,N_9423,N_9374);
nand U14245 (N_14245,N_9138,N_10207);
nor U14246 (N_14246,N_8925,N_8890);
nand U14247 (N_14247,N_9271,N_10824);
nand U14248 (N_14248,N_9033,N_11787);
and U14249 (N_14249,N_9411,N_8090);
or U14250 (N_14250,N_8367,N_10044);
xnor U14251 (N_14251,N_11459,N_9351);
nand U14252 (N_14252,N_9281,N_8944);
xor U14253 (N_14253,N_10301,N_8176);
or U14254 (N_14254,N_8323,N_11418);
and U14255 (N_14255,N_8908,N_11849);
xnor U14256 (N_14256,N_9110,N_10684);
xnor U14257 (N_14257,N_11137,N_10469);
nor U14258 (N_14258,N_9236,N_10129);
nor U14259 (N_14259,N_8256,N_8921);
nand U14260 (N_14260,N_9566,N_11828);
nor U14261 (N_14261,N_11351,N_9675);
and U14262 (N_14262,N_11816,N_9220);
nor U14263 (N_14263,N_9874,N_9637);
nor U14264 (N_14264,N_8035,N_10187);
and U14265 (N_14265,N_8195,N_11086);
nand U14266 (N_14266,N_9409,N_10413);
or U14267 (N_14267,N_11301,N_8839);
nand U14268 (N_14268,N_11089,N_8495);
or U14269 (N_14269,N_11245,N_11892);
and U14270 (N_14270,N_10019,N_10333);
nand U14271 (N_14271,N_10194,N_10673);
xnor U14272 (N_14272,N_9712,N_11192);
xor U14273 (N_14273,N_10324,N_11242);
nand U14274 (N_14274,N_9342,N_10016);
xnor U14275 (N_14275,N_8736,N_8519);
or U14276 (N_14276,N_9954,N_10247);
or U14277 (N_14277,N_9045,N_8931);
nor U14278 (N_14278,N_10297,N_9940);
and U14279 (N_14279,N_10143,N_11468);
and U14280 (N_14280,N_9807,N_11143);
and U14281 (N_14281,N_10489,N_8848);
or U14282 (N_14282,N_10432,N_9316);
or U14283 (N_14283,N_9898,N_9862);
nand U14284 (N_14284,N_11116,N_10396);
or U14285 (N_14285,N_8361,N_11976);
xor U14286 (N_14286,N_10205,N_9937);
nand U14287 (N_14287,N_11746,N_9956);
and U14288 (N_14288,N_8412,N_10885);
nor U14289 (N_14289,N_9382,N_9485);
nor U14290 (N_14290,N_11561,N_10333);
nand U14291 (N_14291,N_11651,N_11507);
xor U14292 (N_14292,N_11990,N_10311);
nand U14293 (N_14293,N_11311,N_10035);
xnor U14294 (N_14294,N_11761,N_8169);
and U14295 (N_14295,N_8457,N_11383);
and U14296 (N_14296,N_11888,N_10985);
or U14297 (N_14297,N_8328,N_9642);
nor U14298 (N_14298,N_10863,N_10945);
nor U14299 (N_14299,N_8346,N_9037);
or U14300 (N_14300,N_10369,N_10254);
and U14301 (N_14301,N_11624,N_8886);
or U14302 (N_14302,N_8854,N_11999);
or U14303 (N_14303,N_10099,N_10439);
or U14304 (N_14304,N_9237,N_9706);
nand U14305 (N_14305,N_9521,N_11786);
and U14306 (N_14306,N_11904,N_9623);
or U14307 (N_14307,N_10938,N_11224);
nand U14308 (N_14308,N_8007,N_9087);
and U14309 (N_14309,N_8086,N_11743);
nand U14310 (N_14310,N_10617,N_8220);
nor U14311 (N_14311,N_9954,N_10964);
and U14312 (N_14312,N_8319,N_10121);
nand U14313 (N_14313,N_10113,N_9014);
nand U14314 (N_14314,N_8493,N_9237);
nor U14315 (N_14315,N_9694,N_8896);
or U14316 (N_14316,N_10141,N_9773);
or U14317 (N_14317,N_9145,N_9996);
xor U14318 (N_14318,N_9390,N_9186);
nand U14319 (N_14319,N_10487,N_8341);
nand U14320 (N_14320,N_10058,N_8795);
nand U14321 (N_14321,N_10978,N_8840);
xor U14322 (N_14322,N_11346,N_10832);
or U14323 (N_14323,N_9122,N_10655);
nor U14324 (N_14324,N_10480,N_10016);
nand U14325 (N_14325,N_11896,N_9660);
and U14326 (N_14326,N_11614,N_9303);
or U14327 (N_14327,N_10564,N_10624);
or U14328 (N_14328,N_9413,N_10026);
or U14329 (N_14329,N_8021,N_9716);
and U14330 (N_14330,N_10823,N_10147);
and U14331 (N_14331,N_9979,N_10770);
nor U14332 (N_14332,N_10679,N_8459);
or U14333 (N_14333,N_9174,N_8952);
xnor U14334 (N_14334,N_10499,N_9115);
nand U14335 (N_14335,N_11195,N_9267);
or U14336 (N_14336,N_8720,N_8075);
nand U14337 (N_14337,N_10433,N_9447);
nor U14338 (N_14338,N_9333,N_11894);
nand U14339 (N_14339,N_9524,N_10506);
or U14340 (N_14340,N_8594,N_11357);
and U14341 (N_14341,N_11017,N_10081);
nand U14342 (N_14342,N_10519,N_10595);
nand U14343 (N_14343,N_11369,N_10406);
or U14344 (N_14344,N_9769,N_8119);
xnor U14345 (N_14345,N_9143,N_9066);
nor U14346 (N_14346,N_11136,N_10486);
and U14347 (N_14347,N_10234,N_8574);
and U14348 (N_14348,N_11703,N_11244);
and U14349 (N_14349,N_9835,N_9242);
nor U14350 (N_14350,N_10045,N_10429);
or U14351 (N_14351,N_11957,N_8837);
or U14352 (N_14352,N_11207,N_9282);
xor U14353 (N_14353,N_10361,N_10138);
xnor U14354 (N_14354,N_8407,N_10362);
xnor U14355 (N_14355,N_8912,N_11328);
and U14356 (N_14356,N_11342,N_9905);
nor U14357 (N_14357,N_10242,N_11729);
nand U14358 (N_14358,N_8169,N_10693);
nor U14359 (N_14359,N_8925,N_8098);
or U14360 (N_14360,N_11867,N_8665);
and U14361 (N_14361,N_9068,N_10931);
xnor U14362 (N_14362,N_8680,N_9144);
or U14363 (N_14363,N_11746,N_8766);
nand U14364 (N_14364,N_8526,N_11583);
and U14365 (N_14365,N_9814,N_11984);
nor U14366 (N_14366,N_11750,N_10831);
or U14367 (N_14367,N_10587,N_10037);
nor U14368 (N_14368,N_8580,N_8802);
xor U14369 (N_14369,N_11522,N_9999);
nand U14370 (N_14370,N_8100,N_8658);
and U14371 (N_14371,N_11771,N_8021);
or U14372 (N_14372,N_11384,N_10677);
and U14373 (N_14373,N_9582,N_9339);
or U14374 (N_14374,N_10883,N_8462);
xor U14375 (N_14375,N_11647,N_11813);
nor U14376 (N_14376,N_11212,N_11673);
nand U14377 (N_14377,N_9892,N_11822);
nor U14378 (N_14378,N_10015,N_9196);
nand U14379 (N_14379,N_11847,N_10746);
or U14380 (N_14380,N_8464,N_10995);
nor U14381 (N_14381,N_10877,N_10164);
nor U14382 (N_14382,N_11398,N_8367);
nand U14383 (N_14383,N_9716,N_9990);
nor U14384 (N_14384,N_8555,N_9488);
and U14385 (N_14385,N_9727,N_10928);
and U14386 (N_14386,N_8764,N_8749);
or U14387 (N_14387,N_8491,N_10367);
nand U14388 (N_14388,N_8856,N_8428);
nand U14389 (N_14389,N_9603,N_10033);
xor U14390 (N_14390,N_10571,N_11764);
nor U14391 (N_14391,N_9895,N_11352);
or U14392 (N_14392,N_9611,N_8437);
nor U14393 (N_14393,N_8912,N_10580);
nor U14394 (N_14394,N_8316,N_9450);
or U14395 (N_14395,N_10198,N_10974);
nor U14396 (N_14396,N_8966,N_9742);
nand U14397 (N_14397,N_10632,N_10201);
nor U14398 (N_14398,N_10992,N_8953);
and U14399 (N_14399,N_8897,N_10336);
xor U14400 (N_14400,N_10228,N_8394);
xor U14401 (N_14401,N_10032,N_9481);
nor U14402 (N_14402,N_11966,N_9957);
nand U14403 (N_14403,N_11591,N_11659);
xor U14404 (N_14404,N_11523,N_8349);
or U14405 (N_14405,N_10488,N_11357);
and U14406 (N_14406,N_9303,N_8708);
nand U14407 (N_14407,N_9885,N_9276);
xnor U14408 (N_14408,N_8187,N_10050);
or U14409 (N_14409,N_10074,N_8785);
nand U14410 (N_14410,N_11154,N_11629);
or U14411 (N_14411,N_11057,N_10869);
nor U14412 (N_14412,N_11970,N_10687);
nor U14413 (N_14413,N_9834,N_8858);
or U14414 (N_14414,N_9020,N_9009);
nor U14415 (N_14415,N_11579,N_11652);
nand U14416 (N_14416,N_9020,N_9405);
nor U14417 (N_14417,N_11679,N_9163);
or U14418 (N_14418,N_10496,N_10105);
or U14419 (N_14419,N_11796,N_11441);
xnor U14420 (N_14420,N_9678,N_9981);
nand U14421 (N_14421,N_8467,N_10617);
xor U14422 (N_14422,N_11429,N_11672);
nor U14423 (N_14423,N_8582,N_11874);
xor U14424 (N_14424,N_9622,N_10004);
nand U14425 (N_14425,N_10827,N_11606);
and U14426 (N_14426,N_11983,N_9240);
xor U14427 (N_14427,N_9910,N_10114);
xor U14428 (N_14428,N_8322,N_8641);
or U14429 (N_14429,N_11919,N_9065);
or U14430 (N_14430,N_11133,N_11434);
xor U14431 (N_14431,N_8171,N_11025);
nand U14432 (N_14432,N_11177,N_11362);
or U14433 (N_14433,N_8690,N_8085);
or U14434 (N_14434,N_9907,N_9234);
or U14435 (N_14435,N_8756,N_8690);
xnor U14436 (N_14436,N_10342,N_11459);
nor U14437 (N_14437,N_10721,N_10108);
or U14438 (N_14438,N_9667,N_8065);
and U14439 (N_14439,N_11706,N_9415);
xor U14440 (N_14440,N_9201,N_10919);
or U14441 (N_14441,N_11261,N_11414);
nor U14442 (N_14442,N_9130,N_10159);
xnor U14443 (N_14443,N_11959,N_8286);
xnor U14444 (N_14444,N_8260,N_11413);
or U14445 (N_14445,N_11635,N_9397);
and U14446 (N_14446,N_10019,N_8243);
nand U14447 (N_14447,N_8650,N_8473);
nand U14448 (N_14448,N_9153,N_10361);
xor U14449 (N_14449,N_8737,N_8336);
or U14450 (N_14450,N_11202,N_10320);
xor U14451 (N_14451,N_8093,N_8058);
xnor U14452 (N_14452,N_10604,N_11028);
nand U14453 (N_14453,N_8616,N_10555);
or U14454 (N_14454,N_11864,N_11537);
nor U14455 (N_14455,N_10963,N_9041);
nand U14456 (N_14456,N_10898,N_10426);
nor U14457 (N_14457,N_11238,N_8070);
xnor U14458 (N_14458,N_11679,N_8747);
xnor U14459 (N_14459,N_9710,N_9842);
or U14460 (N_14460,N_9385,N_11126);
nor U14461 (N_14461,N_10030,N_10294);
or U14462 (N_14462,N_11314,N_10440);
nand U14463 (N_14463,N_8706,N_9622);
xnor U14464 (N_14464,N_8143,N_9390);
nand U14465 (N_14465,N_10910,N_8065);
xnor U14466 (N_14466,N_9889,N_8265);
nor U14467 (N_14467,N_9036,N_8325);
and U14468 (N_14468,N_8088,N_11320);
xor U14469 (N_14469,N_9338,N_8441);
nor U14470 (N_14470,N_8741,N_10915);
nand U14471 (N_14471,N_10332,N_10434);
nand U14472 (N_14472,N_9963,N_11155);
or U14473 (N_14473,N_11638,N_8669);
nand U14474 (N_14474,N_9346,N_9798);
nor U14475 (N_14475,N_9925,N_9914);
nand U14476 (N_14476,N_10101,N_8131);
xor U14477 (N_14477,N_9543,N_10413);
or U14478 (N_14478,N_9865,N_10146);
nand U14479 (N_14479,N_8750,N_8076);
xor U14480 (N_14480,N_8019,N_10539);
nand U14481 (N_14481,N_10590,N_9954);
or U14482 (N_14482,N_9669,N_10584);
nor U14483 (N_14483,N_9344,N_10293);
or U14484 (N_14484,N_11200,N_8712);
xor U14485 (N_14485,N_10845,N_8800);
xnor U14486 (N_14486,N_10530,N_8313);
nand U14487 (N_14487,N_11746,N_10968);
xor U14488 (N_14488,N_8223,N_10296);
or U14489 (N_14489,N_8372,N_8729);
or U14490 (N_14490,N_10715,N_9133);
or U14491 (N_14491,N_10922,N_9370);
xnor U14492 (N_14492,N_10614,N_10944);
or U14493 (N_14493,N_9957,N_8296);
nor U14494 (N_14494,N_8710,N_9573);
and U14495 (N_14495,N_8430,N_10128);
nor U14496 (N_14496,N_9006,N_11991);
xor U14497 (N_14497,N_9217,N_10032);
or U14498 (N_14498,N_10688,N_9185);
or U14499 (N_14499,N_11658,N_9459);
and U14500 (N_14500,N_11152,N_9013);
nor U14501 (N_14501,N_9208,N_9879);
nor U14502 (N_14502,N_10616,N_9996);
nand U14503 (N_14503,N_11248,N_11618);
nor U14504 (N_14504,N_10943,N_11843);
and U14505 (N_14505,N_11288,N_8832);
nand U14506 (N_14506,N_8655,N_8946);
nor U14507 (N_14507,N_10035,N_11263);
nand U14508 (N_14508,N_11936,N_9197);
and U14509 (N_14509,N_10860,N_10118);
and U14510 (N_14510,N_11170,N_8723);
nand U14511 (N_14511,N_8698,N_9394);
xnor U14512 (N_14512,N_10954,N_8900);
nor U14513 (N_14513,N_11956,N_11722);
nand U14514 (N_14514,N_9987,N_8932);
or U14515 (N_14515,N_10551,N_11640);
xnor U14516 (N_14516,N_8713,N_9020);
nand U14517 (N_14517,N_10388,N_9456);
nand U14518 (N_14518,N_8359,N_10642);
or U14519 (N_14519,N_9958,N_9896);
nand U14520 (N_14520,N_9811,N_9353);
or U14521 (N_14521,N_11630,N_9220);
and U14522 (N_14522,N_8319,N_10641);
nor U14523 (N_14523,N_8584,N_11257);
nand U14524 (N_14524,N_8595,N_11551);
and U14525 (N_14525,N_9663,N_8659);
and U14526 (N_14526,N_8199,N_9668);
xor U14527 (N_14527,N_11376,N_10664);
or U14528 (N_14528,N_8696,N_11974);
xor U14529 (N_14529,N_8151,N_8762);
nand U14530 (N_14530,N_11744,N_11136);
and U14531 (N_14531,N_10102,N_8838);
or U14532 (N_14532,N_9644,N_9486);
or U14533 (N_14533,N_9095,N_8127);
or U14534 (N_14534,N_9090,N_8787);
xor U14535 (N_14535,N_8367,N_10486);
nor U14536 (N_14536,N_10633,N_11419);
and U14537 (N_14537,N_8759,N_10128);
nor U14538 (N_14538,N_10072,N_9775);
nor U14539 (N_14539,N_9138,N_10690);
nor U14540 (N_14540,N_10534,N_9734);
and U14541 (N_14541,N_9451,N_9588);
nand U14542 (N_14542,N_11401,N_8279);
nor U14543 (N_14543,N_8646,N_10775);
and U14544 (N_14544,N_9170,N_9009);
xor U14545 (N_14545,N_11919,N_8819);
xor U14546 (N_14546,N_8087,N_10162);
nor U14547 (N_14547,N_9211,N_10511);
nand U14548 (N_14548,N_10154,N_10217);
nand U14549 (N_14549,N_8783,N_9472);
nand U14550 (N_14550,N_11526,N_11707);
and U14551 (N_14551,N_9811,N_8929);
or U14552 (N_14552,N_8443,N_9373);
or U14553 (N_14553,N_11895,N_9572);
nand U14554 (N_14554,N_10118,N_9948);
xor U14555 (N_14555,N_9413,N_11869);
nand U14556 (N_14556,N_8880,N_10113);
or U14557 (N_14557,N_8345,N_9007);
nor U14558 (N_14558,N_10892,N_9639);
and U14559 (N_14559,N_9855,N_10600);
or U14560 (N_14560,N_9220,N_11310);
nor U14561 (N_14561,N_11660,N_10540);
nand U14562 (N_14562,N_9063,N_11406);
nor U14563 (N_14563,N_10169,N_9558);
or U14564 (N_14564,N_8853,N_10071);
nor U14565 (N_14565,N_10127,N_11538);
nand U14566 (N_14566,N_9156,N_10882);
nand U14567 (N_14567,N_11593,N_11485);
and U14568 (N_14568,N_11941,N_11278);
or U14569 (N_14569,N_11941,N_10593);
nor U14570 (N_14570,N_10203,N_10219);
nor U14571 (N_14571,N_9375,N_8160);
and U14572 (N_14572,N_9953,N_10344);
and U14573 (N_14573,N_9065,N_8519);
xor U14574 (N_14574,N_11815,N_8309);
nand U14575 (N_14575,N_9990,N_9382);
nor U14576 (N_14576,N_10890,N_8311);
or U14577 (N_14577,N_11444,N_11127);
nand U14578 (N_14578,N_11645,N_10673);
nor U14579 (N_14579,N_8884,N_9464);
and U14580 (N_14580,N_8611,N_9916);
nand U14581 (N_14581,N_10546,N_9108);
or U14582 (N_14582,N_10394,N_10573);
xor U14583 (N_14583,N_10457,N_8095);
xor U14584 (N_14584,N_9747,N_8170);
nand U14585 (N_14585,N_9460,N_11429);
nand U14586 (N_14586,N_9065,N_10751);
xnor U14587 (N_14587,N_9950,N_9476);
and U14588 (N_14588,N_11906,N_11405);
or U14589 (N_14589,N_10732,N_10374);
nand U14590 (N_14590,N_11196,N_9938);
or U14591 (N_14591,N_11635,N_8466);
nand U14592 (N_14592,N_8108,N_9480);
nand U14593 (N_14593,N_8370,N_10077);
xnor U14594 (N_14594,N_10531,N_9147);
nor U14595 (N_14595,N_8410,N_11627);
nor U14596 (N_14596,N_10741,N_11198);
or U14597 (N_14597,N_9148,N_11971);
nor U14598 (N_14598,N_9945,N_10773);
nand U14599 (N_14599,N_8198,N_11589);
nand U14600 (N_14600,N_8527,N_9680);
or U14601 (N_14601,N_10881,N_11517);
nand U14602 (N_14602,N_8179,N_10311);
xor U14603 (N_14603,N_9096,N_8733);
xnor U14604 (N_14604,N_11099,N_11798);
nor U14605 (N_14605,N_9947,N_9806);
nor U14606 (N_14606,N_10220,N_11031);
xor U14607 (N_14607,N_9304,N_11406);
nor U14608 (N_14608,N_9326,N_11217);
and U14609 (N_14609,N_8393,N_11505);
nor U14610 (N_14610,N_8457,N_9095);
nor U14611 (N_14611,N_8704,N_11010);
xnor U14612 (N_14612,N_10252,N_11870);
nor U14613 (N_14613,N_9204,N_9537);
nand U14614 (N_14614,N_8417,N_11336);
nor U14615 (N_14615,N_9257,N_10473);
xor U14616 (N_14616,N_11530,N_9317);
and U14617 (N_14617,N_8165,N_11722);
or U14618 (N_14618,N_9262,N_10679);
and U14619 (N_14619,N_9398,N_9115);
xor U14620 (N_14620,N_10999,N_8980);
and U14621 (N_14621,N_9535,N_9337);
or U14622 (N_14622,N_8929,N_10025);
or U14623 (N_14623,N_11256,N_9775);
or U14624 (N_14624,N_9479,N_11462);
and U14625 (N_14625,N_11904,N_8714);
and U14626 (N_14626,N_10298,N_10388);
or U14627 (N_14627,N_9703,N_8872);
and U14628 (N_14628,N_11469,N_10753);
or U14629 (N_14629,N_9302,N_11505);
nand U14630 (N_14630,N_8060,N_9903);
or U14631 (N_14631,N_9322,N_11462);
or U14632 (N_14632,N_10894,N_10025);
and U14633 (N_14633,N_10395,N_10718);
or U14634 (N_14634,N_11437,N_11360);
or U14635 (N_14635,N_9874,N_10201);
nand U14636 (N_14636,N_10707,N_11142);
nand U14637 (N_14637,N_8204,N_11178);
nor U14638 (N_14638,N_10657,N_10246);
nand U14639 (N_14639,N_8372,N_9461);
nor U14640 (N_14640,N_8883,N_9962);
nand U14641 (N_14641,N_9059,N_9865);
or U14642 (N_14642,N_11867,N_11161);
nor U14643 (N_14643,N_11138,N_8775);
nor U14644 (N_14644,N_11408,N_11372);
or U14645 (N_14645,N_10556,N_9903);
nand U14646 (N_14646,N_11955,N_10073);
or U14647 (N_14647,N_9778,N_10755);
and U14648 (N_14648,N_9538,N_9204);
nor U14649 (N_14649,N_8423,N_9489);
nor U14650 (N_14650,N_10180,N_11408);
and U14651 (N_14651,N_11022,N_10707);
xnor U14652 (N_14652,N_11341,N_10425);
and U14653 (N_14653,N_11973,N_9986);
or U14654 (N_14654,N_10665,N_9982);
nor U14655 (N_14655,N_11502,N_9832);
and U14656 (N_14656,N_11196,N_8850);
nand U14657 (N_14657,N_11680,N_10932);
and U14658 (N_14658,N_9059,N_11458);
nand U14659 (N_14659,N_8874,N_10392);
nor U14660 (N_14660,N_10392,N_8665);
and U14661 (N_14661,N_8352,N_11945);
and U14662 (N_14662,N_11169,N_9531);
nand U14663 (N_14663,N_11868,N_8840);
xor U14664 (N_14664,N_9022,N_10342);
and U14665 (N_14665,N_8360,N_8629);
nand U14666 (N_14666,N_11506,N_10364);
xnor U14667 (N_14667,N_11732,N_8291);
nand U14668 (N_14668,N_9271,N_8483);
nand U14669 (N_14669,N_8024,N_9035);
or U14670 (N_14670,N_8357,N_8114);
xnor U14671 (N_14671,N_9144,N_10465);
or U14672 (N_14672,N_9769,N_9041);
nor U14673 (N_14673,N_11948,N_10828);
nand U14674 (N_14674,N_10758,N_10053);
nand U14675 (N_14675,N_10243,N_9379);
xnor U14676 (N_14676,N_10519,N_11381);
nand U14677 (N_14677,N_10929,N_8886);
and U14678 (N_14678,N_10060,N_11623);
and U14679 (N_14679,N_9238,N_10507);
nor U14680 (N_14680,N_10952,N_11736);
nor U14681 (N_14681,N_10538,N_8201);
and U14682 (N_14682,N_8708,N_10224);
or U14683 (N_14683,N_8986,N_8031);
nor U14684 (N_14684,N_8612,N_8521);
or U14685 (N_14685,N_10777,N_9107);
xnor U14686 (N_14686,N_8911,N_10821);
nand U14687 (N_14687,N_10083,N_10121);
or U14688 (N_14688,N_11374,N_11311);
nor U14689 (N_14689,N_9902,N_9540);
or U14690 (N_14690,N_11910,N_9130);
or U14691 (N_14691,N_8375,N_10784);
nor U14692 (N_14692,N_11282,N_10974);
or U14693 (N_14693,N_9506,N_8581);
nand U14694 (N_14694,N_9957,N_9304);
xnor U14695 (N_14695,N_8226,N_9402);
nor U14696 (N_14696,N_10109,N_11942);
nor U14697 (N_14697,N_10208,N_9267);
and U14698 (N_14698,N_10030,N_10006);
xnor U14699 (N_14699,N_9883,N_8602);
and U14700 (N_14700,N_11338,N_8025);
or U14701 (N_14701,N_9914,N_8200);
xor U14702 (N_14702,N_10618,N_8894);
nor U14703 (N_14703,N_10507,N_10630);
or U14704 (N_14704,N_10005,N_9271);
xor U14705 (N_14705,N_10582,N_11047);
nor U14706 (N_14706,N_11373,N_8646);
nand U14707 (N_14707,N_8619,N_9955);
and U14708 (N_14708,N_8974,N_9857);
nor U14709 (N_14709,N_11633,N_10087);
xnor U14710 (N_14710,N_10097,N_9687);
nand U14711 (N_14711,N_11537,N_9786);
and U14712 (N_14712,N_10373,N_8727);
or U14713 (N_14713,N_8720,N_8128);
nand U14714 (N_14714,N_11895,N_8814);
xor U14715 (N_14715,N_9794,N_9999);
xor U14716 (N_14716,N_9708,N_8336);
or U14717 (N_14717,N_10332,N_10767);
nor U14718 (N_14718,N_9187,N_11770);
nand U14719 (N_14719,N_8196,N_8332);
or U14720 (N_14720,N_9912,N_9459);
nand U14721 (N_14721,N_9074,N_10126);
nand U14722 (N_14722,N_11915,N_11715);
xor U14723 (N_14723,N_8419,N_9891);
xnor U14724 (N_14724,N_11224,N_8019);
or U14725 (N_14725,N_10108,N_11216);
or U14726 (N_14726,N_10241,N_9734);
nand U14727 (N_14727,N_9697,N_11214);
nor U14728 (N_14728,N_11555,N_10352);
nand U14729 (N_14729,N_8524,N_9529);
nand U14730 (N_14730,N_9931,N_9682);
xnor U14731 (N_14731,N_9971,N_10036);
or U14732 (N_14732,N_11565,N_11779);
and U14733 (N_14733,N_8439,N_11533);
nor U14734 (N_14734,N_8026,N_8266);
nand U14735 (N_14735,N_9982,N_8177);
and U14736 (N_14736,N_9050,N_9271);
and U14737 (N_14737,N_9493,N_9929);
or U14738 (N_14738,N_10756,N_8382);
or U14739 (N_14739,N_9121,N_8362);
and U14740 (N_14740,N_10338,N_11447);
xor U14741 (N_14741,N_9724,N_10791);
nor U14742 (N_14742,N_10223,N_9774);
nor U14743 (N_14743,N_9624,N_10415);
and U14744 (N_14744,N_9876,N_10168);
nor U14745 (N_14745,N_8836,N_8258);
xnor U14746 (N_14746,N_9145,N_11062);
nand U14747 (N_14747,N_9437,N_10403);
nor U14748 (N_14748,N_10265,N_9194);
xor U14749 (N_14749,N_10943,N_11031);
xor U14750 (N_14750,N_8040,N_10701);
and U14751 (N_14751,N_11119,N_8172);
xnor U14752 (N_14752,N_10048,N_9877);
and U14753 (N_14753,N_9827,N_11679);
or U14754 (N_14754,N_10926,N_11232);
nand U14755 (N_14755,N_11729,N_11171);
and U14756 (N_14756,N_9223,N_11195);
xor U14757 (N_14757,N_9104,N_9839);
nor U14758 (N_14758,N_9286,N_10627);
nor U14759 (N_14759,N_10791,N_8042);
xor U14760 (N_14760,N_11661,N_9136);
nor U14761 (N_14761,N_10271,N_10876);
xor U14762 (N_14762,N_10196,N_8490);
and U14763 (N_14763,N_10834,N_9121);
nand U14764 (N_14764,N_11130,N_11267);
nor U14765 (N_14765,N_9072,N_10757);
nand U14766 (N_14766,N_8864,N_8623);
and U14767 (N_14767,N_10874,N_9280);
nor U14768 (N_14768,N_11309,N_9921);
xor U14769 (N_14769,N_11975,N_8707);
nor U14770 (N_14770,N_8071,N_11715);
or U14771 (N_14771,N_9663,N_11113);
xor U14772 (N_14772,N_8878,N_10947);
and U14773 (N_14773,N_9761,N_9827);
and U14774 (N_14774,N_9347,N_10706);
or U14775 (N_14775,N_9636,N_8522);
nor U14776 (N_14776,N_11534,N_11200);
or U14777 (N_14777,N_9014,N_10147);
nor U14778 (N_14778,N_11321,N_9574);
and U14779 (N_14779,N_10310,N_11225);
xnor U14780 (N_14780,N_10479,N_9083);
xor U14781 (N_14781,N_8782,N_8063);
nor U14782 (N_14782,N_11080,N_8294);
and U14783 (N_14783,N_9380,N_10648);
nand U14784 (N_14784,N_9123,N_8201);
nor U14785 (N_14785,N_8839,N_8681);
nor U14786 (N_14786,N_10689,N_11794);
nor U14787 (N_14787,N_8178,N_8902);
nand U14788 (N_14788,N_11738,N_11554);
nor U14789 (N_14789,N_8672,N_10174);
and U14790 (N_14790,N_11922,N_10954);
nor U14791 (N_14791,N_8850,N_9078);
nand U14792 (N_14792,N_11526,N_11075);
nor U14793 (N_14793,N_8240,N_11545);
and U14794 (N_14794,N_10673,N_10945);
nand U14795 (N_14795,N_9248,N_10408);
nor U14796 (N_14796,N_11419,N_8222);
nand U14797 (N_14797,N_10777,N_10066);
or U14798 (N_14798,N_11678,N_9690);
nor U14799 (N_14799,N_9595,N_9351);
or U14800 (N_14800,N_10286,N_8633);
nand U14801 (N_14801,N_8835,N_9456);
nand U14802 (N_14802,N_10197,N_9252);
and U14803 (N_14803,N_9685,N_9468);
or U14804 (N_14804,N_8088,N_8232);
and U14805 (N_14805,N_9330,N_8602);
nor U14806 (N_14806,N_9992,N_10966);
or U14807 (N_14807,N_9773,N_10320);
xor U14808 (N_14808,N_9755,N_9347);
and U14809 (N_14809,N_11486,N_10769);
or U14810 (N_14810,N_10553,N_11836);
and U14811 (N_14811,N_10254,N_8442);
nor U14812 (N_14812,N_9807,N_8290);
or U14813 (N_14813,N_11100,N_10708);
nor U14814 (N_14814,N_11862,N_8315);
and U14815 (N_14815,N_8337,N_8514);
or U14816 (N_14816,N_8745,N_9197);
or U14817 (N_14817,N_11500,N_11640);
or U14818 (N_14818,N_9635,N_8985);
or U14819 (N_14819,N_11524,N_11831);
and U14820 (N_14820,N_8190,N_8904);
nor U14821 (N_14821,N_9900,N_8429);
xnor U14822 (N_14822,N_8003,N_11991);
xnor U14823 (N_14823,N_10062,N_8111);
or U14824 (N_14824,N_8354,N_8891);
xnor U14825 (N_14825,N_10413,N_11843);
and U14826 (N_14826,N_10129,N_11968);
nor U14827 (N_14827,N_9127,N_10593);
nor U14828 (N_14828,N_11873,N_11971);
xnor U14829 (N_14829,N_8794,N_10262);
or U14830 (N_14830,N_10448,N_11951);
xnor U14831 (N_14831,N_10260,N_9755);
nor U14832 (N_14832,N_10481,N_8476);
nor U14833 (N_14833,N_8909,N_8905);
nand U14834 (N_14834,N_8320,N_8188);
xor U14835 (N_14835,N_10270,N_11152);
nand U14836 (N_14836,N_11946,N_10405);
nand U14837 (N_14837,N_9211,N_8447);
nand U14838 (N_14838,N_11872,N_8507);
or U14839 (N_14839,N_8573,N_8476);
nor U14840 (N_14840,N_10985,N_10012);
nand U14841 (N_14841,N_10459,N_8596);
or U14842 (N_14842,N_11745,N_11853);
nor U14843 (N_14843,N_9622,N_11253);
xor U14844 (N_14844,N_8276,N_8083);
nand U14845 (N_14845,N_9278,N_10913);
nor U14846 (N_14846,N_11692,N_10827);
nand U14847 (N_14847,N_8400,N_10415);
xnor U14848 (N_14848,N_8571,N_11406);
or U14849 (N_14849,N_11485,N_8662);
or U14850 (N_14850,N_8971,N_11601);
xnor U14851 (N_14851,N_11364,N_11912);
or U14852 (N_14852,N_9331,N_9057);
and U14853 (N_14853,N_10657,N_10346);
and U14854 (N_14854,N_11911,N_10724);
xor U14855 (N_14855,N_8347,N_9113);
and U14856 (N_14856,N_11828,N_9354);
and U14857 (N_14857,N_9520,N_9931);
xnor U14858 (N_14858,N_11934,N_11808);
nand U14859 (N_14859,N_11183,N_10839);
xor U14860 (N_14860,N_10421,N_8649);
nand U14861 (N_14861,N_8897,N_10229);
or U14862 (N_14862,N_8432,N_10100);
nor U14863 (N_14863,N_10155,N_9005);
xnor U14864 (N_14864,N_10366,N_8639);
xor U14865 (N_14865,N_10477,N_10602);
xor U14866 (N_14866,N_9404,N_8158);
nor U14867 (N_14867,N_11530,N_11286);
and U14868 (N_14868,N_8075,N_10505);
or U14869 (N_14869,N_11987,N_10040);
nor U14870 (N_14870,N_10826,N_8807);
or U14871 (N_14871,N_11873,N_10521);
nand U14872 (N_14872,N_9624,N_10640);
nor U14873 (N_14873,N_9598,N_9615);
nor U14874 (N_14874,N_10368,N_8170);
xnor U14875 (N_14875,N_11299,N_10032);
nand U14876 (N_14876,N_10057,N_10518);
nand U14877 (N_14877,N_10345,N_9242);
nor U14878 (N_14878,N_9116,N_8209);
nand U14879 (N_14879,N_10091,N_11391);
xnor U14880 (N_14880,N_10600,N_8769);
and U14881 (N_14881,N_9781,N_9337);
nor U14882 (N_14882,N_8271,N_9043);
nor U14883 (N_14883,N_11990,N_11029);
nand U14884 (N_14884,N_8890,N_8779);
or U14885 (N_14885,N_11669,N_10050);
and U14886 (N_14886,N_11359,N_11969);
and U14887 (N_14887,N_9470,N_10934);
and U14888 (N_14888,N_11138,N_10206);
and U14889 (N_14889,N_11442,N_8175);
or U14890 (N_14890,N_8862,N_10174);
nor U14891 (N_14891,N_9080,N_8581);
nand U14892 (N_14892,N_8812,N_10518);
nand U14893 (N_14893,N_8413,N_10863);
nand U14894 (N_14894,N_9619,N_10750);
nand U14895 (N_14895,N_11123,N_8023);
or U14896 (N_14896,N_9784,N_9975);
xnor U14897 (N_14897,N_10146,N_8508);
and U14898 (N_14898,N_10734,N_8812);
and U14899 (N_14899,N_11485,N_8809);
xor U14900 (N_14900,N_9009,N_10925);
nor U14901 (N_14901,N_10725,N_8374);
xor U14902 (N_14902,N_11233,N_9905);
and U14903 (N_14903,N_8398,N_11914);
nor U14904 (N_14904,N_8256,N_11775);
nand U14905 (N_14905,N_10343,N_9919);
xnor U14906 (N_14906,N_9950,N_11280);
xnor U14907 (N_14907,N_11445,N_8242);
or U14908 (N_14908,N_10005,N_9783);
nand U14909 (N_14909,N_8034,N_10215);
or U14910 (N_14910,N_11424,N_9167);
and U14911 (N_14911,N_11696,N_8201);
and U14912 (N_14912,N_8244,N_11433);
or U14913 (N_14913,N_9484,N_8150);
or U14914 (N_14914,N_9681,N_11327);
and U14915 (N_14915,N_11007,N_8210);
and U14916 (N_14916,N_11713,N_11779);
xnor U14917 (N_14917,N_10613,N_10955);
and U14918 (N_14918,N_11243,N_10289);
and U14919 (N_14919,N_11806,N_10212);
nand U14920 (N_14920,N_9301,N_8282);
nand U14921 (N_14921,N_11196,N_9845);
or U14922 (N_14922,N_8515,N_10132);
nor U14923 (N_14923,N_8279,N_11950);
nor U14924 (N_14924,N_10681,N_8333);
and U14925 (N_14925,N_8946,N_9307);
or U14926 (N_14926,N_9093,N_11997);
and U14927 (N_14927,N_9064,N_10617);
xor U14928 (N_14928,N_11325,N_9847);
xnor U14929 (N_14929,N_9311,N_11890);
nand U14930 (N_14930,N_10008,N_8390);
or U14931 (N_14931,N_8129,N_10733);
xnor U14932 (N_14932,N_8036,N_11401);
and U14933 (N_14933,N_8959,N_11968);
xor U14934 (N_14934,N_10863,N_10062);
xnor U14935 (N_14935,N_8671,N_9359);
nand U14936 (N_14936,N_11013,N_9967);
xor U14937 (N_14937,N_10586,N_9536);
nor U14938 (N_14938,N_9073,N_10437);
nand U14939 (N_14939,N_11409,N_9406);
nand U14940 (N_14940,N_10498,N_8355);
xnor U14941 (N_14941,N_11764,N_9344);
and U14942 (N_14942,N_8719,N_10177);
nand U14943 (N_14943,N_9139,N_9942);
nor U14944 (N_14944,N_9270,N_10117);
nand U14945 (N_14945,N_11900,N_9899);
nor U14946 (N_14946,N_11679,N_11297);
nand U14947 (N_14947,N_9209,N_8701);
nor U14948 (N_14948,N_11040,N_10679);
nand U14949 (N_14949,N_10932,N_11764);
or U14950 (N_14950,N_9257,N_10680);
or U14951 (N_14951,N_11520,N_11346);
and U14952 (N_14952,N_9950,N_8337);
xnor U14953 (N_14953,N_9484,N_9451);
xnor U14954 (N_14954,N_11304,N_11011);
or U14955 (N_14955,N_9357,N_9704);
nand U14956 (N_14956,N_9246,N_11584);
nand U14957 (N_14957,N_9677,N_10930);
and U14958 (N_14958,N_10953,N_11851);
nor U14959 (N_14959,N_9382,N_11989);
or U14960 (N_14960,N_10990,N_9047);
or U14961 (N_14961,N_9497,N_8678);
nor U14962 (N_14962,N_11681,N_8106);
and U14963 (N_14963,N_11630,N_9824);
nor U14964 (N_14964,N_8273,N_10358);
and U14965 (N_14965,N_8148,N_8218);
and U14966 (N_14966,N_10674,N_11938);
and U14967 (N_14967,N_9753,N_11295);
xnor U14968 (N_14968,N_11639,N_8461);
and U14969 (N_14969,N_10598,N_9640);
nor U14970 (N_14970,N_10635,N_9332);
xnor U14971 (N_14971,N_8644,N_11416);
xor U14972 (N_14972,N_11073,N_10670);
nor U14973 (N_14973,N_10960,N_8226);
xnor U14974 (N_14974,N_11744,N_10467);
and U14975 (N_14975,N_11434,N_11009);
and U14976 (N_14976,N_11865,N_9473);
and U14977 (N_14977,N_10651,N_8116);
xor U14978 (N_14978,N_11828,N_11076);
and U14979 (N_14979,N_8942,N_11659);
and U14980 (N_14980,N_9307,N_9453);
nor U14981 (N_14981,N_11217,N_8174);
nand U14982 (N_14982,N_8746,N_10014);
or U14983 (N_14983,N_9690,N_8571);
nor U14984 (N_14984,N_8290,N_8969);
and U14985 (N_14985,N_8194,N_8104);
xor U14986 (N_14986,N_9152,N_10483);
nand U14987 (N_14987,N_10070,N_11370);
or U14988 (N_14988,N_10132,N_8754);
and U14989 (N_14989,N_9880,N_8331);
and U14990 (N_14990,N_9185,N_9205);
or U14991 (N_14991,N_9441,N_10659);
nor U14992 (N_14992,N_10739,N_8443);
nor U14993 (N_14993,N_8915,N_8419);
nand U14994 (N_14994,N_11102,N_10799);
or U14995 (N_14995,N_9248,N_10109);
xor U14996 (N_14996,N_8715,N_8968);
xor U14997 (N_14997,N_9778,N_11365);
or U14998 (N_14998,N_10492,N_10923);
and U14999 (N_14999,N_10684,N_11021);
and U15000 (N_15000,N_10769,N_9266);
nand U15001 (N_15001,N_11249,N_10469);
nor U15002 (N_15002,N_10254,N_8517);
and U15003 (N_15003,N_9055,N_8393);
or U15004 (N_15004,N_9153,N_11440);
nor U15005 (N_15005,N_10818,N_10898);
or U15006 (N_15006,N_9536,N_11648);
nand U15007 (N_15007,N_8653,N_10718);
or U15008 (N_15008,N_10112,N_11722);
xnor U15009 (N_15009,N_11030,N_8762);
nand U15010 (N_15010,N_10698,N_10871);
or U15011 (N_15011,N_9535,N_11954);
or U15012 (N_15012,N_8218,N_10975);
and U15013 (N_15013,N_8109,N_11249);
xnor U15014 (N_15014,N_11678,N_9807);
xnor U15015 (N_15015,N_10057,N_10797);
xor U15016 (N_15016,N_11415,N_8836);
or U15017 (N_15017,N_10273,N_11041);
and U15018 (N_15018,N_9093,N_9147);
nor U15019 (N_15019,N_11979,N_10274);
nand U15020 (N_15020,N_9188,N_11901);
xnor U15021 (N_15021,N_10382,N_9935);
nand U15022 (N_15022,N_10059,N_8567);
nor U15023 (N_15023,N_9661,N_9095);
nand U15024 (N_15024,N_9651,N_9022);
or U15025 (N_15025,N_8304,N_8362);
nand U15026 (N_15026,N_9339,N_8894);
and U15027 (N_15027,N_10121,N_9752);
xor U15028 (N_15028,N_8101,N_8303);
nand U15029 (N_15029,N_9701,N_9473);
and U15030 (N_15030,N_10614,N_10174);
nand U15031 (N_15031,N_9472,N_8468);
nor U15032 (N_15032,N_9927,N_9074);
or U15033 (N_15033,N_8700,N_8383);
nand U15034 (N_15034,N_10869,N_10301);
or U15035 (N_15035,N_10929,N_8459);
nor U15036 (N_15036,N_8863,N_11681);
xor U15037 (N_15037,N_8976,N_9198);
xnor U15038 (N_15038,N_8632,N_10052);
and U15039 (N_15039,N_10143,N_9474);
xnor U15040 (N_15040,N_9878,N_9432);
or U15041 (N_15041,N_9534,N_10801);
and U15042 (N_15042,N_10919,N_10933);
nor U15043 (N_15043,N_9123,N_9416);
nand U15044 (N_15044,N_8992,N_10928);
nand U15045 (N_15045,N_9010,N_9765);
or U15046 (N_15046,N_8118,N_8537);
and U15047 (N_15047,N_9987,N_9783);
or U15048 (N_15048,N_10066,N_10124);
nand U15049 (N_15049,N_8052,N_8022);
and U15050 (N_15050,N_11045,N_10083);
nand U15051 (N_15051,N_11272,N_8490);
and U15052 (N_15052,N_9340,N_8513);
and U15053 (N_15053,N_11844,N_8837);
nand U15054 (N_15054,N_9599,N_8366);
nand U15055 (N_15055,N_9584,N_11038);
nand U15056 (N_15056,N_11479,N_9154);
or U15057 (N_15057,N_9499,N_9739);
nor U15058 (N_15058,N_10460,N_9934);
or U15059 (N_15059,N_11035,N_9297);
xor U15060 (N_15060,N_9868,N_11204);
nor U15061 (N_15061,N_8957,N_10020);
or U15062 (N_15062,N_11142,N_10920);
nor U15063 (N_15063,N_10643,N_9483);
and U15064 (N_15064,N_9489,N_10270);
nor U15065 (N_15065,N_11227,N_9871);
and U15066 (N_15066,N_10572,N_8749);
and U15067 (N_15067,N_8158,N_8122);
nor U15068 (N_15068,N_8920,N_11283);
and U15069 (N_15069,N_8835,N_9009);
and U15070 (N_15070,N_10788,N_10998);
nand U15071 (N_15071,N_10642,N_11235);
or U15072 (N_15072,N_8470,N_9369);
nand U15073 (N_15073,N_8702,N_10689);
and U15074 (N_15074,N_9355,N_10703);
nor U15075 (N_15075,N_9445,N_9597);
xor U15076 (N_15076,N_10629,N_9584);
or U15077 (N_15077,N_10800,N_10591);
or U15078 (N_15078,N_8894,N_9317);
or U15079 (N_15079,N_11598,N_11042);
nor U15080 (N_15080,N_11208,N_10346);
nand U15081 (N_15081,N_10185,N_8746);
xnor U15082 (N_15082,N_10150,N_11521);
xnor U15083 (N_15083,N_10762,N_9645);
or U15084 (N_15084,N_8593,N_9613);
xnor U15085 (N_15085,N_11102,N_8110);
nand U15086 (N_15086,N_10555,N_11579);
nand U15087 (N_15087,N_11355,N_11985);
or U15088 (N_15088,N_10107,N_8970);
nand U15089 (N_15089,N_9948,N_10948);
xor U15090 (N_15090,N_10373,N_8330);
xor U15091 (N_15091,N_8082,N_11346);
xor U15092 (N_15092,N_10867,N_11159);
and U15093 (N_15093,N_8197,N_11874);
nor U15094 (N_15094,N_10112,N_9571);
and U15095 (N_15095,N_8806,N_8431);
nor U15096 (N_15096,N_11809,N_9870);
xnor U15097 (N_15097,N_11737,N_11895);
nor U15098 (N_15098,N_8962,N_9706);
xnor U15099 (N_15099,N_9782,N_11993);
nand U15100 (N_15100,N_10713,N_10650);
nor U15101 (N_15101,N_8631,N_8871);
nand U15102 (N_15102,N_11242,N_11125);
nand U15103 (N_15103,N_9180,N_8119);
or U15104 (N_15104,N_9379,N_8777);
or U15105 (N_15105,N_10298,N_10362);
nor U15106 (N_15106,N_8463,N_9838);
nand U15107 (N_15107,N_10477,N_9361);
or U15108 (N_15108,N_11567,N_10010);
and U15109 (N_15109,N_8612,N_8597);
or U15110 (N_15110,N_11219,N_9650);
or U15111 (N_15111,N_9068,N_11394);
or U15112 (N_15112,N_10052,N_8682);
and U15113 (N_15113,N_11809,N_10012);
nand U15114 (N_15114,N_11270,N_11848);
nand U15115 (N_15115,N_8228,N_9904);
nor U15116 (N_15116,N_11194,N_11570);
or U15117 (N_15117,N_10502,N_8288);
nand U15118 (N_15118,N_10139,N_11807);
or U15119 (N_15119,N_11300,N_9350);
and U15120 (N_15120,N_11062,N_11411);
nor U15121 (N_15121,N_8641,N_10878);
nand U15122 (N_15122,N_10676,N_9543);
nand U15123 (N_15123,N_10675,N_11296);
and U15124 (N_15124,N_10642,N_8801);
and U15125 (N_15125,N_8212,N_11408);
and U15126 (N_15126,N_10522,N_11824);
and U15127 (N_15127,N_8875,N_11367);
nand U15128 (N_15128,N_11686,N_10011);
nor U15129 (N_15129,N_8969,N_10155);
or U15130 (N_15130,N_10950,N_8811);
or U15131 (N_15131,N_11785,N_11930);
xnor U15132 (N_15132,N_8361,N_11663);
nor U15133 (N_15133,N_9386,N_9452);
xor U15134 (N_15134,N_10492,N_11971);
or U15135 (N_15135,N_8939,N_8185);
nor U15136 (N_15136,N_9044,N_8557);
nand U15137 (N_15137,N_11247,N_10377);
and U15138 (N_15138,N_10704,N_10868);
or U15139 (N_15139,N_9422,N_11756);
or U15140 (N_15140,N_9947,N_9178);
and U15141 (N_15141,N_9509,N_11874);
nor U15142 (N_15142,N_10347,N_10957);
and U15143 (N_15143,N_9470,N_11420);
nand U15144 (N_15144,N_8772,N_10027);
or U15145 (N_15145,N_11077,N_10514);
nor U15146 (N_15146,N_10973,N_9369);
or U15147 (N_15147,N_9757,N_11120);
nand U15148 (N_15148,N_9838,N_10163);
nand U15149 (N_15149,N_9106,N_9818);
nor U15150 (N_15150,N_9235,N_9419);
and U15151 (N_15151,N_10733,N_11325);
or U15152 (N_15152,N_10672,N_10485);
or U15153 (N_15153,N_11339,N_8418);
nand U15154 (N_15154,N_9563,N_10282);
nor U15155 (N_15155,N_10462,N_10313);
xor U15156 (N_15156,N_11704,N_9380);
xnor U15157 (N_15157,N_8363,N_11041);
nand U15158 (N_15158,N_11731,N_9143);
nand U15159 (N_15159,N_8048,N_9009);
or U15160 (N_15160,N_8265,N_8193);
or U15161 (N_15161,N_9267,N_11718);
nor U15162 (N_15162,N_8241,N_8634);
nand U15163 (N_15163,N_9379,N_10141);
nor U15164 (N_15164,N_11469,N_9939);
or U15165 (N_15165,N_8343,N_11340);
xor U15166 (N_15166,N_11725,N_11586);
or U15167 (N_15167,N_8977,N_10176);
nor U15168 (N_15168,N_10395,N_11715);
xnor U15169 (N_15169,N_11137,N_10180);
xor U15170 (N_15170,N_10533,N_11055);
nor U15171 (N_15171,N_11222,N_11371);
nor U15172 (N_15172,N_8827,N_11101);
xor U15173 (N_15173,N_10956,N_9466);
or U15174 (N_15174,N_9728,N_10933);
nand U15175 (N_15175,N_10058,N_9774);
and U15176 (N_15176,N_8919,N_10003);
or U15177 (N_15177,N_8427,N_11787);
and U15178 (N_15178,N_8471,N_11136);
nand U15179 (N_15179,N_9609,N_11652);
nor U15180 (N_15180,N_8831,N_8417);
nor U15181 (N_15181,N_10772,N_9357);
nor U15182 (N_15182,N_9079,N_10986);
and U15183 (N_15183,N_8828,N_10769);
or U15184 (N_15184,N_8200,N_11097);
xnor U15185 (N_15185,N_9046,N_11491);
xnor U15186 (N_15186,N_9776,N_9068);
or U15187 (N_15187,N_10327,N_9818);
xor U15188 (N_15188,N_8324,N_9436);
nor U15189 (N_15189,N_10722,N_11828);
or U15190 (N_15190,N_9449,N_8973);
or U15191 (N_15191,N_9703,N_8812);
nor U15192 (N_15192,N_8055,N_8439);
nor U15193 (N_15193,N_10377,N_11020);
or U15194 (N_15194,N_11460,N_9045);
nand U15195 (N_15195,N_10031,N_9609);
nand U15196 (N_15196,N_8761,N_8813);
or U15197 (N_15197,N_10493,N_11016);
xnor U15198 (N_15198,N_9657,N_9165);
xnor U15199 (N_15199,N_11228,N_11880);
nand U15200 (N_15200,N_9534,N_9331);
or U15201 (N_15201,N_10361,N_8547);
nor U15202 (N_15202,N_11525,N_8077);
xnor U15203 (N_15203,N_8290,N_8087);
nor U15204 (N_15204,N_8990,N_9673);
or U15205 (N_15205,N_9746,N_11782);
and U15206 (N_15206,N_10241,N_8946);
xor U15207 (N_15207,N_11872,N_8326);
nor U15208 (N_15208,N_10867,N_10695);
xor U15209 (N_15209,N_10400,N_8168);
and U15210 (N_15210,N_11969,N_8173);
nor U15211 (N_15211,N_8888,N_10239);
or U15212 (N_15212,N_11825,N_10336);
nor U15213 (N_15213,N_8396,N_8102);
and U15214 (N_15214,N_11429,N_8345);
or U15215 (N_15215,N_11279,N_9333);
and U15216 (N_15216,N_9112,N_8518);
and U15217 (N_15217,N_8689,N_9617);
xnor U15218 (N_15218,N_9387,N_10175);
nand U15219 (N_15219,N_8564,N_9434);
and U15220 (N_15220,N_8635,N_9658);
or U15221 (N_15221,N_11342,N_10629);
nor U15222 (N_15222,N_9699,N_10727);
xnor U15223 (N_15223,N_10541,N_8476);
and U15224 (N_15224,N_8680,N_11607);
nor U15225 (N_15225,N_10822,N_9679);
and U15226 (N_15226,N_11711,N_11479);
nand U15227 (N_15227,N_8558,N_11825);
or U15228 (N_15228,N_9094,N_8730);
and U15229 (N_15229,N_8585,N_8249);
xnor U15230 (N_15230,N_11149,N_8510);
nor U15231 (N_15231,N_8792,N_11929);
nand U15232 (N_15232,N_8042,N_10024);
and U15233 (N_15233,N_8981,N_11018);
xnor U15234 (N_15234,N_9346,N_11812);
nand U15235 (N_15235,N_8189,N_11199);
or U15236 (N_15236,N_9519,N_11565);
nor U15237 (N_15237,N_9981,N_9976);
xor U15238 (N_15238,N_9070,N_10779);
xnor U15239 (N_15239,N_10399,N_8912);
xor U15240 (N_15240,N_10837,N_8928);
or U15241 (N_15241,N_11976,N_11936);
or U15242 (N_15242,N_10475,N_8691);
nor U15243 (N_15243,N_9921,N_11589);
nor U15244 (N_15244,N_9929,N_10846);
nand U15245 (N_15245,N_9070,N_8668);
and U15246 (N_15246,N_9386,N_8257);
nand U15247 (N_15247,N_11113,N_9253);
xor U15248 (N_15248,N_8737,N_9481);
nor U15249 (N_15249,N_8687,N_9620);
nor U15250 (N_15250,N_8884,N_9934);
xor U15251 (N_15251,N_8924,N_10518);
nor U15252 (N_15252,N_11451,N_10638);
nor U15253 (N_15253,N_10680,N_9898);
and U15254 (N_15254,N_8689,N_9876);
nor U15255 (N_15255,N_8840,N_10936);
nand U15256 (N_15256,N_11739,N_8460);
nor U15257 (N_15257,N_8766,N_11711);
and U15258 (N_15258,N_10860,N_9099);
xor U15259 (N_15259,N_11928,N_11391);
or U15260 (N_15260,N_10153,N_10233);
nand U15261 (N_15261,N_9856,N_11824);
nand U15262 (N_15262,N_10593,N_9065);
xor U15263 (N_15263,N_10285,N_11117);
or U15264 (N_15264,N_9979,N_10165);
nand U15265 (N_15265,N_10443,N_9018);
nand U15266 (N_15266,N_8094,N_8916);
or U15267 (N_15267,N_10921,N_10514);
and U15268 (N_15268,N_9908,N_9160);
and U15269 (N_15269,N_8480,N_11265);
and U15270 (N_15270,N_11356,N_11810);
and U15271 (N_15271,N_8197,N_10424);
nand U15272 (N_15272,N_11912,N_9228);
xor U15273 (N_15273,N_11680,N_8849);
nor U15274 (N_15274,N_9842,N_8699);
nand U15275 (N_15275,N_9746,N_8157);
or U15276 (N_15276,N_11824,N_11973);
nand U15277 (N_15277,N_11611,N_10491);
xor U15278 (N_15278,N_9405,N_8623);
nor U15279 (N_15279,N_9371,N_11219);
nor U15280 (N_15280,N_10388,N_11605);
or U15281 (N_15281,N_11911,N_10735);
nand U15282 (N_15282,N_9652,N_11101);
or U15283 (N_15283,N_8242,N_8926);
nand U15284 (N_15284,N_10055,N_10520);
nor U15285 (N_15285,N_11171,N_8529);
xnor U15286 (N_15286,N_10083,N_8369);
nor U15287 (N_15287,N_8686,N_10360);
or U15288 (N_15288,N_8690,N_9950);
xor U15289 (N_15289,N_9560,N_10537);
nand U15290 (N_15290,N_11521,N_11438);
xnor U15291 (N_15291,N_11310,N_8402);
xnor U15292 (N_15292,N_9289,N_11071);
and U15293 (N_15293,N_9230,N_11691);
xor U15294 (N_15294,N_8415,N_9103);
nor U15295 (N_15295,N_8103,N_10544);
nor U15296 (N_15296,N_11061,N_9797);
xnor U15297 (N_15297,N_9123,N_10783);
nor U15298 (N_15298,N_10142,N_8721);
and U15299 (N_15299,N_10556,N_9305);
xor U15300 (N_15300,N_11115,N_11433);
or U15301 (N_15301,N_10389,N_9997);
nor U15302 (N_15302,N_10459,N_10195);
or U15303 (N_15303,N_8043,N_11260);
xnor U15304 (N_15304,N_10809,N_10897);
xor U15305 (N_15305,N_11989,N_9144);
nor U15306 (N_15306,N_8289,N_8059);
nor U15307 (N_15307,N_11923,N_8088);
nor U15308 (N_15308,N_10399,N_8726);
and U15309 (N_15309,N_10075,N_11404);
and U15310 (N_15310,N_9535,N_9013);
nor U15311 (N_15311,N_8984,N_8874);
or U15312 (N_15312,N_10552,N_8220);
xor U15313 (N_15313,N_9112,N_9128);
nand U15314 (N_15314,N_8590,N_11002);
nor U15315 (N_15315,N_9259,N_8132);
xnor U15316 (N_15316,N_11335,N_10732);
or U15317 (N_15317,N_10087,N_9887);
nor U15318 (N_15318,N_9724,N_11779);
or U15319 (N_15319,N_10835,N_9726);
and U15320 (N_15320,N_9723,N_10728);
or U15321 (N_15321,N_8013,N_11986);
and U15322 (N_15322,N_10445,N_10242);
and U15323 (N_15323,N_10826,N_9188);
nor U15324 (N_15324,N_8611,N_8920);
nor U15325 (N_15325,N_10836,N_9787);
nand U15326 (N_15326,N_9910,N_8101);
nor U15327 (N_15327,N_10800,N_9376);
xor U15328 (N_15328,N_8202,N_9981);
xnor U15329 (N_15329,N_10594,N_9053);
nor U15330 (N_15330,N_11007,N_11714);
nand U15331 (N_15331,N_11008,N_8125);
nor U15332 (N_15332,N_9220,N_9955);
or U15333 (N_15333,N_8756,N_10106);
nand U15334 (N_15334,N_10667,N_10079);
nand U15335 (N_15335,N_9658,N_11767);
xor U15336 (N_15336,N_8283,N_10582);
and U15337 (N_15337,N_10257,N_10555);
or U15338 (N_15338,N_8558,N_9849);
nor U15339 (N_15339,N_8534,N_8450);
nand U15340 (N_15340,N_11849,N_8813);
and U15341 (N_15341,N_10959,N_11447);
nor U15342 (N_15342,N_10330,N_10825);
or U15343 (N_15343,N_9439,N_8836);
nor U15344 (N_15344,N_9280,N_8692);
nand U15345 (N_15345,N_10109,N_10467);
nor U15346 (N_15346,N_10201,N_9465);
xnor U15347 (N_15347,N_10753,N_10795);
nand U15348 (N_15348,N_11433,N_8115);
or U15349 (N_15349,N_9468,N_9937);
or U15350 (N_15350,N_8273,N_10618);
nand U15351 (N_15351,N_9665,N_9688);
xor U15352 (N_15352,N_9923,N_10801);
and U15353 (N_15353,N_9175,N_8254);
and U15354 (N_15354,N_11994,N_9193);
nor U15355 (N_15355,N_11585,N_9424);
or U15356 (N_15356,N_11805,N_9049);
and U15357 (N_15357,N_9223,N_9266);
and U15358 (N_15358,N_10620,N_8899);
or U15359 (N_15359,N_10605,N_10394);
xor U15360 (N_15360,N_8850,N_10665);
or U15361 (N_15361,N_9804,N_9991);
and U15362 (N_15362,N_9411,N_8199);
nand U15363 (N_15363,N_8038,N_11592);
xor U15364 (N_15364,N_8511,N_9818);
nand U15365 (N_15365,N_11164,N_10022);
nor U15366 (N_15366,N_8297,N_8512);
xnor U15367 (N_15367,N_10845,N_10726);
nor U15368 (N_15368,N_9605,N_10671);
nand U15369 (N_15369,N_8195,N_8068);
and U15370 (N_15370,N_9590,N_11431);
nor U15371 (N_15371,N_8337,N_10122);
nor U15372 (N_15372,N_8439,N_8634);
nand U15373 (N_15373,N_8914,N_9889);
nor U15374 (N_15374,N_10536,N_11548);
nand U15375 (N_15375,N_10594,N_11849);
nand U15376 (N_15376,N_10758,N_11285);
nor U15377 (N_15377,N_9946,N_8775);
nor U15378 (N_15378,N_10390,N_10345);
and U15379 (N_15379,N_11849,N_8418);
xor U15380 (N_15380,N_9333,N_10257);
xor U15381 (N_15381,N_9188,N_8749);
nand U15382 (N_15382,N_10621,N_9630);
nor U15383 (N_15383,N_11441,N_8317);
xor U15384 (N_15384,N_10111,N_8132);
or U15385 (N_15385,N_9340,N_11311);
nor U15386 (N_15386,N_8929,N_11372);
nand U15387 (N_15387,N_9997,N_8488);
or U15388 (N_15388,N_11362,N_11774);
nand U15389 (N_15389,N_11227,N_9329);
and U15390 (N_15390,N_11133,N_11411);
nand U15391 (N_15391,N_10488,N_10065);
nand U15392 (N_15392,N_10913,N_10419);
nand U15393 (N_15393,N_8832,N_10056);
xor U15394 (N_15394,N_10107,N_8012);
and U15395 (N_15395,N_8742,N_11314);
xnor U15396 (N_15396,N_11151,N_8672);
nor U15397 (N_15397,N_9836,N_9565);
nand U15398 (N_15398,N_10212,N_11706);
nand U15399 (N_15399,N_9728,N_10122);
nand U15400 (N_15400,N_9931,N_10487);
and U15401 (N_15401,N_8305,N_11333);
and U15402 (N_15402,N_8890,N_8612);
and U15403 (N_15403,N_9399,N_8852);
and U15404 (N_15404,N_9868,N_9199);
nand U15405 (N_15405,N_10895,N_11634);
nand U15406 (N_15406,N_11714,N_9214);
nor U15407 (N_15407,N_9704,N_9561);
xor U15408 (N_15408,N_11420,N_9240);
xor U15409 (N_15409,N_10043,N_10636);
nand U15410 (N_15410,N_10307,N_8041);
and U15411 (N_15411,N_8347,N_11112);
nand U15412 (N_15412,N_9596,N_8242);
nand U15413 (N_15413,N_8945,N_11411);
or U15414 (N_15414,N_11601,N_10853);
or U15415 (N_15415,N_9469,N_10257);
nor U15416 (N_15416,N_8525,N_11136);
xor U15417 (N_15417,N_10682,N_9239);
nand U15418 (N_15418,N_11618,N_11338);
nor U15419 (N_15419,N_8918,N_9396);
nor U15420 (N_15420,N_11203,N_11184);
nor U15421 (N_15421,N_8000,N_9767);
or U15422 (N_15422,N_11949,N_9029);
or U15423 (N_15423,N_11846,N_11995);
and U15424 (N_15424,N_9908,N_11084);
nand U15425 (N_15425,N_9275,N_10348);
or U15426 (N_15426,N_9038,N_8256);
and U15427 (N_15427,N_11577,N_11526);
nand U15428 (N_15428,N_10629,N_10282);
xor U15429 (N_15429,N_10451,N_10209);
xor U15430 (N_15430,N_10655,N_10754);
or U15431 (N_15431,N_11954,N_8322);
nand U15432 (N_15432,N_10477,N_10841);
nand U15433 (N_15433,N_10481,N_8549);
or U15434 (N_15434,N_11667,N_8283);
nand U15435 (N_15435,N_11280,N_8014);
and U15436 (N_15436,N_11210,N_9072);
or U15437 (N_15437,N_8537,N_11143);
nand U15438 (N_15438,N_8017,N_11290);
nor U15439 (N_15439,N_11249,N_11203);
and U15440 (N_15440,N_11787,N_11742);
nand U15441 (N_15441,N_8977,N_8536);
and U15442 (N_15442,N_11437,N_10174);
or U15443 (N_15443,N_8240,N_11783);
or U15444 (N_15444,N_11279,N_10547);
nor U15445 (N_15445,N_8664,N_8090);
nand U15446 (N_15446,N_10077,N_10034);
or U15447 (N_15447,N_8020,N_11371);
nand U15448 (N_15448,N_10840,N_9133);
or U15449 (N_15449,N_10525,N_10629);
nand U15450 (N_15450,N_11396,N_11374);
or U15451 (N_15451,N_10295,N_11269);
xnor U15452 (N_15452,N_9300,N_8777);
and U15453 (N_15453,N_11816,N_8447);
or U15454 (N_15454,N_8247,N_8796);
nor U15455 (N_15455,N_11853,N_9522);
and U15456 (N_15456,N_8513,N_10299);
nand U15457 (N_15457,N_9461,N_11409);
and U15458 (N_15458,N_11436,N_11274);
and U15459 (N_15459,N_11606,N_10739);
or U15460 (N_15460,N_10453,N_11737);
nand U15461 (N_15461,N_9386,N_9123);
xnor U15462 (N_15462,N_11865,N_10185);
nand U15463 (N_15463,N_9784,N_10803);
and U15464 (N_15464,N_9379,N_8437);
and U15465 (N_15465,N_10440,N_10428);
or U15466 (N_15466,N_10381,N_11344);
xnor U15467 (N_15467,N_8000,N_10959);
and U15468 (N_15468,N_9681,N_8164);
and U15469 (N_15469,N_10005,N_10534);
nand U15470 (N_15470,N_9563,N_10538);
nor U15471 (N_15471,N_11988,N_9275);
xor U15472 (N_15472,N_11668,N_11316);
nand U15473 (N_15473,N_9660,N_8900);
and U15474 (N_15474,N_9937,N_11036);
xor U15475 (N_15475,N_10750,N_10621);
xor U15476 (N_15476,N_8373,N_9595);
xor U15477 (N_15477,N_10655,N_9525);
and U15478 (N_15478,N_10540,N_11894);
nand U15479 (N_15479,N_8807,N_9670);
or U15480 (N_15480,N_11499,N_8356);
nand U15481 (N_15481,N_11238,N_10176);
or U15482 (N_15482,N_10585,N_11424);
nand U15483 (N_15483,N_9709,N_8443);
xor U15484 (N_15484,N_8448,N_11590);
and U15485 (N_15485,N_8327,N_9421);
nor U15486 (N_15486,N_11459,N_11548);
and U15487 (N_15487,N_11352,N_9271);
nand U15488 (N_15488,N_9242,N_8260);
nor U15489 (N_15489,N_10119,N_10586);
nor U15490 (N_15490,N_8021,N_8674);
and U15491 (N_15491,N_9928,N_8935);
nand U15492 (N_15492,N_11265,N_10254);
nor U15493 (N_15493,N_10972,N_9498);
or U15494 (N_15494,N_11658,N_9953);
nand U15495 (N_15495,N_9916,N_8460);
nor U15496 (N_15496,N_9989,N_10097);
xnor U15497 (N_15497,N_9563,N_10902);
or U15498 (N_15498,N_11840,N_10163);
nand U15499 (N_15499,N_8604,N_11836);
xnor U15500 (N_15500,N_9761,N_10058);
nor U15501 (N_15501,N_10517,N_9557);
nand U15502 (N_15502,N_11404,N_11146);
xor U15503 (N_15503,N_11966,N_8595);
xnor U15504 (N_15504,N_8490,N_8382);
nor U15505 (N_15505,N_11835,N_8177);
xor U15506 (N_15506,N_9336,N_8058);
or U15507 (N_15507,N_10788,N_8106);
xnor U15508 (N_15508,N_8956,N_8608);
and U15509 (N_15509,N_11257,N_9192);
nand U15510 (N_15510,N_11572,N_10978);
or U15511 (N_15511,N_9304,N_9625);
nor U15512 (N_15512,N_9030,N_8692);
nand U15513 (N_15513,N_10541,N_11647);
and U15514 (N_15514,N_9334,N_10210);
or U15515 (N_15515,N_9801,N_9910);
and U15516 (N_15516,N_9130,N_10508);
nor U15517 (N_15517,N_8449,N_10400);
nand U15518 (N_15518,N_10398,N_8109);
nor U15519 (N_15519,N_8428,N_11918);
nor U15520 (N_15520,N_9966,N_8041);
or U15521 (N_15521,N_11215,N_9757);
and U15522 (N_15522,N_11466,N_8888);
or U15523 (N_15523,N_8159,N_11553);
nand U15524 (N_15524,N_11728,N_11333);
nand U15525 (N_15525,N_8559,N_8623);
nor U15526 (N_15526,N_8957,N_10219);
nand U15527 (N_15527,N_8305,N_11142);
nor U15528 (N_15528,N_9612,N_11780);
xnor U15529 (N_15529,N_11747,N_8847);
nand U15530 (N_15530,N_10126,N_10859);
nand U15531 (N_15531,N_9970,N_8630);
or U15532 (N_15532,N_10476,N_9388);
nand U15533 (N_15533,N_10026,N_9003);
xnor U15534 (N_15534,N_10186,N_8633);
or U15535 (N_15535,N_11768,N_9403);
nand U15536 (N_15536,N_10183,N_9705);
xor U15537 (N_15537,N_10959,N_8548);
xor U15538 (N_15538,N_9188,N_9023);
xor U15539 (N_15539,N_9246,N_8532);
nor U15540 (N_15540,N_8395,N_8026);
nand U15541 (N_15541,N_11603,N_10441);
xnor U15542 (N_15542,N_8273,N_11152);
nand U15543 (N_15543,N_9725,N_8972);
nor U15544 (N_15544,N_11440,N_8763);
nand U15545 (N_15545,N_10157,N_8267);
nand U15546 (N_15546,N_8659,N_9701);
nand U15547 (N_15547,N_8698,N_11587);
nor U15548 (N_15548,N_10530,N_11612);
nor U15549 (N_15549,N_8843,N_10859);
nand U15550 (N_15550,N_11950,N_9326);
and U15551 (N_15551,N_10044,N_9936);
and U15552 (N_15552,N_10691,N_11329);
and U15553 (N_15553,N_8315,N_11972);
xor U15554 (N_15554,N_11477,N_10979);
or U15555 (N_15555,N_9403,N_9193);
nand U15556 (N_15556,N_9540,N_10652);
and U15557 (N_15557,N_8509,N_9388);
xor U15558 (N_15558,N_8830,N_10511);
and U15559 (N_15559,N_8123,N_10680);
nand U15560 (N_15560,N_8906,N_10196);
or U15561 (N_15561,N_8150,N_11916);
nor U15562 (N_15562,N_10004,N_10491);
nand U15563 (N_15563,N_11448,N_8484);
or U15564 (N_15564,N_8659,N_9605);
nand U15565 (N_15565,N_11448,N_10031);
nor U15566 (N_15566,N_8372,N_8712);
nor U15567 (N_15567,N_10790,N_11857);
nor U15568 (N_15568,N_8139,N_10363);
xor U15569 (N_15569,N_10245,N_8915);
xnor U15570 (N_15570,N_9002,N_10131);
nand U15571 (N_15571,N_8142,N_10277);
and U15572 (N_15572,N_11191,N_8046);
or U15573 (N_15573,N_11748,N_8909);
and U15574 (N_15574,N_8222,N_10384);
nand U15575 (N_15575,N_9415,N_9534);
xnor U15576 (N_15576,N_8845,N_10120);
nor U15577 (N_15577,N_11201,N_9160);
nand U15578 (N_15578,N_11800,N_10988);
or U15579 (N_15579,N_9639,N_10478);
xnor U15580 (N_15580,N_9107,N_8464);
xnor U15581 (N_15581,N_8515,N_9969);
xor U15582 (N_15582,N_9130,N_9625);
and U15583 (N_15583,N_10022,N_11099);
nor U15584 (N_15584,N_11216,N_8112);
xnor U15585 (N_15585,N_8297,N_9541);
nor U15586 (N_15586,N_9507,N_8298);
nor U15587 (N_15587,N_9046,N_11869);
nand U15588 (N_15588,N_8539,N_11668);
or U15589 (N_15589,N_8756,N_8999);
nand U15590 (N_15590,N_8855,N_9612);
and U15591 (N_15591,N_8121,N_11033);
nand U15592 (N_15592,N_11833,N_11862);
nand U15593 (N_15593,N_8101,N_9013);
nor U15594 (N_15594,N_8464,N_10643);
and U15595 (N_15595,N_10555,N_9691);
or U15596 (N_15596,N_9202,N_9646);
or U15597 (N_15597,N_11921,N_8913);
nand U15598 (N_15598,N_8055,N_10404);
xnor U15599 (N_15599,N_8075,N_11559);
or U15600 (N_15600,N_11684,N_8786);
nor U15601 (N_15601,N_9395,N_9807);
nor U15602 (N_15602,N_8577,N_8476);
nand U15603 (N_15603,N_9673,N_10785);
nor U15604 (N_15604,N_8274,N_9437);
and U15605 (N_15605,N_8430,N_10392);
and U15606 (N_15606,N_11398,N_11348);
xnor U15607 (N_15607,N_10962,N_8176);
or U15608 (N_15608,N_10892,N_8288);
nor U15609 (N_15609,N_9730,N_9388);
nor U15610 (N_15610,N_11245,N_11730);
and U15611 (N_15611,N_8353,N_11119);
xor U15612 (N_15612,N_9619,N_11357);
nor U15613 (N_15613,N_9166,N_10164);
or U15614 (N_15614,N_11219,N_11997);
nor U15615 (N_15615,N_8067,N_8529);
nor U15616 (N_15616,N_11922,N_9083);
nand U15617 (N_15617,N_11380,N_10744);
nand U15618 (N_15618,N_11276,N_10820);
nor U15619 (N_15619,N_11395,N_8876);
and U15620 (N_15620,N_9311,N_10089);
and U15621 (N_15621,N_8413,N_8782);
nor U15622 (N_15622,N_11967,N_8226);
nor U15623 (N_15623,N_9787,N_8995);
and U15624 (N_15624,N_9065,N_10957);
and U15625 (N_15625,N_10765,N_8994);
xnor U15626 (N_15626,N_11389,N_10568);
nor U15627 (N_15627,N_11413,N_9043);
and U15628 (N_15628,N_10757,N_9018);
and U15629 (N_15629,N_10268,N_11146);
or U15630 (N_15630,N_11036,N_11328);
or U15631 (N_15631,N_10919,N_9621);
xor U15632 (N_15632,N_10580,N_8865);
nor U15633 (N_15633,N_8466,N_9122);
nor U15634 (N_15634,N_9526,N_10889);
xnor U15635 (N_15635,N_8464,N_10461);
nor U15636 (N_15636,N_10830,N_11821);
xor U15637 (N_15637,N_11311,N_8212);
nor U15638 (N_15638,N_11552,N_8160);
or U15639 (N_15639,N_11956,N_10327);
xnor U15640 (N_15640,N_9510,N_11223);
nand U15641 (N_15641,N_9419,N_10383);
or U15642 (N_15642,N_9935,N_10326);
and U15643 (N_15643,N_8276,N_11137);
or U15644 (N_15644,N_8168,N_10495);
nor U15645 (N_15645,N_8569,N_10653);
nand U15646 (N_15646,N_9002,N_9232);
nand U15647 (N_15647,N_11912,N_8068);
and U15648 (N_15648,N_11283,N_10003);
or U15649 (N_15649,N_9844,N_9572);
nand U15650 (N_15650,N_10047,N_8147);
and U15651 (N_15651,N_8080,N_10536);
and U15652 (N_15652,N_9885,N_8061);
and U15653 (N_15653,N_11569,N_9154);
nor U15654 (N_15654,N_10655,N_10686);
or U15655 (N_15655,N_11805,N_8499);
or U15656 (N_15656,N_10396,N_9210);
or U15657 (N_15657,N_9501,N_11836);
or U15658 (N_15658,N_10792,N_11531);
xor U15659 (N_15659,N_11625,N_11789);
xnor U15660 (N_15660,N_10908,N_10598);
nor U15661 (N_15661,N_10229,N_8009);
xnor U15662 (N_15662,N_11119,N_9783);
and U15663 (N_15663,N_11408,N_11566);
xor U15664 (N_15664,N_11087,N_8676);
or U15665 (N_15665,N_8892,N_10864);
xor U15666 (N_15666,N_9001,N_10033);
or U15667 (N_15667,N_10576,N_9294);
or U15668 (N_15668,N_8597,N_11973);
nand U15669 (N_15669,N_11350,N_11462);
and U15670 (N_15670,N_9291,N_10887);
nand U15671 (N_15671,N_11365,N_10390);
or U15672 (N_15672,N_11177,N_9370);
nand U15673 (N_15673,N_9836,N_8839);
xor U15674 (N_15674,N_11480,N_10625);
xor U15675 (N_15675,N_10179,N_8581);
and U15676 (N_15676,N_8862,N_8344);
or U15677 (N_15677,N_9425,N_9076);
xor U15678 (N_15678,N_8626,N_8189);
nand U15679 (N_15679,N_11872,N_8865);
nand U15680 (N_15680,N_9104,N_9793);
nand U15681 (N_15681,N_8741,N_8602);
xor U15682 (N_15682,N_8105,N_11987);
nand U15683 (N_15683,N_10495,N_9012);
or U15684 (N_15684,N_8233,N_10680);
and U15685 (N_15685,N_8074,N_10969);
nor U15686 (N_15686,N_8123,N_11915);
nor U15687 (N_15687,N_10436,N_9603);
or U15688 (N_15688,N_10630,N_9587);
xnor U15689 (N_15689,N_8967,N_11124);
nor U15690 (N_15690,N_10509,N_9476);
and U15691 (N_15691,N_9231,N_8327);
nor U15692 (N_15692,N_9884,N_8027);
nand U15693 (N_15693,N_11807,N_9996);
nand U15694 (N_15694,N_10379,N_10681);
nand U15695 (N_15695,N_10709,N_10752);
or U15696 (N_15696,N_10259,N_8518);
nor U15697 (N_15697,N_10057,N_10190);
nand U15698 (N_15698,N_9432,N_9216);
and U15699 (N_15699,N_9407,N_11326);
nand U15700 (N_15700,N_11984,N_10808);
nand U15701 (N_15701,N_10172,N_9240);
nand U15702 (N_15702,N_10732,N_10534);
xnor U15703 (N_15703,N_10708,N_11916);
or U15704 (N_15704,N_11673,N_11616);
nor U15705 (N_15705,N_9355,N_11856);
xor U15706 (N_15706,N_8298,N_10473);
nand U15707 (N_15707,N_8933,N_11029);
xnor U15708 (N_15708,N_11468,N_11641);
xnor U15709 (N_15709,N_10934,N_9942);
and U15710 (N_15710,N_11679,N_10231);
and U15711 (N_15711,N_9891,N_9182);
nand U15712 (N_15712,N_8074,N_11767);
xor U15713 (N_15713,N_9411,N_10426);
nor U15714 (N_15714,N_8104,N_9282);
nor U15715 (N_15715,N_10837,N_8486);
nand U15716 (N_15716,N_9471,N_9479);
or U15717 (N_15717,N_8805,N_11929);
xnor U15718 (N_15718,N_10701,N_11293);
and U15719 (N_15719,N_10886,N_10650);
xor U15720 (N_15720,N_9362,N_10019);
nor U15721 (N_15721,N_8064,N_10096);
or U15722 (N_15722,N_9253,N_8839);
nand U15723 (N_15723,N_9382,N_10267);
xnor U15724 (N_15724,N_11541,N_11859);
and U15725 (N_15725,N_9230,N_10850);
xnor U15726 (N_15726,N_10965,N_10128);
nand U15727 (N_15727,N_8379,N_10645);
nand U15728 (N_15728,N_9004,N_10868);
xnor U15729 (N_15729,N_8658,N_8041);
nand U15730 (N_15730,N_9492,N_11553);
nand U15731 (N_15731,N_8481,N_8055);
xnor U15732 (N_15732,N_11566,N_11169);
xnor U15733 (N_15733,N_9298,N_10138);
or U15734 (N_15734,N_8705,N_8989);
and U15735 (N_15735,N_8559,N_11993);
or U15736 (N_15736,N_9773,N_9182);
nand U15737 (N_15737,N_8772,N_9417);
nor U15738 (N_15738,N_8428,N_9805);
and U15739 (N_15739,N_10925,N_10468);
nand U15740 (N_15740,N_11776,N_8521);
xor U15741 (N_15741,N_8161,N_8588);
xor U15742 (N_15742,N_11310,N_9928);
nand U15743 (N_15743,N_11709,N_8033);
nand U15744 (N_15744,N_9290,N_9968);
nor U15745 (N_15745,N_9105,N_9631);
nand U15746 (N_15746,N_8555,N_9784);
nor U15747 (N_15747,N_8243,N_8419);
nand U15748 (N_15748,N_11332,N_11374);
nand U15749 (N_15749,N_9026,N_11250);
xor U15750 (N_15750,N_9513,N_10583);
xnor U15751 (N_15751,N_11726,N_11008);
nand U15752 (N_15752,N_9747,N_8885);
or U15753 (N_15753,N_11571,N_11076);
nand U15754 (N_15754,N_9087,N_11860);
nor U15755 (N_15755,N_11084,N_11510);
or U15756 (N_15756,N_10195,N_11979);
or U15757 (N_15757,N_10194,N_9738);
or U15758 (N_15758,N_10439,N_9606);
or U15759 (N_15759,N_10065,N_9246);
xor U15760 (N_15760,N_10622,N_9344);
nand U15761 (N_15761,N_8955,N_8336);
nor U15762 (N_15762,N_10918,N_10618);
nand U15763 (N_15763,N_10259,N_8578);
nor U15764 (N_15764,N_11560,N_10765);
nand U15765 (N_15765,N_10611,N_11253);
nor U15766 (N_15766,N_9461,N_8016);
or U15767 (N_15767,N_11741,N_11270);
or U15768 (N_15768,N_8640,N_9788);
nand U15769 (N_15769,N_10681,N_8970);
or U15770 (N_15770,N_8814,N_8332);
nand U15771 (N_15771,N_8588,N_10922);
or U15772 (N_15772,N_11864,N_9335);
nor U15773 (N_15773,N_11425,N_9596);
nand U15774 (N_15774,N_10541,N_11753);
nor U15775 (N_15775,N_10382,N_9127);
nand U15776 (N_15776,N_9421,N_11375);
nand U15777 (N_15777,N_11230,N_9290);
xor U15778 (N_15778,N_8457,N_9690);
nor U15779 (N_15779,N_9549,N_9642);
or U15780 (N_15780,N_8725,N_8649);
and U15781 (N_15781,N_11283,N_10102);
nor U15782 (N_15782,N_9171,N_8090);
nor U15783 (N_15783,N_11399,N_10277);
nor U15784 (N_15784,N_11172,N_10054);
nand U15785 (N_15785,N_8326,N_11046);
xor U15786 (N_15786,N_9162,N_9968);
or U15787 (N_15787,N_8143,N_8813);
nand U15788 (N_15788,N_8787,N_9178);
or U15789 (N_15789,N_11590,N_9974);
nor U15790 (N_15790,N_8108,N_9649);
nand U15791 (N_15791,N_8522,N_9086);
nor U15792 (N_15792,N_8054,N_10677);
nor U15793 (N_15793,N_8781,N_9173);
nand U15794 (N_15794,N_9506,N_8473);
nor U15795 (N_15795,N_9493,N_9735);
or U15796 (N_15796,N_9875,N_9451);
and U15797 (N_15797,N_9626,N_9688);
nand U15798 (N_15798,N_8844,N_9629);
or U15799 (N_15799,N_10019,N_10398);
and U15800 (N_15800,N_11941,N_10780);
nand U15801 (N_15801,N_10583,N_9539);
nand U15802 (N_15802,N_9795,N_10544);
nor U15803 (N_15803,N_9338,N_9864);
nor U15804 (N_15804,N_9937,N_8010);
or U15805 (N_15805,N_10790,N_9996);
nand U15806 (N_15806,N_11461,N_8249);
and U15807 (N_15807,N_10927,N_10824);
xor U15808 (N_15808,N_8679,N_9338);
nand U15809 (N_15809,N_9977,N_9698);
and U15810 (N_15810,N_9715,N_11000);
and U15811 (N_15811,N_8293,N_10853);
nand U15812 (N_15812,N_11087,N_8447);
and U15813 (N_15813,N_9380,N_11884);
xor U15814 (N_15814,N_8803,N_9839);
nand U15815 (N_15815,N_8494,N_9738);
and U15816 (N_15816,N_10921,N_10244);
or U15817 (N_15817,N_10045,N_9811);
nand U15818 (N_15818,N_11180,N_8150);
nor U15819 (N_15819,N_11670,N_9978);
and U15820 (N_15820,N_10755,N_10261);
nor U15821 (N_15821,N_10378,N_10180);
or U15822 (N_15822,N_9250,N_9261);
or U15823 (N_15823,N_11309,N_8380);
and U15824 (N_15824,N_11113,N_11267);
and U15825 (N_15825,N_9941,N_8789);
nand U15826 (N_15826,N_11216,N_8036);
or U15827 (N_15827,N_9074,N_9442);
nand U15828 (N_15828,N_11750,N_9069);
or U15829 (N_15829,N_11746,N_11411);
or U15830 (N_15830,N_10522,N_11000);
and U15831 (N_15831,N_11187,N_10999);
xnor U15832 (N_15832,N_9029,N_10694);
xor U15833 (N_15833,N_11918,N_8555);
xnor U15834 (N_15834,N_9085,N_9614);
xor U15835 (N_15835,N_11963,N_9683);
xor U15836 (N_15836,N_10585,N_9079);
nand U15837 (N_15837,N_11415,N_9689);
nor U15838 (N_15838,N_8759,N_11029);
xnor U15839 (N_15839,N_8790,N_11468);
nor U15840 (N_15840,N_10940,N_8825);
nand U15841 (N_15841,N_11298,N_9983);
nand U15842 (N_15842,N_8266,N_11141);
or U15843 (N_15843,N_11721,N_10931);
or U15844 (N_15844,N_11297,N_11085);
nor U15845 (N_15845,N_9392,N_10989);
nor U15846 (N_15846,N_10527,N_8495);
and U15847 (N_15847,N_8818,N_8211);
or U15848 (N_15848,N_11574,N_11887);
nand U15849 (N_15849,N_10518,N_10517);
and U15850 (N_15850,N_11822,N_8702);
xnor U15851 (N_15851,N_11381,N_10323);
xor U15852 (N_15852,N_10973,N_8323);
nand U15853 (N_15853,N_9443,N_10316);
and U15854 (N_15854,N_9785,N_11005);
nand U15855 (N_15855,N_9439,N_9679);
or U15856 (N_15856,N_10328,N_8085);
xor U15857 (N_15857,N_9422,N_9840);
nand U15858 (N_15858,N_9066,N_10105);
or U15859 (N_15859,N_10995,N_11487);
nor U15860 (N_15860,N_10888,N_10518);
nand U15861 (N_15861,N_8351,N_8011);
or U15862 (N_15862,N_10548,N_10635);
nor U15863 (N_15863,N_11887,N_8202);
nor U15864 (N_15864,N_10829,N_8334);
nand U15865 (N_15865,N_11113,N_10051);
nand U15866 (N_15866,N_8254,N_10260);
or U15867 (N_15867,N_11882,N_9365);
and U15868 (N_15868,N_8970,N_11520);
nand U15869 (N_15869,N_9626,N_8795);
or U15870 (N_15870,N_11327,N_9765);
or U15871 (N_15871,N_8045,N_10549);
nand U15872 (N_15872,N_9582,N_8247);
nor U15873 (N_15873,N_11328,N_10137);
xor U15874 (N_15874,N_10599,N_11757);
or U15875 (N_15875,N_9869,N_10779);
and U15876 (N_15876,N_11295,N_10377);
and U15877 (N_15877,N_11683,N_9171);
or U15878 (N_15878,N_11974,N_11301);
xnor U15879 (N_15879,N_9799,N_9178);
nor U15880 (N_15880,N_11276,N_10214);
nand U15881 (N_15881,N_11268,N_11405);
nor U15882 (N_15882,N_9076,N_8392);
xor U15883 (N_15883,N_11865,N_8336);
nand U15884 (N_15884,N_11342,N_9293);
and U15885 (N_15885,N_11952,N_10193);
nor U15886 (N_15886,N_10125,N_10450);
nand U15887 (N_15887,N_10270,N_11883);
and U15888 (N_15888,N_11569,N_9733);
nand U15889 (N_15889,N_8087,N_8965);
xnor U15890 (N_15890,N_8590,N_8945);
and U15891 (N_15891,N_8092,N_8761);
xnor U15892 (N_15892,N_9515,N_10620);
nor U15893 (N_15893,N_10239,N_10383);
xor U15894 (N_15894,N_8199,N_11241);
nand U15895 (N_15895,N_11275,N_8767);
xnor U15896 (N_15896,N_9132,N_10325);
xnor U15897 (N_15897,N_10808,N_11518);
and U15898 (N_15898,N_11218,N_10894);
and U15899 (N_15899,N_10439,N_9061);
nand U15900 (N_15900,N_10008,N_9338);
nor U15901 (N_15901,N_10557,N_10593);
xor U15902 (N_15902,N_11373,N_10741);
nor U15903 (N_15903,N_9415,N_8871);
xnor U15904 (N_15904,N_9055,N_9095);
nor U15905 (N_15905,N_8887,N_9117);
nor U15906 (N_15906,N_9880,N_11768);
nor U15907 (N_15907,N_10581,N_8704);
xnor U15908 (N_15908,N_9573,N_8135);
nand U15909 (N_15909,N_10591,N_8410);
nand U15910 (N_15910,N_8948,N_10423);
and U15911 (N_15911,N_9423,N_8351);
or U15912 (N_15912,N_9458,N_10766);
and U15913 (N_15913,N_11280,N_9788);
nor U15914 (N_15914,N_11402,N_10855);
nor U15915 (N_15915,N_11033,N_9403);
or U15916 (N_15916,N_8914,N_11020);
and U15917 (N_15917,N_10903,N_10663);
xnor U15918 (N_15918,N_10403,N_8115);
and U15919 (N_15919,N_8211,N_11880);
nand U15920 (N_15920,N_11651,N_11913);
xnor U15921 (N_15921,N_8805,N_10527);
nor U15922 (N_15922,N_8746,N_10758);
or U15923 (N_15923,N_8929,N_9167);
nor U15924 (N_15924,N_10137,N_9712);
and U15925 (N_15925,N_10324,N_8011);
xor U15926 (N_15926,N_11529,N_11897);
nor U15927 (N_15927,N_8944,N_10840);
or U15928 (N_15928,N_10642,N_9781);
and U15929 (N_15929,N_9586,N_8525);
nor U15930 (N_15930,N_11386,N_8431);
xnor U15931 (N_15931,N_9128,N_8259);
nor U15932 (N_15932,N_9655,N_8426);
or U15933 (N_15933,N_9992,N_11070);
xnor U15934 (N_15934,N_8889,N_8027);
and U15935 (N_15935,N_10621,N_9974);
or U15936 (N_15936,N_10388,N_9619);
xnor U15937 (N_15937,N_11529,N_10899);
xor U15938 (N_15938,N_10511,N_10741);
and U15939 (N_15939,N_9771,N_9170);
xnor U15940 (N_15940,N_10899,N_8807);
or U15941 (N_15941,N_10397,N_10332);
and U15942 (N_15942,N_10549,N_10245);
and U15943 (N_15943,N_9077,N_9757);
xor U15944 (N_15944,N_8730,N_8887);
and U15945 (N_15945,N_8974,N_10217);
nor U15946 (N_15946,N_8587,N_8152);
or U15947 (N_15947,N_11253,N_11283);
and U15948 (N_15948,N_11572,N_10901);
and U15949 (N_15949,N_9748,N_10728);
or U15950 (N_15950,N_10941,N_10362);
xor U15951 (N_15951,N_8529,N_9089);
nand U15952 (N_15952,N_9026,N_11709);
nor U15953 (N_15953,N_10754,N_9052);
nor U15954 (N_15954,N_9964,N_10456);
nand U15955 (N_15955,N_10859,N_11431);
nor U15956 (N_15956,N_11405,N_11000);
and U15957 (N_15957,N_11392,N_8577);
nand U15958 (N_15958,N_8601,N_9423);
or U15959 (N_15959,N_9484,N_8920);
nor U15960 (N_15960,N_8358,N_10769);
nor U15961 (N_15961,N_10728,N_8203);
nor U15962 (N_15962,N_8862,N_8532);
and U15963 (N_15963,N_9460,N_10232);
nand U15964 (N_15964,N_9668,N_9786);
or U15965 (N_15965,N_8179,N_11220);
or U15966 (N_15966,N_9112,N_10758);
nor U15967 (N_15967,N_9003,N_10015);
xnor U15968 (N_15968,N_11660,N_9721);
or U15969 (N_15969,N_9971,N_9310);
nor U15970 (N_15970,N_10715,N_11813);
xor U15971 (N_15971,N_11712,N_8551);
nor U15972 (N_15972,N_11975,N_11951);
nor U15973 (N_15973,N_10496,N_10351);
and U15974 (N_15974,N_11314,N_9453);
nand U15975 (N_15975,N_10899,N_11245);
nor U15976 (N_15976,N_8410,N_11365);
nand U15977 (N_15977,N_10444,N_11740);
nor U15978 (N_15978,N_10104,N_10375);
xor U15979 (N_15979,N_11044,N_11431);
or U15980 (N_15980,N_10550,N_9197);
and U15981 (N_15981,N_10636,N_10828);
xnor U15982 (N_15982,N_11859,N_9453);
xor U15983 (N_15983,N_10230,N_8503);
nor U15984 (N_15984,N_8018,N_8927);
nor U15985 (N_15985,N_8028,N_9512);
xor U15986 (N_15986,N_9368,N_10104);
nor U15987 (N_15987,N_11335,N_9852);
nand U15988 (N_15988,N_8857,N_8812);
nor U15989 (N_15989,N_10602,N_11057);
xor U15990 (N_15990,N_8401,N_11019);
or U15991 (N_15991,N_11120,N_9990);
or U15992 (N_15992,N_10192,N_9745);
or U15993 (N_15993,N_10300,N_11452);
or U15994 (N_15994,N_8964,N_9344);
and U15995 (N_15995,N_9682,N_10897);
or U15996 (N_15996,N_10918,N_10683);
nand U15997 (N_15997,N_10585,N_11425);
and U15998 (N_15998,N_9275,N_9161);
or U15999 (N_15999,N_11689,N_8653);
xor U16000 (N_16000,N_12882,N_12437);
and U16001 (N_16001,N_12580,N_13287);
xnor U16002 (N_16002,N_15996,N_14245);
nand U16003 (N_16003,N_15771,N_13640);
and U16004 (N_16004,N_12737,N_15080);
xnor U16005 (N_16005,N_15932,N_15150);
nor U16006 (N_16006,N_14926,N_12077);
or U16007 (N_16007,N_12164,N_12664);
nor U16008 (N_16008,N_14846,N_12517);
xor U16009 (N_16009,N_15674,N_13474);
and U16010 (N_16010,N_12106,N_12797);
or U16011 (N_16011,N_12777,N_15900);
nand U16012 (N_16012,N_15459,N_15672);
or U16013 (N_16013,N_12983,N_13830);
nor U16014 (N_16014,N_14840,N_13059);
or U16015 (N_16015,N_12198,N_13022);
or U16016 (N_16016,N_12323,N_15059);
nor U16017 (N_16017,N_15250,N_15078);
nand U16018 (N_16018,N_13184,N_15185);
nand U16019 (N_16019,N_12819,N_13320);
or U16020 (N_16020,N_12014,N_13834);
xor U16021 (N_16021,N_15325,N_15542);
xor U16022 (N_16022,N_13764,N_13898);
and U16023 (N_16023,N_12374,N_12069);
or U16024 (N_16024,N_12821,N_12035);
or U16025 (N_16025,N_14734,N_14346);
or U16026 (N_16026,N_13170,N_13499);
or U16027 (N_16027,N_13351,N_15854);
nand U16028 (N_16028,N_13255,N_14325);
or U16029 (N_16029,N_12783,N_13386);
and U16030 (N_16030,N_12033,N_13759);
nand U16031 (N_16031,N_12370,N_13027);
xor U16032 (N_16032,N_12810,N_14278);
nor U16033 (N_16033,N_13527,N_15329);
xnor U16034 (N_16034,N_12074,N_12185);
nand U16035 (N_16035,N_14945,N_15376);
and U16036 (N_16036,N_13215,N_15193);
nand U16037 (N_16037,N_13089,N_12419);
nand U16038 (N_16038,N_14550,N_15498);
nor U16039 (N_16039,N_12181,N_13677);
or U16040 (N_16040,N_13708,N_14364);
or U16041 (N_16041,N_14866,N_12174);
and U16042 (N_16042,N_14790,N_15825);
nor U16043 (N_16043,N_15195,N_12604);
nand U16044 (N_16044,N_14353,N_14403);
or U16045 (N_16045,N_13581,N_12108);
or U16046 (N_16046,N_13079,N_13591);
xor U16047 (N_16047,N_14586,N_12829);
nand U16048 (N_16048,N_15123,N_13111);
and U16049 (N_16049,N_15983,N_15326);
or U16050 (N_16050,N_14254,N_13707);
and U16051 (N_16051,N_12787,N_15845);
nand U16052 (N_16052,N_15147,N_13706);
nor U16053 (N_16053,N_12274,N_13742);
xnor U16054 (N_16054,N_13995,N_13421);
xnor U16055 (N_16055,N_15443,N_15169);
or U16056 (N_16056,N_12796,N_15275);
nand U16057 (N_16057,N_12582,N_15151);
or U16058 (N_16058,N_15104,N_13092);
nand U16059 (N_16059,N_12977,N_14295);
nand U16060 (N_16060,N_13722,N_15011);
nor U16061 (N_16061,N_14304,N_13655);
nor U16062 (N_16062,N_13376,N_13015);
nand U16063 (N_16063,N_13267,N_14131);
xor U16064 (N_16064,N_15081,N_13976);
and U16065 (N_16065,N_15593,N_14075);
nand U16066 (N_16066,N_14253,N_14532);
or U16067 (N_16067,N_15849,N_12088);
or U16068 (N_16068,N_13378,N_13063);
nor U16069 (N_16069,N_13841,N_15552);
and U16070 (N_16070,N_12639,N_12306);
xor U16071 (N_16071,N_15844,N_15565);
nand U16072 (N_16072,N_12135,N_15263);
or U16073 (N_16073,N_13020,N_14788);
or U16074 (N_16074,N_12467,N_15172);
nand U16075 (N_16075,N_14252,N_12792);
nand U16076 (N_16076,N_15876,N_13446);
xnor U16077 (N_16077,N_12929,N_12315);
and U16078 (N_16078,N_13788,N_15349);
nand U16079 (N_16079,N_12453,N_13264);
and U16080 (N_16080,N_13638,N_15009);
nand U16081 (N_16081,N_12605,N_14031);
or U16082 (N_16082,N_15190,N_12931);
and U16083 (N_16083,N_12556,N_12563);
or U16084 (N_16084,N_12499,N_14578);
xnor U16085 (N_16085,N_15797,N_14663);
nand U16086 (N_16086,N_13644,N_15830);
nand U16087 (N_16087,N_13046,N_12572);
and U16088 (N_16088,N_14225,N_15543);
xnor U16089 (N_16089,N_12846,N_15311);
nand U16090 (N_16090,N_12221,N_12321);
nor U16091 (N_16091,N_13758,N_13136);
and U16092 (N_16092,N_12403,N_12999);
and U16093 (N_16093,N_14391,N_12836);
nor U16094 (N_16094,N_15430,N_12382);
and U16095 (N_16095,N_14545,N_15563);
and U16096 (N_16096,N_14177,N_12466);
nand U16097 (N_16097,N_13394,N_13437);
nor U16098 (N_16098,N_15574,N_14705);
xor U16099 (N_16099,N_15915,N_12512);
nand U16100 (N_16100,N_15236,N_13907);
and U16101 (N_16101,N_13945,N_15020);
or U16102 (N_16102,N_12126,N_12237);
nor U16103 (N_16103,N_13428,N_14222);
and U16104 (N_16104,N_14337,N_13458);
or U16105 (N_16105,N_13879,N_15053);
or U16106 (N_16106,N_13395,N_14009);
and U16107 (N_16107,N_13893,N_12099);
nor U16108 (N_16108,N_15513,N_13712);
xor U16109 (N_16109,N_15972,N_14236);
nor U16110 (N_16110,N_12723,N_12114);
xnor U16111 (N_16111,N_12961,N_13539);
and U16112 (N_16112,N_15790,N_12579);
nor U16113 (N_16113,N_12417,N_15656);
or U16114 (N_16114,N_15105,N_14292);
or U16115 (N_16115,N_15731,N_12061);
nand U16116 (N_16116,N_15526,N_13784);
or U16117 (N_16117,N_12474,N_15499);
xor U16118 (N_16118,N_15461,N_12159);
nand U16119 (N_16119,N_15170,N_13142);
nor U16120 (N_16120,N_13551,N_13949);
and U16121 (N_16121,N_15088,N_13336);
nand U16122 (N_16122,N_14070,N_15463);
or U16123 (N_16123,N_14171,N_13925);
or U16124 (N_16124,N_13628,N_13082);
nor U16125 (N_16125,N_15562,N_15191);
or U16126 (N_16126,N_15743,N_12113);
or U16127 (N_16127,N_12353,N_14995);
xnor U16128 (N_16128,N_15622,N_12213);
and U16129 (N_16129,N_14659,N_14459);
xor U16130 (N_16130,N_12162,N_12122);
xnor U16131 (N_16131,N_14609,N_13013);
nor U16132 (N_16132,N_15372,N_14849);
xnor U16133 (N_16133,N_14025,N_15717);
nor U16134 (N_16134,N_14821,N_12393);
nor U16135 (N_16135,N_15730,N_13629);
or U16136 (N_16136,N_15165,N_13006);
nor U16137 (N_16137,N_14921,N_12133);
nor U16138 (N_16138,N_13994,N_13980);
or U16139 (N_16139,N_12793,N_13308);
and U16140 (N_16140,N_12594,N_12470);
and U16141 (N_16141,N_12610,N_12085);
and U16142 (N_16142,N_13623,N_12071);
and U16143 (N_16143,N_13954,N_12188);
and U16144 (N_16144,N_12973,N_15576);
or U16145 (N_16145,N_14029,N_13114);
and U16146 (N_16146,N_15440,N_13248);
or U16147 (N_16147,N_15684,N_15164);
or U16148 (N_16148,N_15187,N_15599);
and U16149 (N_16149,N_13097,N_14877);
nor U16150 (N_16150,N_15503,N_15196);
and U16151 (N_16151,N_14049,N_15130);
xor U16152 (N_16152,N_14473,N_15194);
xnor U16153 (N_16153,N_15006,N_15990);
nor U16154 (N_16154,N_13187,N_14852);
and U16155 (N_16155,N_15056,N_13253);
or U16156 (N_16156,N_13525,N_13433);
xor U16157 (N_16157,N_13771,N_13066);
and U16158 (N_16158,N_14328,N_15726);
nand U16159 (N_16159,N_12666,N_12756);
nand U16160 (N_16160,N_15505,N_15457);
or U16161 (N_16161,N_13896,N_12967);
and U16162 (N_16162,N_12290,N_13095);
or U16163 (N_16163,N_13298,N_13178);
xor U16164 (N_16164,N_13947,N_14247);
and U16165 (N_16165,N_14448,N_15560);
nand U16166 (N_16166,N_12758,N_13019);
and U16167 (N_16167,N_12359,N_12506);
and U16168 (N_16168,N_13779,N_13508);
nand U16169 (N_16169,N_13209,N_13807);
nand U16170 (N_16170,N_12678,N_13943);
or U16171 (N_16171,N_12392,N_15813);
and U16172 (N_16172,N_15532,N_14483);
or U16173 (N_16173,N_13414,N_15448);
nor U16174 (N_16174,N_15288,N_14092);
xnor U16175 (N_16175,N_13353,N_13439);
and U16176 (N_16176,N_14434,N_14213);
or U16177 (N_16177,N_15716,N_14149);
nor U16178 (N_16178,N_15154,N_13825);
nor U16179 (N_16179,N_13188,N_15048);
or U16180 (N_16180,N_14676,N_15366);
or U16181 (N_16181,N_14237,N_13148);
or U16182 (N_16182,N_14262,N_13609);
xor U16183 (N_16183,N_12492,N_15284);
nor U16184 (N_16184,N_12719,N_13803);
nand U16185 (N_16185,N_13042,N_12934);
and U16186 (N_16186,N_12441,N_14885);
nand U16187 (N_16187,N_12954,N_13660);
or U16188 (N_16188,N_15874,N_13272);
nand U16189 (N_16189,N_12710,N_14802);
and U16190 (N_16190,N_13300,N_14801);
or U16191 (N_16191,N_14428,N_12505);
xor U16192 (N_16192,N_12659,N_12372);
nand U16193 (N_16193,N_12129,N_15761);
and U16194 (N_16194,N_15801,N_12804);
xor U16195 (N_16195,N_13808,N_14861);
xor U16196 (N_16196,N_12850,N_14842);
and U16197 (N_16197,N_13971,N_15392);
and U16198 (N_16198,N_14670,N_15867);
xor U16199 (N_16199,N_15052,N_15084);
nor U16200 (N_16200,N_14641,N_15939);
xnor U16201 (N_16201,N_12500,N_15507);
and U16202 (N_16202,N_15438,N_13028);
or U16203 (N_16203,N_15781,N_14182);
and U16204 (N_16204,N_12876,N_12769);
nor U16205 (N_16205,N_12620,N_14421);
or U16206 (N_16206,N_14285,N_12540);
and U16207 (N_16207,N_12806,N_12713);
or U16208 (N_16208,N_15571,N_14652);
nand U16209 (N_16209,N_13150,N_14637);
xnor U16210 (N_16210,N_14721,N_14128);
or U16211 (N_16211,N_13423,N_13373);
and U16212 (N_16212,N_12352,N_14186);
or U16213 (N_16213,N_12964,N_15699);
nand U16214 (N_16214,N_15252,N_15749);
xor U16215 (N_16215,N_15493,N_12595);
or U16216 (N_16216,N_15982,N_13494);
nor U16217 (N_16217,N_13674,N_12059);
or U16218 (N_16218,N_12124,N_14927);
or U16219 (N_16219,N_13067,N_13972);
and U16220 (N_16220,N_15295,N_13313);
and U16221 (N_16221,N_14482,N_13231);
xor U16222 (N_16222,N_15721,N_13309);
xnor U16223 (N_16223,N_13648,N_13730);
and U16224 (N_16224,N_15540,N_13192);
and U16225 (N_16225,N_15875,N_13865);
and U16226 (N_16226,N_13147,N_15539);
or U16227 (N_16227,N_14903,N_12823);
xnor U16228 (N_16228,N_14235,N_14754);
and U16229 (N_16229,N_12241,N_13738);
nor U16230 (N_16230,N_13563,N_15551);
nand U16231 (N_16231,N_12468,N_12490);
nor U16232 (N_16232,N_13476,N_13751);
or U16233 (N_16233,N_14430,N_12489);
xnor U16234 (N_16234,N_12337,N_14993);
and U16235 (N_16235,N_13578,N_12178);
nor U16236 (N_16236,N_12865,N_13139);
nor U16237 (N_16237,N_12004,N_13488);
nor U16238 (N_16238,N_14134,N_12996);
nand U16239 (N_16239,N_12867,N_13401);
or U16240 (N_16240,N_15803,N_12825);
nor U16241 (N_16241,N_12957,N_12699);
and U16242 (N_16242,N_12767,N_12084);
xnor U16243 (N_16243,N_13454,N_12495);
nor U16244 (N_16244,N_12502,N_15634);
nor U16245 (N_16245,N_13862,N_12974);
nor U16246 (N_16246,N_12263,N_13535);
xnor U16247 (N_16247,N_14174,N_13832);
or U16248 (N_16248,N_12262,N_14239);
or U16249 (N_16249,N_12948,N_14108);
xnor U16250 (N_16250,N_14716,N_14965);
nor U16251 (N_16251,N_13921,N_14624);
nor U16252 (N_16252,N_12078,N_13164);
nand U16253 (N_16253,N_15695,N_15467);
or U16254 (N_16254,N_12559,N_14494);
xnor U16255 (N_16255,N_15579,N_15268);
xor U16256 (N_16256,N_14739,N_13237);
nand U16257 (N_16257,N_15414,N_14095);
and U16258 (N_16258,N_15024,N_12730);
or U16259 (N_16259,N_14850,N_13393);
or U16260 (N_16260,N_15387,N_15709);
or U16261 (N_16261,N_15863,N_15073);
and U16262 (N_16262,N_14529,N_14071);
and U16263 (N_16263,N_15219,N_13419);
or U16264 (N_16264,N_14557,N_13005);
and U16265 (N_16265,N_15424,N_13033);
or U16266 (N_16266,N_15842,N_14612);
nand U16267 (N_16267,N_13647,N_12802);
or U16268 (N_16268,N_15428,N_12469);
xor U16269 (N_16269,N_12432,N_14859);
nor U16270 (N_16270,N_13791,N_13489);
and U16271 (N_16271,N_12383,N_15008);
xnor U16272 (N_16272,N_13060,N_12038);
nor U16273 (N_16273,N_13854,N_14323);
or U16274 (N_16274,N_15364,N_13641);
nand U16275 (N_16275,N_14013,N_15872);
or U16276 (N_16276,N_12454,N_13897);
and U16277 (N_16277,N_12485,N_12643);
or U16278 (N_16278,N_13481,N_14895);
xnor U16279 (N_16279,N_14643,N_15316);
nor U16280 (N_16280,N_13910,N_13141);
nand U16281 (N_16281,N_14297,N_12048);
or U16282 (N_16282,N_13358,N_12401);
nor U16283 (N_16283,N_15703,N_12458);
nand U16284 (N_16284,N_12310,N_12529);
xnor U16285 (N_16285,N_13314,N_15665);
xor U16286 (N_16286,N_14202,N_14219);
or U16287 (N_16287,N_13661,N_13687);
and U16288 (N_16288,N_14369,N_15332);
nand U16289 (N_16289,N_15969,N_13777);
xor U16290 (N_16290,N_13347,N_13534);
nand U16291 (N_16291,N_15917,N_15533);
nand U16292 (N_16292,N_14540,N_14354);
and U16293 (N_16293,N_13021,N_14246);
and U16294 (N_16294,N_14488,N_14829);
or U16295 (N_16295,N_12155,N_15319);
and U16296 (N_16296,N_14991,N_14521);
or U16297 (N_16297,N_14525,N_13852);
and U16298 (N_16298,N_13983,N_12762);
and U16299 (N_16299,N_12984,N_12227);
nor U16300 (N_16300,N_13953,N_14674);
xnor U16301 (N_16301,N_15553,N_12010);
and U16302 (N_16302,N_14729,N_13658);
nand U16303 (N_16303,N_14946,N_15971);
xnor U16304 (N_16304,N_14610,N_13344);
nor U16305 (N_16305,N_15166,N_15940);
xnor U16306 (N_16306,N_15663,N_15118);
and U16307 (N_16307,N_14874,N_12543);
xnor U16308 (N_16308,N_12438,N_12247);
nor U16309 (N_16309,N_14543,N_13703);
or U16310 (N_16310,N_13819,N_14210);
and U16311 (N_16311,N_12504,N_15698);
nand U16312 (N_16312,N_14294,N_13600);
nand U16313 (N_16313,N_15145,N_13554);
nand U16314 (N_16314,N_13269,N_15348);
or U16315 (N_16315,N_12422,N_12537);
nor U16316 (N_16316,N_15626,N_12591);
or U16317 (N_16317,N_12739,N_15029);
xnor U16318 (N_16318,N_14124,N_15175);
nor U16319 (N_16319,N_12276,N_12457);
nor U16320 (N_16320,N_14644,N_13686);
xnor U16321 (N_16321,N_15235,N_13811);
nand U16322 (N_16322,N_12350,N_13222);
xnor U16323 (N_16323,N_13866,N_12239);
xor U16324 (N_16324,N_15478,N_12363);
nand U16325 (N_16325,N_13895,N_13950);
or U16326 (N_16326,N_13462,N_14417);
and U16327 (N_16327,N_14797,N_15812);
xor U16328 (N_16328,N_15705,N_13726);
nor U16329 (N_16329,N_13176,N_15259);
xor U16330 (N_16330,N_15984,N_15559);
or U16331 (N_16331,N_13933,N_15907);
nor U16332 (N_16332,N_15421,N_13579);
xnor U16333 (N_16333,N_13214,N_14580);
xnor U16334 (N_16334,N_13390,N_14933);
nor U16335 (N_16335,N_15847,N_13472);
nor U16336 (N_16336,N_14238,N_14335);
and U16337 (N_16337,N_15411,N_14197);
nand U16338 (N_16338,N_15327,N_12726);
and U16339 (N_16339,N_13704,N_14456);
nand U16340 (N_16340,N_12448,N_12602);
nor U16341 (N_16341,N_14475,N_15436);
nor U16342 (N_16342,N_13818,N_12011);
xnor U16343 (N_16343,N_15291,N_14605);
and U16344 (N_16344,N_13705,N_12960);
and U16345 (N_16345,N_15470,N_13870);
nand U16346 (N_16346,N_13616,N_13205);
nor U16347 (N_16347,N_15257,N_15851);
nand U16348 (N_16348,N_13285,N_12346);
or U16349 (N_16349,N_14098,N_15342);
xor U16350 (N_16350,N_12523,N_12390);
or U16351 (N_16351,N_13306,N_13786);
xnor U16352 (N_16352,N_12658,N_15535);
or U16353 (N_16353,N_12897,N_13589);
xnor U16354 (N_16354,N_14072,N_13057);
xor U16355 (N_16355,N_14706,N_14195);
and U16356 (N_16356,N_12736,N_13877);
and U16357 (N_16357,N_13682,N_13475);
nand U16358 (N_16358,N_12914,N_13168);
nand U16359 (N_16359,N_15636,N_13024);
nor U16360 (N_16360,N_14748,N_15361);
xnor U16361 (N_16361,N_12808,N_13783);
and U16362 (N_16362,N_12773,N_15811);
nor U16363 (N_16363,N_12298,N_14052);
xnor U16364 (N_16364,N_15210,N_13557);
xor U16365 (N_16365,N_12745,N_15742);
xnor U16366 (N_16366,N_15637,N_13831);
and U16367 (N_16367,N_13604,N_12478);
or U16368 (N_16368,N_15584,N_12528);
nand U16369 (N_16369,N_12901,N_13690);
xor U16370 (N_16370,N_13070,N_15136);
nand U16371 (N_16371,N_12794,N_15287);
or U16372 (N_16372,N_15765,N_12013);
xor U16373 (N_16373,N_14433,N_12105);
or U16374 (N_16374,N_15736,N_13723);
or U16375 (N_16375,N_13460,N_14218);
nand U16376 (N_16376,N_13871,N_12313);
nand U16377 (N_16377,N_14169,N_14374);
or U16378 (N_16378,N_12863,N_13553);
or U16379 (N_16379,N_13915,N_14296);
nand U16380 (N_16380,N_13464,N_15768);
xor U16381 (N_16381,N_14330,N_13729);
nor U16382 (N_16382,N_15920,N_12570);
or U16383 (N_16383,N_14712,N_13333);
nor U16384 (N_16384,N_13103,N_15737);
nand U16385 (N_16385,N_15831,N_12923);
nand U16386 (N_16386,N_14261,N_15102);
nand U16387 (N_16387,N_15955,N_12317);
nor U16388 (N_16388,N_12548,N_12141);
xnor U16389 (N_16389,N_14793,N_14851);
nand U16390 (N_16390,N_12590,N_13328);
or U16391 (N_16391,N_12979,N_13008);
nor U16392 (N_16392,N_15755,N_12307);
xor U16393 (N_16393,N_14227,N_12361);
nand U16394 (N_16394,N_13653,N_15619);
and U16395 (N_16395,N_14603,N_13816);
nor U16396 (N_16396,N_14479,N_12619);
nor U16397 (N_16397,N_15063,N_15594);
or U16398 (N_16398,N_12644,N_13032);
nand U16399 (N_16399,N_13931,N_14023);
xor U16400 (N_16400,N_14981,N_15671);
or U16401 (N_16401,N_15282,N_12456);
nor U16402 (N_16402,N_15077,N_15799);
nand U16403 (N_16403,N_12680,N_15946);
or U16404 (N_16404,N_14176,N_13670);
nand U16405 (N_16405,N_13696,N_15121);
nand U16406 (N_16406,N_13405,N_14002);
or U16407 (N_16407,N_13977,N_14474);
nor U16408 (N_16408,N_14229,N_13829);
xnor U16409 (N_16409,N_14667,N_13463);
xnor U16410 (N_16410,N_15711,N_14635);
xor U16411 (N_16411,N_14458,N_14085);
and U16412 (N_16412,N_13937,N_12925);
nor U16413 (N_16413,N_15837,N_15887);
nor U16414 (N_16414,N_12827,N_12812);
xor U16415 (N_16415,N_12910,N_15167);
nor U16416 (N_16416,N_12172,N_14226);
nor U16417 (N_16417,N_12840,N_15509);
or U16418 (N_16418,N_15527,N_14959);
or U16419 (N_16419,N_15776,N_12640);
or U16420 (N_16420,N_12215,N_12732);
and U16421 (N_16421,N_13480,N_12053);
or U16422 (N_16422,N_12279,N_13238);
nor U16423 (N_16423,N_13608,N_15089);
nand U16424 (N_16424,N_15477,N_12131);
and U16425 (N_16425,N_14552,N_14028);
and U16426 (N_16426,N_13580,N_15489);
xnor U16427 (N_16427,N_14898,N_14435);
nand U16428 (N_16428,N_12801,N_13040);
nand U16429 (N_16429,N_13860,N_12212);
xnor U16430 (N_16430,N_14655,N_15877);
or U16431 (N_16431,N_14107,N_14708);
xor U16432 (N_16432,N_13531,N_14463);
or U16433 (N_16433,N_13888,N_15404);
nor U16434 (N_16434,N_12180,N_13257);
or U16435 (N_16435,N_13851,N_13117);
nor U16436 (N_16436,N_15740,N_13266);
nand U16437 (N_16437,N_13668,N_15353);
and U16438 (N_16438,N_15680,N_12627);
xor U16439 (N_16439,N_13193,N_15836);
nand U16440 (N_16440,N_12667,N_12638);
or U16441 (N_16441,N_15787,N_15292);
nor U16442 (N_16442,N_12729,N_13802);
xor U16443 (N_16443,N_13391,N_15788);
xnor U16444 (N_16444,N_13767,N_15521);
xnor U16445 (N_16445,N_14614,N_13043);
xnor U16446 (N_16446,N_15143,N_13076);
and U16447 (N_16447,N_13339,N_13913);
xor U16448 (N_16448,N_15911,N_13512);
nand U16449 (N_16449,N_12975,N_14478);
xor U16450 (N_16450,N_13191,N_15065);
nand U16451 (N_16451,N_15902,N_14162);
or U16452 (N_16452,N_12988,N_12269);
xnor U16453 (N_16453,N_12338,N_12883);
nand U16454 (N_16454,N_14810,N_13382);
nor U16455 (N_16455,N_13836,N_12717);
nand U16456 (N_16456,N_15176,N_12246);
or U16457 (N_16457,N_12872,N_14172);
xnor U16458 (N_16458,N_15979,N_15639);
and U16459 (N_16459,N_13217,N_14639);
and U16460 (N_16460,N_15265,N_13226);
nand U16461 (N_16461,N_12508,N_13543);
and U16462 (N_16462,N_12308,N_14066);
and U16463 (N_16463,N_14394,N_12847);
or U16464 (N_16464,N_12301,N_15091);
nor U16465 (N_16465,N_13304,N_14350);
xor U16466 (N_16466,N_13235,N_12642);
nor U16467 (N_16467,N_13855,N_13485);
nor U16468 (N_16468,N_12860,N_12493);
nand U16469 (N_16469,N_15362,N_12153);
nor U16470 (N_16470,N_13547,N_13922);
nand U16471 (N_16471,N_13174,N_14042);
xnor U16472 (N_16472,N_12054,N_14536);
and U16473 (N_16473,N_14372,N_12754);
nand U16474 (N_16474,N_12685,N_15808);
and U16475 (N_16475,N_14512,N_14707);
and U16476 (N_16476,N_12163,N_15850);
nor U16477 (N_16477,N_14437,N_15100);
nor U16478 (N_16478,N_12597,N_15927);
nand U16479 (N_16479,N_15642,N_14665);
xnor U16480 (N_16480,N_13853,N_13254);
nand U16481 (N_16481,N_14590,N_14560);
nand U16482 (N_16482,N_14228,N_12412);
nand U16483 (N_16483,N_12748,N_13324);
nor U16484 (N_16484,N_13611,N_15388);
nor U16485 (N_16485,N_12603,N_14360);
and U16486 (N_16486,N_15155,N_13530);
or U16487 (N_16487,N_15606,N_13282);
and U16488 (N_16488,N_15465,N_14882);
xnor U16489 (N_16489,N_15464,N_14027);
and U16490 (N_16490,N_13119,N_13582);
and U16491 (N_16491,N_14607,N_13920);
or U16492 (N_16492,N_14104,N_13025);
nor U16493 (N_16493,N_12063,N_12677);
xnor U16494 (N_16494,N_14701,N_14444);
nor U16495 (N_16495,N_14484,N_12583);
or U16496 (N_16496,N_14116,N_15798);
and U16497 (N_16497,N_12574,N_15545);
or U16498 (N_16498,N_12888,N_14975);
nand U16499 (N_16499,N_14264,N_13004);
nand U16500 (N_16500,N_15022,N_15442);
or U16501 (N_16501,N_13216,N_15040);
or U16502 (N_16502,N_14973,N_13612);
xnor U16503 (N_16503,N_15638,N_14997);
or U16504 (N_16504,N_12673,N_15816);
xor U16505 (N_16505,N_14809,N_14731);
nor U16506 (N_16506,N_13121,N_13389);
or U16507 (N_16507,N_14276,N_14367);
xor U16508 (N_16508,N_15108,N_13936);
or U16509 (N_16509,N_14854,N_14280);
nand U16510 (N_16510,N_14400,N_13346);
and U16511 (N_16511,N_12220,N_15094);
and U16512 (N_16512,N_13633,N_12270);
nand U16513 (N_16513,N_15086,N_12446);
or U16514 (N_16514,N_15839,N_13327);
and U16515 (N_16515,N_14196,N_12297);
or U16516 (N_16516,N_12148,N_15242);
nand U16517 (N_16517,N_14971,N_14507);
or U16518 (N_16518,N_13172,N_14918);
xor U16519 (N_16519,N_14121,N_15358);
and U16520 (N_16520,N_14929,N_13160);
or U16521 (N_16521,N_15171,N_12550);
nor U16522 (N_16522,N_12991,N_13984);
xor U16523 (N_16523,N_15814,N_14650);
xor U16524 (N_16524,N_13691,N_12008);
nand U16525 (N_16525,N_13135,N_13597);
nor U16526 (N_16526,N_13881,N_14270);
and U16527 (N_16527,N_15794,N_15449);
nor U16528 (N_16528,N_14782,N_15415);
nand U16529 (N_16529,N_15775,N_12449);
and U16530 (N_16530,N_12959,N_14604);
or U16531 (N_16531,N_15273,N_12027);
xor U16532 (N_16532,N_13289,N_12637);
or U16533 (N_16533,N_13334,N_13843);
nor U16534 (N_16534,N_13856,N_13528);
nand U16535 (N_16535,N_15994,N_13301);
and U16536 (N_16536,N_12036,N_14241);
and U16537 (N_16537,N_15862,N_12322);
or U16538 (N_16538,N_12849,N_12158);
nor U16539 (N_16539,N_14244,N_15061);
nand U16540 (N_16540,N_15588,N_15738);
nand U16541 (N_16541,N_14271,N_14401);
and U16542 (N_16542,N_12562,N_13762);
xor U16543 (N_16543,N_13354,N_14515);
xor U16544 (N_16544,N_12486,N_15031);
nand U16545 (N_16545,N_15756,N_14205);
nor U16546 (N_16546,N_14682,N_15723);
nor U16547 (N_16547,N_12628,N_15913);
nand U16548 (N_16548,N_13569,N_15537);
and U16549 (N_16549,N_14425,N_12521);
and U16550 (N_16550,N_14158,N_14646);
xor U16551 (N_16551,N_14273,N_12705);
or U16552 (N_16552,N_15573,N_15324);
nor U16553 (N_16553,N_14167,N_14907);
nand U16554 (N_16554,N_13912,N_12051);
or U16555 (N_16555,N_15377,N_14648);
nor U16556 (N_16556,N_14690,N_12515);
nand U16557 (N_16557,N_13434,N_13938);
and U16558 (N_16558,N_12039,N_14890);
and U16559 (N_16559,N_14952,N_15728);
xnor U16560 (N_16560,N_15382,N_14187);
and U16561 (N_16561,N_15481,N_13709);
or U16562 (N_16562,N_12940,N_14979);
nor U16563 (N_16563,N_12264,N_13335);
or U16564 (N_16564,N_15531,N_12768);
or U16565 (N_16565,N_12725,N_12389);
xnor U16566 (N_16566,N_14977,N_12171);
nand U16567 (N_16567,N_15959,N_15400);
nor U16568 (N_16568,N_15796,N_15780);
nand U16569 (N_16569,N_15114,N_13908);
or U16570 (N_16570,N_13071,N_15398);
and U16571 (N_16571,N_14151,N_15646);
nor U16572 (N_16572,N_15903,N_15930);
and U16573 (N_16573,N_14626,N_14059);
xnor U16574 (N_16574,N_14137,N_15510);
nor U16575 (N_16575,N_14825,N_12833);
nand U16576 (N_16576,N_12995,N_14404);
or U16577 (N_16577,N_15032,N_12367);
nand U16578 (N_16578,N_14180,N_12214);
or U16579 (N_16579,N_13765,N_14796);
and U16580 (N_16580,N_13650,N_14978);
nand U16581 (N_16581,N_15225,N_13250);
or U16582 (N_16582,N_15654,N_13990);
nor U16583 (N_16583,N_12939,N_12904);
or U16584 (N_16584,N_13167,N_14048);
or U16585 (N_16585,N_14634,N_14514);
nand U16586 (N_16586,N_14054,N_15370);
nor U16587 (N_16587,N_12413,N_15950);
and U16588 (N_16588,N_13133,N_15587);
or U16589 (N_16589,N_15386,N_13228);
xnor U16590 (N_16590,N_14998,N_13755);
nand U16591 (N_16591,N_14198,N_13331);
xnor U16592 (N_16592,N_13903,N_12226);
nor U16593 (N_16593,N_15848,N_15157);
nor U16594 (N_16594,N_14856,N_12139);
nand U16595 (N_16595,N_12165,N_12329);
nand U16596 (N_16596,N_12320,N_12874);
or U16597 (N_16597,N_14365,N_13445);
xor U16598 (N_16598,N_13244,N_12296);
nand U16599 (N_16599,N_15026,N_13370);
nand U16600 (N_16600,N_12411,N_15152);
or U16601 (N_16601,N_15965,N_13737);
or U16602 (N_16602,N_15623,N_14133);
or U16603 (N_16603,N_13520,N_15033);
and U16604 (N_16604,N_15868,N_13630);
xor U16605 (N_16605,N_15318,N_14003);
xor U16606 (N_16606,N_13754,N_13408);
nand U16607 (N_16607,N_14363,N_12324);
xnor U16608 (N_16608,N_13262,N_12044);
nand U16609 (N_16609,N_15251,N_12568);
xnor U16610 (N_16610,N_14622,N_13506);
xor U16611 (N_16611,N_13493,N_12881);
or U16612 (N_16612,N_15581,N_12990);
or U16613 (N_16613,N_13400,N_15653);
nor U16614 (N_16614,N_13441,N_12421);
nor U16615 (N_16615,N_14980,N_12358);
and U16616 (N_16616,N_13030,N_15947);
nor U16617 (N_16617,N_12464,N_13124);
xnor U16618 (N_16618,N_14316,N_15504);
xnor U16619 (N_16619,N_14014,N_15834);
and U16620 (N_16620,N_13247,N_15708);
nor U16621 (N_16621,N_13817,N_12727);
xnor U16622 (N_16622,N_12908,N_13087);
and U16623 (N_16623,N_13500,N_15297);
nand U16624 (N_16624,N_14897,N_13302);
and U16625 (N_16625,N_12192,N_14828);
nor U16626 (N_16626,N_15517,N_13715);
and U16627 (N_16627,N_13727,N_14234);
xnor U16628 (N_16628,N_12652,N_15884);
xnor U16629 (N_16629,N_13397,N_13839);
nand U16630 (N_16630,N_12918,N_12123);
nand U16631 (N_16631,N_15135,N_13521);
or U16632 (N_16632,N_14232,N_12067);
or U16633 (N_16633,N_14383,N_15230);
and U16634 (N_16634,N_14037,N_15394);
or U16635 (N_16635,N_12491,N_15807);
or U16636 (N_16636,N_12657,N_15352);
nand U16637 (N_16637,N_15233,N_14157);
or U16638 (N_16638,N_15981,N_14007);
xnor U16639 (N_16639,N_12462,N_14221);
nor U16640 (N_16640,N_14787,N_12703);
nor U16641 (N_16641,N_13171,N_15338);
nor U16642 (N_16642,N_13774,N_12944);
and U16643 (N_16643,N_12023,N_14672);
nor U16644 (N_16644,N_12613,N_14083);
nor U16645 (N_16645,N_13260,N_13055);
xnor U16646 (N_16646,N_15840,N_12140);
nor U16647 (N_16647,N_12381,N_12718);
nor U16648 (N_16648,N_12744,N_13805);
xor U16649 (N_16649,N_13835,N_13924);
nand U16650 (N_16650,N_15615,N_14230);
xnor U16651 (N_16651,N_15603,N_13740);
and U16652 (N_16652,N_13483,N_14519);
and U16653 (N_16653,N_15929,N_14163);
or U16654 (N_16654,N_15544,N_15514);
and U16655 (N_16655,N_15770,N_13118);
and U16656 (N_16656,N_13126,N_13958);
xor U16657 (N_16657,N_12200,N_14865);
nor U16658 (N_16658,N_14553,N_13477);
and U16659 (N_16659,N_13974,N_12333);
and U16660 (N_16660,N_13091,N_13849);
xor U16661 (N_16661,N_15004,N_14056);
nor U16662 (N_16662,N_14664,N_15924);
xor U16663 (N_16663,N_14284,N_13223);
or U16664 (N_16664,N_12919,N_13820);
and U16665 (N_16665,N_13241,N_14308);
xnor U16666 (N_16666,N_15970,N_14858);
nand U16667 (N_16667,N_14546,N_12423);
and U16668 (N_16668,N_14678,N_15962);
or U16669 (N_16669,N_13096,N_13145);
nor U16670 (N_16670,N_13473,N_15179);
and U16671 (N_16671,N_13775,N_12782);
nand U16672 (N_16672,N_14442,N_13497);
or U16673 (N_16673,N_15492,N_12839);
nor U16674 (N_16674,N_13000,N_13662);
nand U16675 (N_16675,N_15016,N_13471);
nor U16676 (N_16676,N_13252,N_14688);
or U16677 (N_16677,N_13234,N_14853);
nand U16678 (N_16678,N_15043,N_15473);
and U16679 (N_16679,N_12343,N_15616);
xnor U16680 (N_16680,N_15309,N_14733);
nor U16681 (N_16681,N_13542,N_12184);
and U16682 (N_16682,N_14772,N_13678);
nor U16683 (N_16683,N_14875,N_15870);
or U16684 (N_16684,N_14508,N_14936);
or U16685 (N_16685,N_14632,N_12197);
xnor U16686 (N_16686,N_12609,N_15676);
or U16687 (N_16687,N_15068,N_12647);
or U16688 (N_16688,N_12848,N_12895);
or U16689 (N_16689,N_14776,N_13794);
nand U16690 (N_16690,N_14347,N_15330);
and U16691 (N_16691,N_14982,N_12788);
xnor U16692 (N_16692,N_13567,N_12784);
nand U16693 (N_16693,N_15751,N_12554);
nor U16694 (N_16694,N_14331,N_13203);
xnor U16695 (N_16695,N_12127,N_13149);
or U16696 (N_16696,N_14375,N_15036);
and U16697 (N_16697,N_12626,N_15023);
nor U16698 (N_16698,N_15450,N_13402);
or U16699 (N_16699,N_12708,N_15206);
nand U16700 (N_16700,N_15437,N_12532);
nor U16701 (N_16701,N_15451,N_15276);
and U16702 (N_16702,N_13200,N_12599);
and U16703 (N_16703,N_14393,N_12531);
and U16704 (N_16704,N_13761,N_14361);
or U16705 (N_16705,N_12080,N_14556);
xor U16706 (N_16706,N_15446,N_14267);
nand U16707 (N_16707,N_13699,N_12786);
xnor U16708 (N_16708,N_15296,N_15246);
nor U16709 (N_16709,N_14723,N_14913);
or U16710 (N_16710,N_14935,N_13568);
nor U16711 (N_16711,N_14817,N_14832);
or U16712 (N_16712,N_14891,N_13470);
nor U16713 (N_16713,N_14358,N_15058);
xor U16714 (N_16714,N_14275,N_13337);
and U16715 (N_16715,N_15395,N_12955);
xnor U16716 (N_16716,N_12146,N_15051);
nor U16717 (N_16717,N_15878,N_15585);
and U16718 (N_16718,N_13105,N_15216);
nor U16719 (N_16719,N_15713,N_14770);
nand U16720 (N_16720,N_15298,N_12488);
nand U16721 (N_16721,N_14283,N_14340);
and U16722 (N_16722,N_15772,N_12404);
and U16723 (N_16723,N_13261,N_14565);
xnor U16724 (N_16724,N_14505,N_15957);
or U16725 (N_16725,N_13078,N_15027);
and U16726 (N_16726,N_15733,N_12096);
and U16727 (N_16727,N_12230,N_15696);
or U16728 (N_16728,N_12968,N_15591);
and U16729 (N_16729,N_15126,N_13982);
and U16730 (N_16730,N_13695,N_12541);
or U16731 (N_16731,N_15312,N_14461);
xor U16732 (N_16732,N_13173,N_12418);
nand U16733 (N_16733,N_13772,N_14287);
xnor U16734 (N_16734,N_13763,N_13750);
or U16735 (N_16735,N_13332,N_13281);
nor U16736 (N_16736,N_15555,N_15958);
nand U16737 (N_16737,N_14203,N_13606);
nor U16738 (N_16738,N_12378,N_15439);
nor U16739 (N_16739,N_15764,N_14577);
nand U16740 (N_16740,N_15754,N_12302);
xnor U16741 (N_16741,N_12779,N_14735);
nor U16742 (N_16742,N_14411,N_14179);
and U16743 (N_16743,N_13587,N_15163);
or U16744 (N_16744,N_14055,N_12345);
nor U16745 (N_16745,N_13352,N_14691);
and U16746 (N_16746,N_14068,N_12526);
nor U16747 (N_16747,N_14117,N_12932);
or U16748 (N_16748,N_12208,N_13955);
nand U16749 (N_16749,N_12982,N_13544);
or U16750 (N_16750,N_12107,N_15782);
and U16751 (N_16751,N_13728,N_15628);
and U16752 (N_16752,N_13486,N_12497);
and U16753 (N_16753,N_14570,N_12408);
or U16754 (N_16754,N_12190,N_12356);
or U16755 (N_16755,N_13733,N_14497);
nand U16756 (N_16756,N_14291,N_13665);
or U16757 (N_16757,N_13109,N_13080);
xor U16758 (N_16758,N_12871,N_14061);
or U16759 (N_16759,N_12242,N_15524);
nand U16760 (N_16760,N_15487,N_12130);
nand U16761 (N_16761,N_15741,N_12072);
and U16762 (N_16762,N_14129,N_13054);
nand U16763 (N_16763,N_13128,N_15883);
xor U16764 (N_16764,N_12785,N_13194);
nor U16765 (N_16765,N_14593,N_15144);
or U16766 (N_16766,N_13689,N_12075);
and U16767 (N_16767,N_12906,N_14764);
nand U16768 (N_16768,N_14113,N_13996);
nor U16769 (N_16769,N_14259,N_13732);
nor U16770 (N_16770,N_15334,N_15986);
and U16771 (N_16771,N_12941,N_15631);
or U16772 (N_16772,N_15538,N_15759);
xor U16773 (N_16773,N_13154,N_14348);
nor U16774 (N_16774,N_13566,N_14420);
xnor U16775 (N_16775,N_15098,N_15383);
xnor U16776 (N_16776,N_15718,N_12318);
nor U16777 (N_16777,N_15855,N_13813);
nand U16778 (N_16778,N_15649,N_14847);
or U16779 (N_16779,N_12924,N_15692);
and U16780 (N_16780,N_12444,N_15534);
and U16781 (N_16781,N_14034,N_15746);
nand U16782 (N_16782,N_12300,N_15315);
nand U16783 (N_16783,N_14964,N_13536);
nor U16784 (N_16784,N_15014,N_14894);
and U16785 (N_16785,N_14301,N_13987);
nor U16786 (N_16786,N_15888,N_12168);
and U16787 (N_16787,N_15906,N_12753);
xor U16788 (N_16788,N_13964,N_12520);
nor U16789 (N_16789,N_13277,N_15270);
xor U16790 (N_16790,N_13669,N_14551);
nor U16791 (N_16791,N_15668,N_12873);
and U16792 (N_16792,N_13985,N_15462);
nand U16793 (N_16793,N_14492,N_12326);
xor U16794 (N_16794,N_14763,N_14917);
or U16795 (N_16795,N_14862,N_14101);
nor U16796 (N_16796,N_12878,N_13409);
xor U16797 (N_16797,N_14974,N_12953);
or U16798 (N_16798,N_14940,N_13828);
xnor U16799 (N_16799,N_13529,N_12435);
or U16800 (N_16800,N_12020,N_15496);
nand U16801 (N_16801,N_14265,N_12890);
nor U16802 (N_16802,N_13886,N_12357);
or U16803 (N_16803,N_13622,N_13946);
nand U16804 (N_16804,N_12342,N_12985);
nand U16805 (N_16805,N_15218,N_15502);
nand U16806 (N_16806,N_14146,N_14144);
xor U16807 (N_16807,N_15281,N_12549);
nor U16808 (N_16808,N_15627,N_14876);
nand U16809 (N_16809,N_14190,N_13181);
or U16810 (N_16810,N_15600,N_12701);
nand U16811 (N_16811,N_15116,N_14341);
nand U16812 (N_16812,N_15486,N_13288);
nor U16813 (N_16813,N_15002,N_14681);
xor U16814 (N_16814,N_15497,N_13496);
or U16815 (N_16815,N_15217,N_12898);
and U16816 (N_16816,N_13701,N_15344);
nor U16817 (N_16817,N_15208,N_15601);
xor U16818 (N_16818,N_13204,N_13432);
xor U16819 (N_16819,N_14385,N_13939);
nor U16820 (N_16820,N_13891,N_15892);
xnor U16821 (N_16821,N_14078,N_15419);
xnor U16822 (N_16822,N_13052,N_13069);
or U16823 (N_16823,N_13369,N_15640);
nand U16824 (N_16824,N_12058,N_12943);
nand U16825 (N_16825,N_12219,N_12687);
nand U16826 (N_16826,N_15985,N_13371);
nand U16827 (N_16827,N_12905,N_12187);
and U16828 (N_16828,N_13273,N_13420);
nor U16829 (N_16829,N_12671,N_12410);
nor U16830 (N_16830,N_13848,N_14126);
and U16831 (N_16831,N_12837,N_14490);
nor U16832 (N_16832,N_14692,N_15858);
and U16833 (N_16833,N_15952,N_13916);
xor U16834 (N_16834,N_15258,N_15659);
nand U16835 (N_16835,N_15598,N_12917);
nand U16836 (N_16836,N_12025,N_15547);
nor U16837 (N_16837,N_14414,N_14019);
or U16838 (N_16838,N_14093,N_13444);
and U16839 (N_16839,N_14452,N_12894);
and U16840 (N_16840,N_12956,N_15919);
and U16841 (N_16841,N_15160,N_15247);
or U16842 (N_16842,N_12632,N_15610);
and U16843 (N_16843,N_13700,N_13430);
and U16844 (N_16844,N_12695,N_12679);
xor U16845 (N_16845,N_14527,N_15980);
xor U16846 (N_16846,N_14836,N_12433);
and U16847 (N_16847,N_13411,N_14807);
nor U16848 (N_16848,N_15278,N_15030);
nor U16849 (N_16849,N_14878,N_13721);
xor U16850 (N_16850,N_12655,N_13417);
nand U16851 (N_16851,N_14791,N_15212);
or U16852 (N_16852,N_15678,N_13846);
and U16853 (N_16853,N_15909,N_13944);
and U16854 (N_16854,N_15829,N_14596);
and U16855 (N_16855,N_12341,N_14021);
xor U16856 (N_16856,N_15704,N_12201);
and U16857 (N_16857,N_15922,N_12049);
or U16858 (N_16858,N_12484,N_12682);
or U16859 (N_16859,N_13159,N_15120);
xnor U16860 (N_16860,N_14968,N_15752);
and U16861 (N_16861,N_14313,N_13110);
xor U16862 (N_16862,N_13012,N_15113);
nor U16863 (N_16863,N_14937,N_15396);
and U16864 (N_16864,N_15904,N_14906);
nand U16865 (N_16865,N_15577,N_15241);
and U16866 (N_16866,N_14119,N_14255);
or U16867 (N_16867,N_13796,N_12875);
and U16868 (N_16868,N_14757,N_15856);
or U16869 (N_16869,N_13249,N_13962);
nand U16870 (N_16870,N_13447,N_14783);
and U16871 (N_16871,N_15248,N_12115);
and U16872 (N_16872,N_13679,N_13123);
xnor U16873 (N_16873,N_15357,N_15694);
xnor U16874 (N_16874,N_14224,N_13384);
xor U16875 (N_16875,N_12702,N_15139);
nor U16876 (N_16876,N_13448,N_14067);
nor U16877 (N_16877,N_15378,N_13365);
or U16878 (N_16878,N_13725,N_14611);
nand U16879 (N_16879,N_14679,N_15019);
or U16880 (N_16880,N_14649,N_12711);
and U16881 (N_16881,N_15895,N_12391);
xnor U16882 (N_16882,N_15923,N_13106);
xnor U16883 (N_16883,N_15605,N_13319);
nor U16884 (N_16884,N_12952,N_15597);
and U16885 (N_16885,N_13410,N_12094);
or U16886 (N_16886,N_13966,N_13575);
nand U16887 (N_16887,N_13935,N_15054);
nand U16888 (N_16888,N_15228,N_14951);
xor U16889 (N_16889,N_14511,N_12081);
or U16890 (N_16890,N_15596,N_13094);
nor U16891 (N_16891,N_12288,N_12843);
nor U16892 (N_16892,N_14863,N_14164);
and U16893 (N_16893,N_15321,N_14522);
nor U16894 (N_16894,N_12623,N_13072);
nand U16895 (N_16895,N_15107,N_12877);
nand U16896 (N_16896,N_14418,N_12476);
nor U16897 (N_16897,N_14784,N_15355);
and U16898 (N_16898,N_14110,N_12720);
and U16899 (N_16899,N_15766,N_13062);
and U16900 (N_16900,N_12199,N_12573);
and U16901 (N_16901,N_12304,N_14953);
nand U16902 (N_16902,N_14251,N_15789);
xor U16903 (N_16903,N_15455,N_14105);
xor U16904 (N_16904,N_12615,N_15015);
xnor U16905 (N_16905,N_12646,N_15912);
and U16906 (N_16906,N_14156,N_15471);
xor U16907 (N_16907,N_15891,N_13498);
and U16908 (N_16908,N_14893,N_13710);
nor U16909 (N_16909,N_12805,N_15975);
nor U16910 (N_16910,N_14911,N_14476);
xor U16911 (N_16911,N_15200,N_12625);
xnor U16912 (N_16912,N_15062,N_12947);
and U16913 (N_16913,N_12291,N_13605);
and U16914 (N_16914,N_15528,N_12024);
nand U16915 (N_16915,N_14727,N_12507);
xor U16916 (N_16916,N_13374,N_14600);
nand U16917 (N_16917,N_15520,N_13993);
and U16918 (N_16918,N_14256,N_15548);
nor U16919 (N_16919,N_14063,N_14145);
xnor U16920 (N_16920,N_15760,N_12156);
or U16921 (N_16921,N_14837,N_14333);
and U16922 (N_16922,N_14769,N_15685);
nor U16923 (N_16923,N_13735,N_14109);
xnor U16924 (N_16924,N_15215,N_12480);
xnor U16925 (N_16925,N_12684,N_13904);
or U16926 (N_16926,N_13745,N_13736);
and U16927 (N_16927,N_13436,N_12405);
xor U16928 (N_16928,N_15485,N_14300);
xor U16929 (N_16929,N_15133,N_12299);
and U16930 (N_16930,N_15429,N_15192);
nor U16931 (N_16931,N_13023,N_14949);
and U16932 (N_16932,N_14468,N_13693);
nor U16933 (N_16933,N_15050,N_15951);
xnor U16934 (N_16934,N_13917,N_12083);
or U16935 (N_16935,N_14491,N_14819);
nor U16936 (N_16936,N_12056,N_13601);
nor U16937 (N_16937,N_12813,N_13659);
and U16938 (N_16938,N_14958,N_13284);
xor U16939 (N_16939,N_12551,N_12969);
xor U16940 (N_16940,N_14223,N_12029);
nor U16941 (N_16941,N_14057,N_15001);
nand U16942 (N_16942,N_12752,N_14206);
or U16943 (N_16943,N_12795,N_15592);
nor U16944 (N_16944,N_14755,N_13814);
nor U16945 (N_16945,N_13631,N_14138);
or U16946 (N_16946,N_12309,N_14058);
nor U16947 (N_16947,N_15447,N_12635);
nor U16948 (N_16948,N_13934,N_12330);
xor U16949 (N_16949,N_12774,N_15112);
nor U16950 (N_16950,N_15719,N_13636);
and U16951 (N_16951,N_14920,N_12818);
nor U16952 (N_16952,N_12009,N_15987);
xor U16953 (N_16953,N_13999,N_14415);
or U16954 (N_16954,N_14480,N_15161);
nand U16955 (N_16955,N_15034,N_12889);
or U16956 (N_16956,N_13942,N_14409);
nor U16957 (N_16957,N_15522,N_14413);
or U16958 (N_16958,N_15445,N_12116);
nand U16959 (N_16959,N_13102,N_14467);
and U16960 (N_16960,N_13887,N_13642);
or U16961 (N_16961,N_12397,N_15097);
or U16962 (N_16962,N_15468,N_13713);
nor U16963 (N_16963,N_14142,N_14657);
or U16964 (N_16964,N_12565,N_12050);
nor U16965 (N_16965,N_13517,N_13156);
xnor U16966 (N_16966,N_14886,N_13305);
xnor U16967 (N_16967,N_12380,N_15385);
or U16968 (N_16968,N_13211,N_12790);
nand U16969 (N_16969,N_14349,N_12003);
or U16970 (N_16970,N_14322,N_13413);
and U16971 (N_16971,N_12387,N_13009);
or U16972 (N_16972,N_13003,N_15253);
xnor U16973 (N_16973,N_13290,N_14562);
or U16974 (N_16974,N_12617,N_13624);
or U16975 (N_16975,N_13422,N_14460);
xnor U16976 (N_16976,N_14344,N_13714);
and U16977 (N_16977,N_13595,N_14778);
and U16978 (N_16978,N_15916,N_13815);
nor U16979 (N_16979,N_15586,N_12278);
nor U16980 (N_16980,N_14957,N_12674);
xor U16981 (N_16981,N_14249,N_13504);
or U16982 (N_16982,N_13240,N_12348);
and U16983 (N_16983,N_12471,N_12102);
or U16984 (N_16984,N_13427,N_14768);
xor U16985 (N_16985,N_15261,N_15558);
and U16986 (N_16986,N_14613,N_14888);
nor U16987 (N_16987,N_15648,N_12396);
xor U16988 (N_16988,N_15272,N_13928);
nand U16989 (N_16989,N_14212,N_13514);
and U16990 (N_16990,N_12355,N_12314);
nor U16991 (N_16991,N_14153,N_15038);
xnor U16992 (N_16992,N_13482,N_13799);
or U16993 (N_16993,N_15967,N_12360);
nor U16994 (N_16994,N_15379,N_12121);
nor U16995 (N_16995,N_12858,N_13884);
and U16996 (N_16996,N_15683,N_14694);
and U16997 (N_16997,N_15774,N_13385);
or U16998 (N_16998,N_13592,N_14711);
and U16999 (N_16999,N_13233,N_12152);
nand U17000 (N_17000,N_15025,N_14481);
or U17001 (N_17001,N_14844,N_13560);
or U17002 (N_17002,N_14915,N_15852);
and U17003 (N_17003,N_15283,N_13468);
xnor U17004 (N_17004,N_15184,N_13664);
or U17005 (N_17005,N_14767,N_13398);
nand U17006 (N_17006,N_13524,N_12803);
xor U17007 (N_17007,N_15697,N_12807);
nor U17008 (N_17008,N_15314,N_15590);
and U17009 (N_17009,N_15938,N_13909);
nor U17010 (N_17010,N_12052,N_13435);
xnor U17011 (N_17011,N_15220,N_12240);
xor U17012 (N_17012,N_15110,N_12203);
nand U17013 (N_17013,N_15655,N_15403);
nor U17014 (N_17014,N_13926,N_14760);
and U17015 (N_17015,N_12236,N_13963);
nand U17016 (N_17016,N_13822,N_14438);
xnor U17017 (N_17017,N_13875,N_12349);
and U17018 (N_17018,N_14963,N_15211);
or U17019 (N_17019,N_13509,N_12287);
xnor U17020 (N_17020,N_14306,N_14209);
nor U17021 (N_17021,N_15942,N_13085);
and U17022 (N_17022,N_15823,N_15550);
and U17023 (N_17023,N_12950,N_12416);
xnor U17024 (N_17024,N_12743,N_14450);
xor U17025 (N_17025,N_12651,N_13614);
or U17026 (N_17026,N_12958,N_12327);
nor U17027 (N_17027,N_13165,N_13086);
and U17028 (N_17028,N_14307,N_13724);
nand U17029 (N_17029,N_12527,N_14535);
and U17030 (N_17030,N_13268,N_15607);
or U17031 (N_17031,N_12255,N_13487);
xor U17032 (N_17032,N_15783,N_15341);
nor U17033 (N_17033,N_14388,N_13698);
and U17034 (N_17034,N_13230,N_14091);
xor U17035 (N_17035,N_15222,N_14193);
nor U17036 (N_17036,N_12245,N_12442);
nand U17037 (N_17037,N_13343,N_12728);
nor U17038 (N_17038,N_13583,N_14518);
nand U17039 (N_17039,N_14321,N_14879);
nand U17040 (N_17040,N_12740,N_15374);
nor U17041 (N_17041,N_13511,N_14956);
or U17042 (N_17042,N_13315,N_13768);
xor U17043 (N_17043,N_15936,N_12379);
nand U17044 (N_17044,N_12893,N_12196);
or U17045 (N_17045,N_12641,N_15417);
and U17046 (N_17046,N_12388,N_13465);
or U17047 (N_17047,N_14889,N_12057);
and U17048 (N_17048,N_15964,N_14568);
nor U17049 (N_17049,N_12430,N_13952);
nand U17050 (N_17050,N_12335,N_14088);
xor U17051 (N_17051,N_15997,N_13166);
xnor U17052 (N_17052,N_13731,N_13270);
or U17053 (N_17053,N_13491,N_14039);
nor U17054 (N_17054,N_12585,N_13861);
nor U17055 (N_17055,N_12661,N_15495);
xnor U17056 (N_17056,N_15734,N_12972);
nor U17057 (N_17057,N_14211,N_15418);
or U17058 (N_17058,N_12971,N_14334);
nand U17059 (N_17059,N_15013,N_14873);
xnor U17060 (N_17060,N_14887,N_15087);
nand U17061 (N_17061,N_15931,N_14719);
or U17062 (N_17062,N_14451,N_13317);
nand U17063 (N_17063,N_13570,N_14561);
nor U17064 (N_17064,N_14645,N_14074);
nor U17065 (N_17065,N_14398,N_14495);
xnor U17066 (N_17066,N_13367,N_12046);
xor U17067 (N_17067,N_15083,N_14455);
nand U17068 (N_17068,N_12426,N_12564);
or U17069 (N_17069,N_13161,N_13804);
or U17070 (N_17070,N_13598,N_14185);
or U17071 (N_17071,N_14010,N_12177);
or U17072 (N_17072,N_13366,N_12831);
or U17073 (N_17073,N_12451,N_14326);
nand U17074 (N_17074,N_14317,N_12093);
nor U17075 (N_17075,N_13675,N_13271);
nor U17076 (N_17076,N_13901,N_13785);
nor U17077 (N_17077,N_13890,N_15213);
nand U17078 (N_17078,N_14728,N_13051);
and U17079 (N_17079,N_15224,N_14766);
or U17080 (N_17080,N_13286,N_15099);
xor U17081 (N_17081,N_12109,N_13001);
nand U17082 (N_17082,N_12676,N_13274);
and U17083 (N_17083,N_13863,N_12189);
xnor U17084 (N_17084,N_12228,N_15153);
and U17085 (N_17085,N_13349,N_13869);
or U17086 (N_17086,N_13769,N_14082);
nor U17087 (N_17087,N_15508,N_13157);
nand U17088 (N_17088,N_14779,N_15182);
nor U17089 (N_17089,N_14542,N_12373);
xor U17090 (N_17090,N_13292,N_13189);
nand U17091 (N_17091,N_12281,N_12271);
nor U17092 (N_17092,N_14309,N_14118);
nand U17093 (N_17093,N_15625,N_12631);
or U17094 (N_17094,N_15406,N_13618);
or U17095 (N_17095,N_15748,N_13146);
xnor U17096 (N_17096,N_13294,N_14743);
xor U17097 (N_17097,N_15460,N_14831);
or U17098 (N_17098,N_13797,N_13559);
or U17099 (N_17099,N_12016,N_13036);
xnor U17100 (N_17100,N_14258,N_14725);
nor U17101 (N_17101,N_14756,N_14633);
nand U17102 (N_17102,N_15427,N_12994);
xnor U17103 (N_17103,N_13518,N_13175);
nand U17104 (N_17104,N_14263,N_13948);
xor U17105 (N_17105,N_15343,N_13927);
and U17106 (N_17106,N_15747,N_15687);
and U17107 (N_17107,N_15995,N_14834);
xor U17108 (N_17108,N_13795,N_14405);
nor U17109 (N_17109,N_13245,N_12689);
nor U17110 (N_17110,N_13050,N_14332);
or U17111 (N_17111,N_12294,N_14399);
xor U17112 (N_17112,N_13047,N_13571);
nor U17113 (N_17113,N_13429,N_12055);
nor U17114 (N_17114,N_14136,N_14342);
and U17115 (N_17115,N_13478,N_13719);
nand U17116 (N_17116,N_12511,N_14454);
nand U17117 (N_17117,N_14384,N_15433);
xnor U17118 (N_17118,N_14574,N_13757);
xor U17119 (N_17119,N_13068,N_12145);
nand U17120 (N_17120,N_15549,N_14751);
nor U17121 (N_17121,N_15368,N_13991);
and U17122 (N_17122,N_13275,N_14726);
and U17123 (N_17123,N_13143,N_13857);
or U17124 (N_17124,N_14022,N_12098);
and U17125 (N_17125,N_12110,N_14319);
nor U17126 (N_17126,N_12285,N_12073);
or U17127 (N_17127,N_14395,N_15841);
xnor U17128 (N_17128,N_15673,N_15199);
or U17129 (N_17129,N_12154,N_14011);
xnor U17130 (N_17130,N_15715,N_14703);
or U17131 (N_17131,N_15667,N_15289);
xor U17132 (N_17132,N_13495,N_12415);
and U17133 (N_17133,N_13590,N_14419);
or U17134 (N_17134,N_12976,N_12334);
xor U17135 (N_17135,N_14962,N_12862);
or U17136 (N_17136,N_15624,N_14640);
xnor U17137 (N_17137,N_13507,N_15804);
and U17138 (N_17138,N_12630,N_15162);
and U17139 (N_17139,N_12566,N_12369);
nand U17140 (N_17140,N_12928,N_13760);
nor U17141 (N_17141,N_14824,N_14084);
and U17142 (N_17142,N_13809,N_13064);
nand U17143 (N_17143,N_12993,N_14583);
or U17144 (N_17144,N_13355,N_13685);
and U17145 (N_17145,N_13646,N_13449);
and U17146 (N_17146,N_14416,N_12892);
nand U17147 (N_17147,N_15943,N_13607);
or U17148 (N_17148,N_14141,N_15262);
xnor U17149 (N_17149,N_12400,N_14710);
nor U17150 (N_17150,N_14123,N_12407);
nand U17151 (N_17151,N_15589,N_12277);
or U17152 (N_17152,N_14277,N_12533);
nor U17153 (N_17153,N_15611,N_15047);
and U17154 (N_17154,N_13697,N_13716);
and U17155 (N_17155,N_13416,N_15865);
nor U17156 (N_17156,N_15677,N_13224);
or U17157 (N_17157,N_13403,N_14045);
and U17158 (N_17158,N_13210,N_14934);
nor U17159 (N_17159,N_14902,N_12179);
nand U17160 (N_17160,N_15886,N_12567);
nor U17161 (N_17161,N_13885,N_12428);
nand U17162 (N_17162,N_12978,N_12714);
or U17163 (N_17163,N_13541,N_13065);
nand U17164 (N_17164,N_14771,N_15556);
and U17165 (N_17165,N_13965,N_14742);
or U17166 (N_17166,N_12319,N_13666);
xnor U17167 (N_17167,N_14533,N_15407);
or U17168 (N_17168,N_14090,N_12607);
nor U17169 (N_17169,N_13596,N_12621);
and U17170 (N_17170,N_12645,N_13100);
xor U17171 (N_17171,N_13988,N_14581);
xnor U17172 (N_17172,N_15239,N_13061);
and U17173 (N_17173,N_13717,N_12759);
xor U17174 (N_17174,N_15244,N_12763);
or U17175 (N_17175,N_12394,N_15431);
nor U17176 (N_17176,N_15712,N_12137);
nor U17177 (N_17177,N_13577,N_13951);
nor U17178 (N_17178,N_15777,N_12138);
and U17179 (N_17179,N_12606,N_13362);
or U17180 (N_17180,N_14200,N_15998);
and U17181 (N_17181,N_13821,N_13155);
xnor U17182 (N_17182,N_15838,N_15529);
nand U17183 (N_17183,N_12362,N_15898);
nand U17184 (N_17184,N_14579,N_15279);
nand U17185 (N_17185,N_15072,N_12596);
nand U17186 (N_17186,N_15686,N_14392);
nand U17187 (N_17187,N_15389,N_15896);
or U17188 (N_17188,N_13056,N_14502);
nor U17189 (N_17189,N_14872,N_14426);
and U17190 (N_17190,N_14922,N_13565);
xnor U17191 (N_17191,N_13198,N_12949);
and U17192 (N_17192,N_14178,N_14595);
or U17193 (N_17193,N_14380,N_13031);
nor U17194 (N_17194,N_12524,N_13548);
or U17195 (N_17195,N_14924,N_14352);
or U17196 (N_17196,N_14638,N_15792);
and U17197 (N_17197,N_14587,N_15953);
and U17198 (N_17198,N_14038,N_14100);
and U17199 (N_17199,N_13516,N_15675);
nor U17200 (N_17200,N_15234,N_12828);
xor U17201 (N_17201,N_14656,N_13969);
and U17202 (N_17202,N_14619,N_13291);
nor U17203 (N_17203,N_13753,N_14314);
nand U17204 (N_17204,N_13637,N_14356);
nor U17205 (N_17205,N_13045,N_12142);
nand U17206 (N_17206,N_14250,N_13455);
or U17207 (N_17207,N_12293,N_12191);
or U17208 (N_17208,N_13450,N_13654);
and U17209 (N_17209,N_14623,N_15308);
and U17210 (N_17210,N_14943,N_14445);
and U17211 (N_17211,N_15806,N_12542);
or U17212 (N_17212,N_12149,N_12586);
or U17213 (N_17213,N_13671,N_14806);
or U17214 (N_17214,N_12577,N_15479);
and U17215 (N_17215,N_15079,N_13026);
or U17216 (N_17216,N_12144,N_13741);
nand U17217 (N_17217,N_15255,N_14046);
nor U17218 (N_17218,N_14983,N_15189);
nand U17219 (N_17219,N_12809,N_13169);
xnor U17220 (N_17220,N_15826,N_14548);
xor U17221 (N_17221,N_14373,N_12692);
xor U17222 (N_17222,N_15753,N_13002);
or U17223 (N_17223,N_15963,N_15643);
or U17224 (N_17224,N_12575,N_14869);
or U17225 (N_17225,N_14785,N_14818);
or U17226 (N_17226,N_15561,N_15630);
xor U17227 (N_17227,N_12151,N_15149);
xor U17228 (N_17228,N_14441,N_15541);
or U17229 (N_17229,N_14660,N_14429);
nor U17230 (N_17230,N_14781,N_13550);
or U17231 (N_17231,N_14112,N_12820);
nor U17232 (N_17232,N_14081,N_12424);
or U17233 (N_17233,N_12260,N_13610);
nor U17234 (N_17234,N_12377,N_14279);
and U17235 (N_17235,N_12694,N_14588);
nor U17236 (N_17236,N_13220,N_13115);
or U17237 (N_17237,N_12354,N_13899);
and U17238 (N_17238,N_12761,N_12561);
and U17239 (N_17239,N_12731,N_14357);
nand U17240 (N_17240,N_13221,N_15408);
xor U17241 (N_17241,N_15515,N_15331);
nor U17242 (N_17242,N_15480,N_14089);
nor U17243 (N_17243,N_12854,N_14462);
nor U17244 (N_17244,N_14696,N_13392);
and U17245 (N_17245,N_15795,N_12896);
and U17246 (N_17246,N_13201,N_15323);
and U17247 (N_17247,N_12344,N_12167);
nand U17248 (N_17248,N_14466,N_12693);
and U17249 (N_17249,N_15669,N_13049);
and U17250 (N_17250,N_12834,N_15237);
nand U17251 (N_17251,N_12028,N_14155);
xor U17252 (N_17252,N_13350,N_13265);
or U17253 (N_17253,N_13162,N_14242);
xor U17254 (N_17254,N_13152,N_12560);
nor U17255 (N_17255,N_12328,N_13108);
xnor U17256 (N_17256,N_13229,N_15635);
xor U17257 (N_17257,N_14762,N_13789);
and U17258 (N_17258,N_12665,N_14833);
and U17259 (N_17259,N_14504,N_15350);
and U17260 (N_17260,N_14747,N_15227);
or U17261 (N_17261,N_12656,N_15609);
nor U17262 (N_17262,N_12030,N_12842);
xnor U17263 (N_17263,N_13663,N_14569);
xor U17264 (N_17264,N_14871,N_13132);
and U17265 (N_17265,N_13782,N_13357);
or U17266 (N_17266,N_14503,N_13379);
or U17267 (N_17267,N_14839,N_15564);
nor U17268 (N_17268,N_14389,N_12518);
nand U17269 (N_17269,N_13973,N_14571);
and U17270 (N_17270,N_13833,N_13902);
xor U17271 (N_17271,N_12989,N_13467);
and U17272 (N_17272,N_13515,N_14549);
and U17273 (N_17273,N_12365,N_14012);
nor U17274 (N_17274,N_14086,N_12733);
and U17275 (N_17275,N_13456,N_12614);
or U17276 (N_17276,N_12311,N_15992);
xnor U17277 (N_17277,N_15441,N_13914);
nand U17278 (N_17278,N_14714,N_13882);
xnor U17279 (N_17279,N_13766,N_12885);
nand U17280 (N_17280,N_13998,N_14544);
or U17281 (N_17281,N_15682,N_14816);
nand U17282 (N_17282,N_14984,N_15307);
and U17283 (N_17283,N_13883,N_12800);
xor U17284 (N_17284,N_14486,N_13981);
and U17285 (N_17285,N_15435,N_15041);
xnor U17286 (N_17286,N_12838,N_12545);
xnor U17287 (N_17287,N_14457,N_14685);
xnor U17288 (N_17288,N_12552,N_15335);
or U17289 (N_17289,N_15977,N_13572);
nor U17290 (N_17290,N_12019,N_14183);
and U17291 (N_17291,N_13532,N_15679);
xnor U17292 (N_17292,N_14970,N_14967);
xnor U17293 (N_17293,N_14775,N_15879);
or U17294 (N_17294,N_13702,N_13093);
or U17295 (N_17295,N_15817,N_12704);
and U17296 (N_17296,N_13199,N_15146);
and U17297 (N_17297,N_14191,N_13845);
nor U17298 (N_17298,N_14827,N_13177);
and U17299 (N_17299,N_12516,N_14950);
and U17300 (N_17300,N_13932,N_12267);
or U17301 (N_17301,N_12780,N_15156);
and U17302 (N_17302,N_15518,N_14030);
xor U17303 (N_17303,N_13415,N_15140);
or U17304 (N_17304,N_12249,N_14260);
xnor U17305 (N_17305,N_14900,N_13127);
and U17306 (N_17306,N_13970,N_13440);
xnor U17307 (N_17307,N_12232,N_12868);
xnor U17308 (N_17308,N_12992,N_14387);
and U17309 (N_17309,N_15620,N_12447);
xor U17310 (N_17310,N_13978,N_14896);
and U17311 (N_17311,N_13453,N_14315);
or U17312 (N_17312,N_12022,N_13263);
nor U17313 (N_17313,N_13986,N_13081);
nand U17314 (N_17314,N_14811,N_14449);
or U17315 (N_17315,N_14812,N_12707);
and U17316 (N_17316,N_14720,N_13151);
and U17317 (N_17317,N_13734,N_15045);
nand U17318 (N_17318,N_13625,N_15822);
nor U17319 (N_17319,N_14281,N_14487);
or U17320 (N_17320,N_12915,N_15304);
nand U17321 (N_17321,N_14986,N_12935);
xor U17322 (N_17322,N_15360,N_15075);
nand U17323 (N_17323,N_15458,N_13526);
xor U17324 (N_17324,N_14041,N_12624);
and U17325 (N_17325,N_15757,N_12649);
nand U17326 (N_17326,N_13375,N_12653);
nor U17327 (N_17327,N_14396,N_14599);
xor U17328 (N_17328,N_12589,N_14954);
or U17329 (N_17329,N_15925,N_12092);
xor U17330 (N_17330,N_12913,N_14753);
and U17331 (N_17331,N_12166,N_15238);
or U17332 (N_17332,N_13038,N_14608);
or U17333 (N_17333,N_13452,N_14947);
and U17334 (N_17334,N_12134,N_12275);
and U17335 (N_17335,N_15310,N_12427);
xnor U17336 (N_17336,N_12207,N_14699);
and U17337 (N_17337,N_13673,N_12963);
and U17338 (N_17338,N_12012,N_14972);
and U17339 (N_17339,N_14606,N_15401);
xnor U17340 (N_17340,N_13461,N_14555);
nor U17341 (N_17341,N_14199,N_13316);
and U17342 (N_17342,N_13968,N_12936);
and U17343 (N_17343,N_12569,N_13556);
nor U17344 (N_17344,N_12258,N_12234);
or U17345 (N_17345,N_14381,N_14440);
or U17346 (N_17346,N_14987,N_14288);
nand U17347 (N_17347,N_14628,N_12857);
nor U17348 (N_17348,N_14680,N_14266);
or U17349 (N_17349,N_12845,N_12475);
nor U17350 (N_17350,N_15482,N_12186);
and U17351 (N_17351,N_13207,N_12660);
or U17352 (N_17352,N_15941,N_13479);
or U17353 (N_17353,N_15049,N_14732);
and U17354 (N_17354,N_13806,N_13635);
and U17355 (N_17355,N_15286,N_15828);
nand U17356 (N_17356,N_14472,N_14018);
nand U17357 (N_17357,N_14161,N_13667);
nand U17358 (N_17358,N_13599,N_14408);
nor U17359 (N_17359,N_14517,N_12132);
xnor U17360 (N_17360,N_14575,N_15861);
nand U17361 (N_17361,N_13007,N_13656);
or U17362 (N_17362,N_15375,N_14485);
xnor U17363 (N_17363,N_15632,N_15999);
or U17364 (N_17364,N_15989,N_13202);
nor U17365 (N_17365,N_15889,N_13125);
nor U17366 (N_17366,N_13356,N_13232);
and U17367 (N_17367,N_14848,N_15044);
and U17368 (N_17368,N_12261,N_13243);
or U17369 (N_17369,N_12672,N_13466);
xnor U17370 (N_17370,N_15991,N_15070);
nand U17371 (N_17371,N_13219,N_15580);
nand U17372 (N_17372,N_12079,N_13776);
nand U17373 (N_17373,N_12980,N_15506);
nor U17374 (N_17374,N_15267,N_12909);
xnor U17375 (N_17375,N_14822,N_15207);
nor U17376 (N_17376,N_14704,N_12498);
nand U17377 (N_17377,N_14616,N_12455);
and U17378 (N_17378,N_15111,N_15007);
nand U17379 (N_17379,N_14738,N_15727);
nor U17380 (N_17380,N_12460,N_15948);
xnor U17381 (N_17381,N_14969,N_15369);
nand U17382 (N_17382,N_13258,N_13280);
xor U17383 (N_17383,N_12538,N_14804);
nor U17384 (N_17384,N_12248,N_12238);
nand U17385 (N_17385,N_13684,N_15134);
xnor U17386 (N_17386,N_14774,N_15512);
and U17387 (N_17387,N_14715,N_12481);
nor U17388 (N_17388,N_15785,N_13129);
and U17389 (N_17389,N_15256,N_14168);
nand U17390 (N_17390,N_15472,N_14005);
or U17391 (N_17391,N_12305,N_14004);
or U17392 (N_17392,N_13632,N_13113);
nand U17393 (N_17393,N_12216,N_13594);
nor U17394 (N_17394,N_15095,N_15570);
nand U17395 (N_17395,N_14204,N_13979);
or U17396 (N_17396,N_15739,N_12032);
nand U17397 (N_17397,N_12922,N_13501);
and U17398 (N_17398,N_12539,N_14740);
xor U17399 (N_17399,N_15578,N_13195);
or U17400 (N_17400,N_14192,N_15434);
and U17401 (N_17401,N_12755,N_14697);
nor U17402 (N_17402,N_14053,N_15003);
xnor U17403 (N_17403,N_15356,N_12937);
or U17404 (N_17404,N_14752,N_12853);
xor U17405 (N_17405,N_12951,N_13279);
xor U17406 (N_17406,N_13034,N_12712);
nand U17407 (N_17407,N_12005,N_12530);
and U17408 (N_17408,N_13683,N_15873);
xor U17409 (N_17409,N_15651,N_13404);
and U17410 (N_17410,N_13122,N_13425);
xor U17411 (N_17411,N_14629,N_14371);
and U17412 (N_17412,N_14033,N_13377);
nor U17413 (N_17413,N_13906,N_13523);
or U17414 (N_17414,N_15345,N_14538);
nand U17415 (N_17415,N_14000,N_12525);
nand U17416 (N_17416,N_14528,N_14761);
xnor U17417 (N_17417,N_12715,N_15010);
or U17418 (N_17418,N_15490,N_14453);
or U17419 (N_17419,N_14173,N_12662);
or U17420 (N_17420,N_13310,N_13345);
or U17421 (N_17421,N_15093,N_14303);
xnor U17422 (N_17422,N_13545,N_15405);
xnor U17423 (N_17423,N_15583,N_13639);
or U17424 (N_17424,N_12250,N_12015);
xnor U17425 (N_17425,N_14597,N_14377);
nand U17426 (N_17426,N_12926,N_12087);
nor U17427 (N_17427,N_13396,N_13163);
nor U17428 (N_17428,N_12265,N_15203);
xor U17429 (N_17429,N_15131,N_14496);
nand U17430 (N_17430,N_14724,N_12633);
xnor U17431 (N_17431,N_15380,N_14423);
and U17432 (N_17432,N_12284,N_13182);
nand U17433 (N_17433,N_12514,N_15893);
nand U17434 (N_17434,N_13562,N_15390);
nand U17435 (N_17435,N_15483,N_14410);
or U17436 (N_17436,N_12128,N_15488);
xor U17437 (N_17437,N_13747,N_14948);
and U17438 (N_17438,N_13492,N_15141);
and U17439 (N_17439,N_12295,N_13801);
or U17440 (N_17440,N_12043,N_15106);
nand U17441 (N_17441,N_12064,N_13099);
or U17442 (N_17442,N_13459,N_15618);
nor U17443 (N_17443,N_12339,N_15305);
nor U17444 (N_17444,N_14282,N_15260);
and U17445 (N_17445,N_14220,N_14976);
nand U17446 (N_17446,N_15993,N_14636);
and U17447 (N_17447,N_15397,N_13073);
and U17448 (N_17448,N_12312,N_13619);
xnor U17449 (N_17449,N_14499,N_13348);
nor U17450 (N_17450,N_14576,N_13824);
xor U17451 (N_17451,N_14087,N_12832);
nor U17452 (N_17452,N_15042,N_12775);
xor U17453 (N_17453,N_15961,N_14501);
and U17454 (N_17454,N_14814,N_12835);
or U17455 (N_17455,N_15954,N_15303);
xor U17456 (N_17456,N_13399,N_15866);
or U17457 (N_17457,N_14841,N_15425);
and U17458 (N_17458,N_15232,N_14698);
and U17459 (N_17459,N_15956,N_14620);
xor U17460 (N_17460,N_14443,N_15071);
nor U17461 (N_17461,N_12268,N_12316);
xor U17462 (N_17462,N_12824,N_13361);
nand U17463 (N_17463,N_15767,N_12479);
or U17464 (N_17464,N_13615,N_14122);
xor U17465 (N_17465,N_15557,N_12942);
nor U17466 (N_17466,N_13672,N_14602);
xnor U17467 (N_17467,N_13873,N_14582);
nand U17468 (N_17468,N_15871,N_15271);
nor U17469 (N_17469,N_12420,N_14541);
and U17470 (N_17470,N_15722,N_12496);
and U17471 (N_17471,N_15328,N_12986);
and U17472 (N_17472,N_12691,N_14043);
xor U17473 (N_17473,N_15691,N_14217);
or U17474 (N_17474,N_15926,N_12183);
or U17475 (N_17475,N_13185,N_12143);
nand U17476 (N_17476,N_15129,N_13739);
and U17477 (N_17477,N_14431,N_12587);
nand U17478 (N_17478,N_14154,N_13457);
and U17479 (N_17479,N_13329,N_12225);
xor U17480 (N_17480,N_13864,N_12930);
xnor U17481 (N_17481,N_13749,N_12772);
nand U17482 (N_17482,N_14960,N_15762);
nand U17483 (N_17483,N_14789,N_12218);
and U17484 (N_17484,N_12781,N_12815);
nand U17485 (N_17485,N_14184,N_12830);
xor U17486 (N_17486,N_12041,N_15910);
nor U17487 (N_17487,N_13011,N_13744);
or U17488 (N_17488,N_12091,N_13692);
or U17489 (N_17489,N_12789,N_14881);
nand U17490 (N_17490,N_15519,N_14077);
or U17491 (N_17491,N_15988,N_15452);
and U17492 (N_17492,N_15381,N_14961);
or U17493 (N_17493,N_13812,N_15254);
and U17494 (N_17494,N_15264,N_14955);
and U17495 (N_17495,N_14805,N_14563);
or U17496 (N_17496,N_14051,N_12211);
xnor U17497 (N_17497,N_12921,N_15652);
or U17498 (N_17498,N_12663,N_14592);
and U17499 (N_17499,N_15525,N_13018);
nor U17500 (N_17500,N_14298,N_13876);
xor U17501 (N_17501,N_12503,N_12060);
xor U17502 (N_17502,N_14170,N_12946);
nor U17503 (N_17503,N_13989,N_12204);
or U17504 (N_17504,N_12547,N_14722);
nand U17505 (N_17505,N_15018,N_14653);
or U17506 (N_17506,N_13889,N_12482);
nand U17507 (N_17507,N_14746,N_15231);
and U17508 (N_17508,N_14718,N_13645);
nand U17509 (N_17509,N_15612,N_14097);
or U17510 (N_17510,N_15453,N_15494);
xor U17511 (N_17511,N_14589,N_14148);
nand U17512 (N_17512,N_13756,N_15249);
nor U17513 (N_17513,N_12571,N_13330);
nor U17514 (N_17514,N_12576,N_14938);
and U17515 (N_17515,N_13406,N_12368);
or U17516 (N_17516,N_12706,N_15921);
and U17517 (N_17517,N_12244,N_15186);
xor U17518 (N_17518,N_13484,N_14152);
xor U17519 (N_17519,N_14520,N_12738);
and U17520 (N_17520,N_13792,N_13424);
xor U17521 (N_17521,N_14289,N_13438);
and U17522 (N_17522,N_15614,N_12735);
nor U17523 (N_17523,N_15899,N_13967);
xnor U17524 (N_17524,N_13326,N_12095);
xnor U17525 (N_17525,N_14677,N_15317);
and U17526 (N_17526,N_12724,N_15602);
xnor U17527 (N_17527,N_15974,N_14684);
nand U17528 (N_17528,N_14654,N_13443);
and U17529 (N_17529,N_14096,N_12434);
and U17530 (N_17530,N_13130,N_12042);
or U17531 (N_17531,N_15511,N_15960);
nand U17532 (N_17532,N_15821,N_15159);
nand U17533 (N_17533,N_13617,N_14702);
nand U17534 (N_17534,N_13868,N_15067);
nand U17535 (N_17535,N_12398,N_15688);
or U17536 (N_17536,N_12283,N_15201);
nand U17537 (N_17537,N_14864,N_12557);
nand U17538 (N_17538,N_14362,N_15729);
xor U17539 (N_17539,N_14815,N_12402);
nand U17540 (N_17540,N_14274,N_15183);
nor U17541 (N_17541,N_12062,N_12938);
and U17542 (N_17542,N_12650,N_13359);
nor U17543 (N_17543,N_15820,N_14594);
and U17544 (N_17544,N_14166,N_12902);
nand U17545 (N_17545,N_12173,N_13083);
nor U17546 (N_17546,N_15466,N_15645);
nand U17547 (N_17547,N_14780,N_13017);
xnor U17548 (N_17548,N_13388,N_12161);
nand U17549 (N_17549,N_14006,N_14513);
or U17550 (N_17550,N_12544,N_12160);
and U17551 (N_17551,N_14062,N_13296);
and U17552 (N_17552,N_14302,N_12068);
xor U17553 (N_17553,N_13593,N_12588);
and U17554 (N_17554,N_13900,N_13850);
or U17555 (N_17555,N_14040,N_12243);
nor U17556 (N_17556,N_14689,N_14572);
and U17557 (N_17557,N_15791,N_12100);
xnor U17558 (N_17558,N_15650,N_12217);
xnor U17559 (N_17559,N_13867,N_15060);
nor U17560 (N_17560,N_12450,N_14498);
and U17561 (N_17561,N_15475,N_12465);
or U17562 (N_17562,N_13251,N_12376);
nand U17563 (N_17563,N_13621,N_14231);
nor U17564 (N_17564,N_13627,N_15432);
or U17565 (N_17565,N_13688,N_13519);
nand U17566 (N_17566,N_12385,N_14999);
or U17567 (N_17567,N_15198,N_12366);
xnor U17568 (N_17568,N_14312,N_14658);
and U17569 (N_17569,N_14305,N_14709);
xor U17570 (N_17570,N_15604,N_14379);
and U17571 (N_17571,N_15132,N_15516);
and U17572 (N_17572,N_14564,N_14272);
nor U17573 (N_17573,N_13919,N_15945);
nor U17574 (N_17574,N_14627,N_14286);
nor U17575 (N_17575,N_13183,N_13363);
or U17576 (N_17576,N_12683,N_13694);
nor U17577 (N_17577,N_12741,N_12210);
or U17578 (N_17578,N_12425,N_15818);
and U17579 (N_17579,N_15365,N_13584);
xnor U17580 (N_17580,N_14439,N_14695);
xnor U17581 (N_17581,N_14795,N_13746);
nand U17582 (N_17582,N_12776,N_13929);
or U17583 (N_17583,N_15934,N_13613);
or U17584 (N_17584,N_14992,N_13075);
nand U17585 (N_17585,N_14942,N_13180);
nor U17586 (N_17586,N_15410,N_15978);
xnor U17587 (N_17587,N_13711,N_12170);
nand U17588 (N_17588,N_14509,N_13823);
or U17589 (N_17589,N_15621,N_14397);
or U17590 (N_17590,N_15188,N_13923);
nand U17591 (N_17591,N_15351,N_15005);
and U17592 (N_17592,N_12598,N_12747);
nor U17593 (N_17593,N_13651,N_12103);
nand U17594 (N_17594,N_12760,N_15968);
nor U17595 (N_17595,N_14996,N_12669);
or U17596 (N_17596,N_15037,N_12618);
xor U17597 (N_17597,N_12371,N_14741);
or U17598 (N_17598,N_14573,N_12340);
nor U17599 (N_17599,N_14106,N_13720);
nand U17600 (N_17600,N_12770,N_14857);
and U17601 (N_17601,N_14489,N_12331);
and U17602 (N_17602,N_12884,N_14099);
xnor U17603 (N_17603,N_15832,N_15918);
or U17604 (N_17604,N_12907,N_14207);
and U17605 (N_17605,N_12816,N_12611);
nand U17606 (N_17606,N_12864,N_13259);
and U17607 (N_17607,N_12771,N_14060);
nor U17608 (N_17608,N_12670,N_12811);
and U17609 (N_17609,N_15484,N_15566);
nand U17610 (N_17610,N_15245,N_12534);
and U17611 (N_17611,N_14376,N_14765);
nand U17612 (N_17612,N_15012,N_12887);
nor U17613 (N_17613,N_15769,N_14598);
xnor U17614 (N_17614,N_12169,N_12443);
nor U17615 (N_17615,N_15702,N_12233);
or U17616 (N_17616,N_14823,N_13318);
nand U17617 (N_17617,N_15976,N_13649);
and U17618 (N_17618,N_13325,N_15689);
and U17619 (N_17619,N_15168,N_15064);
nor U17620 (N_17620,N_12076,N_15897);
nand U17621 (N_17621,N_15572,N_15122);
nor U17622 (N_17622,N_12206,N_15057);
nor U17623 (N_17623,N_15409,N_13225);
nor U17624 (N_17624,N_14432,N_12757);
and U17625 (N_17625,N_12920,N_13412);
nand U17626 (N_17626,N_15221,N_12034);
nand U17627 (N_17627,N_15890,N_12933);
and U17628 (N_17628,N_15474,N_12125);
nor U17629 (N_17629,N_13451,N_14064);
xnor U17630 (N_17630,N_12998,N_13743);
nand U17631 (N_17631,N_14181,N_15613);
and U17632 (N_17632,N_15454,N_12997);
and U17633 (N_17633,N_12224,N_12675);
or U17634 (N_17634,N_15399,N_14749);
nand U17635 (N_17635,N_14799,N_13505);
and U17636 (N_17636,N_15306,N_15894);
nor U17637 (N_17637,N_14257,N_14268);
nand U17638 (N_17638,N_12292,N_14366);
nand U17639 (N_17639,N_13053,N_15546);
and U17640 (N_17640,N_12799,N_15124);
nor U17641 (N_17641,N_13144,N_13826);
nor U17642 (N_17642,N_15860,N_14686);
nand U17643 (N_17643,N_14243,N_14248);
nand U17644 (N_17644,N_13186,N_13039);
nor U17645 (N_17645,N_14786,N_12452);
or U17646 (N_17646,N_14615,N_12021);
and U17647 (N_17647,N_12535,N_14310);
nor U17648 (N_17648,N_14324,N_15069);
or U17649 (N_17649,N_13657,N_13431);
nor U17650 (N_17650,N_13276,N_12742);
or U17651 (N_17651,N_13278,N_12698);
nand U17652 (N_17652,N_13197,N_14359);
or U17653 (N_17653,N_15181,N_12668);
and U17654 (N_17654,N_13752,N_13442);
nand U17655 (N_17655,N_13878,N_13153);
and U17656 (N_17656,N_14147,N_14318);
xnor U17657 (N_17657,N_15214,N_12903);
xnor U17658 (N_17658,N_13918,N_15575);
and U17659 (N_17659,N_12600,N_12472);
nand U17660 (N_17660,N_15758,N_15567);
nor U17661 (N_17661,N_13010,N_12266);
and U17662 (N_17662,N_12082,N_13342);
xnor U17663 (N_17663,N_14530,N_14966);
and U17664 (N_17664,N_14269,N_14826);
nor U17665 (N_17665,N_15720,N_15416);
nand U17666 (N_17666,N_12347,N_15469);
or U17667 (N_17667,N_15835,N_15035);
or U17668 (N_17668,N_13041,N_15180);
and U17669 (N_17669,N_14758,N_14803);
or U17670 (N_17670,N_15881,N_12364);
and U17671 (N_17671,N_15908,N_15693);
or U17672 (N_17672,N_13312,N_15346);
and U17673 (N_17673,N_13131,N_12722);
and U17674 (N_17674,N_12026,N_15681);
and U17675 (N_17675,N_13773,N_12593);
nor U17676 (N_17676,N_14625,N_12205);
nand U17677 (N_17677,N_12157,N_14516);
and U17678 (N_17678,N_14032,N_15690);
nand U17679 (N_17679,N_14909,N_15337);
or U17680 (N_17680,N_14944,N_14327);
or U17681 (N_17681,N_14567,N_13503);
and U17682 (N_17682,N_15779,N_14215);
nand U17683 (N_17683,N_12045,N_15096);
nor U17684 (N_17684,N_15422,N_14351);
and U17685 (N_17685,N_15209,N_15320);
xor U17686 (N_17686,N_14127,N_13787);
nand U17687 (N_17687,N_14447,N_15725);
and U17688 (N_17688,N_12194,N_15302);
and U17689 (N_17689,N_14919,N_15322);
or U17690 (N_17690,N_15423,N_14835);
nand U17691 (N_17691,N_14159,N_12120);
xor U17692 (N_17692,N_15935,N_13558);
or U17693 (N_17693,N_15420,N_15204);
nor U17694 (N_17694,N_15869,N_14901);
nor U17695 (N_17695,N_15859,N_12622);
nor U17696 (N_17696,N_14794,N_12553);
and U17697 (N_17697,N_15371,N_14923);
xor U17698 (N_17698,N_12870,N_12861);
xor U17699 (N_17699,N_13138,N_12001);
or U17700 (N_17700,N_12916,N_15657);
and U17701 (N_17701,N_12253,N_15117);
xor U17702 (N_17702,N_14069,N_15661);
nand U17703 (N_17703,N_13340,N_12002);
and U17704 (N_17704,N_14668,N_12766);
xnor U17705 (N_17705,N_14008,N_12031);
xnor U17706 (N_17706,N_12477,N_15393);
or U17707 (N_17707,N_15301,N_12047);
and U17708 (N_17708,N_12086,N_14188);
nand U17709 (N_17709,N_12822,N_14642);
nand U17710 (N_17710,N_15744,N_12118);
xnor U17711 (N_17711,N_15082,N_15880);
or U17712 (N_17712,N_13387,N_14647);
or U17713 (N_17713,N_14990,N_12945);
or U17714 (N_17714,N_15333,N_12150);
or U17715 (N_17715,N_15664,N_15933);
nor U17716 (N_17716,N_14094,N_13956);
or U17717 (N_17717,N_14800,N_12814);
and U17718 (N_17718,N_12147,N_15660);
and U17719 (N_17719,N_15274,N_14554);
nand U17720 (N_17720,N_13858,N_14932);
nor U17721 (N_17721,N_15629,N_12414);
or U17722 (N_17722,N_14883,N_14630);
and U17723 (N_17723,N_12987,N_14820);
nor U17724 (N_17724,N_13368,N_15109);
xnor U17725 (N_17725,N_14880,N_13992);
nor U17726 (N_17726,N_14566,N_15714);
xor U17727 (N_17727,N_15269,N_13626);
nor U17728 (N_17728,N_14855,N_13297);
xnor U17729 (N_17729,N_15074,N_15864);
or U17730 (N_17730,N_13781,N_14994);
and U17731 (N_17731,N_13790,N_12000);
nor U17732 (N_17732,N_15294,N_14427);
xnor U17733 (N_17733,N_14424,N_12513);
or U17734 (N_17734,N_15000,N_12522);
or U17735 (N_17735,N_13227,N_14675);
or U17736 (N_17736,N_15101,N_14798);
nand U17737 (N_17737,N_13652,N_13975);
nand U17738 (N_17738,N_12375,N_14001);
or U17739 (N_17739,N_15363,N_12431);
or U17740 (N_17740,N_14464,N_13323);
nand U17741 (N_17741,N_15290,N_14745);
and U17742 (N_17742,N_15857,N_13676);
or U17743 (N_17743,N_15617,N_15846);
nor U17744 (N_17744,N_15707,N_14103);
and U17745 (N_17745,N_14446,N_13959);
or U17746 (N_17746,N_14017,N_13101);
and U17747 (N_17747,N_14591,N_14076);
nor U17748 (N_17748,N_15055,N_15666);
or U17749 (N_17749,N_15115,N_12536);
and U17750 (N_17750,N_13778,N_15426);
xor U17751 (N_17751,N_13880,N_12399);
or U17752 (N_17752,N_15809,N_15066);
nor U17753 (N_17753,N_13533,N_14808);
or U17754 (N_17754,N_12558,N_12869);
nor U17755 (N_17755,N_14585,N_13016);
nor U17756 (N_17756,N_15882,N_14669);
nor U17757 (N_17757,N_15701,N_15293);
nand U17758 (N_17758,N_13844,N_14345);
nand U17759 (N_17759,N_12899,N_15793);
xnor U17760 (N_17760,N_15285,N_13837);
and U17761 (N_17761,N_15223,N_12749);
nand U17762 (N_17762,N_12436,N_15300);
or U17763 (N_17763,N_13158,N_13137);
or U17764 (N_17764,N_14160,N_14471);
nand U17765 (N_17765,N_15949,N_13212);
or U17766 (N_17766,N_13293,N_14020);
or U17767 (N_17767,N_12459,N_12879);
nand U17768 (N_17768,N_14683,N_14730);
xor U17769 (N_17769,N_14165,N_13780);
and U17770 (N_17770,N_15240,N_12855);
nor U17771 (N_17771,N_14905,N_14132);
xnor U17772 (N_17772,N_14125,N_15476);
or U17773 (N_17773,N_14050,N_14047);
nor U17774 (N_17774,N_13894,N_12384);
or U17775 (N_17775,N_13770,N_14700);
and U17776 (N_17776,N_15745,N_14651);
nand U17777 (N_17777,N_15046,N_13074);
or U17778 (N_17778,N_15569,N_15784);
and U17779 (N_17779,N_13372,N_14773);
xor U17780 (N_17780,N_14939,N_15905);
nor U17781 (N_17781,N_12007,N_15800);
xnor U17782 (N_17782,N_15647,N_13602);
or U17783 (N_17783,N_14293,N_13037);
or U17784 (N_17784,N_13242,N_12696);
nand U17785 (N_17785,N_12112,N_14912);
xnor U17786 (N_17786,N_14370,N_15710);
or U17787 (N_17787,N_15402,N_13540);
nand U17788 (N_17788,N_14618,N_12117);
xor U17789 (N_17789,N_12648,N_15662);
or U17790 (N_17790,N_12111,N_13239);
xor U17791 (N_17791,N_15277,N_15805);
nand U17792 (N_17792,N_12089,N_14537);
and U17793 (N_17793,N_14407,N_12601);
xor U17794 (N_17794,N_15119,N_12487);
nand U17795 (N_17795,N_12844,N_15843);
or U17796 (N_17796,N_14311,N_13088);
nand U17797 (N_17797,N_15028,N_12351);
nor U17798 (N_17798,N_15724,N_13077);
and U17799 (N_17799,N_12303,N_14617);
or U17800 (N_17800,N_14493,N_12229);
nand U17801 (N_17801,N_15582,N_15137);
xor U17802 (N_17802,N_13930,N_12017);
and U17803 (N_17803,N_14343,N_14737);
nand U17804 (N_17804,N_14436,N_12791);
xnor U17805 (N_17805,N_15039,N_13035);
xnor U17806 (N_17806,N_13538,N_12254);
nand U17807 (N_17807,N_12721,N_12018);
nand U17808 (N_17808,N_13383,N_15901);
nand U17809 (N_17809,N_14904,N_14114);
and U17810 (N_17810,N_15138,N_15142);
nor U17811 (N_17811,N_15354,N_15885);
nor U17812 (N_17812,N_14336,N_13552);
nor U17813 (N_17813,N_14386,N_13847);
and U17814 (N_17814,N_14111,N_12325);
nand U17815 (N_17815,N_15827,N_14687);
and U17816 (N_17816,N_14214,N_15966);
xnor U17817 (N_17817,N_13048,N_13586);
xnor U17818 (N_17818,N_13208,N_12286);
and U17819 (N_17819,N_12841,N_14830);
and U17820 (N_17820,N_12592,N_14016);
nand U17821 (N_17821,N_14736,N_14500);
or U17822 (N_17822,N_15391,N_12510);
nor U17823 (N_17823,N_12852,N_12193);
or U17824 (N_17824,N_13246,N_13522);
and U17825 (N_17825,N_15833,N_13213);
nor U17826 (N_17826,N_12765,N_12866);
nor U17827 (N_17827,N_14194,N_12751);
and U17828 (N_17828,N_12746,N_15501);
xnor U17829 (N_17829,N_12900,N_13236);
or U17830 (N_17830,N_14143,N_15243);
and U17831 (N_17831,N_13218,N_14135);
xor U17832 (N_17832,N_14406,N_12104);
nor U17833 (N_17833,N_14130,N_12817);
xor U17834 (N_17834,N_14930,N_12750);
xnor U17835 (N_17835,N_14547,N_15735);
nand U17836 (N_17836,N_12826,N_12195);
and U17837 (N_17837,N_15641,N_15444);
or U17838 (N_17838,N_13892,N_12231);
or U17839 (N_17839,N_13179,N_13311);
or U17840 (N_17840,N_15810,N_13634);
and U17841 (N_17841,N_12445,N_14201);
nor U17842 (N_17842,N_12332,N_12886);
and U17843 (N_17843,N_12734,N_12629);
and U17844 (N_17844,N_15773,N_14914);
and U17845 (N_17845,N_14916,N_13044);
nor U17846 (N_17846,N_13338,N_14899);
or U17847 (N_17847,N_13014,N_15456);
nand U17848 (N_17848,N_14838,N_14584);
or U17849 (N_17849,N_15021,N_12406);
xnor U17850 (N_17850,N_13196,N_15944);
and U17851 (N_17851,N_15568,N_12584);
xor U17852 (N_17852,N_12429,N_15658);
and U17853 (N_17853,N_13107,N_12066);
nand U17854 (N_17854,N_13058,N_12509);
or U17855 (N_17855,N_14290,N_12336);
nor U17856 (N_17856,N_13469,N_12223);
xnor U17857 (N_17857,N_14175,N_15367);
and U17858 (N_17858,N_12461,N_14150);
nor U17859 (N_17859,N_12697,N_12546);
nor U17860 (N_17860,N_13502,N_14843);
xor U17861 (N_17861,N_14928,N_12202);
and U17862 (N_17862,N_13140,N_15824);
xnor U17863 (N_17863,N_14526,N_14036);
or U17864 (N_17864,N_14355,N_13957);
or U17865 (N_17865,N_12289,N_14140);
nand U17866 (N_17866,N_14534,N_13555);
or U17867 (N_17867,N_15914,N_13341);
nand U17868 (N_17868,N_14792,N_12395);
nor U17869 (N_17869,N_12912,N_15339);
xor U17870 (N_17870,N_12981,N_15706);
nor U17871 (N_17871,N_13299,N_13364);
nand U17872 (N_17872,N_12891,N_13961);
or U17873 (N_17873,N_14673,N_15177);
nor U17874 (N_17874,N_13549,N_13680);
nor U17875 (N_17875,N_13322,N_15670);
nand U17876 (N_17876,N_15412,N_15336);
nor U17877 (N_17877,N_12634,N_14558);
and U17878 (N_17878,N_12608,N_13546);
and U17879 (N_17879,N_12101,N_13718);
or U17880 (N_17880,N_13112,N_12251);
and U17881 (N_17881,N_12581,N_15266);
xor U17882 (N_17882,N_13681,N_14339);
nor U17883 (N_17883,N_13838,N_14102);
xnor U17884 (N_17884,N_12798,N_14559);
nor U17885 (N_17885,N_12966,N_13380);
or U17886 (N_17886,N_13564,N_12716);
nand U17887 (N_17887,N_12709,N_12654);
nand U17888 (N_17888,N_13960,N_12097);
nand U17889 (N_17889,N_14079,N_15536);
and U17890 (N_17890,N_14759,N_12235);
nor U17891 (N_17891,N_15173,N_12070);
xor U17892 (N_17892,N_13303,N_13418);
nand U17893 (N_17893,N_14713,N_14390);
xor U17894 (N_17894,N_13116,N_12965);
and U17895 (N_17895,N_14744,N_15937);
nand U17896 (N_17896,N_13997,N_12859);
and U17897 (N_17897,N_14860,N_13941);
and U17898 (N_17898,N_14120,N_13905);
or U17899 (N_17899,N_13098,N_14621);
nand U17900 (N_17900,N_13643,N_12681);
and U17901 (N_17901,N_14531,N_14524);
xnor U17902 (N_17902,N_15340,N_12282);
xnor U17903 (N_17903,N_15017,N_12136);
xor U17904 (N_17904,N_14693,N_13859);
or U17905 (N_17905,N_13134,N_15778);
xor U17906 (N_17906,N_14985,N_13490);
or U17907 (N_17907,N_14368,N_12222);
nor U17908 (N_17908,N_12778,N_14892);
xor U17909 (N_17909,N_15313,N_12252);
nand U17910 (N_17910,N_13537,N_13748);
nand U17911 (N_17911,N_15226,N_12690);
or U17912 (N_17912,N_15633,N_12209);
or U17913 (N_17913,N_15384,N_15500);
or U17914 (N_17914,N_15174,N_14510);
nand U17915 (N_17915,N_14631,N_13283);
nand U17916 (N_17916,N_14320,N_13840);
and U17917 (N_17917,N_13104,N_13561);
or U17918 (N_17918,N_14469,N_12280);
nor U17919 (N_17919,N_12006,N_14026);
nand U17920 (N_17920,N_12386,N_12494);
nand U17921 (N_17921,N_14477,N_13620);
or U17922 (N_17922,N_13573,N_15373);
xor U17923 (N_17923,N_15530,N_14015);
nor U17924 (N_17924,N_13800,N_14989);
and U17925 (N_17925,N_12856,N_12851);
xor U17926 (N_17926,N_13206,N_14506);
xnor U17927 (N_17927,N_14139,N_15280);
nor U17928 (N_17928,N_15523,N_12259);
xnor U17929 (N_17929,N_13084,N_13842);
nand U17930 (N_17930,N_12065,N_13576);
nand U17931 (N_17931,N_14813,N_12257);
or U17932 (N_17932,N_14338,N_15178);
xor U17933 (N_17933,N_14382,N_14233);
xor U17934 (N_17934,N_14208,N_14988);
nand U17935 (N_17935,N_14666,N_14470);
nor U17936 (N_17936,N_14523,N_12272);
xor U17937 (N_17937,N_14080,N_12409);
and U17938 (N_17938,N_15148,N_12463);
and U17939 (N_17939,N_13585,N_12483);
nor U17940 (N_17940,N_12578,N_14539);
nand U17941 (N_17941,N_13360,N_13029);
xor U17942 (N_17942,N_13381,N_15413);
xnor U17943 (N_17943,N_12256,N_15491);
or U17944 (N_17944,N_14329,N_12273);
and U17945 (N_17945,N_15158,N_14044);
xor U17946 (N_17946,N_15786,N_14908);
or U17947 (N_17947,N_12612,N_13321);
nand U17948 (N_17948,N_14750,N_15750);
and U17949 (N_17949,N_15763,N_15085);
nand U17950 (N_17950,N_14465,N_15092);
nor U17951 (N_17951,N_15125,N_12764);
or U17952 (N_17952,N_15732,N_12501);
and U17953 (N_17953,N_15128,N_14925);
xnor U17954 (N_17954,N_12555,N_14299);
xnor U17955 (N_17955,N_14035,N_14662);
xor U17956 (N_17956,N_13407,N_12962);
xor U17957 (N_17957,N_14845,N_12636);
or U17958 (N_17958,N_14910,N_12440);
xnor U17959 (N_17959,N_12700,N_12175);
or U17960 (N_17960,N_15076,N_14216);
or U17961 (N_17961,N_12880,N_14661);
nor U17962 (N_17962,N_15127,N_14412);
nor U17963 (N_17963,N_15700,N_13940);
or U17964 (N_17964,N_15299,N_12473);
nand U17965 (N_17965,N_13090,N_15347);
nand U17966 (N_17966,N_15802,N_15819);
nor U17967 (N_17967,N_14024,N_12182);
nand U17968 (N_17968,N_12176,N_15205);
nand U17969 (N_17969,N_15644,N_14601);
nor U17970 (N_17970,N_15554,N_12519);
xnor U17971 (N_17971,N_14378,N_13588);
or U17972 (N_17972,N_12911,N_12439);
and U17973 (N_17973,N_15595,N_12616);
nor U17974 (N_17974,N_14870,N_13603);
xnor U17975 (N_17975,N_13874,N_14422);
nand U17976 (N_17976,N_14777,N_14941);
xor U17977 (N_17977,N_13827,N_12040);
or U17978 (N_17978,N_13510,N_14402);
or U17979 (N_17979,N_14115,N_15973);
xnor U17980 (N_17980,N_13793,N_13256);
or U17981 (N_17981,N_12927,N_14717);
nor U17982 (N_17982,N_12688,N_13120);
xor U17983 (N_17983,N_14868,N_12119);
nand U17984 (N_17984,N_13911,N_14073);
nor U17985 (N_17985,N_13295,N_13574);
and U17986 (N_17986,N_15229,N_15815);
nor U17987 (N_17987,N_15928,N_14867);
xnor U17988 (N_17988,N_12686,N_14189);
nand U17989 (N_17989,N_15197,N_13426);
and U17990 (N_17990,N_13307,N_15090);
and U17991 (N_17991,N_13810,N_15103);
or U17992 (N_17992,N_13798,N_15853);
nand U17993 (N_17993,N_12090,N_14240);
nor U17994 (N_17994,N_13872,N_14931);
nand U17995 (N_17995,N_12970,N_12037);
nor U17996 (N_17996,N_15359,N_14065);
or U17997 (N_17997,N_15202,N_14671);
nand U17998 (N_17998,N_15608,N_14884);
xor U17999 (N_17999,N_13190,N_13513);
and U18000 (N_18000,N_13953,N_14148);
nor U18001 (N_18001,N_14188,N_12437);
and U18002 (N_18002,N_15498,N_13076);
nor U18003 (N_18003,N_12052,N_15357);
or U18004 (N_18004,N_15145,N_15116);
or U18005 (N_18005,N_15849,N_13102);
nor U18006 (N_18006,N_13058,N_15216);
xor U18007 (N_18007,N_15839,N_12765);
nand U18008 (N_18008,N_15529,N_15158);
nor U18009 (N_18009,N_13890,N_15439);
or U18010 (N_18010,N_13043,N_13011);
xnor U18011 (N_18011,N_15987,N_12252);
xor U18012 (N_18012,N_13267,N_13562);
nand U18013 (N_18013,N_15405,N_13946);
or U18014 (N_18014,N_14170,N_13497);
nand U18015 (N_18015,N_14255,N_12557);
nor U18016 (N_18016,N_15686,N_14832);
and U18017 (N_18017,N_13274,N_15269);
and U18018 (N_18018,N_14977,N_12342);
xnor U18019 (N_18019,N_13851,N_12211);
or U18020 (N_18020,N_15729,N_15969);
and U18021 (N_18021,N_14745,N_15980);
nor U18022 (N_18022,N_12161,N_15810);
xor U18023 (N_18023,N_13836,N_14183);
xnor U18024 (N_18024,N_13545,N_13751);
nand U18025 (N_18025,N_14117,N_14569);
nand U18026 (N_18026,N_13524,N_13478);
xor U18027 (N_18027,N_15482,N_13658);
or U18028 (N_18028,N_14827,N_15566);
nand U18029 (N_18029,N_15840,N_12975);
xor U18030 (N_18030,N_15561,N_12610);
nor U18031 (N_18031,N_15076,N_12130);
nor U18032 (N_18032,N_14691,N_14946);
nand U18033 (N_18033,N_12775,N_15743);
or U18034 (N_18034,N_14209,N_15469);
nand U18035 (N_18035,N_14726,N_14322);
or U18036 (N_18036,N_12171,N_14873);
nor U18037 (N_18037,N_15133,N_14540);
xnor U18038 (N_18038,N_13251,N_13707);
and U18039 (N_18039,N_14199,N_12720);
nand U18040 (N_18040,N_15223,N_15773);
and U18041 (N_18041,N_15997,N_12638);
or U18042 (N_18042,N_15704,N_15551);
xor U18043 (N_18043,N_12634,N_12956);
nand U18044 (N_18044,N_14720,N_12470);
nand U18045 (N_18045,N_12797,N_12377);
nand U18046 (N_18046,N_15566,N_15559);
nand U18047 (N_18047,N_14858,N_12823);
or U18048 (N_18048,N_12132,N_15224);
or U18049 (N_18049,N_14341,N_13696);
or U18050 (N_18050,N_13716,N_12593);
xor U18051 (N_18051,N_14828,N_15914);
xnor U18052 (N_18052,N_12938,N_14724);
xnor U18053 (N_18053,N_15627,N_15739);
and U18054 (N_18054,N_12207,N_14072);
or U18055 (N_18055,N_13650,N_15332);
xor U18056 (N_18056,N_14855,N_12274);
or U18057 (N_18057,N_12036,N_15456);
nor U18058 (N_18058,N_15268,N_14189);
and U18059 (N_18059,N_12865,N_15501);
nor U18060 (N_18060,N_14857,N_15913);
xor U18061 (N_18061,N_13360,N_13881);
nand U18062 (N_18062,N_12325,N_14768);
or U18063 (N_18063,N_15078,N_14277);
or U18064 (N_18064,N_14528,N_12248);
nand U18065 (N_18065,N_12481,N_12750);
nor U18066 (N_18066,N_13506,N_13018);
nand U18067 (N_18067,N_15153,N_14010);
or U18068 (N_18068,N_12735,N_15119);
nor U18069 (N_18069,N_13321,N_12752);
and U18070 (N_18070,N_13701,N_13414);
xor U18071 (N_18071,N_13090,N_12089);
xnor U18072 (N_18072,N_12593,N_12825);
and U18073 (N_18073,N_14992,N_14124);
nor U18074 (N_18074,N_14268,N_13869);
xor U18075 (N_18075,N_13472,N_13144);
nand U18076 (N_18076,N_14101,N_12022);
nor U18077 (N_18077,N_14756,N_12718);
xnor U18078 (N_18078,N_14609,N_12469);
and U18079 (N_18079,N_13380,N_13713);
or U18080 (N_18080,N_15013,N_13799);
nor U18081 (N_18081,N_12612,N_13591);
xor U18082 (N_18082,N_14863,N_14040);
nor U18083 (N_18083,N_14407,N_14659);
and U18084 (N_18084,N_15430,N_13010);
or U18085 (N_18085,N_14517,N_13503);
nand U18086 (N_18086,N_12573,N_14102);
nor U18087 (N_18087,N_15971,N_13290);
xor U18088 (N_18088,N_13582,N_14817);
xnor U18089 (N_18089,N_12117,N_14559);
nor U18090 (N_18090,N_13266,N_15254);
and U18091 (N_18091,N_15670,N_12984);
xnor U18092 (N_18092,N_14044,N_15656);
and U18093 (N_18093,N_12935,N_13085);
or U18094 (N_18094,N_15168,N_13811);
and U18095 (N_18095,N_13412,N_13313);
nand U18096 (N_18096,N_15644,N_13253);
xnor U18097 (N_18097,N_15718,N_12358);
xor U18098 (N_18098,N_13258,N_15118);
or U18099 (N_18099,N_14776,N_15860);
nand U18100 (N_18100,N_14870,N_14156);
xnor U18101 (N_18101,N_15950,N_15039);
or U18102 (N_18102,N_12674,N_12218);
or U18103 (N_18103,N_15409,N_15195);
nand U18104 (N_18104,N_12547,N_13310);
nand U18105 (N_18105,N_14152,N_13957);
and U18106 (N_18106,N_13388,N_14288);
nand U18107 (N_18107,N_15910,N_15003);
or U18108 (N_18108,N_15826,N_14169);
xor U18109 (N_18109,N_14540,N_13424);
or U18110 (N_18110,N_12763,N_15837);
nor U18111 (N_18111,N_13750,N_15251);
and U18112 (N_18112,N_14535,N_12149);
xnor U18113 (N_18113,N_15894,N_14680);
or U18114 (N_18114,N_14611,N_15758);
nand U18115 (N_18115,N_15179,N_13892);
and U18116 (N_18116,N_15216,N_14124);
or U18117 (N_18117,N_14860,N_12078);
and U18118 (N_18118,N_14773,N_15387);
xor U18119 (N_18119,N_14686,N_14678);
nand U18120 (N_18120,N_15944,N_14898);
and U18121 (N_18121,N_13013,N_14451);
nand U18122 (N_18122,N_13390,N_12548);
nor U18123 (N_18123,N_13085,N_13868);
nand U18124 (N_18124,N_13722,N_13653);
or U18125 (N_18125,N_14197,N_14330);
or U18126 (N_18126,N_15185,N_15446);
or U18127 (N_18127,N_14038,N_15408);
nor U18128 (N_18128,N_15737,N_12928);
xor U18129 (N_18129,N_15556,N_12259);
xnor U18130 (N_18130,N_12465,N_13285);
nor U18131 (N_18131,N_15538,N_13351);
nand U18132 (N_18132,N_14267,N_15280);
xor U18133 (N_18133,N_15573,N_13774);
nor U18134 (N_18134,N_13513,N_14153);
xor U18135 (N_18135,N_14875,N_15208);
nand U18136 (N_18136,N_12722,N_15736);
nor U18137 (N_18137,N_13141,N_15925);
nand U18138 (N_18138,N_15879,N_12114);
or U18139 (N_18139,N_14635,N_12421);
and U18140 (N_18140,N_12964,N_13790);
xor U18141 (N_18141,N_12891,N_12013);
nand U18142 (N_18142,N_13484,N_15829);
and U18143 (N_18143,N_15310,N_14214);
and U18144 (N_18144,N_15834,N_13152);
xnor U18145 (N_18145,N_15092,N_13554);
xor U18146 (N_18146,N_13173,N_13051);
nand U18147 (N_18147,N_12200,N_12685);
nor U18148 (N_18148,N_12530,N_15274);
or U18149 (N_18149,N_15269,N_14687);
or U18150 (N_18150,N_15277,N_13911);
or U18151 (N_18151,N_13123,N_14910);
and U18152 (N_18152,N_14655,N_14471);
and U18153 (N_18153,N_15257,N_12399);
or U18154 (N_18154,N_12761,N_12776);
or U18155 (N_18155,N_12423,N_14163);
nor U18156 (N_18156,N_14522,N_12020);
nor U18157 (N_18157,N_15546,N_14899);
or U18158 (N_18158,N_15548,N_12153);
nor U18159 (N_18159,N_13805,N_15312);
and U18160 (N_18160,N_12791,N_13551);
nand U18161 (N_18161,N_15526,N_12463);
or U18162 (N_18162,N_15970,N_13444);
xor U18163 (N_18163,N_14544,N_12394);
nor U18164 (N_18164,N_14770,N_14627);
and U18165 (N_18165,N_15521,N_13440);
or U18166 (N_18166,N_14737,N_15654);
or U18167 (N_18167,N_14974,N_14523);
xnor U18168 (N_18168,N_15780,N_14984);
nand U18169 (N_18169,N_14833,N_14702);
nand U18170 (N_18170,N_14020,N_15775);
xor U18171 (N_18171,N_14167,N_13625);
xnor U18172 (N_18172,N_14620,N_15046);
and U18173 (N_18173,N_13344,N_14842);
nand U18174 (N_18174,N_14888,N_15639);
nand U18175 (N_18175,N_15106,N_13990);
xnor U18176 (N_18176,N_15647,N_14182);
nor U18177 (N_18177,N_12251,N_15824);
nor U18178 (N_18178,N_15128,N_14773);
or U18179 (N_18179,N_13863,N_15811);
nand U18180 (N_18180,N_15561,N_13886);
and U18181 (N_18181,N_13367,N_13340);
and U18182 (N_18182,N_14298,N_14736);
and U18183 (N_18183,N_12137,N_13592);
or U18184 (N_18184,N_14315,N_15362);
nor U18185 (N_18185,N_13757,N_12976);
xnor U18186 (N_18186,N_15156,N_12019);
nand U18187 (N_18187,N_15530,N_12755);
xnor U18188 (N_18188,N_12102,N_12116);
nor U18189 (N_18189,N_15189,N_13925);
nor U18190 (N_18190,N_12692,N_15777);
and U18191 (N_18191,N_13038,N_12282);
nor U18192 (N_18192,N_15374,N_15399);
or U18193 (N_18193,N_13570,N_12133);
nand U18194 (N_18194,N_13126,N_13209);
nand U18195 (N_18195,N_14999,N_12388);
nand U18196 (N_18196,N_15437,N_14060);
nor U18197 (N_18197,N_14110,N_13408);
or U18198 (N_18198,N_12810,N_13919);
nand U18199 (N_18199,N_14349,N_13669);
nor U18200 (N_18200,N_13949,N_13176);
nor U18201 (N_18201,N_15452,N_13443);
and U18202 (N_18202,N_15881,N_15288);
nand U18203 (N_18203,N_13926,N_13801);
or U18204 (N_18204,N_14661,N_14204);
and U18205 (N_18205,N_12557,N_12936);
nor U18206 (N_18206,N_15124,N_13981);
nor U18207 (N_18207,N_15227,N_13813);
nor U18208 (N_18208,N_14420,N_14757);
nor U18209 (N_18209,N_13609,N_14075);
or U18210 (N_18210,N_12245,N_13093);
xnor U18211 (N_18211,N_14954,N_13372);
nand U18212 (N_18212,N_15718,N_13366);
and U18213 (N_18213,N_13466,N_13213);
nor U18214 (N_18214,N_14257,N_14686);
nor U18215 (N_18215,N_14906,N_13104);
xor U18216 (N_18216,N_14690,N_14098);
xor U18217 (N_18217,N_14347,N_13278);
xor U18218 (N_18218,N_14942,N_15297);
or U18219 (N_18219,N_14157,N_13186);
and U18220 (N_18220,N_14543,N_13442);
or U18221 (N_18221,N_12616,N_13085);
nor U18222 (N_18222,N_14991,N_13057);
and U18223 (N_18223,N_14361,N_12206);
nand U18224 (N_18224,N_15325,N_15394);
and U18225 (N_18225,N_15003,N_12371);
or U18226 (N_18226,N_14582,N_12628);
nand U18227 (N_18227,N_14978,N_14633);
or U18228 (N_18228,N_13158,N_12982);
and U18229 (N_18229,N_14758,N_13512);
and U18230 (N_18230,N_13417,N_15058);
xor U18231 (N_18231,N_14635,N_14803);
and U18232 (N_18232,N_15754,N_14248);
and U18233 (N_18233,N_13361,N_13026);
xnor U18234 (N_18234,N_15970,N_12029);
nand U18235 (N_18235,N_12850,N_12338);
and U18236 (N_18236,N_14497,N_12572);
or U18237 (N_18237,N_12120,N_15937);
nor U18238 (N_18238,N_14740,N_12651);
nand U18239 (N_18239,N_15268,N_13298);
and U18240 (N_18240,N_14642,N_13219);
xor U18241 (N_18241,N_13322,N_15650);
nand U18242 (N_18242,N_12709,N_13074);
nand U18243 (N_18243,N_12845,N_12439);
and U18244 (N_18244,N_15292,N_15525);
and U18245 (N_18245,N_14488,N_13050);
nand U18246 (N_18246,N_13712,N_15566);
or U18247 (N_18247,N_15541,N_15927);
nand U18248 (N_18248,N_14757,N_12624);
and U18249 (N_18249,N_14544,N_12052);
xor U18250 (N_18250,N_12494,N_12697);
xor U18251 (N_18251,N_12429,N_13292);
nor U18252 (N_18252,N_15954,N_15369);
nor U18253 (N_18253,N_13489,N_13921);
nor U18254 (N_18254,N_12620,N_13079);
nor U18255 (N_18255,N_13736,N_12995);
xor U18256 (N_18256,N_13024,N_14486);
and U18257 (N_18257,N_12957,N_15462);
nand U18258 (N_18258,N_12270,N_13432);
nand U18259 (N_18259,N_15451,N_12984);
xnor U18260 (N_18260,N_15543,N_13252);
and U18261 (N_18261,N_12337,N_15773);
nand U18262 (N_18262,N_13142,N_14728);
nand U18263 (N_18263,N_14432,N_12154);
xor U18264 (N_18264,N_13453,N_14250);
nor U18265 (N_18265,N_14104,N_15005);
nand U18266 (N_18266,N_15317,N_12926);
nand U18267 (N_18267,N_13325,N_13699);
and U18268 (N_18268,N_15025,N_15341);
xor U18269 (N_18269,N_13602,N_15544);
nor U18270 (N_18270,N_15765,N_14146);
nand U18271 (N_18271,N_14870,N_13023);
or U18272 (N_18272,N_13292,N_15073);
nor U18273 (N_18273,N_14127,N_14942);
nand U18274 (N_18274,N_15340,N_15454);
nor U18275 (N_18275,N_15203,N_15133);
and U18276 (N_18276,N_13523,N_12224);
nor U18277 (N_18277,N_12810,N_12881);
or U18278 (N_18278,N_13685,N_13948);
xnor U18279 (N_18279,N_12329,N_14399);
nor U18280 (N_18280,N_12967,N_12613);
or U18281 (N_18281,N_12102,N_15849);
nor U18282 (N_18282,N_13069,N_12777);
xnor U18283 (N_18283,N_14695,N_14666);
or U18284 (N_18284,N_15630,N_15024);
or U18285 (N_18285,N_14900,N_15994);
nand U18286 (N_18286,N_14302,N_13517);
nand U18287 (N_18287,N_14636,N_15481);
and U18288 (N_18288,N_13886,N_14363);
or U18289 (N_18289,N_14694,N_12517);
and U18290 (N_18290,N_13362,N_14143);
nor U18291 (N_18291,N_12635,N_15127);
nand U18292 (N_18292,N_13801,N_15137);
nand U18293 (N_18293,N_15423,N_15061);
and U18294 (N_18294,N_15893,N_12076);
nor U18295 (N_18295,N_14818,N_12638);
or U18296 (N_18296,N_13452,N_13267);
nand U18297 (N_18297,N_15085,N_12466);
nand U18298 (N_18298,N_12382,N_14684);
and U18299 (N_18299,N_12591,N_14328);
nand U18300 (N_18300,N_15176,N_13231);
xor U18301 (N_18301,N_14407,N_15100);
xnor U18302 (N_18302,N_15407,N_15615);
nand U18303 (N_18303,N_14635,N_15752);
nor U18304 (N_18304,N_14889,N_13627);
xnor U18305 (N_18305,N_14289,N_13962);
nand U18306 (N_18306,N_12790,N_13733);
xnor U18307 (N_18307,N_13950,N_12161);
xnor U18308 (N_18308,N_13300,N_15008);
xnor U18309 (N_18309,N_15861,N_15419);
nor U18310 (N_18310,N_14296,N_14896);
or U18311 (N_18311,N_15080,N_14083);
or U18312 (N_18312,N_13475,N_13162);
or U18313 (N_18313,N_13018,N_13722);
or U18314 (N_18314,N_14105,N_14967);
nor U18315 (N_18315,N_15779,N_13357);
or U18316 (N_18316,N_14614,N_14180);
nor U18317 (N_18317,N_12285,N_13123);
xnor U18318 (N_18318,N_14074,N_12731);
xor U18319 (N_18319,N_14865,N_12241);
and U18320 (N_18320,N_15174,N_13824);
nand U18321 (N_18321,N_13214,N_14670);
or U18322 (N_18322,N_12657,N_15517);
xor U18323 (N_18323,N_15677,N_14138);
and U18324 (N_18324,N_14962,N_14019);
nand U18325 (N_18325,N_13128,N_13334);
xor U18326 (N_18326,N_14932,N_12088);
or U18327 (N_18327,N_14774,N_13735);
or U18328 (N_18328,N_13390,N_15888);
or U18329 (N_18329,N_13153,N_15657);
and U18330 (N_18330,N_13367,N_13712);
and U18331 (N_18331,N_14489,N_12400);
nor U18332 (N_18332,N_15239,N_13610);
or U18333 (N_18333,N_15170,N_15240);
or U18334 (N_18334,N_12002,N_12038);
xnor U18335 (N_18335,N_12211,N_13019);
or U18336 (N_18336,N_13844,N_14480);
nor U18337 (N_18337,N_13739,N_15066);
nor U18338 (N_18338,N_12859,N_15780);
or U18339 (N_18339,N_13821,N_12810);
nor U18340 (N_18340,N_15672,N_14624);
or U18341 (N_18341,N_14181,N_14338);
and U18342 (N_18342,N_14626,N_15247);
and U18343 (N_18343,N_12964,N_12893);
nor U18344 (N_18344,N_14258,N_14229);
xnor U18345 (N_18345,N_13381,N_12791);
and U18346 (N_18346,N_14802,N_14081);
nor U18347 (N_18347,N_15898,N_14451);
nor U18348 (N_18348,N_14703,N_15191);
nor U18349 (N_18349,N_15894,N_15982);
nand U18350 (N_18350,N_14784,N_15860);
or U18351 (N_18351,N_12584,N_12003);
nand U18352 (N_18352,N_14301,N_15561);
nor U18353 (N_18353,N_14442,N_14563);
xnor U18354 (N_18354,N_14196,N_12166);
or U18355 (N_18355,N_15807,N_14601);
nand U18356 (N_18356,N_12214,N_13294);
xor U18357 (N_18357,N_14485,N_15486);
nor U18358 (N_18358,N_15795,N_15013);
nor U18359 (N_18359,N_14430,N_12191);
xor U18360 (N_18360,N_15722,N_14343);
xor U18361 (N_18361,N_14699,N_12891);
nand U18362 (N_18362,N_13630,N_14887);
and U18363 (N_18363,N_13382,N_13930);
nand U18364 (N_18364,N_14255,N_12424);
nor U18365 (N_18365,N_12926,N_13431);
nor U18366 (N_18366,N_15648,N_15331);
and U18367 (N_18367,N_13863,N_13107);
nor U18368 (N_18368,N_14588,N_14610);
nor U18369 (N_18369,N_14213,N_13538);
and U18370 (N_18370,N_15343,N_15549);
nand U18371 (N_18371,N_15883,N_15841);
or U18372 (N_18372,N_13326,N_13097);
nor U18373 (N_18373,N_14373,N_15264);
nand U18374 (N_18374,N_14139,N_12131);
nand U18375 (N_18375,N_14780,N_15366);
nor U18376 (N_18376,N_15298,N_12769);
nand U18377 (N_18377,N_14488,N_15094);
and U18378 (N_18378,N_12401,N_13282);
nor U18379 (N_18379,N_15792,N_15156);
or U18380 (N_18380,N_14488,N_13996);
or U18381 (N_18381,N_12836,N_14047);
xnor U18382 (N_18382,N_14345,N_13347);
nand U18383 (N_18383,N_14875,N_13223);
or U18384 (N_18384,N_14644,N_13817);
and U18385 (N_18385,N_13647,N_13050);
xnor U18386 (N_18386,N_15681,N_12759);
nor U18387 (N_18387,N_12289,N_14135);
and U18388 (N_18388,N_13657,N_14069);
xnor U18389 (N_18389,N_15320,N_13712);
or U18390 (N_18390,N_13927,N_12209);
or U18391 (N_18391,N_15258,N_14224);
and U18392 (N_18392,N_14280,N_15795);
nor U18393 (N_18393,N_13675,N_15734);
nand U18394 (N_18394,N_15738,N_12025);
nand U18395 (N_18395,N_12913,N_15849);
or U18396 (N_18396,N_12589,N_14867);
and U18397 (N_18397,N_13817,N_15034);
nor U18398 (N_18398,N_12690,N_14517);
and U18399 (N_18399,N_14191,N_15582);
or U18400 (N_18400,N_14550,N_14190);
and U18401 (N_18401,N_13143,N_14025);
or U18402 (N_18402,N_14064,N_12568);
nand U18403 (N_18403,N_13997,N_15876);
and U18404 (N_18404,N_12472,N_15439);
nand U18405 (N_18405,N_12792,N_12318);
xor U18406 (N_18406,N_14042,N_13216);
xor U18407 (N_18407,N_14163,N_12275);
xor U18408 (N_18408,N_15406,N_14248);
nor U18409 (N_18409,N_14083,N_12047);
and U18410 (N_18410,N_14969,N_15660);
xor U18411 (N_18411,N_14977,N_12102);
xor U18412 (N_18412,N_14848,N_14265);
nor U18413 (N_18413,N_13983,N_12341);
nor U18414 (N_18414,N_13405,N_12018);
nor U18415 (N_18415,N_12614,N_13910);
or U18416 (N_18416,N_12366,N_14162);
and U18417 (N_18417,N_15185,N_15438);
xor U18418 (N_18418,N_14979,N_15776);
xnor U18419 (N_18419,N_13708,N_13439);
xnor U18420 (N_18420,N_14672,N_13495);
xor U18421 (N_18421,N_15512,N_15131);
and U18422 (N_18422,N_14266,N_13980);
or U18423 (N_18423,N_13431,N_13052);
and U18424 (N_18424,N_13719,N_15726);
xnor U18425 (N_18425,N_15516,N_14594);
nand U18426 (N_18426,N_14113,N_14762);
or U18427 (N_18427,N_14478,N_15701);
nand U18428 (N_18428,N_12471,N_12307);
nand U18429 (N_18429,N_15191,N_15450);
nor U18430 (N_18430,N_14671,N_15262);
nor U18431 (N_18431,N_14833,N_12961);
xnor U18432 (N_18432,N_13468,N_13008);
nand U18433 (N_18433,N_15765,N_13885);
nand U18434 (N_18434,N_13135,N_13060);
or U18435 (N_18435,N_13621,N_13508);
or U18436 (N_18436,N_15415,N_14417);
xnor U18437 (N_18437,N_15074,N_14915);
and U18438 (N_18438,N_12926,N_13904);
nor U18439 (N_18439,N_13941,N_14534);
or U18440 (N_18440,N_12364,N_13499);
and U18441 (N_18441,N_15112,N_12171);
nor U18442 (N_18442,N_12393,N_14054);
and U18443 (N_18443,N_15043,N_13282);
nor U18444 (N_18444,N_14681,N_13532);
or U18445 (N_18445,N_15291,N_14524);
xor U18446 (N_18446,N_13230,N_15302);
nand U18447 (N_18447,N_12339,N_14005);
or U18448 (N_18448,N_14519,N_15856);
xor U18449 (N_18449,N_12763,N_13431);
nor U18450 (N_18450,N_12111,N_15031);
nand U18451 (N_18451,N_12669,N_14124);
and U18452 (N_18452,N_13420,N_15775);
and U18453 (N_18453,N_14331,N_14329);
nor U18454 (N_18454,N_13378,N_13766);
nand U18455 (N_18455,N_13271,N_12447);
and U18456 (N_18456,N_12221,N_15755);
and U18457 (N_18457,N_13675,N_13473);
nor U18458 (N_18458,N_15407,N_15746);
or U18459 (N_18459,N_13945,N_13289);
and U18460 (N_18460,N_12199,N_13066);
and U18461 (N_18461,N_15126,N_13052);
or U18462 (N_18462,N_13193,N_13796);
xnor U18463 (N_18463,N_15087,N_15386);
nand U18464 (N_18464,N_13061,N_15929);
nand U18465 (N_18465,N_14176,N_12928);
xnor U18466 (N_18466,N_14996,N_15598);
and U18467 (N_18467,N_13193,N_14678);
nand U18468 (N_18468,N_12347,N_12032);
and U18469 (N_18469,N_13894,N_13222);
nor U18470 (N_18470,N_14248,N_15402);
xnor U18471 (N_18471,N_12285,N_14075);
and U18472 (N_18472,N_12870,N_15376);
or U18473 (N_18473,N_13781,N_14622);
nand U18474 (N_18474,N_13749,N_12063);
or U18475 (N_18475,N_15350,N_13133);
and U18476 (N_18476,N_14075,N_12060);
and U18477 (N_18477,N_15558,N_13153);
xor U18478 (N_18478,N_14886,N_14147);
and U18479 (N_18479,N_15544,N_13451);
nor U18480 (N_18480,N_15632,N_13777);
or U18481 (N_18481,N_13948,N_13932);
nor U18482 (N_18482,N_14480,N_13062);
or U18483 (N_18483,N_12824,N_12357);
nor U18484 (N_18484,N_14682,N_12300);
xnor U18485 (N_18485,N_14382,N_14806);
nor U18486 (N_18486,N_14784,N_13570);
and U18487 (N_18487,N_14872,N_15043);
xor U18488 (N_18488,N_15278,N_12466);
nor U18489 (N_18489,N_15907,N_14333);
nor U18490 (N_18490,N_15991,N_12549);
xor U18491 (N_18491,N_13695,N_15157);
nor U18492 (N_18492,N_14324,N_14736);
and U18493 (N_18493,N_15142,N_13345);
nand U18494 (N_18494,N_12714,N_12793);
or U18495 (N_18495,N_14748,N_15222);
nand U18496 (N_18496,N_13672,N_13634);
and U18497 (N_18497,N_14220,N_12437);
or U18498 (N_18498,N_12669,N_12975);
and U18499 (N_18499,N_12371,N_15481);
or U18500 (N_18500,N_14459,N_14511);
xor U18501 (N_18501,N_12298,N_12465);
xor U18502 (N_18502,N_12740,N_12179);
xnor U18503 (N_18503,N_12935,N_14444);
nor U18504 (N_18504,N_13802,N_13251);
nor U18505 (N_18505,N_13478,N_15666);
and U18506 (N_18506,N_13545,N_13998);
xor U18507 (N_18507,N_15135,N_12726);
nand U18508 (N_18508,N_15097,N_15303);
nor U18509 (N_18509,N_14576,N_15745);
and U18510 (N_18510,N_12896,N_12773);
or U18511 (N_18511,N_15487,N_15267);
nand U18512 (N_18512,N_14711,N_14342);
xor U18513 (N_18513,N_14615,N_13285);
nand U18514 (N_18514,N_14775,N_12073);
xnor U18515 (N_18515,N_14299,N_13036);
nor U18516 (N_18516,N_13309,N_15581);
xor U18517 (N_18517,N_12656,N_13041);
or U18518 (N_18518,N_13370,N_12379);
or U18519 (N_18519,N_12391,N_15073);
nor U18520 (N_18520,N_13300,N_13924);
xnor U18521 (N_18521,N_12783,N_15787);
nand U18522 (N_18522,N_14358,N_14041);
and U18523 (N_18523,N_14451,N_14131);
or U18524 (N_18524,N_13981,N_14468);
nor U18525 (N_18525,N_15166,N_13526);
and U18526 (N_18526,N_12426,N_13509);
and U18527 (N_18527,N_12843,N_14439);
nand U18528 (N_18528,N_15080,N_15741);
or U18529 (N_18529,N_15681,N_15893);
nand U18530 (N_18530,N_15288,N_15548);
nor U18531 (N_18531,N_12606,N_12301);
and U18532 (N_18532,N_13282,N_12472);
nor U18533 (N_18533,N_12234,N_14645);
nor U18534 (N_18534,N_13311,N_15701);
nand U18535 (N_18535,N_12753,N_12277);
and U18536 (N_18536,N_13504,N_15461);
xor U18537 (N_18537,N_14115,N_14973);
and U18538 (N_18538,N_14937,N_13352);
nand U18539 (N_18539,N_13232,N_12229);
nor U18540 (N_18540,N_12030,N_12620);
or U18541 (N_18541,N_15224,N_13837);
nand U18542 (N_18542,N_14846,N_13585);
nor U18543 (N_18543,N_12056,N_13525);
nor U18544 (N_18544,N_14509,N_14207);
xnor U18545 (N_18545,N_13732,N_13485);
nor U18546 (N_18546,N_13970,N_14571);
or U18547 (N_18547,N_14188,N_14686);
and U18548 (N_18548,N_15698,N_13795);
nor U18549 (N_18549,N_13602,N_15181);
nand U18550 (N_18550,N_14810,N_13628);
xnor U18551 (N_18551,N_12474,N_14507);
nand U18552 (N_18552,N_12130,N_13619);
or U18553 (N_18553,N_13717,N_14809);
nand U18554 (N_18554,N_15639,N_15251);
xor U18555 (N_18555,N_14557,N_13520);
and U18556 (N_18556,N_14583,N_12903);
and U18557 (N_18557,N_14857,N_12899);
or U18558 (N_18558,N_14655,N_14036);
or U18559 (N_18559,N_15014,N_15155);
xnor U18560 (N_18560,N_15819,N_15013);
and U18561 (N_18561,N_15599,N_14031);
and U18562 (N_18562,N_13842,N_12678);
xnor U18563 (N_18563,N_12323,N_15650);
nand U18564 (N_18564,N_13026,N_12510);
or U18565 (N_18565,N_15247,N_15792);
and U18566 (N_18566,N_15772,N_13136);
nor U18567 (N_18567,N_14388,N_12702);
nand U18568 (N_18568,N_13754,N_14474);
and U18569 (N_18569,N_15959,N_13476);
nor U18570 (N_18570,N_12692,N_12919);
nor U18571 (N_18571,N_12875,N_12574);
xnor U18572 (N_18572,N_12260,N_15033);
nor U18573 (N_18573,N_12996,N_14265);
nand U18574 (N_18574,N_14222,N_15196);
and U18575 (N_18575,N_12720,N_15234);
and U18576 (N_18576,N_15214,N_13760);
or U18577 (N_18577,N_12057,N_13780);
or U18578 (N_18578,N_12728,N_13451);
and U18579 (N_18579,N_13215,N_12349);
xnor U18580 (N_18580,N_12419,N_12661);
nand U18581 (N_18581,N_14615,N_15227);
xnor U18582 (N_18582,N_15900,N_15233);
or U18583 (N_18583,N_12689,N_12313);
xnor U18584 (N_18584,N_14905,N_15515);
and U18585 (N_18585,N_13713,N_14645);
nor U18586 (N_18586,N_14165,N_14033);
or U18587 (N_18587,N_14507,N_12825);
nand U18588 (N_18588,N_15500,N_14754);
nand U18589 (N_18589,N_13758,N_13458);
nand U18590 (N_18590,N_15806,N_13343);
xor U18591 (N_18591,N_12475,N_12571);
and U18592 (N_18592,N_14187,N_12101);
and U18593 (N_18593,N_15669,N_12364);
xnor U18594 (N_18594,N_15022,N_12191);
or U18595 (N_18595,N_12137,N_12703);
nor U18596 (N_18596,N_14151,N_15912);
nor U18597 (N_18597,N_13079,N_12147);
and U18598 (N_18598,N_13613,N_13293);
nand U18599 (N_18599,N_15079,N_12305);
xnor U18600 (N_18600,N_14347,N_13143);
and U18601 (N_18601,N_14215,N_13064);
xnor U18602 (N_18602,N_12539,N_15646);
or U18603 (N_18603,N_14555,N_12337);
xor U18604 (N_18604,N_12671,N_14488);
and U18605 (N_18605,N_12544,N_12839);
nor U18606 (N_18606,N_15893,N_12571);
xnor U18607 (N_18607,N_14669,N_15324);
nor U18608 (N_18608,N_14993,N_13490);
xnor U18609 (N_18609,N_15833,N_14013);
or U18610 (N_18610,N_14166,N_13339);
or U18611 (N_18611,N_12431,N_13948);
xor U18612 (N_18612,N_12971,N_12052);
xnor U18613 (N_18613,N_14832,N_13991);
nand U18614 (N_18614,N_12658,N_14184);
or U18615 (N_18615,N_12700,N_13993);
nor U18616 (N_18616,N_12599,N_12187);
nor U18617 (N_18617,N_12528,N_13330);
nand U18618 (N_18618,N_15062,N_14476);
nor U18619 (N_18619,N_13038,N_14068);
nand U18620 (N_18620,N_15936,N_13950);
or U18621 (N_18621,N_14512,N_15321);
nand U18622 (N_18622,N_13162,N_12132);
nor U18623 (N_18623,N_15807,N_12302);
and U18624 (N_18624,N_12564,N_12161);
or U18625 (N_18625,N_14400,N_13356);
or U18626 (N_18626,N_12222,N_13263);
or U18627 (N_18627,N_13004,N_13761);
and U18628 (N_18628,N_13467,N_12067);
nor U18629 (N_18629,N_13190,N_14536);
nand U18630 (N_18630,N_12972,N_14694);
nor U18631 (N_18631,N_12279,N_14318);
nor U18632 (N_18632,N_13256,N_13350);
and U18633 (N_18633,N_13272,N_13646);
nor U18634 (N_18634,N_14487,N_12054);
nor U18635 (N_18635,N_14974,N_15770);
or U18636 (N_18636,N_12309,N_15385);
nand U18637 (N_18637,N_15209,N_13131);
nor U18638 (N_18638,N_13643,N_15975);
nor U18639 (N_18639,N_13050,N_13325);
or U18640 (N_18640,N_13805,N_12612);
xnor U18641 (N_18641,N_14674,N_14398);
and U18642 (N_18642,N_14247,N_14609);
xor U18643 (N_18643,N_14053,N_13492);
nor U18644 (N_18644,N_12430,N_13608);
nand U18645 (N_18645,N_13427,N_14992);
nand U18646 (N_18646,N_14498,N_15058);
nand U18647 (N_18647,N_15521,N_13715);
and U18648 (N_18648,N_13453,N_15093);
or U18649 (N_18649,N_15447,N_15810);
nor U18650 (N_18650,N_12803,N_12424);
and U18651 (N_18651,N_13650,N_12388);
or U18652 (N_18652,N_15398,N_12411);
nand U18653 (N_18653,N_13555,N_14661);
xnor U18654 (N_18654,N_14120,N_15835);
nor U18655 (N_18655,N_15329,N_12158);
nor U18656 (N_18656,N_15841,N_15205);
and U18657 (N_18657,N_13135,N_12313);
nor U18658 (N_18658,N_14209,N_13890);
xor U18659 (N_18659,N_14676,N_14536);
or U18660 (N_18660,N_15182,N_15198);
nand U18661 (N_18661,N_15419,N_14086);
and U18662 (N_18662,N_12738,N_12138);
xnor U18663 (N_18663,N_14374,N_13928);
or U18664 (N_18664,N_15501,N_14821);
and U18665 (N_18665,N_14256,N_14770);
nand U18666 (N_18666,N_15267,N_15966);
and U18667 (N_18667,N_13743,N_15497);
and U18668 (N_18668,N_15521,N_14386);
and U18669 (N_18669,N_14163,N_12617);
nand U18670 (N_18670,N_14547,N_15429);
nand U18671 (N_18671,N_15317,N_15096);
xnor U18672 (N_18672,N_15833,N_14129);
xor U18673 (N_18673,N_14587,N_12177);
nand U18674 (N_18674,N_15777,N_14675);
xnor U18675 (N_18675,N_12548,N_14621);
xor U18676 (N_18676,N_13977,N_15326);
xor U18677 (N_18677,N_14753,N_14841);
nor U18678 (N_18678,N_13772,N_14971);
or U18679 (N_18679,N_12636,N_13277);
xor U18680 (N_18680,N_14569,N_13230);
nand U18681 (N_18681,N_12786,N_13760);
nor U18682 (N_18682,N_15887,N_13889);
and U18683 (N_18683,N_13488,N_14461);
xnor U18684 (N_18684,N_12777,N_13414);
nand U18685 (N_18685,N_12501,N_15019);
nand U18686 (N_18686,N_12331,N_13556);
or U18687 (N_18687,N_14552,N_12210);
nor U18688 (N_18688,N_15166,N_13737);
nor U18689 (N_18689,N_15934,N_14374);
and U18690 (N_18690,N_15759,N_15910);
xnor U18691 (N_18691,N_12469,N_15895);
and U18692 (N_18692,N_14082,N_13939);
nor U18693 (N_18693,N_13945,N_13218);
xnor U18694 (N_18694,N_14134,N_12761);
or U18695 (N_18695,N_14946,N_13523);
and U18696 (N_18696,N_15222,N_13985);
xnor U18697 (N_18697,N_15348,N_12785);
or U18698 (N_18698,N_15110,N_15129);
or U18699 (N_18699,N_15796,N_14649);
and U18700 (N_18700,N_14026,N_15048);
xor U18701 (N_18701,N_15161,N_12790);
nor U18702 (N_18702,N_13109,N_15247);
nor U18703 (N_18703,N_13318,N_15944);
xnor U18704 (N_18704,N_13608,N_15354);
or U18705 (N_18705,N_14568,N_13081);
nand U18706 (N_18706,N_15170,N_14839);
xor U18707 (N_18707,N_13807,N_12229);
and U18708 (N_18708,N_15209,N_13674);
nand U18709 (N_18709,N_13143,N_13337);
and U18710 (N_18710,N_12617,N_13804);
or U18711 (N_18711,N_14122,N_12544);
nor U18712 (N_18712,N_14085,N_12242);
nor U18713 (N_18713,N_15964,N_13764);
xnor U18714 (N_18714,N_12010,N_12330);
nand U18715 (N_18715,N_14177,N_13062);
xor U18716 (N_18716,N_15955,N_12395);
xnor U18717 (N_18717,N_15761,N_12582);
xnor U18718 (N_18718,N_12242,N_14345);
nor U18719 (N_18719,N_14969,N_15982);
and U18720 (N_18720,N_12629,N_13905);
and U18721 (N_18721,N_14010,N_15831);
nand U18722 (N_18722,N_14231,N_14912);
or U18723 (N_18723,N_15502,N_14915);
or U18724 (N_18724,N_15796,N_13600);
xor U18725 (N_18725,N_15415,N_15221);
nand U18726 (N_18726,N_15382,N_14904);
and U18727 (N_18727,N_13072,N_12352);
nand U18728 (N_18728,N_13093,N_13741);
nor U18729 (N_18729,N_14785,N_14515);
nor U18730 (N_18730,N_13358,N_13208);
nand U18731 (N_18731,N_12431,N_15195);
nor U18732 (N_18732,N_14274,N_13245);
nand U18733 (N_18733,N_12289,N_12893);
xnor U18734 (N_18734,N_14802,N_14672);
and U18735 (N_18735,N_13288,N_14844);
nand U18736 (N_18736,N_14828,N_13112);
nor U18737 (N_18737,N_15607,N_12506);
nand U18738 (N_18738,N_15176,N_13880);
xor U18739 (N_18739,N_14779,N_13126);
or U18740 (N_18740,N_12763,N_15617);
or U18741 (N_18741,N_15652,N_15435);
nand U18742 (N_18742,N_12669,N_13775);
xnor U18743 (N_18743,N_12131,N_14950);
nand U18744 (N_18744,N_15175,N_12977);
nand U18745 (N_18745,N_15142,N_13344);
or U18746 (N_18746,N_12870,N_13176);
nor U18747 (N_18747,N_15748,N_15409);
xor U18748 (N_18748,N_12815,N_15242);
xnor U18749 (N_18749,N_13091,N_15891);
xnor U18750 (N_18750,N_13368,N_14133);
nand U18751 (N_18751,N_15999,N_15534);
nand U18752 (N_18752,N_12843,N_13061);
and U18753 (N_18753,N_13949,N_14832);
xnor U18754 (N_18754,N_12079,N_14965);
or U18755 (N_18755,N_13024,N_12866);
or U18756 (N_18756,N_15380,N_14228);
nand U18757 (N_18757,N_14542,N_14933);
nor U18758 (N_18758,N_14058,N_14561);
and U18759 (N_18759,N_15365,N_14828);
nor U18760 (N_18760,N_12773,N_12595);
nor U18761 (N_18761,N_15065,N_13156);
and U18762 (N_18762,N_14594,N_12412);
and U18763 (N_18763,N_13395,N_13228);
nand U18764 (N_18764,N_13716,N_14198);
xnor U18765 (N_18765,N_14483,N_15373);
and U18766 (N_18766,N_13734,N_13876);
nor U18767 (N_18767,N_15598,N_12587);
or U18768 (N_18768,N_14328,N_12348);
xor U18769 (N_18769,N_14686,N_15099);
nor U18770 (N_18770,N_15776,N_14828);
or U18771 (N_18771,N_15529,N_13503);
and U18772 (N_18772,N_12268,N_14652);
nand U18773 (N_18773,N_15022,N_15631);
and U18774 (N_18774,N_14769,N_15615);
xnor U18775 (N_18775,N_15157,N_14274);
and U18776 (N_18776,N_15131,N_14926);
xor U18777 (N_18777,N_15632,N_12460);
nor U18778 (N_18778,N_13586,N_15682);
and U18779 (N_18779,N_12949,N_13928);
xor U18780 (N_18780,N_12085,N_15060);
and U18781 (N_18781,N_15638,N_12765);
and U18782 (N_18782,N_15264,N_12628);
nor U18783 (N_18783,N_13000,N_13660);
or U18784 (N_18784,N_13400,N_12396);
nand U18785 (N_18785,N_15395,N_13801);
and U18786 (N_18786,N_15234,N_14475);
and U18787 (N_18787,N_13752,N_12093);
nand U18788 (N_18788,N_13561,N_15236);
xnor U18789 (N_18789,N_14112,N_13993);
or U18790 (N_18790,N_12363,N_14313);
nand U18791 (N_18791,N_13627,N_13536);
nand U18792 (N_18792,N_12482,N_14779);
nor U18793 (N_18793,N_14136,N_12362);
xor U18794 (N_18794,N_14447,N_12454);
or U18795 (N_18795,N_15481,N_15660);
nor U18796 (N_18796,N_12113,N_13327);
xnor U18797 (N_18797,N_13379,N_15565);
and U18798 (N_18798,N_14774,N_15033);
nor U18799 (N_18799,N_12802,N_15286);
nor U18800 (N_18800,N_13132,N_14586);
nand U18801 (N_18801,N_13750,N_13224);
xor U18802 (N_18802,N_15517,N_15346);
xor U18803 (N_18803,N_15879,N_12675);
xor U18804 (N_18804,N_13128,N_14825);
or U18805 (N_18805,N_12137,N_12219);
or U18806 (N_18806,N_12374,N_14215);
xor U18807 (N_18807,N_15103,N_15813);
or U18808 (N_18808,N_15844,N_15551);
or U18809 (N_18809,N_14816,N_12944);
nor U18810 (N_18810,N_12532,N_15240);
or U18811 (N_18811,N_13911,N_12914);
nand U18812 (N_18812,N_15789,N_15339);
nor U18813 (N_18813,N_12610,N_12377);
xor U18814 (N_18814,N_14597,N_12314);
and U18815 (N_18815,N_13583,N_13135);
nand U18816 (N_18816,N_13690,N_12838);
nor U18817 (N_18817,N_12231,N_12138);
or U18818 (N_18818,N_13547,N_13750);
and U18819 (N_18819,N_13295,N_14108);
and U18820 (N_18820,N_14694,N_12661);
or U18821 (N_18821,N_15783,N_13460);
or U18822 (N_18822,N_13080,N_14379);
nor U18823 (N_18823,N_14009,N_13527);
and U18824 (N_18824,N_14304,N_15516);
nor U18825 (N_18825,N_13816,N_13446);
nor U18826 (N_18826,N_13215,N_13533);
xor U18827 (N_18827,N_12470,N_13129);
or U18828 (N_18828,N_15608,N_13692);
nor U18829 (N_18829,N_13857,N_12992);
and U18830 (N_18830,N_14425,N_14119);
nand U18831 (N_18831,N_14088,N_14926);
nor U18832 (N_18832,N_13539,N_14621);
xnor U18833 (N_18833,N_12370,N_14524);
xnor U18834 (N_18834,N_14756,N_13160);
xor U18835 (N_18835,N_14071,N_13162);
and U18836 (N_18836,N_12615,N_13625);
nand U18837 (N_18837,N_12715,N_12853);
xnor U18838 (N_18838,N_12649,N_15351);
and U18839 (N_18839,N_12620,N_15498);
nor U18840 (N_18840,N_15714,N_14542);
nand U18841 (N_18841,N_12376,N_14745);
or U18842 (N_18842,N_12609,N_13353);
nand U18843 (N_18843,N_12706,N_12122);
nor U18844 (N_18844,N_14115,N_15392);
or U18845 (N_18845,N_13931,N_14723);
xnor U18846 (N_18846,N_14757,N_12184);
nor U18847 (N_18847,N_15282,N_12260);
nor U18848 (N_18848,N_13906,N_15850);
or U18849 (N_18849,N_14937,N_14973);
nand U18850 (N_18850,N_14213,N_14694);
xor U18851 (N_18851,N_12037,N_12558);
and U18852 (N_18852,N_13817,N_14907);
nor U18853 (N_18853,N_13996,N_12566);
xnor U18854 (N_18854,N_12086,N_13784);
or U18855 (N_18855,N_12768,N_12414);
and U18856 (N_18856,N_15791,N_14664);
or U18857 (N_18857,N_12679,N_14257);
or U18858 (N_18858,N_14776,N_13419);
or U18859 (N_18859,N_14180,N_13628);
and U18860 (N_18860,N_14150,N_12134);
nand U18861 (N_18861,N_15669,N_12413);
nand U18862 (N_18862,N_12950,N_15885);
and U18863 (N_18863,N_12592,N_13128);
nor U18864 (N_18864,N_14271,N_15311);
and U18865 (N_18865,N_12882,N_14833);
nand U18866 (N_18866,N_12727,N_14048);
nor U18867 (N_18867,N_13226,N_13659);
and U18868 (N_18868,N_13638,N_12926);
nand U18869 (N_18869,N_15971,N_12174);
nand U18870 (N_18870,N_12093,N_13974);
nand U18871 (N_18871,N_13247,N_13626);
nor U18872 (N_18872,N_15878,N_14469);
and U18873 (N_18873,N_14243,N_14720);
nor U18874 (N_18874,N_14773,N_12449);
nand U18875 (N_18875,N_15857,N_15311);
or U18876 (N_18876,N_12131,N_14987);
nand U18877 (N_18877,N_13038,N_12434);
or U18878 (N_18878,N_14416,N_15155);
nand U18879 (N_18879,N_14001,N_13619);
or U18880 (N_18880,N_14336,N_15666);
nor U18881 (N_18881,N_13308,N_15922);
nand U18882 (N_18882,N_13340,N_14463);
and U18883 (N_18883,N_15744,N_12208);
xnor U18884 (N_18884,N_13621,N_15139);
xnor U18885 (N_18885,N_12313,N_15039);
or U18886 (N_18886,N_12557,N_14648);
nand U18887 (N_18887,N_14430,N_12083);
or U18888 (N_18888,N_13235,N_15417);
or U18889 (N_18889,N_13194,N_13429);
nor U18890 (N_18890,N_13914,N_15897);
and U18891 (N_18891,N_12049,N_14034);
and U18892 (N_18892,N_15131,N_15824);
or U18893 (N_18893,N_12830,N_12096);
and U18894 (N_18894,N_14575,N_15292);
xor U18895 (N_18895,N_14178,N_15728);
and U18896 (N_18896,N_12772,N_12858);
or U18897 (N_18897,N_12239,N_13795);
nand U18898 (N_18898,N_14750,N_14918);
xnor U18899 (N_18899,N_15223,N_13919);
xnor U18900 (N_18900,N_12603,N_15154);
xnor U18901 (N_18901,N_14755,N_12486);
nor U18902 (N_18902,N_15551,N_12558);
xor U18903 (N_18903,N_15794,N_15962);
and U18904 (N_18904,N_15594,N_14945);
and U18905 (N_18905,N_12940,N_14739);
or U18906 (N_18906,N_12899,N_13564);
nand U18907 (N_18907,N_13571,N_12249);
nand U18908 (N_18908,N_15852,N_12214);
xnor U18909 (N_18909,N_14980,N_13596);
nand U18910 (N_18910,N_14056,N_15577);
nor U18911 (N_18911,N_13538,N_15562);
nor U18912 (N_18912,N_12175,N_14551);
or U18913 (N_18913,N_13420,N_13608);
or U18914 (N_18914,N_14345,N_12414);
nor U18915 (N_18915,N_13411,N_14603);
nor U18916 (N_18916,N_14909,N_14380);
nand U18917 (N_18917,N_14256,N_12607);
nor U18918 (N_18918,N_13638,N_15894);
or U18919 (N_18919,N_15270,N_15535);
nand U18920 (N_18920,N_12590,N_14426);
xor U18921 (N_18921,N_12790,N_14295);
or U18922 (N_18922,N_14596,N_14094);
and U18923 (N_18923,N_13247,N_12630);
nor U18924 (N_18924,N_13963,N_12007);
xor U18925 (N_18925,N_15216,N_13616);
nor U18926 (N_18926,N_14263,N_15690);
nand U18927 (N_18927,N_15986,N_14864);
nand U18928 (N_18928,N_15779,N_12913);
xnor U18929 (N_18929,N_13428,N_12708);
xnor U18930 (N_18930,N_15184,N_14144);
xnor U18931 (N_18931,N_15124,N_15669);
xor U18932 (N_18932,N_12193,N_15551);
nand U18933 (N_18933,N_14341,N_13879);
nand U18934 (N_18934,N_14934,N_15346);
nor U18935 (N_18935,N_15893,N_15292);
xor U18936 (N_18936,N_15160,N_15248);
and U18937 (N_18937,N_15407,N_12418);
nand U18938 (N_18938,N_14376,N_13951);
and U18939 (N_18939,N_14485,N_15449);
nand U18940 (N_18940,N_13088,N_13905);
or U18941 (N_18941,N_15401,N_15949);
or U18942 (N_18942,N_12357,N_15712);
xnor U18943 (N_18943,N_12689,N_14979);
nand U18944 (N_18944,N_14212,N_14960);
or U18945 (N_18945,N_15050,N_15004);
or U18946 (N_18946,N_12525,N_12926);
xor U18947 (N_18947,N_15545,N_12830);
nor U18948 (N_18948,N_14447,N_15246);
or U18949 (N_18949,N_14235,N_13721);
or U18950 (N_18950,N_14641,N_14449);
nor U18951 (N_18951,N_15265,N_12734);
or U18952 (N_18952,N_13210,N_13142);
nor U18953 (N_18953,N_14480,N_13892);
nand U18954 (N_18954,N_12562,N_15980);
xor U18955 (N_18955,N_12442,N_12347);
nand U18956 (N_18956,N_14884,N_13580);
and U18957 (N_18957,N_14287,N_15228);
and U18958 (N_18958,N_12421,N_14875);
xnor U18959 (N_18959,N_13499,N_12091);
nand U18960 (N_18960,N_14310,N_15020);
xnor U18961 (N_18961,N_12177,N_15021);
nor U18962 (N_18962,N_14081,N_13789);
nand U18963 (N_18963,N_15843,N_12676);
or U18964 (N_18964,N_13027,N_13743);
xnor U18965 (N_18965,N_14645,N_12554);
xor U18966 (N_18966,N_15701,N_12358);
and U18967 (N_18967,N_15055,N_14647);
nand U18968 (N_18968,N_15364,N_15955);
and U18969 (N_18969,N_14877,N_12652);
nand U18970 (N_18970,N_12260,N_12187);
or U18971 (N_18971,N_14773,N_12716);
xnor U18972 (N_18972,N_12317,N_14185);
nand U18973 (N_18973,N_13132,N_14255);
nand U18974 (N_18974,N_14445,N_13527);
xnor U18975 (N_18975,N_15343,N_13891);
xor U18976 (N_18976,N_15604,N_12216);
and U18977 (N_18977,N_15475,N_15154);
xor U18978 (N_18978,N_12561,N_14158);
xnor U18979 (N_18979,N_13484,N_14084);
nand U18980 (N_18980,N_13076,N_12457);
and U18981 (N_18981,N_14270,N_15150);
or U18982 (N_18982,N_15925,N_12692);
and U18983 (N_18983,N_15965,N_15661);
or U18984 (N_18984,N_12862,N_12977);
nor U18985 (N_18985,N_13228,N_13953);
nand U18986 (N_18986,N_15031,N_14728);
nor U18987 (N_18987,N_14601,N_13652);
and U18988 (N_18988,N_14782,N_15399);
nor U18989 (N_18989,N_15089,N_13255);
nand U18990 (N_18990,N_12406,N_12109);
nand U18991 (N_18991,N_15383,N_14223);
and U18992 (N_18992,N_13792,N_12330);
nor U18993 (N_18993,N_12704,N_13098);
nor U18994 (N_18994,N_12499,N_12772);
nand U18995 (N_18995,N_14364,N_15114);
xor U18996 (N_18996,N_12240,N_14484);
or U18997 (N_18997,N_12330,N_14667);
and U18998 (N_18998,N_15784,N_14665);
and U18999 (N_18999,N_12415,N_12139);
nor U19000 (N_19000,N_12054,N_12400);
nand U19001 (N_19001,N_12205,N_14673);
and U19002 (N_19002,N_13201,N_15671);
xor U19003 (N_19003,N_12501,N_15550);
nand U19004 (N_19004,N_14125,N_14569);
or U19005 (N_19005,N_12720,N_13899);
or U19006 (N_19006,N_13494,N_14767);
nor U19007 (N_19007,N_12831,N_13648);
nand U19008 (N_19008,N_13350,N_14922);
and U19009 (N_19009,N_14354,N_14280);
nor U19010 (N_19010,N_13533,N_13335);
nand U19011 (N_19011,N_13822,N_13249);
nand U19012 (N_19012,N_15160,N_15274);
nor U19013 (N_19013,N_14186,N_14535);
or U19014 (N_19014,N_12674,N_15544);
and U19015 (N_19015,N_12865,N_13766);
nor U19016 (N_19016,N_12417,N_14275);
or U19017 (N_19017,N_14277,N_13020);
and U19018 (N_19018,N_14231,N_13829);
xor U19019 (N_19019,N_12497,N_15475);
or U19020 (N_19020,N_14428,N_13940);
and U19021 (N_19021,N_13138,N_12927);
and U19022 (N_19022,N_12038,N_14996);
or U19023 (N_19023,N_14417,N_15709);
nand U19024 (N_19024,N_13476,N_15647);
and U19025 (N_19025,N_15946,N_14399);
and U19026 (N_19026,N_12362,N_13813);
nor U19027 (N_19027,N_13485,N_12606);
xnor U19028 (N_19028,N_12054,N_14471);
nor U19029 (N_19029,N_15814,N_15043);
nand U19030 (N_19030,N_14237,N_13156);
xnor U19031 (N_19031,N_15553,N_13081);
xor U19032 (N_19032,N_14790,N_12819);
nand U19033 (N_19033,N_13314,N_15576);
or U19034 (N_19034,N_12002,N_12222);
and U19035 (N_19035,N_13422,N_13081);
nor U19036 (N_19036,N_15378,N_15526);
nand U19037 (N_19037,N_14523,N_13892);
and U19038 (N_19038,N_14043,N_13431);
or U19039 (N_19039,N_12955,N_15662);
nor U19040 (N_19040,N_12414,N_14014);
and U19041 (N_19041,N_12166,N_13963);
or U19042 (N_19042,N_12910,N_12233);
nand U19043 (N_19043,N_14512,N_12313);
or U19044 (N_19044,N_15631,N_14073);
nand U19045 (N_19045,N_15517,N_12726);
and U19046 (N_19046,N_12859,N_14587);
nor U19047 (N_19047,N_12010,N_13477);
nand U19048 (N_19048,N_15697,N_14984);
nand U19049 (N_19049,N_14871,N_12699);
and U19050 (N_19050,N_12460,N_14222);
nand U19051 (N_19051,N_14907,N_14235);
nand U19052 (N_19052,N_14537,N_15781);
nand U19053 (N_19053,N_12173,N_12207);
and U19054 (N_19054,N_12362,N_15665);
nor U19055 (N_19055,N_14442,N_14002);
xnor U19056 (N_19056,N_14244,N_14567);
and U19057 (N_19057,N_13233,N_12361);
and U19058 (N_19058,N_13105,N_12565);
xor U19059 (N_19059,N_14640,N_13599);
xnor U19060 (N_19060,N_14791,N_13535);
nor U19061 (N_19061,N_14524,N_13297);
and U19062 (N_19062,N_15600,N_14147);
and U19063 (N_19063,N_12163,N_12278);
and U19064 (N_19064,N_12993,N_12117);
xor U19065 (N_19065,N_14043,N_15252);
xor U19066 (N_19066,N_12213,N_14872);
nand U19067 (N_19067,N_15930,N_14037);
nand U19068 (N_19068,N_15080,N_14187);
nor U19069 (N_19069,N_13566,N_15865);
xor U19070 (N_19070,N_15179,N_14482);
and U19071 (N_19071,N_13055,N_14282);
nor U19072 (N_19072,N_15681,N_14865);
nand U19073 (N_19073,N_12331,N_15443);
nor U19074 (N_19074,N_12311,N_12091);
nand U19075 (N_19075,N_12860,N_15537);
xor U19076 (N_19076,N_15994,N_15912);
and U19077 (N_19077,N_13433,N_15319);
and U19078 (N_19078,N_14706,N_14149);
xor U19079 (N_19079,N_13388,N_14904);
nand U19080 (N_19080,N_14608,N_14478);
nor U19081 (N_19081,N_14830,N_13970);
or U19082 (N_19082,N_13570,N_12312);
nand U19083 (N_19083,N_14577,N_12945);
or U19084 (N_19084,N_15250,N_14579);
or U19085 (N_19085,N_13412,N_14823);
nand U19086 (N_19086,N_14473,N_13937);
and U19087 (N_19087,N_13753,N_15669);
nor U19088 (N_19088,N_12007,N_12688);
nor U19089 (N_19089,N_13001,N_12319);
and U19090 (N_19090,N_14379,N_15423);
nor U19091 (N_19091,N_15364,N_14937);
nor U19092 (N_19092,N_13362,N_15203);
xnor U19093 (N_19093,N_15957,N_15975);
and U19094 (N_19094,N_12502,N_14094);
or U19095 (N_19095,N_13212,N_14217);
nand U19096 (N_19096,N_15304,N_15877);
nor U19097 (N_19097,N_12990,N_13243);
or U19098 (N_19098,N_12266,N_15011);
or U19099 (N_19099,N_13420,N_14487);
and U19100 (N_19100,N_15343,N_13435);
nand U19101 (N_19101,N_15915,N_13381);
nor U19102 (N_19102,N_12374,N_15619);
and U19103 (N_19103,N_14262,N_12394);
or U19104 (N_19104,N_12649,N_12038);
nand U19105 (N_19105,N_12101,N_12447);
xnor U19106 (N_19106,N_13406,N_14733);
nor U19107 (N_19107,N_14360,N_13300);
xor U19108 (N_19108,N_15024,N_14071);
and U19109 (N_19109,N_13850,N_12482);
or U19110 (N_19110,N_12440,N_12325);
or U19111 (N_19111,N_14062,N_15035);
and U19112 (N_19112,N_12560,N_12591);
nor U19113 (N_19113,N_12536,N_13241);
and U19114 (N_19114,N_12592,N_15794);
and U19115 (N_19115,N_13216,N_12689);
or U19116 (N_19116,N_15020,N_13194);
or U19117 (N_19117,N_14157,N_15107);
nand U19118 (N_19118,N_12248,N_12680);
or U19119 (N_19119,N_14726,N_12549);
nand U19120 (N_19120,N_14322,N_13352);
nand U19121 (N_19121,N_15865,N_12889);
or U19122 (N_19122,N_13639,N_13859);
nand U19123 (N_19123,N_13858,N_12072);
and U19124 (N_19124,N_15439,N_13031);
xnor U19125 (N_19125,N_15917,N_15685);
or U19126 (N_19126,N_14381,N_13327);
or U19127 (N_19127,N_13407,N_14020);
xnor U19128 (N_19128,N_15023,N_14029);
xor U19129 (N_19129,N_15416,N_12349);
nand U19130 (N_19130,N_13691,N_14830);
nand U19131 (N_19131,N_13472,N_12588);
nor U19132 (N_19132,N_15966,N_12223);
nor U19133 (N_19133,N_13844,N_14432);
and U19134 (N_19134,N_12380,N_14770);
and U19135 (N_19135,N_13928,N_15306);
xnor U19136 (N_19136,N_15696,N_12860);
xor U19137 (N_19137,N_14862,N_14509);
nor U19138 (N_19138,N_13796,N_15638);
xor U19139 (N_19139,N_14930,N_15108);
or U19140 (N_19140,N_15074,N_12758);
nand U19141 (N_19141,N_14302,N_14292);
nor U19142 (N_19142,N_15594,N_14411);
nand U19143 (N_19143,N_14662,N_14385);
or U19144 (N_19144,N_14019,N_12464);
or U19145 (N_19145,N_12669,N_12364);
xor U19146 (N_19146,N_15144,N_15238);
nor U19147 (N_19147,N_13498,N_12528);
nand U19148 (N_19148,N_14166,N_13890);
or U19149 (N_19149,N_12715,N_12088);
and U19150 (N_19150,N_15172,N_15798);
nor U19151 (N_19151,N_15532,N_14941);
and U19152 (N_19152,N_13433,N_15895);
nor U19153 (N_19153,N_13533,N_15138);
and U19154 (N_19154,N_14471,N_14483);
nand U19155 (N_19155,N_14872,N_12332);
and U19156 (N_19156,N_12765,N_14440);
or U19157 (N_19157,N_14148,N_14895);
or U19158 (N_19158,N_13744,N_15833);
or U19159 (N_19159,N_14704,N_14414);
or U19160 (N_19160,N_13245,N_14228);
and U19161 (N_19161,N_13338,N_12221);
and U19162 (N_19162,N_12454,N_13973);
nand U19163 (N_19163,N_14543,N_14431);
nor U19164 (N_19164,N_15737,N_15991);
or U19165 (N_19165,N_14738,N_13499);
or U19166 (N_19166,N_12595,N_14980);
and U19167 (N_19167,N_15348,N_14976);
nand U19168 (N_19168,N_13637,N_15187);
or U19169 (N_19169,N_13078,N_13812);
nand U19170 (N_19170,N_13526,N_14919);
nand U19171 (N_19171,N_12874,N_13459);
nor U19172 (N_19172,N_12536,N_13020);
nor U19173 (N_19173,N_13182,N_13350);
xnor U19174 (N_19174,N_12759,N_13115);
and U19175 (N_19175,N_12880,N_14546);
nor U19176 (N_19176,N_12232,N_14397);
xnor U19177 (N_19177,N_12297,N_13857);
nand U19178 (N_19178,N_15915,N_13012);
or U19179 (N_19179,N_15430,N_15299);
and U19180 (N_19180,N_15515,N_13764);
or U19181 (N_19181,N_14397,N_12551);
or U19182 (N_19182,N_15407,N_14892);
and U19183 (N_19183,N_15554,N_15539);
nand U19184 (N_19184,N_13159,N_12139);
or U19185 (N_19185,N_14293,N_13083);
and U19186 (N_19186,N_12754,N_13675);
and U19187 (N_19187,N_14993,N_14248);
nor U19188 (N_19188,N_13460,N_13873);
and U19189 (N_19189,N_14381,N_14541);
nor U19190 (N_19190,N_12695,N_14788);
xnor U19191 (N_19191,N_14584,N_12017);
nand U19192 (N_19192,N_13931,N_12730);
nor U19193 (N_19193,N_14541,N_13345);
nand U19194 (N_19194,N_12800,N_14280);
xnor U19195 (N_19195,N_13653,N_12907);
and U19196 (N_19196,N_13691,N_15112);
xnor U19197 (N_19197,N_15750,N_14337);
xnor U19198 (N_19198,N_12515,N_15799);
xnor U19199 (N_19199,N_13548,N_15011);
or U19200 (N_19200,N_12815,N_14170);
or U19201 (N_19201,N_13816,N_13440);
or U19202 (N_19202,N_12920,N_13048);
and U19203 (N_19203,N_14622,N_15757);
nand U19204 (N_19204,N_15032,N_15135);
nand U19205 (N_19205,N_15960,N_14655);
nor U19206 (N_19206,N_15818,N_15858);
nor U19207 (N_19207,N_15611,N_15516);
and U19208 (N_19208,N_12967,N_14121);
nor U19209 (N_19209,N_12394,N_12595);
nand U19210 (N_19210,N_14264,N_15398);
or U19211 (N_19211,N_12455,N_14048);
or U19212 (N_19212,N_15666,N_13943);
or U19213 (N_19213,N_14876,N_12689);
xnor U19214 (N_19214,N_13053,N_15195);
nor U19215 (N_19215,N_14515,N_14257);
and U19216 (N_19216,N_14186,N_13532);
nand U19217 (N_19217,N_14940,N_15403);
and U19218 (N_19218,N_15379,N_12125);
xor U19219 (N_19219,N_12207,N_13651);
nand U19220 (N_19220,N_13625,N_12476);
or U19221 (N_19221,N_13821,N_12097);
nor U19222 (N_19222,N_12773,N_14017);
nand U19223 (N_19223,N_12528,N_13882);
and U19224 (N_19224,N_14997,N_14970);
nor U19225 (N_19225,N_12350,N_13341);
nor U19226 (N_19226,N_12784,N_14792);
xor U19227 (N_19227,N_13908,N_13918);
xor U19228 (N_19228,N_12944,N_15829);
and U19229 (N_19229,N_14739,N_15979);
nor U19230 (N_19230,N_14793,N_13607);
and U19231 (N_19231,N_13403,N_14159);
nor U19232 (N_19232,N_15844,N_13544);
nor U19233 (N_19233,N_12096,N_15013);
xnor U19234 (N_19234,N_14479,N_12631);
xnor U19235 (N_19235,N_14561,N_15485);
and U19236 (N_19236,N_15556,N_12883);
or U19237 (N_19237,N_15322,N_14273);
nand U19238 (N_19238,N_14406,N_12803);
or U19239 (N_19239,N_15091,N_13675);
xor U19240 (N_19240,N_14918,N_12059);
or U19241 (N_19241,N_12003,N_12396);
and U19242 (N_19242,N_14258,N_12529);
or U19243 (N_19243,N_13443,N_13577);
nor U19244 (N_19244,N_13351,N_13787);
and U19245 (N_19245,N_14042,N_14850);
and U19246 (N_19246,N_12788,N_12992);
and U19247 (N_19247,N_12067,N_15810);
or U19248 (N_19248,N_13281,N_14759);
xor U19249 (N_19249,N_12459,N_15157);
and U19250 (N_19250,N_14464,N_13318);
and U19251 (N_19251,N_13560,N_13122);
xnor U19252 (N_19252,N_15737,N_13111);
or U19253 (N_19253,N_14567,N_13970);
xor U19254 (N_19254,N_14928,N_13604);
and U19255 (N_19255,N_13351,N_14569);
nand U19256 (N_19256,N_15266,N_12606);
or U19257 (N_19257,N_13996,N_14337);
and U19258 (N_19258,N_13137,N_12089);
or U19259 (N_19259,N_12631,N_14672);
xor U19260 (N_19260,N_14280,N_15082);
xnor U19261 (N_19261,N_12696,N_14868);
xor U19262 (N_19262,N_14574,N_14365);
nand U19263 (N_19263,N_12794,N_13753);
nand U19264 (N_19264,N_12098,N_13257);
nor U19265 (N_19265,N_13806,N_12142);
nand U19266 (N_19266,N_12873,N_14537);
nor U19267 (N_19267,N_13419,N_13275);
xnor U19268 (N_19268,N_14556,N_14147);
and U19269 (N_19269,N_14336,N_14964);
and U19270 (N_19270,N_13293,N_14768);
or U19271 (N_19271,N_13077,N_12442);
nand U19272 (N_19272,N_13802,N_13663);
xnor U19273 (N_19273,N_14933,N_12204);
nand U19274 (N_19274,N_14754,N_15120);
nor U19275 (N_19275,N_12820,N_14060);
nor U19276 (N_19276,N_12930,N_12858);
nand U19277 (N_19277,N_14318,N_12878);
or U19278 (N_19278,N_12454,N_15369);
nor U19279 (N_19279,N_15306,N_13060);
nor U19280 (N_19280,N_15687,N_15956);
xor U19281 (N_19281,N_13546,N_13030);
or U19282 (N_19282,N_13499,N_14526);
or U19283 (N_19283,N_14980,N_14179);
xnor U19284 (N_19284,N_14454,N_13526);
nor U19285 (N_19285,N_13646,N_13608);
nand U19286 (N_19286,N_12345,N_13916);
xor U19287 (N_19287,N_13610,N_13216);
nor U19288 (N_19288,N_12582,N_15428);
and U19289 (N_19289,N_13314,N_15729);
nor U19290 (N_19290,N_13459,N_14067);
and U19291 (N_19291,N_12628,N_15607);
nor U19292 (N_19292,N_14182,N_14379);
or U19293 (N_19293,N_13104,N_13882);
xnor U19294 (N_19294,N_12896,N_15870);
nor U19295 (N_19295,N_13494,N_13988);
xor U19296 (N_19296,N_15054,N_14073);
or U19297 (N_19297,N_13963,N_14208);
or U19298 (N_19298,N_13184,N_15825);
nor U19299 (N_19299,N_13803,N_12028);
or U19300 (N_19300,N_13952,N_13588);
xnor U19301 (N_19301,N_12480,N_13415);
nor U19302 (N_19302,N_14005,N_15240);
or U19303 (N_19303,N_13754,N_15834);
xnor U19304 (N_19304,N_12748,N_13811);
nand U19305 (N_19305,N_14510,N_12389);
and U19306 (N_19306,N_13098,N_14413);
or U19307 (N_19307,N_13874,N_12517);
and U19308 (N_19308,N_13115,N_13645);
and U19309 (N_19309,N_12049,N_13026);
nor U19310 (N_19310,N_14176,N_15429);
nor U19311 (N_19311,N_14902,N_14016);
xnor U19312 (N_19312,N_14807,N_14809);
xor U19313 (N_19313,N_15355,N_15466);
or U19314 (N_19314,N_15346,N_12312);
nor U19315 (N_19315,N_14343,N_14036);
and U19316 (N_19316,N_12208,N_12561);
or U19317 (N_19317,N_14964,N_14389);
xnor U19318 (N_19318,N_15043,N_13075);
xnor U19319 (N_19319,N_13511,N_14787);
nor U19320 (N_19320,N_13723,N_15788);
nand U19321 (N_19321,N_14802,N_14139);
nand U19322 (N_19322,N_15379,N_12598);
or U19323 (N_19323,N_13688,N_15775);
or U19324 (N_19324,N_15067,N_15338);
nor U19325 (N_19325,N_15063,N_14958);
xor U19326 (N_19326,N_12825,N_12016);
nand U19327 (N_19327,N_14015,N_12598);
and U19328 (N_19328,N_13211,N_13396);
and U19329 (N_19329,N_13167,N_13534);
nor U19330 (N_19330,N_14024,N_13545);
or U19331 (N_19331,N_14793,N_13085);
nor U19332 (N_19332,N_12191,N_14489);
and U19333 (N_19333,N_12414,N_14982);
nand U19334 (N_19334,N_12641,N_12462);
and U19335 (N_19335,N_13688,N_12837);
xnor U19336 (N_19336,N_14251,N_13997);
and U19337 (N_19337,N_12166,N_13066);
nand U19338 (N_19338,N_15661,N_12418);
and U19339 (N_19339,N_15207,N_14586);
or U19340 (N_19340,N_12902,N_13940);
nand U19341 (N_19341,N_12003,N_12068);
xnor U19342 (N_19342,N_14995,N_13620);
nand U19343 (N_19343,N_14334,N_14972);
or U19344 (N_19344,N_15253,N_12668);
and U19345 (N_19345,N_13263,N_12000);
and U19346 (N_19346,N_15688,N_12921);
xnor U19347 (N_19347,N_13975,N_15066);
nor U19348 (N_19348,N_12220,N_15831);
nand U19349 (N_19349,N_13971,N_12863);
nor U19350 (N_19350,N_14305,N_12957);
or U19351 (N_19351,N_14732,N_13881);
xnor U19352 (N_19352,N_12532,N_14210);
nor U19353 (N_19353,N_15238,N_15402);
or U19354 (N_19354,N_14978,N_15443);
or U19355 (N_19355,N_15257,N_12558);
nand U19356 (N_19356,N_14609,N_14299);
nor U19357 (N_19357,N_12996,N_13748);
nand U19358 (N_19358,N_12736,N_12132);
nor U19359 (N_19359,N_12720,N_12126);
xor U19360 (N_19360,N_15512,N_14464);
nand U19361 (N_19361,N_14148,N_14286);
nor U19362 (N_19362,N_13254,N_15949);
and U19363 (N_19363,N_14444,N_13207);
nand U19364 (N_19364,N_12465,N_13216);
nand U19365 (N_19365,N_13622,N_15544);
nand U19366 (N_19366,N_15606,N_14980);
and U19367 (N_19367,N_15432,N_13212);
or U19368 (N_19368,N_12424,N_15116);
or U19369 (N_19369,N_15197,N_13387);
nor U19370 (N_19370,N_14915,N_14745);
nand U19371 (N_19371,N_13531,N_14574);
nand U19372 (N_19372,N_15015,N_15489);
or U19373 (N_19373,N_15061,N_14526);
and U19374 (N_19374,N_14407,N_13744);
nor U19375 (N_19375,N_15559,N_12772);
nand U19376 (N_19376,N_13240,N_12120);
nand U19377 (N_19377,N_14822,N_15438);
xnor U19378 (N_19378,N_12434,N_14090);
xor U19379 (N_19379,N_12215,N_14804);
nor U19380 (N_19380,N_12042,N_14800);
and U19381 (N_19381,N_12158,N_12371);
and U19382 (N_19382,N_14159,N_14867);
nand U19383 (N_19383,N_13212,N_14630);
nor U19384 (N_19384,N_15465,N_12839);
and U19385 (N_19385,N_12659,N_12114);
xnor U19386 (N_19386,N_13104,N_13739);
xnor U19387 (N_19387,N_12905,N_15271);
or U19388 (N_19388,N_14491,N_12165);
or U19389 (N_19389,N_13816,N_13318);
and U19390 (N_19390,N_14928,N_15308);
nor U19391 (N_19391,N_15934,N_15752);
and U19392 (N_19392,N_12128,N_12068);
nand U19393 (N_19393,N_14944,N_14499);
and U19394 (N_19394,N_14608,N_13543);
and U19395 (N_19395,N_13010,N_13800);
or U19396 (N_19396,N_15130,N_14330);
and U19397 (N_19397,N_15981,N_14267);
or U19398 (N_19398,N_14144,N_14430);
and U19399 (N_19399,N_14693,N_12352);
and U19400 (N_19400,N_14310,N_12950);
nand U19401 (N_19401,N_13737,N_13758);
xor U19402 (N_19402,N_13359,N_12257);
nor U19403 (N_19403,N_13775,N_13427);
nand U19404 (N_19404,N_13218,N_15852);
or U19405 (N_19405,N_14158,N_15811);
xnor U19406 (N_19406,N_12514,N_15275);
nand U19407 (N_19407,N_15188,N_12281);
and U19408 (N_19408,N_13488,N_15680);
and U19409 (N_19409,N_15359,N_12401);
nor U19410 (N_19410,N_15142,N_15999);
nor U19411 (N_19411,N_15916,N_13981);
nor U19412 (N_19412,N_12814,N_12712);
xnor U19413 (N_19413,N_15077,N_14410);
or U19414 (N_19414,N_12148,N_12695);
xnor U19415 (N_19415,N_14431,N_15355);
or U19416 (N_19416,N_13274,N_13723);
nand U19417 (N_19417,N_14950,N_15031);
xor U19418 (N_19418,N_12820,N_14385);
nand U19419 (N_19419,N_15458,N_15245);
nand U19420 (N_19420,N_13320,N_13520);
xnor U19421 (N_19421,N_14965,N_15473);
nor U19422 (N_19422,N_15050,N_15475);
and U19423 (N_19423,N_12879,N_15638);
xnor U19424 (N_19424,N_12858,N_12874);
or U19425 (N_19425,N_14914,N_15976);
xnor U19426 (N_19426,N_13959,N_12636);
xnor U19427 (N_19427,N_12461,N_15133);
or U19428 (N_19428,N_14993,N_12382);
or U19429 (N_19429,N_15877,N_14251);
nand U19430 (N_19430,N_15704,N_15665);
xor U19431 (N_19431,N_12674,N_15016);
or U19432 (N_19432,N_13012,N_13680);
nand U19433 (N_19433,N_13704,N_14869);
xor U19434 (N_19434,N_15672,N_15071);
or U19435 (N_19435,N_14199,N_12818);
or U19436 (N_19436,N_15994,N_14650);
nand U19437 (N_19437,N_14455,N_13162);
or U19438 (N_19438,N_15517,N_13813);
and U19439 (N_19439,N_14952,N_15493);
nor U19440 (N_19440,N_14775,N_13571);
or U19441 (N_19441,N_12263,N_15758);
xor U19442 (N_19442,N_13019,N_12355);
or U19443 (N_19443,N_12520,N_14620);
or U19444 (N_19444,N_14014,N_14004);
or U19445 (N_19445,N_15847,N_12988);
xnor U19446 (N_19446,N_13895,N_12310);
nand U19447 (N_19447,N_12577,N_13451);
nand U19448 (N_19448,N_13201,N_14615);
nor U19449 (N_19449,N_14389,N_13869);
or U19450 (N_19450,N_15936,N_13261);
and U19451 (N_19451,N_15976,N_13927);
and U19452 (N_19452,N_12034,N_15679);
nand U19453 (N_19453,N_15762,N_14729);
nor U19454 (N_19454,N_13562,N_15197);
xnor U19455 (N_19455,N_14030,N_12772);
and U19456 (N_19456,N_14769,N_13243);
and U19457 (N_19457,N_13696,N_15523);
or U19458 (N_19458,N_14229,N_12085);
and U19459 (N_19459,N_14733,N_13233);
and U19460 (N_19460,N_13295,N_15254);
and U19461 (N_19461,N_15485,N_15878);
and U19462 (N_19462,N_12702,N_15866);
or U19463 (N_19463,N_12280,N_13201);
nor U19464 (N_19464,N_12044,N_15583);
and U19465 (N_19465,N_13835,N_13451);
or U19466 (N_19466,N_13818,N_13676);
and U19467 (N_19467,N_15801,N_12592);
and U19468 (N_19468,N_14144,N_15844);
or U19469 (N_19469,N_15665,N_13577);
or U19470 (N_19470,N_12549,N_15727);
and U19471 (N_19471,N_15721,N_15210);
nand U19472 (N_19472,N_13702,N_12411);
and U19473 (N_19473,N_12188,N_14960);
nor U19474 (N_19474,N_15617,N_12128);
nor U19475 (N_19475,N_15356,N_12639);
nand U19476 (N_19476,N_13870,N_13872);
nor U19477 (N_19477,N_12311,N_14452);
nand U19478 (N_19478,N_15436,N_12871);
and U19479 (N_19479,N_12198,N_12115);
nor U19480 (N_19480,N_13947,N_13886);
or U19481 (N_19481,N_15246,N_14552);
nor U19482 (N_19482,N_14669,N_14950);
or U19483 (N_19483,N_14403,N_13040);
nor U19484 (N_19484,N_15328,N_13500);
or U19485 (N_19485,N_15711,N_15769);
and U19486 (N_19486,N_14104,N_12144);
nand U19487 (N_19487,N_12873,N_14494);
and U19488 (N_19488,N_14769,N_15422);
nand U19489 (N_19489,N_15771,N_12103);
and U19490 (N_19490,N_12911,N_12915);
or U19491 (N_19491,N_14720,N_14417);
xnor U19492 (N_19492,N_13095,N_13154);
nand U19493 (N_19493,N_13210,N_13608);
or U19494 (N_19494,N_13080,N_13644);
xnor U19495 (N_19495,N_14414,N_13941);
nand U19496 (N_19496,N_12374,N_12014);
xor U19497 (N_19497,N_14757,N_12735);
or U19498 (N_19498,N_12784,N_13583);
or U19499 (N_19499,N_14161,N_12108);
or U19500 (N_19500,N_12034,N_12498);
xor U19501 (N_19501,N_12364,N_13258);
nand U19502 (N_19502,N_14396,N_15551);
or U19503 (N_19503,N_14372,N_15914);
or U19504 (N_19504,N_15206,N_15637);
and U19505 (N_19505,N_12079,N_12068);
nand U19506 (N_19506,N_15848,N_14218);
and U19507 (N_19507,N_12380,N_14798);
nand U19508 (N_19508,N_14907,N_12077);
nor U19509 (N_19509,N_12097,N_13668);
xor U19510 (N_19510,N_15998,N_12001);
or U19511 (N_19511,N_12328,N_12079);
nand U19512 (N_19512,N_13713,N_12890);
xnor U19513 (N_19513,N_15276,N_14632);
or U19514 (N_19514,N_15800,N_13398);
nor U19515 (N_19515,N_15944,N_14735);
and U19516 (N_19516,N_13055,N_13224);
or U19517 (N_19517,N_14865,N_12818);
or U19518 (N_19518,N_12470,N_12480);
xor U19519 (N_19519,N_13451,N_13093);
nor U19520 (N_19520,N_14476,N_15262);
or U19521 (N_19521,N_15910,N_13644);
or U19522 (N_19522,N_15431,N_13418);
or U19523 (N_19523,N_12203,N_14967);
and U19524 (N_19524,N_12322,N_12415);
or U19525 (N_19525,N_13236,N_15616);
xor U19526 (N_19526,N_14147,N_15353);
nand U19527 (N_19527,N_14871,N_13403);
xnor U19528 (N_19528,N_14452,N_13212);
nor U19529 (N_19529,N_14303,N_13883);
xnor U19530 (N_19530,N_14279,N_14825);
nor U19531 (N_19531,N_12764,N_12614);
nand U19532 (N_19532,N_14017,N_13750);
nor U19533 (N_19533,N_12002,N_15788);
and U19534 (N_19534,N_13442,N_15398);
or U19535 (N_19535,N_13769,N_13355);
xnor U19536 (N_19536,N_12985,N_12568);
and U19537 (N_19537,N_12657,N_12806);
and U19538 (N_19538,N_12135,N_14181);
nor U19539 (N_19539,N_14273,N_14743);
nand U19540 (N_19540,N_15313,N_12385);
or U19541 (N_19541,N_12950,N_12445);
or U19542 (N_19542,N_12801,N_15995);
xor U19543 (N_19543,N_12588,N_13515);
xnor U19544 (N_19544,N_13251,N_13304);
xor U19545 (N_19545,N_13684,N_14398);
or U19546 (N_19546,N_13911,N_14963);
nor U19547 (N_19547,N_12549,N_14096);
and U19548 (N_19548,N_15073,N_14178);
or U19549 (N_19549,N_12310,N_12043);
or U19550 (N_19550,N_12390,N_15686);
xnor U19551 (N_19551,N_15073,N_15261);
and U19552 (N_19552,N_15186,N_15873);
xor U19553 (N_19553,N_15503,N_12436);
and U19554 (N_19554,N_14158,N_14243);
and U19555 (N_19555,N_12365,N_14105);
or U19556 (N_19556,N_15031,N_14991);
xnor U19557 (N_19557,N_15504,N_15570);
xnor U19558 (N_19558,N_15257,N_12371);
or U19559 (N_19559,N_13863,N_15639);
or U19560 (N_19560,N_14534,N_14673);
and U19561 (N_19561,N_15182,N_15043);
xnor U19562 (N_19562,N_12384,N_15109);
or U19563 (N_19563,N_13516,N_13571);
and U19564 (N_19564,N_13798,N_15549);
nand U19565 (N_19565,N_15986,N_13384);
or U19566 (N_19566,N_15807,N_12459);
or U19567 (N_19567,N_12077,N_13073);
nor U19568 (N_19568,N_15761,N_15948);
or U19569 (N_19569,N_15601,N_15527);
xor U19570 (N_19570,N_15073,N_15225);
nand U19571 (N_19571,N_12901,N_13599);
nor U19572 (N_19572,N_12948,N_14231);
xor U19573 (N_19573,N_14713,N_13958);
and U19574 (N_19574,N_14880,N_12127);
xor U19575 (N_19575,N_14001,N_13921);
nor U19576 (N_19576,N_12149,N_12311);
or U19577 (N_19577,N_13564,N_14933);
xnor U19578 (N_19578,N_12279,N_14960);
nor U19579 (N_19579,N_14724,N_14539);
nand U19580 (N_19580,N_14852,N_15242);
and U19581 (N_19581,N_13011,N_15488);
xor U19582 (N_19582,N_13730,N_13310);
or U19583 (N_19583,N_15294,N_14846);
and U19584 (N_19584,N_14539,N_14288);
nand U19585 (N_19585,N_12041,N_12803);
and U19586 (N_19586,N_13115,N_13706);
and U19587 (N_19587,N_15643,N_13136);
nor U19588 (N_19588,N_15034,N_13446);
xnor U19589 (N_19589,N_12240,N_12889);
xor U19590 (N_19590,N_15486,N_14888);
nor U19591 (N_19591,N_12853,N_14095);
xnor U19592 (N_19592,N_13604,N_15199);
nor U19593 (N_19593,N_14679,N_12029);
or U19594 (N_19594,N_14290,N_15750);
nor U19595 (N_19595,N_14858,N_14281);
xor U19596 (N_19596,N_14402,N_13821);
or U19597 (N_19597,N_15077,N_12939);
nor U19598 (N_19598,N_14082,N_13528);
nor U19599 (N_19599,N_14482,N_12299);
nand U19600 (N_19600,N_12002,N_15205);
and U19601 (N_19601,N_14260,N_15639);
nor U19602 (N_19602,N_14457,N_13720);
and U19603 (N_19603,N_13905,N_15422);
xor U19604 (N_19604,N_14998,N_14370);
nor U19605 (N_19605,N_15292,N_15425);
and U19606 (N_19606,N_12187,N_13227);
nor U19607 (N_19607,N_13751,N_14487);
xnor U19608 (N_19608,N_14126,N_13643);
nand U19609 (N_19609,N_14774,N_14356);
or U19610 (N_19610,N_15581,N_15486);
xnor U19611 (N_19611,N_14068,N_12744);
and U19612 (N_19612,N_13496,N_12998);
and U19613 (N_19613,N_14181,N_12861);
nor U19614 (N_19614,N_13824,N_15883);
and U19615 (N_19615,N_13843,N_13753);
xnor U19616 (N_19616,N_12876,N_15679);
nor U19617 (N_19617,N_14273,N_15369);
or U19618 (N_19618,N_13458,N_13914);
xnor U19619 (N_19619,N_12104,N_13832);
nor U19620 (N_19620,N_12412,N_12422);
and U19621 (N_19621,N_15428,N_13003);
nor U19622 (N_19622,N_15754,N_14676);
nor U19623 (N_19623,N_14152,N_13421);
nand U19624 (N_19624,N_12969,N_14177);
or U19625 (N_19625,N_12278,N_15359);
and U19626 (N_19626,N_12285,N_15128);
nor U19627 (N_19627,N_12440,N_12473);
nand U19628 (N_19628,N_12546,N_14542);
nor U19629 (N_19629,N_15175,N_13326);
xor U19630 (N_19630,N_13131,N_12776);
xnor U19631 (N_19631,N_15097,N_13371);
or U19632 (N_19632,N_12420,N_13362);
xor U19633 (N_19633,N_15601,N_14175);
nor U19634 (N_19634,N_15153,N_12394);
and U19635 (N_19635,N_13235,N_13089);
nor U19636 (N_19636,N_14439,N_13352);
and U19637 (N_19637,N_14514,N_13676);
nand U19638 (N_19638,N_13080,N_15894);
nand U19639 (N_19639,N_12208,N_12889);
and U19640 (N_19640,N_14024,N_15833);
xnor U19641 (N_19641,N_15570,N_12702);
xnor U19642 (N_19642,N_15458,N_14023);
nor U19643 (N_19643,N_13857,N_14558);
nor U19644 (N_19644,N_13564,N_13437);
xor U19645 (N_19645,N_15934,N_13476);
xnor U19646 (N_19646,N_15159,N_14028);
or U19647 (N_19647,N_13915,N_15106);
xor U19648 (N_19648,N_12333,N_14972);
or U19649 (N_19649,N_13022,N_14620);
nand U19650 (N_19650,N_15935,N_14192);
or U19651 (N_19651,N_15909,N_13254);
nor U19652 (N_19652,N_12301,N_14265);
xnor U19653 (N_19653,N_15144,N_15665);
xnor U19654 (N_19654,N_12112,N_14852);
or U19655 (N_19655,N_14160,N_13913);
nand U19656 (N_19656,N_15865,N_12112);
nand U19657 (N_19657,N_12200,N_13456);
or U19658 (N_19658,N_14427,N_12701);
nand U19659 (N_19659,N_14818,N_13947);
nor U19660 (N_19660,N_15698,N_13586);
and U19661 (N_19661,N_14429,N_12594);
nor U19662 (N_19662,N_15454,N_12112);
xor U19663 (N_19663,N_15179,N_13709);
and U19664 (N_19664,N_14671,N_13735);
or U19665 (N_19665,N_12542,N_12487);
xnor U19666 (N_19666,N_12396,N_13555);
nand U19667 (N_19667,N_13930,N_13128);
nand U19668 (N_19668,N_13633,N_12577);
or U19669 (N_19669,N_14709,N_13353);
or U19670 (N_19670,N_12832,N_14783);
and U19671 (N_19671,N_12137,N_14816);
and U19672 (N_19672,N_15465,N_15856);
or U19673 (N_19673,N_12512,N_13331);
nor U19674 (N_19674,N_12290,N_15408);
or U19675 (N_19675,N_13188,N_13847);
or U19676 (N_19676,N_15033,N_12788);
or U19677 (N_19677,N_14388,N_13166);
nand U19678 (N_19678,N_13578,N_12699);
and U19679 (N_19679,N_12037,N_13617);
and U19680 (N_19680,N_13189,N_14437);
or U19681 (N_19681,N_13233,N_15526);
nand U19682 (N_19682,N_15087,N_14253);
xnor U19683 (N_19683,N_12886,N_12863);
xor U19684 (N_19684,N_12743,N_14628);
or U19685 (N_19685,N_13914,N_14323);
or U19686 (N_19686,N_14502,N_13777);
or U19687 (N_19687,N_14641,N_13147);
xor U19688 (N_19688,N_13011,N_14197);
nor U19689 (N_19689,N_12549,N_12836);
or U19690 (N_19690,N_14771,N_13257);
or U19691 (N_19691,N_12101,N_12907);
nand U19692 (N_19692,N_15065,N_15638);
and U19693 (N_19693,N_13345,N_12668);
or U19694 (N_19694,N_12108,N_15439);
xor U19695 (N_19695,N_15456,N_12152);
nor U19696 (N_19696,N_14577,N_13446);
or U19697 (N_19697,N_12517,N_15195);
xor U19698 (N_19698,N_15852,N_14865);
xor U19699 (N_19699,N_12724,N_14911);
and U19700 (N_19700,N_14301,N_12820);
nand U19701 (N_19701,N_14728,N_14784);
nand U19702 (N_19702,N_15445,N_12305);
or U19703 (N_19703,N_14982,N_13186);
or U19704 (N_19704,N_14151,N_12134);
xnor U19705 (N_19705,N_14223,N_12674);
and U19706 (N_19706,N_15356,N_15446);
or U19707 (N_19707,N_12668,N_13642);
and U19708 (N_19708,N_13419,N_15495);
nor U19709 (N_19709,N_14525,N_15599);
nor U19710 (N_19710,N_14486,N_15054);
and U19711 (N_19711,N_13586,N_15268);
nand U19712 (N_19712,N_13411,N_12825);
xnor U19713 (N_19713,N_14053,N_12664);
xnor U19714 (N_19714,N_13329,N_12287);
nand U19715 (N_19715,N_14775,N_13196);
nor U19716 (N_19716,N_13382,N_13610);
xnor U19717 (N_19717,N_12457,N_14189);
xor U19718 (N_19718,N_12339,N_13829);
and U19719 (N_19719,N_14420,N_12892);
xnor U19720 (N_19720,N_14618,N_15081);
or U19721 (N_19721,N_15038,N_14963);
or U19722 (N_19722,N_14209,N_12226);
nor U19723 (N_19723,N_14985,N_12782);
or U19724 (N_19724,N_13459,N_13869);
nand U19725 (N_19725,N_14353,N_15070);
nand U19726 (N_19726,N_14666,N_12628);
nor U19727 (N_19727,N_13579,N_13317);
nand U19728 (N_19728,N_13176,N_14559);
and U19729 (N_19729,N_14100,N_14208);
nor U19730 (N_19730,N_12621,N_13183);
xnor U19731 (N_19731,N_15042,N_14412);
nor U19732 (N_19732,N_13081,N_13949);
or U19733 (N_19733,N_12376,N_13437);
nand U19734 (N_19734,N_13320,N_13090);
or U19735 (N_19735,N_14328,N_13519);
and U19736 (N_19736,N_15416,N_13887);
nor U19737 (N_19737,N_12907,N_12540);
nand U19738 (N_19738,N_15435,N_12094);
or U19739 (N_19739,N_12108,N_14225);
xnor U19740 (N_19740,N_14221,N_12160);
nor U19741 (N_19741,N_13365,N_14232);
nand U19742 (N_19742,N_13532,N_15985);
nand U19743 (N_19743,N_13058,N_15913);
xnor U19744 (N_19744,N_13774,N_12394);
nor U19745 (N_19745,N_15004,N_14680);
nand U19746 (N_19746,N_14093,N_12279);
nand U19747 (N_19747,N_14904,N_14127);
nor U19748 (N_19748,N_13751,N_13797);
or U19749 (N_19749,N_14444,N_12181);
and U19750 (N_19750,N_13388,N_13309);
nor U19751 (N_19751,N_12264,N_15004);
or U19752 (N_19752,N_15055,N_14722);
or U19753 (N_19753,N_14948,N_15733);
xor U19754 (N_19754,N_15601,N_12140);
and U19755 (N_19755,N_15483,N_14969);
or U19756 (N_19756,N_14065,N_13589);
nor U19757 (N_19757,N_14785,N_14339);
nand U19758 (N_19758,N_12723,N_15940);
or U19759 (N_19759,N_13041,N_14893);
or U19760 (N_19760,N_13536,N_14946);
xor U19761 (N_19761,N_13591,N_13628);
nor U19762 (N_19762,N_15033,N_13857);
xnor U19763 (N_19763,N_15611,N_13747);
or U19764 (N_19764,N_12463,N_15176);
or U19765 (N_19765,N_14303,N_14988);
nand U19766 (N_19766,N_15477,N_12076);
and U19767 (N_19767,N_13181,N_15975);
nor U19768 (N_19768,N_14514,N_13851);
and U19769 (N_19769,N_13049,N_12936);
or U19770 (N_19770,N_13973,N_13093);
or U19771 (N_19771,N_14447,N_12781);
xor U19772 (N_19772,N_15580,N_13164);
nor U19773 (N_19773,N_13339,N_12782);
nor U19774 (N_19774,N_12525,N_14901);
xnor U19775 (N_19775,N_14757,N_15920);
and U19776 (N_19776,N_14526,N_15383);
nor U19777 (N_19777,N_13108,N_13976);
nor U19778 (N_19778,N_15453,N_15589);
xnor U19779 (N_19779,N_13781,N_14419);
nand U19780 (N_19780,N_14359,N_14136);
nor U19781 (N_19781,N_13633,N_13802);
nand U19782 (N_19782,N_14979,N_15706);
nand U19783 (N_19783,N_14931,N_12272);
or U19784 (N_19784,N_13757,N_13091);
nand U19785 (N_19785,N_15441,N_14223);
and U19786 (N_19786,N_12200,N_14988);
and U19787 (N_19787,N_15004,N_13144);
or U19788 (N_19788,N_12435,N_14530);
nand U19789 (N_19789,N_13792,N_13027);
nor U19790 (N_19790,N_15781,N_15104);
and U19791 (N_19791,N_13468,N_14041);
nor U19792 (N_19792,N_13315,N_14285);
nand U19793 (N_19793,N_12766,N_15426);
xnor U19794 (N_19794,N_14661,N_12844);
or U19795 (N_19795,N_15891,N_12103);
and U19796 (N_19796,N_15714,N_15253);
nor U19797 (N_19797,N_14735,N_15888);
and U19798 (N_19798,N_14979,N_13336);
nand U19799 (N_19799,N_12601,N_14698);
nand U19800 (N_19800,N_13438,N_15168);
and U19801 (N_19801,N_12982,N_14249);
xnor U19802 (N_19802,N_12971,N_15109);
xnor U19803 (N_19803,N_15198,N_15561);
or U19804 (N_19804,N_14658,N_14492);
or U19805 (N_19805,N_14591,N_12146);
or U19806 (N_19806,N_15662,N_13891);
xor U19807 (N_19807,N_14198,N_12267);
xnor U19808 (N_19808,N_14268,N_14195);
xor U19809 (N_19809,N_13736,N_15241);
xor U19810 (N_19810,N_13366,N_12904);
xnor U19811 (N_19811,N_12107,N_14375);
or U19812 (N_19812,N_13871,N_14580);
xor U19813 (N_19813,N_13537,N_13045);
and U19814 (N_19814,N_13963,N_12725);
nor U19815 (N_19815,N_14938,N_12754);
and U19816 (N_19816,N_13941,N_15081);
or U19817 (N_19817,N_14777,N_13762);
xor U19818 (N_19818,N_15351,N_14767);
nor U19819 (N_19819,N_12207,N_15388);
xor U19820 (N_19820,N_15893,N_12418);
nand U19821 (N_19821,N_13990,N_13548);
and U19822 (N_19822,N_15516,N_15495);
xor U19823 (N_19823,N_12828,N_15277);
xnor U19824 (N_19824,N_12361,N_12111);
nor U19825 (N_19825,N_15803,N_13360);
nor U19826 (N_19826,N_13759,N_13024);
and U19827 (N_19827,N_15928,N_15604);
or U19828 (N_19828,N_13477,N_14827);
and U19829 (N_19829,N_12523,N_15177);
nand U19830 (N_19830,N_15530,N_12612);
xor U19831 (N_19831,N_14690,N_12552);
nor U19832 (N_19832,N_14629,N_14051);
or U19833 (N_19833,N_12154,N_14233);
nand U19834 (N_19834,N_13158,N_14652);
nor U19835 (N_19835,N_15018,N_14416);
xor U19836 (N_19836,N_12045,N_13548);
or U19837 (N_19837,N_12797,N_15973);
xor U19838 (N_19838,N_12277,N_15537);
xnor U19839 (N_19839,N_13156,N_14300);
nand U19840 (N_19840,N_13297,N_14364);
and U19841 (N_19841,N_13578,N_15662);
or U19842 (N_19842,N_15615,N_14218);
nand U19843 (N_19843,N_13874,N_13669);
nor U19844 (N_19844,N_15906,N_15018);
and U19845 (N_19845,N_15181,N_15145);
nand U19846 (N_19846,N_13888,N_14788);
and U19847 (N_19847,N_12348,N_13492);
xnor U19848 (N_19848,N_12341,N_12778);
nor U19849 (N_19849,N_14357,N_15378);
nand U19850 (N_19850,N_15783,N_12196);
nand U19851 (N_19851,N_15868,N_15078);
xnor U19852 (N_19852,N_12580,N_15489);
nand U19853 (N_19853,N_12528,N_14246);
nor U19854 (N_19854,N_12973,N_13554);
xor U19855 (N_19855,N_13455,N_15918);
xor U19856 (N_19856,N_13904,N_15300);
nor U19857 (N_19857,N_13640,N_15467);
nor U19858 (N_19858,N_12143,N_12908);
nor U19859 (N_19859,N_15054,N_14981);
and U19860 (N_19860,N_14110,N_14620);
nor U19861 (N_19861,N_14910,N_13567);
nand U19862 (N_19862,N_14484,N_15956);
nor U19863 (N_19863,N_14584,N_15844);
xnor U19864 (N_19864,N_15102,N_14775);
nor U19865 (N_19865,N_15862,N_15733);
xnor U19866 (N_19866,N_13952,N_14219);
or U19867 (N_19867,N_15877,N_13053);
or U19868 (N_19868,N_15640,N_14467);
nor U19869 (N_19869,N_13275,N_15697);
nand U19870 (N_19870,N_13514,N_13450);
xor U19871 (N_19871,N_14674,N_13662);
and U19872 (N_19872,N_15698,N_13473);
nand U19873 (N_19873,N_13766,N_12083);
xnor U19874 (N_19874,N_14515,N_12499);
nand U19875 (N_19875,N_15127,N_12138);
or U19876 (N_19876,N_13386,N_12345);
xor U19877 (N_19877,N_14747,N_13777);
xor U19878 (N_19878,N_12768,N_14188);
and U19879 (N_19879,N_14045,N_14708);
and U19880 (N_19880,N_14838,N_14777);
and U19881 (N_19881,N_12793,N_14585);
or U19882 (N_19882,N_12900,N_15389);
and U19883 (N_19883,N_14936,N_12098);
nand U19884 (N_19884,N_15225,N_12327);
and U19885 (N_19885,N_14091,N_14912);
xnor U19886 (N_19886,N_12694,N_12071);
and U19887 (N_19887,N_15524,N_15586);
or U19888 (N_19888,N_13043,N_15115);
nor U19889 (N_19889,N_12055,N_15980);
nand U19890 (N_19890,N_13019,N_15575);
nand U19891 (N_19891,N_15147,N_14429);
or U19892 (N_19892,N_12485,N_15813);
or U19893 (N_19893,N_12927,N_12970);
or U19894 (N_19894,N_14966,N_15187);
nand U19895 (N_19895,N_14883,N_13952);
or U19896 (N_19896,N_13642,N_15770);
and U19897 (N_19897,N_14882,N_13054);
nor U19898 (N_19898,N_14132,N_15774);
nor U19899 (N_19899,N_12944,N_15325);
and U19900 (N_19900,N_13314,N_13866);
xor U19901 (N_19901,N_13417,N_14466);
and U19902 (N_19902,N_13814,N_15865);
and U19903 (N_19903,N_13700,N_14650);
nor U19904 (N_19904,N_14860,N_14886);
nand U19905 (N_19905,N_13222,N_14295);
xnor U19906 (N_19906,N_12540,N_15125);
nand U19907 (N_19907,N_14245,N_13952);
or U19908 (N_19908,N_15225,N_12348);
nand U19909 (N_19909,N_15521,N_12590);
nor U19910 (N_19910,N_12673,N_12715);
and U19911 (N_19911,N_12489,N_15564);
nor U19912 (N_19912,N_12639,N_13651);
nor U19913 (N_19913,N_13376,N_15874);
xnor U19914 (N_19914,N_13095,N_15495);
nor U19915 (N_19915,N_12175,N_12701);
nor U19916 (N_19916,N_15672,N_14494);
nor U19917 (N_19917,N_13400,N_12970);
nand U19918 (N_19918,N_15970,N_15153);
or U19919 (N_19919,N_14736,N_14067);
xnor U19920 (N_19920,N_14287,N_14728);
or U19921 (N_19921,N_15821,N_14751);
and U19922 (N_19922,N_15033,N_13535);
or U19923 (N_19923,N_14734,N_13121);
nand U19924 (N_19924,N_12836,N_12420);
xor U19925 (N_19925,N_14832,N_13482);
nand U19926 (N_19926,N_13387,N_13449);
and U19927 (N_19927,N_12557,N_15995);
and U19928 (N_19928,N_12655,N_15372);
and U19929 (N_19929,N_12541,N_15840);
nand U19930 (N_19930,N_15803,N_14426);
and U19931 (N_19931,N_13861,N_14696);
or U19932 (N_19932,N_15090,N_13412);
or U19933 (N_19933,N_15093,N_13588);
and U19934 (N_19934,N_15623,N_15038);
nor U19935 (N_19935,N_14513,N_15320);
and U19936 (N_19936,N_13109,N_15220);
or U19937 (N_19937,N_13264,N_14099);
nand U19938 (N_19938,N_12258,N_12440);
and U19939 (N_19939,N_12335,N_14571);
nor U19940 (N_19940,N_13766,N_15610);
nand U19941 (N_19941,N_13924,N_14567);
xor U19942 (N_19942,N_12626,N_12279);
and U19943 (N_19943,N_13107,N_12885);
or U19944 (N_19944,N_12101,N_12747);
and U19945 (N_19945,N_15645,N_14175);
xnor U19946 (N_19946,N_13084,N_14075);
nand U19947 (N_19947,N_13849,N_14321);
nor U19948 (N_19948,N_15602,N_15648);
xnor U19949 (N_19949,N_14460,N_13584);
nor U19950 (N_19950,N_14117,N_14437);
nor U19951 (N_19951,N_12462,N_12834);
nor U19952 (N_19952,N_12812,N_12757);
xor U19953 (N_19953,N_14820,N_13549);
nor U19954 (N_19954,N_14044,N_15364);
xor U19955 (N_19955,N_13258,N_14778);
and U19956 (N_19956,N_15783,N_14424);
or U19957 (N_19957,N_15265,N_13577);
xnor U19958 (N_19958,N_13693,N_14998);
xnor U19959 (N_19959,N_13481,N_12559);
and U19960 (N_19960,N_14559,N_14149);
nand U19961 (N_19961,N_15243,N_13974);
or U19962 (N_19962,N_12193,N_14513);
or U19963 (N_19963,N_15209,N_15551);
and U19964 (N_19964,N_13896,N_12010);
nand U19965 (N_19965,N_13998,N_15126);
or U19966 (N_19966,N_14463,N_15563);
or U19967 (N_19967,N_12838,N_12988);
xnor U19968 (N_19968,N_15693,N_14556);
and U19969 (N_19969,N_12902,N_15086);
or U19970 (N_19970,N_14905,N_13825);
nor U19971 (N_19971,N_14653,N_12404);
or U19972 (N_19972,N_15628,N_15262);
xnor U19973 (N_19973,N_14618,N_13927);
xnor U19974 (N_19974,N_13426,N_15567);
nor U19975 (N_19975,N_12097,N_15252);
and U19976 (N_19976,N_13564,N_12967);
xor U19977 (N_19977,N_14979,N_12117);
xor U19978 (N_19978,N_15588,N_14868);
nand U19979 (N_19979,N_15237,N_12625);
or U19980 (N_19980,N_15934,N_15132);
or U19981 (N_19981,N_14243,N_12321);
or U19982 (N_19982,N_12680,N_14826);
or U19983 (N_19983,N_12378,N_15504);
and U19984 (N_19984,N_12158,N_14707);
or U19985 (N_19985,N_13058,N_13572);
nor U19986 (N_19986,N_14699,N_13017);
or U19987 (N_19987,N_15324,N_14802);
xnor U19988 (N_19988,N_15622,N_12106);
and U19989 (N_19989,N_14524,N_13987);
xor U19990 (N_19990,N_13632,N_13882);
xnor U19991 (N_19991,N_14564,N_14740);
and U19992 (N_19992,N_13964,N_15523);
or U19993 (N_19993,N_14542,N_12627);
nor U19994 (N_19994,N_15502,N_15610);
or U19995 (N_19995,N_13652,N_15010);
xor U19996 (N_19996,N_15964,N_15493);
or U19997 (N_19997,N_14476,N_15548);
nor U19998 (N_19998,N_14049,N_15401);
xor U19999 (N_19999,N_14811,N_14496);
nor UO_0 (O_0,N_17240,N_18528);
xor UO_1 (O_1,N_17335,N_17539);
and UO_2 (O_2,N_16490,N_18133);
and UO_3 (O_3,N_17914,N_16540);
xnor UO_4 (O_4,N_17724,N_17264);
nor UO_5 (O_5,N_18939,N_19662);
nor UO_6 (O_6,N_16979,N_18204);
nand UO_7 (O_7,N_17963,N_16534);
and UO_8 (O_8,N_18048,N_16643);
nand UO_9 (O_9,N_19119,N_19982);
nor UO_10 (O_10,N_17956,N_17518);
nor UO_11 (O_11,N_19410,N_19405);
or UO_12 (O_12,N_18598,N_16424);
nor UO_13 (O_13,N_18056,N_17633);
and UO_14 (O_14,N_19913,N_16998);
and UO_15 (O_15,N_18146,N_19866);
nand UO_16 (O_16,N_18454,N_16138);
nor UO_17 (O_17,N_17226,N_17986);
xor UO_18 (O_18,N_19779,N_18444);
and UO_19 (O_19,N_16429,N_16835);
nor UO_20 (O_20,N_19892,N_19879);
nor UO_21 (O_21,N_16282,N_19669);
nand UO_22 (O_22,N_16633,N_19602);
and UO_23 (O_23,N_17588,N_19003);
xor UO_24 (O_24,N_19332,N_18777);
nor UO_25 (O_25,N_16740,N_18693);
nand UO_26 (O_26,N_19382,N_19352);
xnor UO_27 (O_27,N_18807,N_19624);
nand UO_28 (O_28,N_18360,N_17464);
xor UO_29 (O_29,N_16386,N_18695);
nor UO_30 (O_30,N_17296,N_18317);
nor UO_31 (O_31,N_17402,N_16045);
xor UO_32 (O_32,N_18069,N_18718);
nand UO_33 (O_33,N_19653,N_17259);
nand UO_34 (O_34,N_16018,N_19776);
nor UO_35 (O_35,N_19823,N_17883);
xor UO_36 (O_36,N_17526,N_19907);
nor UO_37 (O_37,N_17272,N_17218);
xor UO_38 (O_38,N_18944,N_17051);
nor UO_39 (O_39,N_19145,N_16013);
nand UO_40 (O_40,N_18858,N_16396);
xnor UO_41 (O_41,N_16972,N_18117);
and UO_42 (O_42,N_18565,N_18438);
and UO_43 (O_43,N_16954,N_19717);
nor UO_44 (O_44,N_16789,N_18713);
xor UO_45 (O_45,N_18123,N_17144);
xnor UO_46 (O_46,N_19308,N_17171);
nand UO_47 (O_47,N_17784,N_18768);
nand UO_48 (O_48,N_17931,N_18918);
nand UO_49 (O_49,N_17911,N_16044);
and UO_50 (O_50,N_16901,N_19791);
xnor UO_51 (O_51,N_19001,N_19836);
or UO_52 (O_52,N_17720,N_16423);
nand UO_53 (O_53,N_17418,N_19680);
nor UO_54 (O_54,N_18689,N_18924);
nor UO_55 (O_55,N_18983,N_17180);
or UO_56 (O_56,N_17184,N_16022);
or UO_57 (O_57,N_19048,N_19707);
nor UO_58 (O_58,N_18011,N_17777);
and UO_59 (O_59,N_17554,N_16582);
nand UO_60 (O_60,N_18063,N_17389);
nand UO_61 (O_61,N_18461,N_16058);
nand UO_62 (O_62,N_19792,N_18813);
nand UO_63 (O_63,N_17160,N_18422);
nand UO_64 (O_64,N_16447,N_19325);
or UO_65 (O_65,N_18266,N_18946);
nand UO_66 (O_66,N_18212,N_19129);
nor UO_67 (O_67,N_19128,N_17620);
xnor UO_68 (O_68,N_17982,N_16186);
nand UO_69 (O_69,N_18760,N_18530);
or UO_70 (O_70,N_17084,N_17006);
nor UO_71 (O_71,N_16555,N_19206);
nor UO_72 (O_72,N_16224,N_16362);
and UO_73 (O_73,N_16001,N_19856);
xnor UO_74 (O_74,N_18774,N_18242);
xnor UO_75 (O_75,N_18451,N_16295);
and UO_76 (O_76,N_17353,N_16933);
xor UO_77 (O_77,N_16188,N_18080);
nor UO_78 (O_78,N_19234,N_18670);
xnor UO_79 (O_79,N_17043,N_18015);
or UO_80 (O_80,N_19545,N_17081);
xnor UO_81 (O_81,N_18331,N_19241);
xnor UO_82 (O_82,N_17415,N_18111);
nand UO_83 (O_83,N_18648,N_18621);
or UO_84 (O_84,N_18855,N_17717);
or UO_85 (O_85,N_17749,N_19228);
or UO_86 (O_86,N_17099,N_19588);
xor UO_87 (O_87,N_17787,N_18909);
xor UO_88 (O_88,N_16808,N_19712);
and UO_89 (O_89,N_16019,N_18580);
or UO_90 (O_90,N_19273,N_16779);
xor UO_91 (O_91,N_17541,N_17205);
nor UO_92 (O_92,N_16595,N_17332);
and UO_93 (O_93,N_19829,N_18634);
or UO_94 (O_94,N_17623,N_17384);
and UO_95 (O_95,N_17577,N_19028);
nand UO_96 (O_96,N_17169,N_17894);
and UO_97 (O_97,N_17879,N_17374);
xor UO_98 (O_98,N_18669,N_16104);
nand UO_99 (O_99,N_18059,N_19231);
or UO_100 (O_100,N_18746,N_18811);
nand UO_101 (O_101,N_17032,N_16590);
nor UO_102 (O_102,N_19905,N_18841);
or UO_103 (O_103,N_19630,N_16002);
or UO_104 (O_104,N_19572,N_16800);
xor UO_105 (O_105,N_17165,N_17131);
and UO_106 (O_106,N_18042,N_16694);
nand UO_107 (O_107,N_19169,N_16689);
and UO_108 (O_108,N_19350,N_19246);
nor UO_109 (O_109,N_16365,N_18865);
xor UO_110 (O_110,N_17738,N_17729);
nor UO_111 (O_111,N_19432,N_18299);
or UO_112 (O_112,N_17714,N_19867);
nor UO_113 (O_113,N_17731,N_18156);
and UO_114 (O_114,N_16241,N_19938);
nand UO_115 (O_115,N_18455,N_19392);
xor UO_116 (O_116,N_17115,N_17311);
nor UO_117 (O_117,N_16531,N_19356);
nor UO_118 (O_118,N_19488,N_19577);
nor UO_119 (O_119,N_19262,N_18894);
nor UO_120 (O_120,N_18880,N_19207);
xnor UO_121 (O_121,N_17613,N_16654);
nor UO_122 (O_122,N_16341,N_16592);
nor UO_123 (O_123,N_18188,N_18263);
or UO_124 (O_124,N_17549,N_19966);
nand UO_125 (O_125,N_17647,N_18002);
nor UO_126 (O_126,N_19529,N_19973);
and UO_127 (O_127,N_19265,N_16803);
nor UO_128 (O_128,N_19211,N_16255);
nand UO_129 (O_129,N_17905,N_17453);
xnor UO_130 (O_130,N_19366,N_18546);
or UO_131 (O_131,N_17095,N_19322);
nor UO_132 (O_132,N_16619,N_16561);
nor UO_133 (O_133,N_18883,N_17182);
xnor UO_134 (O_134,N_16693,N_19161);
nand UO_135 (O_135,N_16776,N_17460);
nand UO_136 (O_136,N_17536,N_19224);
nor UO_137 (O_137,N_17607,N_18071);
and UO_138 (O_138,N_19491,N_17591);
and UO_139 (O_139,N_19301,N_18707);
or UO_140 (O_140,N_16005,N_16785);
or UO_141 (O_141,N_18549,N_16956);
or UO_142 (O_142,N_17364,N_19705);
nand UO_143 (O_143,N_19138,N_18493);
and UO_144 (O_144,N_16538,N_19203);
xnor UO_145 (O_145,N_18917,N_18976);
and UO_146 (O_146,N_18828,N_16210);
nor UO_147 (O_147,N_18110,N_19004);
nor UO_148 (O_148,N_18936,N_19385);
nand UO_149 (O_149,N_19146,N_16218);
xor UO_150 (O_150,N_17912,N_18605);
nor UO_151 (O_151,N_16705,N_16037);
xor UO_152 (O_152,N_16411,N_18325);
xnor UO_153 (O_153,N_18866,N_16317);
and UO_154 (O_154,N_19337,N_16075);
nor UO_155 (O_155,N_17725,N_17370);
nand UO_156 (O_156,N_17423,N_19578);
xor UO_157 (O_157,N_19828,N_19798);
nor UO_158 (O_158,N_17028,N_18700);
xor UO_159 (O_159,N_18393,N_19525);
or UO_160 (O_160,N_19674,N_19271);
nand UO_161 (O_161,N_19100,N_19341);
or UO_162 (O_162,N_19476,N_19888);
and UO_163 (O_163,N_19229,N_18950);
nor UO_164 (O_164,N_17576,N_19903);
xnor UO_165 (O_165,N_18642,N_17452);
nand UO_166 (O_166,N_16986,N_18414);
nand UO_167 (O_167,N_17501,N_19898);
nand UO_168 (O_168,N_17571,N_17929);
nor UO_169 (O_169,N_19771,N_18968);
xor UO_170 (O_170,N_19761,N_19181);
nand UO_171 (O_171,N_19453,N_19740);
nor UO_172 (O_172,N_16105,N_18376);
nor UO_173 (O_173,N_16134,N_17872);
or UO_174 (O_174,N_16818,N_16527);
xor UO_175 (O_175,N_18398,N_18551);
and UO_176 (O_176,N_19825,N_16680);
nand UO_177 (O_177,N_19643,N_19818);
xnor UO_178 (O_178,N_18726,N_18388);
and UO_179 (O_179,N_18929,N_17835);
xor UO_180 (O_180,N_19451,N_16865);
nor UO_181 (O_181,N_16358,N_17818);
xnor UO_182 (O_182,N_19162,N_18137);
and UO_183 (O_183,N_19500,N_16128);
xnor UO_184 (O_184,N_17420,N_19587);
and UO_185 (O_185,N_16982,N_18629);
nor UO_186 (O_186,N_18336,N_19394);
or UO_187 (O_187,N_19296,N_18674);
nor UO_188 (O_188,N_16565,N_17670);
xor UO_189 (O_189,N_16398,N_16057);
nor UO_190 (O_190,N_19507,N_19749);
nand UO_191 (O_191,N_19232,N_19972);
nor UO_192 (O_192,N_16922,N_16859);
nor UO_193 (O_193,N_16618,N_17637);
nand UO_194 (O_194,N_19302,N_17298);
nor UO_195 (O_195,N_19091,N_18692);
nor UO_196 (O_196,N_19046,N_19713);
xor UO_197 (O_197,N_16043,N_16091);
nor UO_198 (O_198,N_17207,N_18226);
nor UO_199 (O_199,N_18282,N_17992);
xnor UO_200 (O_200,N_19196,N_19735);
and UO_201 (O_201,N_18889,N_19163);
nor UO_202 (O_202,N_18129,N_16383);
xor UO_203 (O_203,N_18098,N_19878);
xnor UO_204 (O_204,N_19359,N_16127);
xnor UO_205 (O_205,N_16431,N_19011);
nand UO_206 (O_206,N_16201,N_18119);
or UO_207 (O_207,N_18443,N_18966);
xor UO_208 (O_208,N_19752,N_18736);
xor UO_209 (O_209,N_18538,N_19005);
nand UO_210 (O_210,N_18987,N_18440);
and UO_211 (O_211,N_19992,N_19147);
and UO_212 (O_212,N_19266,N_17122);
and UO_213 (O_213,N_19851,N_17831);
xor UO_214 (O_214,N_16941,N_17202);
nand UO_215 (O_215,N_18036,N_18646);
xor UO_216 (O_216,N_19695,N_19551);
and UO_217 (O_217,N_18896,N_19516);
and UO_218 (O_218,N_17926,N_16962);
nand UO_219 (O_219,N_16376,N_16292);
or UO_220 (O_220,N_16512,N_17054);
xnor UO_221 (O_221,N_18751,N_18039);
nand UO_222 (O_222,N_18506,N_18554);
nor UO_223 (O_223,N_18402,N_19092);
xor UO_224 (O_224,N_17543,N_18279);
nand UO_225 (O_225,N_16525,N_19137);
or UO_226 (O_226,N_17373,N_19700);
or UO_227 (O_227,N_17474,N_19801);
nor UO_228 (O_228,N_19351,N_18053);
and UO_229 (O_229,N_16288,N_17398);
nand UO_230 (O_230,N_17593,N_17712);
and UO_231 (O_231,N_17563,N_19861);
xor UO_232 (O_232,N_18335,N_18609);
or UO_233 (O_233,N_17651,N_18151);
nand UO_234 (O_234,N_17938,N_16416);
xor UO_235 (O_235,N_16316,N_19974);
nor UO_236 (O_236,N_16794,N_18179);
xor UO_237 (O_237,N_17959,N_18711);
and UO_238 (O_238,N_18259,N_18287);
and UO_239 (O_239,N_17442,N_17354);
nor UO_240 (O_240,N_19919,N_18734);
and UO_241 (O_241,N_19843,N_16486);
xnor UO_242 (O_242,N_19074,N_16250);
and UO_243 (O_243,N_19789,N_16484);
xnor UO_244 (O_244,N_18367,N_18787);
and UO_245 (O_245,N_19720,N_16896);
nor UO_246 (O_246,N_18792,N_16636);
or UO_247 (O_247,N_18116,N_19734);
or UO_248 (O_248,N_18931,N_17570);
or UO_249 (O_249,N_18547,N_17198);
or UO_250 (O_250,N_18427,N_18076);
and UO_251 (O_251,N_17290,N_16456);
and UO_252 (O_252,N_18521,N_17251);
and UO_253 (O_253,N_16517,N_18384);
and UO_254 (O_254,N_19256,N_16994);
xor UO_255 (O_255,N_17341,N_16702);
nor UO_256 (O_256,N_18884,N_17275);
xnor UO_257 (O_257,N_18213,N_19540);
or UO_258 (O_258,N_19418,N_17928);
or UO_259 (O_259,N_16603,N_18871);
or UO_260 (O_260,N_17621,N_17252);
xor UO_261 (O_261,N_18344,N_19809);
or UO_262 (O_262,N_19200,N_16237);
or UO_263 (O_263,N_18560,N_19514);
nand UO_264 (O_264,N_18687,N_19444);
or UO_265 (O_265,N_16844,N_18870);
and UO_266 (O_266,N_16627,N_16821);
xor UO_267 (O_267,N_19549,N_18254);
and UO_268 (O_268,N_17480,N_17089);
or UO_269 (O_269,N_17346,N_17137);
nand UO_270 (O_270,N_17261,N_17628);
and UO_271 (O_271,N_17987,N_19284);
and UO_272 (O_272,N_18714,N_16165);
nor UO_273 (O_273,N_17219,N_18963);
and UO_274 (O_274,N_16784,N_17098);
xnor UO_275 (O_275,N_16169,N_18154);
and UO_276 (O_276,N_17827,N_17408);
xor UO_277 (O_277,N_16069,N_18186);
nor UO_278 (O_278,N_17005,N_17826);
nand UO_279 (O_279,N_18847,N_19413);
nor UO_280 (O_280,N_17737,N_19852);
or UO_281 (O_281,N_16573,N_18780);
and UO_282 (O_282,N_18334,N_19032);
xnor UO_283 (O_283,N_16378,N_16185);
xnor UO_284 (O_284,N_19821,N_16810);
nand UO_285 (O_285,N_16052,N_18663);
xor UO_286 (O_286,N_18104,N_18737);
and UO_287 (O_287,N_18868,N_16966);
or UO_288 (O_288,N_17136,N_16737);
nor UO_289 (O_289,N_19227,N_17813);
and UO_290 (O_290,N_16629,N_19885);
nor UO_291 (O_291,N_18550,N_16747);
xor UO_292 (O_292,N_18201,N_17154);
nor UO_293 (O_293,N_16602,N_17096);
and UO_294 (O_294,N_19567,N_19117);
xor UO_295 (O_295,N_16313,N_18057);
or UO_296 (O_296,N_19044,N_18582);
nor UO_297 (O_297,N_17328,N_18743);
nand UO_298 (O_298,N_16920,N_19558);
or UO_299 (O_299,N_16154,N_17809);
or UO_300 (O_300,N_19564,N_16221);
xnor UO_301 (O_301,N_16940,N_19378);
nand UO_302 (O_302,N_16196,N_18407);
and UO_303 (O_303,N_17432,N_17677);
xor UO_304 (O_304,N_19718,N_16068);
nand UO_305 (O_305,N_17605,N_19927);
nand UO_306 (O_306,N_18463,N_19306);
or UO_307 (O_307,N_19945,N_18522);
and UO_308 (O_308,N_18300,N_17515);
nand UO_309 (O_309,N_18476,N_18128);
nand UO_310 (O_310,N_16858,N_19434);
and UO_311 (O_311,N_17072,N_17307);
nor UO_312 (O_312,N_18851,N_16906);
or UO_313 (O_313,N_17074,N_18971);
nor UO_314 (O_314,N_18712,N_18650);
xnor UO_315 (O_315,N_19840,N_16804);
or UO_316 (O_316,N_19493,N_18516);
nor UO_317 (O_317,N_19357,N_19371);
nand UO_318 (O_318,N_18890,N_16216);
and UO_319 (O_319,N_16539,N_16728);
or UO_320 (O_320,N_19115,N_19743);
or UO_321 (O_321,N_16989,N_17498);
nand UO_322 (O_322,N_16209,N_16333);
nand UO_323 (O_323,N_17260,N_16511);
and UO_324 (O_324,N_18906,N_17998);
xnor UO_325 (O_325,N_18704,N_18728);
nor UO_326 (O_326,N_17547,N_17049);
or UO_327 (O_327,N_16682,N_17550);
nand UO_328 (O_328,N_17492,N_16349);
xor UO_329 (O_329,N_16913,N_16921);
and UO_330 (O_330,N_16118,N_18796);
xnor UO_331 (O_331,N_18849,N_16515);
xnor UO_332 (O_332,N_19621,N_18784);
nand UO_333 (O_333,N_18068,N_19395);
xor UO_334 (O_334,N_16519,N_17068);
and UO_335 (O_335,N_16208,N_19501);
or UO_336 (O_336,N_18120,N_17933);
and UO_337 (O_337,N_17750,N_18031);
nand UO_338 (O_338,N_18218,N_16971);
nor UO_339 (O_339,N_17875,N_18830);
xor UO_340 (O_340,N_17435,N_18486);
nand UO_341 (O_341,N_16371,N_18881);
or UO_342 (O_342,N_18556,N_19573);
and UO_343 (O_343,N_17339,N_16271);
nand UO_344 (O_344,N_19531,N_18477);
nor UO_345 (O_345,N_17473,N_19650);
xnor UO_346 (O_346,N_17782,N_17097);
xor UO_347 (O_347,N_17196,N_19639);
xnor UO_348 (O_348,N_16688,N_19424);
or UO_349 (O_349,N_19830,N_16968);
xor UO_350 (O_350,N_16748,N_17342);
nor UO_351 (O_351,N_19566,N_19505);
xor UO_352 (O_352,N_19054,N_17610);
nor UO_353 (O_353,N_18769,N_16268);
xnor UO_354 (O_354,N_16026,N_19177);
nand UO_355 (O_355,N_19841,N_16132);
nor UO_356 (O_356,N_16676,N_19297);
or UO_357 (O_357,N_16622,N_19871);
nand UO_358 (O_358,N_16556,N_16440);
nand UO_359 (O_359,N_18318,N_17412);
xor UO_360 (O_360,N_18954,N_18583);
xnor UO_361 (O_361,N_16963,N_16325);
or UO_362 (O_362,N_19504,N_17425);
nor UO_363 (O_363,N_19310,N_18150);
xnor UO_364 (O_364,N_18144,N_18786);
nand UO_365 (O_365,N_16551,N_17399);
nor UO_366 (O_366,N_16934,N_17112);
nand UO_367 (O_367,N_18366,N_18724);
xnor UO_368 (O_368,N_19216,N_19819);
nor UO_369 (O_369,N_17681,N_19187);
xor UO_370 (O_370,N_19971,N_16893);
or UO_371 (O_371,N_16217,N_16323);
nor UO_372 (O_372,N_17836,N_18635);
nor UO_373 (O_373,N_18018,N_17313);
nand UO_374 (O_374,N_17271,N_17619);
nand UO_375 (O_375,N_19375,N_16892);
or UO_376 (O_376,N_18311,N_16399);
and UO_377 (O_377,N_16171,N_19085);
nor UO_378 (O_378,N_16331,N_18241);
xnor UO_379 (O_379,N_17214,N_19008);
xor UO_380 (O_380,N_17463,N_18716);
nand UO_381 (O_381,N_17618,N_19321);
nand UO_382 (O_382,N_18973,N_19406);
xor UO_383 (O_383,N_16266,N_18248);
nand UO_384 (O_384,N_19784,N_19666);
xnor UO_385 (O_385,N_19688,N_16811);
or UO_386 (O_386,N_17643,N_19484);
xor UO_387 (O_387,N_19243,N_16360);
or UO_388 (O_388,N_18874,N_16572);
or UO_389 (O_389,N_16103,N_18878);
nand UO_390 (O_390,N_19539,N_18288);
xnor UO_391 (O_391,N_18345,N_16228);
nor UO_392 (O_392,N_19726,N_19594);
nand UO_393 (O_393,N_16273,N_19926);
xnor UO_394 (O_394,N_19454,N_18000);
xor UO_395 (O_395,N_19031,N_17736);
and UO_396 (O_396,N_16015,N_19407);
nor UO_397 (O_397,N_17053,N_16798);
nand UO_398 (O_398,N_16687,N_18508);
nand UO_399 (O_399,N_18932,N_17730);
xnor UO_400 (O_400,N_16970,N_16377);
nand UO_401 (O_401,N_17728,N_16326);
xor UO_402 (O_402,N_17641,N_18072);
nor UO_403 (O_403,N_17696,N_19433);
nor UO_404 (O_404,N_17804,N_17400);
or UO_405 (O_405,N_17691,N_17548);
xor UO_406 (O_406,N_19738,N_16063);
or UO_407 (O_407,N_17520,N_17297);
xor UO_408 (O_408,N_19584,N_18591);
nand UO_409 (O_409,N_19535,N_16183);
nor UO_410 (O_410,N_17267,N_19027);
and UO_411 (O_411,N_18449,N_18023);
nand UO_412 (O_412,N_19127,N_19609);
xnor UO_413 (O_413,N_19481,N_17322);
or UO_414 (O_414,N_17756,N_18548);
xor UO_415 (O_415,N_18417,N_18996);
nor UO_416 (O_416,N_17350,N_17088);
nor UO_417 (O_417,N_17598,N_16385);
and UO_418 (O_418,N_18439,N_16916);
nor UO_419 (O_419,N_18075,N_17486);
nand UO_420 (O_420,N_17236,N_19999);
or UO_421 (O_421,N_19736,N_17540);
nand UO_422 (O_422,N_18938,N_18596);
or UO_423 (O_423,N_19732,N_17438);
xnor UO_424 (O_424,N_19358,N_18638);
or UO_425 (O_425,N_18239,N_17557);
and UO_426 (O_426,N_18719,N_17357);
nand UO_427 (O_427,N_18586,N_18765);
xor UO_428 (O_428,N_19274,N_17461);
or UO_429 (O_429,N_16656,N_17496);
or UO_430 (O_430,N_18662,N_17531);
nor UO_431 (O_431,N_19426,N_17795);
nor UO_432 (O_432,N_17101,N_16032);
nor UO_433 (O_433,N_19061,N_19388);
xnor UO_434 (O_434,N_16501,N_16885);
nand UO_435 (O_435,N_18357,N_16991);
xor UO_436 (O_436,N_16530,N_17909);
xor UO_437 (O_437,N_16235,N_19197);
nand UO_438 (O_438,N_17482,N_18065);
nor UO_439 (O_439,N_19403,N_19618);
nand UO_440 (O_440,N_16696,N_18130);
nand UO_441 (O_441,N_17866,N_18660);
nor UO_442 (O_442,N_18183,N_17674);
or UO_443 (O_443,N_16131,N_16367);
xnor UO_444 (O_444,N_16929,N_16820);
xnor UO_445 (O_445,N_16151,N_18616);
nand UO_446 (O_446,N_18727,N_16806);
nor UO_447 (O_447,N_16842,N_19282);
xnor UO_448 (O_448,N_18386,N_19910);
nor UO_449 (O_449,N_17033,N_17778);
or UO_450 (O_450,N_19544,N_16566);
nor UO_451 (O_451,N_19521,N_18602);
or UO_452 (O_452,N_19253,N_19922);
nor UO_453 (O_453,N_16099,N_19016);
and UO_454 (O_454,N_17390,N_18415);
nand UO_455 (O_455,N_19414,N_17881);
nand UO_456 (O_456,N_17856,N_17740);
and UO_457 (O_457,N_17152,N_19112);
nand UO_458 (O_458,N_18904,N_18778);
and UO_459 (O_459,N_19116,N_16608);
and UO_460 (O_460,N_18572,N_19023);
xnor UO_461 (O_461,N_16562,N_16559);
or UO_462 (O_462,N_19637,N_19155);
xnor UO_463 (O_463,N_19951,N_16236);
and UO_464 (O_464,N_17355,N_18803);
and UO_465 (O_465,N_19619,N_17832);
xnor UO_466 (O_466,N_17414,N_16056);
nor UO_467 (O_467,N_19546,N_19548);
nor UO_468 (O_468,N_19002,N_17661);
nand UO_469 (O_469,N_18462,N_18585);
or UO_470 (O_470,N_18636,N_19045);
nor UO_471 (O_471,N_18615,N_18731);
xor UO_472 (O_472,N_18394,N_17424);
or UO_473 (O_473,N_18289,N_19209);
nand UO_474 (O_474,N_18752,N_19880);
nor UO_475 (O_475,N_19402,N_18515);
and UO_476 (O_476,N_16615,N_18715);
or UO_477 (O_477,N_18445,N_17493);
nor UO_478 (O_478,N_17940,N_18058);
xor UO_479 (O_479,N_16073,N_17284);
and UO_480 (O_480,N_18303,N_19171);
nand UO_481 (O_481,N_17253,N_18665);
or UO_482 (O_482,N_19050,N_17821);
nor UO_483 (O_483,N_18606,N_19029);
and UO_484 (O_484,N_19042,N_18702);
xnor UO_485 (O_485,N_17601,N_18683);
nor UO_486 (O_486,N_17734,N_17319);
or UO_487 (O_487,N_17041,N_17283);
or UO_488 (O_488,N_16050,N_19205);
nand UO_489 (O_489,N_17727,N_17504);
xnor UO_490 (O_490,N_17212,N_18514);
and UO_491 (O_491,N_18922,N_16348);
xor UO_492 (O_492,N_17221,N_17062);
nor UO_493 (O_493,N_17715,N_19086);
nor UO_494 (O_494,N_19716,N_16462);
nor UO_495 (O_495,N_19364,N_19160);
or UO_496 (O_496,N_18399,N_18389);
or UO_497 (O_497,N_17953,N_18518);
or UO_498 (O_498,N_19467,N_17170);
nand UO_499 (O_499,N_18603,N_18519);
or UO_500 (O_500,N_19708,N_18975);
nor UO_501 (O_501,N_17890,N_19455);
and UO_502 (O_502,N_18396,N_19849);
xnor UO_503 (O_503,N_17814,N_16049);
and UO_504 (O_504,N_19777,N_18159);
and UO_505 (O_505,N_19431,N_16795);
nor UO_506 (O_506,N_16552,N_19220);
nor UO_507 (O_507,N_17201,N_17361);
xor UO_508 (O_508,N_17565,N_17604);
and UO_509 (O_509,N_19826,N_18017);
and UO_510 (O_510,N_19928,N_19118);
nand UO_511 (O_511,N_17120,N_18475);
nor UO_512 (O_512,N_18779,N_16352);
nand UO_513 (O_513,N_18005,N_19477);
nand UO_514 (O_514,N_16079,N_16409);
xnor UO_515 (O_515,N_17823,N_18206);
xor UO_516 (O_516,N_16897,N_16489);
nand UO_517 (O_517,N_16197,N_17747);
nand UO_518 (O_518,N_18485,N_18649);
and UO_519 (O_519,N_19485,N_18267);
nor UO_520 (O_520,N_19842,N_18272);
and UO_521 (O_521,N_16576,N_17981);
nor UO_522 (O_522,N_18595,N_19874);
and UO_523 (O_523,N_16786,N_19377);
xnor UO_524 (O_524,N_17553,N_16825);
xnor UO_525 (O_525,N_17710,N_16353);
nor UO_526 (O_526,N_16711,N_19676);
xor UO_527 (O_527,N_18413,N_17944);
xor UO_528 (O_528,N_19664,N_17882);
nand UO_529 (O_529,N_18369,N_18102);
or UO_530 (O_530,N_17693,N_18943);
nand UO_531 (O_531,N_16279,N_17016);
or UO_532 (O_532,N_18380,N_18322);
xnor UO_533 (O_533,N_16291,N_16771);
or UO_534 (O_534,N_18576,N_19503);
or UO_535 (O_535,N_18542,N_16443);
nand UO_536 (O_536,N_19096,N_18895);
nand UO_537 (O_537,N_18094,N_18927);
and UO_538 (O_538,N_16524,N_16114);
nor UO_539 (O_539,N_16952,N_16589);
xnor UO_540 (O_540,N_18658,N_19298);
nand UO_541 (O_541,N_19361,N_16713);
and UO_542 (O_542,N_18555,N_19869);
or UO_543 (O_543,N_18494,N_18620);
and UO_544 (O_544,N_16332,N_18378);
or UO_545 (O_545,N_17491,N_16115);
or UO_546 (O_546,N_18819,N_17837);
xnor UO_547 (O_547,N_17979,N_19190);
or UO_548 (O_548,N_19144,N_16650);
nand UO_549 (O_549,N_19678,N_16659);
nand UO_550 (O_550,N_16174,N_19191);
xor UO_551 (O_551,N_18982,N_16983);
nor UO_552 (O_552,N_19863,N_19975);
and UO_553 (O_553,N_16846,N_18006);
nor UO_554 (O_554,N_18492,N_17830);
and UO_555 (O_555,N_19911,N_17676);
and UO_556 (O_556,N_18243,N_16756);
nand UO_557 (O_557,N_17690,N_18544);
and UO_558 (O_558,N_18738,N_18479);
xnor UO_559 (O_559,N_18139,N_16280);
or UO_560 (O_560,N_19935,N_17181);
nor UO_561 (O_561,N_18437,N_18203);
and UO_562 (O_562,N_17349,N_18846);
and UO_563 (O_563,N_16974,N_18260);
nand UO_564 (O_564,N_18409,N_17927);
nor UO_565 (O_565,N_17285,N_18008);
and UO_566 (O_566,N_19834,N_16296);
and UO_567 (O_567,N_17059,N_19675);
or UO_568 (O_568,N_17429,N_17910);
or UO_569 (O_569,N_18788,N_17472);
xor UO_570 (O_570,N_18410,N_17907);
nand UO_571 (O_571,N_19342,N_16701);
and UO_572 (O_572,N_19183,N_19906);
nor UO_573 (O_573,N_18362,N_18392);
nor UO_574 (O_574,N_18534,N_19955);
nor UO_575 (O_575,N_16910,N_17187);
nand UO_576 (O_576,N_17644,N_16354);
xor UO_577 (O_577,N_16621,N_18319);
nor UO_578 (O_578,N_19550,N_17047);
and UO_579 (O_579,N_19288,N_19984);
nor UO_580 (O_580,N_19170,N_17073);
nand UO_581 (O_581,N_18153,N_17692);
nor UO_582 (O_582,N_16598,N_17085);
nand UO_583 (O_583,N_16330,N_19645);
nand UO_584 (O_584,N_16090,N_16415);
nor UO_585 (O_585,N_17538,N_19790);
xnor UO_586 (O_586,N_18705,N_17695);
nor UO_587 (O_587,N_17569,N_18651);
nor UO_588 (O_588,N_18834,N_17764);
or UO_589 (O_589,N_16731,N_18165);
xnor UO_590 (O_590,N_19583,N_16500);
xor UO_591 (O_591,N_19865,N_19895);
nand UO_592 (O_592,N_18377,N_19679);
xnor UO_593 (O_593,N_16967,N_17451);
nor UO_594 (O_594,N_16136,N_18135);
xnor UO_595 (O_595,N_17190,N_17393);
nor UO_596 (O_596,N_18875,N_18052);
nand UO_597 (O_597,N_16109,N_18220);
xnor UO_598 (O_598,N_18090,N_17840);
nand UO_599 (O_599,N_16987,N_17254);
nor UO_600 (O_600,N_19745,N_17642);
xnor UO_601 (O_601,N_19750,N_16493);
xnor UO_602 (O_602,N_18639,N_16907);
nor UO_603 (O_603,N_18945,N_17228);
and UO_604 (O_604,N_17365,N_17572);
nor UO_605 (O_605,N_16708,N_16211);
and UO_606 (O_606,N_16071,N_19596);
nor UO_607 (O_607,N_17363,N_17266);
nor UO_608 (O_608,N_17176,N_18678);
xnor UO_609 (O_609,N_17743,N_18114);
nor UO_610 (O_610,N_16240,N_17010);
or UO_611 (O_611,N_16230,N_17675);
nor UO_612 (O_612,N_16850,N_17971);
and UO_613 (O_613,N_16849,N_17525);
nand UO_614 (O_614,N_16666,N_18593);
or UO_615 (O_615,N_16944,N_16600);
nand UO_616 (O_616,N_19056,N_16597);
xnor UO_617 (O_617,N_18049,N_17257);
xor UO_618 (O_618,N_18653,N_19239);
and UO_619 (O_619,N_16557,N_16528);
or UO_620 (O_620,N_19519,N_19252);
nand UO_621 (O_621,N_19079,N_18148);
and UO_622 (O_622,N_19773,N_18891);
or UO_623 (O_623,N_18446,N_17215);
or UO_624 (O_624,N_17519,N_16476);
nor UO_625 (O_625,N_17323,N_19512);
or UO_626 (O_626,N_17029,N_18327);
xor UO_627 (O_627,N_18295,N_19595);
nand UO_628 (O_628,N_16664,N_19698);
xnor UO_629 (O_629,N_18900,N_16100);
xnor UO_630 (O_630,N_17789,N_18914);
or UO_631 (O_631,N_17773,N_16554);
nor UO_632 (O_632,N_19510,N_16229);
and UO_633 (O_633,N_18789,N_16965);
and UO_634 (O_634,N_16772,N_18235);
nand UO_635 (O_635,N_19261,N_18127);
nand UO_636 (O_636,N_17769,N_19552);
or UO_637 (O_637,N_17699,N_18109);
nand UO_638 (O_638,N_18214,N_16652);
or UO_639 (O_639,N_17058,N_19916);
xor UO_640 (O_640,N_18027,N_16898);
nor UO_641 (O_641,N_16274,N_17380);
and UO_642 (O_642,N_19782,N_16226);
xnor UO_643 (O_643,N_19173,N_19221);
or UO_644 (O_644,N_16678,N_17024);
and UO_645 (O_645,N_19800,N_17700);
xor UO_646 (O_646,N_19327,N_18338);
and UO_647 (O_647,N_18368,N_19757);
and UO_648 (O_648,N_17457,N_16436);
nor UO_649 (O_649,N_16380,N_17327);
and UO_650 (O_650,N_19279,N_17044);
nor UO_651 (O_651,N_18569,N_18785);
nand UO_652 (O_652,N_17497,N_18482);
nand UO_653 (O_653,N_17100,N_17110);
xnor UO_654 (O_654,N_17975,N_19381);
xor UO_655 (O_655,N_18088,N_19741);
nand UO_656 (O_656,N_17687,N_19360);
and UO_657 (O_657,N_18628,N_17801);
and UO_658 (O_658,N_17552,N_17511);
and UO_659 (O_659,N_19425,N_19242);
or UO_660 (O_660,N_17149,N_16588);
or UO_661 (O_661,N_17159,N_19036);
xor UO_662 (O_662,N_16408,N_16427);
or UO_663 (O_663,N_18339,N_18820);
xnor UO_664 (O_664,N_18459,N_19538);
nor UO_665 (O_665,N_16361,N_16061);
nand UO_666 (O_666,N_17802,N_18232);
nor UO_667 (O_667,N_19677,N_19661);
nor UO_668 (O_668,N_19847,N_16072);
nor UO_669 (O_669,N_16060,N_19670);
or UO_670 (O_670,N_16135,N_17812);
and UO_671 (O_671,N_17820,N_18771);
xnor UO_672 (O_672,N_16222,N_17537);
nor UO_673 (O_673,N_19130,N_16485);
nand UO_674 (O_674,N_19139,N_18258);
and UO_675 (O_675,N_17761,N_17846);
and UO_676 (O_676,N_17065,N_17023);
nor UO_677 (O_677,N_19769,N_19199);
xnor UO_678 (O_678,N_17061,N_18543);
nor UO_679 (O_679,N_19272,N_18997);
xnor UO_680 (O_680,N_18035,N_17413);
xnor UO_681 (O_681,N_18503,N_18955);
and UO_682 (O_682,N_17488,N_16094);
nor UO_683 (O_683,N_16699,N_17817);
nand UO_684 (O_684,N_17475,N_18313);
nand UO_685 (O_685,N_19462,N_18019);
or UO_686 (O_686,N_16190,N_19165);
nor UO_687 (O_687,N_17983,N_19915);
nor UO_688 (O_688,N_18013,N_16640);
or UO_689 (O_689,N_17039,N_17955);
nor UO_690 (O_690,N_16162,N_18096);
or UO_691 (O_691,N_19835,N_18395);
and UO_692 (O_692,N_18876,N_18189);
nand UO_693 (O_693,N_17031,N_19083);
nand UO_694 (O_694,N_16807,N_19568);
or UO_695 (O_695,N_18202,N_17440);
nand UO_696 (O_696,N_18773,N_16570);
nor UO_697 (O_697,N_17108,N_19959);
nor UO_698 (O_698,N_16924,N_18330);
xor UO_699 (O_699,N_19706,N_17993);
nand UO_700 (O_700,N_16116,N_19991);
nor UO_701 (O_701,N_19946,N_19084);
nand UO_702 (O_702,N_19390,N_18902);
xor UO_703 (O_703,N_18046,N_16203);
or UO_704 (O_704,N_19456,N_19179);
and UO_705 (O_705,N_18020,N_19469);
or UO_706 (O_706,N_16492,N_16382);
and UO_707 (O_707,N_18452,N_18898);
nand UO_708 (O_708,N_19174,N_16591);
or UO_709 (O_709,N_19125,N_16774);
nor UO_710 (O_710,N_18775,N_18761);
and UO_711 (O_711,N_18540,N_17166);
or UO_712 (O_712,N_18122,N_17523);
or UO_713 (O_713,N_19058,N_19543);
xor UO_714 (O_714,N_19641,N_17600);
and UO_715 (O_715,N_16064,N_18942);
and UO_716 (O_716,N_17450,N_16142);
or UO_717 (O_717,N_18610,N_17426);
xnor UO_718 (O_718,N_16080,N_19654);
xor UO_719 (O_719,N_18745,N_18222);
nor UO_720 (O_720,N_18614,N_17204);
nor UO_721 (O_721,N_19124,N_18541);
xor UO_722 (O_722,N_16945,N_18175);
or UO_723 (O_723,N_17238,N_17337);
or UO_724 (O_724,N_18372,N_19472);
nor UO_725 (O_725,N_17078,N_18294);
and UO_726 (O_726,N_17954,N_16390);
nor UO_727 (O_727,N_17776,N_17209);
xor UO_728 (O_728,N_17002,N_18199);
nand UO_729 (O_729,N_17855,N_19471);
and UO_730 (O_730,N_18753,N_17864);
nor UO_731 (O_731,N_18986,N_16757);
nand UO_732 (O_732,N_16445,N_16872);
nor UO_733 (O_733,N_16370,N_16984);
and UO_734 (O_734,N_17663,N_19513);
nor UO_735 (O_735,N_19153,N_18456);
or UO_736 (O_736,N_18265,N_16959);
or UO_737 (O_737,N_18984,N_19475);
nor UO_738 (O_738,N_16477,N_18161);
and UO_739 (O_739,N_19020,N_18879);
nand UO_740 (O_740,N_17850,N_16874);
nor UO_741 (O_741,N_17624,N_17703);
and UO_742 (O_742,N_18101,N_18517);
or UO_743 (O_743,N_18843,N_17237);
nor UO_744 (O_744,N_16192,N_17711);
and UO_745 (O_745,N_16722,N_16902);
or UO_746 (O_746,N_18717,N_17913);
nand UO_747 (O_747,N_17227,N_17035);
nand UO_748 (O_748,N_17401,N_17915);
and UO_749 (O_749,N_16307,N_17106);
and UO_750 (O_750,N_19593,N_19435);
xnor UO_751 (O_751,N_16815,N_16366);
nor UO_752 (O_752,N_17682,N_18873);
nor UO_753 (O_753,N_16147,N_18081);
nor UO_754 (O_754,N_18525,N_19289);
nor UO_755 (O_755,N_19035,N_16294);
xnor UO_756 (O_756,N_19646,N_19275);
or UO_757 (O_757,N_19260,N_18860);
and UO_758 (O_758,N_19401,N_16721);
xnor UO_759 (O_759,N_18115,N_16579);
xnor UO_760 (O_760,N_19293,N_19794);
and UO_761 (O_761,N_16939,N_18346);
and UO_762 (O_762,N_16133,N_17510);
and UO_763 (O_763,N_18965,N_16498);
and UO_764 (O_764,N_16834,N_18297);
and UO_765 (O_765,N_16882,N_19796);
xor UO_766 (O_766,N_18215,N_19520);
nor UO_767 (O_767,N_16177,N_16990);
and UO_768 (O_768,N_16782,N_18928);
and UO_769 (O_769,N_18552,N_19159);
xor UO_770 (O_770,N_16000,N_17324);
and UO_771 (O_771,N_19121,N_17362);
and UO_772 (O_772,N_19532,N_19857);
and UO_773 (O_773,N_16642,N_19620);
nor UO_774 (O_774,N_16251,N_17147);
nor UO_775 (O_775,N_17532,N_18723);
nand UO_776 (O_776,N_17021,N_16523);
nand UO_777 (O_777,N_17871,N_18558);
nand UO_778 (O_778,N_19443,N_19255);
nor UO_779 (O_779,N_18822,N_17990);
or UO_780 (O_780,N_16337,N_16698);
nand UO_781 (O_781,N_19250,N_18656);
nand UO_782 (O_782,N_18009,N_19576);
or UO_783 (O_783,N_16793,N_18797);
nand UO_784 (O_784,N_18487,N_17976);
and UO_785 (O_785,N_17128,N_18430);
nand UO_786 (O_786,N_16723,N_17854);
and UO_787 (O_787,N_18249,N_16690);
nand UO_788 (O_788,N_17920,N_18520);
xnor UO_789 (O_789,N_19057,N_16156);
or UO_790 (O_790,N_18221,N_18074);
and UO_791 (O_791,N_18489,N_17718);
nand UO_792 (O_792,N_17825,N_16168);
or UO_793 (O_793,N_19126,N_16848);
nand UO_794 (O_794,N_19904,N_19730);
xor UO_795 (O_795,N_17951,N_17046);
xor UO_796 (O_796,N_18974,N_16213);
xnor UO_797 (O_797,N_17943,N_17111);
nor UO_798 (O_798,N_19466,N_18252);
nor UO_799 (O_799,N_16727,N_16242);
or UO_800 (O_800,N_16558,N_17013);
xor UO_801 (O_801,N_19108,N_16706);
or UO_802 (O_802,N_19832,N_16263);
nand UO_803 (O_803,N_16843,N_18281);
and UO_804 (O_804,N_17326,N_16150);
xor UO_805 (O_805,N_19803,N_18298);
or UO_806 (O_806,N_17431,N_16027);
nor UO_807 (O_807,N_17994,N_16277);
or UO_808 (O_808,N_19248,N_19506);
nor UO_809 (O_809,N_19634,N_16641);
or UO_810 (O_810,N_19862,N_19983);
or UO_811 (O_811,N_16146,N_19683);
nand UO_812 (O_812,N_19617,N_18448);
or UO_813 (O_813,N_17458,N_19071);
xnor UO_814 (O_814,N_16092,N_16117);
or UO_815 (O_815,N_17751,N_16021);
nor UO_816 (O_816,N_16181,N_16450);
or UO_817 (O_817,N_16504,N_19235);
nor UO_818 (O_818,N_19940,N_17811);
nor UO_819 (O_819,N_16683,N_17242);
xnor UO_820 (O_820,N_16571,N_19814);
and UO_821 (O_821,N_19783,N_19051);
or UO_822 (O_822,N_17507,N_16860);
and UO_823 (O_823,N_18809,N_16497);
nor UO_824 (O_824,N_16220,N_18207);
or UO_825 (O_825,N_17991,N_17512);
nand UO_826 (O_826,N_16459,N_16502);
nand UO_827 (O_827,N_19611,N_16086);
nand UO_828 (O_828,N_16112,N_16074);
or UO_829 (O_829,N_16452,N_17148);
nand UO_830 (O_830,N_16904,N_16261);
nand UO_831 (O_831,N_17125,N_18379);
nor UO_832 (O_832,N_17145,N_18633);
and UO_833 (O_833,N_17842,N_19626);
xor UO_834 (O_834,N_17211,N_16649);
or UO_835 (O_835,N_19816,N_19331);
nand UO_836 (O_836,N_18132,N_17247);
xor UO_837 (O_837,N_19167,N_18385);
nor UO_838 (O_838,N_19684,N_16300);
or UO_839 (O_839,N_16870,N_19665);
and UO_840 (O_840,N_16679,N_16616);
nor UO_841 (O_841,N_18805,N_19022);
nor UO_842 (O_842,N_19509,N_19257);
or UO_843 (O_843,N_18697,N_18733);
xor UO_844 (O_844,N_17839,N_17753);
xnor UO_845 (O_845,N_16460,N_17580);
nand UO_846 (O_846,N_17726,N_16194);
nand UO_847 (O_847,N_19148,N_18067);
xor UO_848 (O_848,N_19936,N_17092);
and UO_849 (O_849,N_17224,N_18190);
and UO_850 (O_850,N_18824,N_17645);
or UO_851 (O_851,N_19368,N_19797);
nor UO_852 (O_852,N_17172,N_18040);
xnor UO_853 (O_853,N_16249,N_17606);
or UO_854 (O_854,N_19349,N_17419);
nand UO_855 (O_855,N_16110,N_17015);
nand UO_856 (O_856,N_16960,N_16516);
nand UO_857 (O_857,N_16101,N_17217);
and UO_858 (O_858,N_18168,N_17916);
nor UO_859 (O_859,N_19963,N_19440);
xnor UO_860 (O_860,N_17347,N_16388);
nor UO_861 (O_861,N_19460,N_16631);
nor UO_862 (O_862,N_17430,N_16033);
and UO_863 (O_863,N_17888,N_19579);
xor UO_864 (O_864,N_17609,N_17014);
nor UO_865 (O_865,N_18526,N_19912);
or UO_866 (O_866,N_16007,N_17596);
nand UO_867 (O_867,N_18370,N_16827);
nor UO_868 (O_868,N_17707,N_19561);
nor UO_869 (O_869,N_17573,N_19762);
xnor UO_870 (O_870,N_16265,N_16144);
xnor UO_871 (O_871,N_17278,N_16947);
or UO_872 (O_872,N_17103,N_18277);
or UO_873 (O_873,N_16905,N_17294);
nand UO_874 (O_874,N_18003,N_16880);
nand UO_875 (O_875,N_18250,N_19182);
xnor UO_876 (O_876,N_19222,N_19311);
xor UO_877 (O_877,N_16368,N_16439);
nand UO_878 (O_878,N_16816,N_18862);
nor UO_879 (O_879,N_18253,N_19268);
and UO_880 (O_880,N_19977,N_19799);
xor UO_881 (O_881,N_17077,N_18619);
nor UO_882 (O_882,N_16886,N_17367);
xnor UO_883 (O_883,N_18886,N_18960);
xor UO_884 (O_884,N_18237,N_17716);
and UO_885 (O_885,N_16547,N_16845);
or UO_886 (O_886,N_16179,N_19449);
and UO_887 (O_887,N_18501,N_17742);
or UO_888 (O_888,N_18699,N_19536);
or UO_889 (O_889,N_17411,N_19994);
nand UO_890 (O_890,N_16707,N_18529);
nor UO_891 (O_891,N_17075,N_17834);
nand UO_892 (O_892,N_17004,N_18907);
and UO_893 (O_893,N_18622,N_17667);
xor UO_894 (O_894,N_19062,N_18913);
xnor UO_895 (O_895,N_19369,N_16760);
xor UO_896 (O_896,N_18729,N_16766);
and UO_897 (O_897,N_18859,N_16900);
nor UO_898 (O_898,N_18453,N_16077);
nand UO_899 (O_899,N_17568,N_17303);
nand UO_900 (O_900,N_17048,N_17459);
nand UO_901 (O_901,N_17168,N_17527);
or UO_902 (O_902,N_16184,N_19416);
xor UO_903 (O_903,N_18999,N_19140);
nor UO_904 (O_904,N_19237,N_17932);
and UO_905 (O_905,N_16343,N_16620);
and UO_906 (O_906,N_19423,N_16106);
nand UO_907 (O_907,N_17891,N_18269);
xor UO_908 (O_908,N_18613,N_16927);
or UO_909 (O_909,N_16036,N_17433);
and UO_910 (O_910,N_16324,N_16735);
nor UO_911 (O_911,N_16734,N_18831);
and UO_912 (O_912,N_17615,N_19158);
or UO_913 (O_913,N_16047,N_16507);
xor UO_914 (O_914,N_18022,N_17011);
xnor UO_915 (O_915,N_17599,N_19212);
and UO_916 (O_916,N_16374,N_19530);
or UO_917 (O_917,N_19647,N_16862);
and UO_918 (O_918,N_17263,N_18892);
or UO_919 (O_919,N_18138,N_19452);
nor UO_920 (O_920,N_16297,N_19802);
nor UO_921 (O_921,N_19658,N_17250);
xnor UO_922 (O_922,N_18872,N_18178);
and UO_923 (O_923,N_19353,N_19601);
nor UO_924 (O_924,N_16888,N_19597);
xor UO_925 (O_925,N_16076,N_18381);
and UO_926 (O_926,N_16876,N_16883);
or UO_927 (O_927,N_16160,N_16028);
xnor UO_928 (O_928,N_17865,N_19240);
or UO_929 (O_929,N_19422,N_16457);
xor UO_930 (O_930,N_16668,N_16334);
nor UO_931 (O_931,N_16344,N_19877);
or UO_932 (O_932,N_17318,N_19287);
and UO_933 (O_933,N_18869,N_17387);
or UO_934 (O_934,N_16606,N_17852);
nand UO_935 (O_935,N_19427,N_16494);
and UO_936 (O_936,N_19109,N_19515);
nand UO_937 (O_937,N_18044,N_18937);
or UO_938 (O_938,N_16428,N_19891);
nand UO_939 (O_939,N_19330,N_16270);
and UO_940 (O_940,N_16234,N_16412);
nand UO_941 (O_941,N_19026,N_18659);
nor UO_942 (O_942,N_19953,N_17967);
xnor UO_943 (O_943,N_16891,N_16646);
nor UO_944 (O_944,N_16543,N_16444);
xnor UO_945 (O_945,N_17985,N_16012);
or UO_946 (O_946,N_16373,N_18577);
nand UO_947 (O_947,N_17611,N_19105);
or UO_948 (O_948,N_17001,N_18755);
xor UO_949 (O_949,N_16899,N_18837);
or UO_950 (O_950,N_18238,N_18416);
or UO_951 (O_951,N_18306,N_19204);
or UO_952 (O_952,N_16473,N_16903);
nor UO_953 (O_953,N_16536,N_17356);
and UO_954 (O_954,N_16081,N_18836);
and UO_955 (O_955,N_18425,N_18496);
and UO_956 (O_956,N_19316,N_17973);
nor UO_957 (O_957,N_16335,N_16070);
and UO_958 (O_958,N_17919,N_18539);
and UO_959 (O_959,N_17105,N_19728);
nor UO_960 (O_960,N_17772,N_19565);
nand UO_961 (O_961,N_19122,N_19582);
or UO_962 (O_962,N_16948,N_17258);
nand UO_963 (O_963,N_18495,N_19157);
nor UO_964 (O_964,N_17797,N_16066);
and UO_965 (O_965,N_17779,N_16215);
and UO_966 (O_966,N_17841,N_16435);
xnor UO_967 (O_967,N_17868,N_18012);
and UO_968 (O_968,N_19043,N_17545);
or UO_969 (O_969,N_18645,N_18802);
or UO_970 (O_970,N_16006,N_18618);
nand UO_971 (O_971,N_16346,N_17317);
nand UO_972 (O_972,N_16338,N_16879);
or UO_973 (O_973,N_19724,N_16763);
nor UO_974 (O_974,N_19136,N_19194);
xor UO_975 (O_975,N_18350,N_16189);
nand UO_976 (O_976,N_18435,N_18845);
and UO_977 (O_977,N_17900,N_19793);
nor UO_978 (O_978,N_17456,N_18498);
or UO_979 (O_979,N_18483,N_19556);
and UO_980 (O_980,N_16624,N_19884);
xor UO_981 (O_981,N_17295,N_19059);
nor UO_982 (O_982,N_17646,N_19875);
and UO_983 (O_983,N_16446,N_16283);
nand UO_984 (O_984,N_18562,N_19908);
or UO_985 (O_985,N_18940,N_17397);
nand UO_986 (O_986,N_19924,N_18608);
nand UO_987 (O_987,N_17689,N_19693);
and UO_988 (O_988,N_16644,N_18838);
xnor UO_989 (O_989,N_17358,N_18172);
nor UO_990 (O_990,N_16394,N_18283);
nor UO_991 (O_991,N_19754,N_16675);
and UO_992 (O_992,N_16736,N_19956);
nor UO_993 (O_993,N_18045,N_18037);
and UO_994 (O_994,N_18107,N_17583);
nor UO_995 (O_995,N_18432,N_17476);
xnor UO_996 (O_996,N_17197,N_17608);
xor UO_997 (O_997,N_17612,N_18225);
xnor UO_998 (O_998,N_17381,N_18864);
xnor UO_999 (O_999,N_17581,N_17308);
xnor UO_1000 (O_1000,N_19859,N_17558);
nand UO_1001 (O_1001,N_18781,N_17586);
or UO_1002 (O_1002,N_17860,N_16065);
or UO_1003 (O_1003,N_19547,N_18887);
nand UO_1004 (O_1004,N_19208,N_16468);
and UO_1005 (O_1005,N_16946,N_18034);
nor UO_1006 (O_1006,N_17406,N_16509);
nor UO_1007 (O_1007,N_18978,N_17026);
xor UO_1008 (O_1008,N_18812,N_16632);
and UO_1009 (O_1009,N_19101,N_19671);
nand UO_1010 (O_1010,N_19813,N_19882);
nor UO_1011 (O_1011,N_19723,N_17819);
or UO_1012 (O_1012,N_18234,N_19886);
nand UO_1013 (O_1013,N_17359,N_16741);
nand UO_1014 (O_1014,N_16973,N_17575);
or UO_1015 (O_1015,N_16395,N_19111);
nor UO_1016 (O_1016,N_16742,N_19499);
nor UO_1017 (O_1017,N_17897,N_16700);
and UO_1018 (O_1018,N_18793,N_19172);
or UO_1019 (O_1019,N_16980,N_19719);
or UO_1020 (O_1020,N_17874,N_18302);
nand UO_1021 (O_1021,N_17396,N_16364);
nor UO_1022 (O_1022,N_16025,N_17063);
and UO_1023 (O_1023,N_18491,N_19017);
and UO_1024 (O_1024,N_18991,N_17564);
and UO_1025 (O_1025,N_19968,N_19292);
or UO_1026 (O_1026,N_18979,N_17680);
and UO_1027 (O_1027,N_17947,N_17709);
nand UO_1028 (O_1028,N_17562,N_19178);
nor UO_1029 (O_1029,N_16267,N_16778);
and UO_1030 (O_1030,N_17306,N_19746);
xnor UO_1031 (O_1031,N_16098,N_18070);
and UO_1032 (O_1032,N_19603,N_19442);
nor UO_1033 (O_1033,N_17952,N_17560);
and UO_1034 (O_1034,N_17770,N_19733);
and UO_1035 (O_1035,N_19264,N_18043);
or UO_1036 (O_1036,N_18176,N_17405);
xnor UO_1037 (O_1037,N_18861,N_17514);
or UO_1038 (O_1038,N_16674,N_18196);
or UO_1039 (O_1039,N_19563,N_16139);
and UO_1040 (O_1040,N_16754,N_16293);
nand UO_1041 (O_1041,N_16269,N_19489);
xnor UO_1042 (O_1042,N_17566,N_17853);
or UO_1043 (O_1043,N_16159,N_19612);
or UO_1044 (O_1044,N_16120,N_16738);
or UO_1045 (O_1045,N_19598,N_17210);
nor UO_1046 (O_1046,N_16123,N_16895);
nand UO_1047 (O_1047,N_16464,N_19694);
or UO_1048 (O_1048,N_19533,N_19483);
and UO_1049 (O_1049,N_16938,N_16083);
xor UO_1050 (O_1050,N_16248,N_16153);
nor UO_1051 (O_1051,N_16491,N_19554);
nand UO_1052 (O_1052,N_19397,N_19482);
nor UO_1053 (O_1053,N_19021,N_19555);
or UO_1054 (O_1054,N_19018,N_16029);
nor UO_1055 (O_1055,N_17701,N_18850);
or UO_1056 (O_1056,N_17765,N_19347);
and UO_1057 (O_1057,N_19040,N_16628);
and UO_1058 (O_1058,N_18305,N_19372);
or UO_1059 (O_1059,N_17194,N_17638);
nand UO_1060 (O_1060,N_17045,N_19295);
and UO_1061 (O_1061,N_17500,N_19756);
nor UO_1062 (O_1062,N_17922,N_16759);
nor UO_1063 (O_1063,N_18497,N_18276);
or UO_1064 (O_1064,N_18682,N_17655);
or UO_1065 (O_1065,N_19323,N_17071);
nor UO_1066 (O_1066,N_19063,N_18291);
nand UO_1067 (O_1067,N_16286,N_16670);
nor UO_1068 (O_1068,N_19259,N_16585);
and UO_1069 (O_1069,N_18270,N_17659);
nand UO_1070 (O_1070,N_17372,N_18170);
nor UO_1071 (O_1071,N_17862,N_18532);
or UO_1072 (O_1072,N_18320,N_19103);
or UO_1073 (O_1073,N_17119,N_18352);
xor UO_1074 (O_1074,N_17849,N_17027);
nor UO_1075 (O_1075,N_17945,N_17410);
and UO_1076 (O_1076,N_16129,N_18143);
xnor UO_1077 (O_1077,N_18066,N_19186);
nand UO_1078 (O_1078,N_19254,N_18750);
nor UO_1079 (O_1079,N_17561,N_16908);
and UO_1080 (O_1080,N_18739,N_19419);
or UO_1081 (O_1081,N_17653,N_18762);
nand UO_1082 (O_1082,N_17052,N_19786);
or UO_1083 (O_1083,N_17631,N_17138);
xnor UO_1084 (O_1084,N_18640,N_19623);
and UO_1085 (O_1085,N_16121,N_17587);
and UO_1086 (O_1086,N_16137,N_19511);
nand UO_1087 (O_1087,N_16564,N_19969);
nand UO_1088 (O_1088,N_17383,N_16692);
or UO_1089 (O_1089,N_16088,N_18329);
and UO_1090 (O_1090,N_16881,N_18989);
xor UO_1091 (O_1091,N_16051,N_17213);
xor UO_1092 (O_1092,N_19391,N_16004);
nand UO_1093 (O_1093,N_17114,N_18599);
nand UO_1094 (O_1094,N_16569,N_16828);
or UO_1095 (O_1095,N_18054,N_17767);
or UO_1096 (O_1096,N_16802,N_17269);
xnor UO_1097 (O_1097,N_18563,N_17234);
xor UO_1098 (O_1098,N_18564,N_19285);
nor UO_1099 (O_1099,N_17183,N_16752);
and UO_1100 (O_1100,N_16733,N_17340);
or UO_1101 (O_1101,N_16812,N_18934);
xor UO_1102 (O_1102,N_17386,N_17754);
nor UO_1103 (O_1103,N_17844,N_18356);
xor UO_1104 (O_1104,N_19490,N_17344);
nor UO_1105 (O_1105,N_18696,N_19810);
and UO_1106 (O_1106,N_17529,N_16658);
or UO_1107 (O_1107,N_16481,N_18754);
nor UO_1108 (O_1108,N_19436,N_17961);
xor UO_1109 (O_1109,N_18839,N_17533);
or UO_1110 (O_1110,N_18464,N_16739);
nor UO_1111 (O_1111,N_17535,N_18655);
nor UO_1112 (O_1112,N_19649,N_19223);
nor UO_1113 (O_1113,N_16729,N_19614);
nand UO_1114 (O_1114,N_19458,N_18574);
nor UO_1115 (O_1115,N_19329,N_16375);
or UO_1116 (O_1116,N_17329,N_16955);
and UO_1117 (O_1117,N_17925,N_18588);
nor UO_1118 (O_1118,N_18155,N_19751);
and UO_1119 (O_1119,N_19067,N_17177);
nor UO_1120 (O_1120,N_18527,N_19943);
and UO_1121 (O_1121,N_16191,N_18568);
nor UO_1122 (O_1122,N_17434,N_18721);
and UO_1123 (O_1123,N_19428,N_16298);
nor UO_1124 (O_1124,N_16392,N_17816);
xor UO_1125 (O_1125,N_19412,N_16677);
xor UO_1126 (O_1126,N_17936,N_16758);
nand UO_1127 (O_1127,N_19106,N_16890);
xnor UO_1128 (O_1128,N_16568,N_19648);
xor UO_1129 (O_1129,N_19772,N_19858);
or UO_1130 (O_1130,N_17625,N_17799);
nand UO_1131 (O_1131,N_19947,N_17069);
or UO_1132 (O_1132,N_19077,N_18064);
nand UO_1133 (O_1133,N_17091,N_16545);
nand UO_1134 (O_1134,N_17678,N_17489);
nor UO_1135 (O_1135,N_17878,N_17530);
or UO_1136 (O_1136,N_19758,N_18332);
nor UO_1137 (O_1137,N_16084,N_18631);
xor UO_1138 (O_1138,N_17648,N_18083);
xor UO_1139 (O_1139,N_19976,N_17265);
nand UO_1140 (O_1140,N_17783,N_16691);
or UO_1141 (O_1141,N_19659,N_17233);
and UO_1142 (O_1142,N_18992,N_18361);
and UO_1143 (O_1143,N_16480,N_18612);
or UO_1144 (O_1144,N_18835,N_16278);
or UO_1145 (O_1145,N_16257,N_17241);
or UO_1146 (O_1146,N_19217,N_16567);
nand UO_1147 (O_1147,N_16857,N_18092);
and UO_1148 (O_1148,N_18594,N_18808);
nand UO_1149 (O_1149,N_19355,N_19523);
nor UO_1150 (O_1150,N_16609,N_18028);
nand UO_1151 (O_1151,N_16164,N_18694);
and UO_1152 (O_1152,N_18307,N_16108);
nand UO_1153 (O_1153,N_16141,N_19334);
and UO_1154 (O_1154,N_16949,N_17857);
nand UO_1155 (O_1155,N_16514,N_16214);
or UO_1156 (O_1156,N_18829,N_19313);
and UO_1157 (O_1157,N_18210,N_19640);
and UO_1158 (O_1158,N_18166,N_17188);
xor UO_1159 (O_1159,N_18597,N_19774);
or UO_1160 (O_1160,N_17771,N_17243);
and UO_1161 (O_1161,N_19494,N_19303);
nor UO_1162 (O_1162,N_18426,N_17889);
nor UO_1163 (O_1163,N_19149,N_18958);
xnor UO_1164 (O_1164,N_16964,N_16513);
nor UO_1165 (O_1165,N_19870,N_17030);
and UO_1166 (O_1166,N_19997,N_18480);
and UO_1167 (O_1167,N_18024,N_18590);
or UO_1168 (O_1168,N_18535,N_19527);
nor UO_1169 (O_1169,N_16761,N_16372);
and UO_1170 (O_1170,N_16814,N_17281);
nor UO_1171 (O_1171,N_19949,N_16167);
nor UO_1172 (O_1172,N_17239,N_19094);
nand UO_1173 (O_1173,N_19290,N_16918);
nor UO_1174 (O_1174,N_16008,N_19655);
nand UO_1175 (O_1175,N_18977,N_19929);
nand UO_1176 (O_1176,N_19233,N_17086);
or UO_1177 (O_1177,N_18359,N_16697);
nor UO_1178 (O_1178,N_17067,N_16560);
nor UO_1179 (O_1179,N_18625,N_16796);
and UO_1180 (O_1180,N_18078,N_16801);
nor UO_1181 (O_1181,N_18412,N_17179);
and UO_1182 (O_1182,N_19868,N_16580);
and UO_1183 (O_1183,N_16645,N_16635);
nor UO_1184 (O_1184,N_17630,N_17590);
or UO_1185 (O_1185,N_18961,N_16839);
xnor UO_1186 (O_1186,N_19781,N_17904);
nand UO_1187 (O_1187,N_17230,N_19376);
and UO_1188 (O_1188,N_16775,N_16877);
nor UO_1189 (O_1189,N_17542,N_19214);
and UO_1190 (O_1190,N_18857,N_18848);
and UO_1191 (O_1191,N_19317,N_17158);
xor UO_1192 (O_1192,N_16009,N_16584);
and UO_1193 (O_1193,N_17222,N_16102);
nand UO_1194 (O_1194,N_18371,N_18041);
xor UO_1195 (O_1195,N_17918,N_16767);
nor UO_1196 (O_1196,N_18926,N_19202);
and UO_1197 (O_1197,N_16838,N_18293);
nand UO_1198 (O_1198,N_16011,N_17300);
and UO_1199 (O_1199,N_16470,N_18915);
or UO_1200 (O_1200,N_16351,N_19652);
and UO_1201 (O_1201,N_18671,N_16871);
and UO_1202 (O_1202,N_19247,N_17658);
nor UO_1203 (O_1203,N_16244,N_17191);
nor UO_1204 (O_1204,N_16686,N_17064);
and UO_1205 (O_1205,N_17055,N_16479);
nand UO_1206 (O_1206,N_17937,N_16662);
nor UO_1207 (O_1207,N_17360,N_17255);
nand UO_1208 (O_1208,N_18280,N_16503);
and UO_1209 (O_1209,N_18423,N_18511);
xnor UO_1210 (O_1210,N_17417,N_18164);
xnor UO_1211 (O_1211,N_18140,N_19663);
nor UO_1212 (O_1212,N_16085,N_17007);
nand UO_1213 (O_1213,N_17060,N_18589);
or UO_1214 (O_1214,N_19979,N_16357);
or UO_1215 (O_1215,N_17721,N_19379);
xor UO_1216 (O_1216,N_16599,N_17758);
nand UO_1217 (O_1217,N_16822,N_17315);
or UO_1218 (O_1218,N_17487,N_19387);
and UO_1219 (O_1219,N_16661,N_16861);
and UO_1220 (O_1220,N_16985,N_17908);
xor UO_1221 (O_1221,N_18180,N_18434);
nand UO_1222 (O_1222,N_16788,N_18405);
nand UO_1223 (O_1223,N_19930,N_16059);
or UO_1224 (O_1224,N_19478,N_19307);
nand UO_1225 (O_1225,N_17467,N_17164);
xnor UO_1226 (O_1226,N_16207,N_18106);
and UO_1227 (O_1227,N_17578,N_16533);
nor UO_1228 (O_1228,N_18471,N_17395);
or UO_1229 (O_1229,N_19812,N_16634);
or UO_1230 (O_1230,N_17174,N_19656);
nor UO_1231 (O_1231,N_16894,N_18200);
xnor UO_1232 (O_1232,N_19934,N_19699);
and UO_1233 (O_1233,N_19110,N_17126);
or UO_1234 (O_1234,N_19690,N_16483);
nand UO_1235 (O_1235,N_19873,N_18664);
nand UO_1236 (O_1236,N_19636,N_16202);
nor UO_1237 (O_1237,N_19987,N_16887);
nor UO_1238 (O_1238,N_16506,N_19833);
xnor UO_1239 (O_1239,N_16339,N_18149);
nand UO_1240 (O_1240,N_19389,N_17478);
nor UO_1241 (O_1241,N_16981,N_18001);
nor UO_1242 (O_1242,N_17705,N_17697);
nand UO_1243 (O_1243,N_16259,N_17722);
nand UO_1244 (O_1244,N_18198,N_19225);
or UO_1245 (O_1245,N_18801,N_16449);
and UO_1246 (O_1246,N_19487,N_17942);
and UO_1247 (O_1247,N_16791,N_19421);
nand UO_1248 (O_1248,N_19038,N_16301);
xnor UO_1249 (O_1249,N_18256,N_18343);
nand UO_1250 (O_1250,N_18766,N_16943);
nor UO_1251 (O_1251,N_18191,N_17768);
nand UO_1252 (O_1252,N_19685,N_16496);
nor UO_1253 (O_1253,N_18136,N_16655);
xor UO_1254 (O_1254,N_19988,N_16455);
or UO_1255 (O_1255,N_19398,N_18810);
xor UO_1256 (O_1256,N_17017,N_19463);
nand UO_1257 (O_1257,N_17083,N_16406);
xor UO_1258 (O_1258,N_18676,N_16797);
nor UO_1259 (O_1259,N_16178,N_18772);
xnor UO_1260 (O_1260,N_16384,N_17546);
xor UO_1261 (O_1261,N_16749,N_17132);
and UO_1262 (O_1262,N_19037,N_19270);
and UO_1263 (O_1263,N_16285,N_16227);
nand UO_1264 (O_1264,N_16953,N_17949);
and UO_1265 (O_1265,N_19065,N_19610);
xor UO_1266 (O_1266,N_19300,N_17443);
nand UO_1267 (O_1267,N_18326,N_16024);
and UO_1268 (O_1268,N_18691,N_16720);
or UO_1269 (O_1269,N_17744,N_16389);
nand UO_1270 (O_1270,N_18261,N_16833);
nor UO_1271 (O_1271,N_16851,N_19263);
or UO_1272 (O_1272,N_16653,N_18157);
xor UO_1273 (O_1273,N_16799,N_17124);
or UO_1274 (O_1274,N_17851,N_19702);
nor UO_1275 (O_1275,N_18758,N_18867);
nor UO_1276 (O_1276,N_18184,N_18466);
nor UO_1277 (O_1277,N_19932,N_17806);
or UO_1278 (O_1278,N_18790,N_17388);
nor UO_1279 (O_1279,N_19107,N_17848);
and UO_1280 (O_1280,N_18833,N_17469);
and UO_1281 (O_1281,N_16755,N_18424);
or UO_1282 (O_1282,N_17161,N_18500);
or UO_1283 (O_1283,N_18748,N_19185);
and UO_1284 (O_1284,N_19464,N_19657);
nand UO_1285 (O_1285,N_19249,N_19367);
nand UO_1286 (O_1286,N_19339,N_17427);
xor UO_1287 (O_1287,N_18182,N_16322);
nand UO_1288 (O_1288,N_17127,N_19386);
nand UO_1289 (O_1289,N_16508,N_19152);
nand UO_1290 (O_1290,N_17958,N_18925);
nor UO_1291 (O_1291,N_17288,N_16309);
nor UO_1292 (O_1292,N_17671,N_18791);
and UO_1293 (O_1293,N_19616,N_18601);
xor UO_1294 (O_1294,N_16193,N_17713);
nor UO_1295 (O_1295,N_18854,N_19280);
nor UO_1296 (O_1296,N_17808,N_19314);
nand UO_1297 (O_1297,N_18524,N_19672);
or UO_1298 (O_1298,N_16931,N_17025);
and UO_1299 (O_1299,N_18611,N_17277);
nand UO_1300 (O_1300,N_16671,N_18124);
or UO_1301 (O_1301,N_17377,N_16448);
nand UO_1302 (O_1302,N_17941,N_19635);
or UO_1303 (O_1303,N_19788,N_18703);
xor UO_1304 (O_1304,N_18531,N_16031);
nor UO_1305 (O_1305,N_17102,N_19937);
nor UO_1306 (O_1306,N_16342,N_19742);
and UO_1307 (O_1307,N_16245,N_18952);
or UO_1308 (O_1308,N_18337,N_18014);
xnor UO_1309 (O_1309,N_18885,N_16321);
and UO_1310 (O_1310,N_16030,N_16923);
nand UO_1311 (O_1311,N_19604,N_19831);
nor UO_1312 (O_1312,N_16532,N_19184);
and UO_1313 (O_1313,N_19811,N_17022);
nand UO_1314 (O_1314,N_19195,N_16199);
nor UO_1315 (O_1315,N_17167,N_19909);
or UO_1316 (O_1316,N_16837,N_17118);
xor UO_1317 (O_1317,N_19143,N_16410);
and UO_1318 (O_1318,N_16817,N_18460);
and UO_1319 (O_1319,N_17616,N_16474);
nand UO_1320 (O_1320,N_19760,N_16526);
xnor UO_1321 (O_1321,N_19215,N_18505);
nor UO_1322 (O_1322,N_17752,N_17662);
nand UO_1323 (O_1323,N_17683,N_19725);
xnor UO_1324 (O_1324,N_17534,N_18347);
nor UO_1325 (O_1325,N_19780,N_19580);
xnor UO_1326 (O_1326,N_18458,N_18685);
or UO_1327 (O_1327,N_17392,N_18626);
nand UO_1328 (O_1328,N_17262,N_19737);
nor UO_1329 (O_1329,N_18905,N_18255);
xnor UO_1330 (O_1330,N_18029,N_18882);
and UO_1331 (O_1331,N_18033,N_19559);
and UO_1332 (O_1332,N_19522,N_16329);
xor UO_1333 (O_1333,N_18167,N_19541);
or UO_1334 (O_1334,N_16995,N_17505);
or UO_1335 (O_1335,N_17946,N_19853);
nand UO_1336 (O_1336,N_18411,N_19459);
and UO_1337 (O_1337,N_16936,N_16161);
xnor UO_1338 (O_1338,N_19052,N_19560);
and UO_1339 (O_1339,N_18355,N_19589);
and UO_1340 (O_1340,N_18720,N_16769);
and UO_1341 (O_1341,N_16175,N_18472);
and UO_1342 (O_1342,N_19286,N_17886);
or UO_1343 (O_1343,N_17178,N_16166);
nor UO_1344 (O_1344,N_16704,N_18584);
and UO_1345 (O_1345,N_19731,N_17666);
or UO_1346 (O_1346,N_16915,N_17800);
nor UO_1347 (O_1347,N_16206,N_18941);
nor UO_1348 (O_1348,N_16400,N_19763);
xnor UO_1349 (O_1349,N_19188,N_17996);
xor UO_1350 (O_1350,N_17409,N_16614);
nand UO_1351 (O_1351,N_16868,N_17762);
nor UO_1352 (O_1352,N_19714,N_18972);
xor UO_1353 (O_1353,N_19508,N_17815);
or UO_1354 (O_1354,N_17984,N_16308);
and UO_1355 (O_1355,N_18060,N_16663);
or UO_1356 (O_1356,N_19625,N_16111);
or UO_1357 (O_1357,N_17153,N_18478);
or UO_1358 (O_1358,N_19854,N_16911);
nand UO_1359 (O_1359,N_16430,N_17020);
xnor UO_1360 (O_1360,N_19998,N_19902);
xnor UO_1361 (O_1361,N_18353,N_16119);
or UO_1362 (O_1362,N_16437,N_18406);
nor UO_1363 (O_1363,N_19312,N_18825);
nor UO_1364 (O_1364,N_16425,N_19667);
or UO_1365 (O_1365,N_17471,N_19627);
and UO_1366 (O_1366,N_19012,N_18400);
nor UO_1367 (O_1367,N_17235,N_17556);
and UO_1368 (O_1368,N_19304,N_16093);
and UO_1369 (O_1369,N_19328,N_18910);
nand UO_1370 (O_1370,N_17629,N_19586);
xor UO_1371 (O_1371,N_18641,N_17042);
xnor UO_1372 (O_1372,N_17301,N_16212);
nand UO_1373 (O_1373,N_16522,N_17343);
xnor UO_1374 (O_1374,N_16841,N_16312);
nor UO_1375 (O_1375,N_17416,N_18193);
nand UO_1376 (O_1376,N_16426,N_19348);
and UO_1377 (O_1377,N_16660,N_18245);
nor UO_1378 (O_1378,N_17479,N_16864);
nand UO_1379 (O_1379,N_16612,N_19309);
and UO_1380 (O_1380,N_17366,N_19964);
nand UO_1381 (O_1381,N_18217,N_19574);
nand UO_1382 (O_1382,N_16596,N_19542);
nand UO_1383 (O_1383,N_19495,N_18100);
and UO_1384 (O_1384,N_17887,N_19437);
nor UO_1385 (O_1385,N_18948,N_16988);
or UO_1386 (O_1386,N_19123,N_18823);
nand UO_1387 (O_1387,N_17466,N_19176);
and UO_1388 (O_1388,N_17352,N_16873);
and UO_1389 (O_1389,N_19474,N_16715);
nor UO_1390 (O_1390,N_17589,N_19528);
or UO_1391 (O_1391,N_18079,N_16204);
xnor UO_1392 (O_1392,N_18262,N_17038);
and UO_1393 (O_1393,N_17066,N_18431);
xor UO_1394 (O_1394,N_18290,N_17018);
and UO_1395 (O_1395,N_16126,N_18637);
or UO_1396 (O_1396,N_19827,N_19817);
or UO_1397 (O_1397,N_16717,N_17454);
or UO_1398 (O_1398,N_17876,N_19570);
or UO_1399 (O_1399,N_18205,N_18404);
and UO_1400 (O_1400,N_16393,N_18545);
nor UO_1401 (O_1401,N_16097,N_18981);
nor UO_1402 (O_1402,N_17382,N_18349);
nand UO_1403 (O_1403,N_16926,N_16287);
and UO_1404 (O_1404,N_16992,N_18647);
or UO_1405 (O_1405,N_17477,N_16418);
and UO_1406 (O_1406,N_16957,N_19517);
nor UO_1407 (O_1407,N_17203,N_18681);
xor UO_1408 (O_1408,N_17934,N_17968);
nor UO_1409 (O_1409,N_18567,N_18271);
xnor UO_1410 (O_1410,N_16856,N_16889);
or UO_1411 (O_1411,N_16272,N_18842);
nand UO_1412 (O_1412,N_17798,N_17008);
nand UO_1413 (O_1413,N_16466,N_19768);
and UO_1414 (O_1414,N_18985,N_19068);
nor UO_1415 (O_1415,N_19088,N_16884);
xnor UO_1416 (O_1416,N_18933,N_19201);
or UO_1417 (O_1417,N_19860,N_18273);
xor UO_1418 (O_1418,N_18419,N_16932);
nand UO_1419 (O_1419,N_16753,N_16284);
nor UO_1420 (O_1420,N_16275,N_18877);
xnor UO_1421 (O_1421,N_16852,N_16475);
or UO_1422 (O_1422,N_17000,N_17792);
xnor UO_1423 (O_1423,N_18216,N_17080);
and UO_1424 (O_1424,N_17483,N_19553);
or UO_1425 (O_1425,N_16639,N_18158);
nor UO_1426 (O_1426,N_16751,N_18888);
xnor UO_1427 (O_1427,N_16417,N_19887);
and UO_1428 (O_1428,N_18470,N_18759);
nand UO_1429 (O_1429,N_19954,N_19691);
xor UO_1430 (O_1430,N_18732,N_17930);
and UO_1431 (O_1431,N_18988,N_19950);
xor UO_1432 (O_1432,N_17231,N_17867);
nor UO_1433 (O_1433,N_18710,N_16363);
nor UO_1434 (O_1434,N_16016,N_19985);
nor UO_1435 (O_1435,N_17939,N_17708);
or UO_1436 (O_1436,N_17584,N_17279);
or UO_1437 (O_1437,N_17336,N_18089);
or UO_1438 (O_1438,N_16014,N_17079);
and UO_1439 (O_1439,N_17070,N_16062);
nand UO_1440 (O_1440,N_19446,N_16124);
nor UO_1441 (O_1441,N_17321,N_17966);
xnor UO_1442 (O_1442,N_19236,N_16305);
and UO_1443 (O_1443,N_16125,N_19411);
and UO_1444 (O_1444,N_18763,N_17873);
xnor UO_1445 (O_1445,N_19785,N_18474);
nand UO_1446 (O_1446,N_19590,N_17229);
nor UO_1447 (O_1447,N_18795,N_19066);
xnor UO_1448 (O_1448,N_17668,N_16613);
and UO_1449 (O_1449,N_16813,N_16909);
xnor UO_1450 (O_1450,N_19080,N_17977);
or UO_1451 (O_1451,N_19569,N_17892);
nor UO_1452 (O_1452,N_16048,N_18197);
xor UO_1453 (O_1453,N_19000,N_18513);
xor UO_1454 (O_1454,N_18581,N_16281);
nand UO_1455 (O_1455,N_19218,N_16594);
nand UO_1456 (O_1456,N_16746,N_16601);
nand UO_1457 (O_1457,N_19010,N_19429);
nand UO_1458 (O_1458,N_19030,N_16563);
or UO_1459 (O_1459,N_17309,N_16381);
nor UO_1460 (O_1460,N_16379,N_16180);
and UO_1461 (O_1461,N_16441,N_16327);
nand UO_1462 (O_1462,N_18364,N_17962);
nand UO_1463 (O_1463,N_16544,N_16355);
xnor UO_1464 (O_1464,N_18490,N_19305);
nand UO_1465 (O_1465,N_17603,N_18920);
and UO_1466 (O_1466,N_19343,N_18268);
or UO_1467 (O_1467,N_17056,N_16853);
nor UO_1468 (O_1468,N_18382,N_16969);
xor UO_1469 (O_1469,N_18304,N_18510);
and UO_1470 (O_1470,N_16935,N_19957);
nand UO_1471 (O_1471,N_18308,N_19668);
xor UO_1472 (O_1472,N_17447,N_17320);
nand UO_1473 (O_1473,N_17185,N_19855);
or UO_1474 (O_1474,N_17232,N_16770);
xnor UO_1475 (O_1475,N_16574,N_17407);
nor UO_1476 (O_1476,N_18108,N_18921);
and UO_1477 (O_1477,N_16826,N_18097);
nor UO_1478 (O_1478,N_17293,N_19962);
and UO_1479 (O_1479,N_19804,N_18644);
xor UO_1480 (O_1480,N_18450,N_16254);
and UO_1481 (O_1481,N_19033,N_17652);
nand UO_1482 (O_1482,N_17869,N_16404);
xnor UO_1483 (O_1483,N_18826,N_19660);
nor UO_1484 (O_1484,N_19715,N_17155);
xor UO_1485 (O_1485,N_19775,N_17775);
nand UO_1486 (O_1486,N_18420,N_17516);
nand UO_1487 (O_1487,N_19344,N_16350);
nor UO_1488 (O_1488,N_17960,N_19073);
xnor UO_1489 (O_1489,N_18632,N_18668);
or UO_1490 (O_1490,N_18990,N_19399);
xnor UO_1491 (O_1491,N_16482,N_18231);
and UO_1492 (O_1492,N_19748,N_16745);
nand UO_1493 (O_1493,N_16340,N_16414);
nor UO_1494 (O_1494,N_18436,N_16832);
nand UO_1495 (O_1495,N_17877,N_17950);
or UO_1496 (O_1496,N_16054,N_17163);
nor UO_1497 (O_1497,N_19473,N_17755);
nand UO_1498 (O_1498,N_19055,N_19320);
and UO_1499 (O_1499,N_19479,N_16863);
nor UO_1500 (O_1500,N_16253,N_18085);
nor UO_1501 (O_1501,N_17256,N_16529);
nand UO_1502 (O_1502,N_17757,N_17702);
xor UO_1503 (O_1503,N_19408,N_19806);
nor UO_1504 (O_1504,N_17134,N_16172);
nand UO_1505 (O_1505,N_18916,N_19961);
nand UO_1506 (O_1506,N_19069,N_18192);
nor UO_1507 (O_1507,N_16607,N_19315);
nor UO_1508 (O_1508,N_17268,N_18604);
and UO_1509 (O_1509,N_17582,N_17788);
nand UO_1510 (O_1510,N_19978,N_19409);
xnor UO_1511 (O_1511,N_17057,N_18113);
or UO_1512 (O_1512,N_19850,N_16130);
nand UO_1513 (O_1513,N_19213,N_18903);
or UO_1514 (O_1514,N_17732,N_19192);
and UO_1515 (O_1515,N_17490,N_18844);
nor UO_1516 (O_1516,N_18093,N_17763);
and UO_1517 (O_1517,N_19014,N_18174);
xor UO_1518 (O_1518,N_19134,N_19899);
and UO_1519 (O_1519,N_19989,N_16518);
nor UO_1520 (O_1520,N_18827,N_16302);
and UO_1521 (O_1521,N_17923,N_19920);
or UO_1522 (O_1522,N_17379,N_17921);
or UO_1523 (O_1523,N_19089,N_17704);
or UO_1524 (O_1524,N_18799,N_18062);
xor UO_1525 (O_1525,N_19013,N_16182);
or UO_1526 (O_1526,N_19632,N_17223);
xor UO_1527 (O_1527,N_18160,N_16505);
nand UO_1528 (O_1528,N_19113,N_16432);
nand UO_1529 (O_1529,N_19897,N_19673);
nand UO_1530 (O_1530,N_19881,N_16306);
or UO_1531 (O_1531,N_19384,N_16187);
xor UO_1532 (O_1532,N_19721,N_18315);
nand UO_1533 (O_1533,N_17310,N_18559);
nor UO_1534 (O_1534,N_18740,N_17521);
or UO_1535 (O_1535,N_17759,N_19151);
nor UO_1536 (O_1536,N_18469,N_16878);
and UO_1537 (O_1537,N_16665,N_17838);
and UO_1538 (O_1538,N_17660,N_18312);
nor UO_1539 (O_1539,N_19518,N_16537);
nand UO_1540 (O_1540,N_17274,N_19470);
and UO_1541 (O_1541,N_16829,N_16488);
and UO_1542 (O_1542,N_19034,N_16158);
xor UO_1543 (O_1543,N_17121,N_16919);
nor UO_1544 (O_1544,N_16067,N_17829);
or UO_1545 (O_1545,N_18686,N_19039);
nand UO_1546 (O_1546,N_19622,N_19335);
or UO_1547 (O_1547,N_17087,N_16320);
nor UO_1548 (O_1548,N_16231,N_18677);
or UO_1549 (O_1549,N_19075,N_17186);
or UO_1550 (O_1550,N_19164,N_19986);
nand UO_1551 (O_1551,N_16391,N_17679);
and UO_1552 (O_1552,N_16718,N_18228);
nor UO_1553 (O_1553,N_18484,N_16657);
nor UO_1554 (O_1554,N_17494,N_18912);
nor UO_1555 (O_1555,N_16581,N_16937);
nand UO_1556 (O_1556,N_18051,N_17216);
or UO_1557 (O_1557,N_16461,N_16546);
and UO_1558 (O_1558,N_18757,N_16042);
or UO_1559 (O_1559,N_16593,N_19889);
and UO_1560 (O_1560,N_19417,N_18185);
or UO_1561 (O_1561,N_19354,N_18342);
and UO_1562 (O_1562,N_18227,N_18967);
nor UO_1563 (O_1563,N_16623,N_19600);
xor UO_1564 (O_1564,N_17972,N_18652);
or UO_1565 (O_1565,N_17917,N_16163);
or UO_1566 (O_1566,N_19534,N_19438);
or UO_1567 (O_1567,N_19078,N_17694);
or UO_1568 (O_1568,N_16402,N_19053);
nor UO_1569 (O_1569,N_16673,N_18397);
or UO_1570 (O_1570,N_17481,N_16232);
and UO_1571 (O_1571,N_17142,N_17499);
xnor UO_1572 (O_1572,N_16685,N_17135);
nor UO_1573 (O_1573,N_18969,N_16290);
xor UO_1574 (O_1574,N_19441,N_18147);
or UO_1575 (O_1575,N_18679,N_19651);
and UO_1576 (O_1576,N_16978,N_19019);
nand UO_1577 (O_1577,N_19318,N_16520);
and UO_1578 (O_1578,N_18666,N_18930);
xnor UO_1579 (O_1579,N_16869,N_18630);
xnor UO_1580 (O_1580,N_18465,N_17391);
and UO_1581 (O_1581,N_16744,N_17997);
nand UO_1582 (O_1582,N_19778,N_19345);
or UO_1583 (O_1583,N_17455,N_19281);
or UO_1584 (O_1584,N_16648,N_19942);
nand UO_1585 (O_1585,N_17200,N_18561);
xnor UO_1586 (O_1586,N_18557,N_19838);
nand UO_1587 (O_1587,N_19461,N_16143);
and UO_1588 (O_1588,N_17506,N_17330);
nand UO_1589 (O_1589,N_16604,N_18575);
and UO_1590 (O_1590,N_19340,N_18240);
nor UO_1591 (O_1591,N_17302,N_18853);
and UO_1592 (O_1592,N_17422,N_19258);
or UO_1593 (O_1593,N_17495,N_18208);
xnor UO_1594 (O_1594,N_19095,N_16407);
nor UO_1595 (O_1595,N_19439,N_18086);
xor UO_1596 (O_1596,N_17441,N_19759);
xnor UO_1597 (O_1597,N_16403,N_18171);
xor UO_1598 (O_1598,N_19336,N_16422);
xor UO_1599 (O_1599,N_17741,N_17371);
nand UO_1600 (O_1600,N_19189,N_19591);
nand UO_1601 (O_1601,N_19981,N_17376);
xnor UO_1602 (O_1602,N_19883,N_17592);
and UO_1603 (O_1603,N_18142,N_17394);
nand UO_1604 (O_1604,N_19064,N_18275);
nor UO_1605 (O_1605,N_18587,N_17935);
xnor UO_1606 (O_1606,N_16730,N_17130);
xnor UO_1607 (O_1607,N_19952,N_17748);
and UO_1608 (O_1608,N_19370,N_17009);
xnor UO_1609 (O_1609,N_19606,N_18418);
nand UO_1610 (O_1610,N_19082,N_19970);
xnor UO_1611 (O_1611,N_17893,N_19901);
nor UO_1612 (O_1612,N_19990,N_17948);
nand UO_1613 (O_1613,N_17706,N_18804);
nand UO_1614 (O_1614,N_17502,N_17685);
and UO_1615 (O_1615,N_19585,N_18776);
xor UO_1616 (O_1616,N_17369,N_16252);
nor UO_1617 (O_1617,N_17485,N_19537);
xnor UO_1618 (O_1618,N_19931,N_18504);
nor UO_1619 (O_1619,N_16311,N_17965);
nand UO_1620 (O_1620,N_17436,N_16942);
xnor UO_1621 (O_1621,N_18949,N_17859);
nand UO_1622 (O_1622,N_17446,N_19890);
nor UO_1623 (O_1623,N_19480,N_17559);
and UO_1624 (O_1624,N_16773,N_18578);
nor UO_1625 (O_1625,N_17034,N_18537);
and UO_1626 (O_1626,N_19396,N_16276);
xor UO_1627 (O_1627,N_17385,N_18211);
nand UO_1628 (O_1628,N_16553,N_16419);
xor UO_1629 (O_1629,N_18264,N_18314);
or UO_1630 (O_1630,N_17845,N_19175);
and UO_1631 (O_1631,N_17289,N_19102);
xnor UO_1632 (O_1632,N_17449,N_16454);
nor UO_1633 (O_1633,N_19445,N_19571);
nand UO_1634 (O_1634,N_17325,N_17368);
xnor UO_1635 (O_1635,N_18230,N_18667);
nor UO_1636 (O_1636,N_19365,N_18901);
nand UO_1637 (O_1637,N_19430,N_16148);
xor UO_1638 (O_1638,N_16637,N_18021);
xnor UO_1639 (O_1639,N_19041,N_18993);
or UO_1640 (O_1640,N_17036,N_18038);
and UO_1641 (O_1641,N_19876,N_17634);
and UO_1642 (O_1642,N_16096,N_18229);
xor UO_1643 (O_1643,N_18082,N_19765);
and UO_1644 (O_1644,N_19900,N_18709);
and UO_1645 (O_1645,N_16264,N_16521);
xor UO_1646 (O_1646,N_19015,N_16258);
or UO_1647 (O_1647,N_18429,N_16611);
nand UO_1648 (O_1648,N_18162,N_19845);
nor UO_1649 (O_1649,N_16356,N_16433);
xor UO_1650 (O_1650,N_18852,N_19338);
and UO_1651 (O_1651,N_16246,N_16830);
nand UO_1652 (O_1652,N_18169,N_19090);
nor UO_1653 (O_1653,N_16205,N_19006);
xnor UO_1654 (O_1654,N_19526,N_17225);
nor UO_1655 (O_1655,N_19808,N_19689);
nor UO_1656 (O_1656,N_19498,N_17076);
nand UO_1657 (O_1657,N_19007,N_18223);
nor UO_1658 (O_1658,N_16405,N_18351);
nand UO_1659 (O_1659,N_17146,N_19822);
xnor UO_1660 (O_1660,N_19383,N_19244);
nor UO_1661 (O_1661,N_19701,N_18553);
xnor UO_1662 (O_1662,N_17899,N_17632);
xor UO_1663 (O_1663,N_16289,N_17597);
or UO_1664 (O_1664,N_18617,N_18087);
and UO_1665 (O_1665,N_18246,N_17195);
nand UO_1666 (O_1666,N_18145,N_19238);
or UO_1667 (O_1667,N_17626,N_17863);
xor UO_1668 (O_1668,N_17314,N_18623);
and UO_1669 (O_1669,N_17617,N_17544);
nor UO_1670 (O_1670,N_19681,N_17334);
or UO_1671 (O_1671,N_19739,N_18722);
xnor UO_1672 (O_1672,N_17140,N_16465);
and UO_1673 (O_1673,N_18923,N_16359);
nand UO_1674 (O_1674,N_17614,N_17785);
xor UO_1675 (O_1675,N_18953,N_19278);
xor UO_1676 (O_1676,N_17654,N_19846);
and UO_1677 (O_1677,N_16053,N_19373);
xor UO_1678 (O_1678,N_18324,N_17903);
nand UO_1679 (O_1679,N_18428,N_17780);
and UO_1680 (O_1680,N_16401,N_18814);
xnor UO_1681 (O_1681,N_18328,N_19047);
and UO_1682 (O_1682,N_19965,N_19404);
and UO_1683 (O_1683,N_18964,N_16499);
or UO_1684 (O_1684,N_17649,N_17208);
nor UO_1685 (O_1685,N_16605,N_16089);
xor UO_1686 (O_1686,N_16764,N_19872);
xor UO_1687 (O_1687,N_16855,N_18375);
nor UO_1688 (O_1688,N_17270,N_19025);
and UO_1689 (O_1689,N_16223,N_17192);
nand UO_1690 (O_1690,N_16478,N_18391);
nor UO_1691 (O_1691,N_18095,N_18821);
nand UO_1692 (O_1692,N_17037,N_17766);
nor UO_1693 (O_1693,N_16472,N_17602);
nand UO_1694 (O_1694,N_19193,N_16831);
xnor UO_1695 (O_1695,N_18970,N_16458);
nand UO_1696 (O_1696,N_18507,N_16587);
nor UO_1697 (O_1697,N_16421,N_17895);
and UO_1698 (O_1698,N_17286,N_17193);
or UO_1699 (O_1699,N_18998,N_17012);
xnor UO_1700 (O_1700,N_18103,N_18030);
nor UO_1701 (O_1701,N_16726,N_16977);
nand UO_1702 (O_1702,N_16487,N_17669);
nand UO_1703 (O_1703,N_19770,N_16610);
nor UO_1704 (O_1704,N_16453,N_18091);
and UO_1705 (O_1705,N_16819,N_18675);
nand UO_1706 (O_1706,N_17822,N_17484);
and UO_1707 (O_1707,N_18284,N_18570);
and UO_1708 (O_1708,N_16328,N_16575);
or UO_1709 (O_1709,N_16930,N_19198);
nor UO_1710 (O_1710,N_17672,N_19104);
and UO_1711 (O_1711,N_16577,N_19628);
nor UO_1712 (O_1712,N_19894,N_18365);
nand UO_1713 (O_1713,N_19524,N_18794);
or UO_1714 (O_1714,N_18708,N_17901);
nor UO_1715 (O_1715,N_16950,N_17445);
nor UO_1716 (O_1716,N_17421,N_16140);
xor UO_1717 (O_1717,N_16438,N_16765);
xor UO_1718 (O_1718,N_18292,N_16710);
nand UO_1719 (O_1719,N_18951,N_18742);
xnor UO_1720 (O_1720,N_16790,N_19939);
nor UO_1721 (O_1721,N_17885,N_18806);
xnor UO_1722 (O_1722,N_18690,N_16651);
nand UO_1723 (O_1723,N_19219,N_18358);
nand UO_1724 (O_1724,N_18340,N_19615);
nand UO_1725 (O_1725,N_18741,N_16792);
or UO_1726 (O_1726,N_17719,N_16840);
nand UO_1727 (O_1727,N_18800,N_19642);
nand UO_1728 (O_1728,N_18815,N_18730);
nor UO_1729 (O_1729,N_18512,N_17880);
or UO_1730 (O_1730,N_16716,N_16951);
nor UO_1731 (O_1731,N_18321,N_17964);
nor UO_1732 (O_1732,N_18084,N_16809);
xnor UO_1733 (O_1733,N_17574,N_17508);
nand UO_1734 (O_1734,N_17884,N_19210);
xor UO_1735 (O_1735,N_16914,N_16238);
and UO_1736 (O_1736,N_18195,N_18980);
or UO_1737 (O_1737,N_17082,N_17988);
xnor UO_1738 (O_1738,N_19362,N_18523);
xor UO_1739 (O_1739,N_19097,N_17316);
nand UO_1740 (O_1740,N_18899,N_18447);
and UO_1741 (O_1741,N_19168,N_18363);
and UO_1742 (O_1742,N_16768,N_17995);
nor UO_1743 (O_1743,N_19081,N_19704);
nor UO_1744 (O_1744,N_19226,N_17906);
nor UO_1745 (O_1745,N_19230,N_16198);
nor UO_1746 (O_1746,N_17331,N_16041);
or UO_1747 (O_1747,N_19764,N_16510);
nand UO_1748 (O_1748,N_19156,N_18897);
or UO_1749 (O_1749,N_17898,N_18856);
or UO_1750 (O_1750,N_16122,N_18383);
or UO_1751 (O_1751,N_19921,N_18403);
xnor UO_1752 (O_1752,N_17291,N_17957);
and UO_1753 (O_1753,N_16777,N_17684);
nor UO_1754 (O_1754,N_19415,N_16684);
and UO_1755 (O_1755,N_19276,N_17040);
nand UO_1756 (O_1756,N_18592,N_19465);
nand UO_1757 (O_1757,N_16975,N_16023);
or UO_1758 (O_1758,N_16993,N_17517);
nand UO_1759 (O_1759,N_19960,N_17723);
nand UO_1760 (O_1760,N_19380,N_18187);
or UO_1761 (O_1761,N_16917,N_16542);
xor UO_1762 (O_1762,N_19918,N_19923);
nand UO_1763 (O_1763,N_17688,N_16495);
and UO_1764 (O_1764,N_16170,N_18055);
or UO_1765 (O_1765,N_18607,N_19363);
and UO_1766 (O_1766,N_16709,N_18105);
nand UO_1767 (O_1767,N_19114,N_18764);
xnor UO_1768 (O_1768,N_17509,N_19142);
or UO_1769 (O_1769,N_16469,N_16055);
or UO_1770 (O_1770,N_19087,N_17664);
and UO_1771 (O_1771,N_17969,N_19755);
xnor UO_1772 (O_1772,N_19815,N_18744);
or UO_1773 (O_1773,N_16149,N_17305);
xnor UO_1774 (O_1774,N_18285,N_19837);
nor UO_1775 (O_1775,N_17733,N_19575);
xor UO_1776 (O_1776,N_18032,N_16762);
xor UO_1777 (O_1777,N_18947,N_16583);
or UO_1778 (O_1778,N_18118,N_16703);
xor UO_1779 (O_1779,N_18112,N_18387);
nor UO_1780 (O_1780,N_16020,N_18126);
nand UO_1781 (O_1781,N_17902,N_17189);
xnor UO_1782 (O_1782,N_16867,N_17745);
nor UO_1783 (O_1783,N_18251,N_18442);
nor UO_1784 (O_1784,N_18706,N_17116);
nand UO_1785 (O_1785,N_16256,N_16549);
or UO_1786 (O_1786,N_18301,N_16387);
and UO_1787 (O_1787,N_17843,N_19133);
nand UO_1788 (O_1788,N_16625,N_16550);
xor UO_1789 (O_1789,N_18481,N_18783);
xnor UO_1790 (O_1790,N_18627,N_18224);
nor UO_1791 (O_1791,N_16999,N_17861);
xnor UO_1792 (O_1792,N_18309,N_16442);
and UO_1793 (O_1793,N_18286,N_19766);
nor UO_1794 (O_1794,N_16824,N_19607);
nand UO_1795 (O_1795,N_16145,N_17555);
or UO_1796 (O_1796,N_17141,N_18782);
and UO_1797 (O_1797,N_18701,N_18333);
xor UO_1798 (O_1798,N_17746,N_19638);
nand UO_1799 (O_1799,N_19497,N_17803);
nand UO_1800 (O_1800,N_19150,N_17810);
nor UO_1801 (O_1801,N_18121,N_17156);
or UO_1802 (O_1802,N_18573,N_19333);
or UO_1803 (O_1803,N_17657,N_19592);
xor UO_1804 (O_1804,N_18025,N_16672);
or UO_1805 (O_1805,N_16958,N_17094);
xnor UO_1806 (O_1806,N_18010,N_19820);
or UO_1807 (O_1807,N_17348,N_16017);
and UO_1808 (O_1808,N_19166,N_17594);
nand UO_1809 (O_1809,N_18571,N_19980);
nor UO_1810 (O_1810,N_17249,N_17870);
nand UO_1811 (O_1811,N_17686,N_16225);
xnor UO_1812 (O_1812,N_18840,N_16626);
and UO_1813 (O_1813,N_17465,N_17989);
and UO_1814 (O_1814,N_17206,N_19933);
nand UO_1815 (O_1815,N_17345,N_17287);
xnor UO_1816 (O_1816,N_17292,N_19131);
nor UO_1817 (O_1817,N_17781,N_18341);
xor UO_1818 (O_1818,N_17133,N_16695);
xnor UO_1819 (O_1819,N_18995,N_16732);
or UO_1820 (O_1820,N_19420,N_17665);
nor UO_1821 (O_1821,N_17245,N_18672);
nor UO_1822 (O_1822,N_18908,N_19319);
nand UO_1823 (O_1823,N_18141,N_18194);
or UO_1824 (O_1824,N_19787,N_19154);
and UO_1825 (O_1825,N_17338,N_16586);
nand UO_1826 (O_1826,N_17462,N_18643);
or UO_1827 (O_1827,N_19251,N_17980);
and UO_1828 (O_1828,N_19267,N_18134);
xor UO_1829 (O_1829,N_17793,N_19711);
or UO_1830 (O_1830,N_17551,N_16925);
or UO_1831 (O_1831,N_17276,N_16434);
and UO_1832 (O_1832,N_16854,N_18173);
xnor UO_1833 (O_1833,N_17595,N_17151);
xnor UO_1834 (O_1834,N_19581,N_16152);
and UO_1835 (O_1835,N_19848,N_17157);
nand UO_1836 (O_1836,N_19753,N_17627);
or UO_1837 (O_1837,N_19492,N_17978);
and UO_1838 (O_1838,N_19839,N_19967);
nand UO_1839 (O_1839,N_18163,N_19076);
xor UO_1840 (O_1840,N_17656,N_19944);
or UO_1841 (O_1841,N_16961,N_18244);
nor UO_1842 (O_1842,N_17974,N_16034);
or UO_1843 (O_1843,N_19631,N_19024);
nand UO_1844 (O_1844,N_18893,N_17760);
or UO_1845 (O_1845,N_19896,N_18919);
nor UO_1846 (O_1846,N_17635,N_19099);
or UO_1847 (O_1847,N_16243,N_16369);
and UO_1848 (O_1848,N_16451,N_19709);
nor UO_1849 (O_1849,N_19072,N_16003);
xor UO_1850 (O_1850,N_18468,N_19729);
and UO_1851 (O_1851,N_17199,N_19120);
or UO_1852 (O_1852,N_17175,N_17698);
and UO_1853 (O_1853,N_19996,N_16039);
and UO_1854 (O_1854,N_17528,N_16046);
or UO_1855 (O_1855,N_17248,N_19644);
xor UO_1856 (O_1856,N_19049,N_18956);
or UO_1857 (O_1857,N_18688,N_18316);
nor UO_1858 (O_1858,N_18181,N_19605);
and UO_1859 (O_1859,N_19141,N_19767);
and UO_1860 (O_1860,N_17828,N_16781);
or UO_1861 (O_1861,N_17143,N_17790);
and UO_1862 (O_1862,N_19448,N_16038);
nor UO_1863 (O_1863,N_16345,N_18131);
nor UO_1864 (O_1864,N_18152,N_18684);
nand UO_1865 (O_1865,N_18962,N_17123);
nor UO_1866 (O_1866,N_19686,N_19283);
xnor UO_1867 (O_1867,N_18457,N_16195);
nor UO_1868 (O_1868,N_17524,N_19245);
nand UO_1869 (O_1869,N_18818,N_16928);
nand UO_1870 (O_1870,N_17735,N_18061);
nand UO_1871 (O_1871,N_18247,N_17375);
xnor UO_1872 (O_1872,N_16669,N_18026);
nor UO_1873 (O_1873,N_16260,N_18994);
nor UO_1874 (O_1874,N_19703,N_17304);
or UO_1875 (O_1875,N_16157,N_16823);
and UO_1876 (O_1876,N_17774,N_18959);
or UO_1877 (O_1877,N_18473,N_19291);
xnor UO_1878 (O_1878,N_16719,N_16219);
nor UO_1879 (O_1879,N_19925,N_19562);
nor UO_1880 (O_1880,N_17244,N_16336);
nor UO_1881 (O_1881,N_19917,N_17639);
or UO_1882 (O_1882,N_18390,N_17093);
and UO_1883 (O_1883,N_16315,N_17794);
and UO_1884 (O_1884,N_16304,N_18047);
nand UO_1885 (O_1885,N_17428,N_18421);
and UO_1886 (O_1886,N_17003,N_19269);
xnor UO_1887 (O_1887,N_17162,N_17786);
nand UO_1888 (O_1888,N_18680,N_19795);
nor UO_1889 (O_1889,N_16107,N_19682);
nor UO_1890 (O_1890,N_18654,N_17833);
nand UO_1891 (O_1891,N_18566,N_16996);
or UO_1892 (O_1892,N_17970,N_17470);
nand UO_1893 (O_1893,N_16078,N_16082);
nor UO_1894 (O_1894,N_16836,N_18749);
and UO_1895 (O_1895,N_17378,N_18957);
nand UO_1896 (O_1896,N_18579,N_19864);
xnor UO_1897 (O_1897,N_17129,N_18236);
nand UO_1898 (O_1898,N_16638,N_19060);
nor UO_1899 (O_1899,N_17220,N_18099);
and UO_1900 (O_1900,N_16314,N_18756);
nor UO_1901 (O_1901,N_18296,N_16647);
nand UO_1902 (O_1902,N_19468,N_16866);
or UO_1903 (O_1903,N_18624,N_19697);
xnor UO_1904 (O_1904,N_17924,N_17896);
nor UO_1905 (O_1905,N_18374,N_18533);
xor UO_1906 (O_1906,N_19744,N_17019);
or UO_1907 (O_1907,N_16787,N_19958);
xor UO_1908 (O_1908,N_18007,N_19941);
nor UO_1909 (O_1909,N_19687,N_19993);
and UO_1910 (O_1910,N_16318,N_17107);
or UO_1911 (O_1911,N_19447,N_18747);
or UO_1912 (O_1912,N_18863,N_16743);
nor UO_1913 (O_1913,N_16780,N_17791);
nor UO_1914 (O_1914,N_19294,N_16847);
xor UO_1915 (O_1915,N_17273,N_18816);
or UO_1916 (O_1916,N_19326,N_18661);
or UO_1917 (O_1917,N_19132,N_16233);
nor UO_1918 (O_1918,N_17673,N_19629);
and UO_1919 (O_1919,N_19722,N_16010);
xnor UO_1920 (O_1920,N_16681,N_18077);
and UO_1921 (O_1921,N_16783,N_16912);
and UO_1922 (O_1922,N_18274,N_18323);
xor UO_1923 (O_1923,N_19346,N_16299);
nand UO_1924 (O_1924,N_16667,N_17404);
xor UO_1925 (O_1925,N_16548,N_18509);
nor UO_1926 (O_1926,N_17280,N_17650);
or UO_1927 (O_1927,N_17444,N_17807);
and UO_1928 (O_1928,N_16578,N_17104);
xnor UO_1929 (O_1929,N_17117,N_16035);
and UO_1930 (O_1930,N_18016,N_17246);
xor UO_1931 (O_1931,N_18310,N_16413);
xnor UO_1932 (O_1932,N_16471,N_19374);
xor UO_1933 (O_1933,N_18401,N_18832);
and UO_1934 (O_1934,N_17579,N_18348);
nand UO_1935 (O_1935,N_18657,N_18767);
nor UO_1936 (O_1936,N_18770,N_16262);
xor UO_1937 (O_1937,N_17282,N_16310);
nor UO_1938 (O_1938,N_19093,N_16095);
or UO_1939 (O_1939,N_17173,N_19496);
nand UO_1940 (O_1940,N_16319,N_17503);
nand UO_1941 (O_1941,N_17824,N_17513);
nor UO_1942 (O_1942,N_19557,N_17333);
or UO_1943 (O_1943,N_17847,N_18373);
and UO_1944 (O_1944,N_19807,N_18050);
nand UO_1945 (O_1945,N_19009,N_18488);
nor UO_1946 (O_1946,N_16347,N_19393);
nand UO_1947 (O_1947,N_18354,N_19692);
nor UO_1948 (O_1948,N_16420,N_16630);
nor UO_1949 (O_1949,N_18257,N_16997);
xnor UO_1950 (O_1950,N_19710,N_16875);
nor UO_1951 (O_1951,N_19914,N_19180);
or UO_1952 (O_1952,N_18467,N_19299);
xnor UO_1953 (O_1953,N_16040,N_17622);
or UO_1954 (O_1954,N_18219,N_19696);
nand UO_1955 (O_1955,N_16087,N_19599);
nand UO_1956 (O_1956,N_18209,N_18433);
nor UO_1957 (O_1957,N_18125,N_17150);
or UO_1958 (O_1958,N_18278,N_17109);
nor UO_1959 (O_1959,N_18798,N_18817);
xor UO_1960 (O_1960,N_17448,N_17640);
nand UO_1961 (O_1961,N_19613,N_16463);
xor UO_1962 (O_1962,N_16397,N_19486);
or UO_1963 (O_1963,N_19805,N_19400);
or UO_1964 (O_1964,N_16467,N_19135);
and UO_1965 (O_1965,N_16173,N_19995);
and UO_1966 (O_1966,N_18408,N_16976);
xnor UO_1967 (O_1967,N_16714,N_18935);
xnor UO_1968 (O_1968,N_19948,N_17796);
or UO_1969 (O_1969,N_18073,N_19070);
and UO_1970 (O_1970,N_17805,N_18673);
or UO_1971 (O_1971,N_18177,N_16750);
nor UO_1972 (O_1972,N_16805,N_17585);
nand UO_1973 (O_1973,N_17739,N_16303);
nand UO_1974 (O_1974,N_18502,N_16113);
and UO_1975 (O_1975,N_19747,N_16617);
or UO_1976 (O_1976,N_18004,N_19633);
nor UO_1977 (O_1977,N_19277,N_17999);
xnor UO_1978 (O_1978,N_17437,N_18911);
nand UO_1979 (O_1979,N_17403,N_17139);
nor UO_1980 (O_1980,N_18600,N_17113);
and UO_1981 (O_1981,N_16541,N_18698);
xnor UO_1982 (O_1982,N_17858,N_19098);
xor UO_1983 (O_1983,N_16176,N_17636);
or UO_1984 (O_1984,N_19844,N_19893);
and UO_1985 (O_1985,N_17468,N_18233);
or UO_1986 (O_1986,N_18735,N_19324);
xor UO_1987 (O_1987,N_16239,N_18536);
and UO_1988 (O_1988,N_19457,N_16535);
nor UO_1989 (O_1989,N_16200,N_16712);
nand UO_1990 (O_1990,N_17567,N_17050);
nand UO_1991 (O_1991,N_17090,N_16247);
and UO_1992 (O_1992,N_19727,N_16724);
nor UO_1993 (O_1993,N_17351,N_19450);
or UO_1994 (O_1994,N_16155,N_19608);
nor UO_1995 (O_1995,N_17439,N_17312);
nand UO_1996 (O_1996,N_18725,N_19502);
or UO_1997 (O_1997,N_16725,N_18499);
nor UO_1998 (O_1998,N_18441,N_17299);
or UO_1999 (O_1999,N_19824,N_17522);
or UO_2000 (O_2000,N_16318,N_19939);
or UO_2001 (O_2001,N_19386,N_19021);
and UO_2002 (O_2002,N_18791,N_17681);
and UO_2003 (O_2003,N_18366,N_18955);
nand UO_2004 (O_2004,N_17389,N_17164);
nand UO_2005 (O_2005,N_19448,N_17805);
xnor UO_2006 (O_2006,N_19599,N_17618);
or UO_2007 (O_2007,N_19349,N_16826);
xnor UO_2008 (O_2008,N_17185,N_19068);
xnor UO_2009 (O_2009,N_17528,N_17379);
xor UO_2010 (O_2010,N_17055,N_16088);
nand UO_2011 (O_2011,N_19148,N_17287);
or UO_2012 (O_2012,N_17524,N_19599);
and UO_2013 (O_2013,N_18373,N_17901);
nor UO_2014 (O_2014,N_19601,N_17398);
and UO_2015 (O_2015,N_16171,N_18614);
nor UO_2016 (O_2016,N_18122,N_16999);
nor UO_2017 (O_2017,N_17290,N_18265);
or UO_2018 (O_2018,N_19838,N_19265);
or UO_2019 (O_2019,N_18126,N_19310);
nand UO_2020 (O_2020,N_17571,N_18033);
or UO_2021 (O_2021,N_18866,N_19048);
and UO_2022 (O_2022,N_18331,N_16786);
and UO_2023 (O_2023,N_16938,N_18902);
or UO_2024 (O_2024,N_19149,N_16289);
xor UO_2025 (O_2025,N_16754,N_18598);
xor UO_2026 (O_2026,N_16436,N_19333);
nand UO_2027 (O_2027,N_17760,N_19999);
or UO_2028 (O_2028,N_18945,N_17560);
xnor UO_2029 (O_2029,N_18018,N_18453);
xor UO_2030 (O_2030,N_16238,N_17729);
nor UO_2031 (O_2031,N_17819,N_18494);
and UO_2032 (O_2032,N_18162,N_17808);
and UO_2033 (O_2033,N_17792,N_19719);
and UO_2034 (O_2034,N_17955,N_19818);
xnor UO_2035 (O_2035,N_16732,N_19685);
nand UO_2036 (O_2036,N_19071,N_16452);
and UO_2037 (O_2037,N_18706,N_18108);
nor UO_2038 (O_2038,N_18718,N_17091);
nand UO_2039 (O_2039,N_18885,N_17224);
nand UO_2040 (O_2040,N_18240,N_18827);
and UO_2041 (O_2041,N_18748,N_17331);
nand UO_2042 (O_2042,N_18192,N_18713);
nand UO_2043 (O_2043,N_19931,N_19575);
and UO_2044 (O_2044,N_19170,N_16764);
nor UO_2045 (O_2045,N_19644,N_19153);
xor UO_2046 (O_2046,N_18684,N_19798);
nand UO_2047 (O_2047,N_18649,N_17593);
and UO_2048 (O_2048,N_17033,N_16471);
xnor UO_2049 (O_2049,N_16643,N_18877);
nand UO_2050 (O_2050,N_17693,N_19954);
or UO_2051 (O_2051,N_19066,N_16756);
xnor UO_2052 (O_2052,N_16498,N_19910);
nand UO_2053 (O_2053,N_18665,N_19691);
xnor UO_2054 (O_2054,N_16547,N_16714);
xor UO_2055 (O_2055,N_19464,N_19722);
nand UO_2056 (O_2056,N_19686,N_17074);
nor UO_2057 (O_2057,N_18093,N_16573);
or UO_2058 (O_2058,N_17990,N_18807);
nor UO_2059 (O_2059,N_19819,N_19813);
nor UO_2060 (O_2060,N_17413,N_16978);
or UO_2061 (O_2061,N_18685,N_17712);
xor UO_2062 (O_2062,N_18331,N_16583);
or UO_2063 (O_2063,N_17638,N_19176);
and UO_2064 (O_2064,N_17860,N_18092);
nor UO_2065 (O_2065,N_18131,N_16350);
nand UO_2066 (O_2066,N_16117,N_19692);
xnor UO_2067 (O_2067,N_18205,N_16933);
nand UO_2068 (O_2068,N_16959,N_19309);
nor UO_2069 (O_2069,N_19911,N_17925);
nand UO_2070 (O_2070,N_19590,N_18198);
or UO_2071 (O_2071,N_18996,N_16924);
or UO_2072 (O_2072,N_16325,N_16790);
xor UO_2073 (O_2073,N_19407,N_19788);
and UO_2074 (O_2074,N_19618,N_18391);
xnor UO_2075 (O_2075,N_16247,N_17354);
nand UO_2076 (O_2076,N_17038,N_19558);
nor UO_2077 (O_2077,N_17169,N_18180);
or UO_2078 (O_2078,N_16182,N_18261);
xnor UO_2079 (O_2079,N_19227,N_19381);
and UO_2080 (O_2080,N_16829,N_17777);
xor UO_2081 (O_2081,N_17997,N_17635);
or UO_2082 (O_2082,N_18230,N_17706);
xor UO_2083 (O_2083,N_16939,N_18987);
and UO_2084 (O_2084,N_16252,N_19141);
nor UO_2085 (O_2085,N_19571,N_16406);
nor UO_2086 (O_2086,N_17540,N_19399);
or UO_2087 (O_2087,N_16320,N_16720);
nor UO_2088 (O_2088,N_18159,N_17126);
and UO_2089 (O_2089,N_16133,N_17051);
xnor UO_2090 (O_2090,N_17069,N_17788);
nor UO_2091 (O_2091,N_19241,N_17941);
nor UO_2092 (O_2092,N_19988,N_17885);
and UO_2093 (O_2093,N_19905,N_19555);
and UO_2094 (O_2094,N_19498,N_16883);
or UO_2095 (O_2095,N_19285,N_16499);
and UO_2096 (O_2096,N_18272,N_16926);
or UO_2097 (O_2097,N_19047,N_16752);
xor UO_2098 (O_2098,N_19277,N_19086);
nand UO_2099 (O_2099,N_16176,N_18690);
nand UO_2100 (O_2100,N_18637,N_19849);
and UO_2101 (O_2101,N_18308,N_16646);
xor UO_2102 (O_2102,N_16003,N_18678);
and UO_2103 (O_2103,N_17642,N_17530);
and UO_2104 (O_2104,N_19715,N_19000);
or UO_2105 (O_2105,N_16857,N_16593);
nor UO_2106 (O_2106,N_19460,N_18194);
and UO_2107 (O_2107,N_16580,N_17997);
nor UO_2108 (O_2108,N_19370,N_19368);
nor UO_2109 (O_2109,N_18949,N_17240);
nand UO_2110 (O_2110,N_18002,N_17078);
nor UO_2111 (O_2111,N_17010,N_18888);
xor UO_2112 (O_2112,N_16045,N_16930);
and UO_2113 (O_2113,N_18438,N_18683);
or UO_2114 (O_2114,N_18891,N_19569);
xnor UO_2115 (O_2115,N_17363,N_19430);
and UO_2116 (O_2116,N_19305,N_19250);
nand UO_2117 (O_2117,N_16625,N_19598);
or UO_2118 (O_2118,N_16830,N_18596);
nand UO_2119 (O_2119,N_17067,N_18033);
and UO_2120 (O_2120,N_19567,N_17756);
xor UO_2121 (O_2121,N_19035,N_17815);
nand UO_2122 (O_2122,N_18461,N_18259);
xor UO_2123 (O_2123,N_19306,N_19521);
nor UO_2124 (O_2124,N_18112,N_16694);
or UO_2125 (O_2125,N_17115,N_19958);
nand UO_2126 (O_2126,N_19668,N_17162);
and UO_2127 (O_2127,N_18214,N_18967);
xor UO_2128 (O_2128,N_17762,N_18944);
and UO_2129 (O_2129,N_16171,N_16312);
nand UO_2130 (O_2130,N_18187,N_19632);
xnor UO_2131 (O_2131,N_17038,N_16150);
nand UO_2132 (O_2132,N_19843,N_18951);
nand UO_2133 (O_2133,N_19243,N_16152);
xnor UO_2134 (O_2134,N_19965,N_19375);
nor UO_2135 (O_2135,N_17021,N_19075);
or UO_2136 (O_2136,N_18846,N_18840);
nor UO_2137 (O_2137,N_18878,N_16307);
nand UO_2138 (O_2138,N_18696,N_18005);
or UO_2139 (O_2139,N_17564,N_19487);
or UO_2140 (O_2140,N_16470,N_17082);
nor UO_2141 (O_2141,N_17057,N_17892);
xor UO_2142 (O_2142,N_18470,N_16083);
nand UO_2143 (O_2143,N_17704,N_18052);
nor UO_2144 (O_2144,N_17000,N_18249);
or UO_2145 (O_2145,N_16603,N_16673);
nor UO_2146 (O_2146,N_17629,N_17888);
and UO_2147 (O_2147,N_19368,N_19202);
xor UO_2148 (O_2148,N_17990,N_16210);
or UO_2149 (O_2149,N_16661,N_19441);
and UO_2150 (O_2150,N_18969,N_18422);
nor UO_2151 (O_2151,N_19213,N_16290);
nand UO_2152 (O_2152,N_19443,N_18805);
or UO_2153 (O_2153,N_19546,N_18362);
xor UO_2154 (O_2154,N_16128,N_18517);
or UO_2155 (O_2155,N_18264,N_18996);
or UO_2156 (O_2156,N_19267,N_16697);
or UO_2157 (O_2157,N_16898,N_18136);
and UO_2158 (O_2158,N_18877,N_16693);
nor UO_2159 (O_2159,N_16243,N_18086);
xnor UO_2160 (O_2160,N_19187,N_18742);
or UO_2161 (O_2161,N_18207,N_16526);
or UO_2162 (O_2162,N_18510,N_16471);
and UO_2163 (O_2163,N_17892,N_19275);
nor UO_2164 (O_2164,N_18966,N_18690);
nand UO_2165 (O_2165,N_19054,N_17320);
nand UO_2166 (O_2166,N_18004,N_19667);
xor UO_2167 (O_2167,N_19903,N_18106);
nand UO_2168 (O_2168,N_16236,N_17478);
or UO_2169 (O_2169,N_19999,N_17916);
nand UO_2170 (O_2170,N_19177,N_17920);
or UO_2171 (O_2171,N_18880,N_18323);
xor UO_2172 (O_2172,N_19233,N_18309);
and UO_2173 (O_2173,N_16437,N_17190);
xnor UO_2174 (O_2174,N_16705,N_16622);
nand UO_2175 (O_2175,N_19301,N_16197);
and UO_2176 (O_2176,N_17531,N_16668);
xnor UO_2177 (O_2177,N_19641,N_18300);
nor UO_2178 (O_2178,N_16954,N_19542);
and UO_2179 (O_2179,N_16687,N_16050);
and UO_2180 (O_2180,N_16094,N_18076);
or UO_2181 (O_2181,N_19844,N_16878);
nand UO_2182 (O_2182,N_19314,N_19960);
nand UO_2183 (O_2183,N_17951,N_17319);
nor UO_2184 (O_2184,N_18027,N_16230);
nand UO_2185 (O_2185,N_18839,N_18569);
nand UO_2186 (O_2186,N_17415,N_18074);
or UO_2187 (O_2187,N_16119,N_18466);
or UO_2188 (O_2188,N_17355,N_19331);
xor UO_2189 (O_2189,N_18864,N_16038);
or UO_2190 (O_2190,N_17654,N_17355);
or UO_2191 (O_2191,N_17293,N_16330);
xor UO_2192 (O_2192,N_17037,N_16729);
xor UO_2193 (O_2193,N_16860,N_18839);
nand UO_2194 (O_2194,N_17496,N_18749);
xnor UO_2195 (O_2195,N_16018,N_17165);
or UO_2196 (O_2196,N_17765,N_19572);
nor UO_2197 (O_2197,N_17726,N_17639);
nor UO_2198 (O_2198,N_17187,N_18718);
nor UO_2199 (O_2199,N_17042,N_17452);
and UO_2200 (O_2200,N_17628,N_18379);
nor UO_2201 (O_2201,N_18417,N_18813);
or UO_2202 (O_2202,N_18375,N_19975);
nor UO_2203 (O_2203,N_17627,N_18144);
xor UO_2204 (O_2204,N_19494,N_17533);
nor UO_2205 (O_2205,N_18119,N_18767);
and UO_2206 (O_2206,N_17555,N_19005);
xor UO_2207 (O_2207,N_19668,N_17730);
nor UO_2208 (O_2208,N_16078,N_19613);
xnor UO_2209 (O_2209,N_16952,N_17751);
xnor UO_2210 (O_2210,N_17345,N_18708);
nand UO_2211 (O_2211,N_19474,N_19694);
nor UO_2212 (O_2212,N_19508,N_16586);
xor UO_2213 (O_2213,N_16051,N_17117);
or UO_2214 (O_2214,N_19600,N_19716);
and UO_2215 (O_2215,N_16414,N_17819);
and UO_2216 (O_2216,N_16146,N_18320);
or UO_2217 (O_2217,N_16825,N_16920);
nand UO_2218 (O_2218,N_16994,N_17377);
or UO_2219 (O_2219,N_17863,N_19589);
nand UO_2220 (O_2220,N_18016,N_19048);
and UO_2221 (O_2221,N_19317,N_16073);
nand UO_2222 (O_2222,N_18861,N_17441);
or UO_2223 (O_2223,N_17130,N_18467);
nor UO_2224 (O_2224,N_18512,N_18178);
nor UO_2225 (O_2225,N_16969,N_16179);
or UO_2226 (O_2226,N_16027,N_16934);
or UO_2227 (O_2227,N_16271,N_16042);
or UO_2228 (O_2228,N_18944,N_18416);
or UO_2229 (O_2229,N_19204,N_18863);
nor UO_2230 (O_2230,N_18733,N_17816);
and UO_2231 (O_2231,N_16437,N_18974);
or UO_2232 (O_2232,N_19101,N_19470);
xnor UO_2233 (O_2233,N_16070,N_19678);
xnor UO_2234 (O_2234,N_16396,N_18952);
nor UO_2235 (O_2235,N_18587,N_18388);
nor UO_2236 (O_2236,N_16225,N_16147);
xnor UO_2237 (O_2237,N_17688,N_17625);
and UO_2238 (O_2238,N_19940,N_16137);
and UO_2239 (O_2239,N_17334,N_17597);
xnor UO_2240 (O_2240,N_19426,N_19651);
nor UO_2241 (O_2241,N_17945,N_17712);
xor UO_2242 (O_2242,N_17530,N_19759);
nor UO_2243 (O_2243,N_19028,N_17918);
nand UO_2244 (O_2244,N_17810,N_18575);
or UO_2245 (O_2245,N_17484,N_16987);
xor UO_2246 (O_2246,N_16238,N_18190);
nand UO_2247 (O_2247,N_19297,N_19683);
nor UO_2248 (O_2248,N_16812,N_16575);
nand UO_2249 (O_2249,N_17786,N_16815);
nand UO_2250 (O_2250,N_17159,N_19719);
or UO_2251 (O_2251,N_18059,N_16292);
and UO_2252 (O_2252,N_19039,N_16057);
nand UO_2253 (O_2253,N_16541,N_18740);
and UO_2254 (O_2254,N_17523,N_16534);
nor UO_2255 (O_2255,N_19871,N_18082);
nand UO_2256 (O_2256,N_18141,N_18522);
nand UO_2257 (O_2257,N_19220,N_18095);
nor UO_2258 (O_2258,N_18254,N_17023);
or UO_2259 (O_2259,N_16449,N_16249);
nor UO_2260 (O_2260,N_16979,N_19675);
xnor UO_2261 (O_2261,N_16066,N_16579);
xor UO_2262 (O_2262,N_17498,N_16902);
nand UO_2263 (O_2263,N_17104,N_19905);
nor UO_2264 (O_2264,N_18312,N_16683);
and UO_2265 (O_2265,N_17059,N_18596);
nand UO_2266 (O_2266,N_16505,N_19025);
nand UO_2267 (O_2267,N_19194,N_16638);
nor UO_2268 (O_2268,N_18689,N_16670);
or UO_2269 (O_2269,N_17400,N_18104);
nor UO_2270 (O_2270,N_19982,N_17147);
nor UO_2271 (O_2271,N_18240,N_17065);
nand UO_2272 (O_2272,N_16678,N_17681);
nor UO_2273 (O_2273,N_18700,N_18071);
and UO_2274 (O_2274,N_17626,N_16340);
xnor UO_2275 (O_2275,N_18665,N_17643);
or UO_2276 (O_2276,N_16758,N_16595);
nand UO_2277 (O_2277,N_19458,N_19327);
and UO_2278 (O_2278,N_18066,N_18874);
nor UO_2279 (O_2279,N_19147,N_17573);
nor UO_2280 (O_2280,N_17697,N_16481);
and UO_2281 (O_2281,N_17956,N_19230);
nor UO_2282 (O_2282,N_19844,N_17101);
and UO_2283 (O_2283,N_19540,N_19397);
xnor UO_2284 (O_2284,N_18370,N_19502);
and UO_2285 (O_2285,N_16816,N_18345);
and UO_2286 (O_2286,N_16097,N_19144);
nand UO_2287 (O_2287,N_18957,N_17065);
nor UO_2288 (O_2288,N_18446,N_19505);
and UO_2289 (O_2289,N_16965,N_16106);
nor UO_2290 (O_2290,N_19048,N_17689);
or UO_2291 (O_2291,N_19039,N_18410);
nand UO_2292 (O_2292,N_19933,N_19328);
nand UO_2293 (O_2293,N_16656,N_17295);
or UO_2294 (O_2294,N_18258,N_19086);
and UO_2295 (O_2295,N_16658,N_19474);
nand UO_2296 (O_2296,N_17195,N_18356);
nand UO_2297 (O_2297,N_17089,N_19363);
nor UO_2298 (O_2298,N_18336,N_18882);
and UO_2299 (O_2299,N_19772,N_16840);
or UO_2300 (O_2300,N_17954,N_16310);
nand UO_2301 (O_2301,N_18426,N_19186);
or UO_2302 (O_2302,N_16098,N_16376);
and UO_2303 (O_2303,N_18997,N_18429);
xor UO_2304 (O_2304,N_19175,N_18304);
or UO_2305 (O_2305,N_16565,N_17022);
and UO_2306 (O_2306,N_16244,N_18071);
and UO_2307 (O_2307,N_16046,N_16501);
and UO_2308 (O_2308,N_16763,N_16553);
nor UO_2309 (O_2309,N_17973,N_18658);
nand UO_2310 (O_2310,N_17808,N_19891);
xor UO_2311 (O_2311,N_16010,N_16933);
and UO_2312 (O_2312,N_18164,N_16517);
xnor UO_2313 (O_2313,N_17926,N_17312);
xor UO_2314 (O_2314,N_19104,N_19462);
nor UO_2315 (O_2315,N_19462,N_16843);
and UO_2316 (O_2316,N_19743,N_19512);
nor UO_2317 (O_2317,N_16777,N_18251);
and UO_2318 (O_2318,N_19859,N_18547);
or UO_2319 (O_2319,N_19908,N_18811);
or UO_2320 (O_2320,N_18337,N_17533);
nor UO_2321 (O_2321,N_18819,N_18608);
nand UO_2322 (O_2322,N_18167,N_17875);
nand UO_2323 (O_2323,N_19980,N_17131);
xnor UO_2324 (O_2324,N_16676,N_18250);
nor UO_2325 (O_2325,N_19032,N_17600);
nand UO_2326 (O_2326,N_18717,N_17196);
nand UO_2327 (O_2327,N_17437,N_19092);
nor UO_2328 (O_2328,N_16738,N_19744);
nand UO_2329 (O_2329,N_19562,N_19765);
xor UO_2330 (O_2330,N_18716,N_16978);
nor UO_2331 (O_2331,N_19853,N_18068);
and UO_2332 (O_2332,N_16331,N_16260);
nor UO_2333 (O_2333,N_16814,N_19796);
or UO_2334 (O_2334,N_17822,N_19341);
nand UO_2335 (O_2335,N_17748,N_19118);
xnor UO_2336 (O_2336,N_18322,N_16470);
xnor UO_2337 (O_2337,N_19366,N_17666);
xor UO_2338 (O_2338,N_18123,N_19164);
nor UO_2339 (O_2339,N_17324,N_16600);
xnor UO_2340 (O_2340,N_19837,N_16663);
and UO_2341 (O_2341,N_19398,N_16849);
nand UO_2342 (O_2342,N_18924,N_18749);
nor UO_2343 (O_2343,N_18642,N_18142);
or UO_2344 (O_2344,N_16345,N_16666);
nor UO_2345 (O_2345,N_16065,N_19796);
or UO_2346 (O_2346,N_17270,N_19387);
nor UO_2347 (O_2347,N_19124,N_17060);
or UO_2348 (O_2348,N_18222,N_18295);
or UO_2349 (O_2349,N_17584,N_16467);
and UO_2350 (O_2350,N_17250,N_17623);
nand UO_2351 (O_2351,N_17619,N_19507);
nand UO_2352 (O_2352,N_19018,N_16541);
or UO_2353 (O_2353,N_17419,N_19705);
nand UO_2354 (O_2354,N_16640,N_16846);
or UO_2355 (O_2355,N_18774,N_19066);
nand UO_2356 (O_2356,N_16677,N_16908);
xor UO_2357 (O_2357,N_18832,N_19241);
nor UO_2358 (O_2358,N_16187,N_17269);
xor UO_2359 (O_2359,N_19553,N_16064);
nor UO_2360 (O_2360,N_16414,N_17132);
and UO_2361 (O_2361,N_16395,N_19486);
nor UO_2362 (O_2362,N_18978,N_18711);
or UO_2363 (O_2363,N_17673,N_18707);
and UO_2364 (O_2364,N_16582,N_18190);
nand UO_2365 (O_2365,N_16018,N_18217);
nor UO_2366 (O_2366,N_18122,N_16166);
nand UO_2367 (O_2367,N_19961,N_16014);
and UO_2368 (O_2368,N_19657,N_18744);
nor UO_2369 (O_2369,N_19733,N_19279);
and UO_2370 (O_2370,N_16010,N_18006);
nand UO_2371 (O_2371,N_17767,N_16598);
nor UO_2372 (O_2372,N_17308,N_18324);
or UO_2373 (O_2373,N_18288,N_17610);
nor UO_2374 (O_2374,N_18897,N_17220);
xnor UO_2375 (O_2375,N_16289,N_19143);
xor UO_2376 (O_2376,N_18392,N_17901);
nor UO_2377 (O_2377,N_18420,N_17512);
or UO_2378 (O_2378,N_19529,N_17248);
xor UO_2379 (O_2379,N_19470,N_18712);
and UO_2380 (O_2380,N_16833,N_19368);
xnor UO_2381 (O_2381,N_16030,N_17332);
or UO_2382 (O_2382,N_17175,N_19537);
nand UO_2383 (O_2383,N_18931,N_17102);
nor UO_2384 (O_2384,N_18228,N_17771);
and UO_2385 (O_2385,N_19716,N_16555);
or UO_2386 (O_2386,N_16604,N_18059);
or UO_2387 (O_2387,N_16371,N_16241);
nor UO_2388 (O_2388,N_16171,N_16466);
and UO_2389 (O_2389,N_19985,N_16414);
xnor UO_2390 (O_2390,N_17308,N_18863);
and UO_2391 (O_2391,N_16275,N_19471);
xnor UO_2392 (O_2392,N_17239,N_18538);
xnor UO_2393 (O_2393,N_16158,N_17246);
or UO_2394 (O_2394,N_18729,N_19070);
and UO_2395 (O_2395,N_17708,N_19663);
and UO_2396 (O_2396,N_16260,N_18607);
nor UO_2397 (O_2397,N_17714,N_17240);
nand UO_2398 (O_2398,N_18305,N_17371);
and UO_2399 (O_2399,N_16246,N_16631);
and UO_2400 (O_2400,N_18642,N_19660);
and UO_2401 (O_2401,N_17168,N_16470);
nand UO_2402 (O_2402,N_18783,N_19345);
nand UO_2403 (O_2403,N_17590,N_19974);
nor UO_2404 (O_2404,N_18325,N_18395);
nor UO_2405 (O_2405,N_16631,N_19851);
and UO_2406 (O_2406,N_17670,N_17974);
nor UO_2407 (O_2407,N_16981,N_16803);
nand UO_2408 (O_2408,N_16595,N_18855);
and UO_2409 (O_2409,N_16897,N_19484);
or UO_2410 (O_2410,N_17673,N_16197);
xnor UO_2411 (O_2411,N_18852,N_16872);
xnor UO_2412 (O_2412,N_18648,N_16186);
nand UO_2413 (O_2413,N_17370,N_19615);
nand UO_2414 (O_2414,N_17623,N_17495);
and UO_2415 (O_2415,N_17298,N_19224);
and UO_2416 (O_2416,N_16277,N_18154);
nand UO_2417 (O_2417,N_19723,N_16407);
nand UO_2418 (O_2418,N_17460,N_17742);
nor UO_2419 (O_2419,N_17420,N_18765);
xnor UO_2420 (O_2420,N_16898,N_17894);
and UO_2421 (O_2421,N_17300,N_17320);
nor UO_2422 (O_2422,N_18971,N_17139);
nand UO_2423 (O_2423,N_17713,N_18820);
and UO_2424 (O_2424,N_16850,N_17926);
or UO_2425 (O_2425,N_16756,N_19793);
nor UO_2426 (O_2426,N_16860,N_17955);
nor UO_2427 (O_2427,N_18565,N_19134);
xnor UO_2428 (O_2428,N_17499,N_18501);
xnor UO_2429 (O_2429,N_16116,N_17761);
and UO_2430 (O_2430,N_17684,N_19629);
and UO_2431 (O_2431,N_18053,N_17948);
nand UO_2432 (O_2432,N_18388,N_19158);
xor UO_2433 (O_2433,N_17031,N_16896);
and UO_2434 (O_2434,N_17534,N_17828);
or UO_2435 (O_2435,N_19543,N_16698);
or UO_2436 (O_2436,N_17974,N_16710);
nor UO_2437 (O_2437,N_16620,N_19736);
nor UO_2438 (O_2438,N_17448,N_16241);
nand UO_2439 (O_2439,N_18310,N_17609);
nor UO_2440 (O_2440,N_19563,N_18359);
or UO_2441 (O_2441,N_18851,N_16141);
and UO_2442 (O_2442,N_17383,N_17592);
and UO_2443 (O_2443,N_18625,N_17624);
and UO_2444 (O_2444,N_19338,N_16453);
nor UO_2445 (O_2445,N_19769,N_18326);
xnor UO_2446 (O_2446,N_18143,N_17145);
and UO_2447 (O_2447,N_19353,N_18305);
or UO_2448 (O_2448,N_16206,N_19954);
nand UO_2449 (O_2449,N_16965,N_16705);
nor UO_2450 (O_2450,N_16825,N_19691);
xor UO_2451 (O_2451,N_18297,N_17814);
xnor UO_2452 (O_2452,N_18060,N_16873);
or UO_2453 (O_2453,N_18137,N_18512);
nand UO_2454 (O_2454,N_19303,N_17387);
nand UO_2455 (O_2455,N_16736,N_17246);
or UO_2456 (O_2456,N_16431,N_19004);
nor UO_2457 (O_2457,N_17715,N_17008);
xor UO_2458 (O_2458,N_18404,N_17256);
and UO_2459 (O_2459,N_18116,N_17113);
nand UO_2460 (O_2460,N_19240,N_16944);
nand UO_2461 (O_2461,N_18528,N_17344);
nand UO_2462 (O_2462,N_17913,N_17198);
nor UO_2463 (O_2463,N_16708,N_19008);
nand UO_2464 (O_2464,N_17232,N_17087);
xnor UO_2465 (O_2465,N_19210,N_17005);
and UO_2466 (O_2466,N_19804,N_17047);
nor UO_2467 (O_2467,N_19131,N_17119);
xor UO_2468 (O_2468,N_19904,N_17949);
nor UO_2469 (O_2469,N_17434,N_17076);
and UO_2470 (O_2470,N_17916,N_19861);
nor UO_2471 (O_2471,N_19148,N_18447);
nor UO_2472 (O_2472,N_17578,N_17069);
or UO_2473 (O_2473,N_19025,N_19669);
nor UO_2474 (O_2474,N_19492,N_16037);
nor UO_2475 (O_2475,N_17240,N_17209);
xor UO_2476 (O_2476,N_19212,N_17175);
xor UO_2477 (O_2477,N_18742,N_18084);
xnor UO_2478 (O_2478,N_19320,N_19988);
or UO_2479 (O_2479,N_19405,N_19716);
nand UO_2480 (O_2480,N_16032,N_16847);
and UO_2481 (O_2481,N_18831,N_19297);
nand UO_2482 (O_2482,N_16431,N_17568);
nand UO_2483 (O_2483,N_16894,N_16466);
or UO_2484 (O_2484,N_18795,N_18811);
nor UO_2485 (O_2485,N_16617,N_17027);
nand UO_2486 (O_2486,N_18610,N_17395);
or UO_2487 (O_2487,N_19526,N_19970);
nand UO_2488 (O_2488,N_17234,N_16435);
nand UO_2489 (O_2489,N_16088,N_19572);
xnor UO_2490 (O_2490,N_16555,N_18155);
and UO_2491 (O_2491,N_17578,N_16924);
xor UO_2492 (O_2492,N_18146,N_18078);
nor UO_2493 (O_2493,N_16174,N_18694);
and UO_2494 (O_2494,N_18117,N_19077);
nand UO_2495 (O_2495,N_16519,N_16240);
or UO_2496 (O_2496,N_19765,N_19342);
nand UO_2497 (O_2497,N_19640,N_18428);
or UO_2498 (O_2498,N_17635,N_17874);
or UO_2499 (O_2499,N_19620,N_18642);
endmodule