module basic_2500_25000_3000_25_levels_10xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
xnor U0 (N_0,In_1543,In_456);
and U1 (N_1,In_1801,In_1035);
and U2 (N_2,In_1684,In_210);
nor U3 (N_3,In_48,In_941);
nor U4 (N_4,In_2010,In_1146);
and U5 (N_5,In_305,In_974);
xnor U6 (N_6,In_1574,In_1904);
or U7 (N_7,In_188,In_814);
xnor U8 (N_8,In_1631,In_564);
and U9 (N_9,In_1996,In_1569);
xor U10 (N_10,In_135,In_2117);
nor U11 (N_11,In_1214,In_866);
and U12 (N_12,In_1320,In_98);
and U13 (N_13,In_2440,In_2339);
and U14 (N_14,In_1940,In_1432);
nand U15 (N_15,In_2093,In_620);
and U16 (N_16,In_375,In_2026);
and U17 (N_17,In_2143,In_2024);
xnor U18 (N_18,In_948,In_2420);
nand U19 (N_19,In_1336,In_1887);
and U20 (N_20,In_813,In_2139);
and U21 (N_21,In_2182,In_1944);
nor U22 (N_22,In_114,In_1341);
xnor U23 (N_23,In_398,In_657);
or U24 (N_24,In_1696,In_1816);
or U25 (N_25,In_736,In_1502);
and U26 (N_26,In_2091,In_651);
nand U27 (N_27,In_47,In_1809);
or U28 (N_28,In_1170,In_1774);
and U29 (N_29,In_95,In_1388);
nor U30 (N_30,In_220,In_1786);
or U31 (N_31,In_1804,In_414);
nor U32 (N_32,In_655,In_1100);
nor U33 (N_33,In_1640,In_998);
xor U34 (N_34,In_1261,In_2307);
nor U35 (N_35,In_827,In_1163);
or U36 (N_36,In_2118,In_1579);
nor U37 (N_37,In_1938,In_1882);
xor U38 (N_38,In_2385,In_2203);
nor U39 (N_39,In_1375,In_1417);
nor U40 (N_40,In_2160,In_1527);
nor U41 (N_41,In_2373,In_1329);
or U42 (N_42,In_1441,In_99);
nor U43 (N_43,In_1557,In_1082);
nand U44 (N_44,In_895,In_1843);
and U45 (N_45,In_1853,In_2430);
nand U46 (N_46,In_1342,In_1354);
xnor U47 (N_47,In_246,In_1326);
or U48 (N_48,In_401,In_692);
nand U49 (N_49,In_1971,In_708);
xnor U50 (N_50,In_275,In_2067);
nor U51 (N_51,In_1637,In_390);
xnor U52 (N_52,In_2011,In_1902);
nor U53 (N_53,In_1202,In_2248);
nand U54 (N_54,In_1443,In_2166);
or U55 (N_55,In_491,In_1067);
xnor U56 (N_56,In_323,In_1888);
nand U57 (N_57,In_1807,In_572);
and U58 (N_58,In_803,In_1611);
nor U59 (N_59,In_1113,In_472);
nor U60 (N_60,In_215,In_1901);
or U61 (N_61,In_2424,In_1681);
xnor U62 (N_62,In_1570,In_1991);
or U63 (N_63,In_1111,In_2333);
and U64 (N_64,In_77,In_820);
and U65 (N_65,In_344,In_2153);
xor U66 (N_66,In_1104,In_1612);
and U67 (N_67,In_1132,In_810);
and U68 (N_68,In_183,In_920);
and U69 (N_69,In_855,In_2382);
and U70 (N_70,In_1366,In_2443);
nor U71 (N_71,In_1437,In_562);
xnor U72 (N_72,In_635,In_962);
nor U73 (N_73,In_806,In_2379);
or U74 (N_74,In_724,In_2049);
nor U75 (N_75,In_501,In_928);
nand U76 (N_76,In_1221,In_662);
xor U77 (N_77,In_451,In_2018);
xor U78 (N_78,In_2051,In_1721);
nand U79 (N_79,In_1308,In_1201);
nor U80 (N_80,In_347,In_85);
nand U81 (N_81,In_417,In_2004);
or U82 (N_82,In_2404,In_2372);
or U83 (N_83,In_990,In_2343);
nand U84 (N_84,In_745,In_882);
nor U85 (N_85,In_1239,In_487);
nor U86 (N_86,In_1302,In_167);
xor U87 (N_87,In_881,In_2208);
nor U88 (N_88,In_2247,In_335);
or U89 (N_89,In_1535,In_2156);
nand U90 (N_90,In_1852,In_113);
and U91 (N_91,In_1226,In_2036);
nand U92 (N_92,In_968,In_252);
nand U93 (N_93,In_2233,In_1572);
xnor U94 (N_94,In_1920,In_1470);
or U95 (N_95,In_25,In_730);
and U96 (N_96,In_2212,In_1649);
nor U97 (N_97,In_823,In_971);
xnor U98 (N_98,In_1269,In_1875);
and U99 (N_99,In_2453,In_1498);
or U100 (N_100,In_1447,In_1032);
nand U101 (N_101,In_1044,In_925);
nand U102 (N_102,In_2187,In_1409);
or U103 (N_103,In_1339,In_303);
nand U104 (N_104,In_2486,In_32);
nand U105 (N_105,In_1648,In_2330);
xor U106 (N_106,In_1069,In_140);
or U107 (N_107,In_461,In_1373);
xnor U108 (N_108,In_269,In_1015);
or U109 (N_109,In_1423,In_1974);
xnor U110 (N_110,In_1322,In_2068);
nor U111 (N_111,In_2371,In_1824);
and U112 (N_112,In_1379,In_1566);
xnor U113 (N_113,In_544,In_294);
xor U114 (N_114,In_2458,In_520);
xnor U115 (N_115,In_763,In_2106);
and U116 (N_116,In_342,In_890);
and U117 (N_117,In_939,In_1957);
xnor U118 (N_118,In_2450,In_2176);
or U119 (N_119,In_2,In_2304);
nor U120 (N_120,In_151,In_1103);
or U121 (N_121,In_2193,In_17);
nor U122 (N_122,In_727,In_673);
and U123 (N_123,In_30,In_1033);
xor U124 (N_124,In_475,In_309);
nor U125 (N_125,In_171,In_1118);
xnor U126 (N_126,In_1003,In_679);
and U127 (N_127,In_2146,In_178);
nor U128 (N_128,In_1532,In_1508);
nor U129 (N_129,In_79,In_63);
and U130 (N_130,In_2188,In_699);
nand U131 (N_131,In_299,In_1390);
xnor U132 (N_132,In_1777,In_1855);
and U133 (N_133,In_450,In_1751);
or U134 (N_134,In_1916,In_2083);
nand U135 (N_135,In_418,In_605);
nor U136 (N_136,In_1711,In_291);
nand U137 (N_137,In_1847,In_1400);
nor U138 (N_138,In_1646,In_1773);
nor U139 (N_139,In_467,In_1465);
or U140 (N_140,In_58,In_731);
nand U141 (N_141,In_365,In_921);
and U142 (N_142,In_903,In_510);
nand U143 (N_143,In_2251,In_1925);
nor U144 (N_144,In_1948,In_1550);
xor U145 (N_145,In_1183,In_283);
xnor U146 (N_146,In_583,In_1909);
or U147 (N_147,In_517,In_872);
and U148 (N_148,In_2115,In_1839);
nand U149 (N_149,In_2417,In_1528);
and U150 (N_150,In_1765,In_1522);
and U151 (N_151,In_2126,In_593);
nand U152 (N_152,In_1401,In_1333);
xor U153 (N_153,In_1934,In_954);
nor U154 (N_154,In_551,In_720);
nand U155 (N_155,In_1635,In_2078);
and U156 (N_156,In_1053,In_650);
nand U157 (N_157,In_1055,In_39);
or U158 (N_158,In_1314,In_908);
nand U159 (N_159,In_2294,In_2214);
nor U160 (N_160,In_1071,In_6);
nand U161 (N_161,In_1052,In_136);
or U162 (N_162,In_652,In_2129);
xnor U163 (N_163,In_691,In_359);
nand U164 (N_164,In_257,In_710);
nor U165 (N_165,In_1304,In_482);
or U166 (N_166,In_1674,In_805);
nor U167 (N_167,In_1990,In_1521);
or U168 (N_168,In_242,In_168);
and U169 (N_169,In_1062,In_2303);
and U170 (N_170,In_350,In_1506);
nor U171 (N_171,In_2386,In_924);
nor U172 (N_172,In_918,In_2133);
nand U173 (N_173,In_555,In_1252);
nand U174 (N_174,In_783,In_2398);
xor U175 (N_175,In_2013,In_1425);
or U176 (N_176,In_1324,In_2215);
nand U177 (N_177,In_221,In_1063);
and U178 (N_178,In_1361,In_513);
and U179 (N_179,In_654,In_1596);
and U180 (N_180,In_1496,In_2088);
or U181 (N_181,In_225,In_486);
nand U182 (N_182,In_849,In_1219);
nor U183 (N_183,In_1802,In_2313);
xnor U184 (N_184,In_1436,In_2235);
or U185 (N_185,In_386,In_802);
nand U186 (N_186,In_1090,In_914);
nand U187 (N_187,In_360,In_1131);
nor U188 (N_188,In_2394,In_277);
or U189 (N_189,In_1414,In_1228);
and U190 (N_190,In_729,In_2295);
xnor U191 (N_191,In_393,In_205);
and U192 (N_192,In_2447,In_818);
nor U193 (N_193,In_2489,In_112);
nand U194 (N_194,In_1884,In_880);
nand U195 (N_195,In_198,In_2270);
nand U196 (N_196,In_674,In_1286);
nand U197 (N_197,In_2042,In_1246);
or U198 (N_198,In_265,In_1293);
nor U199 (N_199,In_644,In_817);
nor U200 (N_200,In_781,In_1505);
or U201 (N_201,In_1583,In_1296);
xor U202 (N_202,In_2292,In_164);
and U203 (N_203,In_1262,In_177);
or U204 (N_204,In_666,In_1735);
xor U205 (N_205,In_1663,In_863);
nand U206 (N_206,In_1150,In_919);
nand U207 (N_207,In_1654,In_1472);
and U208 (N_208,In_2226,In_195);
xnor U209 (N_209,In_1769,In_946);
nor U210 (N_210,In_1958,In_685);
or U211 (N_211,In_1491,In_2100);
nand U212 (N_212,In_535,In_1713);
and U213 (N_213,In_1091,In_1725);
and U214 (N_214,In_1428,In_534);
xor U215 (N_215,In_762,In_2454);
and U216 (N_216,In_1924,In_2211);
or U217 (N_217,In_1985,In_1059);
and U218 (N_218,In_2484,In_922);
and U219 (N_219,In_1970,In_2320);
nand U220 (N_220,In_26,In_1259);
nor U221 (N_221,In_478,In_2259);
xor U222 (N_222,In_2397,In_2273);
and U223 (N_223,In_2015,In_495);
nand U224 (N_224,In_709,In_1374);
or U225 (N_225,In_1551,In_2380);
nand U226 (N_226,In_488,In_1636);
nor U227 (N_227,In_31,In_1714);
and U228 (N_228,In_1471,In_2475);
nor U229 (N_229,In_55,In_256);
nor U230 (N_230,In_1338,In_1863);
and U231 (N_231,In_332,In_4);
or U232 (N_232,In_1627,In_587);
nor U233 (N_233,In_172,In_1619);
nand U234 (N_234,In_851,In_2199);
nand U235 (N_235,In_2198,In_1664);
and U236 (N_236,In_2341,In_1935);
or U237 (N_237,In_841,In_407);
and U238 (N_238,In_1778,In_1537);
and U239 (N_239,In_91,In_1415);
nor U240 (N_240,In_1421,In_1891);
nor U241 (N_241,In_1145,In_2255);
xnor U242 (N_242,In_1832,In_1917);
xor U243 (N_243,In_1364,In_1510);
and U244 (N_244,In_141,In_2094);
nor U245 (N_245,In_696,In_1792);
nor U246 (N_246,In_2002,In_1873);
nand U247 (N_247,In_1668,In_237);
and U248 (N_248,In_774,In_592);
xor U249 (N_249,In_1600,In_473);
xnor U250 (N_250,In_1548,In_1712);
nor U251 (N_251,In_1248,In_664);
nor U252 (N_252,In_1750,In_2201);
and U253 (N_253,In_1656,In_2135);
xor U254 (N_254,In_875,In_2022);
nand U255 (N_255,In_2029,In_1160);
nor U256 (N_256,In_1586,In_2310);
or U257 (N_257,In_1355,In_1556);
or U258 (N_258,In_1467,In_78);
or U259 (N_259,In_485,In_1149);
xnor U260 (N_260,In_1722,In_1495);
and U261 (N_261,In_1965,In_2210);
nand U262 (N_262,In_2406,In_994);
xor U263 (N_263,In_728,In_2033);
and U264 (N_264,In_927,In_1346);
nand U265 (N_265,In_1301,In_1633);
or U266 (N_266,In_412,In_790);
or U267 (N_267,In_111,In_419);
nand U268 (N_268,In_1039,In_1718);
or U269 (N_269,In_1830,In_1729);
nand U270 (N_270,In_978,In_2047);
nand U271 (N_271,In_206,In_1678);
and U272 (N_272,In_2110,In_532);
nor U273 (N_273,In_1607,In_1348);
nand U274 (N_274,In_462,In_445);
xor U275 (N_275,In_93,In_259);
xnor U276 (N_276,In_1024,In_2323);
and U277 (N_277,In_1241,In_2039);
nand U278 (N_278,In_1615,In_293);
and U279 (N_279,In_598,In_1899);
or U280 (N_280,In_1790,In_563);
nand U281 (N_281,In_2085,In_1592);
nor U282 (N_282,In_1780,In_1710);
or U283 (N_283,In_1857,In_886);
nor U284 (N_284,In_23,In_577);
xor U285 (N_285,In_576,In_1726);
xor U286 (N_286,In_744,In_1826);
nand U287 (N_287,In_1240,In_1922);
and U288 (N_288,In_245,In_2261);
and U289 (N_289,In_1290,In_2137);
or U290 (N_290,In_2097,In_239);
xnor U291 (N_291,In_2240,In_1190);
nand U292 (N_292,In_408,In_2321);
nand U293 (N_293,In_1896,In_2325);
or U294 (N_294,In_263,In_1138);
or U295 (N_295,In_1509,In_379);
and U296 (N_296,In_1794,In_2046);
xor U297 (N_297,In_752,In_1672);
xnor U298 (N_298,In_1285,In_972);
nor U299 (N_299,In_898,In_759);
nor U300 (N_300,In_2441,In_2391);
xnor U301 (N_301,In_2482,In_1234);
nor U302 (N_302,In_1859,In_681);
nand U303 (N_303,In_1992,In_1943);
nor U304 (N_304,In_2322,In_1709);
nor U305 (N_305,In_1604,In_2467);
xor U306 (N_306,In_1994,In_527);
nor U307 (N_307,In_1109,In_1599);
nor U308 (N_308,In_270,In_933);
nand U309 (N_309,In_428,In_74);
and U310 (N_310,In_1783,In_2089);
or U311 (N_311,In_2128,In_2206);
nand U312 (N_312,In_279,In_1738);
and U313 (N_313,In_301,In_1087);
xor U314 (N_314,In_1497,In_137);
and U315 (N_315,In_1001,In_1016);
and U316 (N_316,In_2170,In_1143);
or U317 (N_317,In_2412,In_1800);
nor U318 (N_318,In_176,In_628);
and U319 (N_319,In_278,In_1317);
xnor U320 (N_320,In_590,In_2098);
or U321 (N_321,In_33,In_1733);
xnor U322 (N_322,In_1078,In_1838);
and U323 (N_323,In_509,In_2260);
or U324 (N_324,In_484,In_1232);
and U325 (N_325,In_1357,In_2005);
or U326 (N_326,In_497,In_1014);
xnor U327 (N_327,In_1629,In_45);
nor U328 (N_328,In_1533,In_1553);
xor U329 (N_329,In_1979,In_28);
and U330 (N_330,In_2014,In_1785);
or U331 (N_331,In_433,In_857);
nand U332 (N_332,In_16,In_1889);
and U333 (N_333,In_1237,In_2000);
and U334 (N_334,In_1813,In_2328);
nor U335 (N_335,In_159,In_2357);
nand U336 (N_336,In_396,In_846);
xor U337 (N_337,In_815,In_2185);
nor U338 (N_338,In_327,In_1503);
or U339 (N_339,In_798,In_1827);
or U340 (N_340,In_2334,In_2468);
xnor U341 (N_341,In_2369,In_713);
or U342 (N_342,In_334,In_1294);
nand U343 (N_343,In_1748,In_117);
nor U344 (N_344,In_339,In_464);
xnor U345 (N_345,In_333,In_66);
nor U346 (N_346,In_1076,In_394);
nor U347 (N_347,In_1687,In_1139);
nand U348 (N_348,In_2228,In_481);
or U349 (N_349,In_584,In_243);
nor U350 (N_350,In_247,In_1789);
and U351 (N_351,In_330,In_1455);
nor U352 (N_352,In_2315,In_1724);
nand U353 (N_353,In_434,In_411);
and U354 (N_354,In_741,In_2435);
and U355 (N_355,In_2449,In_378);
xor U356 (N_356,In_1265,In_2016);
nand U357 (N_357,In_1677,In_819);
xor U358 (N_358,In_1671,In_435);
or U359 (N_359,In_979,In_2293);
nand U360 (N_360,In_758,In_2058);
nor U361 (N_361,In_2238,In_2352);
and U362 (N_362,In_1110,In_1821);
xor U363 (N_363,In_1263,In_9);
and U364 (N_364,In_1197,In_1225);
xnor U365 (N_365,In_2066,In_530);
nor U366 (N_366,In_2123,In_1288);
and U367 (N_367,In_125,In_825);
xnor U368 (N_368,In_1208,In_697);
nor U369 (N_369,In_2216,In_2145);
xor U370 (N_370,In_1811,In_89);
xor U371 (N_371,In_1079,In_1858);
or U372 (N_372,In_1266,In_490);
or U373 (N_373,In_1999,In_1886);
xnor U374 (N_374,In_1689,In_1108);
and U375 (N_375,In_1484,In_1369);
nand U376 (N_376,In_770,In_2197);
nor U377 (N_377,In_719,In_558);
xnor U378 (N_378,In_2169,In_1845);
and U379 (N_379,In_1158,In_2473);
and U380 (N_380,In_2476,In_97);
and U381 (N_381,In_505,In_1823);
or U382 (N_382,In_1897,In_69);
or U383 (N_383,In_1584,In_1115);
xnor U384 (N_384,In_1960,In_1393);
nor U385 (N_385,In_2076,In_1998);
and U386 (N_386,In_958,In_2263);
or U387 (N_387,In_1861,In_1734);
xor U388 (N_388,In_702,In_2249);
nand U389 (N_389,In_714,In_2241);
and U390 (N_390,In_2130,In_2104);
nor U391 (N_391,In_1289,In_1616);
and U392 (N_392,In_575,In_100);
nand U393 (N_393,In_463,In_1568);
and U394 (N_394,In_284,In_372);
and U395 (N_395,In_694,In_1311);
nand U396 (N_396,In_868,In_1191);
and U397 (N_397,In_1475,In_883);
nand U398 (N_398,In_2237,In_374);
and U399 (N_399,In_1514,In_557);
nand U400 (N_400,In_1921,In_2021);
and U401 (N_401,In_2344,In_1112);
or U402 (N_402,In_2111,In_834);
xor U403 (N_403,In_2256,In_12);
xor U404 (N_404,In_203,In_2008);
nor U405 (N_405,In_2495,In_1731);
xnor U406 (N_406,In_1192,In_952);
xnor U407 (N_407,In_304,In_2455);
and U408 (N_408,In_973,In_2299);
nand U409 (N_409,In_816,In_123);
nor U410 (N_410,In_2102,In_1319);
and U411 (N_411,In_671,In_1647);
xnor U412 (N_412,In_642,In_906);
nand U413 (N_413,In_14,In_292);
nand U414 (N_414,In_2390,In_1590);
or U415 (N_415,In_1661,In_1485);
nor U416 (N_416,In_437,In_1791);
and U417 (N_417,In_355,In_1868);
and U418 (N_418,In_2284,In_2217);
or U419 (N_419,In_104,In_2485);
nand U420 (N_420,In_529,In_603);
or U421 (N_421,In_1385,In_1129);
or U422 (N_422,In_1772,In_1598);
and U423 (N_423,In_2470,In_615);
nor U424 (N_424,In_224,In_2491);
and U425 (N_425,In_452,In_170);
xnor U426 (N_426,In_1490,In_2116);
or U427 (N_427,In_1235,In_1563);
nor U428 (N_428,In_413,In_316);
or U429 (N_429,In_1595,In_1699);
nand U430 (N_430,In_689,In_934);
or U431 (N_431,In_915,In_8);
and U432 (N_432,In_432,In_910);
xor U433 (N_433,In_1565,In_2281);
nand U434 (N_434,In_410,In_1164);
nand U435 (N_435,In_329,In_2297);
and U436 (N_436,In_1309,In_2362);
and U437 (N_437,In_867,In_2223);
or U438 (N_438,In_207,In_2119);
xnor U439 (N_439,In_274,In_879);
and U440 (N_440,In_1907,In_216);
nand U441 (N_441,In_326,In_1941);
nor U442 (N_442,In_780,In_2180);
nor U443 (N_443,In_1058,In_1380);
and U444 (N_444,In_716,In_1492);
nor U445 (N_445,In_596,In_574);
and U446 (N_446,In_1969,In_970);
nor U447 (N_447,In_989,In_1378);
or U448 (N_448,In_465,In_1614);
and U449 (N_449,In_993,In_2426);
and U450 (N_450,In_420,In_2232);
nor U451 (N_451,In_84,In_1439);
nand U452 (N_452,In_13,In_211);
nand U453 (N_453,In_1152,In_982);
nor U454 (N_454,In_766,In_1206);
nand U455 (N_455,In_1976,In_1517);
and U456 (N_456,In_2244,In_1448);
xor U457 (N_457,In_1610,In_610);
nand U458 (N_458,In_425,In_947);
nor U459 (N_459,In_698,In_193);
xnor U460 (N_460,In_202,In_2336);
or U461 (N_461,In_1238,In_1953);
nor U462 (N_462,In_1817,In_373);
or U463 (N_463,In_2353,In_739);
and U464 (N_464,In_764,In_1174);
nand U465 (N_465,In_276,In_767);
or U466 (N_466,In_1165,In_1591);
nor U467 (N_467,In_1315,In_19);
or U468 (N_468,In_352,In_1768);
or U469 (N_469,In_996,In_963);
xor U470 (N_470,In_1363,In_902);
and U471 (N_471,In_2396,In_617);
or U472 (N_472,In_755,In_429);
nor U473 (N_473,In_126,In_663);
and U474 (N_474,In_2282,In_1387);
nor U475 (N_475,In_995,In_442);
nand U476 (N_476,In_320,In_1386);
or U477 (N_477,In_1245,In_155);
nor U478 (N_478,In_1305,In_2254);
or U479 (N_479,In_1267,In_240);
or U480 (N_480,In_254,In_1431);
xor U481 (N_481,In_1114,In_1280);
nand U482 (N_482,In_1870,In_1936);
and U483 (N_483,In_1954,In_2041);
nor U484 (N_484,In_1345,In_1493);
xnor U485 (N_485,In_969,In_1056);
nand U486 (N_486,In_2144,In_271);
xnor U487 (N_487,In_1690,In_2403);
and U488 (N_488,In_2296,In_754);
and U489 (N_489,In_477,In_1593);
nor U490 (N_490,In_397,In_677);
and U491 (N_491,In_2416,In_964);
xnor U492 (N_492,In_884,In_1762);
or U493 (N_493,In_2060,In_784);
nor U494 (N_494,In_680,In_1042);
xnor U495 (N_495,In_1093,In_980);
and U496 (N_496,In_1618,In_2031);
or U497 (N_497,In_2375,In_1107);
xnor U498 (N_498,In_449,In_2179);
and U499 (N_499,In_1539,In_940);
nor U500 (N_500,In_942,In_877);
xnor U501 (N_501,In_5,In_837);
or U502 (N_502,In_2173,In_444);
xnor U503 (N_503,In_458,In_1963);
nand U504 (N_504,In_2465,In_917);
and U505 (N_505,In_1189,In_348);
and U506 (N_506,In_1928,In_1021);
and U507 (N_507,In_961,In_1156);
nand U508 (N_508,In_2483,In_1179);
nor U509 (N_509,In_296,In_547);
xor U510 (N_510,In_1242,In_377);
nor U511 (N_511,In_423,In_1927);
nor U512 (N_512,In_540,In_1915);
nor U513 (N_513,In_1526,In_2040);
nand U514 (N_514,In_1236,In_1360);
nor U515 (N_515,In_992,In_455);
nor U516 (N_516,In_738,In_554);
and U517 (N_517,In_887,In_2457);
or U518 (N_518,In_1002,In_1949);
xor U519 (N_519,In_349,In_1758);
xor U520 (N_520,In_82,In_86);
or U521 (N_521,In_2196,In_1397);
nand U522 (N_522,In_286,In_896);
nor U523 (N_523,In_249,In_1856);
and U524 (N_524,In_1793,In_1602);
xor U525 (N_525,In_2105,In_1086);
nand U526 (N_526,In_1173,In_514);
or U527 (N_527,In_21,In_682);
xnor U528 (N_528,In_1701,In_703);
nor U529 (N_529,In_1133,In_700);
or U530 (N_530,In_2096,In_869);
xor U531 (N_531,In_1653,In_2312);
or U532 (N_532,In_690,In_2246);
or U533 (N_533,In_548,In_1727);
xor U534 (N_534,In_2266,In_600);
nor U535 (N_535,In_187,In_1211);
and U536 (N_536,In_1628,In_400);
xor U537 (N_537,In_1213,In_632);
and U538 (N_538,In_987,In_1119);
or U539 (N_539,In_2363,In_618);
or U540 (N_540,In_1715,In_893);
and U541 (N_541,In_1918,In_2272);
nor U542 (N_542,In_1005,In_1136);
or U543 (N_543,In_1188,In_687);
or U544 (N_544,In_2186,In_2418);
nor U545 (N_545,In_180,In_706);
or U546 (N_546,In_543,In_2032);
xnor U547 (N_547,In_1705,In_538);
or U548 (N_548,In_750,In_732);
or U549 (N_549,In_1271,In_1795);
or U550 (N_550,In_1349,In_158);
nor U551 (N_551,In_53,In_1412);
xor U552 (N_552,In_10,In_956);
and U553 (N_553,In_44,In_403);
xnor U554 (N_554,In_1746,In_2112);
nor U555 (N_555,In_1589,In_230);
or U556 (N_556,In_106,In_1446);
or U557 (N_557,In_1744,In_338);
or U558 (N_558,In_2037,In_2298);
xnor U559 (N_559,In_613,In_1680);
xnor U560 (N_560,In_1942,In_54);
or U561 (N_561,In_2054,In_312);
nor U562 (N_562,In_1613,In_1926);
nor U563 (N_563,In_1023,In_777);
and U564 (N_564,In_2326,In_2084);
nor U565 (N_565,In_1512,In_2439);
xor U566 (N_566,In_772,In_124);
and U567 (N_567,In_197,In_313);
or U568 (N_568,In_787,In_238);
xnor U569 (N_569,In_1862,In_1203);
nand U570 (N_570,In_2389,In_771);
or U571 (N_571,In_1204,In_1453);
or U572 (N_572,In_1452,In_791);
xnor U573 (N_573,In_175,In_2415);
nand U574 (N_574,In_1377,In_438);
and U575 (N_575,In_1913,In_321);
nor U576 (N_576,In_2434,In_1708);
and U577 (N_577,In_422,In_2220);
nand U578 (N_578,In_2149,In_795);
nand U579 (N_579,In_288,In_1728);
and U580 (N_580,In_2264,In_2175);
nor U581 (N_581,In_2121,In_196);
nor U582 (N_582,In_559,In_656);
xor U583 (N_583,In_2493,In_368);
nor U584 (N_584,In_1047,In_1458);
nor U585 (N_585,In_233,In_38);
and U586 (N_586,In_926,In_2350);
and U587 (N_587,In_1413,In_597);
or U588 (N_588,In_361,In_1624);
or U589 (N_589,In_2065,In_1876);
and U590 (N_590,In_2168,In_1457);
nand U591 (N_591,In_388,In_2092);
nand U592 (N_592,In_1122,In_253);
nand U593 (N_593,In_1534,In_404);
xnor U594 (N_594,In_1720,In_1898);
or U595 (N_595,In_2329,In_57);
xor U596 (N_596,In_1273,In_289);
xnor U597 (N_597,In_1767,In_2262);
xnor U598 (N_598,In_2427,In_1930);
xnor U599 (N_599,In_2079,In_1864);
or U600 (N_600,In_566,In_905);
and U601 (N_601,In_2044,In_1487);
or U602 (N_602,In_11,In_1632);
xnor U603 (N_603,In_1513,In_1620);
nor U604 (N_604,In_346,In_2019);
nand U605 (N_605,In_255,In_608);
or U606 (N_606,In_788,In_105);
or U607 (N_607,In_453,In_2057);
nand U608 (N_608,In_371,In_1061);
nand U609 (N_609,In_515,In_1776);
xnor U610 (N_610,In_1040,In_512);
or U611 (N_611,In_2428,In_2279);
nor U612 (N_612,In_878,In_2306);
xnor U613 (N_613,In_1825,In_150);
or U614 (N_614,In_2122,In_1474);
nor U615 (N_615,In_1835,In_415);
or U616 (N_616,In_1967,In_2348);
nor U617 (N_617,In_1576,In_2345);
or U618 (N_618,In_152,In_670);
xnor U619 (N_619,In_1753,In_2157);
xor U620 (N_620,In_2291,In_1194);
and U621 (N_621,In_2429,In_1094);
xnor U622 (N_622,In_1106,In_1064);
nor U623 (N_623,In_102,In_591);
nor U624 (N_624,In_1027,In_2072);
nor U625 (N_625,In_2205,In_1147);
and U626 (N_626,In_616,In_331);
nand U627 (N_627,In_683,In_1088);
nand U628 (N_628,In_1562,In_733);
xnor U629 (N_629,In_1950,In_131);
and U630 (N_630,In_121,In_1833);
nor U631 (N_631,In_1199,In_1742);
nand U632 (N_632,In_1914,In_546);
nor U633 (N_633,In_955,In_594);
or U634 (N_634,In_2001,In_1307);
nor U635 (N_635,In_1703,In_1134);
or U636 (N_636,In_1153,In_1376);
nand U637 (N_637,In_146,In_1224);
nor U638 (N_638,In_357,In_2474);
xnor U639 (N_639,In_2288,In_1831);
xor U640 (N_640,In_2384,In_2161);
nor U641 (N_641,In_1186,In_1365);
and U642 (N_642,In_1454,In_2421);
nor U643 (N_643,In_1281,In_2463);
nand U644 (N_644,In_142,In_1732);
xnor U645 (N_645,In_2269,In_1344);
xnor U646 (N_646,In_2165,In_704);
xnor U647 (N_647,In_149,In_1749);
or U648 (N_648,In_668,In_306);
or U649 (N_649,In_2317,In_601);
or U650 (N_650,In_1988,In_2327);
nand U651 (N_651,In_938,In_1011);
and U652 (N_652,In_768,In_2351);
xor U653 (N_653,In_385,In_430);
xnor U654 (N_654,In_695,In_24);
nand U655 (N_655,In_1193,In_476);
xnor U656 (N_656,In_1196,In_406);
nand U657 (N_657,In_318,In_2480);
xnor U658 (N_658,In_447,In_1895);
nor U659 (N_659,In_2460,In_1679);
nor U660 (N_660,In_773,In_1975);
xor U661 (N_661,In_139,In_2245);
and U662 (N_662,In_340,In_2095);
and U663 (N_663,In_516,In_526);
nor U664 (N_664,In_1404,In_2497);
or U665 (N_665,In_524,In_2388);
nor U666 (N_666,In_907,In_1223);
nor U667 (N_667,In_1356,In_3);
or U668 (N_668,In_1081,In_154);
nor U669 (N_669,In_483,In_2393);
nor U670 (N_670,In_1172,In_1666);
and U671 (N_671,In_43,In_1577);
xor U672 (N_672,In_2402,In_1547);
nand U673 (N_673,In_60,In_838);
or U674 (N_674,In_756,In_860);
nand U675 (N_675,In_1798,In_1844);
nor U676 (N_676,In_1144,In_2354);
xor U677 (N_677,In_300,In_1989);
or U678 (N_678,In_2077,In_1085);
nand U679 (N_679,In_470,In_1573);
and U680 (N_680,In_229,In_626);
or U681 (N_681,In_2140,In_103);
or U682 (N_682,In_1274,In_1638);
nor U683 (N_683,In_1105,In_2381);
or U684 (N_684,In_2451,In_874);
nand U685 (N_685,In_2035,In_185);
xnor U686 (N_686,In_2125,In_358);
or U687 (N_687,In_892,In_448);
xnor U688 (N_688,In_2466,In_1659);
and U689 (N_689,In_199,In_1665);
or U690 (N_690,In_92,In_931);
nand U691 (N_691,In_2316,In_2231);
or U692 (N_692,In_1117,In_1456);
xnor U693 (N_693,In_1588,In_1766);
nand U694 (N_694,In_604,In_1264);
xnor U695 (N_695,In_1559,In_174);
xor U696 (N_696,In_2301,In_1871);
or U697 (N_697,In_2471,In_1478);
xor U698 (N_698,In_1555,In_749);
or U699 (N_699,In_1903,In_2141);
nand U700 (N_700,In_1251,In_364);
nand U701 (N_701,In_1799,In_1961);
xor U702 (N_702,In_2423,In_835);
and U703 (N_703,In_1910,In_2367);
or U704 (N_704,In_73,In_997);
xor U705 (N_705,In_804,In_1151);
and U706 (N_706,In_1982,In_2219);
or U707 (N_707,In_2225,In_1531);
nor U708 (N_708,In_1719,In_1609);
nand U709 (N_709,In_1060,In_1022);
nor U710 (N_710,In_1494,In_1007);
nand U711 (N_711,In_533,In_1254);
and U712 (N_712,In_737,In_2158);
xor U713 (N_713,In_2048,In_912);
nor U714 (N_714,In_61,In_570);
or U715 (N_715,In_1006,In_1464);
and U716 (N_716,In_622,In_440);
and U717 (N_717,In_1250,In_250);
nor U718 (N_718,In_1483,In_953);
nor U719 (N_719,In_1284,In_932);
and U720 (N_720,In_1462,In_1880);
or U721 (N_721,In_2009,In_2478);
and U722 (N_722,In_789,In_1511);
nand U723 (N_723,In_424,In_1540);
xor U724 (N_724,In_2285,In_519);
and U725 (N_725,In_1244,In_1230);
nand U726 (N_726,In_684,In_2496);
nor U727 (N_727,In_1771,In_1740);
xor U728 (N_728,In_888,In_1594);
or U729 (N_729,In_1841,In_653);
or U730 (N_730,In_22,In_2365);
and U731 (N_731,In_1760,In_1997);
nand U732 (N_732,In_1597,In_589);
nand U733 (N_733,In_1383,In_2069);
or U734 (N_734,In_986,In_181);
or U735 (N_735,In_1418,In_138);
and U736 (N_736,In_1630,In_2431);
nor U737 (N_737,In_2400,In_1716);
nor U738 (N_738,In_1438,In_2159);
nand U739 (N_739,In_381,In_87);
nor U740 (N_740,In_1480,In_1479);
or U741 (N_741,In_984,In_208);
and U742 (N_742,In_1737,In_1977);
nand U743 (N_743,In_218,In_369);
xnor U744 (N_744,In_975,In_134);
and U745 (N_745,In_1468,In_1260);
or U746 (N_746,In_1459,In_1984);
and U747 (N_747,In_2408,In_794);
xnor U748 (N_748,In_2374,In_1176);
or U749 (N_749,In_2444,In_1026);
xnor U750 (N_750,In_1031,In_1567);
xnor U751 (N_751,In_778,In_1670);
nand U752 (N_752,In_2172,In_1057);
or U753 (N_753,In_479,In_1482);
xor U754 (N_754,In_40,In_267);
and U755 (N_755,In_341,In_1673);
or U756 (N_756,In_281,In_1587);
and U757 (N_757,In_1606,In_659);
nand U758 (N_758,In_678,In_59);
nand U759 (N_759,In_945,In_943);
xor U760 (N_760,In_1445,In_1168);
nand U761 (N_761,In_2053,In_2425);
and U762 (N_762,In_502,In_1372);
xor U763 (N_763,In_446,In_2227);
or U764 (N_764,In_1652,In_1797);
or U765 (N_765,In_262,In_251);
or U766 (N_766,In_2171,In_828);
and U767 (N_767,In_885,In_2107);
and U768 (N_768,In_2433,In_508);
or U769 (N_769,In_2436,In_2017);
and U770 (N_770,In_119,In_457);
nor U771 (N_771,In_2499,In_1622);
or U772 (N_772,In_2368,In_459);
and U773 (N_773,In_2422,In_1854);
nand U774 (N_774,In_648,In_1310);
nor U775 (N_775,In_223,In_1089);
and U776 (N_776,In_1787,In_190);
nand U777 (N_777,In_582,In_1973);
xor U778 (N_778,In_2003,In_717);
nor U779 (N_779,In_1840,In_725);
and U780 (N_780,In_2242,In_779);
xnor U781 (N_781,In_1217,In_1009);
and U782 (N_782,In_1124,In_1148);
xor U783 (N_783,In_693,In_1050);
or U784 (N_784,In_1912,In_715);
and U785 (N_785,In_831,In_839);
xor U786 (N_786,In_1450,In_64);
or U787 (N_787,In_843,In_2222);
and U788 (N_788,In_268,In_322);
nor U789 (N_789,In_595,In_1321);
or U790 (N_790,In_1306,In_1808);
or U791 (N_791,In_769,In_661);
or U792 (N_792,In_614,In_2358);
nor U793 (N_793,In_2250,In_1278);
nand U794 (N_794,In_1929,In_935);
or U795 (N_795,In_2409,In_356);
and U796 (N_796,In_1177,In_832);
nor U797 (N_797,In_2114,In_1645);
nand U798 (N_798,In_1013,In_1351);
nand U799 (N_799,In_2461,In_1080);
nand U800 (N_800,In_232,In_2359);
nor U801 (N_801,In_2498,In_1848);
nand U802 (N_802,In_56,In_2152);
or U803 (N_803,In_2314,In_1545);
and U804 (N_804,In_2174,In_2305);
or U805 (N_805,In_1788,In_634);
or U806 (N_806,In_285,In_658);
nand U807 (N_807,In_2090,In_173);
nand U808 (N_808,In_864,In_669);
xnor U809 (N_809,In_1779,In_1761);
xnor U810 (N_810,In_1205,In_765);
nand U811 (N_811,In_2027,In_2332);
nand U812 (N_812,In_643,In_1399);
nor U813 (N_813,In_665,In_1391);
nor U814 (N_814,In_2464,In_999);
xnor U815 (N_815,In_2338,In_1764);
or U816 (N_816,In_748,In_1460);
xor U817 (N_817,In_2070,In_861);
nand U818 (N_818,In_1676,In_71);
or U819 (N_819,In_1395,In_2155);
xor U820 (N_820,In_2030,In_2278);
and U821 (N_821,In_959,In_405);
or U822 (N_822,In_228,In_1486);
xnor U823 (N_823,In_2043,In_1693);
nor U824 (N_824,In_1560,In_801);
nor U825 (N_825,In_2148,In_911);
and U826 (N_826,In_2007,In_1166);
nand U827 (N_827,In_1743,In_581);
nand U828 (N_828,In_609,In_51);
or U829 (N_829,In_1381,In_873);
xnor U830 (N_830,In_1077,In_1481);
or U831 (N_831,In_402,In_337);
nand U832 (N_832,In_46,In_1099);
xnor U833 (N_833,In_1028,In_899);
or U834 (N_834,In_611,In_2202);
and U835 (N_835,In_521,In_1065);
xor U836 (N_836,In_182,In_290);
xor U837 (N_837,In_2189,In_950);
nor U838 (N_838,In_49,In_1877);
nand U839 (N_839,In_1803,In_612);
nor U840 (N_840,In_1585,In_231);
and U841 (N_841,In_1215,In_1893);
nand U842 (N_842,In_1874,In_148);
nand U843 (N_843,In_560,In_1410);
nand U844 (N_844,In_2286,In_380);
or U845 (N_845,In_2194,In_1937);
xnor U846 (N_846,In_1187,In_1463);
or U847 (N_847,In_1255,In_1945);
and U848 (N_848,In_2300,In_67);
or U849 (N_849,In_850,In_1966);
xnor U850 (N_850,In_641,In_1126);
and U851 (N_851,In_637,In_949);
or U852 (N_852,In_1987,In_1546);
or U853 (N_853,In_1066,In_836);
or U854 (N_854,In_219,In_1625);
nand U855 (N_855,In_345,In_1634);
nand U856 (N_856,In_2132,In_2364);
nor U857 (N_857,In_2081,In_1865);
xor U858 (N_858,In_751,In_1277);
or U859 (N_859,In_1029,In_2154);
and U860 (N_860,In_1890,In_1227);
and U861 (N_861,In_1155,In_1426);
nor U862 (N_862,In_1461,In_1601);
and U863 (N_863,In_2342,In_2120);
nor U864 (N_864,In_2488,In_1350);
xnor U865 (N_865,In_1872,In_580);
or U866 (N_866,In_2265,In_1688);
xor U867 (N_867,In_1866,In_2162);
and U868 (N_868,In_492,In_1330);
nor U869 (N_869,In_2209,In_1295);
or U870 (N_870,In_1125,In_812);
xnor U871 (N_871,In_536,In_1072);
or U872 (N_872,In_1706,In_2218);
nand U873 (N_873,In_2331,In_1911);
xor U874 (N_874,In_460,In_1739);
xnor U875 (N_875,In_2038,In_1617);
nand U876 (N_876,In_829,In_1012);
nand U877 (N_877,In_1017,In_511);
xnor U878 (N_878,In_2414,In_891);
xnor U879 (N_879,In_1123,In_2136);
or U880 (N_880,In_1698,In_147);
nand U881 (N_881,In_212,In_621);
xor U882 (N_882,In_545,In_1411);
xnor U883 (N_883,In_1102,In_441);
nand U884 (N_884,In_34,In_2419);
nand U885 (N_885,In_189,In_1885);
xnor U886 (N_886,In_118,In_382);
nand U887 (N_887,In_1180,In_15);
and U888 (N_888,In_2050,In_561);
nand U889 (N_889,In_660,In_130);
and U890 (N_890,In_1675,In_1101);
and U891 (N_891,In_1702,In_1256);
xor U892 (N_892,In_217,In_876);
nand U893 (N_893,In_499,In_1552);
and U894 (N_894,In_1207,In_1396);
or U895 (N_895,In_1275,In_1682);
and U896 (N_896,In_2452,In_192);
or U897 (N_897,In_1685,In_957);
xnor U898 (N_898,In_1018,In_1775);
nor U899 (N_899,In_1978,In_1524);
or U900 (N_900,In_1851,In_859);
or U901 (N_901,In_2410,In_688);
or U902 (N_902,In_1276,In_567);
nand U903 (N_903,In_1908,In_2163);
or U904 (N_904,In_528,In_1408);
nor U905 (N_905,In_108,In_631);
and U906 (N_906,In_2052,In_2164);
nand U907 (N_907,In_122,In_1818);
nor U908 (N_908,In_2318,In_1405);
nor U909 (N_909,In_1981,In_916);
xor U910 (N_910,In_646,In_1730);
or U911 (N_911,In_1096,In_1806);
nor U912 (N_912,In_2267,In_2462);
and U913 (N_913,In_169,In_1707);
or U914 (N_914,In_991,In_454);
xor U915 (N_915,In_2045,In_227);
nand U916 (N_916,In_506,In_1074);
nand U917 (N_917,In_1972,In_640);
xnor U918 (N_918,In_1249,In_307);
xnor U919 (N_919,In_143,In_1691);
and U920 (N_920,In_2061,In_2073);
nand U921 (N_921,In_1343,In_988);
nor U922 (N_922,In_2190,In_1530);
nand U923 (N_923,In_2287,In_542);
xnor U924 (N_924,In_858,In_853);
nor U925 (N_925,In_2442,In_844);
xnor U926 (N_926,In_1332,In_493);
nor U927 (N_927,In_2277,In_785);
nand U928 (N_928,In_625,In_1298);
nor U929 (N_929,In_2274,In_145);
or U930 (N_930,In_201,In_1810);
and U931 (N_931,In_735,In_1);
nand U932 (N_932,In_2283,In_1045);
and U933 (N_933,In_1657,In_712);
or U934 (N_934,In_2324,In_1644);
nand U935 (N_935,In_376,In_870);
xnor U936 (N_936,In_742,In_1212);
nand U937 (N_937,In_944,In_897);
nor U938 (N_938,In_909,In_500);
nor U939 (N_939,In_2109,In_52);
and U940 (N_940,In_951,In_2494);
or U941 (N_941,In_2407,In_186);
xor U942 (N_942,In_1347,In_29);
nand U943 (N_943,In_1466,In_854);
xnor U944 (N_944,In_2236,In_1198);
nand U945 (N_945,In_1030,In_1209);
nor U946 (N_946,In_807,In_1523);
xnor U947 (N_947,In_623,In_672);
nor U948 (N_948,In_2349,In_1650);
xor U949 (N_949,In_36,In_913);
and U950 (N_950,In_2124,In_319);
xor U951 (N_951,In_1157,In_2151);
xor U952 (N_952,In_1741,In_523);
and U953 (N_953,In_518,In_362);
xor U954 (N_954,In_845,In_1353);
nand U955 (N_955,In_2127,In_1643);
nand U956 (N_956,In_936,In_1140);
xor U957 (N_957,In_2200,In_2413);
nor U958 (N_958,In_1154,In_1403);
xor U959 (N_959,In_1161,In_1004);
nor U960 (N_960,In_830,In_707);
and U961 (N_961,In_1142,In_1564);
nor U962 (N_962,In_701,In_923);
nand U963 (N_963,In_796,In_1538);
and U964 (N_964,In_1784,In_2401);
xnor U965 (N_965,In_1578,In_191);
nor U966 (N_966,In_2028,In_383);
and U967 (N_967,In_1781,In_1430);
xnor U968 (N_968,In_1956,In_711);
and U969 (N_969,In_480,In_740);
nand U970 (N_970,In_889,In_1686);
nor U971 (N_971,In_163,In_1964);
or U972 (N_972,In_2392,In_1406);
or U973 (N_973,In_1084,In_1892);
or U974 (N_974,In_1700,In_1660);
and U975 (N_975,In_162,In_474);
nor U976 (N_976,In_568,In_234);
and U977 (N_977,In_2437,In_2490);
xnor U978 (N_978,In_852,In_809);
xnor U979 (N_979,In_153,In_1335);
or U980 (N_980,In_2492,In_1175);
xor U981 (N_981,In_1759,In_775);
and U982 (N_982,In_2101,In_1394);
xor U983 (N_983,In_1473,In_1651);
nand U984 (N_984,In_930,In_1233);
nor U985 (N_985,In_101,In_747);
nand U986 (N_986,In_1128,In_1946);
or U987 (N_987,In_2063,In_395);
xnor U988 (N_988,In_392,In_2023);
xnor U989 (N_989,In_1639,In_977);
or U990 (N_990,In_2487,In_1756);
nand U991 (N_991,In_1931,In_1626);
xor U992 (N_992,In_1092,In_1098);
xnor U993 (N_993,In_42,In_2055);
nor U994 (N_994,In_1519,In_1358);
nand U995 (N_995,In_2056,In_2192);
nor U996 (N_996,In_541,In_1292);
and U997 (N_997,In_2138,In_2184);
nand U998 (N_998,In_1127,In_2346);
and U999 (N_999,In_1049,In_2399);
nor U1000 (N_1000,In_606,N_726);
nand U1001 (N_1001,N_36,In_1805);
nand U1002 (N_1002,In_370,N_931);
nor U1003 (N_1003,N_607,N_725);
nand U1004 (N_1004,N_754,In_363);
nor U1005 (N_1005,N_265,In_586);
or U1006 (N_1006,N_997,N_988);
or U1007 (N_1007,In_282,N_278);
xnor U1008 (N_1008,In_244,In_2432);
and U1009 (N_1009,N_955,N_378);
and U1010 (N_1010,N_81,In_1541);
and U1011 (N_1011,N_78,In_676);
nor U1012 (N_1012,In_1476,N_695);
or U1013 (N_1013,N_355,N_461);
nor U1014 (N_1014,N_912,In_1171);
nand U1015 (N_1015,N_519,In_760);
and U1016 (N_1016,In_2356,In_127);
and U1017 (N_1017,In_2086,In_2113);
nand U1018 (N_1018,In_2446,N_432);
nor U1019 (N_1019,N_382,N_350);
nand U1020 (N_1020,N_923,In_800);
and U1021 (N_1021,N_753,N_788);
and U1022 (N_1022,In_273,N_268);
and U1023 (N_1023,N_174,In_1389);
nor U1024 (N_1024,In_1316,N_744);
xnor U1025 (N_1025,N_608,N_430);
and U1026 (N_1026,N_780,N_264);
nand U1027 (N_1027,N_48,N_802);
or U1028 (N_1028,N_653,N_814);
nand U1029 (N_1029,In_2074,In_387);
xnor U1030 (N_1030,In_2150,N_858);
nor U1031 (N_1031,In_1867,N_253);
nor U1032 (N_1032,N_499,N_67);
nor U1033 (N_1033,In_2481,N_700);
and U1034 (N_1034,N_406,N_141);
xnor U1035 (N_1035,N_470,N_513);
or U1036 (N_1036,N_76,In_120);
nor U1037 (N_1037,N_170,N_344);
and U1038 (N_1038,N_976,N_839);
xor U1039 (N_1039,N_11,In_1504);
nor U1040 (N_1040,N_903,In_2147);
nand U1041 (N_1041,In_236,In_2131);
xor U1042 (N_1042,N_301,N_226);
or U1043 (N_1043,In_1407,N_71);
nor U1044 (N_1044,N_148,In_2207);
or U1045 (N_1045,N_186,N_7);
and U1046 (N_1046,N_175,N_545);
nor U1047 (N_1047,N_291,N_940);
nor U1048 (N_1048,N_273,N_512);
and U1049 (N_1049,N_20,N_855);
and U1050 (N_1050,N_866,In_426);
or U1051 (N_1051,In_1268,In_965);
xor U1052 (N_1052,N_690,In_72);
and U1053 (N_1053,In_351,In_1962);
nor U1054 (N_1054,N_567,In_1182);
and U1055 (N_1055,N_999,In_1120);
or U1056 (N_1056,In_1048,N_290);
xnor U1057 (N_1057,In_165,In_343);
nand U1058 (N_1058,N_763,N_692);
or U1059 (N_1059,N_591,In_1571);
nor U1060 (N_1060,In_1433,N_688);
nor U1061 (N_1061,In_2459,N_42);
nor U1062 (N_1062,In_633,N_303);
or U1063 (N_1063,In_248,In_1542);
and U1064 (N_1064,N_901,In_436);
nand U1065 (N_1065,N_498,N_257);
nand U1066 (N_1066,N_585,In_2361);
nor U1067 (N_1067,N_408,N_241);
and U1068 (N_1068,In_1159,N_338);
nand U1069 (N_1069,In_862,N_463);
xor U1070 (N_1070,N_404,N_849);
xnor U1071 (N_1071,In_2080,N_467);
nor U1072 (N_1072,N_589,N_906);
nand U1073 (N_1073,N_320,N_670);
nor U1074 (N_1074,In_1070,N_828);
xor U1075 (N_1075,In_579,N_511);
nor U1076 (N_1076,N_555,N_920);
nor U1077 (N_1077,N_678,N_626);
or U1078 (N_1078,In_1736,In_808);
nor U1079 (N_1079,N_559,N_165);
and U1080 (N_1080,N_538,N_423);
and U1081 (N_1081,In_1025,In_629);
or U1082 (N_1082,N_902,In_1416);
xor U1083 (N_1083,N_407,N_297);
and U1084 (N_1084,N_554,N_664);
nand U1085 (N_1085,N_987,In_639);
or U1086 (N_1086,N_549,N_529);
and U1087 (N_1087,N_333,N_618);
or U1088 (N_1088,N_518,N_40);
nand U1089 (N_1089,N_772,In_27);
xor U1090 (N_1090,N_939,In_317);
nand U1091 (N_1091,N_479,In_2370);
nand U1092 (N_1092,N_65,N_198);
or U1093 (N_1093,N_733,N_287);
nand U1094 (N_1094,N_703,N_525);
nand U1095 (N_1095,In_1020,N_422);
nand U1096 (N_1096,In_116,N_17);
and U1097 (N_1097,N_638,N_23);
or U1098 (N_1098,N_497,In_588);
nand U1099 (N_1099,In_1008,In_1270);
nor U1100 (N_1100,N_798,In_41);
xor U1101 (N_1101,N_601,In_1037);
nand U1102 (N_1102,N_140,N_481);
nand U1103 (N_1103,N_602,N_911);
and U1104 (N_1104,N_950,In_2438);
nor U1105 (N_1105,N_280,N_717);
or U1106 (N_1106,N_654,N_623);
or U1107 (N_1107,In_1822,N_645);
nand U1108 (N_1108,N_635,In_1243);
xor U1109 (N_1109,N_220,N_379);
or U1110 (N_1110,In_1580,In_1558);
or U1111 (N_1111,N_180,N_155);
nor U1112 (N_1112,N_409,N_878);
xnor U1113 (N_1113,N_205,In_2064);
nor U1114 (N_1114,N_677,In_2337);
nand U1115 (N_1115,N_732,In_308);
or U1116 (N_1116,N_989,N_55);
nor U1117 (N_1117,N_310,N_620);
nor U1118 (N_1118,N_416,In_1210);
and U1119 (N_1119,In_295,In_1130);
nand U1120 (N_1120,N_399,N_385);
or U1121 (N_1121,In_1200,N_557);
nor U1122 (N_1122,N_254,In_2472);
nand U1123 (N_1123,In_302,N_977);
or U1124 (N_1124,N_46,In_1983);
or U1125 (N_1125,N_526,N_351);
nand U1126 (N_1126,N_769,N_122);
and U1127 (N_1127,In_619,N_248);
xnor U1128 (N_1128,In_354,N_262);
nor U1129 (N_1129,N_613,In_298);
nor U1130 (N_1130,N_246,In_1178);
xnor U1131 (N_1131,N_390,N_521);
or U1132 (N_1132,In_272,N_172);
and U1133 (N_1133,N_578,N_427);
and U1134 (N_1134,In_1340,In_1279);
and U1135 (N_1135,In_194,N_60);
or U1136 (N_1136,In_287,N_848);
nand U1137 (N_1137,In_1181,N_736);
nor U1138 (N_1138,N_547,N_292);
nor U1139 (N_1139,In_90,N_507);
nor U1140 (N_1140,In_1327,N_985);
or U1141 (N_1141,In_531,N_777);
xor U1142 (N_1142,N_966,In_1313);
nor U1143 (N_1143,N_505,N_307);
xnor U1144 (N_1144,N_656,N_742);
nand U1145 (N_1145,N_84,N_816);
or U1146 (N_1146,In_1282,N_861);
nand U1147 (N_1147,N_238,In_1283);
nor U1148 (N_1148,N_799,In_1318);
and U1149 (N_1149,N_15,In_2034);
or U1150 (N_1150,In_645,N_504);
and U1151 (N_1151,In_1422,N_918);
and U1152 (N_1152,In_35,N_450);
and U1153 (N_1153,In_1046,N_541);
nor U1154 (N_1154,In_1544,N_395);
nand U1155 (N_1155,N_293,N_203);
xor U1156 (N_1156,In_525,N_774);
nand U1157 (N_1157,In_1879,In_1222);
and U1158 (N_1158,N_373,In_585);
or U1159 (N_1159,N_820,N_856);
nand U1160 (N_1160,In_1932,In_2309);
xor U1161 (N_1161,In_280,N_953);
and U1162 (N_1162,N_157,In_552);
and U1163 (N_1163,N_756,In_2243);
xnor U1164 (N_1164,N_580,N_197);
and U1165 (N_1165,N_927,In_496);
xnor U1166 (N_1166,In_894,N_701);
and U1167 (N_1167,In_976,N_974);
or U1168 (N_1168,N_94,N_967);
nand U1169 (N_1169,In_578,N_779);
nor U1170 (N_1170,In_260,N_947);
nand U1171 (N_1171,N_694,N_489);
nor U1172 (N_1172,N_956,N_456);
xor U1173 (N_1173,N_926,N_5);
nor U1174 (N_1174,N_764,In_96);
nand U1175 (N_1175,N_508,N_524);
and U1176 (N_1176,In_1820,N_888);
or U1177 (N_1177,N_149,In_156);
and U1178 (N_1178,N_363,N_343);
or U1179 (N_1179,N_302,N_169);
nor U1180 (N_1180,N_136,In_94);
nor U1181 (N_1181,In_537,In_1253);
or U1182 (N_1182,N_739,In_1162);
or U1183 (N_1183,In_1755,N_884);
xor U1184 (N_1184,In_20,N_551);
or U1185 (N_1185,In_718,In_1869);
or U1186 (N_1186,In_1231,N_396);
nor U1187 (N_1187,N_29,N_542);
nor U1188 (N_1188,N_864,N_641);
nor U1189 (N_1189,N_550,In_1362);
and U1190 (N_1190,N_766,N_791);
nand U1191 (N_1191,N_817,N_924);
nand U1192 (N_1192,In_1980,In_2275);
nor U1193 (N_1193,N_26,In_1947);
or U1194 (N_1194,N_397,In_2191);
and U1195 (N_1195,N_69,N_188);
or U1196 (N_1196,N_546,In_1038);
xor U1197 (N_1197,N_611,N_698);
or U1198 (N_1198,In_1218,N_123);
and U1199 (N_1199,N_332,N_628);
and U1200 (N_1200,N_318,N_672);
nor U1201 (N_1201,N_914,N_812);
nor U1202 (N_1202,N_222,N_862);
nand U1203 (N_1203,N_709,In_336);
xor U1204 (N_1204,N_921,N_109);
xnor U1205 (N_1205,In_1141,N_185);
nand U1206 (N_1206,N_457,In_636);
nand U1207 (N_1207,In_399,N_161);
xnor U1208 (N_1208,N_646,N_274);
nand U1209 (N_1209,N_433,N_751);
nor U1210 (N_1210,In_2253,N_792);
nand U1211 (N_1211,N_894,N_621);
nand U1212 (N_1212,N_622,N_9);
xnor U1213 (N_1213,N_88,In_904);
and U1214 (N_1214,N_680,In_1323);
and U1215 (N_1215,In_310,N_119);
and U1216 (N_1216,N_104,N_305);
or U1217 (N_1217,N_412,In_469);
xor U1218 (N_1218,N_349,N_356);
nor U1219 (N_1219,N_420,N_937);
or U1220 (N_1220,In_1883,N_583);
and U1221 (N_1221,In_1605,N_684);
nand U1222 (N_1222,N_948,N_70);
and U1223 (N_1223,N_929,In_1000);
nor U1224 (N_1224,N_146,In_80);
and U1225 (N_1225,N_539,In_1704);
or U1226 (N_1226,N_340,N_581);
nor U1227 (N_1227,N_886,N_676);
and U1228 (N_1228,In_503,N_568);
nor U1229 (N_1229,N_905,N_750);
nand U1230 (N_1230,In_37,In_1763);
xnor U1231 (N_1231,N_277,N_604);
xor U1232 (N_1232,In_1968,In_753);
nand U1233 (N_1233,N_35,In_1993);
xor U1234 (N_1234,N_32,In_900);
nor U1235 (N_1235,N_990,N_114);
or U1236 (N_1236,N_522,In_2477);
and U1237 (N_1237,N_139,N_770);
or U1238 (N_1238,N_58,In_421);
xor U1239 (N_1239,N_261,N_810);
nand U1240 (N_1240,N_793,In_2178);
nand U1241 (N_1241,N_615,N_313);
nor U1242 (N_1242,In_624,In_1075);
nor U1243 (N_1243,N_917,N_681);
nand U1244 (N_1244,N_111,In_983);
and U1245 (N_1245,In_2383,N_727);
nor U1246 (N_1246,N_919,In_522);
nand U1247 (N_1247,N_757,N_993);
nand U1248 (N_1248,N_478,N_31);
and U1249 (N_1249,In_630,In_2290);
nor U1250 (N_1250,N_740,In_1846);
or U1251 (N_1251,N_804,In_786);
nand U1252 (N_1252,N_421,N_893);
or U1253 (N_1253,N_82,In_160);
xor U1254 (N_1254,N_891,N_468);
nor U1255 (N_1255,N_573,N_825);
xor U1256 (N_1256,N_983,N_288);
nand U1257 (N_1257,N_199,N_201);
nor U1258 (N_1258,N_227,N_658);
and U1259 (N_1259,N_909,In_2469);
nor U1260 (N_1260,N_633,N_177);
xor U1261 (N_1261,In_1325,In_110);
or U1262 (N_1262,N_401,N_25);
xor U1263 (N_1263,N_957,N_244);
nor U1264 (N_1264,In_1520,N_455);
and U1265 (N_1265,In_1043,N_460);
nand U1266 (N_1266,In_431,N_797);
nor U1267 (N_1267,In_833,N_393);
xnor U1268 (N_1268,In_1169,In_848);
nor U1269 (N_1269,N_286,N_495);
xnor U1270 (N_1270,In_793,In_1770);
nor U1271 (N_1271,N_322,N_723);
and U1272 (N_1272,N_366,In_504);
nor U1273 (N_1273,In_129,N_949);
xor U1274 (N_1274,N_721,In_2082);
and U1275 (N_1275,In_161,In_2195);
nand U1276 (N_1276,In_638,N_952);
and U1277 (N_1277,N_217,N_281);
nor U1278 (N_1278,In_1398,N_53);
or U1279 (N_1279,In_1300,In_1623);
and U1280 (N_1280,N_448,N_178);
and U1281 (N_1281,In_1434,In_1420);
nor U1282 (N_1282,N_760,N_3);
and U1283 (N_1283,N_829,In_416);
and U1284 (N_1284,N_729,N_652);
or U1285 (N_1285,In_2395,N_490);
or U1286 (N_1286,N_374,N_610);
or U1287 (N_1287,N_218,N_424);
and U1288 (N_1288,In_1952,N_272);
and U1289 (N_1289,In_1368,N_99);
or U1290 (N_1290,N_335,N_33);
nor U1291 (N_1291,N_179,N_437);
nand U1292 (N_1292,N_182,N_54);
nor U1293 (N_1293,N_276,In_2366);
xnor U1294 (N_1294,N_22,N_711);
and U1295 (N_1295,N_147,N_367);
xor U1296 (N_1296,N_247,In_1923);
and U1297 (N_1297,N_579,N_79);
xnor U1298 (N_1298,N_239,In_83);
nand U1299 (N_1299,In_2445,In_2099);
or U1300 (N_1300,N_206,N_655);
or U1301 (N_1301,N_846,In_1312);
nand U1302 (N_1302,N_782,N_619);
and U1303 (N_1303,N_394,N_986);
nand U1304 (N_1304,N_663,N_741);
xor U1305 (N_1305,In_722,N_969);
and U1306 (N_1306,In_2258,In_1501);
and U1307 (N_1307,N_324,In_1849);
or U1308 (N_1308,N_124,N_150);
nor U1309 (N_1309,N_571,In_1051);
nand U1310 (N_1310,N_958,N_510);
nor U1311 (N_1311,N_767,N_376);
nor U1312 (N_1312,N_631,In_627);
xnor U1313 (N_1313,N_98,N_669);
nor U1314 (N_1314,N_859,N_237);
or U1315 (N_1315,In_1745,N_775);
nor U1316 (N_1316,In_1518,N_240);
or U1317 (N_1317,In_2411,N_108);
nand U1318 (N_1318,N_34,In_1195);
and U1319 (N_1319,In_18,In_1489);
nor U1320 (N_1320,N_458,N_414);
and U1321 (N_1321,N_818,N_661);
or U1322 (N_1322,N_515,N_720);
xnor U1323 (N_1323,In_144,N_130);
and U1324 (N_1324,N_208,N_572);
nand U1325 (N_1325,N_719,N_163);
nor U1326 (N_1326,N_90,N_922);
nor U1327 (N_1327,In_328,N_56);
or U1328 (N_1328,N_734,In_792);
nor U1329 (N_1329,N_59,N_592);
xor U1330 (N_1330,N_689,N_419);
and U1331 (N_1331,N_962,In_1449);
or U1332 (N_1332,N_316,N_260);
xor U1333 (N_1333,N_574,N_215);
nand U1334 (N_1334,N_183,N_128);
nor U1335 (N_1335,N_981,N_38);
and U1336 (N_1336,N_47,In_297);
nand U1337 (N_1337,N_256,N_326);
nand U1338 (N_1338,N_259,N_368);
or U1339 (N_1339,N_135,N_558);
nand U1340 (N_1340,In_966,In_2268);
xnor U1341 (N_1341,N_941,N_282);
or U1342 (N_1342,N_250,N_755);
xor U1343 (N_1343,In_264,N_204);
nand U1344 (N_1344,In_1257,In_166);
xnor U1345 (N_1345,N_713,N_964);
or U1346 (N_1346,In_1359,N_961);
nand U1347 (N_1347,In_200,In_675);
and U1348 (N_1348,N_331,N_834);
or U1349 (N_1349,In_1435,N_115);
or U1350 (N_1350,N_83,N_30);
nor U1351 (N_1351,N_348,In_761);
and U1352 (N_1352,In_2059,N_95);
xor U1353 (N_1353,N_145,N_897);
xnor U1354 (N_1354,N_294,N_907);
or U1355 (N_1355,N_625,In_222);
nor U1356 (N_1356,N_995,N_105);
xor U1357 (N_1357,N_487,In_1034);
xor U1358 (N_1358,N_434,N_934);
nor U1359 (N_1359,In_865,In_226);
nor U1360 (N_1360,N_85,In_599);
nor U1361 (N_1361,N_45,N_892);
or U1362 (N_1362,N_671,N_594);
xor U1363 (N_1363,In_1334,In_209);
or U1364 (N_1364,N_242,N_454);
and U1365 (N_1365,In_133,N_341);
nor U1366 (N_1366,N_133,N_523);
xor U1367 (N_1367,N_860,N_991);
xor U1368 (N_1368,In_1723,N_735);
and U1369 (N_1369,N_100,N_942);
nand U1370 (N_1370,In_2289,In_782);
nand U1371 (N_1371,In_1951,N_899);
or U1372 (N_1372,In_822,In_1073);
nand U1373 (N_1373,N_811,N_271);
and U1374 (N_1374,N_642,N_978);
nor U1375 (N_1375,N_330,N_93);
or U1376 (N_1376,N_552,N_530);
and U1377 (N_1377,N_857,N_992);
nand U1378 (N_1378,N_116,N_979);
or U1379 (N_1379,N_212,N_486);
or U1380 (N_1380,N_968,N_329);
or U1381 (N_1381,N_876,In_1184);
and U1382 (N_1382,In_871,N_304);
xnor U1383 (N_1383,N_963,N_37);
or U1384 (N_1384,N_443,In_1933);
nand U1385 (N_1385,In_258,N_781);
and U1386 (N_1386,N_426,N_63);
nand U1387 (N_1387,N_160,In_1068);
xor U1388 (N_1388,N_319,N_805);
xnor U1389 (N_1389,N_16,N_323);
xor U1390 (N_1390,In_1352,N_609);
xnor U1391 (N_1391,N_617,In_1337);
nand U1392 (N_1392,N_561,In_1444);
xnor U1393 (N_1393,In_1525,N_392);
and U1394 (N_1394,N_439,In_549);
or U1395 (N_1395,N_336,In_427);
xor U1396 (N_1396,N_377,N_747);
and U1397 (N_1397,N_639,N_785);
and U1398 (N_1398,N_269,N_347);
nor U1399 (N_1399,N_138,N_428);
xnor U1400 (N_1400,In_324,N_125);
nor U1401 (N_1401,N_0,In_2302);
or U1402 (N_1402,N_851,N_8);
nor U1403 (N_1403,In_1796,In_311);
or U1404 (N_1404,N_673,In_1955);
nor U1405 (N_1405,N_162,N_771);
and U1406 (N_1406,In_128,N_365);
nand U1407 (N_1407,N_634,In_367);
xnor U1408 (N_1408,N_667,N_562);
nand U1409 (N_1409,In_840,In_1477);
and U1410 (N_1410,N_191,N_66);
nor U1411 (N_1411,N_790,N_371);
nor U1412 (N_1412,In_1299,N_214);
nor U1413 (N_1413,N_875,N_166);
nor U1414 (N_1414,N_606,N_236);
xor U1415 (N_1415,N_266,N_954);
and U1416 (N_1416,In_1536,N_431);
xor U1417 (N_1417,N_898,In_842);
xnor U1418 (N_1418,In_214,N_520);
xor U1419 (N_1419,In_824,N_597);
or U1420 (N_1420,In_1469,In_391);
or U1421 (N_1421,In_366,In_1529);
or U1422 (N_1422,N_548,In_1754);
and U1423 (N_1423,N_706,N_649);
or U1424 (N_1424,In_132,In_826);
xor U1425 (N_1425,N_171,N_630);
or U1426 (N_1426,N_298,N_113);
or U1427 (N_1427,N_500,N_596);
or U1428 (N_1428,In_2335,In_325);
and U1429 (N_1429,N_41,In_471);
xnor U1430 (N_1430,In_213,N_464);
nor U1431 (N_1431,In_1752,N_117);
and U1432 (N_1432,N_636,In_981);
nand U1433 (N_1433,In_569,In_468);
and U1434 (N_1434,N_827,N_582);
nand U1435 (N_1435,N_789,In_821);
nor U1436 (N_1436,N_213,N_106);
and U1437 (N_1437,N_674,In_1642);
and U1438 (N_1438,In_107,N_164);
and U1439 (N_1439,In_1995,N_231);
nand U1440 (N_1440,In_2456,N_192);
or U1441 (N_1441,In_960,N_488);
or U1442 (N_1442,In_443,In_389);
nor U1443 (N_1443,N_91,N_867);
xnor U1444 (N_1444,N_896,In_1247);
nand U1445 (N_1445,In_1135,N_402);
or U1446 (N_1446,N_89,N_575);
or U1447 (N_1447,N_904,N_838);
nor U1448 (N_1448,In_1561,N_436);
or U1449 (N_1449,N_14,N_843);
and U1450 (N_1450,N_945,In_88);
nor U1451 (N_1451,N_446,N_831);
or U1452 (N_1452,In_1747,N_746);
and U1453 (N_1453,In_1488,N_840);
nand U1454 (N_1454,N_930,N_637);
nor U1455 (N_1455,In_1894,In_2271);
nor U1456 (N_1456,N_383,In_1424);
nor U1457 (N_1457,N_758,In_2311);
nor U1458 (N_1458,In_2448,N_599);
nor U1459 (N_1459,In_266,In_1392);
or U1460 (N_1460,N_994,N_28);
nor U1461 (N_1461,N_823,In_1442);
nor U1462 (N_1462,N_143,N_284);
nor U1463 (N_1463,In_1499,In_1860);
nand U1464 (N_1464,In_1881,In_2108);
nor U1465 (N_1465,In_723,N_972);
xnor U1466 (N_1466,N_86,N_534);
and U1467 (N_1467,N_806,N_600);
nand U1468 (N_1468,N_295,In_901);
or U1469 (N_1469,In_2252,In_1010);
xnor U1470 (N_1470,In_1083,N_693);
xor U1471 (N_1471,In_1451,N_787);
or U1472 (N_1472,N_410,In_1782);
or U1473 (N_1473,N_127,N_228);
xnor U1474 (N_1474,N_752,In_1878);
or U1475 (N_1475,N_730,In_1683);
nand U1476 (N_1476,In_1036,N_916);
xor U1477 (N_1477,N_644,In_1582);
and U1478 (N_1478,N_207,N_629);
nor U1479 (N_1479,N_650,N_267);
xor U1480 (N_1480,N_745,N_514);
nand U1481 (N_1481,In_1834,N_996);
xnor U1482 (N_1482,N_200,N_466);
and U1483 (N_1483,N_895,In_929);
and U1484 (N_1484,N_506,N_503);
and U1485 (N_1485,N_325,In_76);
nor U1486 (N_1486,In_1692,N_10);
xor U1487 (N_1487,In_50,N_4);
or U1488 (N_1488,N_716,N_232);
xor U1489 (N_1489,N_142,N_540);
nor U1490 (N_1490,In_1370,N_234);
or U1491 (N_1491,N_632,N_249);
nor U1492 (N_1492,N_296,In_667);
nor U1493 (N_1493,N_360,N_803);
or U1494 (N_1494,N_778,N_190);
nand U1495 (N_1495,N_103,N_317);
nor U1496 (N_1496,In_1507,N_308);
and U1497 (N_1497,N_715,N_309);
and U1498 (N_1498,N_473,In_757);
nor U1499 (N_1499,In_2230,N_476);
xor U1500 (N_1500,N_299,N_80);
xor U1501 (N_1501,N_152,N_445);
and U1502 (N_1502,N_452,N_168);
nor U1503 (N_1503,N_352,In_607);
nand U1504 (N_1504,N_847,In_1919);
xnor U1505 (N_1505,In_1229,N_975);
nand U1506 (N_1506,N_535,N_97);
xor U1507 (N_1507,N_872,In_2405);
and U1508 (N_1508,N_837,In_1515);
nand U1509 (N_1509,In_466,N_531);
nor U1510 (N_1510,N_696,N_651);
or U1511 (N_1511,In_184,In_2181);
xnor U1512 (N_1512,N_944,N_189);
nand U1513 (N_1513,N_532,N_824);
and U1514 (N_1514,N_362,N_588);
xor U1515 (N_1515,In_1516,N_874);
and U1516 (N_1516,N_75,N_275);
or U1517 (N_1517,N_576,N_252);
and U1518 (N_1518,N_666,In_743);
and U1519 (N_1519,N_544,N_270);
xnor U1520 (N_1520,In_1814,N_933);
xnor U1521 (N_1521,N_126,In_2239);
or U1522 (N_1522,N_21,N_151);
and U1523 (N_1523,N_936,N_833);
and U1524 (N_1524,In_2308,N_223);
and U1525 (N_1525,In_1828,N_279);
xor U1526 (N_1526,In_1669,In_937);
or U1527 (N_1527,N_235,N_668);
nor U1528 (N_1528,N_943,In_489);
or U1529 (N_1529,N_900,N_885);
xnor U1530 (N_1530,N_759,N_844);
nor U1531 (N_1531,In_1258,N_440);
or U1532 (N_1532,N_2,N_451);
or U1533 (N_1533,N_194,In_2204);
or U1534 (N_1534,In_1662,In_2075);
xnor U1535 (N_1535,N_403,In_550);
nand U1536 (N_1536,N_784,In_1621);
xor U1537 (N_1537,N_970,In_1137);
nor U1538 (N_1538,N_598,In_1900);
nor U1539 (N_1539,In_1658,N_120);
xnor U1540 (N_1540,In_2340,N_880);
xor U1541 (N_1541,N_112,N_96);
or U1542 (N_1542,In_647,In_573);
or U1543 (N_1543,In_553,In_1694);
or U1544 (N_1544,N_19,N_556);
and U1545 (N_1545,N_74,In_2087);
nor U1546 (N_1546,In_705,N_311);
nor U1547 (N_1547,N_704,N_18);
nand U1548 (N_1548,N_565,N_795);
nor U1549 (N_1549,N_801,In_75);
and U1550 (N_1550,In_1581,In_1272);
xnor U1551 (N_1551,N_643,In_261);
or U1552 (N_1552,N_425,N_159);
nand U1553 (N_1553,In_2360,N_154);
nor U1554 (N_1554,In_315,N_492);
or U1555 (N_1555,In_799,In_2377);
nor U1556 (N_1556,N_221,N_800);
or U1557 (N_1557,N_442,N_219);
nor U1558 (N_1558,In_776,N_564);
or U1559 (N_1559,In_2221,N_167);
nand U1560 (N_1560,In_1371,N_516);
nor U1561 (N_1561,N_543,N_660);
xnor U1562 (N_1562,N_441,N_697);
and U1563 (N_1563,N_211,N_819);
nor U1564 (N_1564,N_761,N_327);
xnor U1565 (N_1565,N_887,N_134);
or U1566 (N_1566,In_1331,In_507);
nand U1567 (N_1567,N_72,In_2355);
xnor U1568 (N_1568,N_683,N_255);
xor U1569 (N_1569,N_850,N_285);
nand U1570 (N_1570,In_1054,In_1608);
and U1571 (N_1571,N_502,In_1384);
or U1572 (N_1572,N_569,N_39);
and U1573 (N_1573,N_195,In_1939);
nor U1574 (N_1574,N_233,N_110);
and U1575 (N_1575,N_263,N_662);
or U1576 (N_1576,N_44,N_405);
nor U1577 (N_1577,N_469,N_158);
and U1578 (N_1578,N_869,N_229);
and U1579 (N_1579,In_856,N_841);
nor U1580 (N_1580,In_2213,In_1697);
nor U1581 (N_1581,N_156,In_109);
nor U1582 (N_1582,N_225,N_61);
and U1583 (N_1583,N_6,N_533);
nor U1584 (N_1584,N_137,In_565);
nand U1585 (N_1585,N_984,N_129);
nor U1586 (N_1586,N_708,N_718);
xnor U1587 (N_1587,N_389,N_603);
or U1588 (N_1588,N_527,In_967);
or U1589 (N_1589,N_648,N_107);
nand U1590 (N_1590,N_853,N_73);
or U1591 (N_1591,In_1667,N_765);
or U1592 (N_1592,In_0,N_768);
xor U1593 (N_1593,N_682,In_2167);
and U1594 (N_1594,In_1303,In_797);
and U1595 (N_1595,N_925,N_822);
or U1596 (N_1596,N_1,N_959);
nand U1597 (N_1597,In_1554,N_707);
and U1598 (N_1598,N_946,N_447);
or U1599 (N_1599,N_132,N_243);
and U1600 (N_1600,In_2103,In_539);
and U1601 (N_1601,N_913,In_2276);
or U1602 (N_1602,In_2234,N_881);
or U1603 (N_1603,N_863,N_657);
or U1604 (N_1604,N_13,In_2012);
and U1605 (N_1605,N_370,In_811);
and U1606 (N_1606,In_1429,N_980);
or U1607 (N_1607,N_877,In_1287);
nor U1608 (N_1608,In_1500,N_449);
nor U1609 (N_1609,N_560,N_43);
xnor U1610 (N_1610,In_439,In_115);
nor U1611 (N_1611,N_193,N_710);
and U1612 (N_1612,N_380,N_369);
xnor U1613 (N_1613,N_647,In_1575);
nand U1614 (N_1614,In_1328,In_2229);
nor U1615 (N_1615,N_686,N_595);
or U1616 (N_1616,In_65,In_1959);
or U1617 (N_1617,N_932,N_587);
and U1618 (N_1618,In_498,In_985);
xor U1619 (N_1619,N_289,N_537);
xor U1620 (N_1620,N_364,In_7);
or U1621 (N_1621,N_131,N_57);
and U1622 (N_1622,N_813,N_52);
or U1623 (N_1623,In_1297,In_70);
nor U1624 (N_1624,In_1116,N_612);
nand U1625 (N_1625,N_444,N_300);
nand U1626 (N_1626,N_346,In_1812);
and U1627 (N_1627,N_938,N_712);
and U1628 (N_1628,In_556,N_372);
nand U1629 (N_1629,N_184,N_665);
nand U1630 (N_1630,N_640,N_971);
or U1631 (N_1631,In_1842,N_738);
nor U1632 (N_1632,N_181,N_321);
xnor U1633 (N_1633,In_1603,N_737);
xor U1634 (N_1634,N_101,N_334);
and U1635 (N_1635,In_649,In_1367);
and U1636 (N_1636,N_314,N_491);
or U1637 (N_1637,N_786,N_384);
or U1638 (N_1638,N_471,N_915);
or U1639 (N_1639,N_224,N_453);
nor U1640 (N_1640,In_2020,N_400);
xor U1641 (N_1641,In_2134,In_1427);
xor U1642 (N_1642,N_328,N_121);
or U1643 (N_1643,In_1655,In_353);
xor U1644 (N_1644,N_748,In_1641);
or U1645 (N_1645,In_2257,In_1549);
xnor U1646 (N_1646,N_494,N_459);
and U1647 (N_1647,N_808,In_602);
or U1648 (N_1648,In_726,N_835);
nand U1649 (N_1649,N_960,N_87);
nor U1650 (N_1650,N_714,N_216);
and U1651 (N_1651,N_312,N_92);
xnor U1652 (N_1652,In_2025,In_1829);
xnor U1653 (N_1653,N_462,N_381);
nor U1654 (N_1654,In_68,In_1815);
and U1655 (N_1655,N_815,N_722);
or U1656 (N_1656,N_563,In_409);
and U1657 (N_1657,N_176,N_359);
xor U1658 (N_1658,N_196,N_702);
or U1659 (N_1659,In_1419,N_465);
nor U1660 (N_1660,N_306,In_2071);
nand U1661 (N_1661,N_315,In_1695);
xnor U1662 (N_1662,N_202,In_1216);
nor U1663 (N_1663,N_496,N_345);
or U1664 (N_1664,In_1185,N_879);
nor U1665 (N_1665,In_1757,N_749);
xor U1666 (N_1666,N_724,N_570);
nand U1667 (N_1667,N_386,N_590);
or U1668 (N_1668,N_472,In_179);
and U1669 (N_1669,In_2347,N_842);
nor U1670 (N_1670,In_241,In_81);
nor U1671 (N_1671,N_475,N_187);
or U1672 (N_1672,In_1836,In_1095);
and U1673 (N_1673,N_870,N_586);
nand U1674 (N_1674,N_593,N_485);
or U1675 (N_1675,In_1019,N_413);
xnor U1676 (N_1676,N_483,N_882);
and U1677 (N_1677,N_616,N_484);
and U1678 (N_1678,In_2479,In_1837);
or U1679 (N_1679,N_418,N_773);
and U1680 (N_1680,N_743,N_342);
nand U1681 (N_1681,N_230,N_118);
nand U1682 (N_1682,N_566,N_998);
xnor U1683 (N_1683,In_384,N_361);
nor U1684 (N_1684,In_2280,N_173);
nor U1685 (N_1685,In_2177,N_245);
nor U1686 (N_1686,N_908,N_482);
nor U1687 (N_1687,N_605,N_68);
or U1688 (N_1688,N_358,N_889);
nor U1689 (N_1689,N_627,N_480);
nor U1690 (N_1690,N_51,N_951);
nor U1691 (N_1691,N_283,In_1819);
xor U1692 (N_1692,N_873,N_536);
nand U1693 (N_1693,N_477,N_77);
or U1694 (N_1694,N_258,N_982);
nor U1695 (N_1695,N_973,N_210);
nor U1696 (N_1696,N_705,N_577);
nand U1697 (N_1697,N_354,In_2376);
and U1698 (N_1698,N_339,N_429);
and U1699 (N_1699,N_731,In_235);
nand U1700 (N_1700,N_832,N_624);
nor U1701 (N_1701,In_1041,N_49);
or U1702 (N_1702,N_438,N_528);
xor U1703 (N_1703,In_2387,N_883);
nor U1704 (N_1704,N_153,N_64);
or U1705 (N_1705,In_1440,N_501);
nand U1706 (N_1706,N_890,N_50);
and U1707 (N_1707,N_826,In_571);
nor U1708 (N_1708,In_62,In_847);
and U1709 (N_1709,N_391,In_1905);
xor U1710 (N_1710,N_809,N_865);
and U1711 (N_1711,N_375,N_691);
and U1712 (N_1712,N_144,N_509);
or U1713 (N_1713,N_776,In_2224);
and U1714 (N_1714,In_2378,In_746);
and U1715 (N_1715,N_24,N_854);
xnor U1716 (N_1716,N_699,N_836);
nor U1717 (N_1717,N_852,N_474);
or U1718 (N_1718,In_2062,In_2006);
nand U1719 (N_1719,N_415,In_1717);
nand U1720 (N_1720,In_734,N_27);
xnor U1721 (N_1721,N_762,N_517);
and U1722 (N_1722,In_1097,N_910);
nand U1723 (N_1723,N_821,N_493);
nand U1724 (N_1724,N_679,N_251);
nor U1725 (N_1725,N_398,N_685);
or U1726 (N_1726,N_845,In_2183);
nor U1727 (N_1727,N_728,N_871);
and U1728 (N_1728,N_417,N_387);
and U1729 (N_1729,In_1382,In_2319);
or U1730 (N_1730,In_2142,In_157);
and U1731 (N_1731,N_62,N_935);
nor U1732 (N_1732,N_807,N_659);
or U1733 (N_1733,In_686,In_1167);
and U1734 (N_1734,N_12,N_209);
or U1735 (N_1735,In_1291,N_794);
xor U1736 (N_1736,N_675,In_494);
or U1737 (N_1737,In_1906,In_1850);
nand U1738 (N_1738,N_102,In_1220);
nand U1739 (N_1739,N_614,In_1121);
and U1740 (N_1740,In_204,In_314);
xnor U1741 (N_1741,N_830,N_388);
or U1742 (N_1742,N_411,N_353);
and U1743 (N_1743,N_435,N_928);
nand U1744 (N_1744,N_553,N_868);
or U1745 (N_1745,N_796,N_584);
and U1746 (N_1746,N_357,N_337);
xor U1747 (N_1747,N_687,N_783);
nor U1748 (N_1748,In_1986,In_1402);
nand U1749 (N_1749,N_965,In_721);
nand U1750 (N_1750,In_1747,N_408);
or U1751 (N_1751,In_2181,In_1200);
or U1752 (N_1752,N_687,N_616);
xnor U1753 (N_1753,N_836,In_1822);
xor U1754 (N_1754,N_117,N_314);
or U1755 (N_1755,N_250,N_371);
nor U1756 (N_1756,In_83,N_291);
and U1757 (N_1757,N_837,In_761);
nand U1758 (N_1758,In_2448,N_693);
xnor U1759 (N_1759,N_525,N_504);
and U1760 (N_1760,N_926,In_833);
and U1761 (N_1761,In_503,In_2340);
nand U1762 (N_1762,In_2271,In_2178);
nand U1763 (N_1763,N_823,N_842);
and U1764 (N_1764,In_1881,In_353);
nor U1765 (N_1765,N_332,N_38);
xnor U1766 (N_1766,N_563,N_438);
and U1767 (N_1767,N_20,N_254);
and U1768 (N_1768,N_661,N_314);
xor U1769 (N_1769,N_516,In_2221);
xnor U1770 (N_1770,N_819,N_536);
xor U1771 (N_1771,N_613,In_565);
nand U1772 (N_1772,N_510,In_2062);
or U1773 (N_1773,N_204,N_246);
nand U1774 (N_1774,N_661,In_573);
nand U1775 (N_1775,In_200,N_199);
or U1776 (N_1776,N_604,N_363);
nor U1777 (N_1777,In_391,N_408);
nand U1778 (N_1778,N_564,In_667);
xnor U1779 (N_1779,N_734,N_343);
xor U1780 (N_1780,In_1894,N_790);
nor U1781 (N_1781,N_102,In_760);
nor U1782 (N_1782,N_996,N_559);
nand U1783 (N_1783,In_272,N_592);
nand U1784 (N_1784,In_1755,N_174);
xor U1785 (N_1785,N_677,N_902);
and U1786 (N_1786,In_50,In_427);
nor U1787 (N_1787,N_759,In_1371);
and U1788 (N_1788,N_415,N_476);
nand U1789 (N_1789,N_660,In_1561);
nor U1790 (N_1790,N_433,N_42);
or U1791 (N_1791,N_613,In_1869);
and U1792 (N_1792,N_55,N_259);
nand U1793 (N_1793,N_126,N_956);
nand U1794 (N_1794,N_656,N_770);
nor U1795 (N_1795,In_2290,N_324);
xor U1796 (N_1796,N_532,N_754);
nand U1797 (N_1797,N_726,In_2289);
or U1798 (N_1798,In_624,In_387);
and U1799 (N_1799,N_303,N_231);
and U1800 (N_1800,N_93,N_602);
or U1801 (N_1801,N_977,In_1182);
and U1802 (N_1802,N_631,N_165);
and U1803 (N_1803,In_1359,N_846);
or U1804 (N_1804,In_1218,In_726);
nand U1805 (N_1805,N_585,In_83);
and U1806 (N_1806,N_438,N_353);
nor U1807 (N_1807,N_695,In_144);
or U1808 (N_1808,N_584,In_2335);
or U1809 (N_1809,N_997,N_791);
nor U1810 (N_1810,N_210,N_45);
nand U1811 (N_1811,In_1757,N_583);
nand U1812 (N_1812,N_280,N_62);
nand U1813 (N_1813,In_1829,N_13);
nand U1814 (N_1814,N_891,N_921);
and U1815 (N_1815,N_398,N_669);
or U1816 (N_1816,N_327,In_107);
and U1817 (N_1817,N_717,In_808);
and U1818 (N_1818,N_121,N_944);
xor U1819 (N_1819,N_277,N_494);
and U1820 (N_1820,In_129,N_14);
or U1821 (N_1821,N_977,N_596);
nand U1822 (N_1822,N_148,In_1655);
xnor U1823 (N_1823,N_323,N_477);
and U1824 (N_1824,In_1371,N_294);
nor U1825 (N_1825,In_1947,N_917);
and U1826 (N_1826,N_765,N_111);
and U1827 (N_1827,In_81,N_352);
nand U1828 (N_1828,N_156,N_910);
nand U1829 (N_1829,N_2,In_504);
nand U1830 (N_1830,N_162,N_712);
xor U1831 (N_1831,N_721,N_201);
and U1832 (N_1832,N_607,N_913);
nor U1833 (N_1833,N_514,N_364);
and U1834 (N_1834,In_1554,N_546);
or U1835 (N_1835,N_371,N_8);
or U1836 (N_1836,N_153,N_996);
nand U1837 (N_1837,N_426,N_235);
and U1838 (N_1838,N_144,N_821);
or U1839 (N_1839,N_400,N_228);
or U1840 (N_1840,In_1952,N_355);
and U1841 (N_1841,N_355,In_1392);
and U1842 (N_1842,N_175,In_856);
nand U1843 (N_1843,N_282,N_177);
and U1844 (N_1844,N_666,N_524);
or U1845 (N_1845,N_29,N_506);
and U1846 (N_1846,N_901,In_498);
nor U1847 (N_1847,N_362,In_705);
xnor U1848 (N_1848,N_54,In_1959);
xnor U1849 (N_1849,N_193,N_138);
nand U1850 (N_1850,N_246,N_35);
nand U1851 (N_1851,N_181,N_760);
or U1852 (N_1852,In_1282,N_216);
nor U1853 (N_1853,In_116,In_1337);
and U1854 (N_1854,In_531,In_627);
or U1855 (N_1855,In_65,In_353);
nor U1856 (N_1856,N_605,In_856);
and U1857 (N_1857,In_399,In_976);
or U1858 (N_1858,N_187,In_967);
nand U1859 (N_1859,In_983,N_415);
nor U1860 (N_1860,N_621,N_472);
nand U1861 (N_1861,In_427,N_819);
or U1862 (N_1862,In_70,N_230);
nand U1863 (N_1863,N_583,N_397);
nor U1864 (N_1864,N_374,In_2361);
and U1865 (N_1865,N_955,In_1362);
or U1866 (N_1866,In_726,N_932);
nor U1867 (N_1867,N_118,N_794);
nor U1868 (N_1868,In_363,N_956);
and U1869 (N_1869,N_864,N_33);
and U1870 (N_1870,N_624,N_661);
or U1871 (N_1871,In_565,N_339);
xor U1872 (N_1872,N_634,N_163);
xor U1873 (N_1873,N_128,N_822);
and U1874 (N_1874,In_2275,N_521);
xor U1875 (N_1875,N_2,N_519);
xnor U1876 (N_1876,N_384,In_1477);
xnor U1877 (N_1877,In_213,N_900);
xor U1878 (N_1878,In_1008,N_310);
nor U1879 (N_1879,In_1869,In_1162);
or U1880 (N_1880,In_1068,In_579);
or U1881 (N_1881,N_73,In_1422);
nor U1882 (N_1882,In_1662,N_151);
or U1883 (N_1883,N_930,N_897);
nand U1884 (N_1884,In_311,N_697);
nand U1885 (N_1885,N_259,In_110);
and U1886 (N_1886,N_708,N_42);
and U1887 (N_1887,N_92,N_362);
nand U1888 (N_1888,N_546,In_399);
xnor U1889 (N_1889,N_271,In_847);
nor U1890 (N_1890,N_8,N_485);
nand U1891 (N_1891,In_1623,In_1442);
xor U1892 (N_1892,In_133,N_417);
nor U1893 (N_1893,N_25,N_434);
and U1894 (N_1894,In_2472,N_940);
and U1895 (N_1895,In_83,N_920);
and U1896 (N_1896,In_2366,N_468);
xor U1897 (N_1897,In_1695,N_449);
xnor U1898 (N_1898,In_793,In_1476);
nand U1899 (N_1899,N_17,N_550);
nor U1900 (N_1900,N_668,N_520);
or U1901 (N_1901,In_1667,N_414);
and U1902 (N_1902,In_7,N_135);
nor U1903 (N_1903,N_647,N_269);
nand U1904 (N_1904,In_1095,In_1282);
and U1905 (N_1905,N_616,N_789);
xnor U1906 (N_1906,N_359,N_390);
nor U1907 (N_1907,In_1182,N_825);
xor U1908 (N_1908,N_425,In_1435);
nand U1909 (N_1909,In_1919,In_1662);
nand U1910 (N_1910,In_983,In_469);
xnor U1911 (N_1911,In_336,N_896);
xnor U1912 (N_1912,N_960,In_2230);
and U1913 (N_1913,N_523,N_468);
nand U1914 (N_1914,N_699,In_1182);
or U1915 (N_1915,N_636,In_328);
nand U1916 (N_1916,N_247,N_777);
xnor U1917 (N_1917,N_670,In_1754);
nor U1918 (N_1918,N_695,In_1520);
or U1919 (N_1919,N_75,N_2);
xor U1920 (N_1920,In_436,N_444);
and U1921 (N_1921,N_60,N_894);
xnor U1922 (N_1922,N_414,In_426);
xnor U1923 (N_1923,N_205,N_317);
nor U1924 (N_1924,In_565,N_746);
nand U1925 (N_1925,N_896,N_533);
nand U1926 (N_1926,N_907,N_872);
nand U1927 (N_1927,N_214,N_468);
nor U1928 (N_1928,N_355,In_1121);
or U1929 (N_1929,N_221,In_2432);
and U1930 (N_1930,In_531,N_676);
and U1931 (N_1931,In_1037,In_2411);
and U1932 (N_1932,N_593,N_662);
xnor U1933 (N_1933,In_1434,N_4);
nor U1934 (N_1934,N_491,N_558);
and U1935 (N_1935,N_994,N_504);
and U1936 (N_1936,N_257,In_753);
and U1937 (N_1937,N_487,N_733);
or U1938 (N_1938,N_442,N_789);
and U1939 (N_1939,In_1846,N_592);
and U1940 (N_1940,N_928,N_496);
or U1941 (N_1941,N_378,In_2481);
nor U1942 (N_1942,N_291,N_980);
and U1943 (N_1943,N_701,N_394);
xor U1944 (N_1944,N_731,N_747);
nand U1945 (N_1945,N_946,N_386);
nand U1946 (N_1946,N_372,In_629);
and U1947 (N_1947,N_259,N_201);
xnor U1948 (N_1948,N_195,In_630);
nor U1949 (N_1949,N_684,N_164);
nor U1950 (N_1950,In_1283,N_345);
xor U1951 (N_1951,N_950,N_47);
nor U1952 (N_1952,N_667,N_597);
xnor U1953 (N_1953,In_753,N_355);
nand U1954 (N_1954,In_1303,In_1641);
and U1955 (N_1955,N_947,N_99);
nand U1956 (N_1956,N_572,N_890);
or U1957 (N_1957,In_1424,In_1041);
or U1958 (N_1958,In_1932,N_693);
nor U1959 (N_1959,N_348,N_939);
nand U1960 (N_1960,N_731,In_343);
nand U1961 (N_1961,N_892,N_598);
or U1962 (N_1962,In_248,In_522);
or U1963 (N_1963,N_379,N_471);
nor U1964 (N_1964,In_1695,In_776);
nand U1965 (N_1965,N_294,In_537);
and U1966 (N_1966,N_188,N_319);
nand U1967 (N_1967,N_329,N_169);
xnor U1968 (N_1968,N_263,N_260);
or U1969 (N_1969,N_591,In_324);
nor U1970 (N_1970,N_139,N_222);
and U1971 (N_1971,In_2448,N_506);
or U1972 (N_1972,In_793,In_1819);
nor U1973 (N_1973,N_808,N_9);
or U1974 (N_1974,N_42,In_2224);
and U1975 (N_1975,N_897,In_1642);
nand U1976 (N_1976,In_1392,N_385);
nand U1977 (N_1977,N_136,N_332);
nor U1978 (N_1978,N_186,N_193);
and U1979 (N_1979,N_879,N_67);
nand U1980 (N_1980,In_2229,In_1554);
or U1981 (N_1981,N_723,N_215);
nand U1982 (N_1982,N_131,In_639);
and U1983 (N_1983,In_439,N_496);
and U1984 (N_1984,In_746,N_966);
and U1985 (N_1985,In_1178,In_821);
nand U1986 (N_1986,In_929,N_671);
xor U1987 (N_1987,N_368,In_1041);
nand U1988 (N_1988,In_1558,N_602);
and U1989 (N_1989,In_2472,N_744);
nor U1990 (N_1990,N_546,In_1075);
and U1991 (N_1991,N_621,N_94);
nor U1992 (N_1992,In_1303,In_619);
or U1993 (N_1993,N_479,N_838);
xor U1994 (N_1994,N_667,N_286);
nand U1995 (N_1995,N_535,N_465);
xor U1996 (N_1996,N_617,In_2271);
or U1997 (N_1997,N_325,N_246);
or U1998 (N_1998,N_373,N_21);
or U1999 (N_1999,N_265,N_53);
nand U2000 (N_2000,N_1500,N_1256);
and U2001 (N_2001,N_1409,N_1945);
nor U2002 (N_2002,N_1644,N_1985);
or U2003 (N_2003,N_1812,N_1461);
and U2004 (N_2004,N_1559,N_1343);
or U2005 (N_2005,N_1841,N_1975);
xor U2006 (N_2006,N_1399,N_1227);
xnor U2007 (N_2007,N_1277,N_1471);
or U2008 (N_2008,N_1745,N_1677);
or U2009 (N_2009,N_1808,N_1322);
and U2010 (N_2010,N_1845,N_1600);
xor U2011 (N_2011,N_1269,N_1806);
or U2012 (N_2012,N_1850,N_1484);
nand U2013 (N_2013,N_1444,N_1382);
nor U2014 (N_2014,N_1619,N_1818);
xor U2015 (N_2015,N_1202,N_1166);
nor U2016 (N_2016,N_1417,N_1012);
or U2017 (N_2017,N_1545,N_1063);
and U2018 (N_2018,N_1878,N_1095);
xnor U2019 (N_2019,N_1756,N_1006);
xnor U2020 (N_2020,N_1740,N_1874);
nor U2021 (N_2021,N_1635,N_1214);
and U2022 (N_2022,N_1879,N_1487);
or U2023 (N_2023,N_1001,N_1198);
nand U2024 (N_2024,N_1733,N_1285);
or U2025 (N_2025,N_1314,N_1104);
or U2026 (N_2026,N_1718,N_1414);
xnor U2027 (N_2027,N_1817,N_1317);
nor U2028 (N_2028,N_1720,N_1569);
xnor U2029 (N_2029,N_1318,N_1250);
nand U2030 (N_2030,N_1467,N_1091);
or U2031 (N_2031,N_1286,N_1290);
nor U2032 (N_2032,N_1955,N_1738);
nand U2033 (N_2033,N_1753,N_1336);
or U2034 (N_2034,N_1491,N_1556);
nand U2035 (N_2035,N_1508,N_1355);
or U2036 (N_2036,N_1296,N_1567);
or U2037 (N_2037,N_1831,N_1557);
nand U2038 (N_2038,N_1777,N_1066);
nor U2039 (N_2039,N_1581,N_1998);
xor U2040 (N_2040,N_1853,N_1389);
and U2041 (N_2041,N_1823,N_1734);
nor U2042 (N_2042,N_1425,N_1043);
nand U2043 (N_2043,N_1013,N_1426);
nand U2044 (N_2044,N_1498,N_1843);
or U2045 (N_2045,N_1136,N_1145);
xnor U2046 (N_2046,N_1502,N_1458);
nand U2047 (N_2047,N_1303,N_1598);
and U2048 (N_2048,N_1297,N_1891);
nor U2049 (N_2049,N_1815,N_1371);
or U2050 (N_2050,N_1231,N_1674);
and U2051 (N_2051,N_1180,N_1531);
nor U2052 (N_2052,N_1613,N_1401);
nand U2053 (N_2053,N_1632,N_1793);
nand U2054 (N_2054,N_1321,N_1931);
nand U2055 (N_2055,N_1939,N_1233);
xnor U2056 (N_2056,N_1763,N_1435);
xnor U2057 (N_2057,N_1093,N_1027);
nand U2058 (N_2058,N_1940,N_1701);
xor U2059 (N_2059,N_1479,N_1108);
nor U2060 (N_2060,N_1102,N_1034);
xor U2061 (N_2061,N_1295,N_1640);
xor U2062 (N_2062,N_1638,N_1342);
nand U2063 (N_2063,N_1418,N_1859);
and U2064 (N_2064,N_1149,N_1407);
nor U2065 (N_2065,N_1751,N_1783);
and U2066 (N_2066,N_1625,N_1482);
xor U2067 (N_2067,N_1030,N_1983);
nand U2068 (N_2068,N_1516,N_1980);
nor U2069 (N_2069,N_1512,N_1488);
and U2070 (N_2070,N_1351,N_1493);
nand U2071 (N_2071,N_1114,N_1921);
nand U2072 (N_2072,N_1714,N_1366);
nor U2073 (N_2073,N_1021,N_1924);
nand U2074 (N_2074,N_1881,N_1055);
and U2075 (N_2075,N_1155,N_1947);
and U2076 (N_2076,N_1449,N_1704);
nand U2077 (N_2077,N_1232,N_1851);
nand U2078 (N_2078,N_1164,N_1253);
xnor U2079 (N_2079,N_1272,N_1292);
and U2080 (N_2080,N_1936,N_1046);
and U2081 (N_2081,N_1995,N_1974);
nand U2082 (N_2082,N_1106,N_1052);
or U2083 (N_2083,N_1561,N_1049);
nand U2084 (N_2084,N_1257,N_1098);
nand U2085 (N_2085,N_1147,N_1773);
nor U2086 (N_2086,N_1293,N_1501);
nor U2087 (N_2087,N_1310,N_1304);
nor U2088 (N_2088,N_1190,N_1544);
nor U2089 (N_2089,N_1040,N_1933);
nor U2090 (N_2090,N_1552,N_1284);
nor U2091 (N_2091,N_1835,N_1270);
or U2092 (N_2092,N_1265,N_1634);
nor U2093 (N_2093,N_1927,N_1421);
or U2094 (N_2094,N_1390,N_1919);
xnor U2095 (N_2095,N_1197,N_1228);
or U2096 (N_2096,N_1967,N_1554);
nand U2097 (N_2097,N_1311,N_1624);
nand U2098 (N_2098,N_1956,N_1490);
and U2099 (N_2099,N_1999,N_1650);
xor U2100 (N_2100,N_1386,N_1210);
or U2101 (N_2101,N_1623,N_1798);
and U2102 (N_2102,N_1660,N_1353);
and U2103 (N_2103,N_1008,N_1805);
nor U2104 (N_2104,N_1587,N_1709);
and U2105 (N_2105,N_1462,N_1577);
and U2106 (N_2106,N_1239,N_1476);
nand U2107 (N_2107,N_1562,N_1679);
nor U2108 (N_2108,N_1123,N_1410);
nand U2109 (N_2109,N_1667,N_1408);
and U2110 (N_2110,N_1339,N_1347);
or U2111 (N_2111,N_1573,N_1657);
and U2112 (N_2112,N_1069,N_1163);
and U2113 (N_2113,N_1977,N_1173);
and U2114 (N_2114,N_1837,N_1222);
xor U2115 (N_2115,N_1363,N_1331);
and U2116 (N_2116,N_1869,N_1176);
nand U2117 (N_2117,N_1968,N_1880);
nor U2118 (N_2118,N_1218,N_1703);
nor U2119 (N_2119,N_1896,N_1494);
and U2120 (N_2120,N_1680,N_1861);
nor U2121 (N_2121,N_1264,N_1535);
xor U2122 (N_2122,N_1464,N_1377);
and U2123 (N_2123,N_1235,N_1706);
nand U2124 (N_2124,N_1928,N_1898);
or U2125 (N_2125,N_1521,N_1656);
xnor U2126 (N_2126,N_1193,N_1972);
nand U2127 (N_2127,N_1060,N_1341);
xor U2128 (N_2128,N_1982,N_1530);
and U2129 (N_2129,N_1450,N_1116);
and U2130 (N_2130,N_1828,N_1492);
xnor U2131 (N_2131,N_1586,N_1456);
or U2132 (N_2132,N_1150,N_1737);
or U2133 (N_2133,N_1796,N_1117);
xor U2134 (N_2134,N_1372,N_1071);
and U2135 (N_2135,N_1255,N_1379);
nand U2136 (N_2136,N_1393,N_1966);
and U2137 (N_2137,N_1662,N_1651);
xnor U2138 (N_2138,N_1094,N_1179);
or U2139 (N_2139,N_1062,N_1959);
nor U2140 (N_2140,N_1378,N_1183);
nor U2141 (N_2141,N_1375,N_1814);
xnor U2142 (N_2142,N_1803,N_1068);
xnor U2143 (N_2143,N_1962,N_1769);
xor U2144 (N_2144,N_1298,N_1663);
and U2145 (N_2145,N_1156,N_1029);
or U2146 (N_2146,N_1139,N_1583);
nor U2147 (N_2147,N_1089,N_1816);
xnor U2148 (N_2148,N_1690,N_1873);
or U2149 (N_2149,N_1597,N_1684);
or U2150 (N_2150,N_1329,N_1267);
or U2151 (N_2151,N_1496,N_1801);
or U2152 (N_2152,N_1246,N_1964);
or U2153 (N_2153,N_1011,N_1100);
nor U2154 (N_2154,N_1137,N_1384);
or U2155 (N_2155,N_1234,N_1746);
or U2156 (N_2156,N_1689,N_1770);
nand U2157 (N_2157,N_1489,N_1398);
nor U2158 (N_2158,N_1154,N_1217);
or U2159 (N_2159,N_1084,N_1802);
or U2160 (N_2160,N_1230,N_1178);
and U2161 (N_2161,N_1839,N_1245);
nand U2162 (N_2162,N_1203,N_1912);
and U2163 (N_2163,N_1065,N_1590);
nor U2164 (N_2164,N_1088,N_1504);
or U2165 (N_2165,N_1799,N_1457);
or U2166 (N_2166,N_1997,N_1037);
and U2167 (N_2167,N_1935,N_1134);
and U2168 (N_2168,N_1993,N_1497);
xor U2169 (N_2169,N_1223,N_1963);
and U2170 (N_2170,N_1887,N_1332);
xor U2171 (N_2171,N_1381,N_1266);
or U2172 (N_2172,N_1905,N_1564);
and U2173 (N_2173,N_1054,N_1141);
nand U2174 (N_2174,N_1129,N_1520);
and U2175 (N_2175,N_1988,N_1362);
nand U2176 (N_2176,N_1300,N_1364);
xor U2177 (N_2177,N_1000,N_1862);
xor U2178 (N_2178,N_1367,N_1143);
and U2179 (N_2179,N_1606,N_1731);
nand U2180 (N_2180,N_1758,N_1821);
nand U2181 (N_2181,N_1238,N_1568);
nor U2182 (N_2182,N_1115,N_1244);
and U2183 (N_2183,N_1495,N_1275);
or U2184 (N_2184,N_1165,N_1610);
and U2185 (N_2185,N_1118,N_1990);
xnor U2186 (N_2186,N_1320,N_1533);
or U2187 (N_2187,N_1026,N_1215);
and U2188 (N_2188,N_1423,N_1876);
and U2189 (N_2189,N_1057,N_1790);
nand U2190 (N_2190,N_1205,N_1757);
nor U2191 (N_2191,N_1648,N_1360);
or U2192 (N_2192,N_1944,N_1468);
nor U2193 (N_2193,N_1161,N_1454);
and U2194 (N_2194,N_1641,N_1101);
nor U2195 (N_2195,N_1965,N_1510);
nand U2196 (N_2196,N_1121,N_1683);
xor U2197 (N_2197,N_1427,N_1306);
xor U2198 (N_2198,N_1728,N_1455);
nor U2199 (N_2199,N_1526,N_1415);
or U2200 (N_2200,N_1283,N_1204);
nor U2201 (N_2201,N_1469,N_1620);
nor U2202 (N_2202,N_1434,N_1185);
and U2203 (N_2203,N_1307,N_1323);
nand U2204 (N_2204,N_1926,N_1614);
nand U2205 (N_2205,N_1044,N_1908);
nand U2206 (N_2206,N_1429,N_1659);
and U2207 (N_2207,N_1574,N_1221);
nor U2208 (N_2208,N_1127,N_1327);
nand U2209 (N_2209,N_1540,N_1888);
or U2210 (N_2210,N_1105,N_1755);
nor U2211 (N_2211,N_1599,N_1394);
or U2212 (N_2212,N_1688,N_1991);
xor U2213 (N_2213,N_1992,N_1181);
xnor U2214 (N_2214,N_1268,N_1133);
nand U2215 (N_2215,N_1396,N_1589);
xnor U2216 (N_2216,N_1788,N_1645);
xor U2217 (N_2217,N_1611,N_1826);
and U2218 (N_2218,N_1092,N_1686);
nor U2219 (N_2219,N_1359,N_1937);
or U2220 (N_2220,N_1082,N_1023);
xnor U2221 (N_2221,N_1830,N_1315);
and U2222 (N_2222,N_1532,N_1595);
nor U2223 (N_2223,N_1505,N_1195);
nor U2224 (N_2224,N_1358,N_1723);
and U2225 (N_2225,N_1833,N_1524);
nand U2226 (N_2226,N_1480,N_1402);
and U2227 (N_2227,N_1829,N_1278);
and U2228 (N_2228,N_1319,N_1741);
nand U2229 (N_2229,N_1333,N_1885);
nand U2230 (N_2230,N_1863,N_1765);
and U2231 (N_2231,N_1537,N_1612);
and U2232 (N_2232,N_1639,N_1099);
or U2233 (N_2233,N_1932,N_1976);
nand U2234 (N_2234,N_1031,N_1499);
or U2235 (N_2235,N_1824,N_1032);
xor U2236 (N_2236,N_1694,N_1249);
and U2237 (N_2237,N_1948,N_1913);
or U2238 (N_2238,N_1525,N_1157);
or U2239 (N_2239,N_1784,N_1602);
nand U2240 (N_2240,N_1097,N_1273);
nand U2241 (N_2241,N_1697,N_1900);
nand U2242 (N_2242,N_1448,N_1445);
xnor U2243 (N_2243,N_1346,N_1670);
and U2244 (N_2244,N_1294,N_1541);
nand U2245 (N_2245,N_1187,N_1513);
or U2246 (N_2246,N_1119,N_1312);
xnor U2247 (N_2247,N_1578,N_1236);
nor U2248 (N_2248,N_1727,N_1328);
or U2249 (N_2249,N_1009,N_1446);
nand U2250 (N_2250,N_1209,N_1387);
nor U2251 (N_2251,N_1039,N_1748);
nand U2252 (N_2252,N_1571,N_1929);
and U2253 (N_2253,N_1515,N_1739);
xor U2254 (N_2254,N_1603,N_1361);
or U2255 (N_2255,N_1804,N_1020);
nor U2256 (N_2256,N_1664,N_1860);
xor U2257 (N_2257,N_1404,N_1820);
nor U2258 (N_2258,N_1374,N_1432);
or U2259 (N_2259,N_1200,N_1871);
and U2260 (N_2260,N_1934,N_1794);
nand U2261 (N_2261,N_1313,N_1855);
nand U2262 (N_2262,N_1685,N_1754);
and U2263 (N_2263,N_1950,N_1917);
nor U2264 (N_2264,N_1325,N_1592);
nand U2265 (N_2265,N_1893,N_1735);
nand U2266 (N_2266,N_1465,N_1813);
or U2267 (N_2267,N_1904,N_1191);
nand U2268 (N_2268,N_1890,N_1609);
and U2269 (N_2269,N_1865,N_1271);
and U2270 (N_2270,N_1546,N_1951);
nand U2271 (N_2271,N_1075,N_1433);
and U2272 (N_2272,N_1768,N_1771);
nand U2273 (N_2273,N_1700,N_1596);
and U2274 (N_2274,N_1128,N_1730);
nor U2275 (N_2275,N_1172,N_1938);
xnor U2276 (N_2276,N_1743,N_1171);
nand U2277 (N_2277,N_1810,N_1014);
or U2278 (N_2278,N_1682,N_1800);
nand U2279 (N_2279,N_1591,N_1665);
xor U2280 (N_2280,N_1693,N_1517);
nand U2281 (N_2281,N_1565,N_1162);
and U2282 (N_2282,N_1710,N_1220);
xor U2283 (N_2283,N_1558,N_1438);
and U2284 (N_2284,N_1615,N_1528);
xor U2285 (N_2285,N_1827,N_1206);
or U2286 (N_2286,N_1047,N_1002);
xnor U2287 (N_2287,N_1241,N_1626);
or U2288 (N_2288,N_1042,N_1543);
nand U2289 (N_2289,N_1698,N_1388);
xnor U2290 (N_2290,N_1169,N_1675);
nand U2291 (N_2291,N_1212,N_1081);
nand U2292 (N_2292,N_1225,N_1949);
or U2293 (N_2293,N_1113,N_1345);
and U2294 (N_2294,N_1668,N_1981);
xnor U2295 (N_2295,N_1629,N_1786);
or U2296 (N_2296,N_1368,N_1208);
or U2297 (N_2297,N_1056,N_1958);
and U2298 (N_2298,N_1906,N_1593);
nand U2299 (N_2299,N_1403,N_1676);
nand U2300 (N_2300,N_1582,N_1848);
nand U2301 (N_2301,N_1005,N_1430);
and U2302 (N_2302,N_1338,N_1666);
or U2303 (N_2303,N_1422,N_1570);
or U2304 (N_2304,N_1192,N_1636);
xor U2305 (N_2305,N_1287,N_1984);
nand U2306 (N_2306,N_1289,N_1673);
nor U2307 (N_2307,N_1144,N_1716);
xor U2308 (N_2308,N_1809,N_1424);
and U2309 (N_2309,N_1542,N_1930);
nand U2310 (N_2310,N_1196,N_1167);
or U2311 (N_2311,N_1715,N_1617);
nor U2312 (N_2312,N_1717,N_1585);
or U2313 (N_2313,N_1922,N_1003);
nand U2314 (N_2314,N_1243,N_1711);
xnor U2315 (N_2315,N_1780,N_1466);
and U2316 (N_2316,N_1892,N_1007);
and U2317 (N_2317,N_1111,N_1080);
and U2318 (N_2318,N_1019,N_1299);
and U2319 (N_2319,N_1400,N_1507);
nor U2320 (N_2320,N_1038,N_1087);
or U2321 (N_2321,N_1254,N_1649);
xor U2322 (N_2322,N_1152,N_1899);
and U2323 (N_2323,N_1376,N_1661);
or U2324 (N_2324,N_1866,N_1782);
and U2325 (N_2325,N_1551,N_1481);
nand U2326 (N_2326,N_1832,N_1691);
and U2327 (N_2327,N_1459,N_1153);
nor U2328 (N_2328,N_1151,N_1344);
xnor U2329 (N_2329,N_1357,N_1696);
nor U2330 (N_2330,N_1405,N_1607);
and U2331 (N_2331,N_1749,N_1015);
nand U2332 (N_2332,N_1064,N_1041);
and U2333 (N_2333,N_1549,N_1048);
nand U2334 (N_2334,N_1872,N_1078);
or U2335 (N_2335,N_1920,N_1889);
nor U2336 (N_2336,N_1261,N_1575);
xor U2337 (N_2337,N_1463,N_1124);
or U2338 (N_2338,N_1781,N_1637);
xnor U2339 (N_2339,N_1747,N_1412);
and U2340 (N_2340,N_1028,N_1252);
nand U2341 (N_2341,N_1907,N_1767);
nor U2342 (N_2342,N_1795,N_1621);
xnor U2343 (N_2343,N_1503,N_1772);
xor U2344 (N_2344,N_1419,N_1122);
xnor U2345 (N_2345,N_1514,N_1447);
nand U2346 (N_2346,N_1941,N_1811);
nand U2347 (N_2347,N_1630,N_1724);
and U2348 (N_2348,N_1761,N_1721);
nand U2349 (N_2349,N_1994,N_1103);
xnor U2350 (N_2350,N_1237,N_1024);
or U2351 (N_2351,N_1112,N_1681);
nand U2352 (N_2352,N_1722,N_1441);
nand U2353 (N_2353,N_1774,N_1061);
nand U2354 (N_2354,N_1588,N_1764);
or U2355 (N_2355,N_1792,N_1548);
nand U2356 (N_2356,N_1168,N_1282);
nor U2357 (N_2357,N_1340,N_1883);
and U2358 (N_2358,N_1655,N_1280);
nand U2359 (N_2359,N_1431,N_1678);
xnor U2360 (N_2360,N_1453,N_1785);
nor U2361 (N_2361,N_1420,N_1506);
nor U2362 (N_2362,N_1652,N_1775);
and U2363 (N_2363,N_1356,N_1518);
nand U2364 (N_2364,N_1182,N_1352);
or U2365 (N_2365,N_1335,N_1536);
nor U2366 (N_2366,N_1132,N_1672);
xor U2367 (N_2367,N_1276,N_1509);
and U2368 (N_2368,N_1109,N_1131);
xor U2369 (N_2369,N_1240,N_1653);
nor U2370 (N_2370,N_1135,N_1527);
or U2371 (N_2371,N_1776,N_1779);
nand U2372 (N_2372,N_1918,N_1671);
or U2373 (N_2373,N_1451,N_1523);
nor U2374 (N_2374,N_1033,N_1560);
and U2375 (N_2375,N_1842,N_1142);
and U2376 (N_2376,N_1291,N_1170);
or U2377 (N_2377,N_1201,N_1973);
or U2378 (N_2378,N_1443,N_1538);
xor U2379 (N_2379,N_1474,N_1628);
xor U2380 (N_2380,N_1742,N_1576);
nor U2381 (N_2381,N_1916,N_1910);
xnor U2382 (N_2382,N_1584,N_1849);
xor U2383 (N_2383,N_1923,N_1566);
or U2384 (N_2384,N_1158,N_1969);
nor U2385 (N_2385,N_1216,N_1107);
xnor U2386 (N_2386,N_1473,N_1213);
nand U2387 (N_2387,N_1699,N_1669);
xnor U2388 (N_2388,N_1018,N_1942);
xnor U2389 (N_2389,N_1010,N_1605);
or U2390 (N_2390,N_1148,N_1369);
and U2391 (N_2391,N_1719,N_1326);
nor U2392 (N_2392,N_1439,N_1380);
nor U2393 (N_2393,N_1349,N_1224);
xor U2394 (N_2394,N_1750,N_1854);
or U2395 (N_2395,N_1440,N_1519);
nor U2396 (N_2396,N_1884,N_1248);
and U2397 (N_2397,N_1687,N_1705);
or U2398 (N_2398,N_1529,N_1778);
xor U2399 (N_2399,N_1016,N_1211);
nor U2400 (N_2400,N_1186,N_1188);
nand U2401 (N_2401,N_1207,N_1911);
or U2402 (N_2402,N_1076,N_1622);
xnor U2403 (N_2403,N_1160,N_1752);
and U2404 (N_2404,N_1631,N_1229);
and U2405 (N_2405,N_1274,N_1350);
nand U2406 (N_2406,N_1580,N_1074);
xor U2407 (N_2407,N_1987,N_1970);
nand U2408 (N_2408,N_1058,N_1413);
or U2409 (N_2409,N_1483,N_1051);
nand U2410 (N_2410,N_1539,N_1791);
xor U2411 (N_2411,N_1022,N_1989);
or U2412 (N_2412,N_1875,N_1288);
nor U2413 (N_2413,N_1083,N_1370);
xnor U2414 (N_2414,N_1259,N_1017);
nand U2415 (N_2415,N_1316,N_1857);
and U2416 (N_2416,N_1914,N_1159);
nor U2417 (N_2417,N_1894,N_1138);
nor U2418 (N_2418,N_1864,N_1647);
xnor U2419 (N_2419,N_1909,N_1125);
nor U2420 (N_2420,N_1086,N_1856);
or U2421 (N_2421,N_1868,N_1819);
nor U2422 (N_2422,N_1242,N_1354);
xnor U2423 (N_2423,N_1486,N_1247);
or U2424 (N_2424,N_1547,N_1695);
and U2425 (N_2425,N_1073,N_1436);
nor U2426 (N_2426,N_1895,N_1608);
nor U2427 (N_2427,N_1726,N_1978);
nor U2428 (N_2428,N_1279,N_1654);
or U2429 (N_2429,N_1762,N_1725);
nand U2430 (N_2430,N_1579,N_1226);
nand U2431 (N_2431,N_1348,N_1199);
nand U2432 (N_2432,N_1807,N_1050);
and U2433 (N_2433,N_1090,N_1120);
nor U2434 (N_2434,N_1787,N_1563);
and U2435 (N_2435,N_1437,N_1692);
xnor U2436 (N_2436,N_1789,N_1903);
xnor U2437 (N_2437,N_1373,N_1219);
nand U2438 (N_2438,N_1146,N_1334);
and U2439 (N_2439,N_1646,N_1258);
or U2440 (N_2440,N_1759,N_1184);
or U2441 (N_2441,N_1365,N_1601);
xnor U2442 (N_2442,N_1834,N_1337);
nand U2443 (N_2443,N_1953,N_1174);
nand U2444 (N_2444,N_1189,N_1475);
or U2445 (N_2445,N_1732,N_1177);
or U2446 (N_2446,N_1572,N_1858);
xor U2447 (N_2447,N_1882,N_1263);
and U2448 (N_2448,N_1996,N_1643);
nor U2449 (N_2449,N_1045,N_1766);
or U2450 (N_2450,N_1301,N_1708);
or U2451 (N_2451,N_1946,N_1260);
xor U2452 (N_2452,N_1392,N_1971);
nand U2453 (N_2453,N_1004,N_1760);
or U2454 (N_2454,N_1096,N_1847);
xor U2455 (N_2455,N_1079,N_1511);
nor U2456 (N_2456,N_1478,N_1840);
nand U2457 (N_2457,N_1846,N_1555);
nor U2458 (N_2458,N_1886,N_1960);
nor U2459 (N_2459,N_1452,N_1943);
nand U2460 (N_2460,N_1979,N_1902);
nor U2461 (N_2461,N_1712,N_1604);
or U2462 (N_2462,N_1485,N_1616);
nand U2463 (N_2463,N_1397,N_1877);
nor U2464 (N_2464,N_1305,N_1729);
nand U2465 (N_2465,N_1395,N_1416);
or U2466 (N_2466,N_1302,N_1036);
and U2467 (N_2467,N_1072,N_1825);
xnor U2468 (N_2468,N_1472,N_1460);
or U2469 (N_2469,N_1961,N_1067);
and U2470 (N_2470,N_1309,N_1550);
xor U2471 (N_2471,N_1822,N_1130);
and U2472 (N_2472,N_1385,N_1836);
or U2473 (N_2473,N_1308,N_1797);
nor U2474 (N_2474,N_1852,N_1901);
xnor U2475 (N_2475,N_1470,N_1085);
or U2476 (N_2476,N_1744,N_1633);
and U2477 (N_2477,N_1059,N_1954);
nor U2478 (N_2478,N_1077,N_1383);
xnor U2479 (N_2479,N_1411,N_1194);
and U2480 (N_2480,N_1642,N_1324);
xor U2481 (N_2481,N_1925,N_1053);
and U2482 (N_2482,N_1110,N_1594);
or U2483 (N_2483,N_1736,N_1844);
nor U2484 (N_2484,N_1025,N_1477);
xor U2485 (N_2485,N_1262,N_1707);
or U2486 (N_2486,N_1428,N_1522);
nor U2487 (N_2487,N_1070,N_1838);
nand U2488 (N_2488,N_1534,N_1126);
and U2489 (N_2489,N_1391,N_1897);
nor U2490 (N_2490,N_1702,N_1627);
xnor U2491 (N_2491,N_1140,N_1330);
xor U2492 (N_2492,N_1867,N_1553);
nor U2493 (N_2493,N_1713,N_1915);
nand U2494 (N_2494,N_1406,N_1618);
xnor U2495 (N_2495,N_1957,N_1035);
xnor U2496 (N_2496,N_1952,N_1658);
nor U2497 (N_2497,N_1251,N_1986);
or U2498 (N_2498,N_1442,N_1175);
nor U2499 (N_2499,N_1281,N_1870);
nand U2500 (N_2500,N_1655,N_1253);
or U2501 (N_2501,N_1706,N_1511);
nand U2502 (N_2502,N_1140,N_1419);
nand U2503 (N_2503,N_1217,N_1783);
or U2504 (N_2504,N_1160,N_1054);
nor U2505 (N_2505,N_1621,N_1253);
xor U2506 (N_2506,N_1274,N_1367);
nor U2507 (N_2507,N_1977,N_1067);
xor U2508 (N_2508,N_1245,N_1075);
nor U2509 (N_2509,N_1844,N_1871);
and U2510 (N_2510,N_1442,N_1492);
xor U2511 (N_2511,N_1296,N_1376);
or U2512 (N_2512,N_1883,N_1685);
or U2513 (N_2513,N_1697,N_1040);
nand U2514 (N_2514,N_1420,N_1906);
nand U2515 (N_2515,N_1867,N_1402);
or U2516 (N_2516,N_1569,N_1882);
nand U2517 (N_2517,N_1823,N_1406);
and U2518 (N_2518,N_1677,N_1151);
xor U2519 (N_2519,N_1579,N_1084);
and U2520 (N_2520,N_1961,N_1782);
nand U2521 (N_2521,N_1161,N_1580);
or U2522 (N_2522,N_1752,N_1309);
xor U2523 (N_2523,N_1122,N_1150);
xor U2524 (N_2524,N_1079,N_1368);
and U2525 (N_2525,N_1620,N_1586);
nand U2526 (N_2526,N_1915,N_1670);
or U2527 (N_2527,N_1385,N_1088);
xnor U2528 (N_2528,N_1408,N_1039);
xnor U2529 (N_2529,N_1270,N_1371);
nand U2530 (N_2530,N_1142,N_1057);
xnor U2531 (N_2531,N_1366,N_1956);
and U2532 (N_2532,N_1023,N_1583);
or U2533 (N_2533,N_1606,N_1103);
nor U2534 (N_2534,N_1489,N_1975);
nand U2535 (N_2535,N_1900,N_1466);
xnor U2536 (N_2536,N_1045,N_1881);
or U2537 (N_2537,N_1861,N_1828);
nor U2538 (N_2538,N_1428,N_1983);
and U2539 (N_2539,N_1547,N_1541);
or U2540 (N_2540,N_1782,N_1293);
and U2541 (N_2541,N_1535,N_1286);
nand U2542 (N_2542,N_1541,N_1649);
or U2543 (N_2543,N_1512,N_1256);
xor U2544 (N_2544,N_1697,N_1936);
or U2545 (N_2545,N_1610,N_1724);
nor U2546 (N_2546,N_1158,N_1102);
nand U2547 (N_2547,N_1063,N_1481);
or U2548 (N_2548,N_1072,N_1416);
and U2549 (N_2549,N_1050,N_1655);
nor U2550 (N_2550,N_1518,N_1505);
xor U2551 (N_2551,N_1749,N_1049);
and U2552 (N_2552,N_1294,N_1288);
and U2553 (N_2553,N_1848,N_1488);
or U2554 (N_2554,N_1160,N_1498);
xor U2555 (N_2555,N_1531,N_1623);
nor U2556 (N_2556,N_1482,N_1283);
nand U2557 (N_2557,N_1824,N_1734);
and U2558 (N_2558,N_1520,N_1231);
xor U2559 (N_2559,N_1020,N_1381);
nand U2560 (N_2560,N_1711,N_1370);
nand U2561 (N_2561,N_1388,N_1975);
or U2562 (N_2562,N_1988,N_1552);
and U2563 (N_2563,N_1117,N_1267);
nand U2564 (N_2564,N_1074,N_1677);
xnor U2565 (N_2565,N_1673,N_1113);
xnor U2566 (N_2566,N_1477,N_1903);
and U2567 (N_2567,N_1668,N_1321);
nor U2568 (N_2568,N_1014,N_1410);
nand U2569 (N_2569,N_1620,N_1961);
or U2570 (N_2570,N_1466,N_1213);
or U2571 (N_2571,N_1160,N_1394);
nor U2572 (N_2572,N_1917,N_1979);
xor U2573 (N_2573,N_1783,N_1711);
nand U2574 (N_2574,N_1098,N_1000);
nor U2575 (N_2575,N_1967,N_1324);
xor U2576 (N_2576,N_1805,N_1288);
and U2577 (N_2577,N_1867,N_1182);
and U2578 (N_2578,N_1712,N_1811);
nor U2579 (N_2579,N_1112,N_1090);
and U2580 (N_2580,N_1670,N_1554);
and U2581 (N_2581,N_1737,N_1324);
or U2582 (N_2582,N_1704,N_1682);
nor U2583 (N_2583,N_1211,N_1495);
nor U2584 (N_2584,N_1967,N_1857);
or U2585 (N_2585,N_1066,N_1676);
nand U2586 (N_2586,N_1140,N_1216);
nand U2587 (N_2587,N_1836,N_1947);
nand U2588 (N_2588,N_1620,N_1450);
and U2589 (N_2589,N_1662,N_1473);
nor U2590 (N_2590,N_1577,N_1817);
or U2591 (N_2591,N_1713,N_1377);
nor U2592 (N_2592,N_1615,N_1091);
nor U2593 (N_2593,N_1701,N_1824);
xnor U2594 (N_2594,N_1751,N_1386);
or U2595 (N_2595,N_1279,N_1591);
nand U2596 (N_2596,N_1432,N_1473);
and U2597 (N_2597,N_1704,N_1792);
nand U2598 (N_2598,N_1285,N_1919);
xor U2599 (N_2599,N_1753,N_1994);
nand U2600 (N_2600,N_1330,N_1813);
nor U2601 (N_2601,N_1782,N_1710);
and U2602 (N_2602,N_1667,N_1947);
and U2603 (N_2603,N_1492,N_1560);
and U2604 (N_2604,N_1454,N_1959);
xor U2605 (N_2605,N_1281,N_1752);
xor U2606 (N_2606,N_1989,N_1202);
nand U2607 (N_2607,N_1968,N_1301);
nor U2608 (N_2608,N_1049,N_1097);
and U2609 (N_2609,N_1974,N_1814);
nor U2610 (N_2610,N_1326,N_1674);
and U2611 (N_2611,N_1263,N_1955);
or U2612 (N_2612,N_1859,N_1626);
nor U2613 (N_2613,N_1233,N_1624);
and U2614 (N_2614,N_1454,N_1455);
xnor U2615 (N_2615,N_1563,N_1717);
nor U2616 (N_2616,N_1007,N_1631);
and U2617 (N_2617,N_1978,N_1081);
or U2618 (N_2618,N_1990,N_1819);
nand U2619 (N_2619,N_1022,N_1787);
nand U2620 (N_2620,N_1231,N_1889);
and U2621 (N_2621,N_1837,N_1688);
nand U2622 (N_2622,N_1223,N_1266);
or U2623 (N_2623,N_1018,N_1190);
xor U2624 (N_2624,N_1784,N_1923);
xnor U2625 (N_2625,N_1204,N_1105);
nor U2626 (N_2626,N_1180,N_1892);
or U2627 (N_2627,N_1738,N_1946);
and U2628 (N_2628,N_1753,N_1648);
xnor U2629 (N_2629,N_1981,N_1190);
nand U2630 (N_2630,N_1051,N_1307);
or U2631 (N_2631,N_1128,N_1356);
xnor U2632 (N_2632,N_1409,N_1086);
xor U2633 (N_2633,N_1366,N_1859);
nor U2634 (N_2634,N_1244,N_1739);
nor U2635 (N_2635,N_1913,N_1004);
xor U2636 (N_2636,N_1354,N_1228);
nand U2637 (N_2637,N_1652,N_1894);
and U2638 (N_2638,N_1856,N_1943);
and U2639 (N_2639,N_1436,N_1547);
and U2640 (N_2640,N_1375,N_1777);
and U2641 (N_2641,N_1105,N_1133);
nand U2642 (N_2642,N_1837,N_1289);
nor U2643 (N_2643,N_1212,N_1868);
nand U2644 (N_2644,N_1831,N_1751);
xor U2645 (N_2645,N_1806,N_1472);
or U2646 (N_2646,N_1587,N_1055);
xnor U2647 (N_2647,N_1819,N_1376);
or U2648 (N_2648,N_1961,N_1888);
nor U2649 (N_2649,N_1792,N_1135);
or U2650 (N_2650,N_1511,N_1806);
nand U2651 (N_2651,N_1082,N_1467);
or U2652 (N_2652,N_1712,N_1899);
nor U2653 (N_2653,N_1823,N_1453);
or U2654 (N_2654,N_1068,N_1919);
nand U2655 (N_2655,N_1441,N_1041);
and U2656 (N_2656,N_1700,N_1309);
and U2657 (N_2657,N_1141,N_1117);
and U2658 (N_2658,N_1051,N_1479);
xor U2659 (N_2659,N_1013,N_1761);
and U2660 (N_2660,N_1552,N_1709);
nand U2661 (N_2661,N_1025,N_1349);
nor U2662 (N_2662,N_1451,N_1022);
or U2663 (N_2663,N_1640,N_1451);
and U2664 (N_2664,N_1484,N_1040);
and U2665 (N_2665,N_1601,N_1670);
and U2666 (N_2666,N_1670,N_1772);
nand U2667 (N_2667,N_1830,N_1063);
and U2668 (N_2668,N_1843,N_1487);
and U2669 (N_2669,N_1759,N_1553);
xor U2670 (N_2670,N_1058,N_1374);
xor U2671 (N_2671,N_1308,N_1780);
nand U2672 (N_2672,N_1489,N_1588);
nor U2673 (N_2673,N_1024,N_1971);
or U2674 (N_2674,N_1108,N_1736);
nor U2675 (N_2675,N_1163,N_1366);
or U2676 (N_2676,N_1700,N_1918);
nor U2677 (N_2677,N_1295,N_1080);
xor U2678 (N_2678,N_1604,N_1472);
and U2679 (N_2679,N_1471,N_1614);
nor U2680 (N_2680,N_1262,N_1265);
nand U2681 (N_2681,N_1427,N_1097);
and U2682 (N_2682,N_1327,N_1827);
xnor U2683 (N_2683,N_1953,N_1354);
nand U2684 (N_2684,N_1765,N_1361);
xnor U2685 (N_2685,N_1822,N_1909);
and U2686 (N_2686,N_1262,N_1833);
or U2687 (N_2687,N_1227,N_1896);
xor U2688 (N_2688,N_1876,N_1307);
and U2689 (N_2689,N_1691,N_1488);
and U2690 (N_2690,N_1942,N_1258);
nand U2691 (N_2691,N_1056,N_1427);
xor U2692 (N_2692,N_1603,N_1919);
nor U2693 (N_2693,N_1859,N_1531);
or U2694 (N_2694,N_1348,N_1016);
xor U2695 (N_2695,N_1659,N_1071);
nor U2696 (N_2696,N_1873,N_1930);
nor U2697 (N_2697,N_1244,N_1127);
nand U2698 (N_2698,N_1552,N_1321);
nand U2699 (N_2699,N_1089,N_1047);
and U2700 (N_2700,N_1580,N_1834);
xnor U2701 (N_2701,N_1799,N_1235);
xnor U2702 (N_2702,N_1109,N_1289);
nor U2703 (N_2703,N_1407,N_1503);
nor U2704 (N_2704,N_1062,N_1464);
or U2705 (N_2705,N_1743,N_1930);
xor U2706 (N_2706,N_1621,N_1850);
or U2707 (N_2707,N_1605,N_1564);
nand U2708 (N_2708,N_1050,N_1716);
or U2709 (N_2709,N_1875,N_1109);
nand U2710 (N_2710,N_1328,N_1190);
nand U2711 (N_2711,N_1508,N_1093);
or U2712 (N_2712,N_1030,N_1991);
or U2713 (N_2713,N_1301,N_1761);
nor U2714 (N_2714,N_1753,N_1863);
nor U2715 (N_2715,N_1896,N_1053);
xnor U2716 (N_2716,N_1936,N_1119);
nand U2717 (N_2717,N_1988,N_1567);
xnor U2718 (N_2718,N_1796,N_1098);
nor U2719 (N_2719,N_1761,N_1609);
or U2720 (N_2720,N_1658,N_1221);
nor U2721 (N_2721,N_1492,N_1833);
or U2722 (N_2722,N_1433,N_1495);
xor U2723 (N_2723,N_1189,N_1270);
nor U2724 (N_2724,N_1336,N_1023);
nor U2725 (N_2725,N_1415,N_1090);
nor U2726 (N_2726,N_1550,N_1473);
nor U2727 (N_2727,N_1822,N_1277);
or U2728 (N_2728,N_1292,N_1346);
or U2729 (N_2729,N_1300,N_1319);
nand U2730 (N_2730,N_1366,N_1986);
nor U2731 (N_2731,N_1891,N_1404);
nor U2732 (N_2732,N_1678,N_1413);
or U2733 (N_2733,N_1305,N_1860);
and U2734 (N_2734,N_1876,N_1979);
nor U2735 (N_2735,N_1684,N_1012);
and U2736 (N_2736,N_1996,N_1188);
or U2737 (N_2737,N_1226,N_1032);
nor U2738 (N_2738,N_1752,N_1239);
nor U2739 (N_2739,N_1108,N_1937);
nand U2740 (N_2740,N_1662,N_1377);
xnor U2741 (N_2741,N_1829,N_1582);
or U2742 (N_2742,N_1352,N_1194);
or U2743 (N_2743,N_1736,N_1620);
and U2744 (N_2744,N_1758,N_1917);
and U2745 (N_2745,N_1216,N_1384);
nand U2746 (N_2746,N_1689,N_1557);
nor U2747 (N_2747,N_1458,N_1469);
and U2748 (N_2748,N_1670,N_1928);
and U2749 (N_2749,N_1372,N_1835);
and U2750 (N_2750,N_1573,N_1455);
and U2751 (N_2751,N_1447,N_1436);
xnor U2752 (N_2752,N_1970,N_1052);
xnor U2753 (N_2753,N_1034,N_1208);
nand U2754 (N_2754,N_1960,N_1311);
nor U2755 (N_2755,N_1601,N_1343);
or U2756 (N_2756,N_1642,N_1678);
or U2757 (N_2757,N_1712,N_1275);
nor U2758 (N_2758,N_1847,N_1623);
nand U2759 (N_2759,N_1051,N_1887);
and U2760 (N_2760,N_1045,N_1787);
nand U2761 (N_2761,N_1932,N_1420);
nand U2762 (N_2762,N_1912,N_1775);
and U2763 (N_2763,N_1111,N_1318);
nand U2764 (N_2764,N_1695,N_1414);
nand U2765 (N_2765,N_1299,N_1783);
xor U2766 (N_2766,N_1966,N_1943);
nor U2767 (N_2767,N_1781,N_1622);
or U2768 (N_2768,N_1612,N_1753);
nor U2769 (N_2769,N_1792,N_1845);
xnor U2770 (N_2770,N_1518,N_1942);
and U2771 (N_2771,N_1641,N_1690);
and U2772 (N_2772,N_1335,N_1526);
or U2773 (N_2773,N_1506,N_1543);
nand U2774 (N_2774,N_1171,N_1386);
and U2775 (N_2775,N_1498,N_1769);
or U2776 (N_2776,N_1308,N_1983);
or U2777 (N_2777,N_1064,N_1047);
and U2778 (N_2778,N_1507,N_1755);
or U2779 (N_2779,N_1272,N_1421);
nor U2780 (N_2780,N_1847,N_1686);
and U2781 (N_2781,N_1878,N_1580);
xnor U2782 (N_2782,N_1765,N_1094);
and U2783 (N_2783,N_1652,N_1439);
or U2784 (N_2784,N_1046,N_1360);
and U2785 (N_2785,N_1966,N_1119);
nand U2786 (N_2786,N_1762,N_1479);
xnor U2787 (N_2787,N_1742,N_1662);
nand U2788 (N_2788,N_1472,N_1851);
or U2789 (N_2789,N_1306,N_1128);
nand U2790 (N_2790,N_1304,N_1590);
nand U2791 (N_2791,N_1637,N_1570);
and U2792 (N_2792,N_1954,N_1219);
nor U2793 (N_2793,N_1387,N_1042);
nor U2794 (N_2794,N_1467,N_1176);
nand U2795 (N_2795,N_1476,N_1283);
xor U2796 (N_2796,N_1302,N_1712);
nor U2797 (N_2797,N_1742,N_1364);
nor U2798 (N_2798,N_1499,N_1586);
and U2799 (N_2799,N_1848,N_1056);
nand U2800 (N_2800,N_1273,N_1751);
nand U2801 (N_2801,N_1528,N_1040);
and U2802 (N_2802,N_1898,N_1791);
xor U2803 (N_2803,N_1124,N_1707);
or U2804 (N_2804,N_1083,N_1642);
nor U2805 (N_2805,N_1481,N_1494);
and U2806 (N_2806,N_1840,N_1690);
or U2807 (N_2807,N_1566,N_1351);
xor U2808 (N_2808,N_1225,N_1009);
or U2809 (N_2809,N_1479,N_1101);
or U2810 (N_2810,N_1276,N_1210);
nor U2811 (N_2811,N_1761,N_1451);
nand U2812 (N_2812,N_1218,N_1579);
and U2813 (N_2813,N_1080,N_1396);
nand U2814 (N_2814,N_1854,N_1312);
nand U2815 (N_2815,N_1856,N_1183);
xnor U2816 (N_2816,N_1828,N_1598);
xor U2817 (N_2817,N_1090,N_1769);
and U2818 (N_2818,N_1089,N_1673);
xnor U2819 (N_2819,N_1245,N_1199);
and U2820 (N_2820,N_1625,N_1346);
xnor U2821 (N_2821,N_1404,N_1760);
nand U2822 (N_2822,N_1523,N_1594);
xnor U2823 (N_2823,N_1394,N_1528);
or U2824 (N_2824,N_1615,N_1086);
xor U2825 (N_2825,N_1787,N_1455);
xnor U2826 (N_2826,N_1971,N_1277);
nand U2827 (N_2827,N_1310,N_1647);
xnor U2828 (N_2828,N_1650,N_1595);
nor U2829 (N_2829,N_1928,N_1097);
and U2830 (N_2830,N_1745,N_1599);
nand U2831 (N_2831,N_1889,N_1315);
or U2832 (N_2832,N_1320,N_1852);
xor U2833 (N_2833,N_1567,N_1843);
and U2834 (N_2834,N_1856,N_1997);
nand U2835 (N_2835,N_1745,N_1513);
nand U2836 (N_2836,N_1707,N_1947);
xor U2837 (N_2837,N_1212,N_1683);
xor U2838 (N_2838,N_1361,N_1057);
nor U2839 (N_2839,N_1614,N_1347);
xor U2840 (N_2840,N_1160,N_1565);
nand U2841 (N_2841,N_1505,N_1934);
nand U2842 (N_2842,N_1131,N_1044);
nand U2843 (N_2843,N_1563,N_1776);
xor U2844 (N_2844,N_1909,N_1756);
or U2845 (N_2845,N_1191,N_1083);
xor U2846 (N_2846,N_1931,N_1437);
xor U2847 (N_2847,N_1028,N_1448);
nor U2848 (N_2848,N_1568,N_1692);
xor U2849 (N_2849,N_1313,N_1271);
and U2850 (N_2850,N_1172,N_1548);
nand U2851 (N_2851,N_1130,N_1596);
or U2852 (N_2852,N_1785,N_1987);
xor U2853 (N_2853,N_1732,N_1841);
or U2854 (N_2854,N_1769,N_1639);
nor U2855 (N_2855,N_1273,N_1289);
and U2856 (N_2856,N_1717,N_1397);
xor U2857 (N_2857,N_1821,N_1743);
xor U2858 (N_2858,N_1682,N_1783);
and U2859 (N_2859,N_1715,N_1151);
nand U2860 (N_2860,N_1968,N_1185);
or U2861 (N_2861,N_1940,N_1722);
xor U2862 (N_2862,N_1634,N_1415);
xnor U2863 (N_2863,N_1496,N_1292);
nor U2864 (N_2864,N_1142,N_1359);
or U2865 (N_2865,N_1185,N_1757);
and U2866 (N_2866,N_1215,N_1259);
nand U2867 (N_2867,N_1391,N_1457);
or U2868 (N_2868,N_1313,N_1038);
nor U2869 (N_2869,N_1296,N_1282);
and U2870 (N_2870,N_1163,N_1713);
or U2871 (N_2871,N_1330,N_1772);
and U2872 (N_2872,N_1403,N_1098);
xnor U2873 (N_2873,N_1748,N_1686);
or U2874 (N_2874,N_1099,N_1772);
nor U2875 (N_2875,N_1521,N_1810);
and U2876 (N_2876,N_1002,N_1933);
nor U2877 (N_2877,N_1310,N_1338);
nor U2878 (N_2878,N_1928,N_1448);
nand U2879 (N_2879,N_1079,N_1437);
and U2880 (N_2880,N_1281,N_1275);
nor U2881 (N_2881,N_1735,N_1946);
nand U2882 (N_2882,N_1775,N_1679);
nand U2883 (N_2883,N_1013,N_1216);
nand U2884 (N_2884,N_1848,N_1527);
nor U2885 (N_2885,N_1214,N_1712);
or U2886 (N_2886,N_1925,N_1344);
or U2887 (N_2887,N_1945,N_1580);
nand U2888 (N_2888,N_1200,N_1663);
xor U2889 (N_2889,N_1725,N_1620);
nand U2890 (N_2890,N_1598,N_1849);
nor U2891 (N_2891,N_1294,N_1434);
and U2892 (N_2892,N_1798,N_1388);
or U2893 (N_2893,N_1260,N_1492);
nor U2894 (N_2894,N_1868,N_1257);
nor U2895 (N_2895,N_1043,N_1871);
xor U2896 (N_2896,N_1279,N_1716);
nor U2897 (N_2897,N_1639,N_1399);
and U2898 (N_2898,N_1942,N_1615);
and U2899 (N_2899,N_1902,N_1950);
or U2900 (N_2900,N_1807,N_1074);
or U2901 (N_2901,N_1910,N_1233);
nor U2902 (N_2902,N_1297,N_1855);
and U2903 (N_2903,N_1366,N_1129);
and U2904 (N_2904,N_1711,N_1495);
and U2905 (N_2905,N_1751,N_1160);
and U2906 (N_2906,N_1267,N_1447);
nand U2907 (N_2907,N_1272,N_1575);
and U2908 (N_2908,N_1355,N_1590);
or U2909 (N_2909,N_1535,N_1792);
and U2910 (N_2910,N_1227,N_1580);
nor U2911 (N_2911,N_1059,N_1211);
or U2912 (N_2912,N_1295,N_1100);
nand U2913 (N_2913,N_1433,N_1920);
nor U2914 (N_2914,N_1213,N_1190);
and U2915 (N_2915,N_1621,N_1493);
or U2916 (N_2916,N_1401,N_1391);
nand U2917 (N_2917,N_1812,N_1701);
or U2918 (N_2918,N_1023,N_1057);
or U2919 (N_2919,N_1723,N_1652);
and U2920 (N_2920,N_1437,N_1336);
nand U2921 (N_2921,N_1551,N_1649);
and U2922 (N_2922,N_1206,N_1730);
or U2923 (N_2923,N_1374,N_1772);
xor U2924 (N_2924,N_1154,N_1549);
nand U2925 (N_2925,N_1496,N_1736);
xnor U2926 (N_2926,N_1275,N_1663);
nor U2927 (N_2927,N_1744,N_1421);
nor U2928 (N_2928,N_1777,N_1541);
nor U2929 (N_2929,N_1434,N_1195);
and U2930 (N_2930,N_1726,N_1177);
xor U2931 (N_2931,N_1795,N_1476);
nand U2932 (N_2932,N_1432,N_1266);
nand U2933 (N_2933,N_1583,N_1573);
nand U2934 (N_2934,N_1716,N_1443);
xnor U2935 (N_2935,N_1927,N_1220);
nand U2936 (N_2936,N_1663,N_1203);
or U2937 (N_2937,N_1716,N_1559);
nor U2938 (N_2938,N_1838,N_1276);
or U2939 (N_2939,N_1664,N_1122);
xor U2940 (N_2940,N_1839,N_1784);
xor U2941 (N_2941,N_1307,N_1714);
xnor U2942 (N_2942,N_1499,N_1190);
or U2943 (N_2943,N_1762,N_1141);
and U2944 (N_2944,N_1407,N_1823);
and U2945 (N_2945,N_1027,N_1447);
and U2946 (N_2946,N_1559,N_1042);
xor U2947 (N_2947,N_1426,N_1364);
nand U2948 (N_2948,N_1040,N_1191);
nor U2949 (N_2949,N_1633,N_1761);
xnor U2950 (N_2950,N_1627,N_1259);
or U2951 (N_2951,N_1395,N_1029);
nor U2952 (N_2952,N_1632,N_1390);
and U2953 (N_2953,N_1066,N_1481);
nand U2954 (N_2954,N_1319,N_1131);
xnor U2955 (N_2955,N_1514,N_1747);
nor U2956 (N_2956,N_1503,N_1393);
nor U2957 (N_2957,N_1783,N_1822);
xor U2958 (N_2958,N_1860,N_1544);
and U2959 (N_2959,N_1791,N_1799);
and U2960 (N_2960,N_1187,N_1098);
nor U2961 (N_2961,N_1982,N_1849);
and U2962 (N_2962,N_1920,N_1300);
or U2963 (N_2963,N_1355,N_1695);
nand U2964 (N_2964,N_1097,N_1270);
or U2965 (N_2965,N_1223,N_1189);
or U2966 (N_2966,N_1390,N_1158);
nand U2967 (N_2967,N_1569,N_1847);
or U2968 (N_2968,N_1793,N_1486);
or U2969 (N_2969,N_1070,N_1488);
nor U2970 (N_2970,N_1668,N_1647);
nor U2971 (N_2971,N_1068,N_1452);
xor U2972 (N_2972,N_1464,N_1855);
xnor U2973 (N_2973,N_1343,N_1842);
nor U2974 (N_2974,N_1843,N_1801);
xnor U2975 (N_2975,N_1279,N_1570);
and U2976 (N_2976,N_1696,N_1245);
or U2977 (N_2977,N_1126,N_1706);
nand U2978 (N_2978,N_1606,N_1517);
nand U2979 (N_2979,N_1733,N_1080);
nor U2980 (N_2980,N_1733,N_1225);
nand U2981 (N_2981,N_1454,N_1853);
nor U2982 (N_2982,N_1527,N_1897);
xnor U2983 (N_2983,N_1203,N_1138);
xnor U2984 (N_2984,N_1454,N_1144);
nand U2985 (N_2985,N_1373,N_1724);
xor U2986 (N_2986,N_1989,N_1561);
xor U2987 (N_2987,N_1189,N_1513);
xor U2988 (N_2988,N_1375,N_1043);
nand U2989 (N_2989,N_1760,N_1593);
xnor U2990 (N_2990,N_1707,N_1828);
xor U2991 (N_2991,N_1695,N_1872);
and U2992 (N_2992,N_1865,N_1217);
nand U2993 (N_2993,N_1883,N_1406);
or U2994 (N_2994,N_1447,N_1734);
xnor U2995 (N_2995,N_1367,N_1267);
nand U2996 (N_2996,N_1204,N_1490);
nor U2997 (N_2997,N_1365,N_1274);
and U2998 (N_2998,N_1610,N_1988);
and U2999 (N_2999,N_1906,N_1660);
and U3000 (N_3000,N_2218,N_2525);
or U3001 (N_3001,N_2216,N_2959);
xor U3002 (N_3002,N_2887,N_2708);
nand U3003 (N_3003,N_2189,N_2357);
xnor U3004 (N_3004,N_2846,N_2409);
xnor U3005 (N_3005,N_2159,N_2332);
or U3006 (N_3006,N_2283,N_2720);
nand U3007 (N_3007,N_2786,N_2209);
nor U3008 (N_3008,N_2370,N_2680);
nand U3009 (N_3009,N_2125,N_2223);
nand U3010 (N_3010,N_2465,N_2580);
xor U3011 (N_3011,N_2647,N_2324);
nor U3012 (N_3012,N_2183,N_2549);
xnor U3013 (N_3013,N_2514,N_2981);
and U3014 (N_3014,N_2446,N_2163);
and U3015 (N_3015,N_2666,N_2805);
xnor U3016 (N_3016,N_2722,N_2906);
nand U3017 (N_3017,N_2946,N_2936);
xor U3018 (N_3018,N_2962,N_2606);
xnor U3019 (N_3019,N_2900,N_2102);
xnor U3020 (N_3020,N_2149,N_2611);
xnor U3021 (N_3021,N_2562,N_2004);
nor U3022 (N_3022,N_2186,N_2416);
and U3023 (N_3023,N_2875,N_2239);
and U3024 (N_3024,N_2983,N_2062);
xor U3025 (N_3025,N_2152,N_2157);
or U3026 (N_3026,N_2038,N_2025);
or U3027 (N_3027,N_2268,N_2154);
xnor U3028 (N_3028,N_2028,N_2200);
xnor U3029 (N_3029,N_2261,N_2964);
xnor U3030 (N_3030,N_2880,N_2018);
nor U3031 (N_3031,N_2527,N_2941);
nand U3032 (N_3032,N_2459,N_2327);
xor U3033 (N_3033,N_2070,N_2642);
xnor U3034 (N_3034,N_2319,N_2422);
nand U3035 (N_3035,N_2289,N_2818);
and U3036 (N_3036,N_2059,N_2405);
xnor U3037 (N_3037,N_2495,N_2453);
or U3038 (N_3038,N_2292,N_2092);
or U3039 (N_3039,N_2048,N_2248);
nand U3040 (N_3040,N_2584,N_2896);
nand U3041 (N_3041,N_2034,N_2693);
and U3042 (N_3042,N_2010,N_2923);
and U3043 (N_3043,N_2297,N_2651);
nor U3044 (N_3044,N_2762,N_2652);
nor U3045 (N_3045,N_2737,N_2541);
and U3046 (N_3046,N_2576,N_2904);
nor U3047 (N_3047,N_2053,N_2995);
xor U3048 (N_3048,N_2953,N_2756);
and U3049 (N_3049,N_2263,N_2598);
or U3050 (N_3050,N_2379,N_2147);
nor U3051 (N_3051,N_2103,N_2745);
or U3052 (N_3052,N_2661,N_2279);
nand U3053 (N_3053,N_2719,N_2231);
and U3054 (N_3054,N_2350,N_2090);
or U3055 (N_3055,N_2631,N_2041);
nor U3056 (N_3056,N_2412,N_2114);
xor U3057 (N_3057,N_2381,N_2858);
or U3058 (N_3058,N_2456,N_2917);
nor U3059 (N_3059,N_2700,N_2049);
and U3060 (N_3060,N_2692,N_2838);
nor U3061 (N_3061,N_2672,N_2957);
or U3062 (N_3062,N_2391,N_2233);
xor U3063 (N_3063,N_2247,N_2673);
nor U3064 (N_3064,N_2641,N_2027);
xor U3065 (N_3065,N_2222,N_2565);
xnor U3066 (N_3066,N_2921,N_2052);
and U3067 (N_3067,N_2282,N_2307);
nand U3068 (N_3068,N_2488,N_2471);
nor U3069 (N_3069,N_2136,N_2971);
xor U3070 (N_3070,N_2889,N_2039);
nor U3071 (N_3071,N_2354,N_2161);
nand U3072 (N_3072,N_2969,N_2945);
and U3073 (N_3073,N_2940,N_2590);
xnor U3074 (N_3074,N_2717,N_2544);
and U3075 (N_3075,N_2845,N_2822);
nor U3076 (N_3076,N_2710,N_2781);
nand U3077 (N_3077,N_2738,N_2285);
and U3078 (N_3078,N_2996,N_2097);
and U3079 (N_3079,N_2395,N_2006);
nand U3080 (N_3080,N_2654,N_2752);
and U3081 (N_3081,N_2689,N_2131);
or U3082 (N_3082,N_2326,N_2081);
xnor U3083 (N_3083,N_2681,N_2221);
xnor U3084 (N_3084,N_2726,N_2943);
or U3085 (N_3085,N_2920,N_2808);
nand U3086 (N_3086,N_2788,N_2392);
nor U3087 (N_3087,N_2867,N_2898);
or U3088 (N_3088,N_2000,N_2045);
or U3089 (N_3089,N_2688,N_2699);
nand U3090 (N_3090,N_2568,N_2629);
nor U3091 (N_3091,N_2547,N_2540);
nand U3092 (N_3092,N_2009,N_2704);
nor U3093 (N_3093,N_2511,N_2759);
nor U3094 (N_3094,N_2162,N_2691);
xnor U3095 (N_3095,N_2106,N_2952);
or U3096 (N_3096,N_2238,N_2243);
xor U3097 (N_3097,N_2587,N_2093);
and U3098 (N_3098,N_2798,N_2076);
or U3099 (N_3099,N_2548,N_2750);
nand U3100 (N_3100,N_2841,N_2733);
and U3101 (N_3101,N_2922,N_2115);
and U3102 (N_3102,N_2120,N_2634);
xor U3103 (N_3103,N_2833,N_2472);
nor U3104 (N_3104,N_2520,N_2187);
nor U3105 (N_3105,N_2690,N_2742);
and U3106 (N_3106,N_2252,N_2537);
nor U3107 (N_3107,N_2826,N_2344);
nor U3108 (N_3108,N_2551,N_2046);
nand U3109 (N_3109,N_2166,N_2881);
nand U3110 (N_3110,N_2172,N_2653);
xor U3111 (N_3111,N_2208,N_2151);
nand U3112 (N_3112,N_2054,N_2224);
nor U3113 (N_3113,N_2650,N_2776);
xor U3114 (N_3114,N_2408,N_2773);
or U3115 (N_3115,N_2080,N_2335);
xnor U3116 (N_3116,N_2134,N_2473);
nand U3117 (N_3117,N_2813,N_2529);
nor U3118 (N_3118,N_2582,N_2804);
or U3119 (N_3119,N_2740,N_2836);
xor U3120 (N_3120,N_2583,N_2121);
and U3121 (N_3121,N_2491,N_2394);
xor U3122 (N_3122,N_2877,N_2293);
xnor U3123 (N_3123,N_2546,N_2791);
or U3124 (N_3124,N_2948,N_2678);
nor U3125 (N_3125,N_2143,N_2821);
nor U3126 (N_3126,N_2814,N_2104);
and U3127 (N_3127,N_2204,N_2847);
and U3128 (N_3128,N_2315,N_2703);
and U3129 (N_3129,N_2257,N_2866);
or U3130 (N_3130,N_2679,N_2269);
and U3131 (N_3131,N_2277,N_2695);
nor U3132 (N_3132,N_2047,N_2452);
or U3133 (N_3133,N_2621,N_2809);
nor U3134 (N_3134,N_2198,N_2368);
xnor U3135 (N_3135,N_2748,N_2270);
xor U3136 (N_3136,N_2155,N_2974);
or U3137 (N_3137,N_2089,N_2637);
or U3138 (N_3138,N_2366,N_2787);
xnor U3139 (N_3139,N_2526,N_2779);
and U3140 (N_3140,N_2212,N_2980);
nor U3141 (N_3141,N_2184,N_2789);
or U3142 (N_3142,N_2913,N_2158);
or U3143 (N_3143,N_2193,N_2604);
or U3144 (N_3144,N_2066,N_2349);
or U3145 (N_3145,N_2820,N_2723);
nand U3146 (N_3146,N_2398,N_2694);
and U3147 (N_3147,N_2873,N_2073);
xor U3148 (N_3148,N_2591,N_2148);
nor U3149 (N_3149,N_2432,N_2840);
xnor U3150 (N_3150,N_2912,N_2676);
nor U3151 (N_3151,N_2975,N_2663);
xor U3152 (N_3152,N_2572,N_2751);
nor U3153 (N_3153,N_2436,N_2301);
xor U3154 (N_3154,N_2088,N_2188);
nand U3155 (N_3155,N_2618,N_2816);
nor U3156 (N_3156,N_2210,N_2852);
or U3157 (N_3157,N_2949,N_2711);
nor U3158 (N_3158,N_2309,N_2707);
nand U3159 (N_3159,N_2785,N_2244);
and U3160 (N_3160,N_2909,N_2013);
or U3161 (N_3161,N_2298,N_2892);
xnor U3162 (N_3162,N_2829,N_2318);
or U3163 (N_3163,N_2987,N_2145);
xor U3164 (N_3164,N_2918,N_2636);
and U3165 (N_3165,N_2518,N_2643);
and U3166 (N_3166,N_2168,N_2775);
nor U3167 (N_3167,N_2571,N_2734);
or U3168 (N_3168,N_2462,N_2044);
xor U3169 (N_3169,N_2192,N_2296);
and U3170 (N_3170,N_2258,N_2033);
and U3171 (N_3171,N_2560,N_2095);
nand U3172 (N_3172,N_2225,N_2487);
nor U3173 (N_3173,N_2599,N_2492);
or U3174 (N_3174,N_2077,N_2063);
or U3175 (N_3175,N_2245,N_2856);
nand U3176 (N_3176,N_2538,N_2721);
or U3177 (N_3177,N_2729,N_2384);
nor U3178 (N_3178,N_2563,N_2494);
or U3179 (N_3179,N_2294,N_2597);
nand U3180 (N_3180,N_2677,N_2174);
and U3181 (N_3181,N_2988,N_2792);
or U3182 (N_3182,N_2557,N_2659);
xor U3183 (N_3183,N_2992,N_2449);
nor U3184 (N_3184,N_2086,N_2317);
and U3185 (N_3185,N_2763,N_2783);
xor U3186 (N_3186,N_2227,N_2810);
and U3187 (N_3187,N_2303,N_2445);
nor U3188 (N_3188,N_2215,N_2393);
xor U3189 (N_3189,N_2182,N_2954);
xnor U3190 (N_3190,N_2385,N_2242);
nor U3191 (N_3191,N_2128,N_2480);
nand U3192 (N_3192,N_2832,N_2116);
xnor U3193 (N_3193,N_2378,N_2057);
nand U3194 (N_3194,N_2108,N_2891);
or U3195 (N_3195,N_2109,N_2023);
nand U3196 (N_3196,N_2765,N_2612);
nor U3197 (N_3197,N_2955,N_2101);
xnor U3198 (N_3198,N_2633,N_2419);
and U3199 (N_3199,N_2534,N_2194);
or U3200 (N_3200,N_2276,N_2731);
nand U3201 (N_3201,N_2835,N_2682);
nand U3202 (N_3202,N_2755,N_2426);
nand U3203 (N_3203,N_2181,N_2757);
xnor U3204 (N_3204,N_2056,N_2404);
xnor U3205 (N_3205,N_2848,N_2937);
nor U3206 (N_3206,N_2342,N_2360);
nor U3207 (N_3207,N_2427,N_2667);
nand U3208 (N_3208,N_2938,N_2589);
xnor U3209 (N_3209,N_2968,N_2005);
and U3210 (N_3210,N_2718,N_2851);
xor U3211 (N_3211,N_2434,N_2535);
or U3212 (N_3212,N_2910,N_2284);
nor U3213 (N_3213,N_2823,N_2645);
and U3214 (N_3214,N_2902,N_2743);
and U3215 (N_3215,N_2908,N_2396);
nor U3216 (N_3216,N_2569,N_2630);
or U3217 (N_3217,N_2761,N_2991);
xnor U3218 (N_3218,N_2064,N_2933);
or U3219 (N_3219,N_2950,N_2735);
or U3220 (N_3220,N_2424,N_2450);
and U3221 (N_3221,N_2112,N_2358);
and U3222 (N_3222,N_2977,N_2577);
or U3223 (N_3223,N_2501,N_2241);
or U3224 (N_3224,N_2457,N_2140);
xnor U3225 (N_3225,N_2346,N_2878);
and U3226 (N_3226,N_2329,N_2367);
or U3227 (N_3227,N_2979,N_2351);
nor U3228 (N_3228,N_2169,N_2972);
xor U3229 (N_3229,N_2435,N_2470);
nor U3230 (N_3230,N_2014,N_2074);
and U3231 (N_3231,N_2803,N_2017);
nor U3232 (N_3232,N_2603,N_2443);
nand U3233 (N_3233,N_2173,N_2096);
nand U3234 (N_3234,N_2469,N_2428);
and U3235 (N_3235,N_2230,N_2288);
or U3236 (N_3236,N_2352,N_2338);
and U3237 (N_3237,N_2963,N_2854);
or U3238 (N_3238,N_2087,N_2850);
or U3239 (N_3239,N_2065,N_2123);
nand U3240 (N_3240,N_2382,N_2749);
and U3241 (N_3241,N_2649,N_2031);
nand U3242 (N_3242,N_2802,N_2022);
nor U3243 (N_3243,N_2040,N_2100);
nor U3244 (N_3244,N_2126,N_2984);
xor U3245 (N_3245,N_2493,N_2331);
xnor U3246 (N_3246,N_2646,N_2219);
nand U3247 (N_3247,N_2895,N_2620);
nor U3248 (N_3248,N_2072,N_2951);
xnor U3249 (N_3249,N_2362,N_2484);
nand U3250 (N_3250,N_2766,N_2439);
xor U3251 (N_3251,N_2475,N_2107);
or U3252 (N_3252,N_2736,N_2760);
nand U3253 (N_3253,N_2579,N_2211);
xnor U3254 (N_3254,N_2947,N_2815);
nand U3255 (N_3255,N_2085,N_2180);
nor U3256 (N_3256,N_2234,N_2516);
or U3257 (N_3257,N_2316,N_2058);
nand U3258 (N_3258,N_2139,N_2674);
nor U3259 (N_3259,N_2118,N_2460);
nand U3260 (N_3260,N_2306,N_2498);
nor U3261 (N_3261,N_2932,N_2573);
nor U3262 (N_3262,N_2373,N_2375);
or U3263 (N_3263,N_2099,N_2978);
or U3264 (N_3264,N_2273,N_2078);
and U3265 (N_3265,N_2595,N_2425);
nor U3266 (N_3266,N_2831,N_2956);
nand U3267 (N_3267,N_2191,N_2849);
and U3268 (N_3268,N_2372,N_2240);
and U3269 (N_3269,N_2132,N_2542);
and U3270 (N_3270,N_2976,N_2506);
or U3271 (N_3271,N_2795,N_2989);
or U3272 (N_3272,N_2935,N_2842);
xor U3273 (N_3273,N_2437,N_2614);
nor U3274 (N_3274,N_2167,N_2037);
and U3275 (N_3275,N_2299,N_2236);
xor U3276 (N_3276,N_2414,N_2176);
nor U3277 (N_3277,N_2146,N_2467);
or U3278 (N_3278,N_2388,N_2837);
nand U3279 (N_3279,N_2926,N_2709);
xnor U3280 (N_3280,N_2638,N_2402);
and U3281 (N_3281,N_2934,N_2746);
or U3282 (N_3282,N_2481,N_2043);
nand U3283 (N_3283,N_2305,N_2628);
or U3284 (N_3284,N_2179,N_2793);
and U3285 (N_3285,N_2725,N_2999);
xnor U3286 (N_3286,N_2207,N_2925);
xor U3287 (N_3287,N_2899,N_2133);
or U3288 (N_3288,N_2203,N_2844);
and U3289 (N_3289,N_2433,N_2429);
or U3290 (N_3290,N_2286,N_2774);
nand U3291 (N_3291,N_2640,N_2615);
nor U3292 (N_3292,N_2337,N_2246);
nor U3293 (N_3293,N_2032,N_2715);
xor U3294 (N_3294,N_2994,N_2220);
nand U3295 (N_3295,N_2780,N_2876);
or U3296 (N_3296,N_2706,N_2359);
nor U3297 (N_3297,N_2929,N_2828);
or U3298 (N_3298,N_2790,N_2250);
and U3299 (N_3299,N_2196,N_2901);
or U3300 (N_3300,N_2778,N_2348);
nand U3301 (N_3301,N_2884,N_2966);
and U3302 (N_3302,N_2769,N_2684);
and U3303 (N_3303,N_2605,N_2254);
xor U3304 (N_3304,N_2624,N_2156);
nand U3305 (N_3305,N_2129,N_2199);
nand U3306 (N_3306,N_2698,N_2782);
nand U3307 (N_3307,N_2019,N_2228);
or U3308 (N_3308,N_2664,N_2530);
and U3309 (N_3309,N_2390,N_2061);
or U3310 (N_3310,N_2532,N_2819);
nor U3311 (N_3311,N_2142,N_2264);
and U3312 (N_3312,N_2237,N_2868);
nand U3313 (N_3313,N_2758,N_2002);
or U3314 (N_3314,N_2593,N_2130);
nor U3315 (N_3315,N_2655,N_2536);
xnor U3316 (N_3316,N_2648,N_2458);
nor U3317 (N_3317,N_2824,N_2185);
or U3318 (N_3318,N_2383,N_2266);
nor U3319 (N_3319,N_2496,N_2229);
nand U3320 (N_3320,N_2644,N_2290);
nor U3321 (N_3321,N_2702,N_2622);
or U3322 (N_3322,N_2539,N_2879);
xnor U3323 (N_3323,N_2524,N_2554);
nand U3324 (N_3324,N_2401,N_2259);
and U3325 (N_3325,N_2202,N_2811);
nor U3326 (N_3326,N_2724,N_2796);
and U3327 (N_3327,N_2497,N_2030);
nand U3328 (N_3328,N_2865,N_2594);
xnor U3329 (N_3329,N_2082,N_2363);
xor U3330 (N_3330,N_2328,N_2967);
and U3331 (N_3331,N_2671,N_2421);
xnor U3332 (N_3332,N_2609,N_2632);
xnor U3333 (N_3333,N_2175,N_2531);
xnor U3334 (N_3334,N_2939,N_2970);
or U3335 (N_3335,N_2320,N_2635);
nand U3336 (N_3336,N_2585,N_2764);
nor U3337 (N_3337,N_2800,N_2965);
or U3338 (N_3338,N_2607,N_2499);
xor U3339 (N_3339,N_2973,N_2007);
xor U3340 (N_3340,N_2924,N_2509);
and U3341 (N_3341,N_2894,N_2275);
nand U3342 (N_3342,N_2701,N_2380);
nand U3343 (N_3343,N_2124,N_2235);
and U3344 (N_3344,N_2336,N_2827);
or U3345 (N_3345,N_2295,N_2197);
xnor U3346 (N_3346,N_2265,N_2623);
or U3347 (N_3347,N_2060,N_2111);
or U3348 (N_3348,N_2696,N_2753);
nor U3349 (N_3349,N_2201,N_2767);
or U3350 (N_3350,N_2574,N_2451);
nand U3351 (N_3351,N_2341,N_2592);
nor U3352 (N_3352,N_2817,N_2857);
xor U3353 (N_3353,N_2727,N_2697);
nor U3354 (N_3354,N_2575,N_2365);
or U3355 (N_3355,N_2411,N_2343);
xor U3356 (N_3356,N_2483,N_2687);
nor U3357 (N_3357,N_2321,N_2993);
xor U3358 (N_3358,N_2812,N_2853);
and U3359 (N_3359,N_2012,N_2015);
or U3360 (N_3360,N_2322,N_2801);
or U3361 (N_3361,N_2355,N_2601);
nor U3362 (N_3362,N_2578,N_2051);
xnor U3363 (N_3363,N_2657,N_2685);
xor U3364 (N_3364,N_2461,N_2474);
and U3365 (N_3365,N_2477,N_2559);
nand U3366 (N_3366,N_2668,N_2190);
or U3367 (N_3367,N_2105,N_2625);
nor U3368 (N_3368,N_2555,N_2008);
xor U3369 (N_3369,N_2165,N_2468);
xnor U3370 (N_3370,N_2675,N_2490);
and U3371 (N_3371,N_2311,N_2374);
nand U3372 (N_3372,N_2503,N_2249);
xnor U3373 (N_3373,N_2280,N_2596);
or U3374 (N_3374,N_2423,N_2430);
and U3375 (N_3375,N_2356,N_2489);
nand U3376 (N_3376,N_2869,N_2001);
or U3377 (N_3377,N_2026,N_2091);
or U3378 (N_3378,N_2170,N_2410);
nand U3379 (N_3379,N_2686,N_2608);
or U3380 (N_3380,N_2806,N_2515);
and U3381 (N_3381,N_2903,N_2916);
nand U3382 (N_3382,N_2500,N_2517);
or U3383 (N_3383,N_2205,N_2413);
and U3384 (N_3384,N_2399,N_2985);
xnor U3385 (N_3385,N_2519,N_2552);
nor U3386 (N_3386,N_2768,N_2874);
and U3387 (N_3387,N_2777,N_2079);
and U3388 (N_3388,N_2464,N_2958);
or U3389 (N_3389,N_2543,N_2098);
nand U3390 (N_3390,N_2915,N_2442);
nor U3391 (N_3391,N_2415,N_2982);
or U3392 (N_3392,N_2420,N_2550);
nand U3393 (N_3393,N_2117,N_2377);
nand U3394 (N_3394,N_2754,N_2930);
nand U3395 (N_3395,N_2581,N_2507);
and U3396 (N_3396,N_2478,N_2226);
and U3397 (N_3397,N_2302,N_2217);
or U3398 (N_3398,N_2942,N_2334);
and U3399 (N_3399,N_2479,N_2020);
nand U3400 (N_3400,N_2113,N_2794);
nor U3401 (N_3401,N_2011,N_2042);
or U3402 (N_3402,N_2586,N_2160);
or U3403 (N_3403,N_2770,N_2897);
xnor U3404 (N_3404,N_2291,N_2400);
nand U3405 (N_3405,N_2418,N_2417);
and U3406 (N_3406,N_2883,N_2262);
and U3407 (N_3407,N_2035,N_2907);
nor U3408 (N_3408,N_2863,N_2890);
or U3409 (N_3409,N_2135,N_2588);
nand U3410 (N_3410,N_2882,N_2799);
nor U3411 (N_3411,N_2029,N_2138);
nand U3412 (N_3412,N_2255,N_2855);
or U3413 (N_3413,N_2144,N_2927);
nor U3414 (N_3414,N_2600,N_2177);
nor U3415 (N_3415,N_2300,N_2616);
and U3416 (N_3416,N_2772,N_2830);
or U3417 (N_3417,N_2504,N_2639);
or U3418 (N_3418,N_2397,N_2325);
and U3419 (N_3419,N_2347,N_2712);
or U3420 (N_3420,N_2068,N_2024);
nor U3421 (N_3421,N_2505,N_2260);
or U3422 (N_3422,N_2705,N_2330);
xnor U3423 (N_3423,N_2308,N_2153);
nand U3424 (N_3424,N_2287,N_2807);
nor U3425 (N_3425,N_2502,N_2508);
or U3426 (N_3426,N_2313,N_2021);
nor U3427 (N_3427,N_2864,N_2084);
nor U3428 (N_3428,N_2050,N_2797);
or U3429 (N_3429,N_2998,N_2986);
xnor U3430 (N_3430,N_2784,N_2127);
xor U3431 (N_3431,N_2825,N_2272);
or U3432 (N_3432,N_2670,N_2067);
or U3433 (N_3433,N_2617,N_2075);
xnor U3434 (N_3434,N_2278,N_2486);
nand U3435 (N_3435,N_2931,N_2438);
nand U3436 (N_3436,N_2376,N_2171);
nand U3437 (N_3437,N_2323,N_2466);
nand U3438 (N_3438,N_2353,N_2602);
and U3439 (N_3439,N_2665,N_2656);
and U3440 (N_3440,N_2619,N_2862);
xor U3441 (N_3441,N_2232,N_2281);
xnor U3442 (N_3442,N_2860,N_2485);
nor U3443 (N_3443,N_2716,N_2310);
nor U3444 (N_3444,N_2110,N_2741);
nand U3445 (N_3445,N_2213,N_2447);
nand U3446 (N_3446,N_2369,N_2304);
or U3447 (N_3447,N_2476,N_2839);
xor U3448 (N_3448,N_2553,N_2339);
and U3449 (N_3449,N_2886,N_2872);
xnor U3450 (N_3450,N_2556,N_2440);
xor U3451 (N_3451,N_2178,N_2431);
or U3452 (N_3452,N_2510,N_2914);
or U3453 (N_3453,N_2885,N_2251);
xor U3454 (N_3454,N_2570,N_2119);
nor U3455 (N_3455,N_2003,N_2137);
and U3456 (N_3456,N_2345,N_2513);
xor U3457 (N_3457,N_2482,N_2094);
xnor U3458 (N_3458,N_2071,N_2403);
nor U3459 (N_3459,N_2150,N_2961);
and U3460 (N_3460,N_2141,N_2610);
xor U3461 (N_3461,N_2455,N_2206);
nor U3462 (N_3462,N_2055,N_2512);
xor U3463 (N_3463,N_2371,N_2960);
or U3464 (N_3464,N_2271,N_2627);
or U3465 (N_3465,N_2566,N_2069);
xor U3466 (N_3466,N_2463,N_2771);
and U3467 (N_3467,N_2448,N_2861);
nand U3468 (N_3468,N_2888,N_2990);
or U3469 (N_3469,N_2613,N_2871);
nand U3470 (N_3470,N_2658,N_2522);
or U3471 (N_3471,N_2997,N_2256);
nand U3472 (N_3472,N_2016,N_2626);
and U3473 (N_3473,N_2122,N_2521);
and U3474 (N_3474,N_2214,N_2545);
and U3475 (N_3475,N_2747,N_2444);
nor U3476 (N_3476,N_2441,N_2859);
nor U3477 (N_3477,N_2928,N_2834);
or U3478 (N_3478,N_2893,N_2364);
nor U3479 (N_3479,N_2389,N_2870);
nand U3480 (N_3480,N_2195,N_2528);
xnor U3481 (N_3481,N_2387,N_2083);
nand U3482 (N_3482,N_2533,N_2744);
nor U3483 (N_3483,N_2314,N_2312);
xnor U3484 (N_3484,N_2036,N_2558);
or U3485 (N_3485,N_2683,N_2274);
nand U3486 (N_3486,N_2253,N_2567);
nand U3487 (N_3487,N_2523,N_2386);
nor U3488 (N_3488,N_2407,N_2564);
nand U3489 (N_3489,N_2333,N_2905);
nand U3490 (N_3490,N_2730,N_2340);
xor U3491 (N_3491,N_2164,N_2454);
xor U3492 (N_3492,N_2732,N_2406);
nand U3493 (N_3493,N_2669,N_2267);
or U3494 (N_3494,N_2713,N_2660);
nand U3495 (N_3495,N_2361,N_2714);
nand U3496 (N_3496,N_2728,N_2662);
xnor U3497 (N_3497,N_2944,N_2561);
or U3498 (N_3498,N_2739,N_2911);
or U3499 (N_3499,N_2843,N_2919);
nor U3500 (N_3500,N_2789,N_2870);
or U3501 (N_3501,N_2681,N_2947);
nand U3502 (N_3502,N_2630,N_2395);
or U3503 (N_3503,N_2087,N_2369);
nand U3504 (N_3504,N_2594,N_2125);
or U3505 (N_3505,N_2418,N_2138);
or U3506 (N_3506,N_2873,N_2274);
nand U3507 (N_3507,N_2128,N_2310);
nor U3508 (N_3508,N_2406,N_2400);
or U3509 (N_3509,N_2455,N_2805);
xor U3510 (N_3510,N_2082,N_2490);
nor U3511 (N_3511,N_2767,N_2558);
and U3512 (N_3512,N_2794,N_2848);
nand U3513 (N_3513,N_2147,N_2767);
xor U3514 (N_3514,N_2534,N_2577);
or U3515 (N_3515,N_2352,N_2952);
nand U3516 (N_3516,N_2081,N_2915);
nor U3517 (N_3517,N_2853,N_2053);
nand U3518 (N_3518,N_2410,N_2962);
xnor U3519 (N_3519,N_2341,N_2669);
nand U3520 (N_3520,N_2692,N_2992);
nor U3521 (N_3521,N_2938,N_2019);
xor U3522 (N_3522,N_2243,N_2741);
nand U3523 (N_3523,N_2877,N_2896);
or U3524 (N_3524,N_2397,N_2827);
xor U3525 (N_3525,N_2267,N_2780);
or U3526 (N_3526,N_2114,N_2163);
xnor U3527 (N_3527,N_2263,N_2248);
nand U3528 (N_3528,N_2995,N_2652);
nand U3529 (N_3529,N_2618,N_2098);
xor U3530 (N_3530,N_2407,N_2341);
xnor U3531 (N_3531,N_2394,N_2770);
nor U3532 (N_3532,N_2260,N_2144);
nand U3533 (N_3533,N_2057,N_2389);
nor U3534 (N_3534,N_2325,N_2107);
nor U3535 (N_3535,N_2045,N_2791);
nor U3536 (N_3536,N_2032,N_2026);
or U3537 (N_3537,N_2667,N_2470);
nand U3538 (N_3538,N_2968,N_2424);
and U3539 (N_3539,N_2135,N_2774);
nand U3540 (N_3540,N_2402,N_2202);
xor U3541 (N_3541,N_2692,N_2237);
xor U3542 (N_3542,N_2926,N_2375);
nand U3543 (N_3543,N_2772,N_2662);
nor U3544 (N_3544,N_2886,N_2005);
or U3545 (N_3545,N_2668,N_2043);
xnor U3546 (N_3546,N_2375,N_2783);
or U3547 (N_3547,N_2142,N_2199);
nand U3548 (N_3548,N_2009,N_2121);
nand U3549 (N_3549,N_2626,N_2787);
nand U3550 (N_3550,N_2520,N_2085);
or U3551 (N_3551,N_2917,N_2415);
nand U3552 (N_3552,N_2470,N_2910);
xor U3553 (N_3553,N_2727,N_2823);
or U3554 (N_3554,N_2124,N_2905);
or U3555 (N_3555,N_2641,N_2733);
xor U3556 (N_3556,N_2440,N_2103);
or U3557 (N_3557,N_2116,N_2080);
nor U3558 (N_3558,N_2259,N_2937);
and U3559 (N_3559,N_2165,N_2306);
or U3560 (N_3560,N_2968,N_2946);
nor U3561 (N_3561,N_2432,N_2580);
nor U3562 (N_3562,N_2216,N_2812);
nand U3563 (N_3563,N_2776,N_2306);
nand U3564 (N_3564,N_2282,N_2417);
nand U3565 (N_3565,N_2516,N_2245);
nand U3566 (N_3566,N_2840,N_2102);
nor U3567 (N_3567,N_2066,N_2168);
xor U3568 (N_3568,N_2472,N_2011);
and U3569 (N_3569,N_2029,N_2054);
nor U3570 (N_3570,N_2926,N_2975);
xnor U3571 (N_3571,N_2596,N_2496);
nand U3572 (N_3572,N_2282,N_2992);
nand U3573 (N_3573,N_2106,N_2354);
xnor U3574 (N_3574,N_2356,N_2959);
or U3575 (N_3575,N_2361,N_2493);
and U3576 (N_3576,N_2210,N_2976);
nor U3577 (N_3577,N_2325,N_2052);
nor U3578 (N_3578,N_2584,N_2137);
or U3579 (N_3579,N_2076,N_2171);
and U3580 (N_3580,N_2955,N_2584);
nand U3581 (N_3581,N_2859,N_2083);
nor U3582 (N_3582,N_2798,N_2787);
nand U3583 (N_3583,N_2431,N_2874);
or U3584 (N_3584,N_2344,N_2226);
nand U3585 (N_3585,N_2985,N_2902);
nand U3586 (N_3586,N_2913,N_2264);
nand U3587 (N_3587,N_2267,N_2894);
xor U3588 (N_3588,N_2044,N_2910);
nand U3589 (N_3589,N_2469,N_2381);
nand U3590 (N_3590,N_2423,N_2138);
nor U3591 (N_3591,N_2583,N_2213);
xor U3592 (N_3592,N_2929,N_2832);
xor U3593 (N_3593,N_2897,N_2996);
nand U3594 (N_3594,N_2762,N_2277);
and U3595 (N_3595,N_2164,N_2942);
or U3596 (N_3596,N_2023,N_2098);
and U3597 (N_3597,N_2013,N_2994);
or U3598 (N_3598,N_2386,N_2487);
or U3599 (N_3599,N_2251,N_2834);
xnor U3600 (N_3600,N_2725,N_2897);
nand U3601 (N_3601,N_2205,N_2015);
and U3602 (N_3602,N_2350,N_2121);
nand U3603 (N_3603,N_2614,N_2509);
and U3604 (N_3604,N_2622,N_2735);
nor U3605 (N_3605,N_2554,N_2750);
xor U3606 (N_3606,N_2720,N_2517);
nor U3607 (N_3607,N_2415,N_2228);
nand U3608 (N_3608,N_2663,N_2768);
xor U3609 (N_3609,N_2078,N_2937);
or U3610 (N_3610,N_2986,N_2298);
or U3611 (N_3611,N_2180,N_2218);
and U3612 (N_3612,N_2858,N_2565);
and U3613 (N_3613,N_2905,N_2798);
nor U3614 (N_3614,N_2941,N_2130);
xnor U3615 (N_3615,N_2769,N_2928);
xnor U3616 (N_3616,N_2256,N_2436);
or U3617 (N_3617,N_2763,N_2093);
nor U3618 (N_3618,N_2098,N_2606);
and U3619 (N_3619,N_2743,N_2176);
xnor U3620 (N_3620,N_2584,N_2731);
nand U3621 (N_3621,N_2960,N_2959);
nor U3622 (N_3622,N_2032,N_2367);
or U3623 (N_3623,N_2230,N_2608);
nor U3624 (N_3624,N_2623,N_2716);
xnor U3625 (N_3625,N_2684,N_2878);
nand U3626 (N_3626,N_2084,N_2619);
and U3627 (N_3627,N_2031,N_2185);
xnor U3628 (N_3628,N_2023,N_2057);
nor U3629 (N_3629,N_2255,N_2704);
nor U3630 (N_3630,N_2859,N_2766);
xor U3631 (N_3631,N_2267,N_2103);
and U3632 (N_3632,N_2120,N_2629);
and U3633 (N_3633,N_2362,N_2140);
or U3634 (N_3634,N_2165,N_2554);
or U3635 (N_3635,N_2710,N_2991);
nor U3636 (N_3636,N_2877,N_2571);
xor U3637 (N_3637,N_2448,N_2401);
or U3638 (N_3638,N_2717,N_2674);
nor U3639 (N_3639,N_2700,N_2818);
nor U3640 (N_3640,N_2881,N_2833);
nand U3641 (N_3641,N_2800,N_2028);
nor U3642 (N_3642,N_2667,N_2924);
or U3643 (N_3643,N_2992,N_2379);
and U3644 (N_3644,N_2649,N_2625);
xor U3645 (N_3645,N_2466,N_2829);
nor U3646 (N_3646,N_2562,N_2650);
and U3647 (N_3647,N_2470,N_2359);
nor U3648 (N_3648,N_2904,N_2212);
nand U3649 (N_3649,N_2618,N_2693);
nor U3650 (N_3650,N_2417,N_2699);
xnor U3651 (N_3651,N_2138,N_2674);
nor U3652 (N_3652,N_2559,N_2773);
or U3653 (N_3653,N_2060,N_2103);
xnor U3654 (N_3654,N_2732,N_2577);
xor U3655 (N_3655,N_2937,N_2772);
nand U3656 (N_3656,N_2351,N_2654);
nand U3657 (N_3657,N_2136,N_2532);
nor U3658 (N_3658,N_2626,N_2445);
nand U3659 (N_3659,N_2788,N_2040);
and U3660 (N_3660,N_2306,N_2157);
xor U3661 (N_3661,N_2321,N_2354);
nor U3662 (N_3662,N_2500,N_2543);
nand U3663 (N_3663,N_2292,N_2792);
or U3664 (N_3664,N_2794,N_2808);
nor U3665 (N_3665,N_2891,N_2361);
and U3666 (N_3666,N_2989,N_2184);
nand U3667 (N_3667,N_2471,N_2991);
nor U3668 (N_3668,N_2702,N_2015);
nor U3669 (N_3669,N_2198,N_2462);
nor U3670 (N_3670,N_2615,N_2274);
xnor U3671 (N_3671,N_2507,N_2537);
nor U3672 (N_3672,N_2823,N_2234);
and U3673 (N_3673,N_2676,N_2096);
nand U3674 (N_3674,N_2784,N_2782);
and U3675 (N_3675,N_2159,N_2928);
or U3676 (N_3676,N_2049,N_2715);
nand U3677 (N_3677,N_2309,N_2598);
and U3678 (N_3678,N_2130,N_2666);
nor U3679 (N_3679,N_2492,N_2989);
xnor U3680 (N_3680,N_2779,N_2003);
nand U3681 (N_3681,N_2327,N_2104);
or U3682 (N_3682,N_2554,N_2360);
and U3683 (N_3683,N_2538,N_2567);
or U3684 (N_3684,N_2549,N_2538);
and U3685 (N_3685,N_2804,N_2167);
and U3686 (N_3686,N_2240,N_2458);
or U3687 (N_3687,N_2617,N_2133);
xnor U3688 (N_3688,N_2184,N_2172);
nor U3689 (N_3689,N_2521,N_2818);
and U3690 (N_3690,N_2881,N_2172);
xnor U3691 (N_3691,N_2080,N_2339);
and U3692 (N_3692,N_2697,N_2099);
or U3693 (N_3693,N_2296,N_2999);
or U3694 (N_3694,N_2970,N_2937);
and U3695 (N_3695,N_2152,N_2884);
xnor U3696 (N_3696,N_2056,N_2795);
nand U3697 (N_3697,N_2045,N_2983);
and U3698 (N_3698,N_2553,N_2376);
and U3699 (N_3699,N_2993,N_2171);
xor U3700 (N_3700,N_2805,N_2334);
and U3701 (N_3701,N_2519,N_2017);
nand U3702 (N_3702,N_2078,N_2806);
or U3703 (N_3703,N_2785,N_2337);
or U3704 (N_3704,N_2937,N_2765);
nand U3705 (N_3705,N_2677,N_2292);
or U3706 (N_3706,N_2947,N_2732);
and U3707 (N_3707,N_2992,N_2521);
nor U3708 (N_3708,N_2707,N_2474);
nor U3709 (N_3709,N_2218,N_2159);
or U3710 (N_3710,N_2113,N_2011);
nor U3711 (N_3711,N_2030,N_2953);
and U3712 (N_3712,N_2827,N_2848);
or U3713 (N_3713,N_2132,N_2511);
and U3714 (N_3714,N_2591,N_2318);
nor U3715 (N_3715,N_2409,N_2136);
xor U3716 (N_3716,N_2966,N_2065);
nor U3717 (N_3717,N_2775,N_2749);
and U3718 (N_3718,N_2401,N_2290);
or U3719 (N_3719,N_2620,N_2388);
nand U3720 (N_3720,N_2681,N_2726);
or U3721 (N_3721,N_2385,N_2279);
nand U3722 (N_3722,N_2779,N_2863);
nand U3723 (N_3723,N_2438,N_2159);
xor U3724 (N_3724,N_2479,N_2548);
or U3725 (N_3725,N_2875,N_2277);
nor U3726 (N_3726,N_2585,N_2681);
and U3727 (N_3727,N_2752,N_2563);
and U3728 (N_3728,N_2028,N_2545);
nor U3729 (N_3729,N_2624,N_2424);
nor U3730 (N_3730,N_2960,N_2106);
nand U3731 (N_3731,N_2911,N_2146);
or U3732 (N_3732,N_2161,N_2749);
nand U3733 (N_3733,N_2531,N_2198);
or U3734 (N_3734,N_2408,N_2818);
xor U3735 (N_3735,N_2852,N_2259);
xnor U3736 (N_3736,N_2098,N_2564);
nand U3737 (N_3737,N_2469,N_2824);
and U3738 (N_3738,N_2884,N_2233);
or U3739 (N_3739,N_2332,N_2324);
nand U3740 (N_3740,N_2469,N_2709);
nor U3741 (N_3741,N_2606,N_2476);
or U3742 (N_3742,N_2710,N_2972);
nand U3743 (N_3743,N_2100,N_2354);
xor U3744 (N_3744,N_2785,N_2211);
or U3745 (N_3745,N_2476,N_2083);
nand U3746 (N_3746,N_2323,N_2880);
or U3747 (N_3747,N_2751,N_2437);
and U3748 (N_3748,N_2401,N_2343);
or U3749 (N_3749,N_2379,N_2722);
and U3750 (N_3750,N_2378,N_2777);
and U3751 (N_3751,N_2086,N_2173);
and U3752 (N_3752,N_2191,N_2293);
and U3753 (N_3753,N_2295,N_2980);
or U3754 (N_3754,N_2994,N_2586);
nand U3755 (N_3755,N_2367,N_2336);
xnor U3756 (N_3756,N_2300,N_2051);
nand U3757 (N_3757,N_2306,N_2361);
nor U3758 (N_3758,N_2774,N_2031);
and U3759 (N_3759,N_2524,N_2150);
nand U3760 (N_3760,N_2424,N_2169);
nand U3761 (N_3761,N_2344,N_2790);
nor U3762 (N_3762,N_2663,N_2181);
and U3763 (N_3763,N_2923,N_2796);
xor U3764 (N_3764,N_2798,N_2978);
nand U3765 (N_3765,N_2429,N_2736);
and U3766 (N_3766,N_2204,N_2817);
and U3767 (N_3767,N_2410,N_2503);
xor U3768 (N_3768,N_2740,N_2143);
and U3769 (N_3769,N_2096,N_2901);
nor U3770 (N_3770,N_2381,N_2390);
xor U3771 (N_3771,N_2567,N_2118);
or U3772 (N_3772,N_2498,N_2883);
xnor U3773 (N_3773,N_2749,N_2822);
nor U3774 (N_3774,N_2015,N_2896);
or U3775 (N_3775,N_2971,N_2226);
or U3776 (N_3776,N_2563,N_2333);
xor U3777 (N_3777,N_2817,N_2985);
or U3778 (N_3778,N_2101,N_2471);
nand U3779 (N_3779,N_2152,N_2668);
nand U3780 (N_3780,N_2119,N_2445);
xnor U3781 (N_3781,N_2397,N_2932);
nand U3782 (N_3782,N_2449,N_2862);
xor U3783 (N_3783,N_2977,N_2873);
or U3784 (N_3784,N_2481,N_2894);
xnor U3785 (N_3785,N_2771,N_2941);
nand U3786 (N_3786,N_2075,N_2175);
nor U3787 (N_3787,N_2267,N_2170);
or U3788 (N_3788,N_2731,N_2708);
xor U3789 (N_3789,N_2106,N_2485);
and U3790 (N_3790,N_2882,N_2642);
xor U3791 (N_3791,N_2834,N_2825);
or U3792 (N_3792,N_2651,N_2677);
and U3793 (N_3793,N_2424,N_2308);
and U3794 (N_3794,N_2605,N_2785);
nor U3795 (N_3795,N_2980,N_2375);
or U3796 (N_3796,N_2340,N_2982);
xnor U3797 (N_3797,N_2270,N_2720);
and U3798 (N_3798,N_2655,N_2685);
and U3799 (N_3799,N_2356,N_2345);
xor U3800 (N_3800,N_2331,N_2765);
or U3801 (N_3801,N_2458,N_2366);
and U3802 (N_3802,N_2601,N_2112);
nor U3803 (N_3803,N_2640,N_2230);
nor U3804 (N_3804,N_2093,N_2972);
or U3805 (N_3805,N_2672,N_2813);
and U3806 (N_3806,N_2945,N_2949);
and U3807 (N_3807,N_2366,N_2652);
and U3808 (N_3808,N_2730,N_2957);
and U3809 (N_3809,N_2254,N_2684);
nor U3810 (N_3810,N_2453,N_2649);
and U3811 (N_3811,N_2439,N_2415);
xnor U3812 (N_3812,N_2460,N_2736);
xor U3813 (N_3813,N_2976,N_2987);
xor U3814 (N_3814,N_2268,N_2339);
or U3815 (N_3815,N_2969,N_2566);
nor U3816 (N_3816,N_2635,N_2864);
and U3817 (N_3817,N_2332,N_2398);
nor U3818 (N_3818,N_2918,N_2712);
nand U3819 (N_3819,N_2418,N_2772);
nand U3820 (N_3820,N_2229,N_2058);
nor U3821 (N_3821,N_2246,N_2906);
nand U3822 (N_3822,N_2036,N_2930);
or U3823 (N_3823,N_2354,N_2926);
or U3824 (N_3824,N_2792,N_2223);
nand U3825 (N_3825,N_2106,N_2289);
xnor U3826 (N_3826,N_2042,N_2440);
and U3827 (N_3827,N_2771,N_2260);
and U3828 (N_3828,N_2157,N_2534);
or U3829 (N_3829,N_2390,N_2602);
xnor U3830 (N_3830,N_2736,N_2945);
nand U3831 (N_3831,N_2147,N_2560);
or U3832 (N_3832,N_2264,N_2896);
and U3833 (N_3833,N_2923,N_2879);
and U3834 (N_3834,N_2657,N_2392);
or U3835 (N_3835,N_2749,N_2279);
nor U3836 (N_3836,N_2398,N_2262);
or U3837 (N_3837,N_2318,N_2753);
xnor U3838 (N_3838,N_2585,N_2205);
nor U3839 (N_3839,N_2925,N_2325);
xnor U3840 (N_3840,N_2441,N_2390);
or U3841 (N_3841,N_2817,N_2290);
and U3842 (N_3842,N_2635,N_2963);
xor U3843 (N_3843,N_2987,N_2647);
nand U3844 (N_3844,N_2415,N_2918);
and U3845 (N_3845,N_2859,N_2525);
nor U3846 (N_3846,N_2603,N_2890);
xor U3847 (N_3847,N_2857,N_2924);
nand U3848 (N_3848,N_2978,N_2510);
nand U3849 (N_3849,N_2247,N_2297);
nor U3850 (N_3850,N_2105,N_2662);
nor U3851 (N_3851,N_2408,N_2555);
or U3852 (N_3852,N_2112,N_2476);
nand U3853 (N_3853,N_2965,N_2589);
xnor U3854 (N_3854,N_2398,N_2020);
nor U3855 (N_3855,N_2005,N_2504);
xor U3856 (N_3856,N_2080,N_2284);
nor U3857 (N_3857,N_2858,N_2612);
nand U3858 (N_3858,N_2065,N_2101);
and U3859 (N_3859,N_2167,N_2313);
xnor U3860 (N_3860,N_2392,N_2779);
or U3861 (N_3861,N_2464,N_2861);
or U3862 (N_3862,N_2763,N_2895);
xor U3863 (N_3863,N_2640,N_2227);
and U3864 (N_3864,N_2656,N_2590);
nand U3865 (N_3865,N_2663,N_2391);
nand U3866 (N_3866,N_2956,N_2039);
nand U3867 (N_3867,N_2820,N_2561);
nor U3868 (N_3868,N_2722,N_2633);
or U3869 (N_3869,N_2122,N_2987);
or U3870 (N_3870,N_2399,N_2200);
or U3871 (N_3871,N_2558,N_2934);
nor U3872 (N_3872,N_2078,N_2503);
and U3873 (N_3873,N_2300,N_2042);
nor U3874 (N_3874,N_2731,N_2768);
nand U3875 (N_3875,N_2096,N_2067);
nor U3876 (N_3876,N_2222,N_2616);
xnor U3877 (N_3877,N_2053,N_2260);
xor U3878 (N_3878,N_2517,N_2058);
and U3879 (N_3879,N_2876,N_2434);
xor U3880 (N_3880,N_2216,N_2068);
xor U3881 (N_3881,N_2533,N_2118);
nand U3882 (N_3882,N_2443,N_2643);
or U3883 (N_3883,N_2496,N_2751);
nand U3884 (N_3884,N_2879,N_2620);
or U3885 (N_3885,N_2133,N_2480);
xor U3886 (N_3886,N_2698,N_2783);
or U3887 (N_3887,N_2187,N_2203);
xnor U3888 (N_3888,N_2992,N_2959);
or U3889 (N_3889,N_2676,N_2475);
nand U3890 (N_3890,N_2044,N_2818);
or U3891 (N_3891,N_2393,N_2829);
nand U3892 (N_3892,N_2311,N_2185);
or U3893 (N_3893,N_2441,N_2557);
and U3894 (N_3894,N_2144,N_2843);
xnor U3895 (N_3895,N_2651,N_2082);
and U3896 (N_3896,N_2368,N_2937);
xor U3897 (N_3897,N_2393,N_2634);
xor U3898 (N_3898,N_2370,N_2081);
or U3899 (N_3899,N_2031,N_2059);
or U3900 (N_3900,N_2159,N_2008);
xor U3901 (N_3901,N_2568,N_2598);
nand U3902 (N_3902,N_2612,N_2805);
or U3903 (N_3903,N_2752,N_2569);
or U3904 (N_3904,N_2965,N_2349);
nand U3905 (N_3905,N_2575,N_2217);
or U3906 (N_3906,N_2839,N_2575);
xor U3907 (N_3907,N_2986,N_2674);
and U3908 (N_3908,N_2486,N_2043);
nor U3909 (N_3909,N_2584,N_2620);
nor U3910 (N_3910,N_2261,N_2852);
xor U3911 (N_3911,N_2516,N_2786);
xor U3912 (N_3912,N_2087,N_2164);
or U3913 (N_3913,N_2285,N_2881);
nor U3914 (N_3914,N_2817,N_2677);
nand U3915 (N_3915,N_2117,N_2019);
nor U3916 (N_3916,N_2272,N_2616);
and U3917 (N_3917,N_2829,N_2161);
nand U3918 (N_3918,N_2488,N_2942);
nand U3919 (N_3919,N_2749,N_2104);
nor U3920 (N_3920,N_2906,N_2504);
nand U3921 (N_3921,N_2136,N_2059);
or U3922 (N_3922,N_2251,N_2799);
or U3923 (N_3923,N_2908,N_2768);
nand U3924 (N_3924,N_2927,N_2166);
and U3925 (N_3925,N_2415,N_2696);
xor U3926 (N_3926,N_2744,N_2646);
nand U3927 (N_3927,N_2332,N_2090);
xnor U3928 (N_3928,N_2627,N_2319);
nor U3929 (N_3929,N_2967,N_2609);
nand U3930 (N_3930,N_2217,N_2885);
or U3931 (N_3931,N_2738,N_2133);
nor U3932 (N_3932,N_2587,N_2109);
nand U3933 (N_3933,N_2733,N_2224);
nor U3934 (N_3934,N_2716,N_2610);
xnor U3935 (N_3935,N_2378,N_2416);
xor U3936 (N_3936,N_2389,N_2884);
nand U3937 (N_3937,N_2200,N_2131);
nor U3938 (N_3938,N_2917,N_2430);
xnor U3939 (N_3939,N_2997,N_2168);
nand U3940 (N_3940,N_2110,N_2609);
nand U3941 (N_3941,N_2826,N_2686);
nand U3942 (N_3942,N_2520,N_2412);
xor U3943 (N_3943,N_2364,N_2879);
and U3944 (N_3944,N_2292,N_2572);
xnor U3945 (N_3945,N_2556,N_2564);
and U3946 (N_3946,N_2498,N_2794);
or U3947 (N_3947,N_2955,N_2767);
xor U3948 (N_3948,N_2081,N_2806);
xor U3949 (N_3949,N_2632,N_2658);
nand U3950 (N_3950,N_2148,N_2478);
nor U3951 (N_3951,N_2316,N_2407);
or U3952 (N_3952,N_2308,N_2084);
and U3953 (N_3953,N_2631,N_2171);
or U3954 (N_3954,N_2774,N_2317);
nand U3955 (N_3955,N_2326,N_2224);
or U3956 (N_3956,N_2574,N_2279);
nor U3957 (N_3957,N_2171,N_2700);
xor U3958 (N_3958,N_2564,N_2428);
nand U3959 (N_3959,N_2677,N_2746);
or U3960 (N_3960,N_2033,N_2725);
nand U3961 (N_3961,N_2063,N_2586);
and U3962 (N_3962,N_2163,N_2643);
nand U3963 (N_3963,N_2379,N_2662);
or U3964 (N_3964,N_2752,N_2400);
or U3965 (N_3965,N_2895,N_2445);
or U3966 (N_3966,N_2042,N_2200);
xnor U3967 (N_3967,N_2792,N_2815);
or U3968 (N_3968,N_2101,N_2295);
xor U3969 (N_3969,N_2917,N_2488);
nor U3970 (N_3970,N_2424,N_2841);
nand U3971 (N_3971,N_2366,N_2906);
and U3972 (N_3972,N_2938,N_2515);
or U3973 (N_3973,N_2101,N_2797);
or U3974 (N_3974,N_2430,N_2727);
and U3975 (N_3975,N_2270,N_2338);
xor U3976 (N_3976,N_2317,N_2721);
xnor U3977 (N_3977,N_2953,N_2341);
or U3978 (N_3978,N_2657,N_2540);
nor U3979 (N_3979,N_2685,N_2410);
xor U3980 (N_3980,N_2485,N_2486);
xor U3981 (N_3981,N_2721,N_2257);
nor U3982 (N_3982,N_2979,N_2930);
and U3983 (N_3983,N_2333,N_2773);
nand U3984 (N_3984,N_2009,N_2122);
nor U3985 (N_3985,N_2134,N_2534);
nand U3986 (N_3986,N_2599,N_2245);
nand U3987 (N_3987,N_2981,N_2175);
nand U3988 (N_3988,N_2904,N_2382);
nand U3989 (N_3989,N_2890,N_2304);
nand U3990 (N_3990,N_2693,N_2134);
xnor U3991 (N_3991,N_2080,N_2007);
and U3992 (N_3992,N_2849,N_2256);
nor U3993 (N_3993,N_2836,N_2046);
nor U3994 (N_3994,N_2476,N_2925);
and U3995 (N_3995,N_2116,N_2657);
xor U3996 (N_3996,N_2746,N_2218);
or U3997 (N_3997,N_2238,N_2522);
nor U3998 (N_3998,N_2396,N_2196);
nand U3999 (N_3999,N_2799,N_2301);
nand U4000 (N_4000,N_3401,N_3454);
nand U4001 (N_4001,N_3906,N_3241);
and U4002 (N_4002,N_3639,N_3201);
or U4003 (N_4003,N_3936,N_3658);
or U4004 (N_4004,N_3573,N_3869);
nand U4005 (N_4005,N_3072,N_3235);
and U4006 (N_4006,N_3593,N_3126);
or U4007 (N_4007,N_3846,N_3723);
and U4008 (N_4008,N_3160,N_3689);
xor U4009 (N_4009,N_3789,N_3890);
nand U4010 (N_4010,N_3910,N_3912);
or U4011 (N_4011,N_3883,N_3775);
nand U4012 (N_4012,N_3803,N_3133);
xor U4013 (N_4013,N_3101,N_3837);
nand U4014 (N_4014,N_3418,N_3546);
nor U4015 (N_4015,N_3635,N_3876);
xnor U4016 (N_4016,N_3048,N_3149);
nor U4017 (N_4017,N_3481,N_3339);
or U4018 (N_4018,N_3698,N_3856);
xnor U4019 (N_4019,N_3419,N_3641);
and U4020 (N_4020,N_3532,N_3547);
and U4021 (N_4021,N_3987,N_3402);
or U4022 (N_4022,N_3839,N_3290);
or U4023 (N_4023,N_3104,N_3902);
nand U4024 (N_4024,N_3759,N_3263);
nand U4025 (N_4025,N_3495,N_3594);
nand U4026 (N_4026,N_3509,N_3446);
nand U4027 (N_4027,N_3304,N_3471);
xor U4028 (N_4028,N_3943,N_3417);
nor U4029 (N_4029,N_3359,N_3988);
nor U4030 (N_4030,N_3390,N_3668);
or U4031 (N_4031,N_3824,N_3199);
nor U4032 (N_4032,N_3962,N_3559);
xor U4033 (N_4033,N_3163,N_3011);
nor U4034 (N_4034,N_3268,N_3203);
and U4035 (N_4035,N_3694,N_3188);
and U4036 (N_4036,N_3574,N_3261);
or U4037 (N_4037,N_3735,N_3485);
xor U4038 (N_4038,N_3817,N_3189);
nand U4039 (N_4039,N_3732,N_3675);
or U4040 (N_4040,N_3851,N_3649);
or U4041 (N_4041,N_3137,N_3042);
or U4042 (N_4042,N_3200,N_3385);
and U4043 (N_4043,N_3174,N_3334);
or U4044 (N_4044,N_3131,N_3752);
and U4045 (N_4045,N_3568,N_3168);
or U4046 (N_4046,N_3034,N_3090);
xor U4047 (N_4047,N_3319,N_3627);
xnor U4048 (N_4048,N_3540,N_3947);
and U4049 (N_4049,N_3143,N_3515);
xnor U4050 (N_4050,N_3792,N_3826);
and U4051 (N_4051,N_3901,N_3862);
nand U4052 (N_4052,N_3640,N_3040);
nor U4053 (N_4053,N_3814,N_3457);
xor U4054 (N_4054,N_3387,N_3172);
or U4055 (N_4055,N_3380,N_3539);
xnor U4056 (N_4056,N_3569,N_3589);
or U4057 (N_4057,N_3891,N_3666);
xnor U4058 (N_4058,N_3108,N_3183);
or U4059 (N_4059,N_3486,N_3468);
xnor U4060 (N_4060,N_3655,N_3415);
or U4061 (N_4061,N_3349,N_3262);
xnor U4062 (N_4062,N_3497,N_3356);
nand U4063 (N_4063,N_3287,N_3626);
nand U4064 (N_4064,N_3941,N_3232);
xor U4065 (N_4065,N_3541,N_3393);
xnor U4066 (N_4066,N_3522,N_3360);
or U4067 (N_4067,N_3351,N_3453);
nor U4068 (N_4068,N_3379,N_3893);
or U4069 (N_4069,N_3771,N_3488);
xor U4070 (N_4070,N_3928,N_3650);
xor U4071 (N_4071,N_3324,N_3282);
nand U4072 (N_4072,N_3612,N_3214);
nor U4073 (N_4073,N_3024,N_3500);
nand U4074 (N_4074,N_3873,N_3633);
nand U4075 (N_4075,N_3676,N_3303);
or U4076 (N_4076,N_3818,N_3507);
nand U4077 (N_4077,N_3805,N_3427);
nand U4078 (N_4078,N_3078,N_3129);
nor U4079 (N_4079,N_3683,N_3397);
nand U4080 (N_4080,N_3562,N_3355);
and U4081 (N_4081,N_3502,N_3520);
or U4082 (N_4082,N_3686,N_3845);
nand U4083 (N_4083,N_3751,N_3727);
nor U4084 (N_4084,N_3472,N_3156);
nor U4085 (N_4085,N_3866,N_3463);
and U4086 (N_4086,N_3622,N_3308);
xnor U4087 (N_4087,N_3075,N_3020);
or U4088 (N_4088,N_3750,N_3055);
nor U4089 (N_4089,N_3644,N_3313);
nor U4090 (N_4090,N_3464,N_3745);
nand U4091 (N_4091,N_3631,N_3151);
nand U4092 (N_4092,N_3190,N_3984);
nor U4093 (N_4093,N_3701,N_3140);
and U4094 (N_4094,N_3504,N_3119);
and U4095 (N_4095,N_3842,N_3062);
nor U4096 (N_4096,N_3396,N_3274);
or U4097 (N_4097,N_3843,N_3492);
and U4098 (N_4098,N_3806,N_3207);
or U4099 (N_4099,N_3616,N_3691);
or U4100 (N_4100,N_3832,N_3022);
and U4101 (N_4101,N_3301,N_3211);
nand U4102 (N_4102,N_3615,N_3587);
nor U4103 (N_4103,N_3852,N_3026);
xnor U4104 (N_4104,N_3804,N_3432);
xnor U4105 (N_4105,N_3760,N_3779);
or U4106 (N_4106,N_3758,N_3498);
nor U4107 (N_4107,N_3565,N_3608);
or U4108 (N_4108,N_3272,N_3307);
nor U4109 (N_4109,N_3868,N_3536);
xor U4110 (N_4110,N_3179,N_3538);
or U4111 (N_4111,N_3619,N_3127);
or U4112 (N_4112,N_3783,N_3479);
nand U4113 (N_4113,N_3958,N_3093);
xnor U4114 (N_4114,N_3850,N_3285);
nor U4115 (N_4115,N_3099,N_3053);
or U4116 (N_4116,N_3659,N_3208);
or U4117 (N_4117,N_3983,N_3312);
or U4118 (N_4118,N_3863,N_3003);
or U4119 (N_4119,N_3624,N_3630);
or U4120 (N_4120,N_3643,N_3667);
nor U4121 (N_4121,N_3726,N_3361);
nand U4122 (N_4122,N_3122,N_3825);
nand U4123 (N_4123,N_3798,N_3348);
or U4124 (N_4124,N_3252,N_3553);
and U4125 (N_4125,N_3341,N_3144);
or U4126 (N_4126,N_3191,N_3524);
nor U4127 (N_4127,N_3311,N_3653);
nor U4128 (N_4128,N_3979,N_3797);
or U4129 (N_4129,N_3166,N_3296);
or U4130 (N_4130,N_3919,N_3749);
or U4131 (N_4131,N_3613,N_3638);
xnor U4132 (N_4132,N_3109,N_3628);
and U4133 (N_4133,N_3972,N_3795);
and U4134 (N_4134,N_3224,N_3147);
or U4135 (N_4135,N_3769,N_3657);
or U4136 (N_4136,N_3281,N_3963);
nor U4137 (N_4137,N_3768,N_3132);
or U4138 (N_4138,N_3332,N_3271);
or U4139 (N_4139,N_3297,N_3091);
and U4140 (N_4140,N_3526,N_3996);
and U4141 (N_4141,N_3169,N_3747);
nor U4142 (N_4142,N_3969,N_3932);
nor U4143 (N_4143,N_3046,N_3244);
nand U4144 (N_4144,N_3784,N_3100);
or U4145 (N_4145,N_3357,N_3823);
nand U4146 (N_4146,N_3094,N_3195);
nor U4147 (N_4147,N_3218,N_3597);
nand U4148 (N_4148,N_3054,N_3865);
nor U4149 (N_4149,N_3314,N_3607);
nor U4150 (N_4150,N_3661,N_3736);
or U4151 (N_4151,N_3455,N_3428);
nor U4152 (N_4152,N_3098,N_3516);
xnor U4153 (N_4153,N_3935,N_3248);
nor U4154 (N_4154,N_3484,N_3346);
and U4155 (N_4155,N_3372,N_3316);
xor U4156 (N_4156,N_3861,N_3813);
or U4157 (N_4157,N_3374,N_3898);
nor U4158 (N_4158,N_3704,N_3197);
nor U4159 (N_4159,N_3702,N_3968);
or U4160 (N_4160,N_3255,N_3210);
nor U4161 (N_4161,N_3302,N_3864);
or U4162 (N_4162,N_3364,N_3422);
xnor U4163 (N_4163,N_3885,N_3378);
xor U4164 (N_4164,N_3579,N_3959);
nand U4165 (N_4165,N_3949,N_3696);
xor U4166 (N_4166,N_3448,N_3796);
xnor U4167 (N_4167,N_3435,N_3693);
and U4168 (N_4168,N_3358,N_3980);
xor U4169 (N_4169,N_3021,N_3494);
or U4170 (N_4170,N_3267,N_3860);
nand U4171 (N_4171,N_3165,N_3008);
xnor U4172 (N_4172,N_3809,N_3050);
and U4173 (N_4173,N_3849,N_3766);
nor U4174 (N_4174,N_3586,N_3025);
or U4175 (N_4175,N_3542,N_3946);
or U4176 (N_4176,N_3529,N_3327);
xor U4177 (N_4177,N_3138,N_3456);
and U4178 (N_4178,N_3872,N_3656);
nor U4179 (N_4179,N_3945,N_3052);
xor U4180 (N_4180,N_3592,N_3337);
and U4181 (N_4181,N_3964,N_3180);
xor U4182 (N_4182,N_3662,N_3373);
nor U4183 (N_4183,N_3181,N_3637);
or U4184 (N_4184,N_3007,N_3317);
or U4185 (N_4185,N_3870,N_3636);
and U4186 (N_4186,N_3037,N_3306);
nand U4187 (N_4187,N_3777,N_3715);
nand U4188 (N_4188,N_3338,N_3714);
or U4189 (N_4189,N_3551,N_3087);
xnor U4190 (N_4190,N_3071,N_3776);
xnor U4191 (N_4191,N_3220,N_3103);
xnor U4192 (N_4192,N_3002,N_3073);
xor U4193 (N_4193,N_3719,N_3343);
nor U4194 (N_4194,N_3383,N_3275);
or U4195 (N_4195,N_3342,N_3107);
and U4196 (N_4196,N_3681,N_3699);
and U4197 (N_4197,N_3413,N_3600);
and U4198 (N_4198,N_3196,N_3773);
or U4199 (N_4199,N_3018,N_3135);
nand U4200 (N_4200,N_3039,N_3533);
or U4201 (N_4201,N_3460,N_3904);
or U4202 (N_4202,N_3781,N_3918);
xnor U4203 (N_4203,N_3903,N_3086);
and U4204 (N_4204,N_3960,N_3505);
and U4205 (N_4205,N_3888,N_3894);
and U4206 (N_4206,N_3116,N_3331);
nor U4207 (N_4207,N_3152,N_3556);
nor U4208 (N_4208,N_3599,N_3377);
or U4209 (N_4209,N_3300,N_3977);
and U4210 (N_4210,N_3223,N_3530);
or U4211 (N_4211,N_3449,N_3175);
xor U4212 (N_4212,N_3482,N_3443);
nor U4213 (N_4213,N_3831,N_3009);
nor U4214 (N_4214,N_3625,N_3060);
nor U4215 (N_4215,N_3618,N_3986);
nand U4216 (N_4216,N_3370,N_3892);
and U4217 (N_4217,N_3206,N_3950);
xor U4218 (N_4218,N_3462,N_3611);
xor U4219 (N_4219,N_3217,N_3077);
nor U4220 (N_4220,N_3142,N_3774);
and U4221 (N_4221,N_3821,N_3971);
nand U4222 (N_4222,N_3162,N_3442);
xnor U4223 (N_4223,N_3209,N_3305);
nand U4224 (N_4224,N_3828,N_3887);
xnor U4225 (N_4225,N_3405,N_3291);
nor U4226 (N_4226,N_3527,N_3257);
or U4227 (N_4227,N_3917,N_3788);
and U4228 (N_4228,N_3731,N_3476);
nor U4229 (N_4229,N_3033,N_3483);
and U4230 (N_4230,N_3391,N_3043);
nand U4231 (N_4231,N_3794,N_3900);
or U4232 (N_4232,N_3877,N_3231);
or U4233 (N_4233,N_3245,N_3822);
and U4234 (N_4234,N_3330,N_3944);
or U4235 (N_4235,N_3115,N_3032);
or U4236 (N_4236,N_3510,N_3858);
or U4237 (N_4237,N_3737,N_3124);
xor U4238 (N_4238,N_3915,N_3215);
xnor U4239 (N_4239,N_3716,N_3645);
xor U4240 (N_4240,N_3085,N_3001);
nor U4241 (N_4241,N_3985,N_3848);
and U4242 (N_4242,N_3519,N_3684);
xnor U4243 (N_4243,N_3561,N_3742);
nor U4244 (N_4244,N_3679,N_3459);
and U4245 (N_4245,N_3786,N_3192);
xor U4246 (N_4246,N_3652,N_3438);
or U4247 (N_4247,N_3256,N_3755);
or U4248 (N_4248,N_3922,N_3929);
or U4249 (N_4249,N_3663,N_3997);
and U4250 (N_4250,N_3924,N_3064);
nor U4251 (N_4251,N_3881,N_3709);
and U4252 (N_4252,N_3315,N_3185);
nand U4253 (N_4253,N_3154,N_3436);
or U4254 (N_4254,N_3738,N_3545);
or U4255 (N_4255,N_3976,N_3725);
xnor U4256 (N_4256,N_3682,N_3280);
xnor U4257 (N_4257,N_3690,N_3672);
or U4258 (N_4258,N_3251,N_3847);
nand U4259 (N_4259,N_3648,N_3764);
and U4260 (N_4260,N_3700,N_3563);
nor U4261 (N_4261,N_3186,N_3182);
nand U4262 (N_4262,N_3925,N_3585);
nor U4263 (N_4263,N_3363,N_3226);
and U4264 (N_4264,N_3184,N_3933);
nor U4265 (N_4265,N_3429,N_3155);
or U4266 (N_4266,N_3230,N_3916);
or U4267 (N_4267,N_3610,N_3820);
nor U4268 (N_4268,N_3952,N_3250);
or U4269 (N_4269,N_3475,N_3581);
or U4270 (N_4270,N_3204,N_3999);
nor U4271 (N_4271,N_3493,N_3733);
nand U4272 (N_4272,N_3309,N_3005);
or U4273 (N_4273,N_3408,N_3221);
and U4274 (N_4274,N_3065,N_3791);
nand U4275 (N_4275,N_3079,N_3970);
and U4276 (N_4276,N_3057,N_3035);
or U4277 (N_4277,N_3596,N_3066);
nor U4278 (N_4278,N_3376,N_3816);
xnor U4279 (N_4279,N_3367,N_3879);
nand U4280 (N_4280,N_3743,N_3673);
nand U4281 (N_4281,N_3978,N_3068);
xor U4282 (N_4282,N_3537,N_3780);
nor U4283 (N_4283,N_3564,N_3395);
or U4284 (N_4284,N_3233,N_3095);
and U4285 (N_4285,N_3006,N_3577);
nand U4286 (N_4286,N_3447,N_3198);
and U4287 (N_4287,N_3259,N_3243);
or U4288 (N_4288,N_3678,N_3354);
and U4289 (N_4289,N_3236,N_3578);
and U4290 (N_4290,N_3807,N_3669);
nand U4291 (N_4291,N_3178,N_3857);
nor U4292 (N_4292,N_3477,N_3421);
nor U4293 (N_4293,N_3310,N_3276);
xnor U4294 (N_4294,N_3121,N_3741);
and U4295 (N_4295,N_3092,N_3246);
or U4296 (N_4296,N_3258,N_3896);
xor U4297 (N_4297,N_3973,N_3609);
nand U4298 (N_4298,N_3111,N_3956);
and U4299 (N_4299,N_3834,N_3134);
nor U4300 (N_4300,N_3712,N_3389);
xnor U4301 (N_4301,N_3028,N_3489);
xnor U4302 (N_4302,N_3753,N_3576);
and U4303 (N_4303,N_3242,N_3139);
and U4304 (N_4304,N_3931,N_3605);
nor U4305 (N_4305,N_3517,N_3323);
nand U4306 (N_4306,N_3480,N_3082);
and U4307 (N_4307,N_3782,N_3404);
nor U4308 (N_4308,N_3031,N_3878);
and U4309 (N_4309,N_3926,N_3710);
and U4310 (N_4310,N_3961,N_3219);
and U4311 (N_4311,N_3023,N_3518);
and U4312 (N_4312,N_3981,N_3029);
nand U4313 (N_4313,N_3664,N_3222);
nand U4314 (N_4314,N_3437,N_3105);
nand U4315 (N_4315,N_3521,N_3874);
xor U4316 (N_4316,N_3030,N_3161);
or U4317 (N_4317,N_3335,N_3765);
and U4318 (N_4318,N_3907,N_3080);
or U4319 (N_4319,N_3705,N_3514);
or U4320 (N_4320,N_3724,N_3920);
nor U4321 (N_4321,N_3473,N_3528);
xor U4322 (N_4322,N_3170,N_3748);
and U4323 (N_4323,N_3239,N_3213);
or U4324 (N_4324,N_3508,N_3899);
nor U4325 (N_4325,N_3014,N_3552);
nand U4326 (N_4326,N_3975,N_3566);
xnor U4327 (N_4327,N_3069,N_3423);
or U4328 (N_4328,N_3583,N_3835);
nor U4329 (N_4329,N_3859,N_3347);
xor U4330 (N_4330,N_3424,N_3365);
nand U4331 (N_4331,N_3466,N_3063);
or U4332 (N_4332,N_3746,N_3772);
or U4333 (N_4333,N_3461,N_3470);
nor U4334 (N_4334,N_3544,N_3757);
or U4335 (N_4335,N_3266,N_3588);
or U4336 (N_4336,N_3793,N_3829);
and U4337 (N_4337,N_3433,N_3017);
xor U4338 (N_4338,N_3270,N_3942);
xnor U4339 (N_4339,N_3164,N_3329);
nand U4340 (N_4340,N_3811,N_3836);
and U4341 (N_4341,N_3416,N_3897);
xnor U4342 (N_4342,N_3875,N_3854);
nand U4343 (N_4343,N_3375,N_3496);
xor U4344 (N_4344,N_3886,N_3591);
and U4345 (N_4345,N_3326,N_3409);
nand U4346 (N_4346,N_3923,N_3440);
or U4347 (N_4347,N_3193,N_3590);
and U4348 (N_4348,N_3411,N_3953);
nor U4349 (N_4349,N_3088,N_3284);
xor U4350 (N_4350,N_3819,N_3934);
xnor U4351 (N_4351,N_3117,N_3734);
nor U4352 (N_4352,N_3812,N_3680);
xnor U4353 (N_4353,N_3989,N_3340);
xor U4354 (N_4354,N_3322,N_3344);
or U4355 (N_4355,N_3499,N_3762);
nor U4356 (N_4356,N_3384,N_3350);
nor U4357 (N_4357,N_3754,N_3167);
or U4358 (N_4358,N_3130,N_3249);
nor U4359 (N_4359,N_3431,N_3927);
nand U4360 (N_4360,N_3620,N_3362);
and U4361 (N_4361,N_3216,N_3808);
nand U4362 (N_4362,N_3112,N_3294);
or U4363 (N_4363,N_3790,N_3056);
xor U4364 (N_4364,N_3228,N_3567);
and U4365 (N_4365,N_3523,N_3212);
xnor U4366 (N_4366,N_3041,N_3720);
or U4367 (N_4367,N_3321,N_3787);
or U4368 (N_4368,N_3102,N_3548);
or U4369 (N_4369,N_3549,N_3279);
or U4370 (N_4370,N_3000,N_3911);
nor U4371 (N_4371,N_3474,N_3913);
and U4372 (N_4372,N_3614,N_3623);
and U4373 (N_4373,N_3067,N_3253);
nand U4374 (N_4374,N_3535,N_3371);
or U4375 (N_4375,N_3019,N_3382);
or U4376 (N_4376,N_3051,N_3265);
or U4377 (N_4377,N_3778,N_3434);
or U4378 (N_4378,N_3908,N_3756);
and U4379 (N_4379,N_3333,N_3237);
xnor U4380 (N_4380,N_3711,N_3110);
and U4381 (N_4381,N_3465,N_3685);
nand U4382 (N_4382,N_3695,N_3293);
or U4383 (N_4383,N_3603,N_3410);
nor U4384 (N_4384,N_3721,N_3491);
xnor U4385 (N_4385,N_3044,N_3706);
and U4386 (N_4386,N_3584,N_3097);
or U4387 (N_4387,N_3642,N_3718);
nor U4388 (N_4388,N_3570,N_3176);
nand U4389 (N_4389,N_3194,N_3801);
nor U4390 (N_4390,N_3286,N_3994);
and U4391 (N_4391,N_3288,N_3406);
nand U4392 (N_4392,N_3511,N_3469);
or U4393 (N_4393,N_3458,N_3036);
or U4394 (N_4394,N_3004,N_3278);
xor U4395 (N_4395,N_3295,N_3074);
xnor U4396 (N_4396,N_3407,N_3660);
nor U4397 (N_4397,N_3954,N_3840);
or U4398 (N_4398,N_3299,N_3744);
nand U4399 (N_4399,N_3697,N_3601);
xor U4400 (N_4400,N_3974,N_3940);
and U4401 (N_4401,N_3114,N_3352);
or U4402 (N_4402,N_3047,N_3081);
or U4403 (N_4403,N_3557,N_3580);
nor U4404 (N_4404,N_3490,N_3990);
or U4405 (N_4405,N_3061,N_3905);
or U4406 (N_4406,N_3830,N_3368);
xnor U4407 (N_4407,N_3070,N_3283);
xor U4408 (N_4408,N_3575,N_3240);
nor U4409 (N_4409,N_3930,N_3513);
nand U4410 (N_4410,N_3717,N_3646);
nor U4411 (N_4411,N_3430,N_3146);
xnor U4412 (N_4412,N_3531,N_3202);
or U4413 (N_4413,N_3739,N_3992);
or U4414 (N_4414,N_3617,N_3158);
nand U4415 (N_4415,N_3965,N_3381);
nor U4416 (N_4416,N_3445,N_3799);
and U4417 (N_4417,N_3414,N_3400);
and U4418 (N_4418,N_3948,N_3487);
nor U4419 (N_4419,N_3534,N_3560);
nand U4420 (N_4420,N_3128,N_3867);
and U4421 (N_4421,N_3298,N_3159);
nand U4422 (N_4422,N_3855,N_3550);
nand U4423 (N_4423,N_3555,N_3571);
nand U4424 (N_4424,N_3123,N_3654);
or U4425 (N_4425,N_3412,N_3016);
and U4426 (N_4426,N_3045,N_3708);
nor U4427 (N_4427,N_3325,N_3844);
and U4428 (N_4428,N_3884,N_3621);
nand U4429 (N_4429,N_3572,N_3722);
and U4430 (N_4430,N_3320,N_3770);
or U4431 (N_4431,N_3478,N_3153);
nand U4432 (N_4432,N_3012,N_3238);
or U4433 (N_4433,N_3394,N_3937);
xnor U4434 (N_4434,N_3802,N_3247);
and U4435 (N_4435,N_3260,N_3728);
or U4436 (N_4436,N_3059,N_3420);
and U4437 (N_4437,N_3670,N_3827);
nor U4438 (N_4438,N_3336,N_3833);
or U4439 (N_4439,N_3229,N_3939);
and U4440 (N_4440,N_3254,N_3076);
xor U4441 (N_4441,N_3089,N_3392);
or U4442 (N_4442,N_3225,N_3399);
nor U4443 (N_4443,N_3058,N_3998);
xor U4444 (N_4444,N_3441,N_3554);
xor U4445 (N_4445,N_3800,N_3558);
xnor U4446 (N_4446,N_3467,N_3853);
nor U4447 (N_4447,N_3525,N_3841);
xnor U4448 (N_4448,N_3692,N_3010);
xnor U4449 (N_4449,N_3677,N_3647);
xor U4450 (N_4450,N_3995,N_3634);
and U4451 (N_4451,N_3703,N_3602);
nor U4452 (N_4452,N_3763,N_3761);
and U4453 (N_4453,N_3740,N_3951);
or U4454 (N_4454,N_3269,N_3403);
or U4455 (N_4455,N_3957,N_3730);
xor U4456 (N_4456,N_3501,N_3688);
nand U4457 (N_4457,N_3038,N_3991);
nand U4458 (N_4458,N_3671,N_3148);
or U4459 (N_4459,N_3083,N_3543);
nor U4460 (N_4460,N_3674,N_3629);
nand U4461 (N_4461,N_3264,N_3815);
nand U4462 (N_4462,N_3729,N_3444);
or U4463 (N_4463,N_3227,N_3150);
nor U4464 (N_4464,N_3665,N_3145);
and U4465 (N_4465,N_3084,N_3120);
nor U4466 (N_4466,N_3582,N_3838);
or U4467 (N_4467,N_3015,N_3451);
and U4468 (N_4468,N_3173,N_3967);
nor U4469 (N_4469,N_3914,N_3921);
nor U4470 (N_4470,N_3966,N_3982);
or U4471 (N_4471,N_3386,N_3450);
nand U4472 (N_4472,N_3187,N_3388);
nor U4473 (N_4473,N_3707,N_3604);
nor U4474 (N_4474,N_3895,N_3328);
and U4475 (N_4475,N_3096,N_3909);
nor U4476 (N_4476,N_3289,N_3606);
and U4477 (N_4477,N_3277,N_3366);
xnor U4478 (N_4478,N_3013,N_3993);
nand U4479 (N_4479,N_3425,N_3353);
xor U4480 (N_4480,N_3439,N_3136);
or U4481 (N_4481,N_3027,N_3234);
nor U4482 (N_4482,N_3512,N_3125);
nand U4483 (N_4483,N_3785,N_3369);
and U4484 (N_4484,N_3651,N_3426);
or U4485 (N_4485,N_3118,N_3318);
nand U4486 (N_4486,N_3141,N_3113);
and U4487 (N_4487,N_3955,N_3205);
nand U4488 (N_4488,N_3595,N_3598);
nand U4489 (N_4489,N_3503,N_3506);
or U4490 (N_4490,N_3880,N_3157);
and U4491 (N_4491,N_3292,N_3345);
and U4492 (N_4492,N_3938,N_3273);
xnor U4493 (N_4493,N_3177,N_3767);
xor U4494 (N_4494,N_3713,N_3810);
and U4495 (N_4495,N_3882,N_3171);
nand U4496 (N_4496,N_3687,N_3049);
nand U4497 (N_4497,N_3106,N_3871);
and U4498 (N_4498,N_3632,N_3452);
and U4499 (N_4499,N_3398,N_3889);
nand U4500 (N_4500,N_3856,N_3068);
xor U4501 (N_4501,N_3638,N_3721);
nor U4502 (N_4502,N_3848,N_3142);
xnor U4503 (N_4503,N_3768,N_3422);
nor U4504 (N_4504,N_3149,N_3627);
and U4505 (N_4505,N_3138,N_3245);
and U4506 (N_4506,N_3817,N_3888);
xnor U4507 (N_4507,N_3450,N_3631);
or U4508 (N_4508,N_3002,N_3807);
nand U4509 (N_4509,N_3017,N_3102);
nor U4510 (N_4510,N_3240,N_3937);
xnor U4511 (N_4511,N_3931,N_3751);
nand U4512 (N_4512,N_3777,N_3412);
or U4513 (N_4513,N_3389,N_3038);
xnor U4514 (N_4514,N_3015,N_3053);
nor U4515 (N_4515,N_3093,N_3125);
xnor U4516 (N_4516,N_3625,N_3496);
or U4517 (N_4517,N_3055,N_3797);
xnor U4518 (N_4518,N_3908,N_3179);
nor U4519 (N_4519,N_3282,N_3260);
nor U4520 (N_4520,N_3492,N_3892);
nand U4521 (N_4521,N_3186,N_3841);
xor U4522 (N_4522,N_3308,N_3884);
nor U4523 (N_4523,N_3638,N_3082);
or U4524 (N_4524,N_3853,N_3427);
or U4525 (N_4525,N_3472,N_3293);
xor U4526 (N_4526,N_3649,N_3363);
or U4527 (N_4527,N_3542,N_3682);
nand U4528 (N_4528,N_3402,N_3541);
nand U4529 (N_4529,N_3770,N_3146);
nor U4530 (N_4530,N_3121,N_3598);
xnor U4531 (N_4531,N_3801,N_3319);
xnor U4532 (N_4532,N_3344,N_3861);
xor U4533 (N_4533,N_3024,N_3231);
or U4534 (N_4534,N_3473,N_3698);
xnor U4535 (N_4535,N_3607,N_3457);
nor U4536 (N_4536,N_3184,N_3934);
or U4537 (N_4537,N_3344,N_3346);
nor U4538 (N_4538,N_3927,N_3715);
and U4539 (N_4539,N_3874,N_3245);
or U4540 (N_4540,N_3310,N_3895);
nor U4541 (N_4541,N_3031,N_3870);
or U4542 (N_4542,N_3416,N_3303);
or U4543 (N_4543,N_3385,N_3186);
nand U4544 (N_4544,N_3622,N_3680);
and U4545 (N_4545,N_3456,N_3679);
and U4546 (N_4546,N_3782,N_3203);
nand U4547 (N_4547,N_3817,N_3244);
nand U4548 (N_4548,N_3638,N_3488);
or U4549 (N_4549,N_3916,N_3801);
xnor U4550 (N_4550,N_3189,N_3330);
nor U4551 (N_4551,N_3470,N_3610);
and U4552 (N_4552,N_3681,N_3688);
nor U4553 (N_4553,N_3464,N_3453);
xnor U4554 (N_4554,N_3382,N_3101);
nand U4555 (N_4555,N_3056,N_3971);
xnor U4556 (N_4556,N_3118,N_3910);
xnor U4557 (N_4557,N_3973,N_3370);
and U4558 (N_4558,N_3654,N_3033);
and U4559 (N_4559,N_3371,N_3179);
nor U4560 (N_4560,N_3980,N_3410);
and U4561 (N_4561,N_3650,N_3517);
or U4562 (N_4562,N_3476,N_3976);
or U4563 (N_4563,N_3061,N_3847);
xor U4564 (N_4564,N_3838,N_3382);
or U4565 (N_4565,N_3072,N_3794);
nor U4566 (N_4566,N_3489,N_3370);
or U4567 (N_4567,N_3933,N_3680);
and U4568 (N_4568,N_3044,N_3511);
nand U4569 (N_4569,N_3792,N_3602);
or U4570 (N_4570,N_3962,N_3383);
or U4571 (N_4571,N_3939,N_3759);
and U4572 (N_4572,N_3021,N_3525);
xor U4573 (N_4573,N_3545,N_3732);
or U4574 (N_4574,N_3091,N_3905);
or U4575 (N_4575,N_3200,N_3173);
and U4576 (N_4576,N_3898,N_3322);
nor U4577 (N_4577,N_3842,N_3912);
nand U4578 (N_4578,N_3648,N_3660);
or U4579 (N_4579,N_3619,N_3495);
xnor U4580 (N_4580,N_3819,N_3541);
nand U4581 (N_4581,N_3958,N_3343);
nor U4582 (N_4582,N_3231,N_3814);
nor U4583 (N_4583,N_3153,N_3412);
or U4584 (N_4584,N_3400,N_3455);
nor U4585 (N_4585,N_3552,N_3239);
and U4586 (N_4586,N_3895,N_3501);
xor U4587 (N_4587,N_3955,N_3470);
or U4588 (N_4588,N_3347,N_3913);
xor U4589 (N_4589,N_3722,N_3447);
xnor U4590 (N_4590,N_3990,N_3299);
and U4591 (N_4591,N_3939,N_3607);
or U4592 (N_4592,N_3299,N_3731);
or U4593 (N_4593,N_3541,N_3533);
nor U4594 (N_4594,N_3822,N_3821);
and U4595 (N_4595,N_3101,N_3867);
xnor U4596 (N_4596,N_3871,N_3371);
or U4597 (N_4597,N_3632,N_3359);
and U4598 (N_4598,N_3809,N_3558);
nor U4599 (N_4599,N_3476,N_3011);
or U4600 (N_4600,N_3537,N_3293);
nand U4601 (N_4601,N_3650,N_3076);
and U4602 (N_4602,N_3977,N_3787);
and U4603 (N_4603,N_3441,N_3610);
and U4604 (N_4604,N_3472,N_3627);
and U4605 (N_4605,N_3353,N_3031);
or U4606 (N_4606,N_3386,N_3020);
xnor U4607 (N_4607,N_3611,N_3955);
xnor U4608 (N_4608,N_3503,N_3528);
nor U4609 (N_4609,N_3467,N_3010);
xor U4610 (N_4610,N_3336,N_3112);
and U4611 (N_4611,N_3662,N_3978);
nand U4612 (N_4612,N_3460,N_3715);
nand U4613 (N_4613,N_3441,N_3808);
or U4614 (N_4614,N_3579,N_3774);
nor U4615 (N_4615,N_3515,N_3950);
xor U4616 (N_4616,N_3306,N_3206);
nor U4617 (N_4617,N_3971,N_3976);
or U4618 (N_4618,N_3640,N_3813);
nor U4619 (N_4619,N_3912,N_3726);
nand U4620 (N_4620,N_3934,N_3177);
xnor U4621 (N_4621,N_3445,N_3337);
or U4622 (N_4622,N_3129,N_3429);
xor U4623 (N_4623,N_3619,N_3330);
xnor U4624 (N_4624,N_3105,N_3477);
nor U4625 (N_4625,N_3910,N_3445);
xor U4626 (N_4626,N_3185,N_3599);
nand U4627 (N_4627,N_3339,N_3878);
and U4628 (N_4628,N_3962,N_3274);
xnor U4629 (N_4629,N_3199,N_3684);
nor U4630 (N_4630,N_3478,N_3617);
xor U4631 (N_4631,N_3135,N_3558);
nor U4632 (N_4632,N_3506,N_3340);
nand U4633 (N_4633,N_3729,N_3205);
or U4634 (N_4634,N_3360,N_3169);
and U4635 (N_4635,N_3812,N_3091);
xor U4636 (N_4636,N_3759,N_3398);
nand U4637 (N_4637,N_3910,N_3469);
nand U4638 (N_4638,N_3779,N_3383);
and U4639 (N_4639,N_3048,N_3993);
nand U4640 (N_4640,N_3625,N_3656);
and U4641 (N_4641,N_3127,N_3368);
nor U4642 (N_4642,N_3948,N_3369);
xor U4643 (N_4643,N_3255,N_3908);
nor U4644 (N_4644,N_3439,N_3388);
nand U4645 (N_4645,N_3229,N_3945);
and U4646 (N_4646,N_3334,N_3151);
xnor U4647 (N_4647,N_3817,N_3646);
xnor U4648 (N_4648,N_3552,N_3458);
and U4649 (N_4649,N_3266,N_3506);
nand U4650 (N_4650,N_3382,N_3220);
nand U4651 (N_4651,N_3485,N_3282);
xnor U4652 (N_4652,N_3767,N_3824);
nor U4653 (N_4653,N_3838,N_3970);
nor U4654 (N_4654,N_3422,N_3117);
and U4655 (N_4655,N_3152,N_3210);
nor U4656 (N_4656,N_3481,N_3611);
or U4657 (N_4657,N_3174,N_3154);
and U4658 (N_4658,N_3477,N_3020);
nand U4659 (N_4659,N_3835,N_3514);
or U4660 (N_4660,N_3359,N_3645);
or U4661 (N_4661,N_3445,N_3423);
nand U4662 (N_4662,N_3411,N_3516);
or U4663 (N_4663,N_3656,N_3585);
nor U4664 (N_4664,N_3510,N_3523);
xnor U4665 (N_4665,N_3314,N_3220);
or U4666 (N_4666,N_3060,N_3543);
or U4667 (N_4667,N_3658,N_3322);
nand U4668 (N_4668,N_3457,N_3011);
nor U4669 (N_4669,N_3797,N_3581);
and U4670 (N_4670,N_3470,N_3552);
and U4671 (N_4671,N_3438,N_3823);
and U4672 (N_4672,N_3280,N_3916);
nand U4673 (N_4673,N_3786,N_3227);
xor U4674 (N_4674,N_3200,N_3967);
and U4675 (N_4675,N_3903,N_3800);
or U4676 (N_4676,N_3411,N_3814);
xnor U4677 (N_4677,N_3246,N_3193);
or U4678 (N_4678,N_3265,N_3736);
nand U4679 (N_4679,N_3133,N_3237);
nor U4680 (N_4680,N_3345,N_3509);
xor U4681 (N_4681,N_3593,N_3167);
and U4682 (N_4682,N_3088,N_3508);
xor U4683 (N_4683,N_3706,N_3247);
nor U4684 (N_4684,N_3964,N_3650);
xor U4685 (N_4685,N_3015,N_3311);
nand U4686 (N_4686,N_3429,N_3738);
xnor U4687 (N_4687,N_3637,N_3925);
and U4688 (N_4688,N_3057,N_3518);
and U4689 (N_4689,N_3608,N_3364);
nor U4690 (N_4690,N_3850,N_3215);
or U4691 (N_4691,N_3753,N_3567);
or U4692 (N_4692,N_3185,N_3822);
xnor U4693 (N_4693,N_3288,N_3950);
or U4694 (N_4694,N_3813,N_3030);
nor U4695 (N_4695,N_3730,N_3519);
nand U4696 (N_4696,N_3727,N_3552);
nor U4697 (N_4697,N_3078,N_3473);
and U4698 (N_4698,N_3789,N_3235);
xnor U4699 (N_4699,N_3765,N_3363);
or U4700 (N_4700,N_3368,N_3666);
xor U4701 (N_4701,N_3489,N_3504);
xor U4702 (N_4702,N_3113,N_3545);
nor U4703 (N_4703,N_3317,N_3201);
nor U4704 (N_4704,N_3172,N_3148);
nand U4705 (N_4705,N_3364,N_3953);
or U4706 (N_4706,N_3736,N_3000);
nor U4707 (N_4707,N_3636,N_3929);
nand U4708 (N_4708,N_3535,N_3983);
and U4709 (N_4709,N_3028,N_3694);
nand U4710 (N_4710,N_3172,N_3567);
xor U4711 (N_4711,N_3088,N_3676);
nand U4712 (N_4712,N_3756,N_3701);
and U4713 (N_4713,N_3817,N_3234);
or U4714 (N_4714,N_3219,N_3353);
nor U4715 (N_4715,N_3677,N_3279);
nor U4716 (N_4716,N_3574,N_3902);
xnor U4717 (N_4717,N_3057,N_3960);
nor U4718 (N_4718,N_3485,N_3533);
or U4719 (N_4719,N_3257,N_3132);
or U4720 (N_4720,N_3626,N_3532);
and U4721 (N_4721,N_3197,N_3863);
nand U4722 (N_4722,N_3450,N_3517);
xor U4723 (N_4723,N_3903,N_3496);
and U4724 (N_4724,N_3968,N_3666);
xor U4725 (N_4725,N_3603,N_3039);
nand U4726 (N_4726,N_3425,N_3899);
xor U4727 (N_4727,N_3014,N_3265);
and U4728 (N_4728,N_3670,N_3322);
and U4729 (N_4729,N_3428,N_3001);
and U4730 (N_4730,N_3860,N_3719);
xor U4731 (N_4731,N_3607,N_3377);
nor U4732 (N_4732,N_3224,N_3350);
nor U4733 (N_4733,N_3413,N_3501);
or U4734 (N_4734,N_3563,N_3056);
nand U4735 (N_4735,N_3634,N_3242);
nor U4736 (N_4736,N_3804,N_3173);
or U4737 (N_4737,N_3495,N_3313);
or U4738 (N_4738,N_3291,N_3499);
nor U4739 (N_4739,N_3726,N_3808);
or U4740 (N_4740,N_3004,N_3777);
xnor U4741 (N_4741,N_3644,N_3756);
xor U4742 (N_4742,N_3071,N_3959);
nand U4743 (N_4743,N_3114,N_3569);
or U4744 (N_4744,N_3207,N_3307);
nor U4745 (N_4745,N_3711,N_3500);
nor U4746 (N_4746,N_3581,N_3665);
xnor U4747 (N_4747,N_3953,N_3323);
xnor U4748 (N_4748,N_3168,N_3808);
nand U4749 (N_4749,N_3190,N_3588);
nor U4750 (N_4750,N_3374,N_3385);
or U4751 (N_4751,N_3146,N_3563);
xnor U4752 (N_4752,N_3262,N_3730);
nor U4753 (N_4753,N_3450,N_3596);
nand U4754 (N_4754,N_3345,N_3418);
and U4755 (N_4755,N_3867,N_3322);
or U4756 (N_4756,N_3019,N_3551);
xor U4757 (N_4757,N_3491,N_3757);
nand U4758 (N_4758,N_3770,N_3394);
nor U4759 (N_4759,N_3406,N_3751);
and U4760 (N_4760,N_3690,N_3667);
nand U4761 (N_4761,N_3732,N_3235);
nand U4762 (N_4762,N_3945,N_3705);
and U4763 (N_4763,N_3534,N_3651);
or U4764 (N_4764,N_3099,N_3568);
and U4765 (N_4765,N_3244,N_3327);
or U4766 (N_4766,N_3848,N_3870);
and U4767 (N_4767,N_3769,N_3821);
and U4768 (N_4768,N_3846,N_3256);
or U4769 (N_4769,N_3698,N_3920);
nand U4770 (N_4770,N_3669,N_3413);
and U4771 (N_4771,N_3347,N_3776);
nand U4772 (N_4772,N_3067,N_3928);
and U4773 (N_4773,N_3775,N_3983);
nor U4774 (N_4774,N_3833,N_3811);
nand U4775 (N_4775,N_3725,N_3486);
and U4776 (N_4776,N_3568,N_3221);
or U4777 (N_4777,N_3348,N_3161);
or U4778 (N_4778,N_3799,N_3520);
nor U4779 (N_4779,N_3838,N_3888);
nor U4780 (N_4780,N_3219,N_3164);
and U4781 (N_4781,N_3821,N_3715);
nor U4782 (N_4782,N_3573,N_3842);
nor U4783 (N_4783,N_3816,N_3375);
or U4784 (N_4784,N_3162,N_3627);
nor U4785 (N_4785,N_3494,N_3235);
or U4786 (N_4786,N_3455,N_3523);
nor U4787 (N_4787,N_3550,N_3172);
nor U4788 (N_4788,N_3611,N_3461);
or U4789 (N_4789,N_3340,N_3384);
and U4790 (N_4790,N_3191,N_3202);
or U4791 (N_4791,N_3228,N_3290);
xor U4792 (N_4792,N_3471,N_3582);
nor U4793 (N_4793,N_3205,N_3608);
xnor U4794 (N_4794,N_3185,N_3581);
nor U4795 (N_4795,N_3609,N_3363);
or U4796 (N_4796,N_3525,N_3177);
or U4797 (N_4797,N_3577,N_3638);
nor U4798 (N_4798,N_3142,N_3391);
nand U4799 (N_4799,N_3402,N_3283);
xnor U4800 (N_4800,N_3961,N_3321);
xor U4801 (N_4801,N_3078,N_3144);
and U4802 (N_4802,N_3183,N_3315);
nor U4803 (N_4803,N_3002,N_3935);
xnor U4804 (N_4804,N_3974,N_3232);
nand U4805 (N_4805,N_3460,N_3283);
nand U4806 (N_4806,N_3953,N_3707);
or U4807 (N_4807,N_3889,N_3616);
or U4808 (N_4808,N_3742,N_3840);
or U4809 (N_4809,N_3832,N_3208);
nand U4810 (N_4810,N_3221,N_3583);
and U4811 (N_4811,N_3514,N_3465);
and U4812 (N_4812,N_3161,N_3422);
and U4813 (N_4813,N_3379,N_3643);
xnor U4814 (N_4814,N_3889,N_3564);
nor U4815 (N_4815,N_3673,N_3044);
xor U4816 (N_4816,N_3870,N_3917);
nand U4817 (N_4817,N_3638,N_3644);
or U4818 (N_4818,N_3293,N_3674);
nand U4819 (N_4819,N_3333,N_3685);
xnor U4820 (N_4820,N_3667,N_3347);
nor U4821 (N_4821,N_3829,N_3385);
and U4822 (N_4822,N_3570,N_3203);
xor U4823 (N_4823,N_3083,N_3165);
xor U4824 (N_4824,N_3392,N_3049);
xor U4825 (N_4825,N_3768,N_3737);
xnor U4826 (N_4826,N_3131,N_3393);
nand U4827 (N_4827,N_3510,N_3160);
nand U4828 (N_4828,N_3857,N_3936);
nand U4829 (N_4829,N_3858,N_3271);
or U4830 (N_4830,N_3925,N_3959);
nand U4831 (N_4831,N_3791,N_3795);
or U4832 (N_4832,N_3285,N_3839);
or U4833 (N_4833,N_3957,N_3219);
nor U4834 (N_4834,N_3639,N_3945);
or U4835 (N_4835,N_3784,N_3880);
or U4836 (N_4836,N_3108,N_3461);
nand U4837 (N_4837,N_3931,N_3477);
xor U4838 (N_4838,N_3718,N_3255);
nor U4839 (N_4839,N_3110,N_3364);
nand U4840 (N_4840,N_3411,N_3871);
and U4841 (N_4841,N_3042,N_3600);
nand U4842 (N_4842,N_3724,N_3085);
nor U4843 (N_4843,N_3732,N_3233);
and U4844 (N_4844,N_3047,N_3607);
nand U4845 (N_4845,N_3468,N_3331);
xnor U4846 (N_4846,N_3654,N_3608);
and U4847 (N_4847,N_3763,N_3928);
and U4848 (N_4848,N_3134,N_3673);
nor U4849 (N_4849,N_3266,N_3420);
nor U4850 (N_4850,N_3802,N_3848);
and U4851 (N_4851,N_3408,N_3364);
nand U4852 (N_4852,N_3763,N_3934);
nand U4853 (N_4853,N_3642,N_3999);
or U4854 (N_4854,N_3146,N_3086);
nand U4855 (N_4855,N_3245,N_3835);
nor U4856 (N_4856,N_3525,N_3110);
nor U4857 (N_4857,N_3418,N_3900);
or U4858 (N_4858,N_3660,N_3345);
xor U4859 (N_4859,N_3757,N_3609);
and U4860 (N_4860,N_3633,N_3759);
xnor U4861 (N_4861,N_3832,N_3986);
or U4862 (N_4862,N_3659,N_3660);
nor U4863 (N_4863,N_3220,N_3401);
and U4864 (N_4864,N_3310,N_3138);
xor U4865 (N_4865,N_3686,N_3883);
nand U4866 (N_4866,N_3809,N_3336);
nor U4867 (N_4867,N_3105,N_3665);
nand U4868 (N_4868,N_3168,N_3111);
nor U4869 (N_4869,N_3751,N_3510);
or U4870 (N_4870,N_3362,N_3230);
nor U4871 (N_4871,N_3246,N_3427);
nand U4872 (N_4872,N_3192,N_3334);
xnor U4873 (N_4873,N_3771,N_3312);
and U4874 (N_4874,N_3820,N_3103);
xnor U4875 (N_4875,N_3445,N_3430);
or U4876 (N_4876,N_3238,N_3999);
xor U4877 (N_4877,N_3005,N_3259);
nor U4878 (N_4878,N_3739,N_3818);
or U4879 (N_4879,N_3148,N_3141);
xor U4880 (N_4880,N_3044,N_3308);
and U4881 (N_4881,N_3486,N_3876);
xnor U4882 (N_4882,N_3829,N_3240);
xnor U4883 (N_4883,N_3488,N_3664);
nor U4884 (N_4884,N_3968,N_3983);
or U4885 (N_4885,N_3796,N_3730);
or U4886 (N_4886,N_3772,N_3280);
xor U4887 (N_4887,N_3674,N_3751);
or U4888 (N_4888,N_3969,N_3565);
and U4889 (N_4889,N_3829,N_3157);
or U4890 (N_4890,N_3087,N_3562);
nor U4891 (N_4891,N_3579,N_3234);
and U4892 (N_4892,N_3768,N_3562);
nor U4893 (N_4893,N_3339,N_3249);
or U4894 (N_4894,N_3884,N_3114);
or U4895 (N_4895,N_3841,N_3706);
nand U4896 (N_4896,N_3455,N_3420);
and U4897 (N_4897,N_3686,N_3249);
or U4898 (N_4898,N_3331,N_3512);
nand U4899 (N_4899,N_3284,N_3484);
xnor U4900 (N_4900,N_3779,N_3623);
xor U4901 (N_4901,N_3441,N_3195);
nand U4902 (N_4902,N_3803,N_3951);
xnor U4903 (N_4903,N_3707,N_3768);
and U4904 (N_4904,N_3376,N_3277);
or U4905 (N_4905,N_3813,N_3436);
nor U4906 (N_4906,N_3898,N_3448);
nor U4907 (N_4907,N_3934,N_3795);
or U4908 (N_4908,N_3157,N_3918);
nor U4909 (N_4909,N_3833,N_3518);
nand U4910 (N_4910,N_3146,N_3814);
xnor U4911 (N_4911,N_3768,N_3867);
and U4912 (N_4912,N_3624,N_3516);
nand U4913 (N_4913,N_3030,N_3223);
xnor U4914 (N_4914,N_3329,N_3640);
nand U4915 (N_4915,N_3151,N_3268);
xnor U4916 (N_4916,N_3226,N_3063);
nand U4917 (N_4917,N_3634,N_3378);
xnor U4918 (N_4918,N_3810,N_3276);
nor U4919 (N_4919,N_3357,N_3143);
xor U4920 (N_4920,N_3503,N_3765);
nand U4921 (N_4921,N_3399,N_3212);
or U4922 (N_4922,N_3825,N_3240);
and U4923 (N_4923,N_3845,N_3956);
or U4924 (N_4924,N_3124,N_3753);
or U4925 (N_4925,N_3274,N_3574);
xnor U4926 (N_4926,N_3981,N_3067);
nor U4927 (N_4927,N_3415,N_3632);
nand U4928 (N_4928,N_3467,N_3728);
and U4929 (N_4929,N_3550,N_3957);
or U4930 (N_4930,N_3084,N_3844);
and U4931 (N_4931,N_3459,N_3536);
nor U4932 (N_4932,N_3095,N_3488);
or U4933 (N_4933,N_3851,N_3762);
xor U4934 (N_4934,N_3606,N_3926);
nor U4935 (N_4935,N_3320,N_3016);
and U4936 (N_4936,N_3998,N_3315);
nor U4937 (N_4937,N_3008,N_3938);
xor U4938 (N_4938,N_3575,N_3282);
or U4939 (N_4939,N_3886,N_3197);
xor U4940 (N_4940,N_3196,N_3482);
xor U4941 (N_4941,N_3901,N_3319);
nor U4942 (N_4942,N_3916,N_3051);
xnor U4943 (N_4943,N_3543,N_3882);
or U4944 (N_4944,N_3749,N_3563);
or U4945 (N_4945,N_3617,N_3911);
xor U4946 (N_4946,N_3502,N_3433);
xnor U4947 (N_4947,N_3739,N_3686);
or U4948 (N_4948,N_3125,N_3604);
xor U4949 (N_4949,N_3306,N_3752);
or U4950 (N_4950,N_3167,N_3670);
nor U4951 (N_4951,N_3312,N_3289);
or U4952 (N_4952,N_3886,N_3387);
nand U4953 (N_4953,N_3312,N_3389);
nand U4954 (N_4954,N_3754,N_3508);
nand U4955 (N_4955,N_3387,N_3904);
and U4956 (N_4956,N_3365,N_3063);
and U4957 (N_4957,N_3744,N_3037);
nand U4958 (N_4958,N_3899,N_3494);
and U4959 (N_4959,N_3754,N_3982);
nor U4960 (N_4960,N_3259,N_3890);
nor U4961 (N_4961,N_3053,N_3709);
or U4962 (N_4962,N_3689,N_3696);
nand U4963 (N_4963,N_3586,N_3903);
or U4964 (N_4964,N_3941,N_3599);
xnor U4965 (N_4965,N_3107,N_3886);
nand U4966 (N_4966,N_3081,N_3900);
or U4967 (N_4967,N_3294,N_3626);
or U4968 (N_4968,N_3636,N_3919);
nand U4969 (N_4969,N_3393,N_3520);
xnor U4970 (N_4970,N_3387,N_3100);
nand U4971 (N_4971,N_3546,N_3721);
nand U4972 (N_4972,N_3543,N_3853);
or U4973 (N_4973,N_3154,N_3097);
xor U4974 (N_4974,N_3867,N_3470);
nor U4975 (N_4975,N_3724,N_3080);
xor U4976 (N_4976,N_3932,N_3170);
nor U4977 (N_4977,N_3890,N_3461);
nand U4978 (N_4978,N_3050,N_3543);
nor U4979 (N_4979,N_3722,N_3294);
nor U4980 (N_4980,N_3026,N_3610);
nor U4981 (N_4981,N_3465,N_3384);
nor U4982 (N_4982,N_3216,N_3996);
nor U4983 (N_4983,N_3370,N_3871);
xor U4984 (N_4984,N_3208,N_3748);
nor U4985 (N_4985,N_3512,N_3842);
nor U4986 (N_4986,N_3356,N_3149);
or U4987 (N_4987,N_3068,N_3090);
xor U4988 (N_4988,N_3270,N_3365);
and U4989 (N_4989,N_3046,N_3577);
or U4990 (N_4990,N_3153,N_3329);
or U4991 (N_4991,N_3272,N_3702);
xor U4992 (N_4992,N_3721,N_3913);
xor U4993 (N_4993,N_3096,N_3437);
nand U4994 (N_4994,N_3118,N_3087);
and U4995 (N_4995,N_3467,N_3074);
nor U4996 (N_4996,N_3012,N_3463);
nand U4997 (N_4997,N_3534,N_3909);
nand U4998 (N_4998,N_3123,N_3524);
nor U4999 (N_4999,N_3430,N_3592);
xnor U5000 (N_5000,N_4304,N_4959);
and U5001 (N_5001,N_4351,N_4328);
and U5002 (N_5002,N_4677,N_4666);
xor U5003 (N_5003,N_4430,N_4603);
nand U5004 (N_5004,N_4403,N_4752);
nand U5005 (N_5005,N_4776,N_4963);
and U5006 (N_5006,N_4179,N_4934);
xnor U5007 (N_5007,N_4923,N_4979);
nor U5008 (N_5008,N_4297,N_4514);
nand U5009 (N_5009,N_4784,N_4726);
xor U5010 (N_5010,N_4830,N_4252);
nor U5011 (N_5011,N_4819,N_4334);
and U5012 (N_5012,N_4417,N_4006);
xor U5013 (N_5013,N_4438,N_4619);
and U5014 (N_5014,N_4922,N_4574);
nand U5015 (N_5015,N_4311,N_4924);
or U5016 (N_5016,N_4333,N_4489);
nor U5017 (N_5017,N_4238,N_4994);
or U5018 (N_5018,N_4378,N_4967);
xor U5019 (N_5019,N_4173,N_4741);
and U5020 (N_5020,N_4267,N_4192);
nor U5021 (N_5021,N_4560,N_4874);
nand U5022 (N_5022,N_4169,N_4082);
and U5023 (N_5023,N_4408,N_4734);
xor U5024 (N_5024,N_4101,N_4626);
nor U5025 (N_5025,N_4010,N_4027);
and U5026 (N_5026,N_4686,N_4866);
or U5027 (N_5027,N_4893,N_4270);
nor U5028 (N_5028,N_4463,N_4385);
and U5029 (N_5029,N_4160,N_4850);
nand U5030 (N_5030,N_4847,N_4371);
nand U5031 (N_5031,N_4436,N_4092);
or U5032 (N_5032,N_4380,N_4142);
nand U5033 (N_5033,N_4155,N_4766);
or U5034 (N_5034,N_4158,N_4234);
nor U5035 (N_5035,N_4835,N_4511);
xnor U5036 (N_5036,N_4901,N_4109);
xor U5037 (N_5037,N_4769,N_4949);
xnor U5038 (N_5038,N_4896,N_4258);
or U5039 (N_5039,N_4903,N_4995);
nand U5040 (N_5040,N_4310,N_4374);
and U5041 (N_5041,N_4865,N_4115);
and U5042 (N_5042,N_4250,N_4411);
and U5043 (N_5043,N_4559,N_4014);
xor U5044 (N_5044,N_4637,N_4879);
xor U5045 (N_5045,N_4080,N_4797);
xor U5046 (N_5046,N_4883,N_4937);
nand U5047 (N_5047,N_4647,N_4163);
nor U5048 (N_5048,N_4294,N_4805);
nor U5049 (N_5049,N_4673,N_4578);
nand U5050 (N_5050,N_4800,N_4357);
or U5051 (N_5051,N_4525,N_4210);
nor U5052 (N_5052,N_4892,N_4118);
or U5053 (N_5053,N_4391,N_4499);
nor U5054 (N_5054,N_4185,N_4206);
nand U5055 (N_5055,N_4887,N_4376);
xor U5056 (N_5056,N_4093,N_4953);
or U5057 (N_5057,N_4672,N_4736);
and U5058 (N_5058,N_4616,N_4406);
nor U5059 (N_5059,N_4941,N_4057);
xor U5060 (N_5060,N_4418,N_4491);
or U5061 (N_5061,N_4951,N_4876);
nand U5062 (N_5062,N_4723,N_4465);
nand U5063 (N_5063,N_4838,N_4220);
and U5064 (N_5064,N_4164,N_4728);
nand U5065 (N_5065,N_4359,N_4003);
nand U5066 (N_5066,N_4244,N_4042);
xor U5067 (N_5067,N_4791,N_4415);
and U5068 (N_5068,N_4447,N_4288);
nor U5069 (N_5069,N_4864,N_4205);
nand U5070 (N_5070,N_4320,N_4638);
nor U5071 (N_5071,N_4226,N_4919);
or U5072 (N_5072,N_4822,N_4177);
nor U5073 (N_5073,N_4579,N_4516);
nand U5074 (N_5074,N_4702,N_4381);
xnor U5075 (N_5075,N_4253,N_4325);
or U5076 (N_5076,N_4631,N_4722);
or U5077 (N_5077,N_4368,N_4668);
or U5078 (N_5078,N_4494,N_4674);
and U5079 (N_5079,N_4824,N_4586);
and U5080 (N_5080,N_4182,N_4028);
xnor U5081 (N_5081,N_4015,N_4571);
or U5082 (N_5082,N_4171,N_4375);
and U5083 (N_5083,N_4984,N_4130);
nor U5084 (N_5084,N_4695,N_4059);
nand U5085 (N_5085,N_4562,N_4506);
nor U5086 (N_5086,N_4920,N_4921);
or U5087 (N_5087,N_4398,N_4435);
or U5088 (N_5088,N_4624,N_4426);
nand U5089 (N_5089,N_4373,N_4821);
xor U5090 (N_5090,N_4277,N_4534);
nor U5091 (N_5091,N_4051,N_4189);
nor U5092 (N_5092,N_4260,N_4476);
xor U5093 (N_5093,N_4157,N_4843);
or U5094 (N_5094,N_4416,N_4399);
xor U5095 (N_5095,N_4862,N_4460);
xor U5096 (N_5096,N_4473,N_4707);
nand U5097 (N_5097,N_4251,N_4369);
xnor U5098 (N_5098,N_4096,N_4214);
or U5099 (N_5099,N_4980,N_4219);
nor U5100 (N_5100,N_4909,N_4973);
and U5101 (N_5101,N_4259,N_4688);
nand U5102 (N_5102,N_4427,N_4105);
xor U5103 (N_5103,N_4040,N_4193);
and U5104 (N_5104,N_4857,N_4946);
xnor U5105 (N_5105,N_4732,N_4318);
nor U5106 (N_5106,N_4029,N_4282);
or U5107 (N_5107,N_4256,N_4993);
nand U5108 (N_5108,N_4429,N_4431);
nor U5109 (N_5109,N_4167,N_4954);
xnor U5110 (N_5110,N_4079,N_4299);
nand U5111 (N_5111,N_4235,N_4420);
and U5112 (N_5112,N_4492,N_4183);
nand U5113 (N_5113,N_4496,N_4224);
nand U5114 (N_5114,N_4787,N_4407);
and U5115 (N_5115,N_4337,N_4263);
nand U5116 (N_5116,N_4948,N_4513);
nand U5117 (N_5117,N_4622,N_4462);
or U5118 (N_5118,N_4454,N_4793);
nand U5119 (N_5119,N_4877,N_4912);
nand U5120 (N_5120,N_4938,N_4504);
xor U5121 (N_5121,N_4257,N_4354);
nand U5122 (N_5122,N_4120,N_4213);
and U5123 (N_5123,N_4097,N_4518);
nor U5124 (N_5124,N_4349,N_4744);
nor U5125 (N_5125,N_4087,N_4607);
nand U5126 (N_5126,N_4820,N_4795);
nand U5127 (N_5127,N_4166,N_4456);
and U5128 (N_5128,N_4414,N_4701);
nand U5129 (N_5129,N_4558,N_4470);
or U5130 (N_5130,N_4340,N_4746);
xor U5131 (N_5131,N_4653,N_4273);
xnor U5132 (N_5132,N_4348,N_4248);
xnor U5133 (N_5133,N_4881,N_4846);
or U5134 (N_5134,N_4030,N_4945);
nand U5135 (N_5135,N_4854,N_4002);
and U5136 (N_5136,N_4670,N_4550);
xor U5137 (N_5137,N_4608,N_4085);
and U5138 (N_5138,N_4988,N_4140);
and U5139 (N_5139,N_4113,N_4347);
nand U5140 (N_5140,N_4405,N_4428);
nor U5141 (N_5141,N_4636,N_4271);
and U5142 (N_5142,N_4577,N_4678);
and U5143 (N_5143,N_4060,N_4186);
xor U5144 (N_5144,N_4992,N_4245);
or U5145 (N_5145,N_4449,N_4927);
or U5146 (N_5146,N_4366,N_4190);
or U5147 (N_5147,N_4291,N_4597);
xor U5148 (N_5148,N_4441,N_4308);
nand U5149 (N_5149,N_4041,N_4543);
and U5150 (N_5150,N_4660,N_4884);
or U5151 (N_5151,N_4545,N_4024);
and U5152 (N_5152,N_4095,N_4900);
xor U5153 (N_5153,N_4471,N_4007);
nand U5154 (N_5154,N_4855,N_4239);
or U5155 (N_5155,N_4018,N_4104);
and U5156 (N_5156,N_4459,N_4032);
nor U5157 (N_5157,N_4084,N_4071);
or U5158 (N_5158,N_4397,N_4585);
nor U5159 (N_5159,N_4554,N_4898);
nand U5160 (N_5160,N_4849,N_4625);
nand U5161 (N_5161,N_4851,N_4590);
and U5162 (N_5162,N_4798,N_4102);
nor U5163 (N_5163,N_4233,N_4268);
and U5164 (N_5164,N_4243,N_4323);
nor U5165 (N_5165,N_4196,N_4069);
xor U5166 (N_5166,N_4989,N_4049);
nor U5167 (N_5167,N_4640,N_4675);
or U5168 (N_5168,N_4394,N_4602);
xnor U5169 (N_5169,N_4487,N_4526);
nor U5170 (N_5170,N_4650,N_4116);
nand U5171 (N_5171,N_4966,N_4977);
and U5172 (N_5172,N_4696,N_4996);
xor U5173 (N_5173,N_4026,N_4284);
nor U5174 (N_5174,N_4731,N_4227);
and U5175 (N_5175,N_4236,N_4469);
nor U5176 (N_5176,N_4161,N_4222);
nand U5177 (N_5177,N_4572,N_4106);
and U5178 (N_5178,N_4779,N_4794);
or U5179 (N_5179,N_4446,N_4532);
nand U5180 (N_5180,N_4745,N_4209);
nand U5181 (N_5181,N_4488,N_4434);
nand U5182 (N_5182,N_4617,N_4567);
xnor U5183 (N_5183,N_4801,N_4187);
and U5184 (N_5184,N_4448,N_4781);
or U5185 (N_5185,N_4017,N_4442);
nor U5186 (N_5186,N_4902,N_4131);
nor U5187 (N_5187,N_4241,N_4422);
nand U5188 (N_5188,N_4601,N_4455);
and U5189 (N_5189,N_4802,N_4181);
or U5190 (N_5190,N_4775,N_4022);
nand U5191 (N_5191,N_4122,N_4149);
xor U5192 (N_5192,N_4302,N_4409);
xnor U5193 (N_5193,N_4552,N_4316);
and U5194 (N_5194,N_4063,N_4721);
or U5195 (N_5195,N_4940,N_4046);
or U5196 (N_5196,N_4144,N_4742);
nor U5197 (N_5197,N_4001,N_4064);
or U5198 (N_5198,N_4971,N_4382);
or U5199 (N_5199,N_4604,N_4778);
or U5200 (N_5200,N_4642,N_4154);
nor U5201 (N_5201,N_4710,N_4869);
xnor U5202 (N_5202,N_4035,N_4012);
or U5203 (N_5203,N_4203,N_4910);
and U5204 (N_5204,N_4107,N_4443);
nand U5205 (N_5205,N_4965,N_4955);
or U5206 (N_5206,N_4648,N_4276);
xor U5207 (N_5207,N_4162,N_4305);
nor U5208 (N_5208,N_4094,N_4174);
or U5209 (N_5209,N_4180,N_4393);
nand U5210 (N_5210,N_4128,N_4699);
and U5211 (N_5211,N_4772,N_4911);
nand U5212 (N_5212,N_4815,N_4062);
and U5213 (N_5213,N_4885,N_4528);
or U5214 (N_5214,N_4451,N_4058);
xnor U5215 (N_5215,N_4468,N_4502);
xor U5216 (N_5216,N_4262,N_4594);
xor U5217 (N_5217,N_4823,N_4090);
xnor U5218 (N_5218,N_4942,N_4292);
or U5219 (N_5219,N_4352,N_4037);
nor U5220 (N_5220,N_4498,N_4467);
xor U5221 (N_5221,N_4837,N_4894);
or U5222 (N_5222,N_4649,N_4845);
and U5223 (N_5223,N_4056,N_4536);
nand U5224 (N_5224,N_4629,N_4561);
xor U5225 (N_5225,N_4384,N_4976);
xor U5226 (N_5226,N_4814,N_4540);
xnor U5227 (N_5227,N_4240,N_4939);
nand U5228 (N_5228,N_4043,N_4520);
nor U5229 (N_5229,N_4524,N_4895);
nor U5230 (N_5230,N_4266,N_4147);
and U5231 (N_5231,N_4669,N_4836);
nor U5232 (N_5232,N_4293,N_4507);
and U5233 (N_5233,N_4098,N_4868);
xnor U5234 (N_5234,N_4537,N_4175);
xnor U5235 (N_5235,N_4970,N_4691);
and U5236 (N_5236,N_4486,N_4685);
and U5237 (N_5237,N_4000,N_4272);
nor U5238 (N_5238,N_4533,N_4423);
nor U5239 (N_5239,N_4176,N_4321);
or U5240 (N_5240,N_4289,N_4480);
or U5241 (N_5241,N_4777,N_4074);
and U5242 (N_5242,N_4553,N_4453);
xor U5243 (N_5243,N_4362,N_4413);
or U5244 (N_5244,N_4360,N_4072);
nand U5245 (N_5245,N_4832,N_4875);
or U5246 (N_5246,N_4091,N_4905);
xnor U5247 (N_5247,N_4729,N_4828);
nand U5248 (N_5248,N_4529,N_4714);
and U5249 (N_5249,N_4719,N_4332);
xnor U5250 (N_5250,N_4872,N_4606);
nor U5251 (N_5251,N_4708,N_4557);
or U5252 (N_5252,N_4681,N_4103);
xnor U5253 (N_5253,N_4197,N_4969);
or U5254 (N_5254,N_4661,N_4576);
xor U5255 (N_5255,N_4662,N_4510);
nand U5256 (N_5256,N_4402,N_4111);
nor U5257 (N_5257,N_4700,N_4134);
or U5258 (N_5258,N_4760,N_4531);
or U5259 (N_5259,N_4275,N_4123);
nor U5260 (N_5260,N_4724,N_4052);
and U5261 (N_5261,N_4365,N_4718);
and U5262 (N_5262,N_4605,N_4265);
nor U5263 (N_5263,N_4750,N_4743);
nand U5264 (N_5264,N_4806,N_4129);
or U5265 (N_5265,N_4314,N_4612);
nor U5266 (N_5266,N_4589,N_4555);
nor U5267 (N_5267,N_4433,N_4034);
and U5268 (N_5268,N_4763,N_4367);
nor U5269 (N_5269,N_4915,N_4931);
and U5270 (N_5270,N_4584,N_4546);
xor U5271 (N_5271,N_4005,N_4740);
nand U5272 (N_5272,N_4983,N_4108);
nand U5273 (N_5273,N_4544,N_4852);
or U5274 (N_5274,N_4148,N_4073);
or U5275 (N_5275,N_4817,N_4986);
nor U5276 (N_5276,N_4457,N_4246);
nand U5277 (N_5277,N_4889,N_4200);
nor U5278 (N_5278,N_4410,N_4466);
xor U5279 (N_5279,N_4503,N_4009);
and U5280 (N_5280,N_4753,N_4549);
nor U5281 (N_5281,N_4419,N_4255);
nand U5282 (N_5282,N_4345,N_4981);
or U5283 (N_5283,N_4008,N_4632);
nor U5284 (N_5284,N_4782,N_4739);
and U5285 (N_5285,N_4364,N_4319);
nor U5286 (N_5286,N_4388,N_4952);
nor U5287 (N_5287,N_4509,N_4278);
or U5288 (N_5288,N_4810,N_4495);
nor U5289 (N_5289,N_4112,N_4644);
and U5290 (N_5290,N_4508,N_4816);
nor U5291 (N_5291,N_4078,N_4930);
xor U5292 (N_5292,N_4482,N_4964);
or U5293 (N_5293,N_4978,N_4517);
and U5294 (N_5294,N_4858,N_4692);
nand U5295 (N_5295,N_4987,N_4860);
or U5296 (N_5296,N_4211,N_4392);
xor U5297 (N_5297,N_4773,N_4218);
nor U5298 (N_5298,N_4296,N_4840);
and U5299 (N_5299,N_4904,N_4725);
xnor U5300 (N_5300,N_4755,N_4358);
xor U5301 (N_5301,N_4627,N_4581);
and U5302 (N_5302,N_4737,N_4790);
nor U5303 (N_5303,N_4556,N_4065);
nor U5304 (N_5304,N_4237,N_4156);
and U5305 (N_5305,N_4929,N_4886);
nand U5306 (N_5306,N_4039,N_4803);
xnor U5307 (N_5307,N_4818,N_4871);
and U5308 (N_5308,N_4269,N_4705);
nand U5309 (N_5309,N_4230,N_4184);
xor U5310 (N_5310,N_4355,N_4826);
nand U5311 (N_5311,N_4135,N_4786);
xnor U5312 (N_5312,N_4379,N_4195);
nand U5313 (N_5313,N_4796,N_4159);
nor U5314 (N_5314,N_4936,N_4165);
nor U5315 (N_5315,N_4335,N_4387);
nor U5316 (N_5316,N_4767,N_4573);
xor U5317 (N_5317,N_4917,N_4050);
nor U5318 (N_5318,N_4813,N_4285);
nand U5319 (N_5319,N_4324,N_4764);
or U5320 (N_5320,N_4950,N_4522);
xor U5321 (N_5321,N_4061,N_4703);
nand U5322 (N_5322,N_4530,N_4596);
or U5323 (N_5323,N_4223,N_4926);
xnor U5324 (N_5324,N_4990,N_4139);
and U5325 (N_5325,N_4483,N_4281);
nor U5326 (N_5326,N_4853,N_4505);
or U5327 (N_5327,N_4036,N_4717);
nand U5328 (N_5328,N_4114,N_4044);
nand U5329 (N_5329,N_4804,N_4761);
nand U5330 (N_5330,N_4315,N_4013);
nand U5331 (N_5331,N_4792,N_4811);
nor U5332 (N_5332,N_4132,N_4338);
and U5333 (N_5333,N_4242,N_4350);
xnor U5334 (N_5334,N_4048,N_4831);
nand U5335 (N_5335,N_4888,N_4848);
xnor U5336 (N_5336,N_4833,N_4143);
nor U5337 (N_5337,N_4309,N_4682);
nor U5338 (N_5338,N_4216,N_4280);
nor U5339 (N_5339,N_4733,N_4783);
nor U5340 (N_5340,N_4582,N_4587);
or U5341 (N_5341,N_4943,N_4444);
nand U5342 (N_5342,N_4329,N_4789);
or U5343 (N_5343,N_4512,N_4152);
xor U5344 (N_5344,N_4346,N_4564);
nand U5345 (N_5345,N_4322,N_4228);
or U5346 (N_5346,N_4464,N_4635);
and U5347 (N_5347,N_4404,N_4809);
or U5348 (N_5348,N_4439,N_4389);
nand U5349 (N_5349,N_4119,N_4974);
nor U5350 (N_5350,N_4599,N_4523);
nor U5351 (N_5351,N_4298,N_4844);
nand U5352 (N_5352,N_4117,N_4829);
or U5353 (N_5353,N_4748,N_4386);
or U5354 (N_5354,N_4501,N_4054);
and U5355 (N_5355,N_4484,N_4053);
nor U5356 (N_5356,N_4654,N_4680);
xor U5357 (N_5357,N_4137,N_4283);
or U5358 (N_5358,N_4639,N_4424);
nand U5359 (N_5359,N_4727,N_4047);
and U5360 (N_5360,N_4339,N_4145);
nand U5361 (N_5361,N_4188,N_4841);
or U5362 (N_5362,N_4747,N_4891);
nor U5363 (N_5363,N_4547,N_4440);
or U5364 (N_5364,N_4201,N_4541);
nand U5365 (N_5365,N_4527,N_4301);
and U5366 (N_5366,N_4207,N_4788);
and U5367 (N_5367,N_4295,N_4706);
nor U5368 (N_5368,N_4264,N_4136);
nor U5369 (N_5369,N_4928,N_4437);
xnor U5370 (N_5370,N_4690,N_4925);
nand U5371 (N_5371,N_4076,N_4618);
xnor U5372 (N_5372,N_4370,N_4671);
and U5373 (N_5373,N_4317,N_4344);
or U5374 (N_5374,N_4225,N_4757);
xor U5375 (N_5375,N_4247,N_4038);
and U5376 (N_5376,N_4842,N_4125);
and U5377 (N_5377,N_4960,N_4957);
xnor U5378 (N_5378,N_4341,N_4490);
or U5379 (N_5379,N_4020,N_4023);
and U5380 (N_5380,N_4890,N_4834);
and U5381 (N_5381,N_4595,N_4356);
or U5382 (N_5382,N_4771,N_4421);
xor U5383 (N_5383,N_4812,N_4548);
and U5384 (N_5384,N_4202,N_4756);
nand U5385 (N_5385,N_4610,N_4372);
xnor U5386 (N_5386,N_4019,N_4127);
nand U5387 (N_5387,N_4799,N_4390);
or U5388 (N_5388,N_4878,N_4655);
or U5389 (N_5389,N_4880,N_4998);
nand U5390 (N_5390,N_4588,N_4713);
or U5391 (N_5391,N_4472,N_4614);
nand U5392 (N_5392,N_4343,N_4307);
or U5393 (N_5393,N_4997,N_4565);
xnor U5394 (N_5394,N_4856,N_4908);
nand U5395 (N_5395,N_4913,N_4765);
or U5396 (N_5396,N_4575,N_4290);
nand U5397 (N_5397,N_4475,N_4651);
nor U5398 (N_5398,N_4172,N_4972);
or U5399 (N_5399,N_4807,N_4198);
xnor U5400 (N_5400,N_4899,N_4539);
and U5401 (N_5401,N_4313,N_4312);
and U5402 (N_5402,N_4306,N_4519);
nand U5403 (N_5403,N_4738,N_4215);
xnor U5404 (N_5404,N_4151,N_4697);
nand U5405 (N_5405,N_4099,N_4944);
xnor U5406 (N_5406,N_4999,N_4363);
or U5407 (N_5407,N_4458,N_4231);
nand U5408 (N_5408,N_4758,N_4535);
and U5409 (N_5409,N_4254,N_4004);
or U5410 (N_5410,N_4825,N_4679);
xor U5411 (N_5411,N_4694,N_4445);
nor U5412 (N_5412,N_4615,N_4538);
xnor U5413 (N_5413,N_4593,N_4657);
and U5414 (N_5414,N_4031,N_4684);
xor U5415 (N_5415,N_4634,N_4759);
or U5416 (N_5416,N_4146,N_4867);
nor U5417 (N_5417,N_4947,N_4432);
and U5418 (N_5418,N_4569,N_4711);
or U5419 (N_5419,N_4478,N_4249);
or U5420 (N_5420,N_4361,N_4591);
nand U5421 (N_5421,N_4652,N_4770);
nor U5422 (N_5422,N_4613,N_4975);
and U5423 (N_5423,N_4481,N_4704);
or U5424 (N_5424,N_4274,N_4474);
xor U5425 (N_5425,N_4641,N_4412);
or U5426 (N_5426,N_4353,N_4914);
and U5427 (N_5427,N_4683,N_4808);
or U5428 (N_5428,N_4935,N_4663);
nor U5429 (N_5429,N_4395,N_4665);
nand U5430 (N_5430,N_4621,N_4982);
and U5431 (N_5431,N_4066,N_4768);
and U5432 (N_5432,N_4628,N_4126);
or U5433 (N_5433,N_4664,N_4124);
nor U5434 (N_5434,N_4086,N_4623);
or U5435 (N_5435,N_4336,N_4331);
xnor U5436 (N_5436,N_4933,N_4170);
nand U5437 (N_5437,N_4121,N_4907);
and U5438 (N_5438,N_4067,N_4991);
xnor U5439 (N_5439,N_4168,N_4055);
nor U5440 (N_5440,N_4958,N_4229);
xnor U5441 (N_5441,N_4780,N_4217);
xor U5442 (N_5442,N_4658,N_4077);
nand U5443 (N_5443,N_4749,N_4859);
nor U5444 (N_5444,N_4968,N_4178);
and U5445 (N_5445,N_4330,N_4754);
nand U5446 (N_5446,N_4089,N_4730);
xnor U5447 (N_5447,N_4400,N_4212);
nor U5448 (N_5448,N_4592,N_4208);
nor U5449 (N_5449,N_4932,N_4656);
nand U5450 (N_5450,N_4630,N_4088);
nand U5451 (N_5451,N_4303,N_4133);
nand U5452 (N_5452,N_4497,N_4110);
or U5453 (N_5453,N_4762,N_4620);
xor U5454 (N_5454,N_4645,N_4081);
or U5455 (N_5455,N_4493,N_4774);
nor U5456 (N_5456,N_4033,N_4450);
xor U5457 (N_5457,N_4286,N_4751);
xor U5458 (N_5458,N_4045,N_4709);
xnor U5459 (N_5459,N_4693,N_4100);
nand U5460 (N_5460,N_4956,N_4138);
and U5461 (N_5461,N_4687,N_4521);
nor U5462 (N_5462,N_4204,N_4083);
xnor U5463 (N_5463,N_4221,N_4070);
xor U5464 (N_5464,N_4785,N_4141);
xor U5465 (N_5465,N_4580,N_4897);
or U5466 (N_5466,N_4479,N_4199);
and U5467 (N_5467,N_4477,N_4667);
or U5468 (N_5468,N_4598,N_4563);
and U5469 (N_5469,N_4191,N_4839);
and U5470 (N_5470,N_4906,N_4643);
nand U5471 (N_5471,N_4153,N_4326);
or U5472 (N_5472,N_4698,N_4232);
nor U5473 (N_5473,N_4377,N_4452);
and U5474 (N_5474,N_4150,N_4611);
nand U5475 (N_5475,N_4720,N_4500);
nand U5476 (N_5476,N_4916,N_4485);
and U5477 (N_5477,N_4712,N_4676);
nor U5478 (N_5478,N_4279,N_4583);
and U5479 (N_5479,N_4300,N_4542);
nor U5480 (N_5480,N_4383,N_4918);
and U5481 (N_5481,N_4401,N_4021);
nor U5482 (N_5482,N_4633,N_4566);
xor U5483 (N_5483,N_4194,N_4025);
or U5484 (N_5484,N_4827,N_4327);
nand U5485 (N_5485,N_4261,N_4646);
xnor U5486 (N_5486,N_4600,N_4735);
and U5487 (N_5487,N_4716,N_4985);
xnor U5488 (N_5488,N_4882,N_4425);
xnor U5489 (N_5489,N_4873,N_4863);
and U5490 (N_5490,N_4287,N_4861);
nor U5491 (N_5491,N_4342,N_4962);
nor U5492 (N_5492,N_4068,N_4689);
nor U5493 (N_5493,N_4870,N_4075);
and U5494 (N_5494,N_4659,N_4011);
xor U5495 (N_5495,N_4551,N_4396);
nor U5496 (N_5496,N_4461,N_4715);
or U5497 (N_5497,N_4515,N_4961);
nand U5498 (N_5498,N_4609,N_4568);
and U5499 (N_5499,N_4570,N_4016);
or U5500 (N_5500,N_4979,N_4175);
nand U5501 (N_5501,N_4948,N_4356);
nor U5502 (N_5502,N_4798,N_4069);
nand U5503 (N_5503,N_4255,N_4699);
nand U5504 (N_5504,N_4875,N_4594);
nand U5505 (N_5505,N_4745,N_4660);
and U5506 (N_5506,N_4195,N_4385);
nand U5507 (N_5507,N_4672,N_4756);
nand U5508 (N_5508,N_4957,N_4454);
nor U5509 (N_5509,N_4042,N_4482);
and U5510 (N_5510,N_4952,N_4561);
and U5511 (N_5511,N_4717,N_4753);
or U5512 (N_5512,N_4548,N_4628);
xnor U5513 (N_5513,N_4140,N_4038);
and U5514 (N_5514,N_4613,N_4003);
and U5515 (N_5515,N_4197,N_4935);
nand U5516 (N_5516,N_4450,N_4007);
nand U5517 (N_5517,N_4722,N_4027);
nand U5518 (N_5518,N_4621,N_4698);
xor U5519 (N_5519,N_4773,N_4071);
nor U5520 (N_5520,N_4844,N_4384);
and U5521 (N_5521,N_4362,N_4496);
and U5522 (N_5522,N_4589,N_4177);
and U5523 (N_5523,N_4729,N_4762);
nand U5524 (N_5524,N_4324,N_4497);
and U5525 (N_5525,N_4498,N_4171);
xor U5526 (N_5526,N_4560,N_4659);
xor U5527 (N_5527,N_4765,N_4082);
nor U5528 (N_5528,N_4171,N_4998);
and U5529 (N_5529,N_4274,N_4232);
xnor U5530 (N_5530,N_4521,N_4590);
or U5531 (N_5531,N_4687,N_4995);
or U5532 (N_5532,N_4782,N_4468);
xor U5533 (N_5533,N_4614,N_4773);
nand U5534 (N_5534,N_4306,N_4090);
and U5535 (N_5535,N_4611,N_4344);
nor U5536 (N_5536,N_4918,N_4754);
xor U5537 (N_5537,N_4296,N_4132);
and U5538 (N_5538,N_4911,N_4013);
xor U5539 (N_5539,N_4941,N_4062);
or U5540 (N_5540,N_4690,N_4462);
nor U5541 (N_5541,N_4002,N_4654);
and U5542 (N_5542,N_4356,N_4299);
or U5543 (N_5543,N_4404,N_4678);
xor U5544 (N_5544,N_4552,N_4481);
xor U5545 (N_5545,N_4031,N_4078);
and U5546 (N_5546,N_4350,N_4618);
nor U5547 (N_5547,N_4194,N_4953);
nand U5548 (N_5548,N_4658,N_4287);
and U5549 (N_5549,N_4784,N_4605);
nor U5550 (N_5550,N_4703,N_4311);
nor U5551 (N_5551,N_4722,N_4616);
xor U5552 (N_5552,N_4502,N_4639);
nor U5553 (N_5553,N_4173,N_4172);
or U5554 (N_5554,N_4874,N_4792);
nor U5555 (N_5555,N_4311,N_4331);
xor U5556 (N_5556,N_4699,N_4257);
and U5557 (N_5557,N_4286,N_4953);
and U5558 (N_5558,N_4144,N_4605);
and U5559 (N_5559,N_4303,N_4486);
and U5560 (N_5560,N_4950,N_4612);
nand U5561 (N_5561,N_4438,N_4268);
and U5562 (N_5562,N_4849,N_4171);
xor U5563 (N_5563,N_4909,N_4258);
nand U5564 (N_5564,N_4302,N_4603);
xor U5565 (N_5565,N_4210,N_4986);
and U5566 (N_5566,N_4032,N_4132);
nor U5567 (N_5567,N_4775,N_4548);
and U5568 (N_5568,N_4083,N_4799);
nor U5569 (N_5569,N_4939,N_4384);
or U5570 (N_5570,N_4671,N_4665);
nor U5571 (N_5571,N_4381,N_4730);
xor U5572 (N_5572,N_4537,N_4162);
and U5573 (N_5573,N_4474,N_4725);
xnor U5574 (N_5574,N_4256,N_4151);
or U5575 (N_5575,N_4306,N_4122);
nand U5576 (N_5576,N_4817,N_4429);
or U5577 (N_5577,N_4989,N_4919);
and U5578 (N_5578,N_4562,N_4899);
nand U5579 (N_5579,N_4302,N_4124);
nand U5580 (N_5580,N_4920,N_4974);
and U5581 (N_5581,N_4895,N_4255);
and U5582 (N_5582,N_4449,N_4007);
or U5583 (N_5583,N_4149,N_4142);
xnor U5584 (N_5584,N_4517,N_4833);
or U5585 (N_5585,N_4956,N_4614);
nor U5586 (N_5586,N_4552,N_4366);
nand U5587 (N_5587,N_4394,N_4135);
nor U5588 (N_5588,N_4590,N_4844);
xor U5589 (N_5589,N_4126,N_4458);
nand U5590 (N_5590,N_4594,N_4724);
or U5591 (N_5591,N_4956,N_4423);
xor U5592 (N_5592,N_4075,N_4436);
nand U5593 (N_5593,N_4896,N_4570);
and U5594 (N_5594,N_4936,N_4245);
nor U5595 (N_5595,N_4092,N_4018);
nand U5596 (N_5596,N_4317,N_4631);
nand U5597 (N_5597,N_4759,N_4998);
and U5598 (N_5598,N_4114,N_4230);
or U5599 (N_5599,N_4654,N_4016);
or U5600 (N_5600,N_4099,N_4100);
or U5601 (N_5601,N_4680,N_4934);
and U5602 (N_5602,N_4344,N_4913);
nand U5603 (N_5603,N_4659,N_4973);
or U5604 (N_5604,N_4101,N_4982);
nor U5605 (N_5605,N_4761,N_4815);
nor U5606 (N_5606,N_4298,N_4593);
or U5607 (N_5607,N_4570,N_4643);
xnor U5608 (N_5608,N_4632,N_4455);
or U5609 (N_5609,N_4068,N_4369);
and U5610 (N_5610,N_4859,N_4792);
and U5611 (N_5611,N_4895,N_4705);
or U5612 (N_5612,N_4121,N_4252);
xor U5613 (N_5613,N_4837,N_4982);
nor U5614 (N_5614,N_4572,N_4440);
nand U5615 (N_5615,N_4806,N_4279);
nand U5616 (N_5616,N_4936,N_4133);
and U5617 (N_5617,N_4501,N_4570);
xor U5618 (N_5618,N_4026,N_4494);
nand U5619 (N_5619,N_4557,N_4401);
xnor U5620 (N_5620,N_4776,N_4200);
and U5621 (N_5621,N_4646,N_4086);
or U5622 (N_5622,N_4641,N_4396);
nor U5623 (N_5623,N_4271,N_4521);
nand U5624 (N_5624,N_4116,N_4567);
xnor U5625 (N_5625,N_4862,N_4609);
and U5626 (N_5626,N_4600,N_4522);
nor U5627 (N_5627,N_4914,N_4597);
or U5628 (N_5628,N_4231,N_4602);
or U5629 (N_5629,N_4505,N_4046);
nand U5630 (N_5630,N_4909,N_4181);
xnor U5631 (N_5631,N_4930,N_4186);
xor U5632 (N_5632,N_4225,N_4537);
and U5633 (N_5633,N_4626,N_4689);
nor U5634 (N_5634,N_4380,N_4410);
xnor U5635 (N_5635,N_4070,N_4873);
nor U5636 (N_5636,N_4523,N_4476);
and U5637 (N_5637,N_4401,N_4031);
xnor U5638 (N_5638,N_4976,N_4592);
nor U5639 (N_5639,N_4145,N_4932);
xor U5640 (N_5640,N_4873,N_4218);
nor U5641 (N_5641,N_4639,N_4439);
nand U5642 (N_5642,N_4890,N_4945);
or U5643 (N_5643,N_4533,N_4838);
xnor U5644 (N_5644,N_4433,N_4964);
nand U5645 (N_5645,N_4573,N_4091);
or U5646 (N_5646,N_4160,N_4923);
or U5647 (N_5647,N_4093,N_4896);
nor U5648 (N_5648,N_4436,N_4872);
and U5649 (N_5649,N_4433,N_4081);
nor U5650 (N_5650,N_4774,N_4879);
xor U5651 (N_5651,N_4649,N_4098);
or U5652 (N_5652,N_4735,N_4721);
and U5653 (N_5653,N_4342,N_4578);
or U5654 (N_5654,N_4966,N_4093);
nor U5655 (N_5655,N_4556,N_4769);
xnor U5656 (N_5656,N_4258,N_4654);
nor U5657 (N_5657,N_4848,N_4240);
nor U5658 (N_5658,N_4310,N_4323);
xnor U5659 (N_5659,N_4405,N_4359);
xnor U5660 (N_5660,N_4645,N_4789);
or U5661 (N_5661,N_4232,N_4318);
nor U5662 (N_5662,N_4639,N_4433);
nor U5663 (N_5663,N_4478,N_4018);
or U5664 (N_5664,N_4237,N_4669);
xnor U5665 (N_5665,N_4391,N_4210);
xnor U5666 (N_5666,N_4610,N_4961);
nor U5667 (N_5667,N_4867,N_4239);
nor U5668 (N_5668,N_4281,N_4316);
nand U5669 (N_5669,N_4506,N_4464);
xor U5670 (N_5670,N_4438,N_4502);
or U5671 (N_5671,N_4365,N_4589);
xnor U5672 (N_5672,N_4282,N_4730);
xnor U5673 (N_5673,N_4820,N_4176);
nor U5674 (N_5674,N_4411,N_4566);
nor U5675 (N_5675,N_4489,N_4042);
nand U5676 (N_5676,N_4986,N_4328);
and U5677 (N_5677,N_4371,N_4137);
and U5678 (N_5678,N_4007,N_4253);
nor U5679 (N_5679,N_4442,N_4818);
or U5680 (N_5680,N_4375,N_4084);
nor U5681 (N_5681,N_4367,N_4568);
and U5682 (N_5682,N_4970,N_4273);
nand U5683 (N_5683,N_4454,N_4472);
and U5684 (N_5684,N_4937,N_4378);
or U5685 (N_5685,N_4056,N_4448);
nor U5686 (N_5686,N_4690,N_4828);
xnor U5687 (N_5687,N_4527,N_4164);
xor U5688 (N_5688,N_4148,N_4998);
or U5689 (N_5689,N_4472,N_4189);
and U5690 (N_5690,N_4117,N_4310);
nand U5691 (N_5691,N_4310,N_4668);
nand U5692 (N_5692,N_4189,N_4469);
xor U5693 (N_5693,N_4462,N_4067);
nor U5694 (N_5694,N_4234,N_4763);
and U5695 (N_5695,N_4291,N_4982);
or U5696 (N_5696,N_4077,N_4713);
nand U5697 (N_5697,N_4409,N_4923);
xor U5698 (N_5698,N_4881,N_4969);
xor U5699 (N_5699,N_4814,N_4358);
and U5700 (N_5700,N_4160,N_4890);
nor U5701 (N_5701,N_4026,N_4352);
nor U5702 (N_5702,N_4181,N_4793);
or U5703 (N_5703,N_4408,N_4310);
or U5704 (N_5704,N_4758,N_4512);
xor U5705 (N_5705,N_4375,N_4350);
nand U5706 (N_5706,N_4915,N_4136);
nand U5707 (N_5707,N_4589,N_4382);
and U5708 (N_5708,N_4464,N_4674);
or U5709 (N_5709,N_4664,N_4659);
xnor U5710 (N_5710,N_4449,N_4193);
xnor U5711 (N_5711,N_4888,N_4364);
nor U5712 (N_5712,N_4855,N_4657);
xnor U5713 (N_5713,N_4063,N_4874);
and U5714 (N_5714,N_4783,N_4739);
and U5715 (N_5715,N_4399,N_4363);
or U5716 (N_5716,N_4779,N_4883);
nor U5717 (N_5717,N_4889,N_4589);
or U5718 (N_5718,N_4087,N_4025);
nor U5719 (N_5719,N_4253,N_4793);
nand U5720 (N_5720,N_4990,N_4983);
nor U5721 (N_5721,N_4021,N_4972);
nand U5722 (N_5722,N_4233,N_4027);
xnor U5723 (N_5723,N_4574,N_4756);
nor U5724 (N_5724,N_4780,N_4603);
xnor U5725 (N_5725,N_4030,N_4066);
and U5726 (N_5726,N_4232,N_4322);
and U5727 (N_5727,N_4480,N_4240);
and U5728 (N_5728,N_4137,N_4696);
xor U5729 (N_5729,N_4311,N_4345);
xnor U5730 (N_5730,N_4697,N_4656);
xnor U5731 (N_5731,N_4575,N_4180);
or U5732 (N_5732,N_4942,N_4161);
nor U5733 (N_5733,N_4886,N_4624);
or U5734 (N_5734,N_4939,N_4075);
nand U5735 (N_5735,N_4029,N_4330);
or U5736 (N_5736,N_4808,N_4174);
and U5737 (N_5737,N_4840,N_4772);
or U5738 (N_5738,N_4635,N_4819);
or U5739 (N_5739,N_4039,N_4266);
nor U5740 (N_5740,N_4461,N_4655);
nor U5741 (N_5741,N_4672,N_4769);
xnor U5742 (N_5742,N_4982,N_4870);
and U5743 (N_5743,N_4980,N_4380);
nor U5744 (N_5744,N_4244,N_4303);
nor U5745 (N_5745,N_4541,N_4835);
nor U5746 (N_5746,N_4378,N_4684);
xor U5747 (N_5747,N_4873,N_4994);
xnor U5748 (N_5748,N_4164,N_4048);
or U5749 (N_5749,N_4696,N_4362);
and U5750 (N_5750,N_4777,N_4864);
nand U5751 (N_5751,N_4462,N_4060);
xor U5752 (N_5752,N_4186,N_4803);
nand U5753 (N_5753,N_4657,N_4673);
and U5754 (N_5754,N_4494,N_4855);
and U5755 (N_5755,N_4623,N_4582);
xnor U5756 (N_5756,N_4102,N_4981);
xnor U5757 (N_5757,N_4693,N_4911);
nor U5758 (N_5758,N_4032,N_4099);
nor U5759 (N_5759,N_4061,N_4727);
xnor U5760 (N_5760,N_4662,N_4203);
or U5761 (N_5761,N_4421,N_4711);
nor U5762 (N_5762,N_4803,N_4899);
or U5763 (N_5763,N_4238,N_4297);
or U5764 (N_5764,N_4950,N_4960);
or U5765 (N_5765,N_4852,N_4296);
nand U5766 (N_5766,N_4897,N_4372);
and U5767 (N_5767,N_4130,N_4949);
nand U5768 (N_5768,N_4618,N_4060);
xnor U5769 (N_5769,N_4994,N_4997);
and U5770 (N_5770,N_4492,N_4827);
nand U5771 (N_5771,N_4787,N_4976);
and U5772 (N_5772,N_4050,N_4038);
or U5773 (N_5773,N_4027,N_4119);
nor U5774 (N_5774,N_4619,N_4027);
or U5775 (N_5775,N_4714,N_4507);
or U5776 (N_5776,N_4003,N_4593);
nor U5777 (N_5777,N_4544,N_4197);
or U5778 (N_5778,N_4471,N_4757);
or U5779 (N_5779,N_4740,N_4221);
and U5780 (N_5780,N_4705,N_4649);
nor U5781 (N_5781,N_4902,N_4350);
nor U5782 (N_5782,N_4213,N_4632);
and U5783 (N_5783,N_4799,N_4945);
nand U5784 (N_5784,N_4350,N_4781);
xnor U5785 (N_5785,N_4957,N_4858);
nand U5786 (N_5786,N_4518,N_4591);
xnor U5787 (N_5787,N_4979,N_4049);
and U5788 (N_5788,N_4010,N_4376);
xor U5789 (N_5789,N_4445,N_4164);
nand U5790 (N_5790,N_4523,N_4973);
or U5791 (N_5791,N_4907,N_4647);
nand U5792 (N_5792,N_4619,N_4189);
or U5793 (N_5793,N_4913,N_4060);
nor U5794 (N_5794,N_4303,N_4496);
xor U5795 (N_5795,N_4818,N_4838);
and U5796 (N_5796,N_4282,N_4959);
and U5797 (N_5797,N_4578,N_4785);
nor U5798 (N_5798,N_4305,N_4695);
and U5799 (N_5799,N_4370,N_4740);
xor U5800 (N_5800,N_4587,N_4501);
nand U5801 (N_5801,N_4807,N_4808);
nand U5802 (N_5802,N_4666,N_4263);
or U5803 (N_5803,N_4783,N_4768);
nor U5804 (N_5804,N_4545,N_4134);
nor U5805 (N_5805,N_4085,N_4995);
and U5806 (N_5806,N_4171,N_4704);
nor U5807 (N_5807,N_4323,N_4341);
and U5808 (N_5808,N_4006,N_4343);
or U5809 (N_5809,N_4810,N_4144);
or U5810 (N_5810,N_4003,N_4422);
and U5811 (N_5811,N_4640,N_4571);
or U5812 (N_5812,N_4923,N_4786);
or U5813 (N_5813,N_4440,N_4624);
xor U5814 (N_5814,N_4994,N_4497);
and U5815 (N_5815,N_4122,N_4892);
nand U5816 (N_5816,N_4825,N_4522);
or U5817 (N_5817,N_4491,N_4096);
and U5818 (N_5818,N_4112,N_4094);
or U5819 (N_5819,N_4183,N_4067);
xnor U5820 (N_5820,N_4116,N_4272);
nand U5821 (N_5821,N_4178,N_4289);
nor U5822 (N_5822,N_4034,N_4777);
and U5823 (N_5823,N_4060,N_4989);
nor U5824 (N_5824,N_4253,N_4871);
and U5825 (N_5825,N_4409,N_4924);
and U5826 (N_5826,N_4045,N_4304);
or U5827 (N_5827,N_4270,N_4959);
xor U5828 (N_5828,N_4902,N_4951);
xor U5829 (N_5829,N_4944,N_4932);
or U5830 (N_5830,N_4009,N_4673);
nand U5831 (N_5831,N_4548,N_4851);
xor U5832 (N_5832,N_4195,N_4173);
xor U5833 (N_5833,N_4902,N_4282);
xor U5834 (N_5834,N_4659,N_4401);
nand U5835 (N_5835,N_4402,N_4736);
xnor U5836 (N_5836,N_4921,N_4688);
or U5837 (N_5837,N_4217,N_4370);
nor U5838 (N_5838,N_4682,N_4041);
xnor U5839 (N_5839,N_4651,N_4931);
and U5840 (N_5840,N_4109,N_4862);
and U5841 (N_5841,N_4931,N_4962);
nand U5842 (N_5842,N_4258,N_4872);
and U5843 (N_5843,N_4391,N_4717);
nor U5844 (N_5844,N_4736,N_4949);
or U5845 (N_5845,N_4547,N_4801);
or U5846 (N_5846,N_4215,N_4375);
nand U5847 (N_5847,N_4085,N_4201);
nor U5848 (N_5848,N_4711,N_4055);
nor U5849 (N_5849,N_4804,N_4083);
xor U5850 (N_5850,N_4485,N_4882);
nand U5851 (N_5851,N_4363,N_4046);
and U5852 (N_5852,N_4166,N_4020);
nor U5853 (N_5853,N_4761,N_4498);
and U5854 (N_5854,N_4825,N_4324);
nand U5855 (N_5855,N_4686,N_4671);
and U5856 (N_5856,N_4737,N_4939);
nand U5857 (N_5857,N_4924,N_4848);
xor U5858 (N_5858,N_4323,N_4037);
xnor U5859 (N_5859,N_4071,N_4535);
nor U5860 (N_5860,N_4825,N_4725);
or U5861 (N_5861,N_4871,N_4722);
or U5862 (N_5862,N_4162,N_4801);
or U5863 (N_5863,N_4152,N_4049);
or U5864 (N_5864,N_4103,N_4980);
nand U5865 (N_5865,N_4732,N_4199);
xnor U5866 (N_5866,N_4157,N_4857);
nand U5867 (N_5867,N_4152,N_4036);
nand U5868 (N_5868,N_4105,N_4875);
xor U5869 (N_5869,N_4705,N_4291);
or U5870 (N_5870,N_4862,N_4087);
nand U5871 (N_5871,N_4005,N_4485);
xnor U5872 (N_5872,N_4708,N_4974);
or U5873 (N_5873,N_4164,N_4233);
or U5874 (N_5874,N_4463,N_4610);
xnor U5875 (N_5875,N_4887,N_4012);
or U5876 (N_5876,N_4136,N_4929);
nand U5877 (N_5877,N_4919,N_4789);
nand U5878 (N_5878,N_4731,N_4035);
nand U5879 (N_5879,N_4252,N_4845);
nor U5880 (N_5880,N_4456,N_4761);
nand U5881 (N_5881,N_4899,N_4549);
and U5882 (N_5882,N_4911,N_4033);
nor U5883 (N_5883,N_4471,N_4640);
and U5884 (N_5884,N_4045,N_4094);
xnor U5885 (N_5885,N_4138,N_4434);
or U5886 (N_5886,N_4781,N_4345);
nand U5887 (N_5887,N_4230,N_4182);
nor U5888 (N_5888,N_4014,N_4372);
and U5889 (N_5889,N_4708,N_4591);
and U5890 (N_5890,N_4546,N_4763);
xor U5891 (N_5891,N_4496,N_4709);
or U5892 (N_5892,N_4761,N_4558);
xor U5893 (N_5893,N_4941,N_4807);
or U5894 (N_5894,N_4136,N_4288);
nor U5895 (N_5895,N_4394,N_4640);
or U5896 (N_5896,N_4329,N_4576);
and U5897 (N_5897,N_4000,N_4059);
or U5898 (N_5898,N_4291,N_4665);
xor U5899 (N_5899,N_4026,N_4715);
xor U5900 (N_5900,N_4641,N_4636);
and U5901 (N_5901,N_4018,N_4234);
and U5902 (N_5902,N_4120,N_4054);
nand U5903 (N_5903,N_4428,N_4483);
nand U5904 (N_5904,N_4547,N_4191);
xor U5905 (N_5905,N_4364,N_4186);
or U5906 (N_5906,N_4744,N_4131);
and U5907 (N_5907,N_4086,N_4842);
nor U5908 (N_5908,N_4229,N_4088);
and U5909 (N_5909,N_4823,N_4383);
nand U5910 (N_5910,N_4107,N_4875);
or U5911 (N_5911,N_4104,N_4700);
nand U5912 (N_5912,N_4039,N_4905);
nand U5913 (N_5913,N_4206,N_4007);
nor U5914 (N_5914,N_4350,N_4240);
xnor U5915 (N_5915,N_4346,N_4312);
xnor U5916 (N_5916,N_4236,N_4947);
nor U5917 (N_5917,N_4431,N_4100);
nor U5918 (N_5918,N_4707,N_4120);
and U5919 (N_5919,N_4235,N_4501);
xor U5920 (N_5920,N_4325,N_4131);
or U5921 (N_5921,N_4375,N_4352);
xnor U5922 (N_5922,N_4820,N_4036);
xnor U5923 (N_5923,N_4461,N_4181);
and U5924 (N_5924,N_4172,N_4182);
and U5925 (N_5925,N_4270,N_4970);
or U5926 (N_5926,N_4198,N_4844);
nor U5927 (N_5927,N_4462,N_4755);
nor U5928 (N_5928,N_4699,N_4635);
nor U5929 (N_5929,N_4924,N_4522);
xor U5930 (N_5930,N_4333,N_4885);
nor U5931 (N_5931,N_4721,N_4282);
nand U5932 (N_5932,N_4436,N_4919);
xor U5933 (N_5933,N_4910,N_4027);
or U5934 (N_5934,N_4589,N_4328);
and U5935 (N_5935,N_4368,N_4699);
and U5936 (N_5936,N_4810,N_4464);
nor U5937 (N_5937,N_4135,N_4241);
and U5938 (N_5938,N_4790,N_4049);
nand U5939 (N_5939,N_4300,N_4008);
and U5940 (N_5940,N_4889,N_4635);
or U5941 (N_5941,N_4472,N_4180);
nor U5942 (N_5942,N_4604,N_4706);
nand U5943 (N_5943,N_4264,N_4718);
xor U5944 (N_5944,N_4788,N_4685);
or U5945 (N_5945,N_4772,N_4452);
xnor U5946 (N_5946,N_4037,N_4469);
or U5947 (N_5947,N_4991,N_4205);
or U5948 (N_5948,N_4184,N_4015);
nor U5949 (N_5949,N_4901,N_4907);
nor U5950 (N_5950,N_4333,N_4599);
nand U5951 (N_5951,N_4410,N_4615);
xnor U5952 (N_5952,N_4247,N_4680);
nand U5953 (N_5953,N_4506,N_4986);
or U5954 (N_5954,N_4021,N_4867);
nor U5955 (N_5955,N_4932,N_4836);
or U5956 (N_5956,N_4351,N_4985);
nand U5957 (N_5957,N_4742,N_4168);
and U5958 (N_5958,N_4451,N_4541);
nor U5959 (N_5959,N_4401,N_4243);
and U5960 (N_5960,N_4322,N_4064);
nor U5961 (N_5961,N_4699,N_4787);
nand U5962 (N_5962,N_4001,N_4998);
nor U5963 (N_5963,N_4286,N_4435);
nand U5964 (N_5964,N_4078,N_4132);
xnor U5965 (N_5965,N_4486,N_4905);
nand U5966 (N_5966,N_4218,N_4136);
or U5967 (N_5967,N_4468,N_4808);
or U5968 (N_5968,N_4257,N_4012);
or U5969 (N_5969,N_4127,N_4712);
and U5970 (N_5970,N_4388,N_4897);
nand U5971 (N_5971,N_4902,N_4889);
nand U5972 (N_5972,N_4711,N_4331);
nand U5973 (N_5973,N_4201,N_4586);
xor U5974 (N_5974,N_4799,N_4692);
or U5975 (N_5975,N_4826,N_4237);
nand U5976 (N_5976,N_4348,N_4244);
nand U5977 (N_5977,N_4364,N_4346);
nand U5978 (N_5978,N_4880,N_4390);
or U5979 (N_5979,N_4280,N_4844);
and U5980 (N_5980,N_4441,N_4445);
xnor U5981 (N_5981,N_4664,N_4716);
nor U5982 (N_5982,N_4288,N_4608);
nand U5983 (N_5983,N_4660,N_4367);
nand U5984 (N_5984,N_4615,N_4576);
and U5985 (N_5985,N_4230,N_4297);
nand U5986 (N_5986,N_4688,N_4289);
and U5987 (N_5987,N_4119,N_4732);
and U5988 (N_5988,N_4184,N_4200);
xnor U5989 (N_5989,N_4709,N_4065);
nor U5990 (N_5990,N_4597,N_4112);
xnor U5991 (N_5991,N_4090,N_4326);
xor U5992 (N_5992,N_4465,N_4650);
nor U5993 (N_5993,N_4158,N_4146);
nor U5994 (N_5994,N_4091,N_4997);
xor U5995 (N_5995,N_4872,N_4908);
xor U5996 (N_5996,N_4635,N_4138);
nand U5997 (N_5997,N_4676,N_4389);
nand U5998 (N_5998,N_4119,N_4314);
or U5999 (N_5999,N_4780,N_4032);
nand U6000 (N_6000,N_5767,N_5170);
nor U6001 (N_6001,N_5242,N_5139);
xor U6002 (N_6002,N_5707,N_5574);
or U6003 (N_6003,N_5416,N_5605);
nor U6004 (N_6004,N_5635,N_5428);
or U6005 (N_6005,N_5035,N_5917);
nor U6006 (N_6006,N_5010,N_5993);
nor U6007 (N_6007,N_5820,N_5697);
xor U6008 (N_6008,N_5183,N_5637);
and U6009 (N_6009,N_5281,N_5771);
or U6010 (N_6010,N_5163,N_5625);
nand U6011 (N_6011,N_5255,N_5476);
nand U6012 (N_6012,N_5586,N_5768);
nand U6013 (N_6013,N_5088,N_5250);
xor U6014 (N_6014,N_5075,N_5162);
or U6015 (N_6015,N_5016,N_5093);
and U6016 (N_6016,N_5916,N_5127);
nor U6017 (N_6017,N_5740,N_5340);
and U6018 (N_6018,N_5152,N_5046);
nor U6019 (N_6019,N_5232,N_5173);
nand U6020 (N_6020,N_5603,N_5188);
nor U6021 (N_6021,N_5439,N_5668);
xor U6022 (N_6022,N_5226,N_5903);
or U6023 (N_6023,N_5462,N_5276);
nand U6024 (N_6024,N_5481,N_5133);
and U6025 (N_6025,N_5224,N_5789);
nor U6026 (N_6026,N_5681,N_5876);
and U6027 (N_6027,N_5632,N_5470);
nor U6028 (N_6028,N_5248,N_5030);
nand U6029 (N_6029,N_5465,N_5736);
or U6030 (N_6030,N_5671,N_5089);
xor U6031 (N_6031,N_5990,N_5940);
nor U6032 (N_6032,N_5260,N_5129);
xnor U6033 (N_6033,N_5848,N_5892);
nand U6034 (N_6034,N_5786,N_5887);
nor U6035 (N_6035,N_5354,N_5832);
nor U6036 (N_6036,N_5794,N_5814);
nor U6037 (N_6037,N_5987,N_5816);
and U6038 (N_6038,N_5756,N_5377);
nor U6039 (N_6039,N_5651,N_5433);
nor U6040 (N_6040,N_5272,N_5639);
nand U6041 (N_6041,N_5414,N_5322);
nor U6042 (N_6042,N_5619,N_5998);
xor U6043 (N_6043,N_5544,N_5883);
nor U6044 (N_6044,N_5002,N_5338);
nand U6045 (N_6045,N_5763,N_5533);
xnor U6046 (N_6046,N_5967,N_5659);
nor U6047 (N_6047,N_5951,N_5634);
and U6048 (N_6048,N_5285,N_5724);
nor U6049 (N_6049,N_5692,N_5385);
nor U6050 (N_6050,N_5191,N_5400);
xor U6051 (N_6051,N_5563,N_5324);
nor U6052 (N_6052,N_5120,N_5755);
nand U6053 (N_6053,N_5304,N_5607);
xnor U6054 (N_6054,N_5980,N_5446);
or U6055 (N_6055,N_5334,N_5395);
nor U6056 (N_6056,N_5690,N_5107);
and U6057 (N_6057,N_5328,N_5040);
xnor U6058 (N_6058,N_5236,N_5508);
or U6059 (N_6059,N_5636,N_5344);
nand U6060 (N_6060,N_5283,N_5259);
and U6061 (N_6061,N_5207,N_5350);
and U6062 (N_6062,N_5512,N_5902);
nand U6063 (N_6063,N_5144,N_5646);
or U6064 (N_6064,N_5971,N_5679);
or U6065 (N_6065,N_5609,N_5796);
nand U6066 (N_6066,N_5238,N_5831);
nand U6067 (N_6067,N_5944,N_5857);
nor U6068 (N_6068,N_5023,N_5538);
nand U6069 (N_6069,N_5332,N_5580);
xor U6070 (N_6070,N_5858,N_5153);
nor U6071 (N_6071,N_5698,N_5743);
nor U6072 (N_6072,N_5026,N_5404);
xnor U6073 (N_6073,N_5059,N_5065);
nand U6074 (N_6074,N_5837,N_5128);
and U6075 (N_6075,N_5329,N_5031);
and U6076 (N_6076,N_5037,N_5119);
or U6077 (N_6077,N_5134,N_5114);
xnor U6078 (N_6078,N_5267,N_5559);
or U6079 (N_6079,N_5291,N_5901);
nand U6080 (N_6080,N_5367,N_5409);
nand U6081 (N_6081,N_5148,N_5199);
or U6082 (N_6082,N_5525,N_5363);
nand U6083 (N_6083,N_5182,N_5005);
nand U6084 (N_6084,N_5009,N_5906);
nor U6085 (N_6085,N_5176,N_5562);
or U6086 (N_6086,N_5561,N_5169);
nand U6087 (N_6087,N_5274,N_5444);
nor U6088 (N_6088,N_5359,N_5012);
or U6089 (N_6089,N_5578,N_5955);
nand U6090 (N_6090,N_5312,N_5209);
nor U6091 (N_6091,N_5801,N_5843);
and U6092 (N_6092,N_5985,N_5706);
and U6093 (N_6093,N_5104,N_5576);
xnor U6094 (N_6094,N_5371,N_5213);
xnor U6095 (N_6095,N_5808,N_5537);
nand U6096 (N_6096,N_5583,N_5131);
xnor U6097 (N_6097,N_5223,N_5598);
and U6098 (N_6098,N_5933,N_5282);
nor U6099 (N_6099,N_5000,N_5770);
nor U6100 (N_6100,N_5369,N_5214);
xnor U6101 (N_6101,N_5926,N_5029);
xor U6102 (N_6102,N_5345,N_5290);
nand U6103 (N_6103,N_5682,N_5752);
xor U6104 (N_6104,N_5667,N_5316);
or U6105 (N_6105,N_5573,N_5534);
nor U6106 (N_6106,N_5022,N_5571);
nor U6107 (N_6107,N_5500,N_5257);
xnor U6108 (N_6108,N_5048,N_5256);
nor U6109 (N_6109,N_5780,N_5092);
xor U6110 (N_6110,N_5785,N_5042);
nand U6111 (N_6111,N_5105,N_5497);
nor U6112 (N_6112,N_5196,N_5287);
xor U6113 (N_6113,N_5504,N_5230);
and U6114 (N_6114,N_5912,N_5301);
nand U6115 (N_6115,N_5723,N_5389);
or U6116 (N_6116,N_5856,N_5125);
or U6117 (N_6117,N_5498,N_5412);
and U6118 (N_6118,N_5014,N_5845);
nand U6119 (N_6119,N_5358,N_5977);
or U6120 (N_6120,N_5063,N_5529);
or U6121 (N_6121,N_5069,N_5479);
nor U6122 (N_6122,N_5981,N_5725);
xnor U6123 (N_6123,N_5013,N_5774);
xnor U6124 (N_6124,N_5860,N_5982);
and U6125 (N_6125,N_5136,N_5159);
and U6126 (N_6126,N_5517,N_5310);
nor U6127 (N_6127,N_5886,N_5746);
or U6128 (N_6128,N_5643,N_5566);
nor U6129 (N_6129,N_5017,N_5346);
or U6130 (N_6130,N_5868,N_5008);
nor U6131 (N_6131,N_5406,N_5383);
nand U6132 (N_6132,N_5070,N_5068);
nor U6133 (N_6133,N_5907,N_5506);
nor U6134 (N_6134,N_5252,N_5791);
nor U6135 (N_6135,N_5325,N_5388);
nor U6136 (N_6136,N_5530,N_5420);
and U6137 (N_6137,N_5920,N_5793);
or U6138 (N_6138,N_5979,N_5271);
nor U6139 (N_6139,N_5772,N_5043);
nor U6140 (N_6140,N_5028,N_5386);
nor U6141 (N_6141,N_5556,N_5937);
nor U6142 (N_6142,N_5600,N_5894);
and U6143 (N_6143,N_5929,N_5469);
nand U6144 (N_6144,N_5673,N_5602);
and U6145 (N_6145,N_5472,N_5364);
and U6146 (N_6146,N_5475,N_5171);
nor U6147 (N_6147,N_5652,N_5074);
or U6148 (N_6148,N_5676,N_5953);
and U6149 (N_6149,N_5132,N_5084);
nor U6150 (N_6150,N_5055,N_5642);
xor U6151 (N_6151,N_5091,N_5211);
xor U6152 (N_6152,N_5590,N_5501);
or U6153 (N_6153,N_5478,N_5052);
nor U6154 (N_6154,N_5448,N_5674);
xnor U6155 (N_6155,N_5391,N_5899);
xnor U6156 (N_6156,N_5370,N_5210);
nor U6157 (N_6157,N_5567,N_5846);
nor U6158 (N_6158,N_5137,N_5935);
nor U6159 (N_6159,N_5644,N_5693);
xnor U6160 (N_6160,N_5594,N_5694);
nand U6161 (N_6161,N_5751,N_5718);
nand U6162 (N_6162,N_5349,N_5288);
or U6163 (N_6163,N_5225,N_5552);
or U6164 (N_6164,N_5417,N_5265);
or U6165 (N_6165,N_5422,N_5266);
and U6166 (N_6166,N_5064,N_5241);
and U6167 (N_6167,N_5721,N_5800);
or U6168 (N_6168,N_5072,N_5108);
xor U6169 (N_6169,N_5557,N_5066);
xor U6170 (N_6170,N_5572,N_5728);
and U6171 (N_6171,N_5057,N_5229);
xnor U6172 (N_6172,N_5313,N_5430);
or U6173 (N_6173,N_5175,N_5585);
nand U6174 (N_6174,N_5934,N_5309);
nor U6175 (N_6175,N_5938,N_5554);
xnor U6176 (N_6176,N_5488,N_5337);
or U6177 (N_6177,N_5696,N_5490);
nand U6178 (N_6178,N_5773,N_5394);
xnor U6179 (N_6179,N_5700,N_5691);
nand U6180 (N_6180,N_5320,N_5833);
and U6181 (N_6181,N_5803,N_5268);
nand U6182 (N_6182,N_5339,N_5398);
nor U6183 (N_6183,N_5976,N_5112);
and U6184 (N_6184,N_5082,N_5081);
or U6185 (N_6185,N_5258,N_5413);
xnor U6186 (N_6186,N_5311,N_5675);
nand U6187 (N_6187,N_5713,N_5822);
nand U6188 (N_6188,N_5071,N_5547);
and U6189 (N_6189,N_5885,N_5434);
nand U6190 (N_6190,N_5405,N_5477);
xnor U6191 (N_6191,N_5300,N_5952);
or U6192 (N_6192,N_5839,N_5307);
and U6193 (N_6193,N_5415,N_5664);
nand U6194 (N_6194,N_5841,N_5879);
or U6195 (N_6195,N_5684,N_5001);
nor U6196 (N_6196,N_5449,N_5924);
xor U6197 (N_6197,N_5034,N_5032);
nor U6198 (N_6198,N_5455,N_5251);
and U6199 (N_6199,N_5519,N_5984);
nand U6200 (N_6200,N_5658,N_5626);
or U6201 (N_6201,N_5106,N_5489);
xnor U6202 (N_6202,N_5466,N_5166);
nor U6203 (N_6203,N_5548,N_5965);
nor U6204 (N_6204,N_5631,N_5510);
or U6205 (N_6205,N_5147,N_5825);
nor U6206 (N_6206,N_5333,N_5592);
or U6207 (N_6207,N_5521,N_5807);
nor U6208 (N_6208,N_5549,N_5897);
nand U6209 (N_6209,N_5970,N_5445);
nand U6210 (N_6210,N_5319,N_5584);
nand U6211 (N_6211,N_5966,N_5184);
or U6212 (N_6212,N_5264,N_5461);
nor U6213 (N_6213,N_5099,N_5550);
xor U6214 (N_6214,N_5427,N_5067);
nand U6215 (N_6215,N_5645,N_5670);
nand U6216 (N_6216,N_5919,N_5859);
nor U6217 (N_6217,N_5918,N_5044);
nand U6218 (N_6218,N_5140,N_5922);
and U6219 (N_6219,N_5453,N_5877);
xnor U6220 (N_6220,N_5587,N_5579);
nor U6221 (N_6221,N_5193,N_5954);
or U6222 (N_6222,N_5121,N_5331);
nand U6223 (N_6223,N_5838,N_5156);
xor U6224 (N_6224,N_5893,N_5408);
nor U6225 (N_6225,N_5353,N_5198);
nand U6226 (N_6226,N_5160,N_5761);
and U6227 (N_6227,N_5185,N_5373);
or U6228 (N_6228,N_5323,N_5737);
nand U6229 (N_6229,N_5376,N_5189);
nand U6230 (N_6230,N_5687,N_5080);
xor U6231 (N_6231,N_5526,N_5486);
and U6232 (N_6232,N_5654,N_5870);
nor U6233 (N_6233,N_5246,N_5588);
or U6234 (N_6234,N_5172,N_5622);
nor U6235 (N_6235,N_5891,N_5298);
xnor U6236 (N_6236,N_5880,N_5399);
nand U6237 (N_6237,N_5220,N_5118);
or U6238 (N_6238,N_5368,N_5834);
nand U6239 (N_6239,N_5003,N_5991);
xor U6240 (N_6240,N_5049,N_5050);
xor U6241 (N_6241,N_5436,N_5491);
xor U6242 (N_6242,N_5380,N_5577);
and U6243 (N_6243,N_5709,N_5511);
nor U6244 (N_6244,N_5753,N_5835);
nor U6245 (N_6245,N_5541,N_5716);
and U6246 (N_6246,N_5969,N_5215);
nor U6247 (N_6247,N_5895,N_5503);
nand U6248 (N_6248,N_5306,N_5722);
nor U6249 (N_6249,N_5624,N_5372);
xnor U6250 (N_6250,N_5757,N_5418);
nand U6251 (N_6251,N_5881,N_5873);
and U6252 (N_6252,N_5532,N_5142);
or U6253 (N_6253,N_5591,N_5423);
or U6254 (N_6254,N_5254,N_5401);
nor U6255 (N_6255,N_5842,N_5620);
nand U6256 (N_6256,N_5115,N_5195);
or U6257 (N_6257,N_5103,N_5811);
nor U6258 (N_6258,N_5779,N_5317);
nand U6259 (N_6259,N_5234,N_5680);
nor U6260 (N_6260,N_5085,N_5174);
and U6261 (N_6261,N_5468,N_5165);
and U6262 (N_6262,N_5126,N_5708);
nand U6263 (N_6263,N_5355,N_5484);
and U6264 (N_6264,N_5109,N_5524);
nor U6265 (N_6265,N_5758,N_5961);
or U6266 (N_6266,N_5715,N_5663);
or U6267 (N_6267,N_5216,N_5357);
and U6268 (N_6268,N_5988,N_5994);
nor U6269 (N_6269,N_5683,N_5218);
nand U6270 (N_6270,N_5792,N_5507);
and U6271 (N_6271,N_5871,N_5456);
xnor U6272 (N_6272,N_5830,N_5205);
and U6273 (N_6273,N_5805,N_5124);
nand U6274 (N_6274,N_5798,N_5151);
xor U6275 (N_6275,N_5492,N_5347);
xnor U6276 (N_6276,N_5235,N_5270);
and U6277 (N_6277,N_5007,N_5949);
or U6278 (N_6278,N_5710,N_5543);
nand U6279 (N_6279,N_5321,N_5932);
nand U6280 (N_6280,N_5914,N_5096);
nand U6281 (N_6281,N_5735,N_5677);
xnor U6282 (N_6282,N_5778,N_5717);
nand U6283 (N_6283,N_5665,N_5204);
xor U6284 (N_6284,N_5520,N_5702);
or U6285 (N_6285,N_5076,N_5844);
nor U6286 (N_6286,N_5326,N_5884);
nand U6287 (N_6287,N_5384,N_5178);
xor U6288 (N_6288,N_5361,N_5719);
xor U6289 (N_6289,N_5123,N_5968);
xor U6290 (N_6290,N_5648,N_5425);
xor U6291 (N_6291,N_5077,N_5806);
nand U6292 (N_6292,N_5228,N_5569);
or U6293 (N_6293,N_5565,N_5872);
nor U6294 (N_6294,N_5041,N_5161);
and U6295 (N_6295,N_5618,N_5983);
or U6296 (N_6296,N_5975,N_5633);
xor U6297 (N_6297,N_5435,N_5273);
and U6298 (N_6298,N_5141,N_5765);
nor U6299 (N_6299,N_5869,N_5177);
and U6300 (N_6300,N_5782,N_5640);
or U6301 (N_6301,N_5164,N_5020);
nor U6302 (N_6302,N_5045,N_5818);
nor U6303 (N_6303,N_5375,N_5056);
and U6304 (N_6304,N_5623,N_5921);
nor U6305 (N_6305,N_5493,N_5303);
nand U6306 (N_6306,N_5996,N_5392);
and U6307 (N_6307,N_5827,N_5777);
and U6308 (N_6308,N_5051,N_5615);
nand U6309 (N_6309,N_5748,N_5720);
nor U6310 (N_6310,N_5038,N_5900);
xor U6311 (N_6311,N_5666,N_5754);
and U6312 (N_6312,N_5402,N_5986);
and U6313 (N_6313,N_5135,N_5947);
and U6314 (N_6314,N_5678,N_5878);
and U6315 (N_6315,N_5011,N_5729);
or U6316 (N_6316,N_5101,N_5540);
or U6317 (N_6317,N_5730,N_5231);
xor U6318 (N_6318,N_5181,N_5604);
nand U6319 (N_6319,N_5711,N_5908);
or U6320 (N_6320,N_5621,N_5851);
and U6321 (N_6321,N_5157,N_5180);
nor U6322 (N_6322,N_5381,N_5387);
xor U6323 (N_6323,N_5458,N_5653);
or U6324 (N_6324,N_5269,N_5245);
xor U6325 (N_6325,N_5025,N_5295);
nand U6326 (N_6326,N_5531,N_5039);
xor U6327 (N_6327,N_5898,N_5352);
xor U6328 (N_6328,N_5581,N_5379);
or U6329 (N_6329,N_5095,N_5518);
and U6330 (N_6330,N_5882,N_5464);
nand U6331 (N_6331,N_5366,N_5611);
and U6332 (N_6332,N_5145,N_5741);
and U6333 (N_6333,N_5528,N_5911);
or U6334 (N_6334,N_5747,N_5558);
or U6335 (N_6335,N_5759,N_5875);
nand U6336 (N_6336,N_5727,N_5515);
nor U6337 (N_6337,N_5610,N_5864);
or U6338 (N_6338,N_5315,N_5452);
nor U6339 (N_6339,N_5546,N_5732);
or U6340 (N_6340,N_5078,N_5606);
or U6341 (N_6341,N_5997,N_5239);
or U6342 (N_6342,N_5424,N_5393);
and U6343 (N_6343,N_5505,N_5201);
or U6344 (N_6344,N_5809,N_5973);
nand U6345 (N_6345,N_5824,N_5314);
and U6346 (N_6346,N_5113,N_5974);
xnor U6347 (N_6347,N_5212,N_5440);
xnor U6348 (N_6348,N_5457,N_5374);
nor U6349 (N_6349,N_5516,N_5942);
and U6350 (N_6350,N_5655,N_5247);
xnor U6351 (N_6351,N_5437,N_5930);
nand U6352 (N_6352,N_5293,N_5155);
and U6353 (N_6353,N_5672,N_5356);
nor U6354 (N_6354,N_5958,N_5249);
and U6355 (N_6355,N_5781,N_5560);
nand U6356 (N_6356,N_5289,N_5502);
and U6357 (N_6357,N_5742,N_5551);
and U6358 (N_6358,N_5382,N_5474);
and U6359 (N_6359,N_5593,N_5927);
nand U6360 (N_6360,N_5233,N_5775);
and U6361 (N_6361,N_5928,N_5866);
and U6362 (N_6362,N_5261,N_5397);
and U6363 (N_6363,N_5278,N_5931);
nor U6364 (N_6364,N_5788,N_5978);
nand U6365 (N_6365,N_5553,N_5483);
and U6366 (N_6366,N_5817,N_5495);
xor U6367 (N_6367,N_5097,N_5616);
and U6368 (N_6368,N_5910,N_5854);
nor U6369 (N_6369,N_5330,N_5150);
or U6370 (N_6370,N_5407,N_5203);
nand U6371 (N_6371,N_5143,N_5826);
or U6372 (N_6372,N_5454,N_5614);
or U6373 (N_6373,N_5061,N_5596);
nor U6374 (N_6374,N_5335,N_5745);
nand U6375 (N_6375,N_5750,N_5744);
nand U6376 (N_6376,N_5760,N_5535);
nand U6377 (N_6377,N_5787,N_5286);
nand U6378 (N_6378,N_5410,N_5989);
xor U6379 (N_6379,N_5460,N_5117);
or U6380 (N_6380,N_5669,N_5904);
xor U6381 (N_6381,N_5925,N_5186);
and U6382 (N_6382,N_5110,N_5130);
xor U6383 (N_6383,N_5053,N_5795);
nor U6384 (N_6384,N_5712,N_5714);
and U6385 (N_6385,N_5154,N_5086);
nor U6386 (N_6386,N_5896,N_5190);
xnor U6387 (N_6387,N_5482,N_5936);
or U6388 (N_6388,N_5451,N_5208);
or U6389 (N_6389,N_5962,N_5487);
and U6390 (N_6390,N_5206,N_5060);
or U6391 (N_6391,N_5194,N_5058);
xor U6392 (N_6392,N_5613,N_5033);
and U6393 (N_6393,N_5699,N_5956);
and U6394 (N_6394,N_5443,N_5221);
or U6395 (N_6395,N_5964,N_5079);
xnor U6396 (N_6396,N_5426,N_5429);
nand U6397 (N_6397,N_5992,N_5810);
or U6398 (N_6398,N_5823,N_5847);
nand U6399 (N_6399,N_5390,N_5701);
or U6400 (N_6400,N_5656,N_5849);
nor U6401 (N_6401,N_5734,N_5284);
nand U6402 (N_6402,N_5187,N_5828);
nor U6403 (N_6403,N_5582,N_5509);
nand U6404 (N_6404,N_5783,N_5850);
nor U6405 (N_6405,N_5015,N_5297);
or U6406 (N_6406,N_5861,N_5705);
nand U6407 (N_6407,N_5018,N_5836);
and U6408 (N_6408,N_5419,N_5815);
nor U6409 (N_6409,N_5308,N_5087);
nand U6410 (N_6410,N_5689,N_5862);
nor U6411 (N_6411,N_5804,N_5629);
or U6412 (N_6412,N_5829,N_5865);
xor U6413 (N_6413,N_5889,N_5733);
nor U6414 (N_6414,N_5122,N_5217);
and U6415 (N_6415,N_5863,N_5950);
nand U6416 (N_6416,N_5336,N_5960);
and U6417 (N_6417,N_5365,N_5473);
or U6418 (N_6418,N_5111,N_5090);
nor U6419 (N_6419,N_5703,N_5463);
and U6420 (N_6420,N_5948,N_5957);
or U6421 (N_6421,N_5351,N_5296);
and U6422 (N_6422,N_5054,N_5294);
xnor U6423 (N_6423,N_5237,N_5943);
xnor U6424 (N_6424,N_5905,N_5738);
xor U6425 (N_6425,N_5471,N_5360);
nor U6426 (N_6426,N_5764,N_5149);
nand U6427 (N_6427,N_5813,N_5802);
nand U6428 (N_6428,N_5945,N_5499);
nor U6429 (N_6429,N_5568,N_5116);
or U6430 (N_6430,N_5403,N_5279);
or U6431 (N_6431,N_5855,N_5972);
nand U6432 (N_6432,N_5447,N_5299);
nor U6433 (N_6433,N_5812,N_5784);
and U6434 (N_6434,N_5853,N_5219);
nand U6435 (N_6435,N_5628,N_5662);
nand U6436 (N_6436,N_5318,N_5343);
nand U6437 (N_6437,N_5601,N_5253);
nor U6438 (N_6438,N_5564,N_5496);
nand U6439 (N_6439,N_5522,N_5545);
and U6440 (N_6440,N_5599,N_5959);
nand U6441 (N_6441,N_5168,N_5004);
xor U6442 (N_6442,N_5467,N_5939);
or U6443 (N_6443,N_5575,N_5686);
nor U6444 (N_6444,N_5342,N_5396);
or U6445 (N_6445,N_5378,N_5913);
xnor U6446 (N_6446,N_5275,N_5612);
or U6447 (N_6447,N_5138,N_5006);
nand U6448 (N_6448,N_5527,N_5450);
nor U6449 (N_6449,N_5589,N_5200);
nor U6450 (N_6450,N_5909,N_5660);
nand U6451 (N_6451,N_5995,N_5421);
or U6452 (N_6452,N_5595,N_5946);
and U6453 (N_6453,N_5021,N_5262);
nor U6454 (N_6454,N_5442,N_5688);
and U6455 (N_6455,N_5874,N_5999);
or U6456 (N_6456,N_5158,N_5570);
xor U6457 (N_6457,N_5766,N_5555);
or U6458 (N_6458,N_5739,N_5852);
or U6459 (N_6459,N_5704,N_5327);
nor U6460 (N_6460,N_5432,N_5731);
or U6461 (N_6461,N_5348,N_5083);
nor U6462 (N_6462,N_5305,N_5819);
xnor U6463 (N_6463,N_5263,N_5202);
nor U6464 (N_6464,N_5536,N_5647);
nor U6465 (N_6465,N_5098,N_5019);
nand U6466 (N_6466,N_5915,N_5431);
nand U6467 (N_6467,N_5438,N_5523);
and U6468 (N_6468,N_5302,N_5100);
xnor U6469 (N_6469,N_5867,N_5179);
or U6470 (N_6470,N_5769,N_5062);
or U6471 (N_6471,N_5726,N_5840);
and U6472 (N_6472,N_5630,N_5441);
or U6473 (N_6473,N_5776,N_5243);
nand U6474 (N_6474,N_5821,N_5597);
nor U6475 (N_6475,N_5649,N_5197);
or U6476 (N_6476,N_5749,N_5341);
xor U6477 (N_6477,N_5799,N_5608);
nor U6478 (N_6478,N_5292,N_5480);
nor U6479 (N_6479,N_5513,N_5024);
or U6480 (N_6480,N_5941,N_5514);
xor U6481 (N_6481,N_5485,N_5227);
nand U6482 (N_6482,N_5638,N_5890);
xor U6483 (N_6483,N_5102,N_5650);
or U6484 (N_6484,N_5494,N_5657);
and U6485 (N_6485,N_5073,N_5459);
or U6486 (N_6486,N_5542,N_5244);
or U6487 (N_6487,N_5036,N_5661);
nand U6488 (N_6488,N_5685,N_5641);
or U6489 (N_6489,N_5617,N_5240);
or U6490 (N_6490,N_5167,N_5923);
xnor U6491 (N_6491,N_5192,N_5790);
or U6492 (N_6492,N_5277,N_5146);
and U6493 (N_6493,N_5094,N_5627);
xnor U6494 (N_6494,N_5222,N_5411);
nor U6495 (N_6495,N_5027,N_5762);
nand U6496 (N_6496,N_5695,N_5362);
and U6497 (N_6497,N_5797,N_5047);
xnor U6498 (N_6498,N_5888,N_5539);
nor U6499 (N_6499,N_5963,N_5280);
and U6500 (N_6500,N_5500,N_5141);
xor U6501 (N_6501,N_5892,N_5075);
or U6502 (N_6502,N_5753,N_5065);
nor U6503 (N_6503,N_5898,N_5845);
and U6504 (N_6504,N_5343,N_5408);
and U6505 (N_6505,N_5415,N_5794);
xnor U6506 (N_6506,N_5166,N_5468);
nor U6507 (N_6507,N_5921,N_5685);
or U6508 (N_6508,N_5875,N_5823);
or U6509 (N_6509,N_5583,N_5999);
nand U6510 (N_6510,N_5889,N_5204);
nand U6511 (N_6511,N_5804,N_5352);
nand U6512 (N_6512,N_5798,N_5076);
and U6513 (N_6513,N_5401,N_5592);
and U6514 (N_6514,N_5546,N_5171);
and U6515 (N_6515,N_5144,N_5751);
xnor U6516 (N_6516,N_5881,N_5070);
nand U6517 (N_6517,N_5810,N_5020);
nand U6518 (N_6518,N_5903,N_5441);
xor U6519 (N_6519,N_5977,N_5374);
nand U6520 (N_6520,N_5678,N_5478);
nand U6521 (N_6521,N_5597,N_5204);
nor U6522 (N_6522,N_5038,N_5617);
nor U6523 (N_6523,N_5130,N_5834);
nor U6524 (N_6524,N_5600,N_5941);
nand U6525 (N_6525,N_5826,N_5763);
nand U6526 (N_6526,N_5569,N_5604);
nand U6527 (N_6527,N_5483,N_5501);
or U6528 (N_6528,N_5369,N_5351);
and U6529 (N_6529,N_5581,N_5322);
and U6530 (N_6530,N_5941,N_5854);
nor U6531 (N_6531,N_5029,N_5042);
nand U6532 (N_6532,N_5081,N_5047);
nor U6533 (N_6533,N_5777,N_5685);
or U6534 (N_6534,N_5748,N_5571);
or U6535 (N_6535,N_5623,N_5809);
xnor U6536 (N_6536,N_5225,N_5609);
nor U6537 (N_6537,N_5764,N_5766);
or U6538 (N_6538,N_5254,N_5614);
xnor U6539 (N_6539,N_5863,N_5935);
xnor U6540 (N_6540,N_5785,N_5739);
and U6541 (N_6541,N_5336,N_5046);
or U6542 (N_6542,N_5149,N_5041);
and U6543 (N_6543,N_5558,N_5305);
and U6544 (N_6544,N_5303,N_5702);
and U6545 (N_6545,N_5544,N_5069);
or U6546 (N_6546,N_5192,N_5160);
and U6547 (N_6547,N_5383,N_5036);
or U6548 (N_6548,N_5537,N_5960);
and U6549 (N_6549,N_5932,N_5637);
or U6550 (N_6550,N_5425,N_5226);
xor U6551 (N_6551,N_5595,N_5646);
or U6552 (N_6552,N_5117,N_5262);
and U6553 (N_6553,N_5753,N_5781);
xnor U6554 (N_6554,N_5277,N_5301);
xnor U6555 (N_6555,N_5126,N_5792);
or U6556 (N_6556,N_5614,N_5858);
nor U6557 (N_6557,N_5034,N_5208);
nor U6558 (N_6558,N_5111,N_5624);
nor U6559 (N_6559,N_5996,N_5083);
nor U6560 (N_6560,N_5283,N_5307);
nand U6561 (N_6561,N_5858,N_5517);
and U6562 (N_6562,N_5022,N_5424);
nor U6563 (N_6563,N_5508,N_5054);
or U6564 (N_6564,N_5339,N_5026);
xnor U6565 (N_6565,N_5257,N_5200);
nand U6566 (N_6566,N_5225,N_5126);
xor U6567 (N_6567,N_5607,N_5511);
nand U6568 (N_6568,N_5985,N_5560);
nand U6569 (N_6569,N_5348,N_5855);
and U6570 (N_6570,N_5730,N_5888);
xor U6571 (N_6571,N_5226,N_5557);
and U6572 (N_6572,N_5753,N_5962);
or U6573 (N_6573,N_5210,N_5533);
nor U6574 (N_6574,N_5874,N_5691);
nand U6575 (N_6575,N_5738,N_5476);
nand U6576 (N_6576,N_5546,N_5525);
nand U6577 (N_6577,N_5924,N_5017);
and U6578 (N_6578,N_5718,N_5895);
and U6579 (N_6579,N_5433,N_5641);
or U6580 (N_6580,N_5828,N_5722);
xor U6581 (N_6581,N_5145,N_5989);
nor U6582 (N_6582,N_5926,N_5850);
and U6583 (N_6583,N_5318,N_5392);
nor U6584 (N_6584,N_5073,N_5984);
nand U6585 (N_6585,N_5724,N_5444);
and U6586 (N_6586,N_5296,N_5273);
xnor U6587 (N_6587,N_5575,N_5598);
and U6588 (N_6588,N_5266,N_5512);
nor U6589 (N_6589,N_5797,N_5407);
and U6590 (N_6590,N_5342,N_5464);
xor U6591 (N_6591,N_5629,N_5251);
and U6592 (N_6592,N_5472,N_5702);
or U6593 (N_6593,N_5600,N_5197);
and U6594 (N_6594,N_5346,N_5426);
or U6595 (N_6595,N_5292,N_5279);
or U6596 (N_6596,N_5796,N_5789);
and U6597 (N_6597,N_5892,N_5050);
or U6598 (N_6598,N_5681,N_5878);
nor U6599 (N_6599,N_5694,N_5440);
and U6600 (N_6600,N_5406,N_5883);
xnor U6601 (N_6601,N_5972,N_5552);
or U6602 (N_6602,N_5987,N_5488);
and U6603 (N_6603,N_5820,N_5932);
nor U6604 (N_6604,N_5659,N_5040);
xnor U6605 (N_6605,N_5769,N_5595);
nand U6606 (N_6606,N_5436,N_5959);
xor U6607 (N_6607,N_5964,N_5183);
or U6608 (N_6608,N_5208,N_5146);
nand U6609 (N_6609,N_5576,N_5898);
and U6610 (N_6610,N_5532,N_5561);
or U6611 (N_6611,N_5324,N_5249);
nor U6612 (N_6612,N_5051,N_5699);
nand U6613 (N_6613,N_5260,N_5712);
or U6614 (N_6614,N_5450,N_5303);
nand U6615 (N_6615,N_5266,N_5670);
xnor U6616 (N_6616,N_5455,N_5022);
xor U6617 (N_6617,N_5398,N_5760);
nand U6618 (N_6618,N_5717,N_5081);
xnor U6619 (N_6619,N_5946,N_5147);
nor U6620 (N_6620,N_5183,N_5442);
nor U6621 (N_6621,N_5202,N_5405);
and U6622 (N_6622,N_5267,N_5257);
or U6623 (N_6623,N_5105,N_5030);
and U6624 (N_6624,N_5224,N_5003);
xnor U6625 (N_6625,N_5822,N_5378);
and U6626 (N_6626,N_5568,N_5859);
nor U6627 (N_6627,N_5670,N_5601);
and U6628 (N_6628,N_5507,N_5081);
and U6629 (N_6629,N_5432,N_5416);
and U6630 (N_6630,N_5564,N_5148);
or U6631 (N_6631,N_5506,N_5251);
nor U6632 (N_6632,N_5729,N_5405);
nand U6633 (N_6633,N_5669,N_5464);
xor U6634 (N_6634,N_5931,N_5894);
nor U6635 (N_6635,N_5746,N_5729);
nand U6636 (N_6636,N_5020,N_5402);
or U6637 (N_6637,N_5884,N_5069);
and U6638 (N_6638,N_5874,N_5510);
or U6639 (N_6639,N_5505,N_5876);
or U6640 (N_6640,N_5935,N_5724);
nor U6641 (N_6641,N_5275,N_5880);
xnor U6642 (N_6642,N_5123,N_5380);
or U6643 (N_6643,N_5271,N_5386);
xnor U6644 (N_6644,N_5400,N_5246);
nor U6645 (N_6645,N_5841,N_5837);
xor U6646 (N_6646,N_5292,N_5159);
xor U6647 (N_6647,N_5252,N_5165);
nand U6648 (N_6648,N_5703,N_5924);
xor U6649 (N_6649,N_5112,N_5859);
nor U6650 (N_6650,N_5059,N_5134);
or U6651 (N_6651,N_5438,N_5684);
or U6652 (N_6652,N_5605,N_5685);
or U6653 (N_6653,N_5569,N_5978);
xor U6654 (N_6654,N_5144,N_5599);
nor U6655 (N_6655,N_5189,N_5734);
xnor U6656 (N_6656,N_5202,N_5501);
nand U6657 (N_6657,N_5152,N_5483);
xor U6658 (N_6658,N_5298,N_5633);
xor U6659 (N_6659,N_5756,N_5384);
and U6660 (N_6660,N_5482,N_5345);
xnor U6661 (N_6661,N_5424,N_5229);
or U6662 (N_6662,N_5821,N_5433);
and U6663 (N_6663,N_5160,N_5584);
or U6664 (N_6664,N_5562,N_5666);
and U6665 (N_6665,N_5141,N_5017);
or U6666 (N_6666,N_5920,N_5908);
nor U6667 (N_6667,N_5811,N_5633);
and U6668 (N_6668,N_5794,N_5685);
nor U6669 (N_6669,N_5598,N_5732);
or U6670 (N_6670,N_5801,N_5563);
nor U6671 (N_6671,N_5392,N_5416);
or U6672 (N_6672,N_5628,N_5965);
xnor U6673 (N_6673,N_5044,N_5375);
nor U6674 (N_6674,N_5891,N_5323);
and U6675 (N_6675,N_5350,N_5198);
or U6676 (N_6676,N_5460,N_5277);
and U6677 (N_6677,N_5758,N_5476);
xnor U6678 (N_6678,N_5459,N_5089);
nand U6679 (N_6679,N_5030,N_5354);
or U6680 (N_6680,N_5335,N_5574);
or U6681 (N_6681,N_5152,N_5175);
nor U6682 (N_6682,N_5370,N_5164);
xor U6683 (N_6683,N_5748,N_5524);
or U6684 (N_6684,N_5334,N_5457);
and U6685 (N_6685,N_5709,N_5875);
or U6686 (N_6686,N_5142,N_5266);
nand U6687 (N_6687,N_5727,N_5951);
xnor U6688 (N_6688,N_5445,N_5179);
or U6689 (N_6689,N_5138,N_5882);
nand U6690 (N_6690,N_5168,N_5950);
nor U6691 (N_6691,N_5738,N_5722);
nor U6692 (N_6692,N_5341,N_5512);
and U6693 (N_6693,N_5260,N_5210);
nor U6694 (N_6694,N_5584,N_5881);
or U6695 (N_6695,N_5681,N_5901);
nor U6696 (N_6696,N_5286,N_5935);
xnor U6697 (N_6697,N_5912,N_5481);
or U6698 (N_6698,N_5907,N_5964);
nand U6699 (N_6699,N_5257,N_5223);
xnor U6700 (N_6700,N_5192,N_5759);
nor U6701 (N_6701,N_5298,N_5833);
nor U6702 (N_6702,N_5471,N_5761);
and U6703 (N_6703,N_5939,N_5826);
and U6704 (N_6704,N_5494,N_5296);
nor U6705 (N_6705,N_5397,N_5679);
nor U6706 (N_6706,N_5927,N_5835);
xnor U6707 (N_6707,N_5789,N_5447);
and U6708 (N_6708,N_5183,N_5293);
xnor U6709 (N_6709,N_5126,N_5596);
and U6710 (N_6710,N_5607,N_5341);
nor U6711 (N_6711,N_5985,N_5635);
nor U6712 (N_6712,N_5887,N_5340);
or U6713 (N_6713,N_5062,N_5470);
or U6714 (N_6714,N_5733,N_5827);
nor U6715 (N_6715,N_5077,N_5102);
or U6716 (N_6716,N_5040,N_5004);
or U6717 (N_6717,N_5884,N_5965);
nand U6718 (N_6718,N_5083,N_5367);
nand U6719 (N_6719,N_5844,N_5896);
nand U6720 (N_6720,N_5693,N_5134);
nand U6721 (N_6721,N_5182,N_5585);
nand U6722 (N_6722,N_5030,N_5412);
xor U6723 (N_6723,N_5601,N_5047);
and U6724 (N_6724,N_5643,N_5542);
nand U6725 (N_6725,N_5894,N_5445);
and U6726 (N_6726,N_5823,N_5708);
nand U6727 (N_6727,N_5747,N_5975);
nand U6728 (N_6728,N_5195,N_5289);
and U6729 (N_6729,N_5235,N_5258);
and U6730 (N_6730,N_5457,N_5324);
nor U6731 (N_6731,N_5574,N_5003);
nand U6732 (N_6732,N_5917,N_5014);
nor U6733 (N_6733,N_5318,N_5448);
or U6734 (N_6734,N_5858,N_5338);
nor U6735 (N_6735,N_5184,N_5209);
or U6736 (N_6736,N_5115,N_5717);
or U6737 (N_6737,N_5708,N_5336);
or U6738 (N_6738,N_5293,N_5968);
and U6739 (N_6739,N_5002,N_5518);
nor U6740 (N_6740,N_5533,N_5708);
nor U6741 (N_6741,N_5981,N_5098);
or U6742 (N_6742,N_5143,N_5145);
nor U6743 (N_6743,N_5080,N_5312);
xor U6744 (N_6744,N_5249,N_5532);
or U6745 (N_6745,N_5471,N_5514);
nand U6746 (N_6746,N_5014,N_5209);
and U6747 (N_6747,N_5181,N_5257);
xnor U6748 (N_6748,N_5809,N_5441);
xnor U6749 (N_6749,N_5273,N_5451);
nand U6750 (N_6750,N_5425,N_5738);
or U6751 (N_6751,N_5271,N_5428);
or U6752 (N_6752,N_5700,N_5675);
and U6753 (N_6753,N_5898,N_5441);
and U6754 (N_6754,N_5536,N_5564);
nor U6755 (N_6755,N_5355,N_5740);
or U6756 (N_6756,N_5053,N_5412);
nor U6757 (N_6757,N_5936,N_5554);
xor U6758 (N_6758,N_5755,N_5875);
or U6759 (N_6759,N_5354,N_5310);
and U6760 (N_6760,N_5384,N_5793);
nor U6761 (N_6761,N_5569,N_5592);
nor U6762 (N_6762,N_5036,N_5589);
or U6763 (N_6763,N_5773,N_5988);
and U6764 (N_6764,N_5291,N_5367);
or U6765 (N_6765,N_5313,N_5261);
nor U6766 (N_6766,N_5848,N_5435);
or U6767 (N_6767,N_5210,N_5045);
nand U6768 (N_6768,N_5264,N_5870);
nor U6769 (N_6769,N_5722,N_5672);
nand U6770 (N_6770,N_5434,N_5408);
nor U6771 (N_6771,N_5708,N_5972);
nand U6772 (N_6772,N_5512,N_5656);
and U6773 (N_6773,N_5229,N_5253);
and U6774 (N_6774,N_5553,N_5929);
and U6775 (N_6775,N_5508,N_5826);
nor U6776 (N_6776,N_5161,N_5571);
xor U6777 (N_6777,N_5584,N_5070);
or U6778 (N_6778,N_5369,N_5790);
and U6779 (N_6779,N_5110,N_5568);
and U6780 (N_6780,N_5587,N_5470);
or U6781 (N_6781,N_5902,N_5696);
and U6782 (N_6782,N_5071,N_5767);
nor U6783 (N_6783,N_5930,N_5318);
xnor U6784 (N_6784,N_5915,N_5574);
nor U6785 (N_6785,N_5830,N_5554);
and U6786 (N_6786,N_5813,N_5631);
or U6787 (N_6787,N_5199,N_5843);
nor U6788 (N_6788,N_5779,N_5436);
nor U6789 (N_6789,N_5157,N_5248);
and U6790 (N_6790,N_5134,N_5071);
or U6791 (N_6791,N_5547,N_5426);
xnor U6792 (N_6792,N_5293,N_5022);
nand U6793 (N_6793,N_5656,N_5457);
xor U6794 (N_6794,N_5542,N_5944);
nand U6795 (N_6795,N_5216,N_5742);
or U6796 (N_6796,N_5856,N_5177);
nand U6797 (N_6797,N_5904,N_5404);
nor U6798 (N_6798,N_5615,N_5176);
xor U6799 (N_6799,N_5511,N_5739);
nor U6800 (N_6800,N_5266,N_5448);
nor U6801 (N_6801,N_5243,N_5001);
or U6802 (N_6802,N_5331,N_5066);
xnor U6803 (N_6803,N_5101,N_5445);
nor U6804 (N_6804,N_5777,N_5461);
and U6805 (N_6805,N_5491,N_5885);
nand U6806 (N_6806,N_5437,N_5531);
xor U6807 (N_6807,N_5995,N_5939);
xnor U6808 (N_6808,N_5956,N_5841);
and U6809 (N_6809,N_5727,N_5372);
xor U6810 (N_6810,N_5160,N_5754);
nor U6811 (N_6811,N_5678,N_5745);
nor U6812 (N_6812,N_5067,N_5931);
xor U6813 (N_6813,N_5671,N_5496);
nand U6814 (N_6814,N_5069,N_5109);
or U6815 (N_6815,N_5913,N_5674);
nor U6816 (N_6816,N_5638,N_5272);
xor U6817 (N_6817,N_5965,N_5243);
nand U6818 (N_6818,N_5851,N_5041);
nor U6819 (N_6819,N_5328,N_5368);
or U6820 (N_6820,N_5217,N_5923);
nand U6821 (N_6821,N_5658,N_5464);
nor U6822 (N_6822,N_5158,N_5849);
and U6823 (N_6823,N_5793,N_5894);
nor U6824 (N_6824,N_5435,N_5174);
and U6825 (N_6825,N_5280,N_5657);
xor U6826 (N_6826,N_5719,N_5935);
xnor U6827 (N_6827,N_5016,N_5749);
and U6828 (N_6828,N_5876,N_5818);
nand U6829 (N_6829,N_5771,N_5220);
nand U6830 (N_6830,N_5149,N_5417);
xor U6831 (N_6831,N_5404,N_5068);
nor U6832 (N_6832,N_5864,N_5224);
or U6833 (N_6833,N_5929,N_5614);
or U6834 (N_6834,N_5549,N_5712);
or U6835 (N_6835,N_5775,N_5366);
xor U6836 (N_6836,N_5297,N_5594);
nand U6837 (N_6837,N_5620,N_5087);
and U6838 (N_6838,N_5530,N_5846);
xor U6839 (N_6839,N_5727,N_5784);
or U6840 (N_6840,N_5015,N_5894);
and U6841 (N_6841,N_5127,N_5684);
or U6842 (N_6842,N_5685,N_5139);
and U6843 (N_6843,N_5657,N_5318);
nor U6844 (N_6844,N_5559,N_5126);
nor U6845 (N_6845,N_5651,N_5973);
xnor U6846 (N_6846,N_5989,N_5583);
nand U6847 (N_6847,N_5437,N_5714);
nand U6848 (N_6848,N_5966,N_5496);
nor U6849 (N_6849,N_5093,N_5279);
or U6850 (N_6850,N_5536,N_5334);
nor U6851 (N_6851,N_5426,N_5382);
and U6852 (N_6852,N_5117,N_5779);
nor U6853 (N_6853,N_5287,N_5255);
and U6854 (N_6854,N_5029,N_5720);
nor U6855 (N_6855,N_5271,N_5836);
or U6856 (N_6856,N_5547,N_5083);
nor U6857 (N_6857,N_5844,N_5861);
nor U6858 (N_6858,N_5624,N_5505);
xor U6859 (N_6859,N_5926,N_5352);
or U6860 (N_6860,N_5367,N_5177);
nand U6861 (N_6861,N_5205,N_5026);
and U6862 (N_6862,N_5021,N_5440);
xnor U6863 (N_6863,N_5044,N_5410);
nand U6864 (N_6864,N_5162,N_5598);
xnor U6865 (N_6865,N_5046,N_5715);
xor U6866 (N_6866,N_5112,N_5770);
xnor U6867 (N_6867,N_5414,N_5884);
or U6868 (N_6868,N_5168,N_5113);
nor U6869 (N_6869,N_5713,N_5203);
xnor U6870 (N_6870,N_5868,N_5786);
nor U6871 (N_6871,N_5882,N_5166);
nand U6872 (N_6872,N_5840,N_5086);
xor U6873 (N_6873,N_5482,N_5323);
and U6874 (N_6874,N_5429,N_5538);
and U6875 (N_6875,N_5497,N_5286);
and U6876 (N_6876,N_5636,N_5729);
nor U6877 (N_6877,N_5089,N_5099);
or U6878 (N_6878,N_5862,N_5109);
nand U6879 (N_6879,N_5286,N_5192);
nand U6880 (N_6880,N_5027,N_5817);
nand U6881 (N_6881,N_5666,N_5037);
xor U6882 (N_6882,N_5071,N_5738);
or U6883 (N_6883,N_5838,N_5360);
xor U6884 (N_6884,N_5440,N_5831);
nor U6885 (N_6885,N_5727,N_5232);
xnor U6886 (N_6886,N_5208,N_5340);
nor U6887 (N_6887,N_5046,N_5309);
nor U6888 (N_6888,N_5941,N_5623);
or U6889 (N_6889,N_5491,N_5187);
and U6890 (N_6890,N_5949,N_5425);
xor U6891 (N_6891,N_5248,N_5703);
xnor U6892 (N_6892,N_5433,N_5567);
or U6893 (N_6893,N_5934,N_5949);
and U6894 (N_6894,N_5485,N_5679);
and U6895 (N_6895,N_5269,N_5181);
xnor U6896 (N_6896,N_5932,N_5152);
nor U6897 (N_6897,N_5985,N_5394);
or U6898 (N_6898,N_5016,N_5702);
xor U6899 (N_6899,N_5120,N_5637);
nand U6900 (N_6900,N_5292,N_5276);
or U6901 (N_6901,N_5962,N_5648);
xnor U6902 (N_6902,N_5120,N_5866);
and U6903 (N_6903,N_5438,N_5685);
nand U6904 (N_6904,N_5134,N_5824);
nand U6905 (N_6905,N_5629,N_5118);
nand U6906 (N_6906,N_5261,N_5705);
xnor U6907 (N_6907,N_5201,N_5159);
xor U6908 (N_6908,N_5535,N_5512);
xnor U6909 (N_6909,N_5699,N_5098);
nand U6910 (N_6910,N_5047,N_5065);
and U6911 (N_6911,N_5829,N_5423);
and U6912 (N_6912,N_5628,N_5102);
or U6913 (N_6913,N_5223,N_5464);
and U6914 (N_6914,N_5691,N_5249);
xor U6915 (N_6915,N_5005,N_5335);
xor U6916 (N_6916,N_5951,N_5095);
nand U6917 (N_6917,N_5350,N_5196);
xnor U6918 (N_6918,N_5474,N_5255);
and U6919 (N_6919,N_5775,N_5738);
xor U6920 (N_6920,N_5062,N_5228);
xor U6921 (N_6921,N_5639,N_5834);
nand U6922 (N_6922,N_5992,N_5038);
xor U6923 (N_6923,N_5557,N_5105);
xnor U6924 (N_6924,N_5742,N_5186);
nand U6925 (N_6925,N_5268,N_5718);
and U6926 (N_6926,N_5623,N_5953);
nor U6927 (N_6927,N_5967,N_5628);
nor U6928 (N_6928,N_5659,N_5632);
nand U6929 (N_6929,N_5160,N_5910);
nor U6930 (N_6930,N_5476,N_5306);
and U6931 (N_6931,N_5530,N_5023);
xor U6932 (N_6932,N_5886,N_5359);
nand U6933 (N_6933,N_5688,N_5831);
nand U6934 (N_6934,N_5443,N_5708);
xor U6935 (N_6935,N_5585,N_5561);
or U6936 (N_6936,N_5047,N_5094);
or U6937 (N_6937,N_5019,N_5476);
nand U6938 (N_6938,N_5957,N_5065);
and U6939 (N_6939,N_5183,N_5310);
or U6940 (N_6940,N_5118,N_5913);
nand U6941 (N_6941,N_5677,N_5878);
xnor U6942 (N_6942,N_5471,N_5809);
or U6943 (N_6943,N_5828,N_5780);
nor U6944 (N_6944,N_5117,N_5038);
or U6945 (N_6945,N_5620,N_5584);
nand U6946 (N_6946,N_5353,N_5701);
nor U6947 (N_6947,N_5281,N_5888);
or U6948 (N_6948,N_5661,N_5944);
xnor U6949 (N_6949,N_5904,N_5205);
xor U6950 (N_6950,N_5834,N_5257);
or U6951 (N_6951,N_5736,N_5144);
and U6952 (N_6952,N_5587,N_5412);
or U6953 (N_6953,N_5868,N_5962);
nand U6954 (N_6954,N_5473,N_5894);
xor U6955 (N_6955,N_5634,N_5263);
or U6956 (N_6956,N_5210,N_5568);
nor U6957 (N_6957,N_5937,N_5065);
xor U6958 (N_6958,N_5558,N_5088);
xnor U6959 (N_6959,N_5371,N_5136);
xnor U6960 (N_6960,N_5369,N_5514);
and U6961 (N_6961,N_5249,N_5948);
and U6962 (N_6962,N_5386,N_5759);
xnor U6963 (N_6963,N_5054,N_5705);
nand U6964 (N_6964,N_5754,N_5114);
or U6965 (N_6965,N_5670,N_5328);
or U6966 (N_6966,N_5994,N_5268);
nand U6967 (N_6967,N_5832,N_5627);
xor U6968 (N_6968,N_5265,N_5635);
or U6969 (N_6969,N_5949,N_5174);
and U6970 (N_6970,N_5127,N_5237);
nand U6971 (N_6971,N_5908,N_5289);
and U6972 (N_6972,N_5344,N_5411);
nand U6973 (N_6973,N_5868,N_5828);
nor U6974 (N_6974,N_5693,N_5968);
and U6975 (N_6975,N_5419,N_5987);
xor U6976 (N_6976,N_5763,N_5036);
nand U6977 (N_6977,N_5441,N_5553);
nand U6978 (N_6978,N_5917,N_5452);
or U6979 (N_6979,N_5455,N_5282);
nand U6980 (N_6980,N_5453,N_5240);
and U6981 (N_6981,N_5257,N_5105);
and U6982 (N_6982,N_5949,N_5407);
nand U6983 (N_6983,N_5210,N_5821);
and U6984 (N_6984,N_5878,N_5134);
xor U6985 (N_6985,N_5836,N_5924);
or U6986 (N_6986,N_5974,N_5996);
or U6987 (N_6987,N_5662,N_5241);
nand U6988 (N_6988,N_5374,N_5674);
nand U6989 (N_6989,N_5173,N_5761);
nor U6990 (N_6990,N_5434,N_5600);
and U6991 (N_6991,N_5969,N_5822);
nor U6992 (N_6992,N_5519,N_5048);
nor U6993 (N_6993,N_5755,N_5029);
xor U6994 (N_6994,N_5058,N_5628);
nand U6995 (N_6995,N_5357,N_5190);
xor U6996 (N_6996,N_5398,N_5311);
and U6997 (N_6997,N_5244,N_5829);
xor U6998 (N_6998,N_5917,N_5428);
and U6999 (N_6999,N_5518,N_5483);
nand U7000 (N_7000,N_6210,N_6713);
or U7001 (N_7001,N_6201,N_6569);
xor U7002 (N_7002,N_6370,N_6507);
or U7003 (N_7003,N_6738,N_6620);
and U7004 (N_7004,N_6492,N_6957);
or U7005 (N_7005,N_6949,N_6032);
nor U7006 (N_7006,N_6482,N_6230);
or U7007 (N_7007,N_6955,N_6020);
nor U7008 (N_7008,N_6191,N_6319);
nor U7009 (N_7009,N_6596,N_6764);
xnor U7010 (N_7010,N_6410,N_6233);
xnor U7011 (N_7011,N_6740,N_6071);
nand U7012 (N_7012,N_6404,N_6649);
nor U7013 (N_7013,N_6617,N_6480);
or U7014 (N_7014,N_6090,N_6054);
and U7015 (N_7015,N_6003,N_6986);
nor U7016 (N_7016,N_6060,N_6842);
nand U7017 (N_7017,N_6262,N_6558);
xor U7018 (N_7018,N_6089,N_6792);
xnor U7019 (N_7019,N_6638,N_6282);
nand U7020 (N_7020,N_6857,N_6280);
nand U7021 (N_7021,N_6696,N_6712);
xor U7022 (N_7022,N_6013,N_6775);
nand U7023 (N_7023,N_6968,N_6747);
or U7024 (N_7024,N_6145,N_6268);
nand U7025 (N_7025,N_6070,N_6913);
nor U7026 (N_7026,N_6841,N_6814);
nor U7027 (N_7027,N_6359,N_6822);
and U7028 (N_7028,N_6880,N_6152);
xor U7029 (N_7029,N_6905,N_6754);
xor U7030 (N_7030,N_6081,N_6932);
and U7031 (N_7031,N_6242,N_6209);
xor U7032 (N_7032,N_6402,N_6748);
and U7033 (N_7033,N_6112,N_6515);
nand U7034 (N_7034,N_6072,N_6142);
xor U7035 (N_7035,N_6449,N_6944);
nand U7036 (N_7036,N_6799,N_6030);
and U7037 (N_7037,N_6690,N_6954);
and U7038 (N_7038,N_6141,N_6065);
nor U7039 (N_7039,N_6837,N_6861);
xnor U7040 (N_7040,N_6196,N_6371);
and U7041 (N_7041,N_6976,N_6945);
xnor U7042 (N_7042,N_6600,N_6828);
nand U7043 (N_7043,N_6715,N_6753);
nand U7044 (N_7044,N_6687,N_6639);
and U7045 (N_7045,N_6217,N_6534);
or U7046 (N_7046,N_6397,N_6719);
nand U7047 (N_7047,N_6961,N_6232);
or U7048 (N_7048,N_6756,N_6667);
nor U7049 (N_7049,N_6500,N_6363);
nor U7050 (N_7050,N_6585,N_6956);
or U7051 (N_7051,N_6646,N_6336);
or U7052 (N_7052,N_6644,N_6931);
nand U7053 (N_7053,N_6628,N_6110);
or U7054 (N_7054,N_6185,N_6975);
and U7055 (N_7055,N_6391,N_6885);
or U7056 (N_7056,N_6203,N_6076);
xnor U7057 (N_7057,N_6736,N_6037);
nand U7058 (N_7058,N_6996,N_6252);
nor U7059 (N_7059,N_6889,N_6940);
xnor U7060 (N_7060,N_6044,N_6181);
xnor U7061 (N_7061,N_6314,N_6487);
nand U7062 (N_7062,N_6321,N_6833);
nor U7063 (N_7063,N_6704,N_6832);
xor U7064 (N_7064,N_6271,N_6007);
nor U7065 (N_7065,N_6139,N_6303);
or U7066 (N_7066,N_6290,N_6286);
nand U7067 (N_7067,N_6711,N_6263);
or U7068 (N_7068,N_6517,N_6730);
nor U7069 (N_7069,N_6016,N_6461);
nand U7070 (N_7070,N_6582,N_6818);
nor U7071 (N_7071,N_6075,N_6510);
xor U7072 (N_7072,N_6923,N_6811);
nand U7073 (N_7073,N_6120,N_6732);
nor U7074 (N_7074,N_6723,N_6679);
nor U7075 (N_7075,N_6265,N_6570);
and U7076 (N_7076,N_6858,N_6838);
xnor U7077 (N_7077,N_6867,N_6989);
and U7078 (N_7078,N_6312,N_6426);
or U7079 (N_7079,N_6465,N_6270);
nor U7080 (N_7080,N_6398,N_6035);
and U7081 (N_7081,N_6459,N_6188);
and U7082 (N_7082,N_6038,N_6572);
and U7083 (N_7083,N_6637,N_6186);
or U7084 (N_7084,N_6636,N_6595);
nor U7085 (N_7085,N_6476,N_6187);
nor U7086 (N_7086,N_6686,N_6538);
nor U7087 (N_7087,N_6731,N_6251);
and U7088 (N_7088,N_6432,N_6539);
and U7089 (N_7089,N_6329,N_6255);
nand U7090 (N_7090,N_6953,N_6702);
or U7091 (N_7091,N_6668,N_6755);
xor U7092 (N_7092,N_6019,N_6721);
nor U7093 (N_7093,N_6938,N_6971);
or U7094 (N_7094,N_6706,N_6729);
or U7095 (N_7095,N_6829,N_6896);
or U7096 (N_7096,N_6026,N_6852);
or U7097 (N_7097,N_6220,N_6962);
and U7098 (N_7098,N_6437,N_6165);
or U7099 (N_7099,N_6279,N_6689);
nand U7100 (N_7100,N_6526,N_6501);
or U7101 (N_7101,N_6119,N_6199);
nor U7102 (N_7102,N_6219,N_6213);
xor U7103 (N_7103,N_6293,N_6490);
nand U7104 (N_7104,N_6088,N_6907);
or U7105 (N_7105,N_6936,N_6769);
or U7106 (N_7106,N_6650,N_6389);
nand U7107 (N_7107,N_6400,N_6425);
nand U7108 (N_7108,N_6422,N_6067);
or U7109 (N_7109,N_6772,N_6888);
and U7110 (N_7110,N_6904,N_6536);
or U7111 (N_7111,N_6077,N_6519);
nand U7112 (N_7112,N_6059,N_6795);
nand U7113 (N_7113,N_6735,N_6560);
nor U7114 (N_7114,N_6415,N_6392);
nor U7115 (N_7115,N_6195,N_6357);
nand U7116 (N_7116,N_6423,N_6597);
and U7117 (N_7117,N_6380,N_6522);
xor U7118 (N_7118,N_6891,N_6894);
nand U7119 (N_7119,N_6578,N_6294);
xnor U7120 (N_7120,N_6918,N_6648);
or U7121 (N_7121,N_6903,N_6151);
nand U7122 (N_7122,N_6250,N_6663);
or U7123 (N_7123,N_6960,N_6296);
nand U7124 (N_7124,N_6374,N_6162);
and U7125 (N_7125,N_6453,N_6605);
nand U7126 (N_7126,N_6523,N_6922);
or U7127 (N_7127,N_6238,N_6691);
xnor U7128 (N_7128,N_6790,N_6847);
and U7129 (N_7129,N_6146,N_6987);
xor U7130 (N_7130,N_6403,N_6793);
and U7131 (N_7131,N_6726,N_6068);
nor U7132 (N_7132,N_6930,N_6566);
nor U7133 (N_7133,N_6514,N_6029);
and U7134 (N_7134,N_6099,N_6700);
xor U7135 (N_7135,N_6051,N_6395);
and U7136 (N_7136,N_6023,N_6479);
and U7137 (N_7137,N_6337,N_6977);
or U7138 (N_7138,N_6601,N_6970);
or U7139 (N_7139,N_6406,N_6789);
or U7140 (N_7140,N_6854,N_6865);
nor U7141 (N_7141,N_6025,N_6207);
nor U7142 (N_7142,N_6509,N_6681);
nand U7143 (N_7143,N_6602,N_6261);
nand U7144 (N_7144,N_6671,N_6697);
xor U7145 (N_7145,N_6419,N_6031);
nand U7146 (N_7146,N_6844,N_6225);
nand U7147 (N_7147,N_6665,N_6535);
and U7148 (N_7148,N_6763,N_6608);
nor U7149 (N_7149,N_6017,N_6157);
nand U7150 (N_7150,N_6766,N_6000);
or U7151 (N_7151,N_6592,N_6291);
and U7152 (N_7152,N_6675,N_6061);
nor U7153 (N_7153,N_6863,N_6401);
and U7154 (N_7154,N_6229,N_6197);
nor U7155 (N_7155,N_6179,N_6817);
xor U7156 (N_7156,N_6607,N_6101);
and U7157 (N_7157,N_6028,N_6272);
or U7158 (N_7158,N_6773,N_6114);
and U7159 (N_7159,N_6184,N_6860);
or U7160 (N_7160,N_6375,N_6626);
nor U7161 (N_7161,N_6576,N_6450);
or U7162 (N_7162,N_6468,N_6338);
or U7163 (N_7163,N_6777,N_6963);
nand U7164 (N_7164,N_6483,N_6149);
or U7165 (N_7165,N_6463,N_6623);
nor U7166 (N_7166,N_6335,N_6881);
or U7167 (N_7167,N_6947,N_6192);
nand U7168 (N_7168,N_6444,N_6757);
or U7169 (N_7169,N_6571,N_6990);
xnor U7170 (N_7170,N_6387,N_6491);
and U7171 (N_7171,N_6385,N_6662);
xnor U7172 (N_7172,N_6231,N_6202);
xor U7173 (N_7173,N_6542,N_6246);
and U7174 (N_7174,N_6992,N_6797);
and U7175 (N_7175,N_6481,N_6369);
nand U7176 (N_7176,N_6666,N_6136);
nor U7177 (N_7177,N_6934,N_6647);
xor U7178 (N_7178,N_6127,N_6868);
nor U7179 (N_7179,N_6830,N_6591);
and U7180 (N_7180,N_6448,N_6762);
and U7181 (N_7181,N_6316,N_6175);
or U7182 (N_7182,N_6234,N_6848);
nor U7183 (N_7183,N_6417,N_6244);
xor U7184 (N_7184,N_6627,N_6485);
nor U7185 (N_7185,N_6456,N_6393);
xor U7186 (N_7186,N_6759,N_6057);
nor U7187 (N_7187,N_6325,N_6150);
nand U7188 (N_7188,N_6734,N_6875);
or U7189 (N_7189,N_6512,N_6362);
nand U7190 (N_7190,N_6086,N_6599);
or U7191 (N_7191,N_6682,N_6058);
nand U7192 (N_7192,N_6741,N_6941);
nand U7193 (N_7193,N_6004,N_6484);
nor U7194 (N_7194,N_6386,N_6914);
or U7195 (N_7195,N_6309,N_6190);
and U7196 (N_7196,N_6356,N_6442);
nor U7197 (N_7197,N_6733,N_6978);
xor U7198 (N_7198,N_6331,N_6606);
and U7199 (N_7199,N_6575,N_6091);
nor U7200 (N_7200,N_6014,N_6147);
nor U7201 (N_7201,N_6341,N_6022);
and U7202 (N_7202,N_6427,N_6494);
nand U7203 (N_7203,N_6916,N_6407);
xnor U7204 (N_7204,N_6586,N_6288);
and U7205 (N_7205,N_6205,N_6641);
xor U7206 (N_7206,N_6455,N_6633);
nand U7207 (N_7207,N_6816,N_6160);
xor U7208 (N_7208,N_6887,N_6778);
and U7209 (N_7209,N_6568,N_6724);
nand U7210 (N_7210,N_6171,N_6438);
nand U7211 (N_7211,N_6812,N_6758);
and U7212 (N_7212,N_6241,N_6069);
or U7213 (N_7213,N_6163,N_6553);
xnor U7214 (N_7214,N_6497,N_6761);
nand U7215 (N_7215,N_6254,N_6504);
nand U7216 (N_7216,N_6172,N_6573);
nor U7217 (N_7217,N_6347,N_6843);
nand U7218 (N_7218,N_6826,N_6717);
nor U7219 (N_7219,N_6053,N_6343);
xnor U7220 (N_7220,N_6693,N_6431);
nor U7221 (N_7221,N_6532,N_6630);
and U7222 (N_7222,N_6364,N_6737);
xnor U7223 (N_7223,N_6477,N_6457);
xor U7224 (N_7224,N_6851,N_6267);
or U7225 (N_7225,N_6452,N_6508);
and U7226 (N_7226,N_6527,N_6259);
or U7227 (N_7227,N_6651,N_6893);
xnor U7228 (N_7228,N_6910,N_6897);
and U7229 (N_7229,N_6593,N_6382);
nand U7230 (N_7230,N_6043,N_6024);
nand U7231 (N_7231,N_6625,N_6440);
and U7232 (N_7232,N_6670,N_6342);
nand U7233 (N_7233,N_6545,N_6531);
and U7234 (N_7234,N_6079,N_6055);
and U7235 (N_7235,N_6496,N_6289);
and U7236 (N_7236,N_6421,N_6036);
or U7237 (N_7237,N_6785,N_6466);
and U7238 (N_7238,N_6111,N_6669);
and U7239 (N_7239,N_6615,N_6302);
nand U7240 (N_7240,N_6106,N_6166);
or U7241 (N_7241,N_6307,N_6159);
nor U7242 (N_7242,N_6584,N_6445);
xnor U7243 (N_7243,N_6249,N_6454);
and U7244 (N_7244,N_6915,N_6654);
nand U7245 (N_7245,N_6499,N_6473);
nand U7246 (N_7246,N_6658,N_6742);
xor U7247 (N_7247,N_6937,N_6656);
nor U7248 (N_7248,N_6684,N_6258);
xnor U7249 (N_7249,N_6581,N_6376);
nor U7250 (N_7250,N_6277,N_6676);
and U7251 (N_7251,N_6332,N_6588);
nor U7252 (N_7252,N_6698,N_6547);
and U7253 (N_7253,N_6413,N_6308);
nand U7254 (N_7254,N_6624,N_6805);
xnor U7255 (N_7255,N_6580,N_6680);
and U7256 (N_7256,N_6178,N_6182);
xor U7257 (N_7257,N_6950,N_6351);
and U7258 (N_7258,N_6618,N_6085);
nor U7259 (N_7259,N_6958,N_6033);
and U7260 (N_7260,N_6056,N_6218);
and U7261 (N_7261,N_6831,N_6103);
nor U7262 (N_7262,N_6474,N_6952);
nor U7263 (N_7263,N_6948,N_6315);
and U7264 (N_7264,N_6983,N_6104);
nand U7265 (N_7265,N_6743,N_6718);
nor U7266 (N_7266,N_6169,N_6604);
xor U7267 (N_7267,N_6621,N_6529);
and U7268 (N_7268,N_6804,N_6379);
nand U7269 (N_7269,N_6353,N_6550);
xnor U7270 (N_7270,N_6720,N_6050);
or U7271 (N_7271,N_6064,N_6489);
or U7272 (N_7272,N_6520,N_6791);
or U7273 (N_7273,N_6609,N_6856);
or U7274 (N_7274,N_6807,N_6672);
or U7275 (N_7275,N_6767,N_6108);
or U7276 (N_7276,N_6722,N_6109);
nor U7277 (N_7277,N_6046,N_6673);
nand U7278 (N_7278,N_6653,N_6800);
xor U7279 (N_7279,N_6939,N_6287);
or U7280 (N_7280,N_6541,N_6040);
nand U7281 (N_7281,N_6619,N_6298);
xnor U7282 (N_7282,N_6123,N_6430);
xnor U7283 (N_7283,N_6925,N_6657);
and U7284 (N_7284,N_6557,N_6200);
or U7285 (N_7285,N_6012,N_6874);
nor U7286 (N_7286,N_6810,N_6911);
or U7287 (N_7287,N_6909,N_6823);
or U7288 (N_7288,N_6222,N_6513);
xor U7289 (N_7289,N_6121,N_6102);
and U7290 (N_7290,N_6340,N_6969);
nor U7291 (N_7291,N_6982,N_6782);
nand U7292 (N_7292,N_6642,N_6048);
xnor U7293 (N_7293,N_6300,N_6746);
nand U7294 (N_7294,N_6269,N_6886);
or U7295 (N_7295,N_6138,N_6324);
nor U7296 (N_7296,N_6629,N_6381);
and U7297 (N_7297,N_6273,N_6943);
nor U7298 (N_7298,N_6168,N_6281);
xor U7299 (N_7299,N_6446,N_6140);
xor U7300 (N_7300,N_6927,N_6212);
nor U7301 (N_7301,N_6835,N_6383);
nor U7302 (N_7302,N_6041,N_6871);
or U7303 (N_7303,N_6635,N_6879);
or U7304 (N_7304,N_6942,N_6420);
nand U7305 (N_7305,N_6564,N_6095);
and U7306 (N_7306,N_6685,N_6745);
or U7307 (N_7307,N_6274,N_6208);
xor U7308 (N_7308,N_6153,N_6228);
and U7309 (N_7309,N_6546,N_6295);
nor U7310 (N_7310,N_6310,N_6148);
nor U7311 (N_7311,N_6248,N_6034);
nor U7312 (N_7312,N_6997,N_6117);
or U7313 (N_7313,N_6326,N_6367);
nor U7314 (N_7314,N_6774,N_6821);
and U7315 (N_7315,N_6890,N_6128);
or U7316 (N_7316,N_6247,N_6236);
nor U7317 (N_7317,N_6562,N_6352);
and U7318 (N_7318,N_6770,N_6808);
xnor U7319 (N_7319,N_6544,N_6396);
xor U7320 (N_7320,N_6906,N_6311);
nor U7321 (N_7321,N_6981,N_6317);
or U7322 (N_7322,N_6333,N_6660);
and U7323 (N_7323,N_6074,N_6974);
nand U7324 (N_7324,N_6873,N_6257);
nor U7325 (N_7325,N_6414,N_6701);
and U7326 (N_7326,N_6714,N_6819);
and U7327 (N_7327,N_6898,N_6092);
and U7328 (N_7328,N_6577,N_6728);
and U7329 (N_7329,N_6809,N_6610);
nand U7330 (N_7330,N_6853,N_6170);
nor U7331 (N_7331,N_6946,N_6622);
xor U7332 (N_7332,N_6908,N_6105);
or U7333 (N_7333,N_6781,N_6827);
nand U7334 (N_7334,N_6411,N_6011);
nand U7335 (N_7335,N_6901,N_6015);
xor U7336 (N_7336,N_6285,N_6365);
nand U7337 (N_7337,N_6643,N_6409);
nand U7338 (N_7338,N_6211,N_6661);
and U7339 (N_7339,N_6846,N_6451);
xor U7340 (N_7340,N_6495,N_6929);
nor U7341 (N_7341,N_6235,N_6801);
nor U7342 (N_7342,N_6436,N_6042);
or U7343 (N_7343,N_6511,N_6134);
nor U7344 (N_7344,N_6707,N_6083);
nand U7345 (N_7345,N_6725,N_6339);
nand U7346 (N_7346,N_6078,N_6613);
xnor U7347 (N_7347,N_6839,N_6471);
xor U7348 (N_7348,N_6328,N_6084);
and U7349 (N_7349,N_6439,N_6330);
xor U7350 (N_7350,N_6788,N_6528);
or U7351 (N_7351,N_6935,N_6469);
xor U7352 (N_7352,N_6695,N_6283);
nor U7353 (N_7353,N_6899,N_6815);
xor U7354 (N_7354,N_6859,N_6405);
or U7355 (N_7355,N_6486,N_6866);
and U7356 (N_7356,N_6921,N_6708);
xor U7357 (N_7357,N_6783,N_6080);
nand U7358 (N_7358,N_6350,N_6598);
nand U7359 (N_7359,N_6750,N_6612);
or U7360 (N_7360,N_6503,N_6559);
and U7361 (N_7361,N_6820,N_6966);
and U7362 (N_7362,N_6964,N_6984);
xor U7363 (N_7363,N_6275,N_6505);
nand U7364 (N_7364,N_6470,N_6073);
nor U7365 (N_7365,N_6928,N_6173);
and U7366 (N_7366,N_6926,N_6441);
or U7367 (N_7367,N_6537,N_6334);
xnor U7368 (N_7368,N_6129,N_6460);
and U7369 (N_7369,N_6845,N_6855);
or U7370 (N_7370,N_6378,N_6998);
and U7371 (N_7371,N_6744,N_6716);
and U7372 (N_7372,N_6204,N_6164);
xnor U7373 (N_7373,N_6253,N_6390);
xnor U7374 (N_7374,N_6118,N_6683);
xor U7375 (N_7375,N_6802,N_6552);
nand U7376 (N_7376,N_6478,N_6399);
xor U7377 (N_7377,N_6739,N_6434);
or U7378 (N_7378,N_6877,N_6779);
and U7379 (N_7379,N_6920,N_6999);
or U7380 (N_7380,N_6433,N_6824);
or U7381 (N_7381,N_6524,N_6297);
and U7382 (N_7382,N_6664,N_6563);
nor U7383 (N_7383,N_6087,N_6749);
nor U7384 (N_7384,N_6752,N_6174);
and U7385 (N_7385,N_6005,N_6227);
or U7386 (N_7386,N_6884,N_6985);
nor U7387 (N_7387,N_6278,N_6292);
and U7388 (N_7388,N_6107,N_6322);
and U7389 (N_7389,N_6919,N_6876);
or U7390 (N_7390,N_6193,N_6358);
nand U7391 (N_7391,N_6346,N_6206);
nor U7392 (N_7392,N_6214,N_6710);
xnor U7393 (N_7393,N_6836,N_6349);
xnor U7394 (N_7394,N_6587,N_6872);
nor U7395 (N_7395,N_6548,N_6096);
nand U7396 (N_7396,N_6786,N_6180);
nor U7397 (N_7397,N_6115,N_6097);
xor U7398 (N_7398,N_6912,N_6703);
nand U7399 (N_7399,N_6549,N_6137);
or U7400 (N_7400,N_6902,N_6533);
or U7401 (N_7401,N_6632,N_6933);
nand U7402 (N_7402,N_6305,N_6047);
or U7403 (N_7403,N_6840,N_6435);
xor U7404 (N_7404,N_6464,N_6768);
xor U7405 (N_7405,N_6883,N_6082);
or U7406 (N_7406,N_6155,N_6878);
nand U7407 (N_7407,N_6645,N_6001);
or U7408 (N_7408,N_6589,N_6260);
or U7409 (N_7409,N_6388,N_6130);
xor U7410 (N_7410,N_6093,N_6424);
and U7411 (N_7411,N_6198,N_6780);
or U7412 (N_7412,N_6488,N_6688);
nand U7413 (N_7413,N_6652,N_6565);
nand U7414 (N_7414,N_6994,N_6125);
or U7415 (N_7415,N_6299,N_6002);
xnor U7416 (N_7416,N_6354,N_6245);
nor U7417 (N_7417,N_6116,N_6458);
nand U7418 (N_7418,N_6784,N_6009);
nor U7419 (N_7419,N_6677,N_6776);
nand U7420 (N_7420,N_6727,N_6443);
and U7421 (N_7421,N_6850,N_6428);
and U7422 (N_7422,N_6062,N_6699);
nor U7423 (N_7423,N_6183,N_6010);
and U7424 (N_7424,N_6751,N_6995);
nand U7425 (N_7425,N_6521,N_6418);
nand U7426 (N_7426,N_6540,N_6771);
nor U7427 (N_7427,N_6813,N_6132);
nor U7428 (N_7428,N_6760,N_6798);
or U7429 (N_7429,N_6320,N_6561);
nand U7430 (N_7430,N_6590,N_6394);
or U7431 (N_7431,N_6177,N_6408);
nand U7432 (N_7432,N_6366,N_6895);
and U7433 (N_7433,N_6659,N_6674);
or U7434 (N_7434,N_6126,N_6027);
and U7435 (N_7435,N_6965,N_6216);
nand U7436 (N_7436,N_6189,N_6063);
and U7437 (N_7437,N_6567,N_6516);
nor U7438 (N_7438,N_6239,N_6039);
nor U7439 (N_7439,N_6045,N_6221);
nor U7440 (N_7440,N_6525,N_6882);
nor U7441 (N_7441,N_6124,N_6530);
and U7442 (N_7442,N_6167,N_6447);
nand U7443 (N_7443,N_6304,N_6256);
and U7444 (N_7444,N_6611,N_6049);
nand U7445 (N_7445,N_6144,N_6543);
or U7446 (N_7446,N_6306,N_6429);
nand U7447 (N_7447,N_6765,N_6869);
nor U7448 (N_7448,N_6006,N_6133);
nand U7449 (N_7449,N_6161,N_6154);
and U7450 (N_7450,N_6870,N_6327);
nor U7451 (N_7451,N_6412,N_6100);
and U7452 (N_7452,N_6556,N_6098);
xor U7453 (N_7453,N_6377,N_6694);
xnor U7454 (N_7454,N_6355,N_6803);
and U7455 (N_7455,N_6892,N_6951);
xnor U7456 (N_7456,N_6917,N_6318);
xnor U7457 (N_7457,N_6967,N_6583);
or U7458 (N_7458,N_6240,N_6709);
or U7459 (N_7459,N_6052,N_6705);
nor U7460 (N_7460,N_6614,N_6373);
or U7461 (N_7461,N_6472,N_6506);
xor U7462 (N_7462,N_6924,N_6493);
or U7463 (N_7463,N_6972,N_6368);
nor U7464 (N_7464,N_6384,N_6634);
or U7465 (N_7465,N_6266,N_6574);
or U7466 (N_7466,N_6135,N_6467);
xor U7467 (N_7467,N_6991,N_6264);
nand U7468 (N_7468,N_6594,N_6988);
nor U7469 (N_7469,N_6361,N_6008);
xnor U7470 (N_7470,N_6502,N_6416);
or U7471 (N_7471,N_6475,N_6113);
xor U7472 (N_7472,N_6579,N_6018);
nor U7473 (N_7473,N_6323,N_6979);
nand U7474 (N_7474,N_6796,N_6176);
and U7475 (N_7475,N_6223,N_6066);
nor U7476 (N_7476,N_6980,N_6900);
nor U7477 (N_7477,N_6237,N_6276);
xnor U7478 (N_7478,N_6498,N_6344);
and U7479 (N_7479,N_6372,N_6806);
nor U7480 (N_7480,N_6959,N_6345);
or U7481 (N_7481,N_6603,N_6640);
or U7482 (N_7482,N_6156,N_6825);
nor U7483 (N_7483,N_6655,N_6555);
nand U7484 (N_7484,N_6864,N_6551);
and U7485 (N_7485,N_6631,N_6973);
and U7486 (N_7486,N_6834,N_6518);
nor U7487 (N_7487,N_6215,N_6360);
nand U7488 (N_7488,N_6678,N_6313);
xnor U7489 (N_7489,N_6862,N_6849);
nor U7490 (N_7490,N_6094,N_6787);
xor U7491 (N_7491,N_6462,N_6194);
nand U7492 (N_7492,N_6794,N_6348);
xnor U7493 (N_7493,N_6143,N_6243);
xor U7494 (N_7494,N_6616,N_6224);
xor U7495 (N_7495,N_6131,N_6021);
xor U7496 (N_7496,N_6122,N_6301);
nor U7497 (N_7497,N_6554,N_6158);
and U7498 (N_7498,N_6692,N_6993);
xor U7499 (N_7499,N_6284,N_6226);
nor U7500 (N_7500,N_6017,N_6282);
and U7501 (N_7501,N_6430,N_6973);
nor U7502 (N_7502,N_6168,N_6999);
nand U7503 (N_7503,N_6040,N_6686);
nor U7504 (N_7504,N_6970,N_6349);
nand U7505 (N_7505,N_6908,N_6790);
xor U7506 (N_7506,N_6650,N_6916);
nand U7507 (N_7507,N_6859,N_6623);
nor U7508 (N_7508,N_6341,N_6762);
xnor U7509 (N_7509,N_6129,N_6135);
nor U7510 (N_7510,N_6039,N_6289);
nor U7511 (N_7511,N_6463,N_6127);
nand U7512 (N_7512,N_6437,N_6111);
or U7513 (N_7513,N_6351,N_6870);
xnor U7514 (N_7514,N_6097,N_6947);
nand U7515 (N_7515,N_6709,N_6231);
nor U7516 (N_7516,N_6377,N_6604);
and U7517 (N_7517,N_6024,N_6388);
xor U7518 (N_7518,N_6669,N_6810);
nand U7519 (N_7519,N_6164,N_6866);
or U7520 (N_7520,N_6774,N_6792);
xnor U7521 (N_7521,N_6271,N_6581);
xnor U7522 (N_7522,N_6175,N_6771);
nor U7523 (N_7523,N_6432,N_6788);
or U7524 (N_7524,N_6254,N_6952);
and U7525 (N_7525,N_6591,N_6075);
or U7526 (N_7526,N_6742,N_6171);
nor U7527 (N_7527,N_6784,N_6334);
or U7528 (N_7528,N_6192,N_6564);
and U7529 (N_7529,N_6925,N_6064);
or U7530 (N_7530,N_6026,N_6425);
or U7531 (N_7531,N_6953,N_6515);
nand U7532 (N_7532,N_6452,N_6936);
nor U7533 (N_7533,N_6994,N_6948);
and U7534 (N_7534,N_6763,N_6779);
xnor U7535 (N_7535,N_6127,N_6551);
or U7536 (N_7536,N_6790,N_6244);
nor U7537 (N_7537,N_6933,N_6887);
xnor U7538 (N_7538,N_6692,N_6559);
xnor U7539 (N_7539,N_6031,N_6139);
and U7540 (N_7540,N_6246,N_6023);
xnor U7541 (N_7541,N_6559,N_6128);
and U7542 (N_7542,N_6106,N_6532);
xnor U7543 (N_7543,N_6445,N_6180);
and U7544 (N_7544,N_6053,N_6042);
or U7545 (N_7545,N_6697,N_6903);
or U7546 (N_7546,N_6447,N_6041);
nand U7547 (N_7547,N_6231,N_6907);
nand U7548 (N_7548,N_6262,N_6688);
nand U7549 (N_7549,N_6673,N_6413);
or U7550 (N_7550,N_6213,N_6053);
nand U7551 (N_7551,N_6710,N_6786);
nor U7552 (N_7552,N_6256,N_6958);
nor U7553 (N_7553,N_6813,N_6069);
nand U7554 (N_7554,N_6163,N_6654);
or U7555 (N_7555,N_6387,N_6190);
nor U7556 (N_7556,N_6707,N_6923);
nand U7557 (N_7557,N_6639,N_6734);
xnor U7558 (N_7558,N_6908,N_6939);
xor U7559 (N_7559,N_6732,N_6444);
xor U7560 (N_7560,N_6294,N_6645);
nor U7561 (N_7561,N_6152,N_6201);
nand U7562 (N_7562,N_6864,N_6657);
xnor U7563 (N_7563,N_6406,N_6759);
xnor U7564 (N_7564,N_6014,N_6952);
xor U7565 (N_7565,N_6130,N_6883);
or U7566 (N_7566,N_6713,N_6311);
xor U7567 (N_7567,N_6876,N_6460);
and U7568 (N_7568,N_6055,N_6327);
and U7569 (N_7569,N_6315,N_6080);
nor U7570 (N_7570,N_6102,N_6125);
and U7571 (N_7571,N_6075,N_6576);
xor U7572 (N_7572,N_6877,N_6588);
nor U7573 (N_7573,N_6508,N_6009);
xnor U7574 (N_7574,N_6511,N_6864);
and U7575 (N_7575,N_6290,N_6384);
or U7576 (N_7576,N_6526,N_6117);
or U7577 (N_7577,N_6329,N_6207);
or U7578 (N_7578,N_6274,N_6093);
and U7579 (N_7579,N_6067,N_6337);
xnor U7580 (N_7580,N_6855,N_6693);
nor U7581 (N_7581,N_6078,N_6264);
nor U7582 (N_7582,N_6662,N_6295);
nand U7583 (N_7583,N_6836,N_6521);
xnor U7584 (N_7584,N_6305,N_6670);
and U7585 (N_7585,N_6009,N_6686);
nand U7586 (N_7586,N_6562,N_6651);
nand U7587 (N_7587,N_6157,N_6400);
nor U7588 (N_7588,N_6155,N_6783);
or U7589 (N_7589,N_6508,N_6121);
nor U7590 (N_7590,N_6323,N_6652);
and U7591 (N_7591,N_6934,N_6257);
xor U7592 (N_7592,N_6775,N_6640);
nand U7593 (N_7593,N_6958,N_6311);
nor U7594 (N_7594,N_6654,N_6036);
or U7595 (N_7595,N_6841,N_6632);
nor U7596 (N_7596,N_6066,N_6180);
xor U7597 (N_7597,N_6081,N_6289);
nand U7598 (N_7598,N_6902,N_6881);
and U7599 (N_7599,N_6710,N_6531);
nand U7600 (N_7600,N_6651,N_6953);
or U7601 (N_7601,N_6274,N_6977);
xor U7602 (N_7602,N_6431,N_6734);
nand U7603 (N_7603,N_6397,N_6177);
xnor U7604 (N_7604,N_6904,N_6268);
nor U7605 (N_7605,N_6979,N_6748);
or U7606 (N_7606,N_6713,N_6039);
and U7607 (N_7607,N_6871,N_6229);
or U7608 (N_7608,N_6070,N_6010);
nand U7609 (N_7609,N_6541,N_6281);
xor U7610 (N_7610,N_6653,N_6496);
nand U7611 (N_7611,N_6958,N_6712);
nor U7612 (N_7612,N_6863,N_6148);
nor U7613 (N_7613,N_6552,N_6347);
or U7614 (N_7614,N_6691,N_6190);
and U7615 (N_7615,N_6421,N_6353);
and U7616 (N_7616,N_6010,N_6494);
nand U7617 (N_7617,N_6964,N_6345);
or U7618 (N_7618,N_6362,N_6223);
or U7619 (N_7619,N_6801,N_6499);
nor U7620 (N_7620,N_6039,N_6187);
or U7621 (N_7621,N_6963,N_6556);
or U7622 (N_7622,N_6945,N_6588);
nor U7623 (N_7623,N_6768,N_6912);
or U7624 (N_7624,N_6921,N_6726);
and U7625 (N_7625,N_6701,N_6622);
xnor U7626 (N_7626,N_6207,N_6614);
nand U7627 (N_7627,N_6738,N_6250);
nor U7628 (N_7628,N_6260,N_6918);
nand U7629 (N_7629,N_6290,N_6039);
nor U7630 (N_7630,N_6030,N_6539);
nor U7631 (N_7631,N_6042,N_6542);
or U7632 (N_7632,N_6757,N_6987);
or U7633 (N_7633,N_6755,N_6056);
nand U7634 (N_7634,N_6356,N_6001);
or U7635 (N_7635,N_6463,N_6752);
or U7636 (N_7636,N_6604,N_6200);
nor U7637 (N_7637,N_6391,N_6131);
nor U7638 (N_7638,N_6646,N_6884);
xor U7639 (N_7639,N_6868,N_6817);
xor U7640 (N_7640,N_6200,N_6587);
nor U7641 (N_7641,N_6779,N_6080);
and U7642 (N_7642,N_6583,N_6812);
or U7643 (N_7643,N_6935,N_6175);
xnor U7644 (N_7644,N_6824,N_6919);
nand U7645 (N_7645,N_6363,N_6635);
nand U7646 (N_7646,N_6900,N_6147);
or U7647 (N_7647,N_6730,N_6556);
nand U7648 (N_7648,N_6540,N_6585);
or U7649 (N_7649,N_6552,N_6043);
and U7650 (N_7650,N_6170,N_6073);
nor U7651 (N_7651,N_6533,N_6027);
xnor U7652 (N_7652,N_6686,N_6109);
or U7653 (N_7653,N_6929,N_6269);
nor U7654 (N_7654,N_6186,N_6625);
nor U7655 (N_7655,N_6890,N_6238);
xnor U7656 (N_7656,N_6391,N_6937);
nand U7657 (N_7657,N_6197,N_6796);
and U7658 (N_7658,N_6851,N_6975);
nand U7659 (N_7659,N_6985,N_6325);
nand U7660 (N_7660,N_6122,N_6191);
and U7661 (N_7661,N_6648,N_6375);
nand U7662 (N_7662,N_6954,N_6121);
or U7663 (N_7663,N_6624,N_6992);
xnor U7664 (N_7664,N_6370,N_6931);
and U7665 (N_7665,N_6970,N_6854);
nand U7666 (N_7666,N_6029,N_6389);
nor U7667 (N_7667,N_6336,N_6344);
xor U7668 (N_7668,N_6339,N_6755);
xnor U7669 (N_7669,N_6570,N_6808);
nand U7670 (N_7670,N_6618,N_6749);
xnor U7671 (N_7671,N_6929,N_6267);
nor U7672 (N_7672,N_6300,N_6191);
or U7673 (N_7673,N_6609,N_6690);
nand U7674 (N_7674,N_6500,N_6598);
xnor U7675 (N_7675,N_6021,N_6016);
or U7676 (N_7676,N_6780,N_6559);
xor U7677 (N_7677,N_6871,N_6546);
xor U7678 (N_7678,N_6139,N_6808);
or U7679 (N_7679,N_6736,N_6211);
nand U7680 (N_7680,N_6043,N_6834);
nor U7681 (N_7681,N_6271,N_6634);
nand U7682 (N_7682,N_6811,N_6725);
and U7683 (N_7683,N_6777,N_6473);
and U7684 (N_7684,N_6163,N_6316);
and U7685 (N_7685,N_6145,N_6651);
or U7686 (N_7686,N_6087,N_6805);
xnor U7687 (N_7687,N_6840,N_6697);
nand U7688 (N_7688,N_6298,N_6305);
xnor U7689 (N_7689,N_6097,N_6544);
or U7690 (N_7690,N_6059,N_6595);
xnor U7691 (N_7691,N_6370,N_6035);
and U7692 (N_7692,N_6666,N_6822);
and U7693 (N_7693,N_6732,N_6447);
xor U7694 (N_7694,N_6331,N_6889);
or U7695 (N_7695,N_6299,N_6645);
xor U7696 (N_7696,N_6954,N_6464);
and U7697 (N_7697,N_6912,N_6753);
nand U7698 (N_7698,N_6168,N_6195);
xor U7699 (N_7699,N_6776,N_6143);
nor U7700 (N_7700,N_6567,N_6342);
nand U7701 (N_7701,N_6408,N_6134);
and U7702 (N_7702,N_6289,N_6481);
nand U7703 (N_7703,N_6503,N_6166);
xor U7704 (N_7704,N_6337,N_6333);
nor U7705 (N_7705,N_6533,N_6883);
xnor U7706 (N_7706,N_6502,N_6496);
nand U7707 (N_7707,N_6388,N_6416);
or U7708 (N_7708,N_6263,N_6435);
xnor U7709 (N_7709,N_6752,N_6170);
and U7710 (N_7710,N_6433,N_6299);
and U7711 (N_7711,N_6613,N_6586);
nand U7712 (N_7712,N_6948,N_6769);
and U7713 (N_7713,N_6416,N_6196);
nand U7714 (N_7714,N_6982,N_6814);
nor U7715 (N_7715,N_6859,N_6461);
nand U7716 (N_7716,N_6486,N_6736);
nand U7717 (N_7717,N_6455,N_6586);
nor U7718 (N_7718,N_6417,N_6976);
nor U7719 (N_7719,N_6781,N_6289);
nor U7720 (N_7720,N_6620,N_6717);
xor U7721 (N_7721,N_6246,N_6564);
and U7722 (N_7722,N_6147,N_6219);
xor U7723 (N_7723,N_6859,N_6249);
nor U7724 (N_7724,N_6045,N_6069);
nand U7725 (N_7725,N_6243,N_6940);
xnor U7726 (N_7726,N_6924,N_6962);
and U7727 (N_7727,N_6155,N_6501);
nand U7728 (N_7728,N_6962,N_6487);
xor U7729 (N_7729,N_6573,N_6294);
xnor U7730 (N_7730,N_6235,N_6456);
and U7731 (N_7731,N_6039,N_6231);
and U7732 (N_7732,N_6073,N_6098);
or U7733 (N_7733,N_6567,N_6133);
and U7734 (N_7734,N_6885,N_6557);
or U7735 (N_7735,N_6944,N_6759);
nor U7736 (N_7736,N_6391,N_6399);
xnor U7737 (N_7737,N_6816,N_6285);
xnor U7738 (N_7738,N_6555,N_6117);
or U7739 (N_7739,N_6775,N_6734);
and U7740 (N_7740,N_6593,N_6226);
nand U7741 (N_7741,N_6613,N_6066);
nand U7742 (N_7742,N_6258,N_6402);
nor U7743 (N_7743,N_6491,N_6606);
xor U7744 (N_7744,N_6731,N_6730);
or U7745 (N_7745,N_6323,N_6715);
nor U7746 (N_7746,N_6269,N_6568);
and U7747 (N_7747,N_6016,N_6471);
nor U7748 (N_7748,N_6821,N_6755);
nand U7749 (N_7749,N_6506,N_6348);
or U7750 (N_7750,N_6096,N_6116);
and U7751 (N_7751,N_6960,N_6929);
and U7752 (N_7752,N_6234,N_6665);
nor U7753 (N_7753,N_6682,N_6626);
and U7754 (N_7754,N_6402,N_6347);
xnor U7755 (N_7755,N_6120,N_6147);
and U7756 (N_7756,N_6646,N_6030);
or U7757 (N_7757,N_6225,N_6108);
nor U7758 (N_7758,N_6102,N_6290);
nor U7759 (N_7759,N_6830,N_6053);
and U7760 (N_7760,N_6448,N_6109);
and U7761 (N_7761,N_6671,N_6256);
or U7762 (N_7762,N_6708,N_6172);
nor U7763 (N_7763,N_6019,N_6164);
nor U7764 (N_7764,N_6613,N_6900);
nand U7765 (N_7765,N_6170,N_6450);
or U7766 (N_7766,N_6246,N_6836);
nand U7767 (N_7767,N_6039,N_6210);
nor U7768 (N_7768,N_6850,N_6920);
and U7769 (N_7769,N_6427,N_6234);
nor U7770 (N_7770,N_6400,N_6424);
xnor U7771 (N_7771,N_6793,N_6834);
nor U7772 (N_7772,N_6216,N_6168);
or U7773 (N_7773,N_6209,N_6198);
nand U7774 (N_7774,N_6215,N_6625);
and U7775 (N_7775,N_6539,N_6932);
xor U7776 (N_7776,N_6195,N_6791);
nand U7777 (N_7777,N_6313,N_6041);
nor U7778 (N_7778,N_6975,N_6609);
nor U7779 (N_7779,N_6402,N_6427);
and U7780 (N_7780,N_6002,N_6190);
nand U7781 (N_7781,N_6709,N_6674);
or U7782 (N_7782,N_6310,N_6263);
nand U7783 (N_7783,N_6245,N_6818);
nand U7784 (N_7784,N_6063,N_6456);
and U7785 (N_7785,N_6631,N_6832);
or U7786 (N_7786,N_6298,N_6697);
nand U7787 (N_7787,N_6363,N_6781);
or U7788 (N_7788,N_6283,N_6054);
xor U7789 (N_7789,N_6536,N_6804);
and U7790 (N_7790,N_6245,N_6949);
nand U7791 (N_7791,N_6916,N_6440);
or U7792 (N_7792,N_6472,N_6579);
or U7793 (N_7793,N_6074,N_6222);
xor U7794 (N_7794,N_6461,N_6415);
xor U7795 (N_7795,N_6533,N_6460);
and U7796 (N_7796,N_6241,N_6637);
xnor U7797 (N_7797,N_6568,N_6758);
nand U7798 (N_7798,N_6484,N_6763);
nor U7799 (N_7799,N_6980,N_6882);
nand U7800 (N_7800,N_6087,N_6471);
or U7801 (N_7801,N_6302,N_6594);
and U7802 (N_7802,N_6708,N_6691);
nor U7803 (N_7803,N_6064,N_6797);
and U7804 (N_7804,N_6227,N_6601);
and U7805 (N_7805,N_6465,N_6272);
or U7806 (N_7806,N_6383,N_6553);
nor U7807 (N_7807,N_6370,N_6793);
nor U7808 (N_7808,N_6195,N_6792);
or U7809 (N_7809,N_6972,N_6453);
and U7810 (N_7810,N_6496,N_6741);
and U7811 (N_7811,N_6881,N_6128);
or U7812 (N_7812,N_6254,N_6777);
xnor U7813 (N_7813,N_6979,N_6819);
nor U7814 (N_7814,N_6356,N_6664);
nor U7815 (N_7815,N_6640,N_6161);
and U7816 (N_7816,N_6381,N_6545);
and U7817 (N_7817,N_6905,N_6817);
and U7818 (N_7818,N_6238,N_6718);
xor U7819 (N_7819,N_6166,N_6641);
nand U7820 (N_7820,N_6860,N_6830);
nor U7821 (N_7821,N_6358,N_6057);
nor U7822 (N_7822,N_6057,N_6586);
nand U7823 (N_7823,N_6145,N_6399);
xnor U7824 (N_7824,N_6663,N_6120);
and U7825 (N_7825,N_6781,N_6372);
or U7826 (N_7826,N_6276,N_6422);
and U7827 (N_7827,N_6110,N_6062);
nor U7828 (N_7828,N_6337,N_6445);
and U7829 (N_7829,N_6202,N_6288);
or U7830 (N_7830,N_6700,N_6309);
nor U7831 (N_7831,N_6043,N_6723);
nor U7832 (N_7832,N_6330,N_6615);
and U7833 (N_7833,N_6105,N_6681);
or U7834 (N_7834,N_6827,N_6033);
or U7835 (N_7835,N_6950,N_6072);
or U7836 (N_7836,N_6924,N_6006);
or U7837 (N_7837,N_6024,N_6951);
and U7838 (N_7838,N_6319,N_6293);
nor U7839 (N_7839,N_6069,N_6468);
or U7840 (N_7840,N_6471,N_6904);
and U7841 (N_7841,N_6139,N_6086);
nor U7842 (N_7842,N_6288,N_6469);
xnor U7843 (N_7843,N_6337,N_6706);
and U7844 (N_7844,N_6800,N_6146);
xor U7845 (N_7845,N_6196,N_6068);
and U7846 (N_7846,N_6986,N_6930);
or U7847 (N_7847,N_6524,N_6770);
xor U7848 (N_7848,N_6202,N_6337);
nor U7849 (N_7849,N_6204,N_6247);
nand U7850 (N_7850,N_6000,N_6118);
nand U7851 (N_7851,N_6194,N_6206);
and U7852 (N_7852,N_6284,N_6704);
nand U7853 (N_7853,N_6937,N_6235);
nand U7854 (N_7854,N_6411,N_6465);
or U7855 (N_7855,N_6443,N_6099);
and U7856 (N_7856,N_6738,N_6645);
or U7857 (N_7857,N_6436,N_6066);
or U7858 (N_7858,N_6749,N_6900);
nand U7859 (N_7859,N_6760,N_6105);
xnor U7860 (N_7860,N_6346,N_6128);
and U7861 (N_7861,N_6830,N_6321);
and U7862 (N_7862,N_6321,N_6202);
nand U7863 (N_7863,N_6673,N_6550);
or U7864 (N_7864,N_6375,N_6605);
xor U7865 (N_7865,N_6047,N_6027);
and U7866 (N_7866,N_6663,N_6929);
nor U7867 (N_7867,N_6470,N_6597);
nor U7868 (N_7868,N_6136,N_6884);
or U7869 (N_7869,N_6890,N_6118);
nand U7870 (N_7870,N_6210,N_6951);
xor U7871 (N_7871,N_6408,N_6417);
xnor U7872 (N_7872,N_6038,N_6273);
or U7873 (N_7873,N_6600,N_6921);
nor U7874 (N_7874,N_6758,N_6289);
nand U7875 (N_7875,N_6291,N_6348);
nor U7876 (N_7876,N_6782,N_6896);
xor U7877 (N_7877,N_6341,N_6591);
nand U7878 (N_7878,N_6391,N_6134);
or U7879 (N_7879,N_6816,N_6746);
nor U7880 (N_7880,N_6384,N_6288);
or U7881 (N_7881,N_6043,N_6508);
nand U7882 (N_7882,N_6303,N_6636);
or U7883 (N_7883,N_6022,N_6071);
nor U7884 (N_7884,N_6955,N_6522);
and U7885 (N_7885,N_6586,N_6067);
nand U7886 (N_7886,N_6279,N_6776);
nand U7887 (N_7887,N_6988,N_6722);
or U7888 (N_7888,N_6311,N_6435);
nand U7889 (N_7889,N_6692,N_6340);
or U7890 (N_7890,N_6855,N_6764);
nand U7891 (N_7891,N_6145,N_6711);
nand U7892 (N_7892,N_6951,N_6760);
nand U7893 (N_7893,N_6349,N_6220);
xor U7894 (N_7894,N_6743,N_6603);
nor U7895 (N_7895,N_6473,N_6452);
xnor U7896 (N_7896,N_6455,N_6167);
or U7897 (N_7897,N_6905,N_6488);
nor U7898 (N_7898,N_6211,N_6636);
nor U7899 (N_7899,N_6878,N_6196);
nor U7900 (N_7900,N_6399,N_6264);
nand U7901 (N_7901,N_6696,N_6389);
nand U7902 (N_7902,N_6433,N_6229);
nand U7903 (N_7903,N_6953,N_6386);
xor U7904 (N_7904,N_6397,N_6928);
nand U7905 (N_7905,N_6277,N_6476);
and U7906 (N_7906,N_6582,N_6139);
or U7907 (N_7907,N_6183,N_6859);
and U7908 (N_7908,N_6648,N_6255);
nand U7909 (N_7909,N_6937,N_6759);
and U7910 (N_7910,N_6211,N_6921);
and U7911 (N_7911,N_6929,N_6233);
xnor U7912 (N_7912,N_6407,N_6256);
or U7913 (N_7913,N_6990,N_6369);
and U7914 (N_7914,N_6047,N_6186);
nand U7915 (N_7915,N_6323,N_6320);
xor U7916 (N_7916,N_6607,N_6247);
xnor U7917 (N_7917,N_6635,N_6766);
and U7918 (N_7918,N_6907,N_6423);
and U7919 (N_7919,N_6912,N_6459);
nor U7920 (N_7920,N_6927,N_6239);
or U7921 (N_7921,N_6856,N_6054);
and U7922 (N_7922,N_6002,N_6119);
nand U7923 (N_7923,N_6952,N_6040);
or U7924 (N_7924,N_6821,N_6218);
nand U7925 (N_7925,N_6194,N_6963);
and U7926 (N_7926,N_6596,N_6294);
nand U7927 (N_7927,N_6285,N_6622);
nor U7928 (N_7928,N_6333,N_6745);
xor U7929 (N_7929,N_6399,N_6480);
nor U7930 (N_7930,N_6392,N_6993);
nand U7931 (N_7931,N_6814,N_6199);
or U7932 (N_7932,N_6001,N_6929);
or U7933 (N_7933,N_6085,N_6776);
and U7934 (N_7934,N_6002,N_6293);
xor U7935 (N_7935,N_6601,N_6698);
xor U7936 (N_7936,N_6162,N_6252);
xor U7937 (N_7937,N_6465,N_6178);
and U7938 (N_7938,N_6142,N_6512);
nand U7939 (N_7939,N_6137,N_6046);
nand U7940 (N_7940,N_6972,N_6328);
and U7941 (N_7941,N_6255,N_6050);
nor U7942 (N_7942,N_6137,N_6069);
or U7943 (N_7943,N_6713,N_6665);
nand U7944 (N_7944,N_6868,N_6687);
nand U7945 (N_7945,N_6328,N_6611);
and U7946 (N_7946,N_6510,N_6584);
and U7947 (N_7947,N_6998,N_6752);
and U7948 (N_7948,N_6494,N_6712);
nand U7949 (N_7949,N_6928,N_6149);
nand U7950 (N_7950,N_6153,N_6595);
xor U7951 (N_7951,N_6749,N_6671);
xor U7952 (N_7952,N_6490,N_6748);
xnor U7953 (N_7953,N_6480,N_6673);
and U7954 (N_7954,N_6029,N_6600);
xnor U7955 (N_7955,N_6966,N_6427);
nand U7956 (N_7956,N_6759,N_6461);
nand U7957 (N_7957,N_6018,N_6194);
or U7958 (N_7958,N_6067,N_6208);
or U7959 (N_7959,N_6148,N_6160);
nand U7960 (N_7960,N_6250,N_6601);
nand U7961 (N_7961,N_6111,N_6780);
nand U7962 (N_7962,N_6760,N_6553);
xnor U7963 (N_7963,N_6597,N_6065);
nor U7964 (N_7964,N_6055,N_6734);
and U7965 (N_7965,N_6689,N_6187);
and U7966 (N_7966,N_6616,N_6493);
or U7967 (N_7967,N_6698,N_6284);
xor U7968 (N_7968,N_6248,N_6813);
nand U7969 (N_7969,N_6880,N_6274);
or U7970 (N_7970,N_6258,N_6693);
nor U7971 (N_7971,N_6516,N_6772);
or U7972 (N_7972,N_6203,N_6141);
and U7973 (N_7973,N_6199,N_6961);
nor U7974 (N_7974,N_6751,N_6433);
and U7975 (N_7975,N_6340,N_6158);
xnor U7976 (N_7976,N_6081,N_6595);
and U7977 (N_7977,N_6344,N_6675);
xor U7978 (N_7978,N_6849,N_6872);
nand U7979 (N_7979,N_6141,N_6392);
xnor U7980 (N_7980,N_6877,N_6819);
nor U7981 (N_7981,N_6381,N_6165);
or U7982 (N_7982,N_6379,N_6326);
or U7983 (N_7983,N_6239,N_6460);
xor U7984 (N_7984,N_6293,N_6846);
nand U7985 (N_7985,N_6595,N_6146);
and U7986 (N_7986,N_6915,N_6627);
nor U7987 (N_7987,N_6831,N_6372);
and U7988 (N_7988,N_6970,N_6105);
or U7989 (N_7989,N_6791,N_6135);
xor U7990 (N_7990,N_6706,N_6575);
and U7991 (N_7991,N_6271,N_6276);
nor U7992 (N_7992,N_6158,N_6929);
nand U7993 (N_7993,N_6774,N_6468);
nor U7994 (N_7994,N_6833,N_6562);
and U7995 (N_7995,N_6392,N_6110);
or U7996 (N_7996,N_6218,N_6966);
xnor U7997 (N_7997,N_6607,N_6289);
nand U7998 (N_7998,N_6135,N_6161);
nand U7999 (N_7999,N_6720,N_6610);
or U8000 (N_8000,N_7882,N_7219);
nor U8001 (N_8001,N_7628,N_7213);
nand U8002 (N_8002,N_7360,N_7676);
nor U8003 (N_8003,N_7016,N_7320);
xor U8004 (N_8004,N_7431,N_7526);
and U8005 (N_8005,N_7761,N_7018);
xnor U8006 (N_8006,N_7606,N_7103);
xnor U8007 (N_8007,N_7138,N_7952);
xor U8008 (N_8008,N_7875,N_7074);
xnor U8009 (N_8009,N_7602,N_7895);
or U8010 (N_8010,N_7722,N_7383);
or U8011 (N_8011,N_7177,N_7989);
or U8012 (N_8012,N_7949,N_7100);
and U8013 (N_8013,N_7155,N_7239);
nor U8014 (N_8014,N_7935,N_7301);
nor U8015 (N_8015,N_7050,N_7559);
nor U8016 (N_8016,N_7695,N_7004);
nor U8017 (N_8017,N_7373,N_7113);
nor U8018 (N_8018,N_7342,N_7404);
and U8019 (N_8019,N_7820,N_7796);
or U8020 (N_8020,N_7554,N_7965);
nand U8021 (N_8021,N_7275,N_7290);
or U8022 (N_8022,N_7326,N_7394);
or U8023 (N_8023,N_7890,N_7261);
nor U8024 (N_8024,N_7444,N_7599);
and U8025 (N_8025,N_7906,N_7202);
or U8026 (N_8026,N_7334,N_7822);
or U8027 (N_8027,N_7963,N_7283);
nand U8028 (N_8028,N_7532,N_7309);
nand U8029 (N_8029,N_7666,N_7530);
and U8030 (N_8030,N_7964,N_7868);
xor U8031 (N_8031,N_7960,N_7860);
and U8032 (N_8032,N_7488,N_7355);
nor U8033 (N_8033,N_7499,N_7614);
xnor U8034 (N_8034,N_7075,N_7749);
or U8035 (N_8035,N_7214,N_7473);
and U8036 (N_8036,N_7484,N_7763);
or U8037 (N_8037,N_7696,N_7790);
or U8038 (N_8038,N_7068,N_7374);
or U8039 (N_8039,N_7748,N_7083);
nor U8040 (N_8040,N_7448,N_7516);
nand U8041 (N_8041,N_7311,N_7997);
or U8042 (N_8042,N_7914,N_7288);
xor U8043 (N_8043,N_7564,N_7338);
and U8044 (N_8044,N_7885,N_7998);
or U8045 (N_8045,N_7871,N_7001);
and U8046 (N_8046,N_7787,N_7793);
or U8047 (N_8047,N_7612,N_7151);
and U8048 (N_8048,N_7992,N_7923);
or U8049 (N_8049,N_7525,N_7318);
nor U8050 (N_8050,N_7678,N_7881);
xor U8051 (N_8051,N_7416,N_7289);
and U8052 (N_8052,N_7717,N_7101);
and U8053 (N_8053,N_7485,N_7972);
and U8054 (N_8054,N_7359,N_7609);
or U8055 (N_8055,N_7682,N_7683);
nor U8056 (N_8056,N_7037,N_7744);
nand U8057 (N_8057,N_7848,N_7560);
or U8058 (N_8058,N_7865,N_7105);
or U8059 (N_8059,N_7694,N_7370);
and U8060 (N_8060,N_7044,N_7066);
nand U8061 (N_8061,N_7421,N_7994);
or U8062 (N_8062,N_7082,N_7122);
nand U8063 (N_8063,N_7139,N_7794);
nand U8064 (N_8064,N_7310,N_7414);
xnor U8065 (N_8065,N_7322,N_7916);
nand U8066 (N_8066,N_7437,N_7670);
or U8067 (N_8067,N_7225,N_7231);
xor U8068 (N_8068,N_7474,N_7733);
nand U8069 (N_8069,N_7805,N_7115);
nor U8070 (N_8070,N_7624,N_7380);
nor U8071 (N_8071,N_7178,N_7942);
and U8072 (N_8072,N_7813,N_7157);
and U8073 (N_8073,N_7986,N_7999);
xor U8074 (N_8074,N_7331,N_7637);
and U8075 (N_8075,N_7280,N_7005);
and U8076 (N_8076,N_7106,N_7343);
or U8077 (N_8077,N_7714,N_7767);
xor U8078 (N_8078,N_7302,N_7097);
or U8079 (N_8079,N_7493,N_7323);
and U8080 (N_8080,N_7388,N_7503);
or U8081 (N_8081,N_7424,N_7956);
nor U8082 (N_8082,N_7366,N_7568);
nor U8083 (N_8083,N_7954,N_7142);
nand U8084 (N_8084,N_7240,N_7440);
nor U8085 (N_8085,N_7341,N_7687);
and U8086 (N_8086,N_7947,N_7596);
or U8087 (N_8087,N_7182,N_7642);
or U8088 (N_8088,N_7222,N_7212);
or U8089 (N_8089,N_7000,N_7060);
nor U8090 (N_8090,N_7974,N_7619);
and U8091 (N_8091,N_7762,N_7009);
or U8092 (N_8092,N_7154,N_7120);
nand U8093 (N_8093,N_7896,N_7041);
nand U8094 (N_8094,N_7920,N_7096);
nand U8095 (N_8095,N_7519,N_7766);
nor U8096 (N_8096,N_7109,N_7057);
or U8097 (N_8097,N_7521,N_7789);
xor U8098 (N_8098,N_7292,N_7938);
nand U8099 (N_8099,N_7317,N_7601);
nand U8100 (N_8100,N_7583,N_7738);
xor U8101 (N_8101,N_7033,N_7778);
or U8102 (N_8102,N_7128,N_7728);
xor U8103 (N_8103,N_7220,N_7582);
xor U8104 (N_8104,N_7853,N_7218);
and U8105 (N_8105,N_7736,N_7287);
nor U8106 (N_8106,N_7681,N_7897);
xnor U8107 (N_8107,N_7915,N_7078);
xnor U8108 (N_8108,N_7032,N_7726);
nor U8109 (N_8109,N_7467,N_7476);
and U8110 (N_8110,N_7648,N_7929);
or U8111 (N_8111,N_7752,N_7135);
and U8112 (N_8112,N_7464,N_7022);
nand U8113 (N_8113,N_7731,N_7818);
nand U8114 (N_8114,N_7544,N_7543);
or U8115 (N_8115,N_7863,N_7198);
nor U8116 (N_8116,N_7812,N_7760);
xor U8117 (N_8117,N_7775,N_7468);
and U8118 (N_8118,N_7158,N_7656);
xnor U8119 (N_8119,N_7659,N_7961);
xnor U8120 (N_8120,N_7828,N_7433);
xor U8121 (N_8121,N_7522,N_7884);
nand U8122 (N_8122,N_7449,N_7143);
xnor U8123 (N_8123,N_7831,N_7256);
nand U8124 (N_8124,N_7791,N_7422);
and U8125 (N_8125,N_7857,N_7201);
nor U8126 (N_8126,N_7644,N_7934);
or U8127 (N_8127,N_7056,N_7372);
and U8128 (N_8128,N_7176,N_7015);
or U8129 (N_8129,N_7846,N_7732);
xnor U8130 (N_8130,N_7181,N_7452);
or U8131 (N_8131,N_7786,N_7930);
and U8132 (N_8132,N_7730,N_7306);
xor U8133 (N_8133,N_7203,N_7608);
and U8134 (N_8134,N_7163,N_7455);
xnor U8135 (N_8135,N_7566,N_7149);
or U8136 (N_8136,N_7921,N_7709);
and U8137 (N_8137,N_7179,N_7579);
xnor U8138 (N_8138,N_7702,N_7506);
nor U8139 (N_8139,N_7209,N_7561);
xnor U8140 (N_8140,N_7210,N_7346);
nor U8141 (N_8141,N_7042,N_7299);
nand U8142 (N_8142,N_7169,N_7011);
nand U8143 (N_8143,N_7739,N_7990);
nor U8144 (N_8144,N_7396,N_7363);
or U8145 (N_8145,N_7505,N_7565);
nor U8146 (N_8146,N_7053,N_7824);
nand U8147 (N_8147,N_7536,N_7978);
or U8148 (N_8148,N_7278,N_7123);
and U8149 (N_8149,N_7577,N_7174);
or U8150 (N_8150,N_7393,N_7862);
xor U8151 (N_8151,N_7040,N_7887);
xor U8152 (N_8152,N_7065,N_7395);
xor U8153 (N_8153,N_7878,N_7495);
or U8154 (N_8154,N_7727,N_7325);
nor U8155 (N_8155,N_7540,N_7126);
nand U8156 (N_8156,N_7980,N_7773);
xor U8157 (N_8157,N_7038,N_7527);
nand U8158 (N_8158,N_7195,N_7783);
or U8159 (N_8159,N_7618,N_7447);
or U8160 (N_8160,N_7951,N_7321);
and U8161 (N_8161,N_7832,N_7651);
or U8162 (N_8162,N_7377,N_7185);
or U8163 (N_8163,N_7962,N_7697);
nand U8164 (N_8164,N_7852,N_7026);
and U8165 (N_8165,N_7246,N_7402);
nor U8166 (N_8166,N_7632,N_7171);
or U8167 (N_8167,N_7861,N_7047);
nor U8168 (N_8168,N_7470,N_7982);
and U8169 (N_8169,N_7584,N_7487);
nor U8170 (N_8170,N_7592,N_7392);
or U8171 (N_8171,N_7339,N_7785);
nor U8172 (N_8172,N_7248,N_7036);
nand U8173 (N_8173,N_7226,N_7273);
nor U8174 (N_8174,N_7084,N_7356);
nand U8175 (N_8175,N_7241,N_7556);
xnor U8176 (N_8176,N_7839,N_7234);
nand U8177 (N_8177,N_7755,N_7443);
nor U8178 (N_8178,N_7415,N_7093);
or U8179 (N_8179,N_7406,N_7446);
or U8180 (N_8180,N_7888,N_7967);
xnor U8181 (N_8181,N_7585,N_7953);
nor U8182 (N_8182,N_7684,N_7511);
nand U8183 (N_8183,N_7939,N_7586);
or U8184 (N_8184,N_7605,N_7199);
xnor U8185 (N_8185,N_7357,N_7686);
and U8186 (N_8186,N_7804,N_7173);
or U8187 (N_8187,N_7305,N_7673);
xnor U8188 (N_8188,N_7408,N_7847);
nor U8189 (N_8189,N_7389,N_7364);
nand U8190 (N_8190,N_7134,N_7611);
xnor U8191 (N_8191,N_7693,N_7379);
xnor U8192 (N_8192,N_7017,N_7335);
or U8193 (N_8193,N_7462,N_7502);
xor U8194 (N_8194,N_7640,N_7898);
nand U8195 (N_8195,N_7515,N_7269);
nor U8196 (N_8196,N_7698,N_7753);
nand U8197 (N_8197,N_7337,N_7734);
xnor U8198 (N_8198,N_7712,N_7039);
or U8199 (N_8199,N_7919,N_7286);
nor U8200 (N_8200,N_7948,N_7984);
or U8201 (N_8201,N_7855,N_7946);
or U8202 (N_8202,N_7168,N_7553);
and U8203 (N_8203,N_7837,N_7808);
nand U8204 (N_8204,N_7798,N_7966);
or U8205 (N_8205,N_7996,N_7977);
or U8206 (N_8206,N_7235,N_7578);
xor U8207 (N_8207,N_7551,N_7161);
xor U8208 (N_8208,N_7439,N_7943);
nand U8209 (N_8209,N_7641,N_7607);
nor U8210 (N_8210,N_7453,N_7080);
nor U8211 (N_8211,N_7192,N_7274);
nor U8212 (N_8212,N_7054,N_7740);
nor U8213 (N_8213,N_7587,N_7297);
nand U8214 (N_8214,N_7830,N_7533);
xnor U8215 (N_8215,N_7649,N_7501);
xnor U8216 (N_8216,N_7816,N_7397);
and U8217 (N_8217,N_7770,N_7588);
nor U8218 (N_8218,N_7165,N_7450);
nor U8219 (N_8219,N_7750,N_7531);
xnor U8220 (N_8220,N_7504,N_7597);
and U8221 (N_8221,N_7567,N_7489);
and U8222 (N_8222,N_7021,N_7757);
and U8223 (N_8223,N_7615,N_7430);
nor U8224 (N_8224,N_7627,N_7937);
nor U8225 (N_8225,N_7995,N_7076);
or U8226 (N_8226,N_7238,N_7023);
nand U8227 (N_8227,N_7051,N_7889);
xnor U8228 (N_8228,N_7549,N_7512);
nand U8229 (N_8229,N_7869,N_7340);
nand U8230 (N_8230,N_7912,N_7542);
or U8231 (N_8231,N_7405,N_7639);
and U8232 (N_8232,N_7482,N_7626);
and U8233 (N_8233,N_7369,N_7224);
xor U8234 (N_8234,N_7715,N_7569);
xnor U8235 (N_8235,N_7826,N_7719);
and U8236 (N_8236,N_7124,N_7441);
and U8237 (N_8237,N_7013,N_7620);
xor U8238 (N_8238,N_7249,N_7776);
nand U8239 (N_8239,N_7186,N_7206);
nor U8240 (N_8240,N_7293,N_7385);
and U8241 (N_8241,N_7253,N_7419);
nor U8242 (N_8242,N_7413,N_7085);
nand U8243 (N_8243,N_7107,N_7062);
xnor U8244 (N_8244,N_7900,N_7008);
xnor U8245 (N_8245,N_7067,N_7159);
nand U8246 (N_8246,N_7049,N_7228);
or U8247 (N_8247,N_7014,N_7130);
xor U8248 (N_8248,N_7811,N_7170);
nor U8249 (N_8249,N_7092,N_7539);
nor U8250 (N_8250,N_7745,N_7409);
xnor U8251 (N_8251,N_7002,N_7870);
or U8252 (N_8252,N_7070,N_7403);
xnor U8253 (N_8253,N_7211,N_7873);
nor U8254 (N_8254,N_7035,N_7891);
nor U8255 (N_8255,N_7230,N_7264);
and U8256 (N_8256,N_7555,N_7970);
nor U8257 (N_8257,N_7010,N_7007);
and U8258 (N_8258,N_7658,N_7490);
and U8259 (N_8259,N_7312,N_7491);
or U8260 (N_8260,N_7645,N_7707);
nor U8261 (N_8261,N_7932,N_7764);
nor U8262 (N_8262,N_7500,N_7316);
or U8263 (N_8263,N_7327,N_7110);
nand U8264 (N_8264,N_7469,N_7215);
and U8265 (N_8265,N_7072,N_7481);
nand U8266 (N_8266,N_7616,N_7460);
xor U8267 (N_8267,N_7432,N_7112);
nand U8268 (N_8268,N_7859,N_7237);
and U8269 (N_8269,N_7095,N_7513);
and U8270 (N_8270,N_7308,N_7933);
nor U8271 (N_8271,N_7164,N_7589);
xnor U8272 (N_8272,N_7271,N_7653);
nand U8273 (N_8273,N_7236,N_7457);
nand U8274 (N_8274,N_7417,N_7114);
or U8275 (N_8275,N_7438,N_7958);
and U8276 (N_8276,N_7917,N_7562);
nor U8277 (N_8277,N_7771,N_7375);
xor U8278 (N_8278,N_7807,N_7523);
xor U8279 (N_8279,N_7260,N_7840);
and U8280 (N_8280,N_7806,N_7418);
xnor U8281 (N_8281,N_7646,N_7675);
or U8282 (N_8282,N_7711,N_7756);
and U8283 (N_8283,N_7779,N_7133);
nand U8284 (N_8284,N_7610,N_7844);
or U8285 (N_8285,N_7028,N_7475);
nor U8286 (N_8286,N_7162,N_7205);
and U8287 (N_8287,N_7911,N_7672);
nand U8288 (N_8288,N_7188,N_7034);
and U8289 (N_8289,N_7196,N_7132);
xnor U8290 (N_8290,N_7747,N_7819);
nand U8291 (N_8291,N_7137,N_7077);
nand U8292 (N_8292,N_7924,N_7843);
or U8293 (N_8293,N_7483,N_7841);
xnor U8294 (N_8294,N_7183,N_7307);
nand U8295 (N_8295,N_7886,N_7091);
or U8296 (N_8296,N_7772,N_7314);
and U8297 (N_8297,N_7063,N_7630);
nor U8298 (N_8298,N_7572,N_7429);
and U8299 (N_8299,N_7621,N_7909);
xor U8300 (N_8300,N_7362,N_7631);
or U8301 (N_8301,N_7720,N_7242);
and U8302 (N_8302,N_7663,N_7398);
nand U8303 (N_8303,N_7765,N_7647);
nor U8304 (N_8304,N_7774,N_7742);
and U8305 (N_8305,N_7668,N_7378);
or U8306 (N_8306,N_7721,N_7250);
nor U8307 (N_8307,N_7976,N_7514);
xor U8308 (N_8308,N_7479,N_7466);
or U8309 (N_8309,N_7401,N_7823);
and U8310 (N_8310,N_7879,N_7581);
and U8311 (N_8311,N_7347,N_7634);
and U8312 (N_8312,N_7781,N_7679);
nor U8313 (N_8313,N_7486,N_7344);
nand U8314 (N_8314,N_7180,N_7061);
and U8315 (N_8315,N_7454,N_7800);
or U8316 (N_8316,N_7175,N_7425);
or U8317 (N_8317,N_7024,N_7907);
nor U8318 (N_8318,N_7427,N_7266);
nor U8319 (N_8319,N_7459,N_7754);
and U8320 (N_8320,N_7296,N_7144);
xnor U8321 (N_8321,N_7724,N_7116);
and U8322 (N_8322,N_7263,N_7277);
and U8323 (N_8323,N_7146,N_7059);
and U8324 (N_8324,N_7777,N_7703);
xnor U8325 (N_8325,N_7187,N_7633);
or U8326 (N_8326,N_7545,N_7494);
nor U8327 (N_8327,N_7193,N_7136);
nand U8328 (N_8328,N_7534,N_7892);
xnor U8329 (N_8329,N_7352,N_7129);
or U8330 (N_8330,N_7768,N_7104);
nor U8331 (N_8331,N_7908,N_7650);
and U8332 (N_8332,N_7876,N_7304);
nand U8333 (N_8333,N_7575,N_7971);
and U8334 (N_8334,N_7387,N_7046);
xor U8335 (N_8335,N_7548,N_7988);
nor U8336 (N_8336,N_7081,N_7901);
and U8337 (N_8337,N_7674,N_7160);
nand U8338 (N_8338,N_7905,N_7893);
nor U8339 (N_8339,N_7636,N_7737);
or U8340 (N_8340,N_7098,N_7625);
nand U8341 (N_8341,N_7243,N_7769);
nand U8342 (N_8342,N_7817,N_7524);
and U8343 (N_8343,N_7458,N_7945);
or U8344 (N_8344,N_7936,N_7156);
nor U8345 (N_8345,N_7167,N_7071);
and U8346 (N_8346,N_7692,N_7300);
and U8347 (N_8347,N_7877,N_7498);
and U8348 (N_8348,N_7247,N_7102);
xor U8349 (N_8349,N_7685,N_7677);
xor U8350 (N_8350,N_7968,N_7699);
and U8351 (N_8351,N_7461,N_7391);
and U8352 (N_8352,N_7617,N_7194);
xor U8353 (N_8353,N_7259,N_7850);
nor U8354 (N_8354,N_7603,N_7520);
xor U8355 (N_8355,N_7701,N_7244);
nand U8356 (N_8356,N_7838,N_7801);
nand U8357 (N_8357,N_7294,N_7279);
nand U8358 (N_8358,N_7073,N_7197);
nor U8359 (N_8359,N_7613,N_7983);
nor U8360 (N_8360,N_7079,N_7842);
xnor U8361 (N_8361,N_7223,N_7688);
or U8362 (N_8362,N_7351,N_7638);
or U8363 (N_8363,N_7189,N_7276);
nor U8364 (N_8364,N_7436,N_7281);
or U8365 (N_8365,N_7782,N_7029);
xnor U8366 (N_8366,N_7324,N_7570);
xnor U8367 (N_8367,N_7574,N_7622);
nor U8368 (N_8368,N_7814,N_7981);
nor U8369 (N_8369,N_7463,N_7797);
and U8370 (N_8370,N_7931,N_7810);
and U8371 (N_8371,N_7232,N_7282);
nor U8372 (N_8372,N_7492,N_7127);
nand U8373 (N_8373,N_7537,N_7552);
and U8374 (N_8374,N_7147,N_7880);
or U8375 (N_8375,N_7657,N_7099);
and U8376 (N_8376,N_7207,N_7904);
nand U8377 (N_8377,N_7845,N_7883);
nor U8378 (N_8378,N_7576,N_7445);
or U8379 (N_8379,N_7595,N_7780);
nand U8380 (N_8380,N_7557,N_7987);
nand U8381 (N_8381,N_7058,N_7086);
xnor U8382 (N_8382,N_7284,N_7689);
and U8383 (N_8383,N_7221,N_7623);
xor U8384 (N_8384,N_7200,N_7872);
xnor U8385 (N_8385,N_7940,N_7451);
xnor U8386 (N_8386,N_7119,N_7713);
or U8387 (N_8387,N_7979,N_7784);
or U8388 (N_8388,N_7407,N_7849);
or U8389 (N_8389,N_7866,N_7348);
xnor U8390 (N_8390,N_7710,N_7538);
and U8391 (N_8391,N_7153,N_7043);
nor U8392 (N_8392,N_7400,N_7048);
nor U8393 (N_8393,N_7517,N_7465);
or U8394 (N_8394,N_7131,N_7345);
and U8395 (N_8395,N_7216,N_7547);
or U8396 (N_8396,N_7354,N_7546);
nor U8397 (N_8397,N_7064,N_7166);
and U8398 (N_8398,N_7723,N_7252);
xnor U8399 (N_8399,N_7864,N_7145);
nor U8400 (N_8400,N_7204,N_7792);
nor U8401 (N_8401,N_7590,N_7172);
or U8402 (N_8402,N_7959,N_7652);
or U8403 (N_8403,N_7856,N_7012);
or U8404 (N_8404,N_7191,N_7361);
and U8405 (N_8405,N_7927,N_7227);
nor U8406 (N_8406,N_7903,N_7661);
and U8407 (N_8407,N_7108,N_7350);
nor U8408 (N_8408,N_7089,N_7148);
nand U8409 (N_8409,N_7125,N_7255);
or U8410 (N_8410,N_7315,N_7558);
nor U8411 (N_8411,N_7665,N_7654);
nor U8412 (N_8412,N_7518,N_7270);
xnor U8413 (N_8413,N_7117,N_7020);
nor U8414 (N_8414,N_7435,N_7836);
or U8415 (N_8415,N_7118,N_7591);
or U8416 (N_8416,N_7390,N_7550);
and U8417 (N_8417,N_7833,N_7141);
nand U8418 (N_8418,N_7941,N_7471);
xnor U8419 (N_8419,N_7088,N_7121);
and U8420 (N_8420,N_7718,N_7535);
or U8421 (N_8421,N_7208,N_7368);
and U8422 (N_8422,N_7851,N_7329);
xnor U8423 (N_8423,N_7478,N_7643);
nand U8424 (N_8424,N_7829,N_7975);
nand U8425 (N_8425,N_7969,N_7664);
xnor U8426 (N_8426,N_7496,N_7573);
nand U8427 (N_8427,N_7834,N_7291);
and U8428 (N_8428,N_7298,N_7867);
and U8429 (N_8429,N_7258,N_7031);
nand U8430 (N_8430,N_7245,N_7957);
nor U8431 (N_8431,N_7690,N_7708);
nand U8432 (N_8432,N_7328,N_7508);
nor U8433 (N_8433,N_7420,N_7358);
nand U8434 (N_8434,N_7019,N_7381);
xor U8435 (N_8435,N_7229,N_7815);
nor U8436 (N_8436,N_7365,N_7944);
nand U8437 (N_8437,N_7313,N_7257);
nor U8438 (N_8438,N_7854,N_7434);
and U8439 (N_8439,N_7926,N_7667);
nor U8440 (N_8440,N_7825,N_7874);
xor U8441 (N_8441,N_7598,N_7993);
nor U8442 (N_8442,N_7412,N_7426);
nand U8443 (N_8443,N_7376,N_7319);
xnor U8444 (N_8444,N_7423,N_7660);
or U8445 (N_8445,N_7442,N_7629);
nand U8446 (N_8446,N_7480,N_7330);
xor U8447 (N_8447,N_7991,N_7955);
nor U8448 (N_8448,N_7254,N_7111);
or U8449 (N_8449,N_7925,N_7827);
nor U8450 (N_8450,N_7265,N_7894);
and U8451 (N_8451,N_7580,N_7922);
and U8452 (N_8452,N_7382,N_7803);
or U8453 (N_8453,N_7006,N_7913);
nor U8454 (N_8454,N_7332,N_7386);
or U8455 (N_8455,N_7333,N_7217);
nor U8456 (N_8456,N_7563,N_7809);
xor U8457 (N_8457,N_7741,N_7593);
xnor U8458 (N_8458,N_7267,N_7662);
nor U8459 (N_8459,N_7353,N_7704);
nand U8460 (N_8460,N_7950,N_7090);
or U8461 (N_8461,N_7152,N_7410);
nand U8462 (N_8462,N_7509,N_7150);
xnor U8463 (N_8463,N_7528,N_7003);
nand U8464 (N_8464,N_7303,N_7902);
or U8465 (N_8465,N_7928,N_7262);
nand U8466 (N_8466,N_7428,N_7985);
and U8467 (N_8467,N_7716,N_7140);
or U8468 (N_8468,N_7973,N_7541);
nor U8469 (N_8469,N_7758,N_7069);
and U8470 (N_8470,N_7045,N_7529);
nor U8471 (N_8471,N_7604,N_7233);
nor U8472 (N_8472,N_7055,N_7705);
and U8473 (N_8473,N_7285,N_7295);
nor U8474 (N_8474,N_7384,N_7399);
nand U8475 (N_8475,N_7858,N_7743);
xnor U8476 (N_8476,N_7472,N_7510);
nand U8477 (N_8477,N_7635,N_7918);
or U8478 (N_8478,N_7087,N_7821);
or U8479 (N_8479,N_7251,N_7184);
nor U8480 (N_8480,N_7371,N_7746);
xnor U8481 (N_8481,N_7336,N_7751);
nor U8482 (N_8482,N_7706,N_7725);
and U8483 (N_8483,N_7349,N_7669);
or U8484 (N_8484,N_7030,N_7272);
xnor U8485 (N_8485,N_7899,N_7027);
xnor U8486 (N_8486,N_7759,N_7507);
and U8487 (N_8487,N_7671,N_7735);
nand U8488 (N_8488,N_7802,N_7456);
xor U8489 (N_8489,N_7795,N_7729);
xnor U8490 (N_8490,N_7052,N_7700);
nand U8491 (N_8491,N_7600,N_7788);
xor U8492 (N_8492,N_7571,N_7477);
xnor U8493 (N_8493,N_7411,N_7799);
xnor U8494 (N_8494,N_7025,N_7835);
xor U8495 (N_8495,N_7367,N_7691);
and U8496 (N_8496,N_7094,N_7910);
or U8497 (N_8497,N_7655,N_7497);
nand U8498 (N_8498,N_7190,N_7594);
xor U8499 (N_8499,N_7268,N_7680);
nand U8500 (N_8500,N_7142,N_7109);
or U8501 (N_8501,N_7810,N_7804);
nand U8502 (N_8502,N_7240,N_7643);
or U8503 (N_8503,N_7822,N_7303);
nor U8504 (N_8504,N_7626,N_7840);
nor U8505 (N_8505,N_7289,N_7622);
xor U8506 (N_8506,N_7453,N_7643);
nand U8507 (N_8507,N_7310,N_7585);
and U8508 (N_8508,N_7167,N_7795);
or U8509 (N_8509,N_7392,N_7799);
or U8510 (N_8510,N_7987,N_7270);
or U8511 (N_8511,N_7738,N_7500);
and U8512 (N_8512,N_7838,N_7764);
nor U8513 (N_8513,N_7745,N_7610);
and U8514 (N_8514,N_7378,N_7256);
or U8515 (N_8515,N_7173,N_7596);
and U8516 (N_8516,N_7067,N_7587);
or U8517 (N_8517,N_7437,N_7399);
nand U8518 (N_8518,N_7188,N_7356);
nor U8519 (N_8519,N_7052,N_7085);
nand U8520 (N_8520,N_7468,N_7373);
nor U8521 (N_8521,N_7785,N_7998);
nand U8522 (N_8522,N_7698,N_7215);
xnor U8523 (N_8523,N_7720,N_7849);
and U8524 (N_8524,N_7585,N_7333);
nand U8525 (N_8525,N_7574,N_7163);
nand U8526 (N_8526,N_7578,N_7049);
or U8527 (N_8527,N_7459,N_7606);
or U8528 (N_8528,N_7787,N_7070);
nand U8529 (N_8529,N_7999,N_7745);
and U8530 (N_8530,N_7228,N_7744);
nand U8531 (N_8531,N_7030,N_7596);
and U8532 (N_8532,N_7545,N_7158);
nor U8533 (N_8533,N_7659,N_7609);
nor U8534 (N_8534,N_7038,N_7851);
or U8535 (N_8535,N_7186,N_7383);
nand U8536 (N_8536,N_7275,N_7348);
or U8537 (N_8537,N_7528,N_7970);
nor U8538 (N_8538,N_7382,N_7968);
xnor U8539 (N_8539,N_7497,N_7153);
nand U8540 (N_8540,N_7484,N_7848);
nor U8541 (N_8541,N_7228,N_7714);
nor U8542 (N_8542,N_7773,N_7331);
nand U8543 (N_8543,N_7019,N_7286);
or U8544 (N_8544,N_7538,N_7758);
or U8545 (N_8545,N_7683,N_7101);
and U8546 (N_8546,N_7538,N_7556);
nand U8547 (N_8547,N_7785,N_7001);
nand U8548 (N_8548,N_7523,N_7501);
nor U8549 (N_8549,N_7727,N_7716);
or U8550 (N_8550,N_7224,N_7058);
and U8551 (N_8551,N_7271,N_7499);
xor U8552 (N_8552,N_7778,N_7747);
nand U8553 (N_8553,N_7988,N_7873);
or U8554 (N_8554,N_7177,N_7510);
nor U8555 (N_8555,N_7116,N_7653);
or U8556 (N_8556,N_7798,N_7350);
and U8557 (N_8557,N_7595,N_7821);
nor U8558 (N_8558,N_7551,N_7845);
nand U8559 (N_8559,N_7619,N_7652);
nor U8560 (N_8560,N_7978,N_7919);
xor U8561 (N_8561,N_7671,N_7715);
nand U8562 (N_8562,N_7377,N_7430);
nand U8563 (N_8563,N_7826,N_7604);
or U8564 (N_8564,N_7620,N_7584);
or U8565 (N_8565,N_7237,N_7416);
nor U8566 (N_8566,N_7486,N_7308);
xor U8567 (N_8567,N_7866,N_7285);
xnor U8568 (N_8568,N_7920,N_7892);
nand U8569 (N_8569,N_7867,N_7134);
xor U8570 (N_8570,N_7702,N_7076);
xnor U8571 (N_8571,N_7324,N_7832);
and U8572 (N_8572,N_7003,N_7847);
nor U8573 (N_8573,N_7928,N_7884);
nand U8574 (N_8574,N_7900,N_7189);
or U8575 (N_8575,N_7380,N_7004);
xnor U8576 (N_8576,N_7483,N_7832);
nand U8577 (N_8577,N_7201,N_7229);
xor U8578 (N_8578,N_7471,N_7014);
nand U8579 (N_8579,N_7796,N_7478);
xor U8580 (N_8580,N_7695,N_7751);
xor U8581 (N_8581,N_7806,N_7814);
nand U8582 (N_8582,N_7646,N_7659);
nor U8583 (N_8583,N_7305,N_7711);
nand U8584 (N_8584,N_7844,N_7701);
xnor U8585 (N_8585,N_7491,N_7903);
or U8586 (N_8586,N_7486,N_7004);
xnor U8587 (N_8587,N_7715,N_7066);
xnor U8588 (N_8588,N_7274,N_7901);
xor U8589 (N_8589,N_7353,N_7437);
nor U8590 (N_8590,N_7456,N_7005);
and U8591 (N_8591,N_7372,N_7416);
xor U8592 (N_8592,N_7291,N_7884);
and U8593 (N_8593,N_7085,N_7640);
and U8594 (N_8594,N_7227,N_7967);
and U8595 (N_8595,N_7500,N_7765);
nor U8596 (N_8596,N_7418,N_7336);
or U8597 (N_8597,N_7664,N_7320);
nor U8598 (N_8598,N_7509,N_7805);
nor U8599 (N_8599,N_7028,N_7819);
xnor U8600 (N_8600,N_7563,N_7804);
or U8601 (N_8601,N_7388,N_7825);
nor U8602 (N_8602,N_7133,N_7626);
and U8603 (N_8603,N_7589,N_7521);
or U8604 (N_8604,N_7431,N_7713);
xor U8605 (N_8605,N_7188,N_7442);
nor U8606 (N_8606,N_7199,N_7847);
or U8607 (N_8607,N_7869,N_7822);
xor U8608 (N_8608,N_7585,N_7358);
nand U8609 (N_8609,N_7214,N_7376);
and U8610 (N_8610,N_7244,N_7312);
and U8611 (N_8611,N_7397,N_7369);
nand U8612 (N_8612,N_7364,N_7712);
and U8613 (N_8613,N_7558,N_7904);
nor U8614 (N_8614,N_7358,N_7537);
xnor U8615 (N_8615,N_7251,N_7012);
nand U8616 (N_8616,N_7505,N_7557);
nor U8617 (N_8617,N_7388,N_7614);
nor U8618 (N_8618,N_7073,N_7920);
and U8619 (N_8619,N_7515,N_7955);
and U8620 (N_8620,N_7502,N_7973);
nor U8621 (N_8621,N_7599,N_7553);
nand U8622 (N_8622,N_7659,N_7592);
nor U8623 (N_8623,N_7133,N_7914);
nand U8624 (N_8624,N_7646,N_7848);
or U8625 (N_8625,N_7387,N_7267);
xor U8626 (N_8626,N_7912,N_7854);
or U8627 (N_8627,N_7026,N_7435);
or U8628 (N_8628,N_7023,N_7559);
nand U8629 (N_8629,N_7245,N_7461);
or U8630 (N_8630,N_7874,N_7849);
nand U8631 (N_8631,N_7301,N_7308);
nor U8632 (N_8632,N_7830,N_7410);
or U8633 (N_8633,N_7717,N_7592);
xnor U8634 (N_8634,N_7600,N_7649);
nor U8635 (N_8635,N_7858,N_7496);
nand U8636 (N_8636,N_7537,N_7357);
and U8637 (N_8637,N_7536,N_7060);
xor U8638 (N_8638,N_7638,N_7175);
nand U8639 (N_8639,N_7427,N_7654);
and U8640 (N_8640,N_7585,N_7779);
and U8641 (N_8641,N_7107,N_7164);
and U8642 (N_8642,N_7919,N_7441);
or U8643 (N_8643,N_7870,N_7050);
and U8644 (N_8644,N_7067,N_7725);
or U8645 (N_8645,N_7648,N_7201);
and U8646 (N_8646,N_7879,N_7014);
and U8647 (N_8647,N_7329,N_7688);
xnor U8648 (N_8648,N_7816,N_7953);
nand U8649 (N_8649,N_7515,N_7222);
nand U8650 (N_8650,N_7334,N_7637);
nor U8651 (N_8651,N_7684,N_7033);
or U8652 (N_8652,N_7903,N_7312);
and U8653 (N_8653,N_7615,N_7109);
xnor U8654 (N_8654,N_7037,N_7261);
nor U8655 (N_8655,N_7274,N_7308);
nand U8656 (N_8656,N_7187,N_7018);
nor U8657 (N_8657,N_7130,N_7941);
nor U8658 (N_8658,N_7680,N_7590);
nand U8659 (N_8659,N_7914,N_7099);
nand U8660 (N_8660,N_7810,N_7414);
xnor U8661 (N_8661,N_7101,N_7090);
and U8662 (N_8662,N_7198,N_7314);
xnor U8663 (N_8663,N_7164,N_7476);
or U8664 (N_8664,N_7677,N_7630);
nand U8665 (N_8665,N_7906,N_7703);
and U8666 (N_8666,N_7569,N_7871);
or U8667 (N_8667,N_7440,N_7672);
or U8668 (N_8668,N_7770,N_7391);
and U8669 (N_8669,N_7657,N_7385);
nor U8670 (N_8670,N_7150,N_7958);
and U8671 (N_8671,N_7398,N_7626);
nand U8672 (N_8672,N_7356,N_7012);
nor U8673 (N_8673,N_7468,N_7357);
or U8674 (N_8674,N_7513,N_7012);
and U8675 (N_8675,N_7515,N_7778);
nand U8676 (N_8676,N_7489,N_7160);
or U8677 (N_8677,N_7888,N_7575);
and U8678 (N_8678,N_7416,N_7515);
and U8679 (N_8679,N_7551,N_7273);
nor U8680 (N_8680,N_7898,N_7317);
or U8681 (N_8681,N_7145,N_7733);
or U8682 (N_8682,N_7511,N_7523);
nand U8683 (N_8683,N_7920,N_7702);
or U8684 (N_8684,N_7953,N_7401);
xnor U8685 (N_8685,N_7764,N_7228);
and U8686 (N_8686,N_7432,N_7631);
and U8687 (N_8687,N_7422,N_7116);
and U8688 (N_8688,N_7317,N_7353);
xnor U8689 (N_8689,N_7841,N_7633);
xnor U8690 (N_8690,N_7780,N_7168);
xnor U8691 (N_8691,N_7741,N_7400);
and U8692 (N_8692,N_7597,N_7056);
or U8693 (N_8693,N_7425,N_7825);
nand U8694 (N_8694,N_7448,N_7344);
nand U8695 (N_8695,N_7279,N_7008);
or U8696 (N_8696,N_7569,N_7832);
xnor U8697 (N_8697,N_7340,N_7387);
nand U8698 (N_8698,N_7821,N_7376);
nand U8699 (N_8699,N_7367,N_7704);
or U8700 (N_8700,N_7012,N_7900);
nand U8701 (N_8701,N_7862,N_7758);
and U8702 (N_8702,N_7781,N_7376);
nand U8703 (N_8703,N_7433,N_7889);
xnor U8704 (N_8704,N_7870,N_7898);
nor U8705 (N_8705,N_7250,N_7665);
xor U8706 (N_8706,N_7833,N_7548);
nand U8707 (N_8707,N_7621,N_7205);
or U8708 (N_8708,N_7500,N_7574);
nor U8709 (N_8709,N_7979,N_7925);
nor U8710 (N_8710,N_7636,N_7137);
and U8711 (N_8711,N_7492,N_7170);
and U8712 (N_8712,N_7843,N_7447);
nor U8713 (N_8713,N_7543,N_7763);
nor U8714 (N_8714,N_7640,N_7926);
nor U8715 (N_8715,N_7665,N_7388);
or U8716 (N_8716,N_7447,N_7331);
xnor U8717 (N_8717,N_7041,N_7788);
and U8718 (N_8718,N_7483,N_7182);
nand U8719 (N_8719,N_7783,N_7265);
xor U8720 (N_8720,N_7851,N_7559);
or U8721 (N_8721,N_7287,N_7048);
or U8722 (N_8722,N_7773,N_7505);
or U8723 (N_8723,N_7014,N_7221);
nand U8724 (N_8724,N_7556,N_7901);
or U8725 (N_8725,N_7941,N_7886);
and U8726 (N_8726,N_7680,N_7273);
nor U8727 (N_8727,N_7409,N_7337);
nor U8728 (N_8728,N_7660,N_7198);
or U8729 (N_8729,N_7608,N_7235);
nand U8730 (N_8730,N_7877,N_7266);
nor U8731 (N_8731,N_7628,N_7425);
or U8732 (N_8732,N_7375,N_7570);
and U8733 (N_8733,N_7117,N_7462);
or U8734 (N_8734,N_7311,N_7990);
nor U8735 (N_8735,N_7225,N_7420);
nor U8736 (N_8736,N_7982,N_7489);
nor U8737 (N_8737,N_7403,N_7059);
nand U8738 (N_8738,N_7331,N_7839);
nand U8739 (N_8739,N_7752,N_7722);
nor U8740 (N_8740,N_7067,N_7265);
nor U8741 (N_8741,N_7257,N_7933);
or U8742 (N_8742,N_7283,N_7718);
or U8743 (N_8743,N_7823,N_7648);
nand U8744 (N_8744,N_7610,N_7765);
xor U8745 (N_8745,N_7476,N_7511);
nand U8746 (N_8746,N_7473,N_7319);
or U8747 (N_8747,N_7455,N_7562);
and U8748 (N_8748,N_7077,N_7279);
xnor U8749 (N_8749,N_7283,N_7011);
or U8750 (N_8750,N_7327,N_7832);
and U8751 (N_8751,N_7957,N_7345);
nor U8752 (N_8752,N_7578,N_7447);
nand U8753 (N_8753,N_7299,N_7948);
and U8754 (N_8754,N_7968,N_7470);
xnor U8755 (N_8755,N_7873,N_7441);
and U8756 (N_8756,N_7816,N_7970);
xnor U8757 (N_8757,N_7220,N_7991);
and U8758 (N_8758,N_7924,N_7712);
nor U8759 (N_8759,N_7848,N_7977);
or U8760 (N_8760,N_7596,N_7921);
xnor U8761 (N_8761,N_7267,N_7901);
xor U8762 (N_8762,N_7818,N_7938);
nor U8763 (N_8763,N_7870,N_7618);
xnor U8764 (N_8764,N_7704,N_7858);
and U8765 (N_8765,N_7649,N_7219);
and U8766 (N_8766,N_7971,N_7959);
xor U8767 (N_8767,N_7053,N_7401);
nand U8768 (N_8768,N_7556,N_7881);
or U8769 (N_8769,N_7226,N_7120);
or U8770 (N_8770,N_7432,N_7650);
or U8771 (N_8771,N_7963,N_7091);
and U8772 (N_8772,N_7413,N_7744);
and U8773 (N_8773,N_7715,N_7028);
or U8774 (N_8774,N_7681,N_7850);
and U8775 (N_8775,N_7975,N_7854);
and U8776 (N_8776,N_7683,N_7605);
or U8777 (N_8777,N_7004,N_7787);
nor U8778 (N_8778,N_7268,N_7678);
and U8779 (N_8779,N_7943,N_7029);
and U8780 (N_8780,N_7557,N_7370);
nand U8781 (N_8781,N_7684,N_7433);
nand U8782 (N_8782,N_7607,N_7782);
nor U8783 (N_8783,N_7027,N_7513);
and U8784 (N_8784,N_7705,N_7317);
nor U8785 (N_8785,N_7727,N_7829);
nor U8786 (N_8786,N_7448,N_7686);
nand U8787 (N_8787,N_7282,N_7974);
nand U8788 (N_8788,N_7487,N_7678);
and U8789 (N_8789,N_7700,N_7372);
nor U8790 (N_8790,N_7611,N_7164);
xnor U8791 (N_8791,N_7060,N_7750);
and U8792 (N_8792,N_7619,N_7395);
nor U8793 (N_8793,N_7530,N_7114);
xnor U8794 (N_8794,N_7714,N_7061);
nand U8795 (N_8795,N_7238,N_7263);
and U8796 (N_8796,N_7945,N_7629);
nand U8797 (N_8797,N_7498,N_7241);
xor U8798 (N_8798,N_7808,N_7707);
nand U8799 (N_8799,N_7853,N_7201);
nand U8800 (N_8800,N_7151,N_7024);
nand U8801 (N_8801,N_7906,N_7002);
and U8802 (N_8802,N_7543,N_7922);
nand U8803 (N_8803,N_7723,N_7186);
xor U8804 (N_8804,N_7879,N_7276);
nand U8805 (N_8805,N_7798,N_7080);
nand U8806 (N_8806,N_7000,N_7034);
nor U8807 (N_8807,N_7229,N_7848);
nand U8808 (N_8808,N_7413,N_7736);
xor U8809 (N_8809,N_7495,N_7928);
nor U8810 (N_8810,N_7065,N_7168);
or U8811 (N_8811,N_7114,N_7162);
or U8812 (N_8812,N_7780,N_7745);
nor U8813 (N_8813,N_7316,N_7911);
xor U8814 (N_8814,N_7286,N_7225);
and U8815 (N_8815,N_7507,N_7983);
nand U8816 (N_8816,N_7454,N_7896);
and U8817 (N_8817,N_7079,N_7966);
or U8818 (N_8818,N_7221,N_7681);
and U8819 (N_8819,N_7918,N_7288);
nand U8820 (N_8820,N_7463,N_7483);
nand U8821 (N_8821,N_7386,N_7873);
nand U8822 (N_8822,N_7388,N_7481);
and U8823 (N_8823,N_7668,N_7376);
or U8824 (N_8824,N_7756,N_7576);
nor U8825 (N_8825,N_7307,N_7322);
and U8826 (N_8826,N_7745,N_7643);
nor U8827 (N_8827,N_7052,N_7060);
or U8828 (N_8828,N_7219,N_7701);
xnor U8829 (N_8829,N_7888,N_7710);
nor U8830 (N_8830,N_7990,N_7551);
nor U8831 (N_8831,N_7977,N_7884);
nand U8832 (N_8832,N_7615,N_7344);
xor U8833 (N_8833,N_7392,N_7866);
xnor U8834 (N_8834,N_7227,N_7717);
nor U8835 (N_8835,N_7443,N_7520);
nor U8836 (N_8836,N_7538,N_7764);
or U8837 (N_8837,N_7182,N_7761);
and U8838 (N_8838,N_7116,N_7250);
xnor U8839 (N_8839,N_7415,N_7430);
nand U8840 (N_8840,N_7671,N_7860);
and U8841 (N_8841,N_7651,N_7992);
nand U8842 (N_8842,N_7969,N_7275);
or U8843 (N_8843,N_7346,N_7318);
nor U8844 (N_8844,N_7168,N_7486);
and U8845 (N_8845,N_7973,N_7988);
xor U8846 (N_8846,N_7058,N_7685);
nand U8847 (N_8847,N_7211,N_7848);
nand U8848 (N_8848,N_7851,N_7541);
nor U8849 (N_8849,N_7052,N_7807);
or U8850 (N_8850,N_7904,N_7419);
or U8851 (N_8851,N_7796,N_7266);
nor U8852 (N_8852,N_7512,N_7878);
xor U8853 (N_8853,N_7988,N_7288);
nor U8854 (N_8854,N_7794,N_7731);
nand U8855 (N_8855,N_7306,N_7516);
xnor U8856 (N_8856,N_7209,N_7368);
and U8857 (N_8857,N_7927,N_7946);
nor U8858 (N_8858,N_7980,N_7770);
or U8859 (N_8859,N_7875,N_7689);
xnor U8860 (N_8860,N_7832,N_7492);
and U8861 (N_8861,N_7718,N_7372);
and U8862 (N_8862,N_7045,N_7363);
nor U8863 (N_8863,N_7909,N_7565);
nand U8864 (N_8864,N_7419,N_7916);
xor U8865 (N_8865,N_7666,N_7548);
nor U8866 (N_8866,N_7914,N_7059);
nand U8867 (N_8867,N_7757,N_7289);
and U8868 (N_8868,N_7489,N_7056);
xnor U8869 (N_8869,N_7421,N_7162);
or U8870 (N_8870,N_7688,N_7313);
xnor U8871 (N_8871,N_7288,N_7098);
nand U8872 (N_8872,N_7008,N_7213);
xnor U8873 (N_8873,N_7199,N_7506);
nor U8874 (N_8874,N_7787,N_7894);
nand U8875 (N_8875,N_7139,N_7297);
nand U8876 (N_8876,N_7422,N_7674);
nand U8877 (N_8877,N_7625,N_7156);
or U8878 (N_8878,N_7396,N_7311);
or U8879 (N_8879,N_7105,N_7035);
or U8880 (N_8880,N_7536,N_7595);
nor U8881 (N_8881,N_7406,N_7388);
nor U8882 (N_8882,N_7960,N_7343);
and U8883 (N_8883,N_7596,N_7857);
xnor U8884 (N_8884,N_7826,N_7035);
or U8885 (N_8885,N_7663,N_7816);
nor U8886 (N_8886,N_7298,N_7286);
nor U8887 (N_8887,N_7254,N_7977);
nand U8888 (N_8888,N_7624,N_7012);
or U8889 (N_8889,N_7398,N_7327);
nand U8890 (N_8890,N_7403,N_7967);
nand U8891 (N_8891,N_7245,N_7335);
xnor U8892 (N_8892,N_7008,N_7456);
xnor U8893 (N_8893,N_7156,N_7553);
nand U8894 (N_8894,N_7791,N_7902);
or U8895 (N_8895,N_7044,N_7446);
nor U8896 (N_8896,N_7060,N_7858);
xor U8897 (N_8897,N_7656,N_7187);
nand U8898 (N_8898,N_7187,N_7322);
and U8899 (N_8899,N_7961,N_7208);
nor U8900 (N_8900,N_7438,N_7546);
and U8901 (N_8901,N_7474,N_7459);
nor U8902 (N_8902,N_7484,N_7834);
nor U8903 (N_8903,N_7442,N_7146);
xnor U8904 (N_8904,N_7393,N_7903);
xnor U8905 (N_8905,N_7044,N_7489);
nand U8906 (N_8906,N_7572,N_7786);
or U8907 (N_8907,N_7580,N_7192);
and U8908 (N_8908,N_7001,N_7180);
xor U8909 (N_8909,N_7089,N_7375);
xor U8910 (N_8910,N_7310,N_7778);
xor U8911 (N_8911,N_7698,N_7154);
nor U8912 (N_8912,N_7282,N_7756);
xnor U8913 (N_8913,N_7033,N_7209);
or U8914 (N_8914,N_7698,N_7584);
nor U8915 (N_8915,N_7352,N_7219);
or U8916 (N_8916,N_7683,N_7806);
or U8917 (N_8917,N_7317,N_7316);
nor U8918 (N_8918,N_7069,N_7862);
nor U8919 (N_8919,N_7363,N_7546);
nand U8920 (N_8920,N_7406,N_7156);
nand U8921 (N_8921,N_7123,N_7552);
nor U8922 (N_8922,N_7212,N_7323);
xnor U8923 (N_8923,N_7129,N_7972);
and U8924 (N_8924,N_7719,N_7530);
xnor U8925 (N_8925,N_7910,N_7542);
or U8926 (N_8926,N_7886,N_7631);
or U8927 (N_8927,N_7262,N_7507);
nor U8928 (N_8928,N_7691,N_7281);
nor U8929 (N_8929,N_7834,N_7873);
or U8930 (N_8930,N_7653,N_7006);
xnor U8931 (N_8931,N_7146,N_7591);
nand U8932 (N_8932,N_7835,N_7472);
nor U8933 (N_8933,N_7600,N_7331);
and U8934 (N_8934,N_7788,N_7724);
nor U8935 (N_8935,N_7515,N_7807);
and U8936 (N_8936,N_7524,N_7006);
nor U8937 (N_8937,N_7137,N_7646);
nor U8938 (N_8938,N_7433,N_7940);
and U8939 (N_8939,N_7903,N_7706);
and U8940 (N_8940,N_7700,N_7046);
or U8941 (N_8941,N_7158,N_7262);
nor U8942 (N_8942,N_7283,N_7018);
and U8943 (N_8943,N_7404,N_7118);
or U8944 (N_8944,N_7298,N_7909);
nor U8945 (N_8945,N_7462,N_7967);
nor U8946 (N_8946,N_7994,N_7143);
or U8947 (N_8947,N_7226,N_7619);
nand U8948 (N_8948,N_7823,N_7940);
nor U8949 (N_8949,N_7413,N_7049);
nor U8950 (N_8950,N_7206,N_7272);
or U8951 (N_8951,N_7043,N_7897);
xnor U8952 (N_8952,N_7730,N_7971);
or U8953 (N_8953,N_7358,N_7831);
nor U8954 (N_8954,N_7435,N_7983);
and U8955 (N_8955,N_7027,N_7920);
nand U8956 (N_8956,N_7277,N_7766);
and U8957 (N_8957,N_7961,N_7343);
nand U8958 (N_8958,N_7103,N_7497);
nand U8959 (N_8959,N_7758,N_7297);
nand U8960 (N_8960,N_7110,N_7465);
nand U8961 (N_8961,N_7883,N_7212);
nor U8962 (N_8962,N_7806,N_7735);
or U8963 (N_8963,N_7978,N_7516);
and U8964 (N_8964,N_7624,N_7171);
nand U8965 (N_8965,N_7947,N_7967);
and U8966 (N_8966,N_7984,N_7519);
nor U8967 (N_8967,N_7105,N_7942);
or U8968 (N_8968,N_7135,N_7081);
xnor U8969 (N_8969,N_7710,N_7024);
and U8970 (N_8970,N_7225,N_7169);
xnor U8971 (N_8971,N_7686,N_7965);
nand U8972 (N_8972,N_7500,N_7914);
xnor U8973 (N_8973,N_7316,N_7006);
xnor U8974 (N_8974,N_7846,N_7907);
and U8975 (N_8975,N_7841,N_7728);
nor U8976 (N_8976,N_7857,N_7329);
and U8977 (N_8977,N_7501,N_7598);
and U8978 (N_8978,N_7578,N_7066);
and U8979 (N_8979,N_7267,N_7532);
xor U8980 (N_8980,N_7937,N_7740);
or U8981 (N_8981,N_7999,N_7661);
nor U8982 (N_8982,N_7626,N_7269);
and U8983 (N_8983,N_7305,N_7057);
and U8984 (N_8984,N_7381,N_7815);
xnor U8985 (N_8985,N_7935,N_7592);
or U8986 (N_8986,N_7498,N_7000);
nand U8987 (N_8987,N_7124,N_7554);
or U8988 (N_8988,N_7000,N_7642);
nor U8989 (N_8989,N_7759,N_7287);
xor U8990 (N_8990,N_7122,N_7193);
nand U8991 (N_8991,N_7701,N_7422);
xor U8992 (N_8992,N_7022,N_7662);
nor U8993 (N_8993,N_7763,N_7806);
xor U8994 (N_8994,N_7973,N_7376);
nand U8995 (N_8995,N_7812,N_7938);
or U8996 (N_8996,N_7954,N_7258);
and U8997 (N_8997,N_7809,N_7438);
or U8998 (N_8998,N_7666,N_7795);
nor U8999 (N_8999,N_7679,N_7333);
or U9000 (N_9000,N_8111,N_8504);
or U9001 (N_9001,N_8522,N_8584);
or U9002 (N_9002,N_8649,N_8748);
nor U9003 (N_9003,N_8172,N_8755);
nand U9004 (N_9004,N_8356,N_8531);
xnor U9005 (N_9005,N_8407,N_8656);
xnor U9006 (N_9006,N_8447,N_8057);
xor U9007 (N_9007,N_8323,N_8231);
xor U9008 (N_9008,N_8920,N_8510);
or U9009 (N_9009,N_8648,N_8156);
or U9010 (N_9010,N_8265,N_8007);
xor U9011 (N_9011,N_8972,N_8024);
or U9012 (N_9012,N_8069,N_8072);
nand U9013 (N_9013,N_8178,N_8555);
nand U9014 (N_9014,N_8880,N_8318);
nand U9015 (N_9015,N_8672,N_8805);
and U9016 (N_9016,N_8518,N_8740);
nand U9017 (N_9017,N_8556,N_8736);
and U9018 (N_9018,N_8128,N_8728);
and U9019 (N_9019,N_8278,N_8257);
nand U9020 (N_9020,N_8874,N_8227);
or U9021 (N_9021,N_8962,N_8803);
and U9022 (N_9022,N_8126,N_8075);
xnor U9023 (N_9023,N_8300,N_8897);
nand U9024 (N_9024,N_8939,N_8524);
nor U9025 (N_9025,N_8485,N_8664);
nor U9026 (N_9026,N_8366,N_8306);
or U9027 (N_9027,N_8309,N_8009);
nor U9028 (N_9028,N_8663,N_8638);
xnor U9029 (N_9029,N_8989,N_8229);
nand U9030 (N_9030,N_8208,N_8877);
or U9031 (N_9031,N_8254,N_8434);
nand U9032 (N_9032,N_8222,N_8351);
nor U9033 (N_9033,N_8170,N_8662);
nand U9034 (N_9034,N_8466,N_8583);
and U9035 (N_9035,N_8054,N_8947);
nand U9036 (N_9036,N_8490,N_8324);
nand U9037 (N_9037,N_8396,N_8281);
xnor U9038 (N_9038,N_8945,N_8688);
nor U9039 (N_9039,N_8997,N_8986);
nor U9040 (N_9040,N_8596,N_8418);
nor U9041 (N_9041,N_8620,N_8034);
nor U9042 (N_9042,N_8330,N_8012);
nor U9043 (N_9043,N_8669,N_8046);
nand U9044 (N_9044,N_8767,N_8798);
nand U9045 (N_9045,N_8785,N_8275);
and U9046 (N_9046,N_8599,N_8980);
or U9047 (N_9047,N_8965,N_8283);
and U9048 (N_9048,N_8975,N_8601);
or U9049 (N_9049,N_8383,N_8723);
nor U9050 (N_9050,N_8180,N_8209);
or U9051 (N_9051,N_8154,N_8704);
or U9052 (N_9052,N_8692,N_8978);
xor U9053 (N_9053,N_8566,N_8731);
nand U9054 (N_9054,N_8863,N_8889);
nor U9055 (N_9055,N_8987,N_8276);
or U9056 (N_9056,N_8578,N_8191);
xor U9057 (N_9057,N_8941,N_8218);
and U9058 (N_9058,N_8899,N_8368);
and U9059 (N_9059,N_8876,N_8480);
nand U9060 (N_9060,N_8791,N_8135);
nand U9061 (N_9061,N_8190,N_8515);
or U9062 (N_9062,N_8977,N_8701);
xor U9063 (N_9063,N_8613,N_8652);
or U9064 (N_9064,N_8326,N_8822);
nand U9065 (N_9065,N_8859,N_8217);
or U9066 (N_9066,N_8079,N_8832);
or U9067 (N_9067,N_8725,N_8151);
nor U9068 (N_9068,N_8677,N_8412);
nor U9069 (N_9069,N_8460,N_8352);
or U9070 (N_9070,N_8838,N_8763);
xnor U9071 (N_9071,N_8471,N_8262);
nand U9072 (N_9072,N_8760,N_8197);
nor U9073 (N_9073,N_8818,N_8703);
or U9074 (N_9074,N_8623,N_8194);
nor U9075 (N_9075,N_8056,N_8631);
nand U9076 (N_9076,N_8006,N_8847);
and U9077 (N_9077,N_8630,N_8071);
nand U9078 (N_9078,N_8973,N_8014);
or U9079 (N_9079,N_8269,N_8158);
or U9080 (N_9080,N_8633,N_8001);
or U9081 (N_9081,N_8761,N_8298);
or U9082 (N_9082,N_8038,N_8572);
and U9083 (N_9083,N_8523,N_8674);
xnor U9084 (N_9084,N_8509,N_8552);
or U9085 (N_9085,N_8422,N_8495);
or U9086 (N_9086,N_8077,N_8095);
xnor U9087 (N_9087,N_8346,N_8427);
nor U9088 (N_9088,N_8195,N_8313);
or U9089 (N_9089,N_8867,N_8308);
nor U9090 (N_9090,N_8148,N_8240);
and U9091 (N_9091,N_8726,N_8105);
and U9092 (N_9092,N_8602,N_8340);
nand U9093 (N_9093,N_8117,N_8409);
nor U9094 (N_9094,N_8234,N_8086);
nor U9095 (N_9095,N_8942,N_8350);
nand U9096 (N_9096,N_8319,N_8051);
nor U9097 (N_9097,N_8931,N_8990);
nor U9098 (N_9098,N_8499,N_8906);
nand U9099 (N_9099,N_8587,N_8059);
or U9100 (N_9100,N_8114,N_8280);
or U9101 (N_9101,N_8415,N_8104);
xnor U9102 (N_9102,N_8616,N_8253);
xor U9103 (N_9103,N_8406,N_8629);
xnor U9104 (N_9104,N_8563,N_8640);
or U9105 (N_9105,N_8299,N_8919);
or U9106 (N_9106,N_8909,N_8457);
and U9107 (N_9107,N_8689,N_8750);
and U9108 (N_9108,N_8696,N_8933);
nor U9109 (N_9109,N_8203,N_8712);
nand U9110 (N_9110,N_8944,N_8545);
or U9111 (N_9111,N_8643,N_8905);
xnor U9112 (N_9112,N_8093,N_8532);
xnor U9113 (N_9113,N_8835,N_8174);
xnor U9114 (N_9114,N_8302,N_8938);
or U9115 (N_9115,N_8742,N_8186);
xor U9116 (N_9116,N_8873,N_8053);
or U9117 (N_9117,N_8327,N_8903);
nor U9118 (N_9118,N_8949,N_8547);
nand U9119 (N_9119,N_8403,N_8379);
nor U9120 (N_9120,N_8013,N_8296);
xor U9121 (N_9121,N_8088,N_8772);
xor U9122 (N_9122,N_8301,N_8746);
nand U9123 (N_9123,N_8168,N_8559);
and U9124 (N_9124,N_8142,N_8189);
and U9125 (N_9125,N_8236,N_8834);
and U9126 (N_9126,N_8811,N_8147);
xnor U9127 (N_9127,N_8162,N_8985);
nor U9128 (N_9128,N_8573,N_8252);
xor U9129 (N_9129,N_8094,N_8386);
nand U9130 (N_9130,N_8400,N_8045);
nor U9131 (N_9131,N_8448,N_8771);
nor U9132 (N_9132,N_8605,N_8914);
and U9133 (N_9133,N_8829,N_8310);
nor U9134 (N_9134,N_8816,N_8894);
xor U9135 (N_9135,N_8442,N_8389);
and U9136 (N_9136,N_8844,N_8597);
nor U9137 (N_9137,N_8200,N_8198);
nor U9138 (N_9138,N_8388,N_8565);
xnor U9139 (N_9139,N_8924,N_8118);
xnor U9140 (N_9140,N_8347,N_8426);
nor U9141 (N_9141,N_8710,N_8671);
nor U9142 (N_9142,N_8372,N_8819);
or U9143 (N_9143,N_8858,N_8477);
xnor U9144 (N_9144,N_8483,N_8193);
xor U9145 (N_9145,N_8064,N_8788);
nor U9146 (N_9146,N_8247,N_8592);
and U9147 (N_9147,N_8183,N_8463);
xor U9148 (N_9148,N_8333,N_8404);
nor U9149 (N_9149,N_8461,N_8697);
nand U9150 (N_9150,N_8435,N_8709);
nand U9151 (N_9151,N_8138,N_8155);
nand U9152 (N_9152,N_8391,N_8925);
nand U9153 (N_9153,N_8784,N_8420);
nor U9154 (N_9154,N_8582,N_8588);
or U9155 (N_9155,N_8224,N_8780);
nor U9156 (N_9156,N_8459,N_8502);
or U9157 (N_9157,N_8487,N_8809);
nor U9158 (N_9158,N_8132,N_8984);
nor U9159 (N_9159,N_8708,N_8845);
or U9160 (N_9160,N_8739,N_8770);
or U9161 (N_9161,N_8624,N_8864);
or U9162 (N_9162,N_8594,N_8440);
and U9163 (N_9163,N_8891,N_8751);
and U9164 (N_9164,N_8016,N_8851);
xor U9165 (N_9165,N_8716,N_8686);
nand U9166 (N_9166,N_8551,N_8453);
and U9167 (N_9167,N_8871,N_8657);
and U9168 (N_9168,N_8113,N_8887);
nor U9169 (N_9169,N_8294,N_8019);
nor U9170 (N_9170,N_8856,N_8872);
and U9171 (N_9171,N_8546,N_8506);
and U9172 (N_9172,N_8316,N_8797);
or U9173 (N_9173,N_8355,N_8033);
nor U9174 (N_9174,N_8707,N_8187);
or U9175 (N_9175,N_8619,N_8215);
nand U9176 (N_9176,N_8026,N_8238);
and U9177 (N_9177,N_8981,N_8370);
nand U9178 (N_9178,N_8982,N_8402);
nor U9179 (N_9179,N_8806,N_8166);
and U9180 (N_9180,N_8954,N_8496);
nor U9181 (N_9181,N_8098,N_8511);
nand U9182 (N_9182,N_8549,N_8272);
nand U9183 (N_9183,N_8207,N_8639);
and U9184 (N_9184,N_8239,N_8047);
and U9185 (N_9185,N_8617,N_8121);
or U9186 (N_9186,N_8206,N_8449);
or U9187 (N_9187,N_8452,N_8843);
and U9188 (N_9188,N_8774,N_8287);
xnor U9189 (N_9189,N_8539,N_8089);
and U9190 (N_9190,N_8083,N_8192);
and U9191 (N_9191,N_8250,N_8003);
and U9192 (N_9192,N_8754,N_8943);
nand U9193 (N_9193,N_8382,N_8825);
or U9194 (N_9194,N_8830,N_8691);
and U9195 (N_9195,N_8397,N_8020);
nor U9196 (N_9196,N_8450,N_8994);
xnor U9197 (N_9197,N_8371,N_8468);
and U9198 (N_9198,N_8794,N_8029);
xor U9199 (N_9199,N_8410,N_8808);
xnor U9200 (N_9200,N_8841,N_8607);
xnor U9201 (N_9201,N_8971,N_8263);
nand U9202 (N_9202,N_8421,N_8651);
and U9203 (N_9203,N_8812,N_8305);
and U9204 (N_9204,N_8277,N_8735);
nor U9205 (N_9205,N_8964,N_8665);
or U9206 (N_9206,N_8585,N_8365);
nand U9207 (N_9207,N_8810,N_8285);
and U9208 (N_9208,N_8885,N_8724);
nand U9209 (N_9209,N_8846,N_8361);
nor U9210 (N_9210,N_8127,N_8557);
xnor U9211 (N_9211,N_8080,N_8364);
xnor U9212 (N_9212,N_8641,N_8926);
nor U9213 (N_9213,N_8439,N_8161);
or U9214 (N_9214,N_8027,N_8800);
and U9215 (N_9215,N_8216,N_8414);
nand U9216 (N_9216,N_8713,N_8456);
and U9217 (N_9217,N_8852,N_8930);
xnor U9218 (N_9218,N_8043,N_8076);
or U9219 (N_9219,N_8011,N_8394);
nand U9220 (N_9220,N_8022,N_8907);
or U9221 (N_9221,N_8659,N_8375);
nand U9222 (N_9222,N_8348,N_8969);
nor U9223 (N_9223,N_8968,N_8918);
or U9224 (N_9224,N_8498,N_8908);
or U9225 (N_9225,N_8110,N_8550);
and U9226 (N_9226,N_8136,N_8598);
and U9227 (N_9227,N_8890,N_8554);
xor U9228 (N_9228,N_8738,N_8513);
or U9229 (N_9229,N_8729,N_8866);
and U9230 (N_9230,N_8184,N_8544);
nor U9231 (N_9231,N_8683,N_8211);
nor U9232 (N_9232,N_8936,N_8827);
nor U9233 (N_9233,N_8727,N_8910);
and U9234 (N_9234,N_8233,N_8343);
and U9235 (N_9235,N_8143,N_8349);
xor U9236 (N_9236,N_8458,N_8214);
or U9237 (N_9237,N_8025,N_8245);
xnor U9238 (N_9238,N_8644,N_8824);
xor U9239 (N_9239,N_8423,N_8654);
and U9240 (N_9240,N_8996,N_8661);
nand U9241 (N_9241,N_8267,N_8823);
nand U9242 (N_9242,N_8658,N_8615);
xnor U9243 (N_9243,N_8469,N_8951);
nor U9244 (N_9244,N_8430,N_8749);
and U9245 (N_9245,N_8955,N_8087);
nor U9246 (N_9246,N_8571,N_8219);
and U9247 (N_9247,N_8486,N_8618);
xnor U9248 (N_9248,N_8646,N_8384);
nand U9249 (N_9249,N_8360,N_8721);
xnor U9250 (N_9250,N_8861,N_8529);
and U9251 (N_9251,N_8374,N_8332);
or U9252 (N_9252,N_8249,N_8106);
nor U9253 (N_9253,N_8482,N_8660);
and U9254 (N_9254,N_8297,N_8437);
nor U9255 (N_9255,N_8917,N_8765);
and U9256 (N_9256,N_8293,N_8625);
or U9257 (N_9257,N_8762,N_8580);
nand U9258 (N_9258,N_8993,N_8501);
nand U9259 (N_9259,N_8553,N_8881);
nand U9260 (N_9260,N_8304,N_8940);
nand U9261 (N_9261,N_8627,N_8579);
or U9262 (N_9262,N_8479,N_8354);
and U9263 (N_9263,N_8979,N_8722);
xor U9264 (N_9264,N_8606,N_8680);
or U9265 (N_9265,N_8611,N_8050);
nor U9266 (N_9266,N_8896,N_8904);
xnor U9267 (N_9267,N_8134,N_8562);
xnor U9268 (N_9268,N_8052,N_8455);
nand U9269 (N_9269,N_8715,N_8787);
nand U9270 (N_9270,N_8232,N_8321);
xor U9271 (N_9271,N_8102,N_8419);
or U9272 (N_9272,N_8109,N_8133);
or U9273 (N_9273,N_8574,N_8884);
xnor U9274 (N_9274,N_8429,N_8900);
or U9275 (N_9275,N_8831,N_8764);
and U9276 (N_9276,N_8150,N_8248);
nand U9277 (N_9277,N_8160,N_8678);
and U9278 (N_9278,N_8328,N_8694);
and U9279 (N_9279,N_8378,N_8115);
nor U9280 (N_9280,N_8078,N_8778);
or U9281 (N_9281,N_8530,N_8065);
nand U9282 (N_9282,N_8693,N_8737);
or U9283 (N_9283,N_8040,N_8878);
xor U9284 (N_9284,N_8882,N_8362);
and U9285 (N_9285,N_8650,N_8091);
and U9286 (N_9286,N_8068,N_8494);
nor U9287 (N_9287,N_8614,N_8817);
nor U9288 (N_9288,N_8451,N_8569);
nor U9289 (N_9289,N_8992,N_8120);
xnor U9290 (N_9290,N_8976,N_8719);
nand U9291 (N_9291,N_8983,N_8789);
nor U9292 (N_9292,N_8303,N_8860);
xnor U9293 (N_9293,N_8066,N_8169);
or U9294 (N_9294,N_8676,N_8063);
nand U9295 (N_9295,N_8934,N_8002);
or U9296 (N_9296,N_8417,N_8698);
and U9297 (N_9297,N_8637,N_8488);
nand U9298 (N_9298,N_8503,N_8315);
nor U9299 (N_9299,N_8815,N_8425);
nor U9300 (N_9300,N_8491,N_8854);
nand U9301 (N_9301,N_8768,N_8892);
and U9302 (N_9302,N_8131,N_8225);
nand U9303 (N_9303,N_8966,N_8901);
or U9304 (N_9304,N_8291,N_8464);
xor U9305 (N_9305,N_8018,N_8230);
nand U9306 (N_9306,N_8935,N_8534);
and U9307 (N_9307,N_8886,N_8632);
nor U9308 (N_9308,N_8341,N_8145);
xor U9309 (N_9309,N_8432,N_8008);
nand U9310 (N_9310,N_8099,N_8141);
or U9311 (N_9311,N_8171,N_8745);
or U9312 (N_9312,N_8685,N_8149);
nor U9313 (N_9313,N_8923,N_8474);
nor U9314 (N_9314,N_8048,N_8416);
or U9315 (N_9315,N_8289,N_8679);
xor U9316 (N_9316,N_8411,N_8339);
xor U9317 (N_9317,N_8668,N_8779);
xnor U9318 (N_9318,N_8220,N_8441);
or U9319 (N_9319,N_8561,N_8288);
xor U9320 (N_9320,N_8733,N_8505);
or U9321 (N_9321,N_8647,N_8591);
nand U9322 (N_9322,N_8957,N_8998);
and U9323 (N_9323,N_8381,N_8140);
or U9324 (N_9324,N_8802,N_8282);
and U9325 (N_9325,N_8857,N_8621);
and U9326 (N_9326,N_8526,N_8177);
nor U9327 (N_9327,N_8176,N_8338);
or U9328 (N_9328,N_8369,N_8813);
nand U9329 (N_9329,N_8271,N_8443);
nor U9330 (N_9330,N_8528,N_8959);
xnor U9331 (N_9331,N_8096,N_8221);
nor U9332 (N_9332,N_8581,N_8775);
nor U9333 (N_9333,N_8137,N_8653);
xor U9334 (N_9334,N_8241,N_8681);
nand U9335 (N_9335,N_8392,N_8270);
or U9336 (N_9336,N_8049,N_8359);
xor U9337 (N_9337,N_8146,N_8720);
or U9338 (N_9338,N_8312,N_8344);
or U9339 (N_9339,N_8521,N_8092);
nand U9340 (N_9340,N_8084,N_8246);
and U9341 (N_9341,N_8055,N_8256);
nor U9342 (N_9342,N_8970,N_8870);
and U9343 (N_9343,N_8636,N_8163);
nand U9344 (N_9344,N_8032,N_8868);
or U9345 (N_9345,N_8100,N_8393);
nand U9346 (N_9346,N_8357,N_8489);
nand U9347 (N_9347,N_8527,N_8380);
nand U9348 (N_9348,N_8165,N_8258);
nand U9349 (N_9349,N_8112,N_8363);
xor U9350 (N_9350,N_8037,N_8237);
nor U9351 (N_9351,N_8311,N_8058);
or U9352 (N_9352,N_8833,N_8385);
and U9353 (N_9353,N_8125,N_8928);
nor U9354 (N_9354,N_8807,N_8937);
xor U9355 (N_9355,N_8929,N_8337);
or U9356 (N_9356,N_8766,N_8465);
xnor U9357 (N_9357,N_8820,N_8950);
nor U9358 (N_9358,N_8181,N_8274);
nor U9359 (N_9359,N_8108,N_8732);
nor U9360 (N_9360,N_8261,N_8999);
and U9361 (N_9361,N_8373,N_8500);
xnor U9362 (N_9362,N_8804,N_8564);
nor U9363 (N_9363,N_8097,N_8307);
xnor U9364 (N_9364,N_8028,N_8292);
nor U9365 (N_9365,N_8044,N_8705);
and U9366 (N_9366,N_8865,N_8548);
nor U9367 (N_9367,N_8666,N_8367);
and U9368 (N_9368,N_8690,N_8525);
nor U9369 (N_9369,N_8687,N_8888);
xor U9370 (N_9370,N_8567,N_8781);
xor U9371 (N_9371,N_8314,N_8558);
nand U9372 (N_9372,N_8744,N_8035);
and U9373 (N_9373,N_8814,N_8946);
or U9374 (N_9374,N_8279,N_8213);
or U9375 (N_9375,N_8634,N_8786);
xnor U9376 (N_9376,N_8535,N_8438);
nor U9377 (N_9377,N_8921,N_8536);
xor U9378 (N_9378,N_8010,N_8960);
or U9379 (N_9379,N_8995,N_8589);
nand U9380 (N_9380,N_8130,N_8387);
or U9381 (N_9381,N_8492,N_8756);
and U9382 (N_9382,N_8799,N_8898);
or U9383 (N_9383,N_8508,N_8152);
nand U9384 (N_9384,N_8462,N_8702);
and U9385 (N_9385,N_8927,N_8390);
xnor U9386 (N_9386,N_8675,N_8073);
or U9387 (N_9387,N_8266,N_8850);
nor U9388 (N_9388,N_8484,N_8948);
nor U9389 (N_9389,N_8205,N_8849);
and U9390 (N_9390,N_8199,N_8988);
nor U9391 (N_9391,N_8902,N_8226);
or U9392 (N_9392,N_8242,N_8542);
nand U9393 (N_9393,N_8793,N_8322);
and U9394 (N_9394,N_8753,N_8023);
xor U9395 (N_9395,N_8202,N_8182);
or U9396 (N_9396,N_8119,N_8541);
nand U9397 (N_9397,N_8295,N_8244);
or U9398 (N_9398,N_8593,N_8185);
nand U9399 (N_9399,N_8626,N_8782);
nand U9400 (N_9400,N_8911,N_8470);
nor U9401 (N_9401,N_8576,N_8129);
xor U9402 (N_9402,N_8481,N_8475);
and U9403 (N_9403,N_8801,N_8967);
nand U9404 (N_9404,N_8604,N_8255);
or U9405 (N_9405,N_8840,N_8699);
xnor U9406 (N_9406,N_8796,N_8575);
xnor U9407 (N_9407,N_8875,N_8061);
nor U9408 (N_9408,N_8446,N_8673);
or U9409 (N_9409,N_8015,N_8413);
xnor U9410 (N_9410,N_8519,N_8655);
nand U9411 (N_9411,N_8395,N_8445);
nand U9412 (N_9412,N_8517,N_8144);
and U9413 (N_9413,N_8004,N_8030);
nand U9414 (N_9414,N_8848,N_8913);
nor U9415 (N_9415,N_8883,N_8961);
nand U9416 (N_9416,N_8264,N_8070);
nand U9417 (N_9417,N_8842,N_8157);
and U9418 (N_9418,N_8538,N_8336);
or U9419 (N_9419,N_8036,N_8122);
and U9420 (N_9420,N_8974,N_8759);
and U9421 (N_9421,N_8700,N_8895);
nor U9422 (N_9422,N_8837,N_8568);
nand U9423 (N_9423,N_8329,N_8752);
nand U9424 (N_9424,N_8345,N_8628);
xnor U9425 (N_9425,N_8717,N_8792);
and U9426 (N_9426,N_8164,N_8684);
nand U9427 (N_9427,N_8916,N_8635);
nand U9428 (N_9428,N_8991,N_8399);
nor U9429 (N_9429,N_8507,N_8714);
xnor U9430 (N_9430,N_8512,N_8963);
and U9431 (N_9431,N_8103,N_8769);
nor U9432 (N_9432,N_8353,N_8869);
nor U9433 (N_9433,N_8711,N_8424);
nand U9434 (N_9434,N_8235,N_8730);
or U9435 (N_9435,N_8777,N_8376);
nor U9436 (N_9436,N_8609,N_8153);
nor U9437 (N_9437,N_8497,N_8000);
nor U9438 (N_9438,N_8667,N_8682);
nand U9439 (N_9439,N_8179,N_8795);
xnor U9440 (N_9440,N_8081,N_8853);
nor U9441 (N_9441,N_8167,N_8821);
nand U9442 (N_9442,N_8953,N_8862);
xor U9443 (N_9443,N_8734,N_8577);
xor U9444 (N_9444,N_8912,N_8377);
nor U9445 (N_9445,N_8645,N_8893);
xor U9446 (N_9446,N_8334,N_8879);
or U9447 (N_9447,N_8783,N_8021);
nand U9448 (N_9448,N_8082,N_8790);
xnor U9449 (N_9449,N_8139,N_8243);
xnor U9450 (N_9450,N_8915,N_8718);
xnor U9451 (N_9451,N_8706,N_8586);
xnor U9452 (N_9452,N_8670,N_8204);
or U9453 (N_9453,N_8335,N_8472);
and U9454 (N_9454,N_8325,N_8473);
or U9455 (N_9455,N_8260,N_8836);
nor U9456 (N_9456,N_8408,N_8467);
nand U9457 (N_9457,N_8537,N_8695);
xnor U9458 (N_9458,N_8210,N_8228);
and U9459 (N_9459,N_8600,N_8223);
or U9460 (N_9460,N_8855,N_8062);
xor U9461 (N_9461,N_8358,N_8039);
and U9462 (N_9462,N_8031,N_8005);
nand U9463 (N_9463,N_8642,N_8042);
xnor U9464 (N_9464,N_8101,N_8493);
xor U9465 (N_9465,N_8570,N_8444);
nor U9466 (N_9466,N_8251,N_8398);
xnor U9467 (N_9467,N_8017,N_8595);
nor U9468 (N_9468,N_8828,N_8952);
and U9469 (N_9469,N_8478,N_8773);
xnor U9470 (N_9470,N_8603,N_8320);
nand U9471 (N_9471,N_8173,N_8196);
or U9472 (N_9472,N_8107,N_8041);
nand U9473 (N_9473,N_8826,N_8543);
xor U9474 (N_9474,N_8610,N_8776);
xnor U9475 (N_9475,N_8608,N_8273);
and U9476 (N_9476,N_8516,N_8060);
nor U9477 (N_9477,N_8124,N_8476);
and U9478 (N_9478,N_8201,N_8090);
nand U9479 (N_9479,N_8922,N_8590);
nand U9480 (N_9480,N_8956,N_8533);
and U9481 (N_9481,N_8741,N_8758);
or U9482 (N_9482,N_8747,N_8743);
nand U9483 (N_9483,N_8188,N_8331);
nor U9484 (N_9484,N_8431,N_8622);
or U9485 (N_9485,N_8290,N_8342);
nand U9486 (N_9486,N_8085,N_8159);
nand U9487 (N_9487,N_8433,N_8116);
or U9488 (N_9488,N_8317,N_8520);
and U9489 (N_9489,N_8958,N_8123);
nand U9490 (N_9490,N_8436,N_8540);
or U9491 (N_9491,N_8284,N_8612);
xor U9492 (N_9492,N_8757,N_8074);
nand U9493 (N_9493,N_8560,N_8932);
nor U9494 (N_9494,N_8175,N_8428);
or U9495 (N_9495,N_8514,N_8405);
nor U9496 (N_9496,N_8454,N_8212);
or U9497 (N_9497,N_8268,N_8259);
and U9498 (N_9498,N_8839,N_8401);
nor U9499 (N_9499,N_8067,N_8286);
and U9500 (N_9500,N_8838,N_8657);
nor U9501 (N_9501,N_8236,N_8034);
nand U9502 (N_9502,N_8818,N_8159);
nor U9503 (N_9503,N_8386,N_8671);
xor U9504 (N_9504,N_8836,N_8041);
or U9505 (N_9505,N_8837,N_8770);
nand U9506 (N_9506,N_8498,N_8484);
xnor U9507 (N_9507,N_8068,N_8344);
nor U9508 (N_9508,N_8793,N_8981);
and U9509 (N_9509,N_8095,N_8074);
nor U9510 (N_9510,N_8867,N_8696);
nor U9511 (N_9511,N_8944,N_8350);
or U9512 (N_9512,N_8314,N_8278);
xnor U9513 (N_9513,N_8641,N_8854);
nor U9514 (N_9514,N_8779,N_8685);
xor U9515 (N_9515,N_8872,N_8136);
and U9516 (N_9516,N_8877,N_8334);
xnor U9517 (N_9517,N_8564,N_8158);
nor U9518 (N_9518,N_8454,N_8327);
nand U9519 (N_9519,N_8776,N_8468);
or U9520 (N_9520,N_8004,N_8378);
or U9521 (N_9521,N_8448,N_8132);
and U9522 (N_9522,N_8827,N_8699);
or U9523 (N_9523,N_8728,N_8208);
and U9524 (N_9524,N_8662,N_8766);
or U9525 (N_9525,N_8930,N_8230);
nor U9526 (N_9526,N_8871,N_8372);
nor U9527 (N_9527,N_8765,N_8093);
or U9528 (N_9528,N_8487,N_8301);
nor U9529 (N_9529,N_8461,N_8384);
xnor U9530 (N_9530,N_8816,N_8942);
nor U9531 (N_9531,N_8210,N_8078);
xnor U9532 (N_9532,N_8513,N_8881);
or U9533 (N_9533,N_8754,N_8349);
or U9534 (N_9534,N_8481,N_8752);
or U9535 (N_9535,N_8111,N_8982);
nor U9536 (N_9536,N_8366,N_8646);
and U9537 (N_9537,N_8565,N_8484);
and U9538 (N_9538,N_8398,N_8962);
nor U9539 (N_9539,N_8350,N_8760);
and U9540 (N_9540,N_8554,N_8301);
nand U9541 (N_9541,N_8238,N_8116);
nand U9542 (N_9542,N_8736,N_8531);
xnor U9543 (N_9543,N_8589,N_8862);
nor U9544 (N_9544,N_8063,N_8846);
nor U9545 (N_9545,N_8598,N_8772);
and U9546 (N_9546,N_8453,N_8538);
nand U9547 (N_9547,N_8806,N_8795);
and U9548 (N_9548,N_8364,N_8136);
xnor U9549 (N_9549,N_8439,N_8472);
xnor U9550 (N_9550,N_8642,N_8192);
and U9551 (N_9551,N_8383,N_8183);
or U9552 (N_9552,N_8105,N_8584);
xor U9553 (N_9553,N_8126,N_8802);
nand U9554 (N_9554,N_8761,N_8426);
nand U9555 (N_9555,N_8904,N_8376);
nand U9556 (N_9556,N_8928,N_8841);
xnor U9557 (N_9557,N_8858,N_8148);
and U9558 (N_9558,N_8757,N_8840);
or U9559 (N_9559,N_8817,N_8338);
and U9560 (N_9560,N_8732,N_8609);
nor U9561 (N_9561,N_8332,N_8021);
nand U9562 (N_9562,N_8703,N_8112);
xnor U9563 (N_9563,N_8124,N_8425);
xor U9564 (N_9564,N_8626,N_8310);
and U9565 (N_9565,N_8403,N_8872);
or U9566 (N_9566,N_8053,N_8016);
nand U9567 (N_9567,N_8162,N_8705);
nor U9568 (N_9568,N_8413,N_8945);
xor U9569 (N_9569,N_8012,N_8713);
xor U9570 (N_9570,N_8059,N_8266);
or U9571 (N_9571,N_8597,N_8088);
nor U9572 (N_9572,N_8030,N_8866);
and U9573 (N_9573,N_8735,N_8695);
and U9574 (N_9574,N_8365,N_8462);
or U9575 (N_9575,N_8963,N_8786);
nand U9576 (N_9576,N_8184,N_8435);
or U9577 (N_9577,N_8943,N_8178);
and U9578 (N_9578,N_8020,N_8539);
xor U9579 (N_9579,N_8796,N_8938);
xnor U9580 (N_9580,N_8966,N_8215);
nor U9581 (N_9581,N_8624,N_8721);
and U9582 (N_9582,N_8148,N_8245);
or U9583 (N_9583,N_8184,N_8593);
or U9584 (N_9584,N_8148,N_8670);
nor U9585 (N_9585,N_8293,N_8661);
and U9586 (N_9586,N_8399,N_8558);
nand U9587 (N_9587,N_8440,N_8230);
xor U9588 (N_9588,N_8340,N_8075);
or U9589 (N_9589,N_8505,N_8351);
xnor U9590 (N_9590,N_8715,N_8923);
nand U9591 (N_9591,N_8028,N_8288);
or U9592 (N_9592,N_8328,N_8531);
xnor U9593 (N_9593,N_8968,N_8929);
nand U9594 (N_9594,N_8242,N_8730);
nor U9595 (N_9595,N_8869,N_8890);
and U9596 (N_9596,N_8834,N_8119);
nand U9597 (N_9597,N_8290,N_8050);
xnor U9598 (N_9598,N_8503,N_8931);
or U9599 (N_9599,N_8917,N_8209);
nand U9600 (N_9600,N_8822,N_8547);
xor U9601 (N_9601,N_8727,N_8979);
nor U9602 (N_9602,N_8414,N_8422);
xor U9603 (N_9603,N_8319,N_8999);
xor U9604 (N_9604,N_8426,N_8350);
and U9605 (N_9605,N_8495,N_8087);
xor U9606 (N_9606,N_8154,N_8803);
or U9607 (N_9607,N_8047,N_8716);
nand U9608 (N_9608,N_8476,N_8699);
xor U9609 (N_9609,N_8988,N_8958);
nand U9610 (N_9610,N_8780,N_8710);
or U9611 (N_9611,N_8883,N_8303);
and U9612 (N_9612,N_8559,N_8878);
nand U9613 (N_9613,N_8730,N_8448);
xnor U9614 (N_9614,N_8136,N_8874);
and U9615 (N_9615,N_8877,N_8817);
nor U9616 (N_9616,N_8063,N_8616);
nor U9617 (N_9617,N_8256,N_8013);
xor U9618 (N_9618,N_8892,N_8596);
nor U9619 (N_9619,N_8251,N_8376);
nor U9620 (N_9620,N_8342,N_8181);
or U9621 (N_9621,N_8406,N_8095);
nand U9622 (N_9622,N_8078,N_8166);
nor U9623 (N_9623,N_8490,N_8920);
nor U9624 (N_9624,N_8906,N_8491);
or U9625 (N_9625,N_8971,N_8713);
nand U9626 (N_9626,N_8471,N_8250);
xnor U9627 (N_9627,N_8657,N_8437);
or U9628 (N_9628,N_8902,N_8593);
nand U9629 (N_9629,N_8588,N_8045);
xnor U9630 (N_9630,N_8654,N_8118);
nand U9631 (N_9631,N_8180,N_8426);
nand U9632 (N_9632,N_8336,N_8640);
nor U9633 (N_9633,N_8017,N_8547);
or U9634 (N_9634,N_8223,N_8624);
xnor U9635 (N_9635,N_8811,N_8697);
and U9636 (N_9636,N_8973,N_8871);
or U9637 (N_9637,N_8437,N_8011);
nand U9638 (N_9638,N_8753,N_8083);
nor U9639 (N_9639,N_8018,N_8542);
xnor U9640 (N_9640,N_8486,N_8796);
nor U9641 (N_9641,N_8175,N_8575);
xnor U9642 (N_9642,N_8696,N_8793);
xnor U9643 (N_9643,N_8434,N_8251);
or U9644 (N_9644,N_8992,N_8799);
nand U9645 (N_9645,N_8432,N_8019);
nor U9646 (N_9646,N_8591,N_8372);
and U9647 (N_9647,N_8505,N_8315);
xor U9648 (N_9648,N_8879,N_8898);
nand U9649 (N_9649,N_8806,N_8168);
and U9650 (N_9650,N_8800,N_8153);
nand U9651 (N_9651,N_8318,N_8700);
or U9652 (N_9652,N_8436,N_8837);
and U9653 (N_9653,N_8112,N_8882);
nand U9654 (N_9654,N_8172,N_8586);
or U9655 (N_9655,N_8967,N_8197);
nor U9656 (N_9656,N_8272,N_8138);
and U9657 (N_9657,N_8217,N_8821);
xnor U9658 (N_9658,N_8440,N_8001);
and U9659 (N_9659,N_8032,N_8344);
xor U9660 (N_9660,N_8699,N_8031);
nor U9661 (N_9661,N_8467,N_8139);
and U9662 (N_9662,N_8512,N_8518);
nor U9663 (N_9663,N_8369,N_8106);
nand U9664 (N_9664,N_8133,N_8077);
xor U9665 (N_9665,N_8366,N_8427);
xor U9666 (N_9666,N_8751,N_8853);
nand U9667 (N_9667,N_8259,N_8522);
xnor U9668 (N_9668,N_8534,N_8900);
nor U9669 (N_9669,N_8469,N_8993);
nor U9670 (N_9670,N_8931,N_8354);
nand U9671 (N_9671,N_8769,N_8857);
nand U9672 (N_9672,N_8369,N_8933);
nor U9673 (N_9673,N_8280,N_8637);
or U9674 (N_9674,N_8484,N_8191);
xor U9675 (N_9675,N_8583,N_8613);
or U9676 (N_9676,N_8690,N_8190);
xor U9677 (N_9677,N_8169,N_8186);
xor U9678 (N_9678,N_8264,N_8579);
or U9679 (N_9679,N_8274,N_8926);
xnor U9680 (N_9680,N_8998,N_8668);
nand U9681 (N_9681,N_8871,N_8018);
and U9682 (N_9682,N_8439,N_8504);
or U9683 (N_9683,N_8013,N_8845);
nand U9684 (N_9684,N_8723,N_8563);
nor U9685 (N_9685,N_8216,N_8815);
nor U9686 (N_9686,N_8074,N_8721);
or U9687 (N_9687,N_8436,N_8421);
xnor U9688 (N_9688,N_8522,N_8795);
or U9689 (N_9689,N_8893,N_8555);
nor U9690 (N_9690,N_8298,N_8794);
nor U9691 (N_9691,N_8784,N_8968);
nor U9692 (N_9692,N_8534,N_8577);
nor U9693 (N_9693,N_8353,N_8504);
xor U9694 (N_9694,N_8458,N_8201);
and U9695 (N_9695,N_8788,N_8837);
xor U9696 (N_9696,N_8509,N_8910);
nand U9697 (N_9697,N_8459,N_8716);
or U9698 (N_9698,N_8676,N_8182);
nand U9699 (N_9699,N_8997,N_8208);
nand U9700 (N_9700,N_8726,N_8866);
or U9701 (N_9701,N_8965,N_8507);
or U9702 (N_9702,N_8583,N_8983);
and U9703 (N_9703,N_8374,N_8031);
nor U9704 (N_9704,N_8417,N_8739);
nand U9705 (N_9705,N_8385,N_8944);
nor U9706 (N_9706,N_8325,N_8542);
xor U9707 (N_9707,N_8626,N_8933);
or U9708 (N_9708,N_8232,N_8486);
and U9709 (N_9709,N_8150,N_8376);
xnor U9710 (N_9710,N_8514,N_8422);
nand U9711 (N_9711,N_8874,N_8238);
nor U9712 (N_9712,N_8529,N_8927);
xor U9713 (N_9713,N_8615,N_8486);
nor U9714 (N_9714,N_8548,N_8724);
or U9715 (N_9715,N_8307,N_8367);
xnor U9716 (N_9716,N_8846,N_8604);
and U9717 (N_9717,N_8214,N_8926);
and U9718 (N_9718,N_8381,N_8915);
nand U9719 (N_9719,N_8161,N_8297);
or U9720 (N_9720,N_8264,N_8369);
nand U9721 (N_9721,N_8167,N_8034);
and U9722 (N_9722,N_8199,N_8182);
and U9723 (N_9723,N_8080,N_8547);
nand U9724 (N_9724,N_8241,N_8232);
nor U9725 (N_9725,N_8008,N_8628);
xnor U9726 (N_9726,N_8545,N_8138);
nor U9727 (N_9727,N_8888,N_8510);
xnor U9728 (N_9728,N_8487,N_8255);
xnor U9729 (N_9729,N_8680,N_8025);
or U9730 (N_9730,N_8019,N_8420);
and U9731 (N_9731,N_8782,N_8369);
nor U9732 (N_9732,N_8570,N_8713);
nand U9733 (N_9733,N_8737,N_8688);
and U9734 (N_9734,N_8767,N_8996);
and U9735 (N_9735,N_8591,N_8549);
nand U9736 (N_9736,N_8119,N_8359);
and U9737 (N_9737,N_8192,N_8239);
or U9738 (N_9738,N_8611,N_8672);
nor U9739 (N_9739,N_8056,N_8161);
and U9740 (N_9740,N_8314,N_8434);
or U9741 (N_9741,N_8703,N_8825);
nand U9742 (N_9742,N_8574,N_8559);
xor U9743 (N_9743,N_8316,N_8588);
nand U9744 (N_9744,N_8273,N_8544);
nor U9745 (N_9745,N_8548,N_8801);
xor U9746 (N_9746,N_8682,N_8413);
nand U9747 (N_9747,N_8449,N_8815);
and U9748 (N_9748,N_8804,N_8867);
and U9749 (N_9749,N_8615,N_8057);
nor U9750 (N_9750,N_8542,N_8489);
xor U9751 (N_9751,N_8456,N_8203);
nor U9752 (N_9752,N_8828,N_8786);
xor U9753 (N_9753,N_8142,N_8000);
nor U9754 (N_9754,N_8424,N_8982);
or U9755 (N_9755,N_8390,N_8289);
nand U9756 (N_9756,N_8155,N_8559);
nor U9757 (N_9757,N_8946,N_8314);
xor U9758 (N_9758,N_8773,N_8151);
nand U9759 (N_9759,N_8730,N_8901);
xnor U9760 (N_9760,N_8217,N_8063);
xnor U9761 (N_9761,N_8029,N_8703);
nand U9762 (N_9762,N_8620,N_8507);
or U9763 (N_9763,N_8531,N_8625);
or U9764 (N_9764,N_8930,N_8795);
nor U9765 (N_9765,N_8273,N_8330);
nand U9766 (N_9766,N_8721,N_8251);
and U9767 (N_9767,N_8359,N_8173);
or U9768 (N_9768,N_8214,N_8947);
nand U9769 (N_9769,N_8962,N_8060);
nand U9770 (N_9770,N_8266,N_8712);
or U9771 (N_9771,N_8697,N_8791);
and U9772 (N_9772,N_8960,N_8466);
nor U9773 (N_9773,N_8032,N_8390);
nand U9774 (N_9774,N_8587,N_8548);
nor U9775 (N_9775,N_8167,N_8227);
nor U9776 (N_9776,N_8311,N_8261);
and U9777 (N_9777,N_8224,N_8668);
nand U9778 (N_9778,N_8408,N_8511);
xnor U9779 (N_9779,N_8269,N_8215);
nand U9780 (N_9780,N_8539,N_8327);
or U9781 (N_9781,N_8639,N_8981);
nand U9782 (N_9782,N_8874,N_8956);
xor U9783 (N_9783,N_8826,N_8279);
or U9784 (N_9784,N_8224,N_8004);
xnor U9785 (N_9785,N_8620,N_8241);
or U9786 (N_9786,N_8587,N_8201);
xnor U9787 (N_9787,N_8292,N_8462);
nor U9788 (N_9788,N_8852,N_8369);
xnor U9789 (N_9789,N_8161,N_8596);
and U9790 (N_9790,N_8053,N_8950);
xor U9791 (N_9791,N_8519,N_8903);
or U9792 (N_9792,N_8456,N_8248);
xor U9793 (N_9793,N_8476,N_8787);
xnor U9794 (N_9794,N_8212,N_8614);
xor U9795 (N_9795,N_8681,N_8900);
nor U9796 (N_9796,N_8289,N_8727);
and U9797 (N_9797,N_8560,N_8309);
or U9798 (N_9798,N_8383,N_8576);
nor U9799 (N_9799,N_8689,N_8737);
or U9800 (N_9800,N_8003,N_8998);
and U9801 (N_9801,N_8862,N_8056);
and U9802 (N_9802,N_8298,N_8574);
xnor U9803 (N_9803,N_8000,N_8697);
or U9804 (N_9804,N_8001,N_8069);
nand U9805 (N_9805,N_8083,N_8311);
and U9806 (N_9806,N_8415,N_8187);
and U9807 (N_9807,N_8174,N_8764);
nor U9808 (N_9808,N_8000,N_8952);
or U9809 (N_9809,N_8932,N_8636);
nand U9810 (N_9810,N_8480,N_8250);
nor U9811 (N_9811,N_8578,N_8754);
or U9812 (N_9812,N_8237,N_8430);
xnor U9813 (N_9813,N_8159,N_8287);
nand U9814 (N_9814,N_8958,N_8745);
and U9815 (N_9815,N_8448,N_8871);
xor U9816 (N_9816,N_8413,N_8289);
or U9817 (N_9817,N_8956,N_8639);
nor U9818 (N_9818,N_8511,N_8268);
or U9819 (N_9819,N_8689,N_8747);
nand U9820 (N_9820,N_8481,N_8338);
xnor U9821 (N_9821,N_8577,N_8889);
nor U9822 (N_9822,N_8374,N_8874);
or U9823 (N_9823,N_8157,N_8147);
nor U9824 (N_9824,N_8699,N_8345);
or U9825 (N_9825,N_8541,N_8132);
nand U9826 (N_9826,N_8192,N_8514);
nand U9827 (N_9827,N_8271,N_8811);
and U9828 (N_9828,N_8290,N_8877);
nor U9829 (N_9829,N_8597,N_8404);
nor U9830 (N_9830,N_8028,N_8707);
and U9831 (N_9831,N_8760,N_8812);
and U9832 (N_9832,N_8623,N_8012);
or U9833 (N_9833,N_8074,N_8037);
and U9834 (N_9834,N_8427,N_8133);
nand U9835 (N_9835,N_8953,N_8347);
nand U9836 (N_9836,N_8248,N_8561);
nor U9837 (N_9837,N_8201,N_8505);
xor U9838 (N_9838,N_8757,N_8018);
nand U9839 (N_9839,N_8148,N_8544);
nand U9840 (N_9840,N_8743,N_8641);
xnor U9841 (N_9841,N_8384,N_8626);
and U9842 (N_9842,N_8664,N_8272);
nor U9843 (N_9843,N_8253,N_8663);
nor U9844 (N_9844,N_8983,N_8168);
and U9845 (N_9845,N_8728,N_8535);
nor U9846 (N_9846,N_8912,N_8742);
nor U9847 (N_9847,N_8596,N_8655);
and U9848 (N_9848,N_8580,N_8240);
xnor U9849 (N_9849,N_8451,N_8402);
nor U9850 (N_9850,N_8381,N_8936);
or U9851 (N_9851,N_8544,N_8523);
and U9852 (N_9852,N_8680,N_8757);
xnor U9853 (N_9853,N_8487,N_8499);
xor U9854 (N_9854,N_8998,N_8892);
and U9855 (N_9855,N_8272,N_8260);
and U9856 (N_9856,N_8334,N_8421);
nand U9857 (N_9857,N_8669,N_8768);
nand U9858 (N_9858,N_8919,N_8085);
xor U9859 (N_9859,N_8391,N_8709);
nor U9860 (N_9860,N_8405,N_8343);
xnor U9861 (N_9861,N_8194,N_8696);
nor U9862 (N_9862,N_8494,N_8325);
xor U9863 (N_9863,N_8922,N_8959);
or U9864 (N_9864,N_8534,N_8452);
xnor U9865 (N_9865,N_8851,N_8620);
and U9866 (N_9866,N_8701,N_8479);
and U9867 (N_9867,N_8005,N_8371);
or U9868 (N_9868,N_8335,N_8212);
nor U9869 (N_9869,N_8353,N_8200);
nor U9870 (N_9870,N_8616,N_8979);
or U9871 (N_9871,N_8532,N_8036);
nor U9872 (N_9872,N_8104,N_8254);
or U9873 (N_9873,N_8022,N_8557);
and U9874 (N_9874,N_8176,N_8446);
xor U9875 (N_9875,N_8777,N_8130);
or U9876 (N_9876,N_8156,N_8231);
and U9877 (N_9877,N_8185,N_8934);
xnor U9878 (N_9878,N_8072,N_8318);
xnor U9879 (N_9879,N_8101,N_8888);
or U9880 (N_9880,N_8402,N_8631);
and U9881 (N_9881,N_8302,N_8540);
or U9882 (N_9882,N_8630,N_8712);
nor U9883 (N_9883,N_8137,N_8394);
xor U9884 (N_9884,N_8338,N_8756);
and U9885 (N_9885,N_8052,N_8491);
nor U9886 (N_9886,N_8468,N_8742);
nand U9887 (N_9887,N_8218,N_8065);
nand U9888 (N_9888,N_8881,N_8566);
xor U9889 (N_9889,N_8860,N_8298);
nor U9890 (N_9890,N_8615,N_8122);
or U9891 (N_9891,N_8996,N_8503);
and U9892 (N_9892,N_8437,N_8770);
xnor U9893 (N_9893,N_8557,N_8661);
nand U9894 (N_9894,N_8034,N_8870);
nor U9895 (N_9895,N_8819,N_8300);
nor U9896 (N_9896,N_8927,N_8157);
xor U9897 (N_9897,N_8997,N_8886);
or U9898 (N_9898,N_8237,N_8285);
nor U9899 (N_9899,N_8882,N_8435);
and U9900 (N_9900,N_8447,N_8623);
xor U9901 (N_9901,N_8670,N_8788);
or U9902 (N_9902,N_8780,N_8672);
nand U9903 (N_9903,N_8775,N_8393);
and U9904 (N_9904,N_8174,N_8296);
xor U9905 (N_9905,N_8076,N_8056);
nand U9906 (N_9906,N_8004,N_8497);
and U9907 (N_9907,N_8082,N_8002);
nand U9908 (N_9908,N_8024,N_8283);
nand U9909 (N_9909,N_8591,N_8996);
nor U9910 (N_9910,N_8264,N_8477);
nand U9911 (N_9911,N_8541,N_8960);
and U9912 (N_9912,N_8070,N_8027);
or U9913 (N_9913,N_8049,N_8788);
nor U9914 (N_9914,N_8207,N_8230);
nand U9915 (N_9915,N_8662,N_8573);
and U9916 (N_9916,N_8582,N_8121);
xor U9917 (N_9917,N_8491,N_8793);
nand U9918 (N_9918,N_8001,N_8788);
or U9919 (N_9919,N_8790,N_8384);
nand U9920 (N_9920,N_8615,N_8471);
or U9921 (N_9921,N_8210,N_8173);
or U9922 (N_9922,N_8104,N_8349);
and U9923 (N_9923,N_8254,N_8207);
nand U9924 (N_9924,N_8575,N_8650);
or U9925 (N_9925,N_8299,N_8689);
nor U9926 (N_9926,N_8982,N_8572);
nand U9927 (N_9927,N_8375,N_8354);
or U9928 (N_9928,N_8627,N_8096);
nor U9929 (N_9929,N_8860,N_8546);
nor U9930 (N_9930,N_8685,N_8186);
nand U9931 (N_9931,N_8738,N_8555);
and U9932 (N_9932,N_8491,N_8423);
nand U9933 (N_9933,N_8461,N_8926);
xnor U9934 (N_9934,N_8150,N_8442);
xnor U9935 (N_9935,N_8842,N_8208);
and U9936 (N_9936,N_8393,N_8079);
xor U9937 (N_9937,N_8010,N_8105);
nand U9938 (N_9938,N_8687,N_8965);
nand U9939 (N_9939,N_8398,N_8577);
nand U9940 (N_9940,N_8442,N_8521);
nor U9941 (N_9941,N_8587,N_8423);
and U9942 (N_9942,N_8160,N_8535);
or U9943 (N_9943,N_8873,N_8049);
xnor U9944 (N_9944,N_8677,N_8904);
nand U9945 (N_9945,N_8100,N_8556);
and U9946 (N_9946,N_8704,N_8358);
nor U9947 (N_9947,N_8836,N_8615);
nand U9948 (N_9948,N_8725,N_8349);
nor U9949 (N_9949,N_8888,N_8802);
xor U9950 (N_9950,N_8860,N_8729);
or U9951 (N_9951,N_8779,N_8691);
and U9952 (N_9952,N_8931,N_8020);
nand U9953 (N_9953,N_8045,N_8517);
nor U9954 (N_9954,N_8363,N_8369);
nor U9955 (N_9955,N_8275,N_8511);
nor U9956 (N_9956,N_8200,N_8464);
and U9957 (N_9957,N_8646,N_8643);
or U9958 (N_9958,N_8897,N_8490);
nand U9959 (N_9959,N_8009,N_8622);
nand U9960 (N_9960,N_8856,N_8613);
nand U9961 (N_9961,N_8845,N_8096);
and U9962 (N_9962,N_8885,N_8386);
nand U9963 (N_9963,N_8298,N_8585);
nand U9964 (N_9964,N_8374,N_8900);
nor U9965 (N_9965,N_8127,N_8071);
xor U9966 (N_9966,N_8670,N_8947);
and U9967 (N_9967,N_8187,N_8283);
nor U9968 (N_9968,N_8905,N_8663);
and U9969 (N_9969,N_8842,N_8546);
nand U9970 (N_9970,N_8712,N_8356);
xor U9971 (N_9971,N_8585,N_8377);
nor U9972 (N_9972,N_8029,N_8526);
and U9973 (N_9973,N_8575,N_8685);
and U9974 (N_9974,N_8761,N_8208);
or U9975 (N_9975,N_8779,N_8775);
nor U9976 (N_9976,N_8729,N_8503);
xnor U9977 (N_9977,N_8086,N_8171);
nor U9978 (N_9978,N_8055,N_8087);
nand U9979 (N_9979,N_8535,N_8163);
or U9980 (N_9980,N_8502,N_8983);
and U9981 (N_9981,N_8916,N_8972);
or U9982 (N_9982,N_8057,N_8499);
xnor U9983 (N_9983,N_8506,N_8669);
or U9984 (N_9984,N_8182,N_8530);
and U9985 (N_9985,N_8460,N_8389);
and U9986 (N_9986,N_8586,N_8610);
and U9987 (N_9987,N_8490,N_8495);
or U9988 (N_9988,N_8904,N_8031);
and U9989 (N_9989,N_8825,N_8386);
nor U9990 (N_9990,N_8134,N_8236);
and U9991 (N_9991,N_8906,N_8247);
xnor U9992 (N_9992,N_8063,N_8832);
nand U9993 (N_9993,N_8537,N_8023);
and U9994 (N_9994,N_8061,N_8252);
xnor U9995 (N_9995,N_8804,N_8864);
xnor U9996 (N_9996,N_8286,N_8575);
xor U9997 (N_9997,N_8725,N_8137);
and U9998 (N_9998,N_8478,N_8888);
nand U9999 (N_9999,N_8915,N_8436);
or U10000 (N_10000,N_9997,N_9364);
xor U10001 (N_10001,N_9657,N_9496);
xnor U10002 (N_10002,N_9709,N_9960);
or U10003 (N_10003,N_9872,N_9635);
nor U10004 (N_10004,N_9253,N_9204);
nor U10005 (N_10005,N_9083,N_9297);
nor U10006 (N_10006,N_9691,N_9039);
or U10007 (N_10007,N_9158,N_9379);
nand U10008 (N_10008,N_9086,N_9862);
and U10009 (N_10009,N_9205,N_9510);
nor U10010 (N_10010,N_9331,N_9559);
and U10011 (N_10011,N_9308,N_9285);
xnor U10012 (N_10012,N_9237,N_9777);
nor U10013 (N_10013,N_9233,N_9725);
nor U10014 (N_10014,N_9455,N_9956);
or U10015 (N_10015,N_9197,N_9181);
nor U10016 (N_10016,N_9921,N_9460);
nand U10017 (N_10017,N_9164,N_9954);
and U10018 (N_10018,N_9342,N_9411);
or U10019 (N_10019,N_9281,N_9433);
nand U10020 (N_10020,N_9151,N_9140);
xnor U10021 (N_10021,N_9974,N_9724);
nand U10022 (N_10022,N_9336,N_9699);
or U10023 (N_10023,N_9917,N_9256);
nand U10024 (N_10024,N_9275,N_9080);
or U10025 (N_10025,N_9525,N_9983);
or U10026 (N_10026,N_9058,N_9685);
nor U10027 (N_10027,N_9044,N_9515);
and U10028 (N_10028,N_9070,N_9671);
and U10029 (N_10029,N_9634,N_9200);
or U10030 (N_10030,N_9560,N_9866);
and U10031 (N_10031,N_9797,N_9268);
xnor U10032 (N_10032,N_9992,N_9792);
xor U10033 (N_10033,N_9823,N_9684);
and U10034 (N_10034,N_9071,N_9130);
nand U10035 (N_10035,N_9841,N_9500);
nor U10036 (N_10036,N_9489,N_9615);
and U10037 (N_10037,N_9776,N_9739);
nor U10038 (N_10038,N_9572,N_9394);
xor U10039 (N_10039,N_9064,N_9891);
nand U10040 (N_10040,N_9230,N_9869);
and U10041 (N_10041,N_9661,N_9113);
nor U10042 (N_10042,N_9479,N_9103);
and U10043 (N_10043,N_9213,N_9734);
nand U10044 (N_10044,N_9410,N_9643);
nor U10045 (N_10045,N_9101,N_9918);
and U10046 (N_10046,N_9073,N_9348);
xnor U10047 (N_10047,N_9024,N_9929);
xor U10048 (N_10048,N_9988,N_9408);
nor U10049 (N_10049,N_9888,N_9374);
or U10050 (N_10050,N_9224,N_9987);
nor U10051 (N_10051,N_9258,N_9371);
and U10052 (N_10052,N_9265,N_9472);
or U10053 (N_10053,N_9690,N_9577);
or U10054 (N_10054,N_9787,N_9782);
or U10055 (N_10055,N_9604,N_9445);
nand U10056 (N_10056,N_9856,N_9404);
or U10057 (N_10057,N_9284,N_9169);
or U10058 (N_10058,N_9074,N_9673);
nand U10059 (N_10059,N_9937,N_9287);
nand U10060 (N_10060,N_9835,N_9764);
xnor U10061 (N_10061,N_9859,N_9844);
or U10062 (N_10062,N_9640,N_9625);
nor U10063 (N_10063,N_9139,N_9023);
nor U10064 (N_10064,N_9380,N_9007);
and U10065 (N_10065,N_9965,N_9104);
and U10066 (N_10066,N_9340,N_9100);
xor U10067 (N_10067,N_9530,N_9332);
or U10068 (N_10068,N_9211,N_9497);
xor U10069 (N_10069,N_9748,N_9943);
nand U10070 (N_10070,N_9566,N_9629);
nor U10071 (N_10071,N_9520,N_9703);
xor U10072 (N_10072,N_9939,N_9273);
and U10073 (N_10073,N_9546,N_9579);
or U10074 (N_10074,N_9850,N_9432);
xor U10075 (N_10075,N_9437,N_9123);
nor U10076 (N_10076,N_9301,N_9522);
and U10077 (N_10077,N_9060,N_9329);
or U10078 (N_10078,N_9675,N_9234);
nor U10079 (N_10079,N_9976,N_9677);
and U10080 (N_10080,N_9318,N_9619);
xor U10081 (N_10081,N_9183,N_9356);
nand U10082 (N_10082,N_9467,N_9786);
or U10083 (N_10083,N_9352,N_9305);
or U10084 (N_10084,N_9798,N_9938);
xor U10085 (N_10085,N_9499,N_9189);
nor U10086 (N_10086,N_9138,N_9470);
nand U10087 (N_10087,N_9621,N_9264);
or U10088 (N_10088,N_9042,N_9680);
nor U10089 (N_10089,N_9879,N_9365);
or U10090 (N_10090,N_9958,N_9814);
and U10091 (N_10091,N_9267,N_9926);
and U10092 (N_10092,N_9737,N_9424);
nand U10093 (N_10093,N_9706,N_9442);
xor U10094 (N_10094,N_9475,N_9541);
nand U10095 (N_10095,N_9434,N_9344);
nor U10096 (N_10096,N_9214,N_9735);
nor U10097 (N_10097,N_9391,N_9067);
nand U10098 (N_10098,N_9209,N_9179);
and U10099 (N_10099,N_9119,N_9679);
nand U10100 (N_10100,N_9807,N_9291);
nor U10101 (N_10101,N_9583,N_9438);
and U10102 (N_10102,N_9127,N_9726);
nand U10103 (N_10103,N_9596,N_9902);
and U10104 (N_10104,N_9381,N_9893);
or U10105 (N_10105,N_9471,N_9000);
xor U10106 (N_10106,N_9802,N_9250);
or U10107 (N_10107,N_9587,N_9370);
nor U10108 (N_10108,N_9999,N_9375);
nand U10109 (N_10109,N_9451,N_9319);
xor U10110 (N_10110,N_9575,N_9242);
and U10111 (N_10111,N_9820,N_9949);
and U10112 (N_10112,N_9132,N_9535);
nand U10113 (N_10113,N_9085,N_9358);
nor U10114 (N_10114,N_9097,N_9576);
nor U10115 (N_10115,N_9474,N_9752);
xor U10116 (N_10116,N_9864,N_9897);
xnor U10117 (N_10117,N_9889,N_9796);
nor U10118 (N_10118,N_9149,N_9322);
nor U10119 (N_10119,N_9808,N_9162);
or U10120 (N_10120,N_9035,N_9638);
xnor U10121 (N_10121,N_9756,N_9563);
or U10122 (N_10122,N_9082,N_9278);
nor U10123 (N_10123,N_9586,N_9591);
and U10124 (N_10124,N_9970,N_9620);
nor U10125 (N_10125,N_9713,N_9075);
nand U10126 (N_10126,N_9747,N_9932);
nor U10127 (N_10127,N_9026,N_9114);
and U10128 (N_10128,N_9836,N_9282);
and U10129 (N_10129,N_9257,N_9210);
nand U10130 (N_10130,N_9649,N_9600);
nand U10131 (N_10131,N_9659,N_9868);
or U10132 (N_10132,N_9360,N_9916);
nor U10133 (N_10133,N_9666,N_9302);
nor U10134 (N_10134,N_9010,N_9505);
nor U10135 (N_10135,N_9186,N_9678);
or U10136 (N_10136,N_9266,N_9829);
nor U10137 (N_10137,N_9373,N_9616);
xnor U10138 (N_10138,N_9429,N_9589);
nor U10139 (N_10139,N_9454,N_9357);
xor U10140 (N_10140,N_9601,N_9229);
nand U10141 (N_10141,N_9495,N_9014);
xnor U10142 (N_10142,N_9885,N_9487);
and U10143 (N_10143,N_9409,N_9800);
or U10144 (N_10144,N_9749,N_9512);
xor U10145 (N_10145,N_9016,N_9066);
or U10146 (N_10146,N_9824,N_9642);
xor U10147 (N_10147,N_9632,N_9919);
nand U10148 (N_10148,N_9338,N_9544);
and U10149 (N_10149,N_9686,N_9660);
or U10150 (N_10150,N_9290,N_9550);
nand U10151 (N_10151,N_9037,N_9681);
and U10152 (N_10152,N_9274,N_9799);
or U10153 (N_10153,N_9165,N_9383);
xnor U10154 (N_10154,N_9193,N_9395);
nor U10155 (N_10155,N_9627,N_9427);
nand U10156 (N_10156,N_9402,N_9368);
nand U10157 (N_10157,N_9805,N_9452);
or U10158 (N_10158,N_9002,N_9372);
or U10159 (N_10159,N_9354,N_9072);
nor U10160 (N_10160,N_9838,N_9157);
nor U10161 (N_10161,N_9184,N_9599);
or U10162 (N_10162,N_9187,N_9767);
xor U10163 (N_10163,N_9602,N_9710);
xnor U10164 (N_10164,N_9081,N_9131);
and U10165 (N_10165,N_9674,N_9166);
or U10166 (N_10166,N_9185,N_9822);
nor U10167 (N_10167,N_9750,N_9975);
or U10168 (N_10168,N_9191,N_9736);
or U10169 (N_10169,N_9953,N_9240);
nand U10170 (N_10170,N_9175,N_9087);
nand U10171 (N_10171,N_9668,N_9387);
and U10172 (N_10172,N_9320,N_9942);
xor U10173 (N_10173,N_9239,N_9339);
and U10174 (N_10174,N_9006,N_9412);
and U10175 (N_10175,N_9911,N_9909);
and U10176 (N_10176,N_9435,N_9262);
and U10177 (N_10177,N_9561,N_9656);
xor U10178 (N_10178,N_9446,N_9245);
or U10179 (N_10179,N_9884,N_9038);
and U10180 (N_10180,N_9436,N_9390);
nor U10181 (N_10181,N_9030,N_9818);
and U10182 (N_10182,N_9098,N_9716);
nand U10183 (N_10183,N_9768,N_9309);
and U10184 (N_10184,N_9207,N_9848);
or U10185 (N_10185,N_9027,N_9948);
xor U10186 (N_10186,N_9813,N_9606);
xor U10187 (N_10187,N_9727,N_9263);
nand U10188 (N_10188,N_9554,N_9057);
nand U10189 (N_10189,N_9697,N_9513);
xor U10190 (N_10190,N_9982,N_9712);
nor U10191 (N_10191,N_9055,N_9251);
xnor U10192 (N_10192,N_9636,N_9746);
or U10193 (N_10193,N_9622,N_9832);
xor U10194 (N_10194,N_9815,N_9144);
nor U10195 (N_10195,N_9386,N_9292);
nor U10196 (N_10196,N_9134,N_9972);
or U10197 (N_10197,N_9047,N_9564);
and U10198 (N_10198,N_9914,N_9286);
and U10199 (N_10199,N_9501,N_9523);
nor U10200 (N_10200,N_9018,N_9664);
nand U10201 (N_10201,N_9102,N_9020);
and U10202 (N_10202,N_9323,N_9477);
xnor U10203 (N_10203,N_9962,N_9195);
nand U10204 (N_10204,N_9524,N_9400);
or U10205 (N_10205,N_9481,N_9056);
nor U10206 (N_10206,N_9088,N_9795);
nand U10207 (N_10207,N_9464,N_9277);
and U10208 (N_10208,N_9069,N_9757);
xnor U10209 (N_10209,N_9901,N_9219);
nor U10210 (N_10210,N_9581,N_9519);
nor U10211 (N_10211,N_9907,N_9248);
and U10212 (N_10212,N_9315,N_9176);
or U10213 (N_10213,N_9842,N_9950);
xor U10214 (N_10214,N_9742,N_9136);
nand U10215 (N_10215,N_9650,N_9778);
nand U10216 (N_10216,N_9578,N_9899);
or U10217 (N_10217,N_9203,N_9269);
and U10218 (N_10218,N_9618,N_9147);
xnor U10219 (N_10219,N_9843,N_9419);
or U10220 (N_10220,N_9817,N_9922);
xor U10221 (N_10221,N_9126,N_9514);
xnor U10222 (N_10222,N_9721,N_9480);
and U10223 (N_10223,N_9755,N_9053);
nand U10224 (N_10224,N_9521,N_9592);
nand U10225 (N_10225,N_9880,N_9019);
and U10226 (N_10226,N_9078,N_9384);
and U10227 (N_10227,N_9051,N_9971);
xnor U10228 (N_10228,N_9562,N_9508);
nor U10229 (N_10229,N_9465,N_9863);
nand U10230 (N_10230,N_9785,N_9012);
or U10231 (N_10231,N_9702,N_9977);
xor U10232 (N_10232,N_9762,N_9857);
xnor U10233 (N_10233,N_9208,N_9852);
nor U10234 (N_10234,N_9468,N_9733);
nor U10235 (N_10235,N_9952,N_9968);
nor U10236 (N_10236,N_9783,N_9784);
and U10237 (N_10237,N_9089,N_9221);
xor U10238 (N_10238,N_9173,N_9667);
nand U10239 (N_10239,N_9486,N_9048);
xnor U10240 (N_10240,N_9973,N_9385);
nand U10241 (N_10241,N_9539,N_9811);
and U10242 (N_10242,N_9672,N_9614);
nand U10243 (N_10243,N_9298,N_9244);
xor U10244 (N_10244,N_9145,N_9017);
nand U10245 (N_10245,N_9025,N_9540);
nor U10246 (N_10246,N_9118,N_9321);
xor U10247 (N_10247,N_9310,N_9156);
nor U10248 (N_10248,N_9993,N_9531);
xnor U10249 (N_10249,N_9655,N_9029);
nor U10250 (N_10250,N_9998,N_9503);
nor U10251 (N_10251,N_9715,N_9426);
and U10252 (N_10252,N_9096,N_9966);
xor U10253 (N_10253,N_9254,N_9738);
nor U10254 (N_10254,N_9683,N_9611);
nand U10255 (N_10255,N_9110,N_9912);
and U10256 (N_10256,N_9790,N_9759);
or U10257 (N_10257,N_9243,N_9718);
and U10258 (N_10258,N_9654,N_9324);
or U10259 (N_10259,N_9865,N_9485);
xor U10260 (N_10260,N_9307,N_9700);
or U10261 (N_10261,N_9517,N_9476);
and U10262 (N_10262,N_9117,N_9398);
and U10263 (N_10263,N_9645,N_9092);
xnor U10264 (N_10264,N_9124,N_9773);
xor U10265 (N_10265,N_9146,N_9719);
xor U10266 (N_10266,N_9353,N_9924);
or U10267 (N_10267,N_9913,N_9927);
or U10268 (N_10268,N_9552,N_9533);
nand U10269 (N_10269,N_9984,N_9416);
nand U10270 (N_10270,N_9760,N_9420);
nor U10271 (N_10271,N_9567,N_9293);
or U10272 (N_10272,N_9803,N_9443);
nor U10273 (N_10273,N_9687,N_9216);
nor U10274 (N_10274,N_9526,N_9624);
nor U10275 (N_10275,N_9448,N_9646);
nor U10276 (N_10276,N_9129,N_9694);
nand U10277 (N_10277,N_9270,N_9652);
nand U10278 (N_10278,N_9717,N_9873);
and U10279 (N_10279,N_9547,N_9417);
nor U10280 (N_10280,N_9036,N_9543);
or U10281 (N_10281,N_9215,N_9780);
or U10282 (N_10282,N_9439,N_9349);
or U10283 (N_10283,N_9283,N_9444);
and U10284 (N_10284,N_9794,N_9722);
nor U10285 (N_10285,N_9663,N_9895);
nand U10286 (N_10286,N_9964,N_9595);
xnor U10287 (N_10287,N_9827,N_9153);
xnor U10288 (N_10288,N_9378,N_9549);
or U10289 (N_10289,N_9731,N_9612);
or U10290 (N_10290,N_9311,N_9994);
nor U10291 (N_10291,N_9705,N_9188);
or U10292 (N_10292,N_9631,N_9137);
nand U10293 (N_10293,N_9641,N_9940);
nand U10294 (N_10294,N_9106,N_9720);
xor U10295 (N_10295,N_9930,N_9633);
or U10296 (N_10296,N_9033,N_9763);
and U10297 (N_10297,N_9676,N_9507);
and U10298 (N_10298,N_9878,N_9708);
and U10299 (N_10299,N_9174,N_9946);
nor U10300 (N_10300,N_9849,N_9986);
nand U10301 (N_10301,N_9238,N_9013);
and U10302 (N_10302,N_9299,N_9545);
or U10303 (N_10303,N_9854,N_9148);
nor U10304 (N_10304,N_9227,N_9090);
nand U10305 (N_10305,N_9682,N_9382);
or U10306 (N_10306,N_9969,N_9537);
nor U10307 (N_10307,N_9594,N_9959);
nor U10308 (N_10308,N_9723,N_9831);
and U10309 (N_10309,N_9774,N_9826);
xnor U10310 (N_10310,N_9816,N_9414);
nor U10311 (N_10311,N_9247,N_9701);
nand U10312 (N_10312,N_9192,N_9294);
nor U10313 (N_10313,N_9839,N_9289);
or U10314 (N_10314,N_9316,N_9259);
xor U10315 (N_10315,N_9121,N_9359);
nor U10316 (N_10316,N_9040,N_9054);
xor U10317 (N_10317,N_9651,N_9143);
and U10318 (N_10318,N_9809,N_9582);
and U10319 (N_10319,N_9711,N_9076);
and U10320 (N_10320,N_9333,N_9226);
or U10321 (N_10321,N_9347,N_9573);
and U10322 (N_10322,N_9833,N_9430);
nor U10323 (N_10323,N_9695,N_9511);
nand U10324 (N_10324,N_9199,N_9473);
nand U10325 (N_10325,N_9367,N_9840);
or U10326 (N_10326,N_9597,N_9167);
xor U10327 (N_10327,N_9637,N_9933);
or U10328 (N_10328,N_9935,N_9330);
nand U10329 (N_10329,N_9551,N_9022);
nand U10330 (N_10330,N_9751,N_9079);
nand U10331 (N_10331,N_9196,N_9847);
and U10332 (N_10332,N_9851,N_9571);
nor U10333 (N_10333,N_9236,N_9190);
xnor U10334 (N_10334,N_9028,N_9198);
or U10335 (N_10335,N_9272,N_9890);
or U10336 (N_10336,N_9772,N_9493);
or U10337 (N_10337,N_9990,N_9376);
or U10338 (N_10338,N_9337,N_9689);
xnor U10339 (N_10339,N_9534,N_9598);
xnor U10340 (N_10340,N_9492,N_9194);
and U10341 (N_10341,N_9279,N_9985);
xor U10342 (N_10342,N_9771,N_9059);
nor U10343 (N_10343,N_9647,N_9328);
xnor U10344 (N_10344,N_9021,N_9154);
xor U10345 (N_10345,N_9418,N_9423);
xnor U10346 (N_10346,N_9008,N_9280);
and U10347 (N_10347,N_9788,N_9335);
xor U10348 (N_10348,N_9482,N_9793);
xor U10349 (N_10349,N_9046,N_9369);
or U10350 (N_10350,N_9955,N_9392);
and U10351 (N_10351,N_9804,N_9920);
and U10352 (N_10352,N_9407,N_9108);
or U10353 (N_10353,N_9052,N_9255);
and U10354 (N_10354,N_9553,N_9334);
xnor U10355 (N_10355,N_9669,N_9812);
nand U10356 (N_10356,N_9142,N_9232);
or U10357 (N_10357,N_9061,N_9312);
nor U10358 (N_10358,N_9111,N_9639);
nor U10359 (N_10359,N_9883,N_9928);
or U10360 (N_10360,N_9249,N_9351);
or U10361 (N_10361,N_9463,N_9317);
nand U10362 (N_10362,N_9483,N_9593);
nor U10363 (N_10363,N_9393,N_9754);
nand U10364 (N_10364,N_9855,N_9590);
nor U10365 (N_10365,N_9903,N_9858);
xnor U10366 (N_10366,N_9488,N_9150);
and U10367 (N_10367,N_9542,N_9355);
nand U10368 (N_10368,N_9484,N_9995);
nor U10369 (N_10369,N_9825,N_9628);
xor U10370 (N_10370,N_9325,N_9957);
or U10371 (N_10371,N_9610,N_9031);
nor U10372 (N_10372,N_9462,N_9456);
or U10373 (N_10373,N_9870,N_9775);
and U10374 (N_10374,N_9961,N_9766);
nand U10375 (N_10375,N_9225,N_9693);
nor U10376 (N_10376,N_9388,N_9876);
nor U10377 (N_10377,N_9177,N_9653);
nor U10378 (N_10378,N_9112,N_9896);
and U10379 (N_10379,N_9877,N_9704);
or U10380 (N_10380,N_9860,N_9658);
nor U10381 (N_10381,N_9504,N_9906);
or U10382 (N_10382,N_9527,N_9529);
and U10383 (N_10383,N_9951,N_9218);
nor U10384 (N_10384,N_9004,N_9396);
or U10385 (N_10385,N_9892,N_9607);
or U10386 (N_10386,N_9261,N_9648);
xnor U10387 (N_10387,N_9967,N_9944);
or U10388 (N_10388,N_9623,N_9401);
or U10389 (N_10389,N_9206,N_9421);
xnor U10390 (N_10390,N_9692,N_9502);
xnor U10391 (N_10391,N_9005,N_9574);
xnor U10392 (N_10392,N_9447,N_9609);
nand U10393 (N_10393,N_9288,N_9898);
nor U10394 (N_10394,N_9001,N_9644);
xor U10395 (N_10395,N_9871,N_9978);
nand U10396 (N_10396,N_9141,N_9923);
or U10397 (N_10397,N_9491,N_9222);
and U10398 (N_10398,N_9980,N_9161);
xor U10399 (N_10399,N_9936,N_9212);
and U10400 (N_10400,N_9761,N_9707);
nand U10401 (N_10401,N_9801,N_9568);
nand U10402 (N_10402,N_9744,N_9518);
xnor U10403 (N_10403,N_9714,N_9116);
nand U10404 (N_10404,N_9934,N_9362);
and U10405 (N_10405,N_9963,N_9729);
and U10406 (N_10406,N_9630,N_9389);
nand U10407 (N_10407,N_9881,N_9182);
or U10408 (N_10408,N_9662,N_9728);
xor U10409 (N_10409,N_9062,N_9989);
or U10410 (N_10410,N_9015,N_9548);
nand U10411 (N_10411,N_9528,N_9745);
and U10412 (N_10412,N_9945,N_9034);
and U10413 (N_10413,N_9867,N_9276);
xor U10414 (N_10414,N_9422,N_9406);
nand U10415 (N_10415,N_9065,N_9125);
nand U10416 (N_10416,N_9556,N_9557);
xnor U10417 (N_10417,N_9861,N_9094);
nor U10418 (N_10418,N_9459,N_9361);
xor U10419 (N_10419,N_9837,N_9350);
or U10420 (N_10420,N_9415,N_9821);
xor U10421 (N_10421,N_9910,N_9122);
nor U10422 (N_10422,N_9296,N_9670);
xnor U10423 (N_10423,N_9770,N_9791);
and U10424 (N_10424,N_9882,N_9915);
nand U10425 (N_10425,N_9584,N_9084);
or U10426 (N_10426,N_9041,N_9458);
nand U10427 (N_10427,N_9580,N_9555);
nand U10428 (N_10428,N_9450,N_9925);
nand U10429 (N_10429,N_9314,N_9397);
and U10430 (N_10430,N_9009,N_9743);
nand U10431 (N_10431,N_9478,N_9941);
nor U10432 (N_10432,N_9688,N_9741);
and U10433 (N_10433,N_9163,N_9095);
nand U10434 (N_10434,N_9343,N_9170);
or U10435 (N_10435,N_9730,N_9769);
xor U10436 (N_10436,N_9180,N_9532);
nand U10437 (N_10437,N_9091,N_9905);
and U10438 (N_10438,N_9516,N_9461);
or U10439 (N_10439,N_9440,N_9758);
or U10440 (N_10440,N_9845,N_9049);
xnor U10441 (N_10441,N_9779,N_9231);
xor U10442 (N_10442,N_9405,N_9753);
nand U10443 (N_10443,N_9223,N_9128);
or U10444 (N_10444,N_9172,N_9449);
nand U10445 (N_10445,N_9133,N_9469);
nor U10446 (N_10446,N_9908,N_9947);
or U10447 (N_10447,N_9931,N_9588);
xnor U10448 (N_10448,N_9453,N_9894);
and U10449 (N_10449,N_9506,N_9295);
xnor U10450 (N_10450,N_9806,N_9991);
and U10451 (N_10451,N_9846,N_9228);
xnor U10452 (N_10452,N_9765,N_9904);
or U10453 (N_10453,N_9109,N_9428);
or U10454 (N_10454,N_9740,N_9304);
xor U10455 (N_10455,N_9886,N_9538);
nor U10456 (N_10456,N_9135,N_9617);
nand U10457 (N_10457,N_9032,N_9099);
nor U10458 (N_10458,N_9810,N_9120);
and U10459 (N_10459,N_9603,N_9171);
nand U10460 (N_10460,N_9271,N_9313);
or U10461 (N_10461,N_9565,N_9698);
nor U10462 (N_10462,N_9490,N_9217);
nand U10463 (N_10463,N_9819,N_9045);
nor U10464 (N_10464,N_9558,N_9326);
or U10465 (N_10465,N_9696,N_9608);
nor U10466 (N_10466,N_9789,N_9900);
xnor U10467 (N_10467,N_9303,N_9246);
xnor U10468 (N_10468,N_9377,N_9996);
xor U10469 (N_10469,N_9235,N_9457);
xor U10470 (N_10470,N_9441,N_9159);
nor U10471 (N_10471,N_9003,N_9252);
or U10472 (N_10472,N_9834,N_9585);
or U10473 (N_10473,N_9241,N_9830);
nand U10474 (N_10474,N_9732,N_9853);
xnor U10475 (N_10475,N_9887,N_9050);
xnor U10476 (N_10476,N_9431,N_9105);
and U10477 (N_10477,N_9498,N_9399);
or U10478 (N_10478,N_9828,N_9068);
nand U10479 (N_10479,N_9363,N_9626);
or U10480 (N_10480,N_9201,N_9494);
or U10481 (N_10481,N_9168,N_9107);
and U10482 (N_10482,N_9981,N_9160);
xnor U10483 (N_10483,N_9466,N_9093);
nor U10484 (N_10484,N_9874,N_9115);
xnor U10485 (N_10485,N_9152,N_9043);
and U10486 (N_10486,N_9260,N_9077);
nand U10487 (N_10487,N_9341,N_9425);
nor U10488 (N_10488,N_9346,N_9979);
xnor U10489 (N_10489,N_9366,N_9155);
nand U10490 (N_10490,N_9345,N_9300);
nand U10491 (N_10491,N_9605,N_9413);
xnor U10492 (N_10492,N_9178,N_9536);
nor U10493 (N_10493,N_9202,N_9327);
and U10494 (N_10494,N_9665,N_9875);
xor U10495 (N_10495,N_9011,N_9509);
and U10496 (N_10496,N_9220,N_9063);
nand U10497 (N_10497,N_9569,N_9781);
or U10498 (N_10498,N_9403,N_9570);
nor U10499 (N_10499,N_9613,N_9306);
xnor U10500 (N_10500,N_9984,N_9851);
and U10501 (N_10501,N_9999,N_9504);
and U10502 (N_10502,N_9423,N_9835);
xor U10503 (N_10503,N_9254,N_9489);
nor U10504 (N_10504,N_9160,N_9389);
xnor U10505 (N_10505,N_9284,N_9125);
xor U10506 (N_10506,N_9376,N_9023);
nor U10507 (N_10507,N_9339,N_9837);
nor U10508 (N_10508,N_9937,N_9738);
and U10509 (N_10509,N_9716,N_9244);
or U10510 (N_10510,N_9357,N_9482);
xnor U10511 (N_10511,N_9457,N_9179);
nand U10512 (N_10512,N_9985,N_9626);
nand U10513 (N_10513,N_9038,N_9573);
nor U10514 (N_10514,N_9061,N_9591);
and U10515 (N_10515,N_9969,N_9390);
and U10516 (N_10516,N_9094,N_9038);
and U10517 (N_10517,N_9013,N_9313);
xor U10518 (N_10518,N_9268,N_9246);
xnor U10519 (N_10519,N_9863,N_9865);
and U10520 (N_10520,N_9193,N_9776);
xnor U10521 (N_10521,N_9770,N_9893);
nand U10522 (N_10522,N_9621,N_9987);
xnor U10523 (N_10523,N_9152,N_9956);
xor U10524 (N_10524,N_9629,N_9532);
xnor U10525 (N_10525,N_9300,N_9274);
nand U10526 (N_10526,N_9348,N_9832);
nand U10527 (N_10527,N_9044,N_9749);
nor U10528 (N_10528,N_9645,N_9912);
or U10529 (N_10529,N_9005,N_9748);
and U10530 (N_10530,N_9981,N_9632);
and U10531 (N_10531,N_9814,N_9871);
xor U10532 (N_10532,N_9876,N_9229);
and U10533 (N_10533,N_9244,N_9073);
nor U10534 (N_10534,N_9648,N_9713);
nor U10535 (N_10535,N_9159,N_9180);
or U10536 (N_10536,N_9797,N_9079);
or U10537 (N_10537,N_9974,N_9741);
nand U10538 (N_10538,N_9408,N_9638);
and U10539 (N_10539,N_9420,N_9414);
nor U10540 (N_10540,N_9328,N_9235);
nor U10541 (N_10541,N_9017,N_9953);
and U10542 (N_10542,N_9505,N_9361);
nand U10543 (N_10543,N_9179,N_9014);
and U10544 (N_10544,N_9216,N_9890);
or U10545 (N_10545,N_9860,N_9643);
nor U10546 (N_10546,N_9132,N_9752);
or U10547 (N_10547,N_9164,N_9146);
and U10548 (N_10548,N_9609,N_9798);
or U10549 (N_10549,N_9998,N_9369);
and U10550 (N_10550,N_9814,N_9261);
nor U10551 (N_10551,N_9921,N_9147);
or U10552 (N_10552,N_9458,N_9498);
xnor U10553 (N_10553,N_9542,N_9397);
and U10554 (N_10554,N_9783,N_9614);
nand U10555 (N_10555,N_9580,N_9417);
and U10556 (N_10556,N_9140,N_9385);
and U10557 (N_10557,N_9104,N_9409);
xor U10558 (N_10558,N_9679,N_9244);
xnor U10559 (N_10559,N_9784,N_9955);
nor U10560 (N_10560,N_9316,N_9855);
or U10561 (N_10561,N_9572,N_9093);
nand U10562 (N_10562,N_9972,N_9919);
and U10563 (N_10563,N_9771,N_9379);
nor U10564 (N_10564,N_9618,N_9580);
nand U10565 (N_10565,N_9565,N_9831);
nand U10566 (N_10566,N_9699,N_9467);
and U10567 (N_10567,N_9817,N_9968);
nand U10568 (N_10568,N_9150,N_9837);
nor U10569 (N_10569,N_9037,N_9438);
nor U10570 (N_10570,N_9135,N_9120);
and U10571 (N_10571,N_9945,N_9700);
nand U10572 (N_10572,N_9262,N_9120);
or U10573 (N_10573,N_9078,N_9863);
nand U10574 (N_10574,N_9510,N_9996);
or U10575 (N_10575,N_9384,N_9233);
nor U10576 (N_10576,N_9231,N_9819);
xnor U10577 (N_10577,N_9086,N_9895);
or U10578 (N_10578,N_9321,N_9626);
and U10579 (N_10579,N_9519,N_9909);
nor U10580 (N_10580,N_9458,N_9849);
nor U10581 (N_10581,N_9222,N_9472);
nand U10582 (N_10582,N_9444,N_9713);
nand U10583 (N_10583,N_9906,N_9759);
or U10584 (N_10584,N_9690,N_9705);
xor U10585 (N_10585,N_9991,N_9036);
nand U10586 (N_10586,N_9540,N_9291);
nor U10587 (N_10587,N_9835,N_9004);
nand U10588 (N_10588,N_9778,N_9961);
nor U10589 (N_10589,N_9497,N_9682);
or U10590 (N_10590,N_9330,N_9975);
xnor U10591 (N_10591,N_9687,N_9430);
nor U10592 (N_10592,N_9851,N_9180);
nor U10593 (N_10593,N_9489,N_9042);
xor U10594 (N_10594,N_9136,N_9610);
nand U10595 (N_10595,N_9050,N_9784);
nor U10596 (N_10596,N_9328,N_9091);
nand U10597 (N_10597,N_9511,N_9710);
and U10598 (N_10598,N_9325,N_9610);
nor U10599 (N_10599,N_9994,N_9496);
nand U10600 (N_10600,N_9829,N_9872);
nand U10601 (N_10601,N_9558,N_9778);
and U10602 (N_10602,N_9420,N_9131);
nand U10603 (N_10603,N_9587,N_9943);
xor U10604 (N_10604,N_9981,N_9813);
nand U10605 (N_10605,N_9840,N_9807);
or U10606 (N_10606,N_9952,N_9243);
and U10607 (N_10607,N_9359,N_9593);
nand U10608 (N_10608,N_9567,N_9525);
or U10609 (N_10609,N_9060,N_9026);
xor U10610 (N_10610,N_9152,N_9666);
nor U10611 (N_10611,N_9609,N_9018);
nor U10612 (N_10612,N_9594,N_9550);
or U10613 (N_10613,N_9770,N_9399);
xor U10614 (N_10614,N_9201,N_9644);
xnor U10615 (N_10615,N_9422,N_9463);
nor U10616 (N_10616,N_9353,N_9211);
and U10617 (N_10617,N_9949,N_9445);
nand U10618 (N_10618,N_9360,N_9163);
xnor U10619 (N_10619,N_9392,N_9126);
nand U10620 (N_10620,N_9180,N_9229);
or U10621 (N_10621,N_9176,N_9911);
nand U10622 (N_10622,N_9380,N_9357);
xor U10623 (N_10623,N_9915,N_9107);
xor U10624 (N_10624,N_9069,N_9475);
or U10625 (N_10625,N_9609,N_9834);
nand U10626 (N_10626,N_9045,N_9860);
nor U10627 (N_10627,N_9267,N_9835);
xnor U10628 (N_10628,N_9400,N_9038);
nand U10629 (N_10629,N_9067,N_9329);
xnor U10630 (N_10630,N_9262,N_9489);
and U10631 (N_10631,N_9291,N_9266);
nor U10632 (N_10632,N_9167,N_9762);
xnor U10633 (N_10633,N_9644,N_9454);
or U10634 (N_10634,N_9392,N_9684);
nor U10635 (N_10635,N_9962,N_9939);
xnor U10636 (N_10636,N_9123,N_9539);
nor U10637 (N_10637,N_9849,N_9974);
xor U10638 (N_10638,N_9491,N_9237);
xnor U10639 (N_10639,N_9023,N_9355);
nand U10640 (N_10640,N_9244,N_9290);
nor U10641 (N_10641,N_9796,N_9322);
nor U10642 (N_10642,N_9698,N_9412);
xor U10643 (N_10643,N_9654,N_9900);
or U10644 (N_10644,N_9657,N_9820);
or U10645 (N_10645,N_9805,N_9351);
or U10646 (N_10646,N_9779,N_9878);
or U10647 (N_10647,N_9321,N_9001);
xnor U10648 (N_10648,N_9319,N_9254);
nand U10649 (N_10649,N_9956,N_9693);
xor U10650 (N_10650,N_9309,N_9334);
or U10651 (N_10651,N_9836,N_9075);
nand U10652 (N_10652,N_9988,N_9003);
nor U10653 (N_10653,N_9634,N_9129);
or U10654 (N_10654,N_9445,N_9264);
nor U10655 (N_10655,N_9528,N_9510);
or U10656 (N_10656,N_9084,N_9387);
xor U10657 (N_10657,N_9666,N_9447);
nand U10658 (N_10658,N_9445,N_9962);
or U10659 (N_10659,N_9339,N_9675);
xnor U10660 (N_10660,N_9375,N_9527);
nor U10661 (N_10661,N_9758,N_9183);
and U10662 (N_10662,N_9043,N_9884);
and U10663 (N_10663,N_9802,N_9715);
nand U10664 (N_10664,N_9562,N_9662);
nand U10665 (N_10665,N_9112,N_9855);
nor U10666 (N_10666,N_9141,N_9850);
or U10667 (N_10667,N_9715,N_9208);
nor U10668 (N_10668,N_9137,N_9440);
xor U10669 (N_10669,N_9487,N_9726);
nand U10670 (N_10670,N_9936,N_9228);
xor U10671 (N_10671,N_9437,N_9921);
or U10672 (N_10672,N_9621,N_9273);
xnor U10673 (N_10673,N_9591,N_9574);
and U10674 (N_10674,N_9235,N_9380);
nor U10675 (N_10675,N_9052,N_9189);
or U10676 (N_10676,N_9869,N_9149);
xor U10677 (N_10677,N_9235,N_9790);
nand U10678 (N_10678,N_9840,N_9222);
nor U10679 (N_10679,N_9806,N_9851);
and U10680 (N_10680,N_9864,N_9033);
or U10681 (N_10681,N_9139,N_9911);
and U10682 (N_10682,N_9188,N_9748);
nand U10683 (N_10683,N_9602,N_9665);
nand U10684 (N_10684,N_9676,N_9111);
xor U10685 (N_10685,N_9771,N_9924);
or U10686 (N_10686,N_9684,N_9996);
xor U10687 (N_10687,N_9349,N_9428);
xnor U10688 (N_10688,N_9486,N_9758);
or U10689 (N_10689,N_9209,N_9854);
nand U10690 (N_10690,N_9049,N_9276);
nor U10691 (N_10691,N_9316,N_9185);
xor U10692 (N_10692,N_9735,N_9071);
or U10693 (N_10693,N_9489,N_9113);
and U10694 (N_10694,N_9521,N_9103);
nor U10695 (N_10695,N_9221,N_9291);
nor U10696 (N_10696,N_9854,N_9551);
or U10697 (N_10697,N_9284,N_9374);
nand U10698 (N_10698,N_9960,N_9276);
xnor U10699 (N_10699,N_9112,N_9190);
or U10700 (N_10700,N_9361,N_9190);
nand U10701 (N_10701,N_9017,N_9286);
and U10702 (N_10702,N_9089,N_9604);
and U10703 (N_10703,N_9357,N_9842);
nor U10704 (N_10704,N_9414,N_9098);
nand U10705 (N_10705,N_9638,N_9732);
xnor U10706 (N_10706,N_9682,N_9692);
xor U10707 (N_10707,N_9649,N_9365);
and U10708 (N_10708,N_9338,N_9356);
nor U10709 (N_10709,N_9460,N_9192);
nand U10710 (N_10710,N_9832,N_9440);
and U10711 (N_10711,N_9517,N_9977);
xor U10712 (N_10712,N_9193,N_9828);
xnor U10713 (N_10713,N_9411,N_9607);
or U10714 (N_10714,N_9246,N_9185);
xnor U10715 (N_10715,N_9881,N_9567);
xnor U10716 (N_10716,N_9730,N_9053);
nand U10717 (N_10717,N_9957,N_9472);
xnor U10718 (N_10718,N_9776,N_9289);
nor U10719 (N_10719,N_9298,N_9393);
or U10720 (N_10720,N_9760,N_9905);
or U10721 (N_10721,N_9676,N_9389);
nor U10722 (N_10722,N_9233,N_9662);
and U10723 (N_10723,N_9147,N_9699);
xnor U10724 (N_10724,N_9967,N_9725);
or U10725 (N_10725,N_9221,N_9082);
nor U10726 (N_10726,N_9708,N_9428);
and U10727 (N_10727,N_9868,N_9166);
xor U10728 (N_10728,N_9866,N_9852);
and U10729 (N_10729,N_9909,N_9448);
nor U10730 (N_10730,N_9303,N_9338);
and U10731 (N_10731,N_9371,N_9131);
and U10732 (N_10732,N_9561,N_9004);
nor U10733 (N_10733,N_9926,N_9058);
xor U10734 (N_10734,N_9040,N_9333);
nand U10735 (N_10735,N_9597,N_9261);
xor U10736 (N_10736,N_9587,N_9706);
xnor U10737 (N_10737,N_9243,N_9453);
xor U10738 (N_10738,N_9822,N_9575);
or U10739 (N_10739,N_9230,N_9019);
xnor U10740 (N_10740,N_9229,N_9158);
xnor U10741 (N_10741,N_9524,N_9750);
and U10742 (N_10742,N_9655,N_9593);
nor U10743 (N_10743,N_9848,N_9997);
nor U10744 (N_10744,N_9108,N_9544);
or U10745 (N_10745,N_9683,N_9536);
nor U10746 (N_10746,N_9923,N_9324);
xnor U10747 (N_10747,N_9005,N_9420);
nand U10748 (N_10748,N_9771,N_9633);
and U10749 (N_10749,N_9904,N_9163);
nand U10750 (N_10750,N_9807,N_9187);
xnor U10751 (N_10751,N_9844,N_9117);
nand U10752 (N_10752,N_9137,N_9257);
nand U10753 (N_10753,N_9762,N_9586);
xnor U10754 (N_10754,N_9901,N_9747);
xnor U10755 (N_10755,N_9334,N_9833);
xor U10756 (N_10756,N_9066,N_9269);
and U10757 (N_10757,N_9844,N_9538);
nor U10758 (N_10758,N_9037,N_9792);
nand U10759 (N_10759,N_9505,N_9563);
or U10760 (N_10760,N_9602,N_9264);
nand U10761 (N_10761,N_9652,N_9123);
xnor U10762 (N_10762,N_9676,N_9762);
or U10763 (N_10763,N_9637,N_9695);
and U10764 (N_10764,N_9676,N_9546);
or U10765 (N_10765,N_9985,N_9804);
xnor U10766 (N_10766,N_9658,N_9820);
nor U10767 (N_10767,N_9975,N_9307);
xor U10768 (N_10768,N_9739,N_9560);
or U10769 (N_10769,N_9998,N_9329);
nand U10770 (N_10770,N_9059,N_9547);
nand U10771 (N_10771,N_9582,N_9312);
nor U10772 (N_10772,N_9971,N_9873);
and U10773 (N_10773,N_9457,N_9982);
nand U10774 (N_10774,N_9578,N_9721);
xnor U10775 (N_10775,N_9646,N_9511);
nand U10776 (N_10776,N_9374,N_9198);
nand U10777 (N_10777,N_9869,N_9089);
and U10778 (N_10778,N_9769,N_9202);
nor U10779 (N_10779,N_9313,N_9363);
nor U10780 (N_10780,N_9391,N_9220);
and U10781 (N_10781,N_9209,N_9477);
nand U10782 (N_10782,N_9145,N_9133);
xor U10783 (N_10783,N_9820,N_9021);
and U10784 (N_10784,N_9230,N_9978);
nand U10785 (N_10785,N_9254,N_9695);
nand U10786 (N_10786,N_9445,N_9159);
and U10787 (N_10787,N_9323,N_9811);
and U10788 (N_10788,N_9671,N_9518);
xnor U10789 (N_10789,N_9155,N_9825);
and U10790 (N_10790,N_9641,N_9467);
nand U10791 (N_10791,N_9028,N_9242);
and U10792 (N_10792,N_9851,N_9469);
nand U10793 (N_10793,N_9735,N_9704);
xor U10794 (N_10794,N_9365,N_9065);
xor U10795 (N_10795,N_9779,N_9010);
xnor U10796 (N_10796,N_9999,N_9526);
or U10797 (N_10797,N_9507,N_9703);
nand U10798 (N_10798,N_9290,N_9266);
nor U10799 (N_10799,N_9232,N_9650);
or U10800 (N_10800,N_9697,N_9169);
nor U10801 (N_10801,N_9610,N_9035);
and U10802 (N_10802,N_9361,N_9903);
nand U10803 (N_10803,N_9950,N_9766);
xnor U10804 (N_10804,N_9903,N_9983);
xnor U10805 (N_10805,N_9434,N_9208);
xor U10806 (N_10806,N_9906,N_9639);
or U10807 (N_10807,N_9553,N_9942);
and U10808 (N_10808,N_9564,N_9227);
nor U10809 (N_10809,N_9853,N_9128);
or U10810 (N_10810,N_9725,N_9902);
and U10811 (N_10811,N_9219,N_9512);
and U10812 (N_10812,N_9487,N_9295);
nor U10813 (N_10813,N_9918,N_9255);
nand U10814 (N_10814,N_9870,N_9575);
or U10815 (N_10815,N_9414,N_9035);
nor U10816 (N_10816,N_9459,N_9551);
xor U10817 (N_10817,N_9535,N_9839);
nand U10818 (N_10818,N_9867,N_9553);
and U10819 (N_10819,N_9942,N_9601);
and U10820 (N_10820,N_9957,N_9551);
or U10821 (N_10821,N_9301,N_9979);
nor U10822 (N_10822,N_9117,N_9541);
nor U10823 (N_10823,N_9525,N_9277);
nand U10824 (N_10824,N_9173,N_9422);
nand U10825 (N_10825,N_9520,N_9720);
nand U10826 (N_10826,N_9900,N_9489);
nand U10827 (N_10827,N_9997,N_9231);
nand U10828 (N_10828,N_9187,N_9848);
nor U10829 (N_10829,N_9841,N_9006);
nor U10830 (N_10830,N_9526,N_9867);
or U10831 (N_10831,N_9586,N_9639);
nor U10832 (N_10832,N_9482,N_9821);
nand U10833 (N_10833,N_9919,N_9333);
nor U10834 (N_10834,N_9919,N_9045);
nand U10835 (N_10835,N_9857,N_9375);
nand U10836 (N_10836,N_9623,N_9691);
xor U10837 (N_10837,N_9192,N_9430);
nand U10838 (N_10838,N_9657,N_9397);
xnor U10839 (N_10839,N_9156,N_9161);
and U10840 (N_10840,N_9856,N_9365);
nor U10841 (N_10841,N_9498,N_9098);
xnor U10842 (N_10842,N_9783,N_9063);
nand U10843 (N_10843,N_9771,N_9906);
nor U10844 (N_10844,N_9415,N_9348);
and U10845 (N_10845,N_9423,N_9411);
nor U10846 (N_10846,N_9805,N_9001);
and U10847 (N_10847,N_9904,N_9040);
or U10848 (N_10848,N_9760,N_9892);
or U10849 (N_10849,N_9618,N_9409);
nor U10850 (N_10850,N_9984,N_9934);
or U10851 (N_10851,N_9564,N_9070);
nand U10852 (N_10852,N_9330,N_9765);
nor U10853 (N_10853,N_9774,N_9208);
or U10854 (N_10854,N_9202,N_9627);
nor U10855 (N_10855,N_9958,N_9396);
nand U10856 (N_10856,N_9454,N_9219);
xor U10857 (N_10857,N_9363,N_9916);
xnor U10858 (N_10858,N_9244,N_9813);
nor U10859 (N_10859,N_9606,N_9823);
xnor U10860 (N_10860,N_9508,N_9733);
xor U10861 (N_10861,N_9416,N_9044);
and U10862 (N_10862,N_9086,N_9789);
nor U10863 (N_10863,N_9073,N_9495);
nand U10864 (N_10864,N_9487,N_9069);
or U10865 (N_10865,N_9992,N_9943);
xnor U10866 (N_10866,N_9996,N_9860);
nand U10867 (N_10867,N_9649,N_9539);
xnor U10868 (N_10868,N_9967,N_9524);
and U10869 (N_10869,N_9614,N_9673);
or U10870 (N_10870,N_9814,N_9402);
and U10871 (N_10871,N_9235,N_9171);
or U10872 (N_10872,N_9944,N_9621);
xnor U10873 (N_10873,N_9727,N_9747);
xnor U10874 (N_10874,N_9817,N_9039);
or U10875 (N_10875,N_9949,N_9352);
nor U10876 (N_10876,N_9101,N_9643);
or U10877 (N_10877,N_9567,N_9730);
or U10878 (N_10878,N_9213,N_9166);
nor U10879 (N_10879,N_9088,N_9862);
and U10880 (N_10880,N_9986,N_9784);
or U10881 (N_10881,N_9630,N_9366);
xor U10882 (N_10882,N_9650,N_9954);
nand U10883 (N_10883,N_9325,N_9145);
or U10884 (N_10884,N_9251,N_9598);
or U10885 (N_10885,N_9574,N_9488);
and U10886 (N_10886,N_9516,N_9008);
xor U10887 (N_10887,N_9639,N_9094);
xor U10888 (N_10888,N_9986,N_9392);
xor U10889 (N_10889,N_9911,N_9037);
or U10890 (N_10890,N_9429,N_9756);
or U10891 (N_10891,N_9091,N_9491);
xor U10892 (N_10892,N_9391,N_9758);
nor U10893 (N_10893,N_9373,N_9755);
nand U10894 (N_10894,N_9056,N_9107);
xnor U10895 (N_10895,N_9407,N_9235);
and U10896 (N_10896,N_9608,N_9530);
or U10897 (N_10897,N_9125,N_9742);
and U10898 (N_10898,N_9696,N_9939);
and U10899 (N_10899,N_9235,N_9808);
and U10900 (N_10900,N_9477,N_9282);
nor U10901 (N_10901,N_9055,N_9119);
nand U10902 (N_10902,N_9826,N_9542);
xor U10903 (N_10903,N_9196,N_9531);
or U10904 (N_10904,N_9806,N_9474);
or U10905 (N_10905,N_9301,N_9555);
xor U10906 (N_10906,N_9134,N_9649);
nor U10907 (N_10907,N_9259,N_9930);
or U10908 (N_10908,N_9639,N_9073);
nand U10909 (N_10909,N_9328,N_9643);
and U10910 (N_10910,N_9464,N_9002);
xnor U10911 (N_10911,N_9712,N_9697);
nand U10912 (N_10912,N_9671,N_9841);
or U10913 (N_10913,N_9174,N_9652);
or U10914 (N_10914,N_9714,N_9829);
xnor U10915 (N_10915,N_9786,N_9234);
and U10916 (N_10916,N_9513,N_9358);
and U10917 (N_10917,N_9361,N_9325);
xor U10918 (N_10918,N_9382,N_9641);
xor U10919 (N_10919,N_9221,N_9542);
or U10920 (N_10920,N_9831,N_9380);
nand U10921 (N_10921,N_9683,N_9334);
or U10922 (N_10922,N_9209,N_9652);
xor U10923 (N_10923,N_9219,N_9642);
xor U10924 (N_10924,N_9276,N_9626);
or U10925 (N_10925,N_9228,N_9191);
nand U10926 (N_10926,N_9913,N_9906);
and U10927 (N_10927,N_9895,N_9844);
or U10928 (N_10928,N_9823,N_9966);
nand U10929 (N_10929,N_9815,N_9728);
nor U10930 (N_10930,N_9764,N_9156);
or U10931 (N_10931,N_9839,N_9744);
and U10932 (N_10932,N_9389,N_9447);
nor U10933 (N_10933,N_9053,N_9734);
and U10934 (N_10934,N_9742,N_9266);
or U10935 (N_10935,N_9938,N_9543);
and U10936 (N_10936,N_9885,N_9546);
xnor U10937 (N_10937,N_9838,N_9070);
nand U10938 (N_10938,N_9038,N_9850);
or U10939 (N_10939,N_9793,N_9354);
xnor U10940 (N_10940,N_9014,N_9358);
and U10941 (N_10941,N_9440,N_9957);
nand U10942 (N_10942,N_9274,N_9314);
xnor U10943 (N_10943,N_9264,N_9186);
or U10944 (N_10944,N_9898,N_9976);
nand U10945 (N_10945,N_9770,N_9615);
xor U10946 (N_10946,N_9706,N_9491);
nand U10947 (N_10947,N_9757,N_9901);
xor U10948 (N_10948,N_9711,N_9865);
and U10949 (N_10949,N_9371,N_9003);
nor U10950 (N_10950,N_9035,N_9257);
and U10951 (N_10951,N_9978,N_9303);
nand U10952 (N_10952,N_9428,N_9506);
nand U10953 (N_10953,N_9017,N_9774);
or U10954 (N_10954,N_9857,N_9622);
or U10955 (N_10955,N_9410,N_9321);
and U10956 (N_10956,N_9927,N_9275);
xnor U10957 (N_10957,N_9456,N_9240);
or U10958 (N_10958,N_9167,N_9571);
nor U10959 (N_10959,N_9536,N_9243);
or U10960 (N_10960,N_9095,N_9827);
nand U10961 (N_10961,N_9147,N_9140);
and U10962 (N_10962,N_9831,N_9134);
nand U10963 (N_10963,N_9231,N_9574);
and U10964 (N_10964,N_9489,N_9278);
or U10965 (N_10965,N_9419,N_9267);
xor U10966 (N_10966,N_9524,N_9838);
nor U10967 (N_10967,N_9628,N_9736);
and U10968 (N_10968,N_9659,N_9413);
nand U10969 (N_10969,N_9749,N_9117);
nor U10970 (N_10970,N_9163,N_9034);
nand U10971 (N_10971,N_9028,N_9581);
nand U10972 (N_10972,N_9351,N_9128);
or U10973 (N_10973,N_9597,N_9589);
xor U10974 (N_10974,N_9044,N_9837);
nand U10975 (N_10975,N_9381,N_9328);
xor U10976 (N_10976,N_9898,N_9732);
xnor U10977 (N_10977,N_9358,N_9096);
and U10978 (N_10978,N_9449,N_9736);
or U10979 (N_10979,N_9060,N_9595);
or U10980 (N_10980,N_9866,N_9981);
nor U10981 (N_10981,N_9715,N_9392);
and U10982 (N_10982,N_9847,N_9789);
nand U10983 (N_10983,N_9323,N_9429);
nand U10984 (N_10984,N_9398,N_9472);
nor U10985 (N_10985,N_9188,N_9838);
nand U10986 (N_10986,N_9699,N_9979);
or U10987 (N_10987,N_9319,N_9753);
and U10988 (N_10988,N_9595,N_9805);
and U10989 (N_10989,N_9532,N_9244);
and U10990 (N_10990,N_9558,N_9445);
and U10991 (N_10991,N_9905,N_9478);
and U10992 (N_10992,N_9257,N_9518);
xnor U10993 (N_10993,N_9984,N_9346);
or U10994 (N_10994,N_9495,N_9094);
nor U10995 (N_10995,N_9737,N_9257);
xor U10996 (N_10996,N_9693,N_9402);
nor U10997 (N_10997,N_9700,N_9706);
and U10998 (N_10998,N_9732,N_9870);
xnor U10999 (N_10999,N_9783,N_9374);
xnor U11000 (N_11000,N_10927,N_10813);
nand U11001 (N_11001,N_10482,N_10791);
nor U11002 (N_11002,N_10284,N_10078);
and U11003 (N_11003,N_10135,N_10553);
nor U11004 (N_11004,N_10726,N_10441);
nor U11005 (N_11005,N_10668,N_10365);
nand U11006 (N_11006,N_10091,N_10342);
and U11007 (N_11007,N_10866,N_10196);
xnor U11008 (N_11008,N_10988,N_10179);
xnor U11009 (N_11009,N_10444,N_10037);
or U11010 (N_11010,N_10887,N_10508);
and U11011 (N_11011,N_10189,N_10242);
xor U11012 (N_11012,N_10624,N_10157);
xor U11013 (N_11013,N_10190,N_10671);
nand U11014 (N_11014,N_10908,N_10042);
nor U11015 (N_11015,N_10236,N_10522);
and U11016 (N_11016,N_10292,N_10552);
nand U11017 (N_11017,N_10298,N_10654);
or U11018 (N_11018,N_10776,N_10960);
nor U11019 (N_11019,N_10762,N_10899);
nor U11020 (N_11020,N_10275,N_10399);
xnor U11021 (N_11021,N_10372,N_10529);
xnor U11022 (N_11022,N_10660,N_10808);
and U11023 (N_11023,N_10128,N_10559);
or U11024 (N_11024,N_10005,N_10652);
nand U11025 (N_11025,N_10537,N_10056);
xnor U11026 (N_11026,N_10006,N_10132);
xor U11027 (N_11027,N_10035,N_10356);
nand U11028 (N_11028,N_10423,N_10057);
and U11029 (N_11029,N_10304,N_10289);
nor U11030 (N_11030,N_10391,N_10947);
nor U11031 (N_11031,N_10390,N_10259);
nand U11032 (N_11032,N_10402,N_10421);
nor U11033 (N_11033,N_10985,N_10212);
nand U11034 (N_11034,N_10566,N_10975);
nor U11035 (N_11035,N_10587,N_10069);
nor U11036 (N_11036,N_10119,N_10570);
nor U11037 (N_11037,N_10155,N_10892);
xor U11038 (N_11038,N_10928,N_10574);
xor U11039 (N_11039,N_10807,N_10987);
nand U11040 (N_11040,N_10471,N_10353);
xor U11041 (N_11041,N_10505,N_10407);
and U11042 (N_11042,N_10816,N_10296);
nor U11043 (N_11043,N_10572,N_10516);
xnor U11044 (N_11044,N_10613,N_10691);
and U11045 (N_11045,N_10163,N_10503);
xor U11046 (N_11046,N_10713,N_10653);
or U11047 (N_11047,N_10938,N_10601);
nor U11048 (N_11048,N_10456,N_10067);
and U11049 (N_11049,N_10405,N_10327);
and U11050 (N_11050,N_10533,N_10578);
nand U11051 (N_11051,N_10074,N_10008);
nor U11052 (N_11052,N_10358,N_10090);
nand U11053 (N_11053,N_10707,N_10571);
xnor U11054 (N_11054,N_10350,N_10429);
nor U11055 (N_11055,N_10095,N_10281);
and U11056 (N_11056,N_10959,N_10945);
nand U11057 (N_11057,N_10513,N_10962);
nand U11058 (N_11058,N_10605,N_10766);
or U11059 (N_11059,N_10100,N_10568);
and U11060 (N_11060,N_10002,N_10169);
and U11061 (N_11061,N_10877,N_10715);
nand U11062 (N_11062,N_10794,N_10337);
xor U11063 (N_11063,N_10839,N_10434);
nand U11064 (N_11064,N_10741,N_10207);
and U11065 (N_11065,N_10549,N_10502);
nand U11066 (N_11066,N_10079,N_10528);
nor U11067 (N_11067,N_10158,N_10428);
nor U11068 (N_11068,N_10795,N_10895);
nand U11069 (N_11069,N_10385,N_10396);
xnor U11070 (N_11070,N_10708,N_10573);
xor U11071 (N_11071,N_10114,N_10956);
xor U11072 (N_11072,N_10551,N_10115);
xnor U11073 (N_11073,N_10021,N_10027);
or U11074 (N_11074,N_10483,N_10595);
or U11075 (N_11075,N_10799,N_10501);
nor U11076 (N_11076,N_10285,N_10151);
and U11077 (N_11077,N_10053,N_10581);
nor U11078 (N_11078,N_10834,N_10847);
and U11079 (N_11079,N_10140,N_10519);
xnor U11080 (N_11080,N_10742,N_10393);
xnor U11081 (N_11081,N_10036,N_10911);
and U11082 (N_11082,N_10981,N_10097);
nand U11083 (N_11083,N_10739,N_10958);
and U11084 (N_11084,N_10143,N_10267);
or U11085 (N_11085,N_10137,N_10585);
xnor U11086 (N_11086,N_10066,N_10303);
xnor U11087 (N_11087,N_10200,N_10355);
nor U11088 (N_11088,N_10125,N_10449);
and U11089 (N_11089,N_10345,N_10375);
or U11090 (N_11090,N_10884,N_10332);
xnor U11091 (N_11091,N_10844,N_10065);
and U11092 (N_11092,N_10435,N_10073);
xnor U11093 (N_11093,N_10917,N_10558);
and U11094 (N_11094,N_10093,N_10469);
and U11095 (N_11095,N_10828,N_10142);
and U11096 (N_11096,N_10545,N_10362);
and U11097 (N_11097,N_10782,N_10602);
or U11098 (N_11098,N_10769,N_10584);
or U11099 (N_11099,N_10670,N_10403);
nor U11100 (N_11100,N_10809,N_10491);
or U11101 (N_11101,N_10961,N_10367);
nand U11102 (N_11102,N_10420,N_10862);
or U11103 (N_11103,N_10339,N_10951);
and U11104 (N_11104,N_10175,N_10824);
and U11105 (N_11105,N_10630,N_10563);
nand U11106 (N_11106,N_10986,N_10171);
or U11107 (N_11107,N_10481,N_10751);
or U11108 (N_11108,N_10667,N_10359);
or U11109 (N_11109,N_10278,N_10397);
and U11110 (N_11110,N_10145,N_10431);
and U11111 (N_11111,N_10025,N_10437);
nor U11112 (N_11112,N_10920,N_10736);
xor U11113 (N_11113,N_10392,N_10673);
xnor U11114 (N_11114,N_10044,N_10024);
xnor U11115 (N_11115,N_10215,N_10229);
or U11116 (N_11116,N_10855,N_10937);
xor U11117 (N_11117,N_10310,N_10497);
xnor U11118 (N_11118,N_10973,N_10634);
and U11119 (N_11119,N_10850,N_10110);
and U11120 (N_11120,N_10331,N_10156);
nor U11121 (N_11121,N_10922,N_10546);
nand U11122 (N_11122,N_10188,N_10849);
or U11123 (N_11123,N_10493,N_10354);
nor U11124 (N_11124,N_10820,N_10120);
nor U11125 (N_11125,N_10206,N_10295);
nand U11126 (N_11126,N_10216,N_10705);
or U11127 (N_11127,N_10921,N_10580);
xor U11128 (N_11128,N_10604,N_10525);
and U11129 (N_11129,N_10576,N_10647);
nand U11130 (N_11130,N_10279,N_10783);
xnor U11131 (N_11131,N_10245,N_10489);
nand U11132 (N_11132,N_10357,N_10733);
nor U11133 (N_11133,N_10796,N_10623);
nor U11134 (N_11134,N_10092,N_10521);
nor U11135 (N_11135,N_10931,N_10617);
nor U11136 (N_11136,N_10637,N_10363);
xor U11137 (N_11137,N_10979,N_10217);
nand U11138 (N_11138,N_10022,N_10995);
or U11139 (N_11139,N_10648,N_10832);
xnor U11140 (N_11140,N_10082,N_10124);
nor U11141 (N_11141,N_10523,N_10954);
nor U11142 (N_11142,N_10257,N_10837);
nand U11143 (N_11143,N_10386,N_10544);
nand U11144 (N_11144,N_10925,N_10107);
nor U11145 (N_11145,N_10511,N_10717);
nor U11146 (N_11146,N_10108,N_10470);
or U11147 (N_11147,N_10994,N_10014);
and U11148 (N_11148,N_10841,N_10174);
and U11149 (N_11149,N_10643,N_10658);
xor U11150 (N_11150,N_10038,N_10699);
and U11151 (N_11151,N_10184,N_10395);
nor U11152 (N_11152,N_10440,N_10308);
nand U11153 (N_11153,N_10446,N_10896);
nor U11154 (N_11154,N_10336,N_10848);
nor U11155 (N_11155,N_10371,N_10790);
xor U11156 (N_11156,N_10910,N_10288);
or U11157 (N_11157,N_10116,N_10556);
xnor U11158 (N_11158,N_10182,N_10944);
nor U11159 (N_11159,N_10716,N_10348);
nor U11160 (N_11160,N_10721,N_10514);
or U11161 (N_11161,N_10205,N_10104);
xnor U11162 (N_11162,N_10183,N_10260);
nand U11163 (N_11163,N_10166,N_10055);
nand U11164 (N_11164,N_10784,N_10023);
nand U11165 (N_11165,N_10932,N_10133);
nand U11166 (N_11166,N_10870,N_10315);
or U11167 (N_11167,N_10261,N_10881);
nor U11168 (N_11168,N_10464,N_10948);
xor U11169 (N_11169,N_10088,N_10126);
or U11170 (N_11170,N_10661,N_10302);
or U11171 (N_11171,N_10187,N_10684);
and U11172 (N_11172,N_10086,N_10410);
xor U11173 (N_11173,N_10377,N_10461);
xnor U11174 (N_11174,N_10010,N_10659);
xor U11175 (N_11175,N_10787,N_10270);
or U11176 (N_11176,N_10081,N_10062);
nor U11177 (N_11177,N_10480,N_10603);
or U11178 (N_11178,N_10111,N_10876);
or U11179 (N_11179,N_10248,N_10968);
or U11180 (N_11180,N_10221,N_10230);
and U11181 (N_11181,N_10639,N_10477);
nand U11182 (N_11182,N_10180,N_10577);
xnor U11183 (N_11183,N_10129,N_10131);
or U11184 (N_11184,N_10101,N_10467);
nand U11185 (N_11185,N_10665,N_10294);
or U11186 (N_11186,N_10411,N_10775);
or U11187 (N_11187,N_10527,N_10340);
nand U11188 (N_11188,N_10413,N_10389);
or U11189 (N_11189,N_10814,N_10700);
and U11190 (N_11190,N_10192,N_10687);
and U11191 (N_11191,N_10490,N_10902);
nor U11192 (N_11192,N_10746,N_10498);
nand U11193 (N_11193,N_10176,N_10380);
nand U11194 (N_11194,N_10701,N_10983);
or U11195 (N_11195,N_10621,N_10596);
and U11196 (N_11196,N_10743,N_10510);
nand U11197 (N_11197,N_10406,N_10426);
nor U11198 (N_11198,N_10299,N_10879);
nor U11199 (N_11199,N_10934,N_10494);
or U11200 (N_11200,N_10277,N_10905);
xor U11201 (N_11201,N_10843,N_10136);
and U11202 (N_11202,N_10823,N_10812);
nand U11203 (N_11203,N_10840,N_10851);
and U11204 (N_11204,N_10589,N_10636);
xnor U11205 (N_11205,N_10955,N_10509);
or U11206 (N_11206,N_10773,N_10015);
or U11207 (N_11207,N_10462,N_10352);
xor U11208 (N_11208,N_10492,N_10641);
nand U11209 (N_11209,N_10400,N_10152);
and U11210 (N_11210,N_10451,N_10874);
xor U11211 (N_11211,N_10990,N_10520);
xnor U11212 (N_11212,N_10307,N_10496);
nand U11213 (N_11213,N_10518,N_10821);
nor U11214 (N_11214,N_10201,N_10320);
nor U11215 (N_11215,N_10677,N_10982);
nor U11216 (N_11216,N_10054,N_10535);
nor U11217 (N_11217,N_10117,N_10838);
nand U11218 (N_11218,N_10225,N_10802);
or U11219 (N_11219,N_10121,N_10542);
xnor U11220 (N_11220,N_10744,N_10311);
and U11221 (N_11221,N_10424,N_10416);
and U11222 (N_11222,N_10476,N_10153);
nand U11223 (N_11223,N_10657,N_10040);
xnor U11224 (N_11224,N_10702,N_10341);
and U11225 (N_11225,N_10329,N_10745);
nor U11226 (N_11226,N_10239,N_10723);
or U11227 (N_11227,N_10147,N_10436);
and U11228 (N_11228,N_10422,N_10919);
and U11229 (N_11229,N_10709,N_10439);
xor U11230 (N_11230,N_10974,N_10728);
nand U11231 (N_11231,N_10692,N_10072);
xnor U11232 (N_11232,N_10629,N_10999);
or U11233 (N_11233,N_10417,N_10050);
xor U11234 (N_11234,N_10255,N_10250);
or U11235 (N_11235,N_10051,N_10433);
or U11236 (N_11236,N_10018,N_10912);
nand U11237 (N_11237,N_10077,N_10244);
and U11238 (N_11238,N_10083,N_10419);
nor U11239 (N_11239,N_10651,N_10247);
and U11240 (N_11240,N_10758,N_10254);
and U11241 (N_11241,N_10076,N_10532);
or U11242 (N_11242,N_10594,N_10202);
and U11243 (N_11243,N_10878,N_10548);
or U11244 (N_11244,N_10941,N_10852);
and U11245 (N_11245,N_10068,N_10645);
or U11246 (N_11246,N_10592,N_10764);
nor U11247 (N_11247,N_10803,N_10442);
nor U11248 (N_11248,N_10526,N_10316);
and U11249 (N_11249,N_10806,N_10893);
nor U11250 (N_11250,N_10562,N_10819);
nand U11251 (N_11251,N_10612,N_10565);
and U11252 (N_11252,N_10626,N_10662);
or U11253 (N_11253,N_10989,N_10048);
nand U11254 (N_11254,N_10678,N_10233);
or U11255 (N_11255,N_10753,N_10628);
nor U11256 (N_11256,N_10167,N_10232);
nor U11257 (N_11257,N_10614,N_10075);
nand U11258 (N_11258,N_10454,N_10058);
xnor U11259 (N_11259,N_10028,N_10213);
xor U11260 (N_11260,N_10500,N_10127);
nand U11261 (N_11261,N_10836,N_10234);
nand U11262 (N_11262,N_10977,N_10041);
or U11263 (N_11263,N_10929,N_10711);
xor U11264 (N_11264,N_10009,N_10379);
nor U11265 (N_11265,N_10757,N_10619);
nor U11266 (N_11266,N_10864,N_10064);
and U11267 (N_11267,N_10432,N_10195);
and U11268 (N_11268,N_10972,N_10251);
xnor U11269 (N_11269,N_10930,N_10474);
nor U11270 (N_11270,N_10243,N_10144);
and U11271 (N_11271,N_10448,N_10863);
nand U11272 (N_11272,N_10324,N_10897);
and U11273 (N_11273,N_10305,N_10923);
or U11274 (N_11274,N_10334,N_10231);
and U11275 (N_11275,N_10869,N_10459);
or U11276 (N_11276,N_10924,N_10282);
nand U11277 (N_11277,N_10750,N_10382);
xnor U11278 (N_11278,N_10891,N_10472);
nand U11279 (N_11279,N_10853,N_10940);
and U11280 (N_11280,N_10971,N_10146);
nor U11281 (N_11281,N_10164,N_10455);
xnor U11282 (N_11282,N_10567,N_10227);
nand U11283 (N_11283,N_10591,N_10583);
xor U11284 (N_11284,N_10674,N_10457);
xnor U11285 (N_11285,N_10204,N_10560);
nor U11286 (N_11286,N_10034,N_10903);
or U11287 (N_11287,N_10725,N_10676);
nand U11288 (N_11288,N_10530,N_10616);
and U11289 (N_11289,N_10906,N_10346);
and U11290 (N_11290,N_10160,N_10867);
nand U11291 (N_11291,N_10096,N_10252);
and U11292 (N_11292,N_10588,N_10268);
nor U11293 (N_11293,N_10777,N_10168);
xor U11294 (N_11294,N_10607,N_10597);
nand U11295 (N_11295,N_10185,N_10756);
nand U11296 (N_11296,N_10409,N_10297);
xor U11297 (N_11297,N_10964,N_10969);
nor U11298 (N_11298,N_10933,N_10842);
and U11299 (N_11299,N_10319,N_10276);
and U11300 (N_11300,N_10384,N_10318);
and U11301 (N_11301,N_10012,N_10789);
xnor U11302 (N_11302,N_10262,N_10858);
xor U11303 (N_11303,N_10935,N_10199);
xnor U11304 (N_11304,N_10734,N_10704);
nor U11305 (N_11305,N_10326,N_10942);
xnor U11306 (N_11306,N_10181,N_10875);
nand U11307 (N_11307,N_10029,N_10317);
nand U11308 (N_11308,N_10030,N_10860);
nand U11309 (N_11309,N_10366,N_10102);
or U11310 (N_11310,N_10197,N_10165);
or U11311 (N_11311,N_10682,N_10767);
xnor U11312 (N_11312,N_10450,N_10918);
nand U11313 (N_11313,N_10554,N_10827);
nor U11314 (N_11314,N_10218,N_10246);
and U11315 (N_11315,N_10538,N_10484);
or U11316 (N_11316,N_10113,N_10415);
and U11317 (N_11317,N_10579,N_10240);
xor U11318 (N_11318,N_10264,N_10963);
or U11319 (N_11319,N_10485,N_10003);
nor U11320 (N_11320,N_10280,N_10001);
nor U11321 (N_11321,N_10656,N_10338);
nand U11322 (N_11322,N_10344,N_10374);
xor U11323 (N_11323,N_10016,N_10575);
xnor U11324 (N_11324,N_10649,N_10007);
nand U11325 (N_11325,N_10335,N_10487);
and U11326 (N_11326,N_10401,N_10237);
or U11327 (N_11327,N_10722,N_10499);
and U11328 (N_11328,N_10598,N_10555);
and U11329 (N_11329,N_10089,N_10625);
or U11330 (N_11330,N_10333,N_10425);
nor U11331 (N_11331,N_10620,N_10752);
nor U11332 (N_11332,N_10238,N_10159);
xnor U11333 (N_11333,N_10473,N_10646);
and U11334 (N_11334,N_10889,N_10321);
nand U11335 (N_11335,N_10780,N_10148);
xnor U11336 (N_11336,N_10730,N_10611);
xnor U11337 (N_11337,N_10263,N_10539);
and U11338 (N_11338,N_10606,N_10664);
xnor U11339 (N_11339,N_10273,N_10943);
or U11340 (N_11340,N_10059,N_10749);
xnor U11341 (N_11341,N_10600,N_10831);
nor U11342 (N_11342,N_10909,N_10993);
nor U11343 (N_11343,N_10666,N_10013);
or U11344 (N_11344,N_10697,N_10387);
or U11345 (N_11345,N_10033,N_10627);
or U11346 (N_11346,N_10203,N_10936);
and U11347 (N_11347,N_10249,N_10872);
xnor U11348 (N_11348,N_10830,N_10063);
and U11349 (N_11349,N_10210,N_10811);
xor U11350 (N_11350,N_10690,N_10609);
and U11351 (N_11351,N_10778,N_10373);
and U11352 (N_11352,N_10714,N_10833);
or U11353 (N_11353,N_10368,N_10512);
nor U11354 (N_11354,N_10898,N_10495);
and U11355 (N_11355,N_10880,N_10031);
and U11356 (N_11356,N_10313,N_10507);
and U11357 (N_11357,N_10286,N_10112);
xnor U11358 (N_11358,N_10978,N_10394);
nor U11359 (N_11359,N_10534,N_10323);
or U11360 (N_11360,N_10301,N_10642);
and U11361 (N_11361,N_10438,N_10991);
and U11362 (N_11362,N_10541,N_10186);
xnor U11363 (N_11363,N_10712,N_10398);
nor U11364 (N_11364,N_10632,N_10586);
xor U11365 (N_11365,N_10045,N_10052);
xnor U11366 (N_11366,N_10222,N_10890);
and U11367 (N_11367,N_10211,N_10219);
and U11368 (N_11368,N_10515,N_10663);
nand U11369 (N_11369,N_10797,N_10378);
nand U11370 (N_11370,N_10300,N_10825);
or U11371 (N_11371,N_10256,N_10779);
nor U11372 (N_11372,N_10443,N_10360);
or U11373 (N_11373,N_10098,N_10771);
nor U11374 (N_11374,N_10888,N_10622);
nor U11375 (N_11375,N_10271,N_10689);
nor U11376 (N_11376,N_10997,N_10805);
nand U11377 (N_11377,N_10011,N_10650);
nand U11378 (N_11378,N_10269,N_10894);
nand U11379 (N_11379,N_10361,N_10283);
nor U11380 (N_11380,N_10191,N_10655);
and U11381 (N_11381,N_10504,N_10845);
nor U11382 (N_11382,N_10099,N_10992);
nand U11383 (N_11383,N_10208,N_10996);
nand U11384 (N_11384,N_10226,N_10915);
and U11385 (N_11385,N_10293,N_10060);
xor U11386 (N_11386,N_10150,N_10347);
xor U11387 (N_11387,N_10458,N_10087);
nand U11388 (N_11388,N_10557,N_10047);
nand U11389 (N_11389,N_10032,N_10291);
or U11390 (N_11390,N_10383,N_10071);
and U11391 (N_11391,N_10118,N_10466);
xor U11392 (N_11392,N_10761,N_10781);
or U11393 (N_11393,N_10856,N_10105);
or U11394 (N_11394,N_10109,N_10475);
or U11395 (N_11395,N_10314,N_10582);
xor U11396 (N_11396,N_10193,N_10859);
or U11397 (N_11397,N_10976,N_10680);
xor U11398 (N_11398,N_10904,N_10177);
and U11399 (N_11399,N_10141,N_10139);
and U11400 (N_11400,N_10000,N_10640);
nor U11401 (N_11401,N_10123,N_10590);
and U11402 (N_11402,N_10759,N_10865);
nor U11403 (N_11403,N_10965,N_10414);
xor U11404 (N_11404,N_10949,N_10453);
nor U11405 (N_11405,N_10727,N_10172);
nor U11406 (N_11406,N_10883,N_10103);
or U11407 (N_11407,N_10290,N_10885);
xor U11408 (N_11408,N_10235,N_10312);
and U11409 (N_11409,N_10735,N_10724);
or U11410 (N_11410,N_10253,N_10325);
and U11411 (N_11411,N_10615,N_10531);
xor U11412 (N_11412,N_10043,N_10085);
nor U11413 (N_11413,N_10149,N_10162);
or U11414 (N_11414,N_10683,N_10980);
and U11415 (N_11415,N_10599,N_10241);
xnor U11416 (N_11416,N_10161,N_10679);
xnor U11417 (N_11417,N_10772,N_10786);
or U11418 (N_11418,N_10669,N_10798);
nor U11419 (N_11419,N_10430,N_10785);
nand U11420 (N_11420,N_10952,N_10550);
nand U11421 (N_11421,N_10408,N_10706);
nor U11422 (N_11422,N_10017,N_10886);
xnor U11423 (N_11423,N_10543,N_10793);
xor U11424 (N_11424,N_10130,N_10287);
xor U11425 (N_11425,N_10792,N_10788);
or U11426 (N_11426,N_10631,N_10369);
xnor U11427 (N_11427,N_10633,N_10194);
xnor U11428 (N_11428,N_10719,N_10061);
nand U11429 (N_11429,N_10228,N_10681);
and U11430 (N_11430,N_10835,N_10731);
xor U11431 (N_11431,N_10258,N_10569);
nand U11432 (N_11432,N_10703,N_10763);
nor U11433 (N_11433,N_10381,N_10351);
nor U11434 (N_11434,N_10729,N_10488);
or U11435 (N_11435,N_10966,N_10364);
or U11436 (N_11436,N_10608,N_10564);
nor U11437 (N_11437,N_10748,N_10309);
or U11438 (N_11438,N_10224,N_10822);
nand U11439 (N_11439,N_10343,N_10998);
nor U11440 (N_11440,N_10349,N_10901);
and U11441 (N_11441,N_10214,N_10644);
and U11442 (N_11442,N_10274,N_10815);
nor U11443 (N_11443,N_10694,N_10468);
and U11444 (N_11444,N_10755,N_10718);
and U11445 (N_11445,N_10122,N_10946);
xor U11446 (N_11446,N_10900,N_10322);
nor U11447 (N_11447,N_10737,N_10804);
xnor U11448 (N_11448,N_10080,N_10635);
nand U11449 (N_11449,N_10861,N_10854);
nor U11450 (N_11450,N_10173,N_10412);
or U11451 (N_11451,N_10084,N_10452);
nor U11452 (N_11452,N_10720,N_10672);
xor U11453 (N_11453,N_10916,N_10198);
nand U11454 (N_11454,N_10070,N_10984);
or U11455 (N_11455,N_10801,N_10134);
nand U11456 (N_11456,N_10675,N_10209);
and U11457 (N_11457,N_10178,N_10768);
and U11458 (N_11458,N_10026,N_10732);
nand U11459 (N_11459,N_10710,N_10826);
or U11460 (N_11460,N_10698,N_10445);
xor U11461 (N_11461,N_10479,N_10857);
xnor U11462 (N_11462,N_10561,N_10967);
nand U11463 (N_11463,N_10817,N_10695);
xnor U11464 (N_11464,N_10593,N_10913);
and U11465 (N_11465,N_10427,N_10049);
or U11466 (N_11466,N_10540,N_10517);
nand U11467 (N_11467,N_10740,N_10810);
xor U11468 (N_11468,N_10370,N_10754);
or U11469 (N_11469,N_10818,N_10170);
and U11470 (N_11470,N_10463,N_10272);
and U11471 (N_11471,N_10376,N_10046);
xnor U11472 (N_11472,N_10220,N_10536);
xor U11473 (N_11473,N_10039,N_10873);
nor U11474 (N_11474,N_10770,N_10547);
and U11475 (N_11475,N_10688,N_10447);
nor U11476 (N_11476,N_10846,N_10638);
xor U11477 (N_11477,N_10404,N_10418);
nor U11478 (N_11478,N_10685,N_10388);
nand U11479 (N_11479,N_10610,N_10330);
nand U11480 (N_11480,N_10154,N_10868);
and U11481 (N_11481,N_10306,N_10926);
and U11482 (N_11482,N_10004,N_10524);
nand U11483 (N_11483,N_10094,N_10953);
nand U11484 (N_11484,N_10138,N_10957);
or U11485 (N_11485,N_10465,N_10696);
or U11486 (N_11486,N_10020,N_10950);
xnor U11487 (N_11487,N_10019,N_10686);
or U11488 (N_11488,N_10106,N_10882);
nand U11489 (N_11489,N_10765,N_10939);
or U11490 (N_11490,N_10478,N_10871);
nand U11491 (N_11491,N_10738,N_10970);
or U11492 (N_11492,N_10907,N_10506);
xor U11493 (N_11493,N_10223,N_10800);
nor U11494 (N_11494,N_10266,N_10829);
or U11495 (N_11495,N_10618,N_10460);
nor U11496 (N_11496,N_10328,N_10486);
or U11497 (N_11497,N_10747,N_10265);
nand U11498 (N_11498,N_10760,N_10693);
xnor U11499 (N_11499,N_10914,N_10774);
or U11500 (N_11500,N_10318,N_10205);
xor U11501 (N_11501,N_10095,N_10509);
nor U11502 (N_11502,N_10007,N_10209);
nor U11503 (N_11503,N_10069,N_10903);
nand U11504 (N_11504,N_10551,N_10479);
and U11505 (N_11505,N_10214,N_10980);
nor U11506 (N_11506,N_10717,N_10898);
xnor U11507 (N_11507,N_10395,N_10655);
nand U11508 (N_11508,N_10543,N_10132);
and U11509 (N_11509,N_10064,N_10296);
xor U11510 (N_11510,N_10190,N_10795);
xor U11511 (N_11511,N_10440,N_10028);
or U11512 (N_11512,N_10024,N_10731);
and U11513 (N_11513,N_10026,N_10389);
nand U11514 (N_11514,N_10196,N_10115);
nor U11515 (N_11515,N_10837,N_10870);
and U11516 (N_11516,N_10329,N_10366);
nor U11517 (N_11517,N_10593,N_10201);
and U11518 (N_11518,N_10175,N_10572);
xnor U11519 (N_11519,N_10047,N_10604);
nand U11520 (N_11520,N_10343,N_10845);
nor U11521 (N_11521,N_10091,N_10664);
nor U11522 (N_11522,N_10535,N_10652);
or U11523 (N_11523,N_10417,N_10782);
nor U11524 (N_11524,N_10317,N_10269);
or U11525 (N_11525,N_10216,N_10418);
or U11526 (N_11526,N_10578,N_10204);
nand U11527 (N_11527,N_10620,N_10990);
nand U11528 (N_11528,N_10305,N_10349);
nand U11529 (N_11529,N_10132,N_10886);
xnor U11530 (N_11530,N_10528,N_10248);
or U11531 (N_11531,N_10223,N_10209);
and U11532 (N_11532,N_10174,N_10764);
xor U11533 (N_11533,N_10581,N_10963);
and U11534 (N_11534,N_10946,N_10452);
nand U11535 (N_11535,N_10680,N_10922);
xnor U11536 (N_11536,N_10168,N_10072);
or U11537 (N_11537,N_10410,N_10835);
nor U11538 (N_11538,N_10096,N_10210);
nand U11539 (N_11539,N_10064,N_10146);
or U11540 (N_11540,N_10099,N_10483);
or U11541 (N_11541,N_10136,N_10510);
or U11542 (N_11542,N_10673,N_10285);
or U11543 (N_11543,N_10346,N_10358);
nor U11544 (N_11544,N_10590,N_10826);
and U11545 (N_11545,N_10137,N_10878);
nand U11546 (N_11546,N_10005,N_10289);
xnor U11547 (N_11547,N_10168,N_10958);
xor U11548 (N_11548,N_10884,N_10190);
nor U11549 (N_11549,N_10371,N_10448);
and U11550 (N_11550,N_10952,N_10109);
nor U11551 (N_11551,N_10232,N_10189);
or U11552 (N_11552,N_10797,N_10900);
and U11553 (N_11553,N_10445,N_10660);
xnor U11554 (N_11554,N_10135,N_10919);
nor U11555 (N_11555,N_10048,N_10802);
xnor U11556 (N_11556,N_10189,N_10360);
nand U11557 (N_11557,N_10018,N_10347);
or U11558 (N_11558,N_10296,N_10098);
xor U11559 (N_11559,N_10347,N_10359);
nor U11560 (N_11560,N_10080,N_10921);
nand U11561 (N_11561,N_10288,N_10750);
nand U11562 (N_11562,N_10821,N_10694);
nand U11563 (N_11563,N_10942,N_10385);
or U11564 (N_11564,N_10125,N_10118);
xnor U11565 (N_11565,N_10291,N_10074);
and U11566 (N_11566,N_10669,N_10188);
and U11567 (N_11567,N_10679,N_10191);
or U11568 (N_11568,N_10445,N_10335);
nand U11569 (N_11569,N_10856,N_10921);
xnor U11570 (N_11570,N_10753,N_10356);
nand U11571 (N_11571,N_10683,N_10787);
xor U11572 (N_11572,N_10382,N_10133);
and U11573 (N_11573,N_10154,N_10912);
xnor U11574 (N_11574,N_10446,N_10423);
or U11575 (N_11575,N_10258,N_10650);
nand U11576 (N_11576,N_10582,N_10760);
or U11577 (N_11577,N_10644,N_10896);
nand U11578 (N_11578,N_10957,N_10016);
nand U11579 (N_11579,N_10845,N_10009);
nor U11580 (N_11580,N_10261,N_10557);
nand U11581 (N_11581,N_10459,N_10340);
nor U11582 (N_11582,N_10551,N_10809);
or U11583 (N_11583,N_10890,N_10030);
and U11584 (N_11584,N_10782,N_10618);
and U11585 (N_11585,N_10860,N_10200);
xnor U11586 (N_11586,N_10815,N_10504);
or U11587 (N_11587,N_10531,N_10395);
or U11588 (N_11588,N_10786,N_10343);
nand U11589 (N_11589,N_10720,N_10804);
or U11590 (N_11590,N_10061,N_10257);
and U11591 (N_11591,N_10676,N_10573);
and U11592 (N_11592,N_10071,N_10481);
xor U11593 (N_11593,N_10450,N_10317);
and U11594 (N_11594,N_10040,N_10991);
xnor U11595 (N_11595,N_10467,N_10793);
or U11596 (N_11596,N_10319,N_10476);
and U11597 (N_11597,N_10262,N_10943);
xor U11598 (N_11598,N_10144,N_10535);
or U11599 (N_11599,N_10472,N_10158);
nand U11600 (N_11600,N_10953,N_10661);
xor U11601 (N_11601,N_10654,N_10071);
nand U11602 (N_11602,N_10480,N_10921);
xor U11603 (N_11603,N_10119,N_10388);
nand U11604 (N_11604,N_10347,N_10780);
and U11605 (N_11605,N_10795,N_10665);
nand U11606 (N_11606,N_10200,N_10015);
nand U11607 (N_11607,N_10145,N_10116);
nand U11608 (N_11608,N_10657,N_10448);
and U11609 (N_11609,N_10675,N_10657);
nand U11610 (N_11610,N_10757,N_10024);
xor U11611 (N_11611,N_10180,N_10232);
or U11612 (N_11612,N_10122,N_10243);
xnor U11613 (N_11613,N_10985,N_10168);
xnor U11614 (N_11614,N_10039,N_10728);
nor U11615 (N_11615,N_10663,N_10032);
nand U11616 (N_11616,N_10895,N_10735);
nand U11617 (N_11617,N_10706,N_10135);
nand U11618 (N_11618,N_10072,N_10298);
and U11619 (N_11619,N_10967,N_10187);
nor U11620 (N_11620,N_10291,N_10175);
nor U11621 (N_11621,N_10930,N_10124);
and U11622 (N_11622,N_10575,N_10208);
or U11623 (N_11623,N_10915,N_10037);
and U11624 (N_11624,N_10015,N_10083);
or U11625 (N_11625,N_10237,N_10193);
xnor U11626 (N_11626,N_10783,N_10444);
nand U11627 (N_11627,N_10297,N_10060);
or U11628 (N_11628,N_10266,N_10989);
or U11629 (N_11629,N_10114,N_10889);
xor U11630 (N_11630,N_10924,N_10681);
and U11631 (N_11631,N_10738,N_10205);
and U11632 (N_11632,N_10474,N_10335);
nor U11633 (N_11633,N_10758,N_10010);
xnor U11634 (N_11634,N_10244,N_10087);
xor U11635 (N_11635,N_10268,N_10418);
xor U11636 (N_11636,N_10017,N_10535);
xnor U11637 (N_11637,N_10765,N_10707);
and U11638 (N_11638,N_10828,N_10069);
or U11639 (N_11639,N_10473,N_10819);
xnor U11640 (N_11640,N_10735,N_10486);
nand U11641 (N_11641,N_10436,N_10940);
xnor U11642 (N_11642,N_10122,N_10344);
and U11643 (N_11643,N_10081,N_10896);
nor U11644 (N_11644,N_10715,N_10796);
xor U11645 (N_11645,N_10072,N_10568);
or U11646 (N_11646,N_10591,N_10405);
nor U11647 (N_11647,N_10892,N_10651);
xnor U11648 (N_11648,N_10447,N_10702);
nor U11649 (N_11649,N_10147,N_10036);
xor U11650 (N_11650,N_10336,N_10346);
nand U11651 (N_11651,N_10172,N_10754);
nand U11652 (N_11652,N_10294,N_10068);
and U11653 (N_11653,N_10804,N_10109);
nor U11654 (N_11654,N_10263,N_10137);
xor U11655 (N_11655,N_10923,N_10847);
or U11656 (N_11656,N_10546,N_10662);
nor U11657 (N_11657,N_10160,N_10666);
and U11658 (N_11658,N_10544,N_10560);
xor U11659 (N_11659,N_10272,N_10367);
xnor U11660 (N_11660,N_10662,N_10760);
xnor U11661 (N_11661,N_10905,N_10305);
nor U11662 (N_11662,N_10650,N_10668);
xnor U11663 (N_11663,N_10331,N_10093);
xor U11664 (N_11664,N_10262,N_10754);
and U11665 (N_11665,N_10417,N_10546);
or U11666 (N_11666,N_10936,N_10628);
or U11667 (N_11667,N_10572,N_10292);
or U11668 (N_11668,N_10487,N_10897);
and U11669 (N_11669,N_10591,N_10861);
nor U11670 (N_11670,N_10705,N_10690);
nand U11671 (N_11671,N_10808,N_10494);
nor U11672 (N_11672,N_10342,N_10066);
and U11673 (N_11673,N_10717,N_10759);
or U11674 (N_11674,N_10716,N_10498);
xor U11675 (N_11675,N_10644,N_10949);
xor U11676 (N_11676,N_10538,N_10292);
nor U11677 (N_11677,N_10278,N_10642);
and U11678 (N_11678,N_10861,N_10487);
and U11679 (N_11679,N_10526,N_10839);
nor U11680 (N_11680,N_10262,N_10671);
nand U11681 (N_11681,N_10573,N_10519);
xnor U11682 (N_11682,N_10079,N_10243);
and U11683 (N_11683,N_10401,N_10990);
or U11684 (N_11684,N_10032,N_10156);
nor U11685 (N_11685,N_10902,N_10593);
nor U11686 (N_11686,N_10394,N_10172);
nand U11687 (N_11687,N_10653,N_10102);
nand U11688 (N_11688,N_10052,N_10577);
nand U11689 (N_11689,N_10377,N_10961);
nor U11690 (N_11690,N_10406,N_10499);
xnor U11691 (N_11691,N_10069,N_10876);
nor U11692 (N_11692,N_10062,N_10999);
nand U11693 (N_11693,N_10904,N_10530);
xor U11694 (N_11694,N_10121,N_10201);
nor U11695 (N_11695,N_10614,N_10642);
nand U11696 (N_11696,N_10500,N_10722);
or U11697 (N_11697,N_10083,N_10659);
nand U11698 (N_11698,N_10563,N_10605);
or U11699 (N_11699,N_10514,N_10498);
nor U11700 (N_11700,N_10356,N_10406);
nor U11701 (N_11701,N_10881,N_10701);
xor U11702 (N_11702,N_10710,N_10659);
and U11703 (N_11703,N_10449,N_10924);
or U11704 (N_11704,N_10104,N_10413);
xnor U11705 (N_11705,N_10932,N_10696);
xnor U11706 (N_11706,N_10418,N_10934);
or U11707 (N_11707,N_10105,N_10585);
xnor U11708 (N_11708,N_10132,N_10222);
or U11709 (N_11709,N_10134,N_10451);
and U11710 (N_11710,N_10730,N_10971);
nor U11711 (N_11711,N_10534,N_10186);
or U11712 (N_11712,N_10904,N_10684);
nand U11713 (N_11713,N_10970,N_10353);
or U11714 (N_11714,N_10435,N_10479);
and U11715 (N_11715,N_10045,N_10626);
nand U11716 (N_11716,N_10964,N_10671);
nand U11717 (N_11717,N_10706,N_10950);
nor U11718 (N_11718,N_10308,N_10350);
nand U11719 (N_11719,N_10767,N_10176);
and U11720 (N_11720,N_10901,N_10734);
nor U11721 (N_11721,N_10477,N_10194);
nor U11722 (N_11722,N_10559,N_10683);
and U11723 (N_11723,N_10549,N_10737);
nor U11724 (N_11724,N_10111,N_10001);
xnor U11725 (N_11725,N_10033,N_10385);
nor U11726 (N_11726,N_10415,N_10624);
nand U11727 (N_11727,N_10431,N_10349);
xnor U11728 (N_11728,N_10552,N_10568);
xor U11729 (N_11729,N_10715,N_10126);
or U11730 (N_11730,N_10698,N_10611);
and U11731 (N_11731,N_10791,N_10031);
and U11732 (N_11732,N_10743,N_10356);
nand U11733 (N_11733,N_10940,N_10938);
or U11734 (N_11734,N_10950,N_10454);
xor U11735 (N_11735,N_10864,N_10558);
xor U11736 (N_11736,N_10107,N_10752);
and U11737 (N_11737,N_10863,N_10733);
xor U11738 (N_11738,N_10965,N_10877);
xnor U11739 (N_11739,N_10020,N_10797);
and U11740 (N_11740,N_10467,N_10368);
and U11741 (N_11741,N_10013,N_10031);
xnor U11742 (N_11742,N_10672,N_10285);
xnor U11743 (N_11743,N_10303,N_10942);
or U11744 (N_11744,N_10294,N_10439);
xor U11745 (N_11745,N_10132,N_10152);
and U11746 (N_11746,N_10152,N_10506);
or U11747 (N_11747,N_10680,N_10517);
xnor U11748 (N_11748,N_10818,N_10350);
nand U11749 (N_11749,N_10402,N_10144);
or U11750 (N_11750,N_10966,N_10895);
nand U11751 (N_11751,N_10549,N_10589);
xnor U11752 (N_11752,N_10286,N_10743);
and U11753 (N_11753,N_10093,N_10003);
nand U11754 (N_11754,N_10795,N_10725);
nand U11755 (N_11755,N_10957,N_10584);
nand U11756 (N_11756,N_10027,N_10569);
and U11757 (N_11757,N_10704,N_10164);
and U11758 (N_11758,N_10513,N_10883);
nor U11759 (N_11759,N_10928,N_10338);
nand U11760 (N_11760,N_10432,N_10318);
nor U11761 (N_11761,N_10409,N_10423);
nor U11762 (N_11762,N_10841,N_10878);
xnor U11763 (N_11763,N_10948,N_10190);
nand U11764 (N_11764,N_10704,N_10956);
nand U11765 (N_11765,N_10039,N_10494);
and U11766 (N_11766,N_10445,N_10316);
xor U11767 (N_11767,N_10732,N_10050);
nand U11768 (N_11768,N_10885,N_10806);
nor U11769 (N_11769,N_10742,N_10427);
and U11770 (N_11770,N_10780,N_10544);
nand U11771 (N_11771,N_10747,N_10684);
xor U11772 (N_11772,N_10123,N_10534);
or U11773 (N_11773,N_10786,N_10980);
and U11774 (N_11774,N_10408,N_10517);
and U11775 (N_11775,N_10061,N_10284);
and U11776 (N_11776,N_10473,N_10239);
and U11777 (N_11777,N_10736,N_10148);
xor U11778 (N_11778,N_10629,N_10983);
and U11779 (N_11779,N_10201,N_10071);
nor U11780 (N_11780,N_10595,N_10493);
and U11781 (N_11781,N_10234,N_10230);
nand U11782 (N_11782,N_10894,N_10501);
nand U11783 (N_11783,N_10838,N_10189);
nor U11784 (N_11784,N_10697,N_10271);
and U11785 (N_11785,N_10187,N_10946);
nand U11786 (N_11786,N_10057,N_10314);
nor U11787 (N_11787,N_10021,N_10896);
and U11788 (N_11788,N_10947,N_10959);
and U11789 (N_11789,N_10560,N_10871);
xnor U11790 (N_11790,N_10532,N_10900);
nand U11791 (N_11791,N_10857,N_10191);
or U11792 (N_11792,N_10567,N_10864);
nand U11793 (N_11793,N_10805,N_10415);
and U11794 (N_11794,N_10395,N_10770);
nand U11795 (N_11795,N_10662,N_10819);
xnor U11796 (N_11796,N_10925,N_10662);
xor U11797 (N_11797,N_10031,N_10112);
nand U11798 (N_11798,N_10661,N_10428);
and U11799 (N_11799,N_10469,N_10816);
nor U11800 (N_11800,N_10625,N_10759);
or U11801 (N_11801,N_10152,N_10140);
nor U11802 (N_11802,N_10559,N_10653);
and U11803 (N_11803,N_10880,N_10646);
or U11804 (N_11804,N_10050,N_10363);
nand U11805 (N_11805,N_10151,N_10513);
and U11806 (N_11806,N_10994,N_10294);
nand U11807 (N_11807,N_10324,N_10097);
and U11808 (N_11808,N_10447,N_10381);
xnor U11809 (N_11809,N_10621,N_10419);
nand U11810 (N_11810,N_10321,N_10639);
nor U11811 (N_11811,N_10531,N_10629);
or U11812 (N_11812,N_10345,N_10835);
and U11813 (N_11813,N_10922,N_10571);
and U11814 (N_11814,N_10981,N_10761);
or U11815 (N_11815,N_10224,N_10469);
nor U11816 (N_11816,N_10545,N_10985);
nor U11817 (N_11817,N_10802,N_10747);
xor U11818 (N_11818,N_10507,N_10864);
nor U11819 (N_11819,N_10069,N_10541);
or U11820 (N_11820,N_10035,N_10767);
nor U11821 (N_11821,N_10857,N_10476);
or U11822 (N_11822,N_10114,N_10405);
nor U11823 (N_11823,N_10016,N_10121);
and U11824 (N_11824,N_10314,N_10157);
xnor U11825 (N_11825,N_10353,N_10487);
or U11826 (N_11826,N_10400,N_10777);
or U11827 (N_11827,N_10387,N_10097);
nand U11828 (N_11828,N_10554,N_10777);
or U11829 (N_11829,N_10473,N_10501);
xor U11830 (N_11830,N_10049,N_10643);
or U11831 (N_11831,N_10767,N_10362);
and U11832 (N_11832,N_10263,N_10892);
nor U11833 (N_11833,N_10257,N_10899);
or U11834 (N_11834,N_10517,N_10343);
nor U11835 (N_11835,N_10402,N_10419);
or U11836 (N_11836,N_10350,N_10098);
nand U11837 (N_11837,N_10879,N_10658);
xnor U11838 (N_11838,N_10476,N_10138);
or U11839 (N_11839,N_10496,N_10075);
nand U11840 (N_11840,N_10095,N_10424);
nand U11841 (N_11841,N_10148,N_10224);
and U11842 (N_11842,N_10523,N_10927);
nor U11843 (N_11843,N_10288,N_10643);
and U11844 (N_11844,N_10997,N_10301);
xnor U11845 (N_11845,N_10741,N_10996);
or U11846 (N_11846,N_10711,N_10824);
and U11847 (N_11847,N_10896,N_10314);
or U11848 (N_11848,N_10073,N_10045);
nor U11849 (N_11849,N_10403,N_10095);
xor U11850 (N_11850,N_10277,N_10585);
nand U11851 (N_11851,N_10320,N_10444);
nand U11852 (N_11852,N_10901,N_10051);
xnor U11853 (N_11853,N_10933,N_10521);
nand U11854 (N_11854,N_10861,N_10936);
nand U11855 (N_11855,N_10507,N_10756);
nand U11856 (N_11856,N_10649,N_10272);
xnor U11857 (N_11857,N_10214,N_10354);
nand U11858 (N_11858,N_10266,N_10876);
and U11859 (N_11859,N_10176,N_10457);
or U11860 (N_11860,N_10884,N_10410);
and U11861 (N_11861,N_10571,N_10595);
nand U11862 (N_11862,N_10278,N_10204);
nor U11863 (N_11863,N_10808,N_10285);
or U11864 (N_11864,N_10434,N_10262);
nand U11865 (N_11865,N_10598,N_10825);
and U11866 (N_11866,N_10878,N_10449);
nor U11867 (N_11867,N_10460,N_10554);
nor U11868 (N_11868,N_10574,N_10636);
nor U11869 (N_11869,N_10026,N_10834);
or U11870 (N_11870,N_10843,N_10027);
or U11871 (N_11871,N_10706,N_10758);
or U11872 (N_11872,N_10662,N_10160);
or U11873 (N_11873,N_10798,N_10915);
or U11874 (N_11874,N_10695,N_10744);
xnor U11875 (N_11875,N_10694,N_10572);
and U11876 (N_11876,N_10738,N_10507);
nor U11877 (N_11877,N_10884,N_10560);
nor U11878 (N_11878,N_10450,N_10734);
xor U11879 (N_11879,N_10674,N_10294);
and U11880 (N_11880,N_10305,N_10427);
nor U11881 (N_11881,N_10280,N_10365);
nor U11882 (N_11882,N_10520,N_10635);
xor U11883 (N_11883,N_10950,N_10184);
nand U11884 (N_11884,N_10821,N_10621);
nand U11885 (N_11885,N_10287,N_10026);
and U11886 (N_11886,N_10954,N_10671);
nand U11887 (N_11887,N_10604,N_10937);
nor U11888 (N_11888,N_10370,N_10059);
and U11889 (N_11889,N_10671,N_10512);
xnor U11890 (N_11890,N_10954,N_10818);
and U11891 (N_11891,N_10457,N_10596);
nor U11892 (N_11892,N_10115,N_10090);
xnor U11893 (N_11893,N_10599,N_10053);
or U11894 (N_11894,N_10859,N_10982);
and U11895 (N_11895,N_10788,N_10968);
nand U11896 (N_11896,N_10698,N_10716);
or U11897 (N_11897,N_10479,N_10374);
or U11898 (N_11898,N_10939,N_10096);
or U11899 (N_11899,N_10935,N_10063);
nor U11900 (N_11900,N_10227,N_10273);
and U11901 (N_11901,N_10244,N_10296);
nor U11902 (N_11902,N_10732,N_10589);
nand U11903 (N_11903,N_10970,N_10316);
nand U11904 (N_11904,N_10151,N_10487);
nand U11905 (N_11905,N_10493,N_10079);
nor U11906 (N_11906,N_10805,N_10911);
or U11907 (N_11907,N_10417,N_10930);
xor U11908 (N_11908,N_10469,N_10723);
and U11909 (N_11909,N_10161,N_10430);
or U11910 (N_11910,N_10314,N_10530);
and U11911 (N_11911,N_10161,N_10702);
nand U11912 (N_11912,N_10605,N_10254);
and U11913 (N_11913,N_10337,N_10095);
xor U11914 (N_11914,N_10638,N_10598);
or U11915 (N_11915,N_10488,N_10968);
nor U11916 (N_11916,N_10126,N_10289);
nor U11917 (N_11917,N_10933,N_10079);
and U11918 (N_11918,N_10560,N_10133);
or U11919 (N_11919,N_10201,N_10161);
or U11920 (N_11920,N_10073,N_10357);
nand U11921 (N_11921,N_10269,N_10530);
xor U11922 (N_11922,N_10086,N_10150);
nand U11923 (N_11923,N_10943,N_10090);
nand U11924 (N_11924,N_10455,N_10959);
nand U11925 (N_11925,N_10865,N_10833);
nand U11926 (N_11926,N_10315,N_10668);
nand U11927 (N_11927,N_10210,N_10365);
or U11928 (N_11928,N_10005,N_10578);
xnor U11929 (N_11929,N_10391,N_10155);
and U11930 (N_11930,N_10988,N_10153);
or U11931 (N_11931,N_10501,N_10442);
and U11932 (N_11932,N_10334,N_10331);
and U11933 (N_11933,N_10996,N_10058);
nor U11934 (N_11934,N_10941,N_10877);
nor U11935 (N_11935,N_10065,N_10622);
nand U11936 (N_11936,N_10871,N_10503);
nand U11937 (N_11937,N_10984,N_10078);
or U11938 (N_11938,N_10140,N_10955);
nand U11939 (N_11939,N_10661,N_10506);
or U11940 (N_11940,N_10853,N_10923);
or U11941 (N_11941,N_10975,N_10181);
nor U11942 (N_11942,N_10290,N_10773);
or U11943 (N_11943,N_10073,N_10621);
and U11944 (N_11944,N_10167,N_10225);
nor U11945 (N_11945,N_10765,N_10215);
xor U11946 (N_11946,N_10666,N_10738);
nor U11947 (N_11947,N_10978,N_10860);
and U11948 (N_11948,N_10284,N_10252);
xnor U11949 (N_11949,N_10751,N_10707);
nand U11950 (N_11950,N_10825,N_10301);
xor U11951 (N_11951,N_10078,N_10732);
nand U11952 (N_11952,N_10630,N_10171);
and U11953 (N_11953,N_10492,N_10240);
or U11954 (N_11954,N_10993,N_10785);
nor U11955 (N_11955,N_10692,N_10725);
or U11956 (N_11956,N_10379,N_10776);
nand U11957 (N_11957,N_10673,N_10341);
nor U11958 (N_11958,N_10041,N_10850);
nor U11959 (N_11959,N_10925,N_10950);
nor U11960 (N_11960,N_10396,N_10468);
nor U11961 (N_11961,N_10738,N_10382);
nand U11962 (N_11962,N_10789,N_10435);
and U11963 (N_11963,N_10449,N_10015);
and U11964 (N_11964,N_10012,N_10499);
nor U11965 (N_11965,N_10938,N_10574);
nand U11966 (N_11966,N_10257,N_10586);
xor U11967 (N_11967,N_10000,N_10402);
and U11968 (N_11968,N_10107,N_10572);
or U11969 (N_11969,N_10723,N_10219);
nand U11970 (N_11970,N_10530,N_10578);
or U11971 (N_11971,N_10624,N_10700);
xnor U11972 (N_11972,N_10163,N_10017);
or U11973 (N_11973,N_10821,N_10556);
nor U11974 (N_11974,N_10627,N_10957);
and U11975 (N_11975,N_10895,N_10605);
nor U11976 (N_11976,N_10868,N_10574);
and U11977 (N_11977,N_10570,N_10800);
nor U11978 (N_11978,N_10405,N_10955);
and U11979 (N_11979,N_10266,N_10726);
nor U11980 (N_11980,N_10430,N_10002);
nand U11981 (N_11981,N_10847,N_10580);
and U11982 (N_11982,N_10898,N_10054);
or U11983 (N_11983,N_10810,N_10197);
nand U11984 (N_11984,N_10380,N_10544);
nand U11985 (N_11985,N_10081,N_10031);
xor U11986 (N_11986,N_10383,N_10245);
nor U11987 (N_11987,N_10893,N_10186);
nand U11988 (N_11988,N_10693,N_10888);
or U11989 (N_11989,N_10352,N_10715);
xor U11990 (N_11990,N_10073,N_10099);
nor U11991 (N_11991,N_10038,N_10376);
xnor U11992 (N_11992,N_10977,N_10146);
and U11993 (N_11993,N_10494,N_10890);
nand U11994 (N_11994,N_10149,N_10207);
nand U11995 (N_11995,N_10379,N_10445);
xor U11996 (N_11996,N_10487,N_10906);
xor U11997 (N_11997,N_10574,N_10296);
xor U11998 (N_11998,N_10685,N_10789);
xnor U11999 (N_11999,N_10085,N_10228);
xor U12000 (N_12000,N_11983,N_11227);
and U12001 (N_12001,N_11899,N_11421);
or U12002 (N_12002,N_11278,N_11438);
xnor U12003 (N_12003,N_11788,N_11253);
and U12004 (N_12004,N_11272,N_11191);
or U12005 (N_12005,N_11600,N_11172);
and U12006 (N_12006,N_11688,N_11626);
or U12007 (N_12007,N_11539,N_11893);
nor U12008 (N_12008,N_11345,N_11282);
xor U12009 (N_12009,N_11632,N_11023);
or U12010 (N_12010,N_11114,N_11873);
and U12011 (N_12011,N_11661,N_11766);
nor U12012 (N_12012,N_11397,N_11540);
and U12013 (N_12013,N_11787,N_11178);
nor U12014 (N_12014,N_11925,N_11263);
nand U12015 (N_12015,N_11024,N_11008);
or U12016 (N_12016,N_11570,N_11556);
nand U12017 (N_12017,N_11380,N_11691);
or U12018 (N_12018,N_11156,N_11753);
nor U12019 (N_12019,N_11927,N_11659);
or U12020 (N_12020,N_11013,N_11603);
and U12021 (N_12021,N_11684,N_11660);
nand U12022 (N_12022,N_11897,N_11929);
and U12023 (N_12023,N_11151,N_11810);
xor U12024 (N_12024,N_11005,N_11273);
or U12025 (N_12025,N_11838,N_11746);
or U12026 (N_12026,N_11905,N_11237);
and U12027 (N_12027,N_11721,N_11548);
nor U12028 (N_12028,N_11938,N_11407);
or U12029 (N_12029,N_11484,N_11128);
nor U12030 (N_12030,N_11664,N_11568);
and U12031 (N_12031,N_11348,N_11624);
and U12032 (N_12032,N_11933,N_11775);
nand U12033 (N_12033,N_11879,N_11696);
nor U12034 (N_12034,N_11141,N_11763);
xor U12035 (N_12035,N_11785,N_11847);
nor U12036 (N_12036,N_11454,N_11119);
nor U12037 (N_12037,N_11990,N_11619);
nand U12038 (N_12038,N_11152,N_11098);
or U12039 (N_12039,N_11492,N_11646);
and U12040 (N_12040,N_11823,N_11994);
xnor U12041 (N_12041,N_11707,N_11728);
xor U12042 (N_12042,N_11804,N_11663);
and U12043 (N_12043,N_11201,N_11911);
or U12044 (N_12044,N_11895,N_11379);
nor U12045 (N_12045,N_11774,N_11786);
nand U12046 (N_12046,N_11778,N_11225);
and U12047 (N_12047,N_11700,N_11986);
xor U12048 (N_12048,N_11850,N_11486);
xor U12049 (N_12049,N_11280,N_11003);
xor U12050 (N_12050,N_11022,N_11683);
nand U12051 (N_12051,N_11388,N_11383);
nand U12052 (N_12052,N_11363,N_11713);
or U12053 (N_12053,N_11184,N_11095);
or U12054 (N_12054,N_11790,N_11306);
and U12055 (N_12055,N_11507,N_11063);
or U12056 (N_12056,N_11127,N_11487);
xor U12057 (N_12057,N_11226,N_11161);
nor U12058 (N_12058,N_11288,N_11192);
nand U12059 (N_12059,N_11997,N_11066);
xor U12060 (N_12060,N_11033,N_11678);
or U12061 (N_12061,N_11049,N_11906);
xnor U12062 (N_12062,N_11185,N_11987);
or U12063 (N_12063,N_11016,N_11674);
or U12064 (N_12064,N_11177,N_11420);
xnor U12065 (N_12065,N_11874,N_11973);
xnor U12066 (N_12066,N_11373,N_11039);
xnor U12067 (N_12067,N_11809,N_11448);
and U12068 (N_12068,N_11031,N_11305);
xnor U12069 (N_12069,N_11569,N_11665);
xnor U12070 (N_12070,N_11070,N_11290);
and U12071 (N_12071,N_11807,N_11189);
and U12072 (N_12072,N_11144,N_11286);
nor U12073 (N_12073,N_11625,N_11992);
xor U12074 (N_12074,N_11356,N_11479);
nand U12075 (N_12075,N_11068,N_11389);
xor U12076 (N_12076,N_11783,N_11137);
xor U12077 (N_12077,N_11795,N_11101);
and U12078 (N_12078,N_11208,N_11621);
or U12079 (N_12079,N_11418,N_11541);
or U12080 (N_12080,N_11223,N_11915);
nor U12081 (N_12081,N_11167,N_11868);
or U12082 (N_12082,N_11681,N_11945);
or U12083 (N_12083,N_11977,N_11452);
or U12084 (N_12084,N_11042,N_11350);
nand U12085 (N_12085,N_11944,N_11731);
and U12086 (N_12086,N_11995,N_11200);
and U12087 (N_12087,N_11030,N_11711);
nand U12088 (N_12088,N_11960,N_11687);
and U12089 (N_12089,N_11595,N_11508);
or U12090 (N_12090,N_11830,N_11322);
or U12091 (N_12091,N_11573,N_11670);
nor U12092 (N_12092,N_11108,N_11160);
xnor U12093 (N_12093,N_11179,N_11917);
and U12094 (N_12094,N_11930,N_11878);
nand U12095 (N_12095,N_11481,N_11920);
or U12096 (N_12096,N_11836,N_11107);
and U12097 (N_12097,N_11343,N_11991);
xor U12098 (N_12098,N_11970,N_11921);
nand U12099 (N_12099,N_11756,N_11637);
and U12100 (N_12100,N_11174,N_11248);
or U12101 (N_12101,N_11551,N_11542);
or U12102 (N_12102,N_11516,N_11327);
nor U12103 (N_12103,N_11502,N_11751);
xnor U12104 (N_12104,N_11186,N_11135);
xnor U12105 (N_12105,N_11017,N_11924);
nor U12106 (N_12106,N_11315,N_11162);
and U12107 (N_12107,N_11442,N_11771);
xnor U12108 (N_12108,N_11907,N_11729);
nor U12109 (N_12109,N_11577,N_11985);
nor U12110 (N_12110,N_11296,N_11193);
or U12111 (N_12111,N_11792,N_11240);
nor U12112 (N_12112,N_11163,N_11028);
and U12113 (N_12113,N_11955,N_11217);
nor U12114 (N_12114,N_11768,N_11045);
nand U12115 (N_12115,N_11565,N_11264);
and U12116 (N_12116,N_11463,N_11277);
nor U12117 (N_12117,N_11514,N_11462);
nor U12118 (N_12118,N_11811,N_11048);
nor U12119 (N_12119,N_11888,N_11863);
xnor U12120 (N_12120,N_11205,N_11939);
nand U12121 (N_12121,N_11824,N_11255);
or U12122 (N_12122,N_11839,N_11735);
xnor U12123 (N_12123,N_11585,N_11697);
xor U12124 (N_12124,N_11342,N_11401);
and U12125 (N_12125,N_11204,N_11057);
or U12126 (N_12126,N_11202,N_11212);
xnor U12127 (N_12127,N_11953,N_11717);
nor U12128 (N_12128,N_11961,N_11040);
or U12129 (N_12129,N_11090,N_11274);
and U12130 (N_12130,N_11267,N_11439);
or U12131 (N_12131,N_11676,N_11337);
or U12132 (N_12132,N_11789,N_11597);
or U12133 (N_12133,N_11269,N_11870);
nor U12134 (N_12134,N_11362,N_11550);
nand U12135 (N_12135,N_11375,N_11392);
or U12136 (N_12136,N_11082,N_11904);
or U12137 (N_12137,N_11294,N_11529);
xor U12138 (N_12138,N_11936,N_11424);
nand U12139 (N_12139,N_11950,N_11050);
nand U12140 (N_12140,N_11468,N_11846);
or U12141 (N_12141,N_11689,N_11330);
and U12142 (N_12142,N_11943,N_11558);
nor U12143 (N_12143,N_11443,N_11601);
nor U12144 (N_12144,N_11406,N_11138);
nand U12145 (N_12145,N_11109,N_11694);
nand U12146 (N_12146,N_11469,N_11909);
nor U12147 (N_12147,N_11417,N_11706);
and U12148 (N_12148,N_11121,N_11669);
nor U12149 (N_12149,N_11476,N_11015);
nor U12150 (N_12150,N_11387,N_11367);
or U12151 (N_12151,N_11826,N_11957);
nor U12152 (N_12152,N_11085,N_11859);
nor U12153 (N_12153,N_11896,N_11764);
nand U12154 (N_12154,N_11318,N_11923);
and U12155 (N_12155,N_11230,N_11941);
or U12156 (N_12156,N_11865,N_11521);
nor U12157 (N_12157,N_11313,N_11236);
xnor U12158 (N_12158,N_11988,N_11289);
xnor U12159 (N_12159,N_11371,N_11962);
or U12160 (N_12160,N_11303,N_11881);
and U12161 (N_12161,N_11599,N_11769);
nand U12162 (N_12162,N_11738,N_11582);
and U12163 (N_12163,N_11522,N_11010);
or U12164 (N_12164,N_11758,N_11472);
nor U12165 (N_12165,N_11773,N_11210);
xor U12166 (N_12166,N_11644,N_11298);
nand U12167 (N_12167,N_11937,N_11954);
nor U12168 (N_12168,N_11596,N_11384);
and U12169 (N_12169,N_11382,N_11858);
and U12170 (N_12170,N_11515,N_11394);
nor U12171 (N_12171,N_11027,N_11351);
nor U12172 (N_12172,N_11216,N_11855);
and U12173 (N_12173,N_11335,N_11475);
or U12174 (N_12174,N_11887,N_11444);
nand U12175 (N_12175,N_11750,N_11094);
and U12176 (N_12176,N_11951,N_11077);
nor U12177 (N_12177,N_11195,N_11630);
or U12178 (N_12178,N_11180,N_11146);
nor U12179 (N_12179,N_11054,N_11817);
xor U12180 (N_12180,N_11198,N_11065);
nand U12181 (N_12181,N_11919,N_11975);
nor U12182 (N_12182,N_11482,N_11651);
nand U12183 (N_12183,N_11203,N_11433);
nor U12184 (N_12184,N_11104,N_11701);
nand U12185 (N_12185,N_11222,N_11812);
nor U12186 (N_12186,N_11880,N_11680);
nand U12187 (N_12187,N_11321,N_11149);
nand U12188 (N_12188,N_11579,N_11485);
and U12189 (N_12189,N_11359,N_11658);
nand U12190 (N_12190,N_11319,N_11587);
and U12191 (N_12191,N_11060,N_11325);
xor U12192 (N_12192,N_11805,N_11358);
and U12193 (N_12193,N_11125,N_11918);
xnor U12194 (N_12194,N_11851,N_11559);
and U12195 (N_12195,N_11368,N_11650);
nand U12196 (N_12196,N_11978,N_11806);
xor U12197 (N_12197,N_11376,N_11281);
and U12198 (N_12198,N_11519,N_11317);
and U12199 (N_12199,N_11329,N_11111);
and U12200 (N_12200,N_11808,N_11260);
and U12201 (N_12201,N_11259,N_11534);
xor U12202 (N_12202,N_11244,N_11395);
xnor U12203 (N_12203,N_11093,N_11366);
xnor U12204 (N_12204,N_11971,N_11547);
xor U12205 (N_12205,N_11693,N_11640);
or U12206 (N_12206,N_11733,N_11869);
nand U12207 (N_12207,N_11390,N_11429);
or U12208 (N_12208,N_11434,N_11455);
nor U12209 (N_12209,N_11739,N_11533);
and U12210 (N_12210,N_11276,N_11526);
xnor U12211 (N_12211,N_11578,N_11912);
and U12212 (N_12212,N_11610,N_11075);
and U12213 (N_12213,N_11431,N_11834);
or U12214 (N_12214,N_11506,N_11500);
nor U12215 (N_12215,N_11842,N_11890);
nor U12216 (N_12216,N_11258,N_11667);
or U12217 (N_12217,N_11947,N_11316);
xor U12218 (N_12218,N_11825,N_11583);
nor U12219 (N_12219,N_11798,N_11471);
or U12220 (N_12220,N_11155,N_11633);
and U12221 (N_12221,N_11145,N_11349);
or U12222 (N_12222,N_11257,N_11352);
xnor U12223 (N_12223,N_11483,N_11554);
nor U12224 (N_12224,N_11903,N_11304);
nand U12225 (N_12225,N_11078,N_11404);
nor U12226 (N_12226,N_11532,N_11702);
and U12227 (N_12227,N_11207,N_11607);
nor U12228 (N_12228,N_11159,N_11037);
and U12229 (N_12229,N_11171,N_11323);
nor U12230 (N_12230,N_11501,N_11211);
or U12231 (N_12231,N_11672,N_11628);
nor U12232 (N_12232,N_11797,N_11365);
xor U12233 (N_12233,N_11690,N_11456);
xor U12234 (N_12234,N_11656,N_11385);
xnor U12235 (N_12235,N_11103,N_11035);
and U12236 (N_12236,N_11196,N_11801);
nand U12237 (N_12237,N_11877,N_11531);
xnor U12238 (N_12238,N_11041,N_11124);
or U12239 (N_12239,N_11402,N_11061);
nand U12240 (N_12240,N_11391,N_11677);
nand U12241 (N_12241,N_11636,N_11723);
nand U12242 (N_12242,N_11139,N_11649);
and U12243 (N_12243,N_11843,N_11291);
nor U12244 (N_12244,N_11736,N_11549);
xor U12245 (N_12245,N_11770,N_11357);
or U12246 (N_12246,N_11283,N_11892);
or U12247 (N_12247,N_11168,N_11898);
or U12248 (N_12248,N_11187,N_11491);
or U12249 (N_12249,N_11642,N_11705);
xor U12250 (N_12250,N_11123,N_11627);
nand U12251 (N_12251,N_11422,N_11076);
nand U12252 (N_12252,N_11328,N_11435);
xor U12253 (N_12253,N_11604,N_11331);
nand U12254 (N_12254,N_11524,N_11361);
xnor U12255 (N_12255,N_11510,N_11726);
xnor U12256 (N_12256,N_11724,N_11436);
nor U12257 (N_12257,N_11232,N_11047);
and U12258 (N_12258,N_11284,N_11464);
xnor U12259 (N_12259,N_11638,N_11183);
xnor U12260 (N_12260,N_11791,N_11635);
and U12261 (N_12261,N_11419,N_11679);
xnor U12262 (N_12262,N_11530,N_11835);
and U12263 (N_12263,N_11307,N_11489);
xor U12264 (N_12264,N_11334,N_11261);
xnor U12265 (N_12265,N_11360,N_11091);
or U12266 (N_12266,N_11935,N_11134);
and U12267 (N_12267,N_11073,N_11279);
or U12268 (N_12268,N_11639,N_11080);
nor U12269 (N_12269,N_11963,N_11575);
and U12270 (N_12270,N_11562,N_11698);
and U12271 (N_12271,N_11221,N_11803);
or U12272 (N_12272,N_11982,N_11512);
nand U12273 (N_12273,N_11250,N_11032);
nand U12274 (N_12274,N_11765,N_11942);
xnor U12275 (N_12275,N_11176,N_11647);
and U12276 (N_12276,N_11249,N_11026);
or U12277 (N_12277,N_11871,N_11719);
xor U12278 (N_12278,N_11214,N_11571);
xor U12279 (N_12279,N_11889,N_11457);
or U12280 (N_12280,N_11019,N_11106);
xnor U12281 (N_12281,N_11598,N_11465);
nor U12282 (N_12282,N_11386,N_11381);
nor U12283 (N_12283,N_11504,N_11007);
and U12284 (N_12284,N_11840,N_11503);
or U12285 (N_12285,N_11996,N_11265);
and U12286 (N_12286,N_11910,N_11984);
or U12287 (N_12287,N_11416,N_11505);
nand U12288 (N_12288,N_11243,N_11355);
nand U12289 (N_12289,N_11520,N_11959);
nand U12290 (N_12290,N_11968,N_11606);
nor U12291 (N_12291,N_11965,N_11685);
or U12292 (N_12292,N_11722,N_11546);
nand U12293 (N_12293,N_11814,N_11062);
xor U12294 (N_12294,N_11654,N_11914);
or U12295 (N_12295,N_11623,N_11164);
nand U12296 (N_12296,N_11841,N_11126);
and U12297 (N_12297,N_11308,N_11777);
and U12298 (N_12298,N_11153,N_11150);
nor U12299 (N_12299,N_11885,N_11580);
xnor U12300 (N_12300,N_11882,N_11784);
xor U12301 (N_12301,N_11451,N_11860);
nor U12302 (N_12302,N_11932,N_11686);
or U12303 (N_12303,N_11209,N_11916);
xnor U12304 (N_12304,N_11802,N_11004);
nand U12305 (N_12305,N_11538,N_11447);
nor U12306 (N_12306,N_11413,N_11372);
nor U12307 (N_12307,N_11856,N_11044);
xor U12308 (N_12308,N_11567,N_11426);
or U12309 (N_12309,N_11310,N_11876);
or U12310 (N_12310,N_11102,N_11354);
xor U12311 (N_12311,N_11643,N_11299);
and U12312 (N_12312,N_11594,N_11006);
nor U12313 (N_12313,N_11154,N_11998);
nand U12314 (N_12314,N_11311,N_11148);
nand U12315 (N_12315,N_11110,N_11561);
xnor U12316 (N_12316,N_11622,N_11097);
nor U12317 (N_12317,N_11088,N_11934);
nand U12318 (N_12318,N_11309,N_11036);
and U12319 (N_12319,N_11981,N_11908);
nand U12320 (N_12320,N_11794,N_11710);
or U12321 (N_12321,N_11602,N_11928);
xnor U12322 (N_12322,N_11175,N_11270);
and U12323 (N_12323,N_11655,N_11374);
nand U12324 (N_12324,N_11776,N_11002);
nand U12325 (N_12325,N_11989,N_11292);
nand U12326 (N_12326,N_11011,N_11588);
xor U12327 (N_12327,N_11618,N_11528);
xor U12328 (N_12328,N_11333,N_11461);
nand U12329 (N_12329,N_11415,N_11875);
nor U12330 (N_12330,N_11014,N_11233);
nor U12331 (N_12331,N_11364,N_11254);
and U12332 (N_12332,N_11611,N_11173);
xnor U12333 (N_12333,N_11112,N_11251);
or U12334 (N_12334,N_11715,N_11682);
and U12335 (N_12335,N_11496,N_11720);
or U12336 (N_12336,N_11215,N_11408);
xnor U12337 (N_12337,N_11862,N_11169);
or U12338 (N_12338,N_11615,N_11662);
or U12339 (N_12339,N_11581,N_11206);
nand U12340 (N_12340,N_11370,N_11752);
xnor U12341 (N_12341,N_11092,N_11832);
and U12342 (N_12342,N_11239,N_11116);
nand U12343 (N_12343,N_11194,N_11182);
or U12344 (N_12344,N_11745,N_11949);
nor U12345 (N_12345,N_11143,N_11046);
nand U12346 (N_12346,N_11170,N_11648);
nand U12347 (N_12347,N_11926,N_11147);
nor U12348 (N_12348,N_11300,N_11730);
nor U12349 (N_12349,N_11132,N_11142);
and U12350 (N_12350,N_11190,N_11861);
or U12351 (N_12351,N_11612,N_11634);
xnor U12352 (N_12352,N_11772,N_11086);
nand U12353 (N_12353,N_11460,N_11445);
xor U12354 (N_12354,N_11453,N_11828);
nand U12355 (N_12355,N_11952,N_11440);
and U12356 (N_12356,N_11754,N_11252);
or U12357 (N_12357,N_11591,N_11574);
nor U12358 (N_12358,N_11131,N_11053);
xor U12359 (N_12359,N_11430,N_11409);
nand U12360 (N_12360,N_11852,N_11902);
nor U12361 (N_12361,N_11199,N_11956);
xnor U12362 (N_12362,N_11837,N_11695);
xor U12363 (N_12363,N_11411,N_11056);
nand U12364 (N_12364,N_11473,N_11913);
nor U12365 (N_12365,N_11742,N_11043);
and U12366 (N_12366,N_11849,N_11703);
xor U12367 (N_12367,N_11495,N_11513);
nor U12368 (N_12368,N_11552,N_11979);
nand U12369 (N_12369,N_11377,N_11423);
nand U12370 (N_12370,N_11712,N_11714);
xor U12371 (N_12371,N_11287,N_11326);
xor U12372 (N_12372,N_11759,N_11235);
xor U12373 (N_12373,N_11242,N_11716);
xnor U12374 (N_12374,N_11247,N_11262);
nand U12375 (N_12375,N_11480,N_11509);
or U12376 (N_12376,N_11657,N_11136);
nor U12377 (N_12377,N_11213,N_11572);
and U12378 (N_12378,N_11692,N_11576);
nand U12379 (N_12379,N_11517,N_11617);
and U12380 (N_12380,N_11120,N_11497);
xnor U12381 (N_12381,N_11340,N_11737);
nand U12382 (N_12382,N_11467,N_11245);
nand U12383 (N_12383,N_11544,N_11450);
nor U12384 (N_12384,N_11320,N_11584);
or U12385 (N_12385,N_11748,N_11867);
nand U12386 (N_12386,N_11645,N_11853);
nand U12387 (N_12387,N_11427,N_11069);
nor U12388 (N_12388,N_11872,N_11332);
nor U12389 (N_12389,N_11089,N_11157);
nor U12390 (N_12390,N_11312,N_11614);
nor U12391 (N_12391,N_11527,N_11285);
nand U12392 (N_12392,N_11498,N_11922);
nand U12393 (N_12393,N_11793,N_11536);
nand U12394 (N_12394,N_11749,N_11563);
xor U12395 (N_12395,N_11819,N_11117);
and U12396 (N_12396,N_11412,N_11557);
nor U12397 (N_12397,N_11018,N_11012);
xnor U12398 (N_12398,N_11609,N_11113);
or U12399 (N_12399,N_11122,N_11757);
nand U12400 (N_12400,N_11446,N_11470);
or U12401 (N_12401,N_11894,N_11827);
xor U12402 (N_12402,N_11555,N_11820);
nor U12403 (N_12403,N_11478,N_11560);
nand U12404 (N_12404,N_11854,N_11238);
nand U12405 (N_12405,N_11900,N_11800);
and U12406 (N_12406,N_11761,N_11074);
nand U12407 (N_12407,N_11523,N_11741);
nand U12408 (N_12408,N_11234,N_11972);
and U12409 (N_12409,N_11616,N_11344);
nand U12410 (N_12410,N_11564,N_11096);
and U12411 (N_12411,N_11105,N_11071);
xor U12412 (N_12412,N_11295,N_11055);
or U12413 (N_12413,N_11458,N_11740);
and U12414 (N_12414,N_11886,N_11009);
and U12415 (N_12415,N_11969,N_11224);
or U12416 (N_12416,N_11428,N_11782);
and U12417 (N_12417,N_11833,N_11449);
xnor U12418 (N_12418,N_11668,N_11796);
nor U12419 (N_12419,N_11845,N_11130);
and U12420 (N_12420,N_11553,N_11133);
and U12421 (N_12421,N_11864,N_11079);
nand U12422 (N_12422,N_11025,N_11369);
or U12423 (N_12423,N_11747,N_11181);
xor U12424 (N_12424,N_11589,N_11545);
xnor U12425 (N_12425,N_11118,N_11620);
and U12426 (N_12426,N_11474,N_11652);
xor U12427 (N_12427,N_11883,N_11813);
nor U12428 (N_12428,N_11543,N_11058);
and U12429 (N_12429,N_11425,N_11020);
nor U12430 (N_12430,N_11566,N_11229);
nor U12431 (N_12431,N_11799,N_11673);
xnor U12432 (N_12432,N_11081,N_11477);
xnor U12433 (N_12433,N_11537,N_11059);
nor U12434 (N_12434,N_11302,N_11718);
nand U12435 (N_12435,N_11940,N_11414);
nor U12436 (N_12436,N_11779,N_11535);
nand U12437 (N_12437,N_11067,N_11744);
or U12438 (N_12438,N_11400,N_11964);
or U12439 (N_12439,N_11490,N_11324);
xnor U12440 (N_12440,N_11115,N_11353);
nor U12441 (N_12441,N_11822,N_11884);
or U12442 (N_12442,N_11396,N_11339);
xor U12443 (N_12443,N_11099,N_11967);
and U12444 (N_12444,N_11641,N_11931);
xor U12445 (N_12445,N_11499,N_11593);
xnor U12446 (N_12446,N_11466,N_11336);
xor U12447 (N_12447,N_11976,N_11980);
nand U12448 (N_12448,N_11100,N_11727);
nor U12449 (N_12449,N_11410,N_11241);
or U12450 (N_12450,N_11605,N_11974);
and U12451 (N_12451,N_11829,N_11000);
and U12452 (N_12452,N_11675,N_11699);
and U12453 (N_12453,N_11818,N_11760);
and U12454 (N_12454,N_11762,N_11494);
nand U12455 (N_12455,N_11891,N_11844);
nand U12456 (N_12456,N_11021,N_11029);
nand U12457 (N_12457,N_11084,N_11653);
or U12458 (N_12458,N_11831,N_11613);
xor U12459 (N_12459,N_11220,N_11034);
nor U12460 (N_12460,N_11338,N_11129);
nand U12461 (N_12461,N_11378,N_11268);
nand U12462 (N_12462,N_11347,N_11780);
nor U12463 (N_12463,N_11608,N_11403);
nand U12464 (N_12464,N_11815,N_11848);
or U12465 (N_12465,N_11293,N_11525);
xor U12466 (N_12466,N_11734,N_11266);
xnor U12467 (N_12467,N_11052,N_11297);
and U12468 (N_12468,N_11432,N_11732);
or U12469 (N_12469,N_11755,N_11631);
xnor U12470 (N_12470,N_11399,N_11437);
nor U12471 (N_12471,N_11767,N_11158);
xor U12472 (N_12472,N_11341,N_11709);
xnor U12473 (N_12473,N_11165,N_11405);
xnor U12474 (N_12474,N_11441,N_11166);
xor U12475 (N_12475,N_11592,N_11518);
xnor U12476 (N_12476,N_11948,N_11140);
xor U12477 (N_12477,N_11743,N_11946);
xor U12478 (N_12478,N_11459,N_11256);
xor U12479 (N_12479,N_11999,N_11083);
xor U12480 (N_12480,N_11586,N_11966);
nand U12481 (N_12481,N_11704,N_11228);
or U12482 (N_12482,N_11901,N_11275);
and U12483 (N_12483,N_11866,N_11725);
nand U12484 (N_12484,N_11781,N_11393);
nor U12485 (N_12485,N_11219,N_11398);
xor U12486 (N_12486,N_11708,N_11246);
xnor U12487 (N_12487,N_11821,N_11666);
nor U12488 (N_12488,N_11511,N_11857);
nor U12489 (N_12489,N_11231,N_11271);
nor U12490 (N_12490,N_11197,N_11218);
or U12491 (N_12491,N_11087,N_11314);
nor U12492 (N_12492,N_11493,N_11346);
nand U12493 (N_12493,N_11188,N_11038);
nor U12494 (N_12494,N_11001,N_11816);
nand U12495 (N_12495,N_11958,N_11671);
nor U12496 (N_12496,N_11064,N_11051);
xor U12497 (N_12497,N_11590,N_11993);
nand U12498 (N_12498,N_11301,N_11629);
nor U12499 (N_12499,N_11488,N_11072);
xor U12500 (N_12500,N_11342,N_11509);
nor U12501 (N_12501,N_11545,N_11998);
xnor U12502 (N_12502,N_11931,N_11583);
and U12503 (N_12503,N_11269,N_11877);
xor U12504 (N_12504,N_11420,N_11196);
xor U12505 (N_12505,N_11428,N_11030);
nand U12506 (N_12506,N_11035,N_11419);
or U12507 (N_12507,N_11049,N_11450);
nand U12508 (N_12508,N_11772,N_11091);
nand U12509 (N_12509,N_11893,N_11890);
and U12510 (N_12510,N_11326,N_11252);
xnor U12511 (N_12511,N_11831,N_11675);
nand U12512 (N_12512,N_11180,N_11784);
nor U12513 (N_12513,N_11871,N_11880);
xnor U12514 (N_12514,N_11811,N_11598);
nand U12515 (N_12515,N_11174,N_11680);
xnor U12516 (N_12516,N_11160,N_11977);
nand U12517 (N_12517,N_11405,N_11671);
nand U12518 (N_12518,N_11804,N_11836);
or U12519 (N_12519,N_11396,N_11423);
nor U12520 (N_12520,N_11133,N_11105);
xnor U12521 (N_12521,N_11873,N_11611);
and U12522 (N_12522,N_11369,N_11630);
or U12523 (N_12523,N_11169,N_11312);
nor U12524 (N_12524,N_11418,N_11634);
nand U12525 (N_12525,N_11282,N_11895);
and U12526 (N_12526,N_11443,N_11819);
or U12527 (N_12527,N_11219,N_11704);
or U12528 (N_12528,N_11186,N_11041);
nor U12529 (N_12529,N_11459,N_11038);
or U12530 (N_12530,N_11136,N_11708);
and U12531 (N_12531,N_11505,N_11892);
xor U12532 (N_12532,N_11180,N_11135);
nor U12533 (N_12533,N_11766,N_11945);
nand U12534 (N_12534,N_11686,N_11181);
nor U12535 (N_12535,N_11199,N_11114);
or U12536 (N_12536,N_11058,N_11367);
or U12537 (N_12537,N_11015,N_11957);
xor U12538 (N_12538,N_11328,N_11388);
or U12539 (N_12539,N_11661,N_11035);
nor U12540 (N_12540,N_11030,N_11766);
nor U12541 (N_12541,N_11014,N_11052);
or U12542 (N_12542,N_11281,N_11780);
nor U12543 (N_12543,N_11411,N_11645);
or U12544 (N_12544,N_11873,N_11070);
nand U12545 (N_12545,N_11677,N_11157);
and U12546 (N_12546,N_11533,N_11747);
and U12547 (N_12547,N_11045,N_11072);
nand U12548 (N_12548,N_11681,N_11251);
or U12549 (N_12549,N_11314,N_11504);
xnor U12550 (N_12550,N_11006,N_11400);
or U12551 (N_12551,N_11582,N_11405);
nor U12552 (N_12552,N_11075,N_11510);
nand U12553 (N_12553,N_11916,N_11460);
nand U12554 (N_12554,N_11286,N_11145);
or U12555 (N_12555,N_11086,N_11405);
nand U12556 (N_12556,N_11363,N_11965);
and U12557 (N_12557,N_11318,N_11794);
or U12558 (N_12558,N_11185,N_11836);
nor U12559 (N_12559,N_11979,N_11407);
and U12560 (N_12560,N_11074,N_11144);
nor U12561 (N_12561,N_11165,N_11997);
and U12562 (N_12562,N_11825,N_11422);
and U12563 (N_12563,N_11208,N_11619);
and U12564 (N_12564,N_11994,N_11211);
nand U12565 (N_12565,N_11680,N_11733);
and U12566 (N_12566,N_11903,N_11540);
and U12567 (N_12567,N_11258,N_11750);
xnor U12568 (N_12568,N_11401,N_11799);
or U12569 (N_12569,N_11692,N_11862);
nor U12570 (N_12570,N_11501,N_11685);
and U12571 (N_12571,N_11742,N_11740);
or U12572 (N_12572,N_11572,N_11846);
or U12573 (N_12573,N_11379,N_11381);
and U12574 (N_12574,N_11579,N_11662);
or U12575 (N_12575,N_11189,N_11975);
or U12576 (N_12576,N_11383,N_11987);
and U12577 (N_12577,N_11620,N_11761);
nor U12578 (N_12578,N_11892,N_11276);
or U12579 (N_12579,N_11579,N_11604);
nor U12580 (N_12580,N_11382,N_11338);
nor U12581 (N_12581,N_11320,N_11218);
nor U12582 (N_12582,N_11331,N_11843);
nand U12583 (N_12583,N_11186,N_11673);
and U12584 (N_12584,N_11189,N_11349);
nand U12585 (N_12585,N_11045,N_11784);
or U12586 (N_12586,N_11524,N_11950);
or U12587 (N_12587,N_11999,N_11662);
and U12588 (N_12588,N_11764,N_11351);
nor U12589 (N_12589,N_11378,N_11428);
or U12590 (N_12590,N_11406,N_11884);
nor U12591 (N_12591,N_11793,N_11140);
xor U12592 (N_12592,N_11431,N_11723);
or U12593 (N_12593,N_11013,N_11790);
xor U12594 (N_12594,N_11871,N_11908);
nor U12595 (N_12595,N_11517,N_11844);
xnor U12596 (N_12596,N_11171,N_11180);
nand U12597 (N_12597,N_11309,N_11908);
or U12598 (N_12598,N_11417,N_11370);
xnor U12599 (N_12599,N_11900,N_11949);
xnor U12600 (N_12600,N_11714,N_11066);
nor U12601 (N_12601,N_11018,N_11835);
or U12602 (N_12602,N_11039,N_11752);
nand U12603 (N_12603,N_11973,N_11868);
or U12604 (N_12604,N_11222,N_11878);
nand U12605 (N_12605,N_11690,N_11672);
nand U12606 (N_12606,N_11488,N_11552);
or U12607 (N_12607,N_11231,N_11170);
xnor U12608 (N_12608,N_11476,N_11195);
nor U12609 (N_12609,N_11019,N_11011);
xnor U12610 (N_12610,N_11658,N_11334);
and U12611 (N_12611,N_11890,N_11123);
xor U12612 (N_12612,N_11006,N_11798);
xnor U12613 (N_12613,N_11871,N_11116);
xnor U12614 (N_12614,N_11690,N_11052);
or U12615 (N_12615,N_11794,N_11950);
and U12616 (N_12616,N_11413,N_11401);
nand U12617 (N_12617,N_11182,N_11786);
nand U12618 (N_12618,N_11895,N_11791);
xor U12619 (N_12619,N_11181,N_11169);
nand U12620 (N_12620,N_11565,N_11457);
nor U12621 (N_12621,N_11520,N_11044);
nand U12622 (N_12622,N_11823,N_11731);
or U12623 (N_12623,N_11753,N_11709);
nor U12624 (N_12624,N_11259,N_11373);
or U12625 (N_12625,N_11109,N_11903);
and U12626 (N_12626,N_11198,N_11627);
nand U12627 (N_12627,N_11820,N_11799);
nand U12628 (N_12628,N_11377,N_11718);
xor U12629 (N_12629,N_11921,N_11133);
nand U12630 (N_12630,N_11957,N_11900);
nor U12631 (N_12631,N_11977,N_11085);
xor U12632 (N_12632,N_11320,N_11313);
nor U12633 (N_12633,N_11718,N_11365);
and U12634 (N_12634,N_11059,N_11716);
nand U12635 (N_12635,N_11541,N_11787);
nand U12636 (N_12636,N_11760,N_11747);
nor U12637 (N_12637,N_11732,N_11429);
nor U12638 (N_12638,N_11266,N_11607);
and U12639 (N_12639,N_11656,N_11401);
nor U12640 (N_12640,N_11059,N_11734);
xnor U12641 (N_12641,N_11492,N_11590);
nor U12642 (N_12642,N_11297,N_11333);
nor U12643 (N_12643,N_11267,N_11152);
nand U12644 (N_12644,N_11148,N_11631);
xor U12645 (N_12645,N_11814,N_11047);
nand U12646 (N_12646,N_11610,N_11226);
xor U12647 (N_12647,N_11166,N_11452);
nand U12648 (N_12648,N_11272,N_11855);
xnor U12649 (N_12649,N_11977,N_11814);
nor U12650 (N_12650,N_11009,N_11959);
or U12651 (N_12651,N_11286,N_11733);
nor U12652 (N_12652,N_11063,N_11412);
nor U12653 (N_12653,N_11485,N_11931);
and U12654 (N_12654,N_11597,N_11036);
and U12655 (N_12655,N_11210,N_11665);
and U12656 (N_12656,N_11134,N_11859);
or U12657 (N_12657,N_11833,N_11205);
nor U12658 (N_12658,N_11893,N_11147);
and U12659 (N_12659,N_11290,N_11907);
or U12660 (N_12660,N_11106,N_11145);
and U12661 (N_12661,N_11694,N_11240);
xnor U12662 (N_12662,N_11720,N_11867);
nor U12663 (N_12663,N_11054,N_11901);
xnor U12664 (N_12664,N_11198,N_11086);
nand U12665 (N_12665,N_11448,N_11427);
or U12666 (N_12666,N_11236,N_11950);
nor U12667 (N_12667,N_11209,N_11757);
xor U12668 (N_12668,N_11533,N_11285);
xor U12669 (N_12669,N_11670,N_11930);
xnor U12670 (N_12670,N_11413,N_11987);
nand U12671 (N_12671,N_11465,N_11285);
nor U12672 (N_12672,N_11426,N_11904);
and U12673 (N_12673,N_11231,N_11212);
xnor U12674 (N_12674,N_11073,N_11812);
and U12675 (N_12675,N_11131,N_11207);
xor U12676 (N_12676,N_11193,N_11707);
xnor U12677 (N_12677,N_11424,N_11264);
or U12678 (N_12678,N_11231,N_11050);
and U12679 (N_12679,N_11251,N_11126);
or U12680 (N_12680,N_11769,N_11839);
nor U12681 (N_12681,N_11752,N_11957);
or U12682 (N_12682,N_11027,N_11718);
xnor U12683 (N_12683,N_11540,N_11281);
xnor U12684 (N_12684,N_11731,N_11832);
nand U12685 (N_12685,N_11349,N_11975);
and U12686 (N_12686,N_11516,N_11028);
nand U12687 (N_12687,N_11917,N_11677);
or U12688 (N_12688,N_11502,N_11855);
nor U12689 (N_12689,N_11663,N_11495);
and U12690 (N_12690,N_11424,N_11647);
and U12691 (N_12691,N_11563,N_11263);
or U12692 (N_12692,N_11537,N_11081);
xor U12693 (N_12693,N_11597,N_11741);
and U12694 (N_12694,N_11818,N_11524);
and U12695 (N_12695,N_11448,N_11894);
and U12696 (N_12696,N_11932,N_11927);
or U12697 (N_12697,N_11048,N_11887);
or U12698 (N_12698,N_11526,N_11443);
nand U12699 (N_12699,N_11529,N_11036);
or U12700 (N_12700,N_11034,N_11891);
nor U12701 (N_12701,N_11217,N_11245);
or U12702 (N_12702,N_11705,N_11468);
nor U12703 (N_12703,N_11295,N_11476);
and U12704 (N_12704,N_11153,N_11039);
and U12705 (N_12705,N_11830,N_11106);
nand U12706 (N_12706,N_11848,N_11441);
nor U12707 (N_12707,N_11715,N_11291);
nor U12708 (N_12708,N_11657,N_11832);
nor U12709 (N_12709,N_11740,N_11828);
nand U12710 (N_12710,N_11576,N_11812);
nand U12711 (N_12711,N_11806,N_11792);
nor U12712 (N_12712,N_11173,N_11438);
xnor U12713 (N_12713,N_11792,N_11079);
xor U12714 (N_12714,N_11691,N_11909);
nor U12715 (N_12715,N_11815,N_11491);
nor U12716 (N_12716,N_11089,N_11286);
and U12717 (N_12717,N_11532,N_11190);
xor U12718 (N_12718,N_11043,N_11199);
and U12719 (N_12719,N_11907,N_11613);
xor U12720 (N_12720,N_11948,N_11006);
nand U12721 (N_12721,N_11787,N_11754);
or U12722 (N_12722,N_11186,N_11015);
and U12723 (N_12723,N_11253,N_11863);
or U12724 (N_12724,N_11864,N_11887);
nor U12725 (N_12725,N_11033,N_11312);
xnor U12726 (N_12726,N_11240,N_11108);
and U12727 (N_12727,N_11380,N_11492);
and U12728 (N_12728,N_11168,N_11321);
nor U12729 (N_12729,N_11604,N_11005);
xnor U12730 (N_12730,N_11529,N_11217);
nand U12731 (N_12731,N_11304,N_11496);
xnor U12732 (N_12732,N_11731,N_11191);
nand U12733 (N_12733,N_11429,N_11567);
or U12734 (N_12734,N_11672,N_11969);
and U12735 (N_12735,N_11445,N_11248);
nand U12736 (N_12736,N_11240,N_11690);
xnor U12737 (N_12737,N_11896,N_11110);
xor U12738 (N_12738,N_11537,N_11512);
and U12739 (N_12739,N_11717,N_11805);
and U12740 (N_12740,N_11897,N_11834);
nand U12741 (N_12741,N_11889,N_11452);
or U12742 (N_12742,N_11428,N_11369);
nand U12743 (N_12743,N_11196,N_11715);
nand U12744 (N_12744,N_11777,N_11488);
nand U12745 (N_12745,N_11622,N_11489);
or U12746 (N_12746,N_11921,N_11639);
nor U12747 (N_12747,N_11297,N_11741);
and U12748 (N_12748,N_11964,N_11546);
nor U12749 (N_12749,N_11385,N_11501);
or U12750 (N_12750,N_11806,N_11705);
xnor U12751 (N_12751,N_11340,N_11600);
and U12752 (N_12752,N_11059,N_11068);
or U12753 (N_12753,N_11558,N_11249);
xor U12754 (N_12754,N_11328,N_11207);
or U12755 (N_12755,N_11093,N_11503);
nor U12756 (N_12756,N_11489,N_11898);
and U12757 (N_12757,N_11814,N_11750);
or U12758 (N_12758,N_11354,N_11512);
nand U12759 (N_12759,N_11813,N_11957);
or U12760 (N_12760,N_11021,N_11723);
and U12761 (N_12761,N_11859,N_11237);
and U12762 (N_12762,N_11789,N_11070);
xnor U12763 (N_12763,N_11440,N_11338);
nand U12764 (N_12764,N_11245,N_11859);
nor U12765 (N_12765,N_11792,N_11034);
xnor U12766 (N_12766,N_11198,N_11664);
nand U12767 (N_12767,N_11255,N_11162);
nor U12768 (N_12768,N_11706,N_11217);
nor U12769 (N_12769,N_11918,N_11817);
or U12770 (N_12770,N_11361,N_11946);
nor U12771 (N_12771,N_11739,N_11074);
nor U12772 (N_12772,N_11398,N_11992);
xor U12773 (N_12773,N_11581,N_11805);
and U12774 (N_12774,N_11683,N_11241);
and U12775 (N_12775,N_11225,N_11227);
or U12776 (N_12776,N_11612,N_11726);
xor U12777 (N_12777,N_11815,N_11236);
nand U12778 (N_12778,N_11245,N_11696);
nand U12779 (N_12779,N_11380,N_11674);
xnor U12780 (N_12780,N_11679,N_11236);
and U12781 (N_12781,N_11264,N_11064);
and U12782 (N_12782,N_11796,N_11165);
xnor U12783 (N_12783,N_11329,N_11999);
nand U12784 (N_12784,N_11332,N_11646);
and U12785 (N_12785,N_11799,N_11336);
xor U12786 (N_12786,N_11059,N_11099);
and U12787 (N_12787,N_11540,N_11852);
and U12788 (N_12788,N_11061,N_11165);
xor U12789 (N_12789,N_11808,N_11343);
and U12790 (N_12790,N_11123,N_11695);
nor U12791 (N_12791,N_11284,N_11312);
or U12792 (N_12792,N_11447,N_11208);
and U12793 (N_12793,N_11080,N_11445);
or U12794 (N_12794,N_11407,N_11473);
or U12795 (N_12795,N_11587,N_11460);
or U12796 (N_12796,N_11727,N_11299);
and U12797 (N_12797,N_11767,N_11376);
nor U12798 (N_12798,N_11056,N_11899);
xor U12799 (N_12799,N_11076,N_11888);
or U12800 (N_12800,N_11509,N_11237);
and U12801 (N_12801,N_11631,N_11312);
or U12802 (N_12802,N_11351,N_11101);
or U12803 (N_12803,N_11653,N_11705);
nor U12804 (N_12804,N_11864,N_11373);
nand U12805 (N_12805,N_11548,N_11738);
xor U12806 (N_12806,N_11119,N_11085);
or U12807 (N_12807,N_11263,N_11943);
and U12808 (N_12808,N_11656,N_11635);
or U12809 (N_12809,N_11970,N_11411);
nand U12810 (N_12810,N_11758,N_11095);
or U12811 (N_12811,N_11762,N_11896);
xor U12812 (N_12812,N_11204,N_11422);
xor U12813 (N_12813,N_11332,N_11647);
xnor U12814 (N_12814,N_11409,N_11741);
xnor U12815 (N_12815,N_11236,N_11235);
nor U12816 (N_12816,N_11731,N_11002);
and U12817 (N_12817,N_11403,N_11729);
nor U12818 (N_12818,N_11108,N_11763);
or U12819 (N_12819,N_11601,N_11492);
nand U12820 (N_12820,N_11434,N_11432);
and U12821 (N_12821,N_11896,N_11973);
xnor U12822 (N_12822,N_11229,N_11041);
nand U12823 (N_12823,N_11847,N_11104);
or U12824 (N_12824,N_11402,N_11415);
or U12825 (N_12825,N_11172,N_11041);
xnor U12826 (N_12826,N_11148,N_11983);
xor U12827 (N_12827,N_11053,N_11708);
xnor U12828 (N_12828,N_11396,N_11667);
or U12829 (N_12829,N_11923,N_11648);
and U12830 (N_12830,N_11343,N_11284);
or U12831 (N_12831,N_11742,N_11991);
xor U12832 (N_12832,N_11948,N_11474);
nand U12833 (N_12833,N_11547,N_11399);
nand U12834 (N_12834,N_11717,N_11399);
xnor U12835 (N_12835,N_11760,N_11361);
and U12836 (N_12836,N_11410,N_11640);
and U12837 (N_12837,N_11645,N_11117);
nor U12838 (N_12838,N_11654,N_11778);
nor U12839 (N_12839,N_11085,N_11642);
and U12840 (N_12840,N_11410,N_11590);
or U12841 (N_12841,N_11550,N_11485);
or U12842 (N_12842,N_11763,N_11239);
nand U12843 (N_12843,N_11832,N_11234);
or U12844 (N_12844,N_11600,N_11477);
or U12845 (N_12845,N_11318,N_11899);
nand U12846 (N_12846,N_11717,N_11796);
nor U12847 (N_12847,N_11097,N_11125);
xnor U12848 (N_12848,N_11534,N_11427);
xnor U12849 (N_12849,N_11620,N_11047);
nand U12850 (N_12850,N_11961,N_11797);
or U12851 (N_12851,N_11383,N_11739);
xnor U12852 (N_12852,N_11711,N_11830);
nor U12853 (N_12853,N_11243,N_11459);
or U12854 (N_12854,N_11555,N_11442);
xnor U12855 (N_12855,N_11015,N_11206);
or U12856 (N_12856,N_11810,N_11711);
nor U12857 (N_12857,N_11428,N_11600);
and U12858 (N_12858,N_11642,N_11852);
or U12859 (N_12859,N_11230,N_11630);
and U12860 (N_12860,N_11896,N_11041);
nor U12861 (N_12861,N_11207,N_11530);
and U12862 (N_12862,N_11027,N_11876);
or U12863 (N_12863,N_11198,N_11897);
nor U12864 (N_12864,N_11394,N_11222);
nor U12865 (N_12865,N_11677,N_11418);
and U12866 (N_12866,N_11382,N_11469);
xor U12867 (N_12867,N_11890,N_11770);
or U12868 (N_12868,N_11022,N_11920);
and U12869 (N_12869,N_11102,N_11318);
xnor U12870 (N_12870,N_11485,N_11147);
xnor U12871 (N_12871,N_11194,N_11742);
nor U12872 (N_12872,N_11107,N_11614);
and U12873 (N_12873,N_11098,N_11702);
xor U12874 (N_12874,N_11580,N_11240);
or U12875 (N_12875,N_11620,N_11370);
nand U12876 (N_12876,N_11526,N_11672);
nor U12877 (N_12877,N_11953,N_11229);
or U12878 (N_12878,N_11363,N_11375);
and U12879 (N_12879,N_11659,N_11193);
nor U12880 (N_12880,N_11004,N_11299);
nand U12881 (N_12881,N_11317,N_11491);
nor U12882 (N_12882,N_11897,N_11871);
nand U12883 (N_12883,N_11204,N_11178);
or U12884 (N_12884,N_11201,N_11885);
or U12885 (N_12885,N_11265,N_11094);
xor U12886 (N_12886,N_11540,N_11546);
and U12887 (N_12887,N_11852,N_11806);
xnor U12888 (N_12888,N_11366,N_11097);
nor U12889 (N_12889,N_11337,N_11951);
and U12890 (N_12890,N_11710,N_11941);
and U12891 (N_12891,N_11707,N_11162);
or U12892 (N_12892,N_11293,N_11896);
nor U12893 (N_12893,N_11171,N_11706);
nand U12894 (N_12894,N_11618,N_11504);
nor U12895 (N_12895,N_11744,N_11301);
nand U12896 (N_12896,N_11085,N_11794);
nand U12897 (N_12897,N_11423,N_11545);
or U12898 (N_12898,N_11899,N_11914);
nand U12899 (N_12899,N_11950,N_11863);
xnor U12900 (N_12900,N_11671,N_11825);
and U12901 (N_12901,N_11382,N_11942);
or U12902 (N_12902,N_11651,N_11939);
or U12903 (N_12903,N_11476,N_11165);
or U12904 (N_12904,N_11562,N_11414);
nand U12905 (N_12905,N_11629,N_11966);
or U12906 (N_12906,N_11506,N_11628);
and U12907 (N_12907,N_11431,N_11303);
nand U12908 (N_12908,N_11580,N_11581);
nand U12909 (N_12909,N_11712,N_11469);
xor U12910 (N_12910,N_11607,N_11203);
or U12911 (N_12911,N_11763,N_11770);
xor U12912 (N_12912,N_11258,N_11091);
nand U12913 (N_12913,N_11069,N_11537);
nor U12914 (N_12914,N_11467,N_11310);
nand U12915 (N_12915,N_11648,N_11299);
nand U12916 (N_12916,N_11065,N_11805);
and U12917 (N_12917,N_11816,N_11485);
nand U12918 (N_12918,N_11258,N_11974);
nor U12919 (N_12919,N_11983,N_11445);
and U12920 (N_12920,N_11129,N_11536);
or U12921 (N_12921,N_11443,N_11465);
xnor U12922 (N_12922,N_11651,N_11813);
xnor U12923 (N_12923,N_11422,N_11265);
nand U12924 (N_12924,N_11032,N_11495);
nand U12925 (N_12925,N_11543,N_11898);
xnor U12926 (N_12926,N_11807,N_11933);
and U12927 (N_12927,N_11699,N_11408);
or U12928 (N_12928,N_11615,N_11464);
xor U12929 (N_12929,N_11706,N_11152);
nor U12930 (N_12930,N_11434,N_11746);
nor U12931 (N_12931,N_11596,N_11832);
and U12932 (N_12932,N_11970,N_11541);
nor U12933 (N_12933,N_11675,N_11688);
or U12934 (N_12934,N_11301,N_11026);
nand U12935 (N_12935,N_11291,N_11345);
nor U12936 (N_12936,N_11617,N_11823);
and U12937 (N_12937,N_11887,N_11080);
nor U12938 (N_12938,N_11303,N_11942);
or U12939 (N_12939,N_11204,N_11497);
nor U12940 (N_12940,N_11613,N_11832);
nand U12941 (N_12941,N_11578,N_11122);
and U12942 (N_12942,N_11030,N_11500);
and U12943 (N_12943,N_11787,N_11700);
nand U12944 (N_12944,N_11713,N_11705);
xor U12945 (N_12945,N_11250,N_11828);
nand U12946 (N_12946,N_11390,N_11161);
xor U12947 (N_12947,N_11139,N_11153);
xor U12948 (N_12948,N_11469,N_11764);
or U12949 (N_12949,N_11134,N_11309);
or U12950 (N_12950,N_11801,N_11015);
xor U12951 (N_12951,N_11734,N_11589);
and U12952 (N_12952,N_11106,N_11472);
nand U12953 (N_12953,N_11456,N_11808);
xnor U12954 (N_12954,N_11835,N_11341);
or U12955 (N_12955,N_11064,N_11661);
nor U12956 (N_12956,N_11362,N_11437);
or U12957 (N_12957,N_11017,N_11863);
or U12958 (N_12958,N_11266,N_11972);
or U12959 (N_12959,N_11571,N_11493);
nor U12960 (N_12960,N_11135,N_11713);
or U12961 (N_12961,N_11298,N_11150);
xnor U12962 (N_12962,N_11618,N_11946);
xor U12963 (N_12963,N_11265,N_11365);
nand U12964 (N_12964,N_11100,N_11045);
xor U12965 (N_12965,N_11292,N_11249);
nand U12966 (N_12966,N_11405,N_11173);
and U12967 (N_12967,N_11834,N_11149);
or U12968 (N_12968,N_11678,N_11089);
and U12969 (N_12969,N_11670,N_11377);
and U12970 (N_12970,N_11531,N_11476);
and U12971 (N_12971,N_11911,N_11549);
and U12972 (N_12972,N_11648,N_11021);
and U12973 (N_12973,N_11396,N_11943);
and U12974 (N_12974,N_11518,N_11018);
nor U12975 (N_12975,N_11425,N_11882);
nor U12976 (N_12976,N_11137,N_11538);
nor U12977 (N_12977,N_11700,N_11004);
nor U12978 (N_12978,N_11490,N_11139);
xnor U12979 (N_12979,N_11784,N_11398);
or U12980 (N_12980,N_11291,N_11753);
xor U12981 (N_12981,N_11036,N_11954);
xnor U12982 (N_12982,N_11126,N_11365);
nand U12983 (N_12983,N_11772,N_11715);
nor U12984 (N_12984,N_11872,N_11643);
xnor U12985 (N_12985,N_11359,N_11477);
nor U12986 (N_12986,N_11187,N_11477);
nor U12987 (N_12987,N_11333,N_11995);
nor U12988 (N_12988,N_11019,N_11415);
xor U12989 (N_12989,N_11708,N_11965);
or U12990 (N_12990,N_11686,N_11464);
nor U12991 (N_12991,N_11364,N_11613);
nand U12992 (N_12992,N_11924,N_11875);
nor U12993 (N_12993,N_11990,N_11653);
and U12994 (N_12994,N_11178,N_11340);
and U12995 (N_12995,N_11592,N_11558);
xor U12996 (N_12996,N_11303,N_11906);
and U12997 (N_12997,N_11764,N_11496);
nor U12998 (N_12998,N_11130,N_11076);
xor U12999 (N_12999,N_11943,N_11300);
xor U13000 (N_13000,N_12762,N_12223);
and U13001 (N_13001,N_12264,N_12962);
nand U13002 (N_13002,N_12084,N_12276);
nand U13003 (N_13003,N_12036,N_12180);
nand U13004 (N_13004,N_12746,N_12459);
xor U13005 (N_13005,N_12199,N_12144);
nor U13006 (N_13006,N_12838,N_12862);
or U13007 (N_13007,N_12267,N_12309);
nand U13008 (N_13008,N_12105,N_12121);
nor U13009 (N_13009,N_12617,N_12437);
nor U13010 (N_13010,N_12989,N_12399);
and U13011 (N_13011,N_12873,N_12371);
nor U13012 (N_13012,N_12648,N_12791);
nand U13013 (N_13013,N_12712,N_12628);
xor U13014 (N_13014,N_12137,N_12204);
and U13015 (N_13015,N_12584,N_12577);
and U13016 (N_13016,N_12759,N_12910);
or U13017 (N_13017,N_12284,N_12176);
nand U13018 (N_13018,N_12509,N_12683);
nor U13019 (N_13019,N_12357,N_12414);
or U13020 (N_13020,N_12187,N_12219);
and U13021 (N_13021,N_12956,N_12739);
or U13022 (N_13022,N_12828,N_12321);
nand U13023 (N_13023,N_12556,N_12716);
and U13024 (N_13024,N_12147,N_12880);
xor U13025 (N_13025,N_12570,N_12040);
nor U13026 (N_13026,N_12390,N_12039);
xnor U13027 (N_13027,N_12374,N_12893);
xnor U13028 (N_13028,N_12749,N_12519);
nor U13029 (N_13029,N_12280,N_12117);
or U13030 (N_13030,N_12170,N_12586);
nor U13031 (N_13031,N_12427,N_12768);
nor U13032 (N_13032,N_12614,N_12361);
and U13033 (N_13033,N_12193,N_12903);
or U13034 (N_13034,N_12423,N_12271);
nor U13035 (N_13035,N_12943,N_12005);
xor U13036 (N_13036,N_12813,N_12241);
and U13037 (N_13037,N_12673,N_12191);
xor U13038 (N_13038,N_12334,N_12709);
or U13039 (N_13039,N_12043,N_12184);
nand U13040 (N_13040,N_12328,N_12960);
nand U13041 (N_13041,N_12559,N_12443);
xnor U13042 (N_13042,N_12386,N_12963);
and U13043 (N_13043,N_12777,N_12343);
xnor U13044 (N_13044,N_12229,N_12984);
or U13045 (N_13045,N_12496,N_12185);
and U13046 (N_13046,N_12831,N_12366);
and U13047 (N_13047,N_12168,N_12534);
or U13048 (N_13048,N_12861,N_12125);
nand U13049 (N_13049,N_12625,N_12832);
xnor U13050 (N_13050,N_12844,N_12634);
or U13051 (N_13051,N_12319,N_12588);
and U13052 (N_13052,N_12133,N_12201);
nand U13053 (N_13053,N_12506,N_12672);
or U13054 (N_13054,N_12476,N_12249);
xor U13055 (N_13055,N_12085,N_12014);
or U13056 (N_13056,N_12292,N_12317);
nand U13057 (N_13057,N_12725,N_12700);
nor U13058 (N_13058,N_12901,N_12327);
xnor U13059 (N_13059,N_12607,N_12801);
and U13060 (N_13060,N_12622,N_12073);
xor U13061 (N_13061,N_12999,N_12858);
or U13062 (N_13062,N_12031,N_12574);
nor U13063 (N_13063,N_12575,N_12590);
and U13064 (N_13064,N_12865,N_12104);
and U13065 (N_13065,N_12348,N_12969);
or U13066 (N_13066,N_12800,N_12430);
xor U13067 (N_13067,N_12044,N_12213);
nor U13068 (N_13068,N_12128,N_12781);
xnor U13069 (N_13069,N_12792,N_12312);
xnor U13070 (N_13070,N_12635,N_12825);
and U13071 (N_13071,N_12473,N_12373);
and U13072 (N_13072,N_12690,N_12340);
nor U13073 (N_13073,N_12680,N_12602);
xnor U13074 (N_13074,N_12410,N_12745);
nor U13075 (N_13075,N_12520,N_12472);
xnor U13076 (N_13076,N_12782,N_12632);
nand U13077 (N_13077,N_12130,N_12262);
or U13078 (N_13078,N_12975,N_12403);
xor U13079 (N_13079,N_12543,N_12909);
xor U13080 (N_13080,N_12216,N_12490);
or U13081 (N_13081,N_12082,N_12756);
nand U13082 (N_13082,N_12726,N_12484);
and U13083 (N_13083,N_12320,N_12057);
xor U13084 (N_13084,N_12046,N_12917);
nand U13085 (N_13085,N_12440,N_12697);
nand U13086 (N_13086,N_12851,N_12879);
and U13087 (N_13087,N_12947,N_12689);
nand U13088 (N_13088,N_12899,N_12863);
or U13089 (N_13089,N_12232,N_12834);
or U13090 (N_13090,N_12286,N_12477);
nand U13091 (N_13091,N_12350,N_12765);
xor U13092 (N_13092,N_12704,N_12686);
or U13093 (N_13093,N_12018,N_12959);
nor U13094 (N_13094,N_12000,N_12172);
and U13095 (N_13095,N_12424,N_12681);
or U13096 (N_13096,N_12101,N_12279);
nor U13097 (N_13097,N_12612,N_12937);
and U13098 (N_13098,N_12110,N_12270);
nand U13099 (N_13099,N_12566,N_12408);
or U13100 (N_13100,N_12954,N_12532);
or U13101 (N_13101,N_12789,N_12278);
xor U13102 (N_13102,N_12338,N_12932);
or U13103 (N_13103,N_12670,N_12449);
or U13104 (N_13104,N_12819,N_12375);
and U13105 (N_13105,N_12458,N_12737);
and U13106 (N_13106,N_12835,N_12273);
nand U13107 (N_13107,N_12568,N_12970);
and U13108 (N_13108,N_12977,N_12684);
nor U13109 (N_13109,N_12126,N_12431);
nand U13110 (N_13110,N_12315,N_12064);
or U13111 (N_13111,N_12478,N_12239);
or U13112 (N_13112,N_12878,N_12849);
and U13113 (N_13113,N_12818,N_12146);
nand U13114 (N_13114,N_12240,N_12339);
and U13115 (N_13115,N_12433,N_12994);
nor U13116 (N_13116,N_12491,N_12485);
and U13117 (N_13117,N_12460,N_12653);
nand U13118 (N_13118,N_12479,N_12981);
xor U13119 (N_13119,N_12305,N_12465);
xnor U13120 (N_13120,N_12163,N_12252);
xnor U13121 (N_13121,N_12961,N_12435);
nand U13122 (N_13122,N_12904,N_12676);
and U13123 (N_13123,N_12812,N_12742);
xnor U13124 (N_13124,N_12771,N_12868);
xnor U13125 (N_13125,N_12086,N_12929);
or U13126 (N_13126,N_12523,N_12513);
nand U13127 (N_13127,N_12560,N_12565);
xnor U13128 (N_13128,N_12102,N_12234);
or U13129 (N_13129,N_12555,N_12717);
and U13130 (N_13130,N_12992,N_12799);
nor U13131 (N_13131,N_12921,N_12035);
xnor U13132 (N_13132,N_12811,N_12946);
nand U13133 (N_13133,N_12729,N_12181);
xnor U13134 (N_13134,N_12200,N_12066);
or U13135 (N_13135,N_12353,N_12949);
nand U13136 (N_13136,N_12720,N_12615);
nand U13137 (N_13137,N_12052,N_12450);
or U13138 (N_13138,N_12311,N_12268);
nand U13139 (N_13139,N_12764,N_12597);
nor U13140 (N_13140,N_12222,N_12561);
xnor U13141 (N_13141,N_12623,N_12175);
nor U13142 (N_13142,N_12074,N_12691);
or U13143 (N_13143,N_12820,N_12659);
nor U13144 (N_13144,N_12083,N_12076);
xnor U13145 (N_13145,N_12197,N_12866);
or U13146 (N_13146,N_12589,N_12242);
or U13147 (N_13147,N_12226,N_12441);
or U13148 (N_13148,N_12337,N_12934);
xor U13149 (N_13149,N_12593,N_12770);
nor U13150 (N_13150,N_12752,N_12613);
or U13151 (N_13151,N_12257,N_12627);
nand U13152 (N_13152,N_12224,N_12688);
and U13153 (N_13153,N_12404,N_12349);
nand U13154 (N_13154,N_12498,N_12088);
nor U13155 (N_13155,N_12302,N_12106);
and U13156 (N_13156,N_12029,N_12362);
or U13157 (N_13157,N_12011,N_12129);
or U13158 (N_13158,N_12833,N_12525);
and U13159 (N_13159,N_12058,N_12930);
nor U13160 (N_13160,N_12378,N_12779);
nor U13161 (N_13161,N_12499,N_12528);
or U13162 (N_13162,N_12401,N_12996);
nor U13163 (N_13163,N_12255,N_12277);
nand U13164 (N_13164,N_12293,N_12107);
nor U13165 (N_13165,N_12753,N_12439);
or U13166 (N_13166,N_12462,N_12758);
nand U13167 (N_13167,N_12853,N_12285);
xnor U13168 (N_13168,N_12755,N_12493);
and U13169 (N_13169,N_12398,N_12396);
and U13170 (N_13170,N_12638,N_12821);
nand U13171 (N_13171,N_12581,N_12884);
xor U13172 (N_13172,N_12671,N_12335);
nor U13173 (N_13173,N_12127,N_12227);
nor U13174 (N_13174,N_12322,N_12616);
and U13175 (N_13175,N_12250,N_12160);
xor U13176 (N_13176,N_12776,N_12900);
or U13177 (N_13177,N_12382,N_12457);
nor U13178 (N_13178,N_12134,N_12301);
or U13179 (N_13179,N_12174,N_12489);
xnor U13180 (N_13180,N_12256,N_12149);
nor U13181 (N_13181,N_12010,N_12206);
xnor U13182 (N_13182,N_12140,N_12931);
nand U13183 (N_13183,N_12436,N_12377);
and U13184 (N_13184,N_12678,N_12657);
nor U13185 (N_13185,N_12093,N_12652);
nor U13186 (N_13186,N_12325,N_12631);
nor U13187 (N_13187,N_12620,N_12468);
and U13188 (N_13188,N_12471,N_12874);
and U13189 (N_13189,N_12721,N_12860);
and U13190 (N_13190,N_12188,N_12952);
and U13191 (N_13191,N_12344,N_12171);
nor U13192 (N_13192,N_12854,N_12601);
and U13193 (N_13193,N_12155,N_12061);
nand U13194 (N_13194,N_12150,N_12856);
and U13195 (N_13195,N_12368,N_12573);
nor U13196 (N_13196,N_12906,N_12815);
nor U13197 (N_13197,N_12016,N_12048);
nor U13198 (N_13198,N_12983,N_12416);
or U13199 (N_13199,N_12669,N_12360);
or U13200 (N_13200,N_12703,N_12069);
and U13201 (N_13201,N_12814,N_12936);
or U13202 (N_13202,N_12907,N_12750);
nand U13203 (N_13203,N_12407,N_12097);
or U13204 (N_13204,N_12922,N_12238);
and U13205 (N_13205,N_12001,N_12384);
nand U13206 (N_13206,N_12194,N_12501);
or U13207 (N_13207,N_12394,N_12599);
and U13208 (N_13208,N_12731,N_12875);
nor U13209 (N_13209,N_12692,N_12215);
xor U13210 (N_13210,N_12650,N_12705);
xnor U13211 (N_13211,N_12979,N_12816);
nor U13212 (N_13212,N_12452,N_12540);
xnor U13213 (N_13213,N_12905,N_12913);
nor U13214 (N_13214,N_12619,N_12365);
xor U13215 (N_13215,N_12817,N_12735);
nor U13216 (N_13216,N_12054,N_12898);
xor U13217 (N_13217,N_12651,N_12920);
and U13218 (N_13218,N_12037,N_12113);
and U13219 (N_13219,N_12667,N_12455);
xor U13220 (N_13220,N_12592,N_12164);
nand U13221 (N_13221,N_12707,N_12748);
nand U13222 (N_13222,N_12537,N_12804);
xor U13223 (N_13223,N_12823,N_12050);
or U13224 (N_13224,N_12557,N_12542);
and U13225 (N_13225,N_12274,N_12767);
and U13226 (N_13226,N_12713,N_12316);
nand U13227 (N_13227,N_12212,N_12159);
nor U13228 (N_13228,N_12299,N_12551);
nand U13229 (N_13229,N_12108,N_12087);
nand U13230 (N_13230,N_12153,N_12971);
or U13231 (N_13231,N_12908,N_12028);
and U13232 (N_13232,N_12095,N_12323);
nor U13233 (N_13233,N_12253,N_12774);
xnor U13234 (N_13234,N_12103,N_12483);
nand U13235 (N_13235,N_12045,N_12847);
or U13236 (N_13236,N_12358,N_12552);
and U13237 (N_13237,N_12497,N_12666);
or U13238 (N_13238,N_12655,N_12926);
nor U13239 (N_13239,N_12702,N_12795);
or U13240 (N_13240,N_12914,N_12892);
and U13241 (N_13241,N_12081,N_12665);
nor U13242 (N_13242,N_12355,N_12114);
nor U13243 (N_13243,N_12985,N_12071);
nand U13244 (N_13244,N_12701,N_12237);
xnor U13245 (N_13245,N_12794,N_12236);
xnor U13246 (N_13246,N_12541,N_12143);
nand U13247 (N_13247,N_12600,N_12090);
nand U13248 (N_13248,N_12165,N_12372);
or U13249 (N_13249,N_12392,N_12100);
or U13250 (N_13250,N_12636,N_12679);
and U13251 (N_13251,N_12883,N_12507);
and U13252 (N_13252,N_12972,N_12529);
nand U13253 (N_13253,N_12549,N_12718);
xor U13254 (N_13254,N_12026,N_12783);
or U13255 (N_13255,N_12220,N_12957);
xor U13256 (N_13256,N_12841,N_12002);
nand U13257 (N_13257,N_12848,N_12051);
nand U13258 (N_13258,N_12790,N_12428);
and U13259 (N_13259,N_12797,N_12411);
or U13260 (N_13260,N_12743,N_12662);
nand U13261 (N_13261,N_12230,N_12456);
nand U13262 (N_13262,N_12508,N_12734);
nand U13263 (N_13263,N_12517,N_12166);
or U13264 (N_13264,N_12775,N_12744);
and U13265 (N_13265,N_12864,N_12708);
or U13266 (N_13266,N_12562,N_12829);
nand U13267 (N_13267,N_12550,N_12080);
nand U13268 (N_13268,N_12730,N_12694);
xnor U13269 (N_13269,N_12710,N_12603);
and U13270 (N_13270,N_12618,N_12151);
nand U13271 (N_13271,N_12885,N_12763);
and U13272 (N_13272,N_12805,N_12604);
xnor U13273 (N_13273,N_12939,N_12007);
nor U13274 (N_13274,N_12682,N_12202);
xor U13275 (N_13275,N_12780,N_12421);
and U13276 (N_13276,N_12675,N_12724);
nand U13277 (N_13277,N_12511,N_12630);
and U13278 (N_13278,N_12925,N_12210);
or U13279 (N_13279,N_12515,N_12228);
or U13280 (N_13280,N_12693,N_12024);
nand U13281 (N_13281,N_12023,N_12099);
nor U13282 (N_13282,N_12927,N_12356);
nand U13283 (N_13283,N_12976,N_12442);
nor U13284 (N_13284,N_12809,N_12233);
or U13285 (N_13285,N_12269,N_12189);
or U13286 (N_13286,N_12587,N_12757);
xor U13287 (N_13287,N_12062,N_12647);
nand U13288 (N_13288,N_12945,N_12564);
xnor U13289 (N_13289,N_12626,N_12260);
or U13290 (N_13290,N_12182,N_12870);
and U13291 (N_13291,N_12563,N_12379);
nor U13292 (N_13292,N_12719,N_12649);
nor U13293 (N_13293,N_12367,N_12296);
xnor U13294 (N_13294,N_12598,N_12214);
nor U13295 (N_13295,N_12263,N_12060);
and U13296 (N_13296,N_12928,N_12915);
and U13297 (N_13297,N_12876,N_12987);
and U13298 (N_13298,N_12890,N_12715);
or U13299 (N_13299,N_12142,N_12723);
and U13300 (N_13300,N_12132,N_12736);
nand U13301 (N_13301,N_12881,N_12843);
and U13302 (N_13302,N_12583,N_12123);
nor U13303 (N_13303,N_12119,N_12406);
xor U13304 (N_13304,N_12807,N_12116);
xor U13305 (N_13305,N_12644,N_12092);
nor U13306 (N_13306,N_12594,N_12530);
or U13307 (N_13307,N_12098,N_12872);
or U13308 (N_13308,N_12124,N_12461);
and U13309 (N_13309,N_12243,N_12289);
and U13310 (N_13310,N_12986,N_12266);
or U13311 (N_13311,N_12967,N_12806);
nand U13312 (N_13312,N_12502,N_12706);
or U13313 (N_13313,N_12246,N_12902);
nor U13314 (N_13314,N_12258,N_12030);
and U13315 (N_13315,N_12778,N_12463);
nor U13316 (N_13316,N_12282,N_12536);
or U13317 (N_13317,N_12432,N_12364);
or U13318 (N_13318,N_12342,N_12827);
xnor U13319 (N_13319,N_12609,N_12389);
nand U13320 (N_13320,N_12221,N_12297);
xnor U13321 (N_13321,N_12621,N_12916);
nand U13322 (N_13322,N_12131,N_12487);
nor U13323 (N_13323,N_12475,N_12973);
nand U13324 (N_13324,N_12381,N_12205);
xor U13325 (N_13325,N_12383,N_12646);
nand U13326 (N_13326,N_12068,N_12547);
nor U13327 (N_13327,N_12624,N_12846);
or U13328 (N_13328,N_12156,N_12740);
and U13329 (N_13329,N_12940,N_12310);
xor U13330 (N_13330,N_12162,N_12504);
and U13331 (N_13331,N_12580,N_12235);
and U13332 (N_13332,N_12259,N_12298);
nand U13333 (N_13333,N_12287,N_12409);
and U13334 (N_13334,N_12447,N_12953);
or U13335 (N_13335,N_12065,N_12741);
and U13336 (N_13336,N_12606,N_12538);
and U13337 (N_13337,N_12351,N_12824);
xor U13338 (N_13338,N_12480,N_12695);
nand U13339 (N_13339,N_12579,N_12505);
nand U13340 (N_13340,N_12516,N_12145);
and U13341 (N_13341,N_12047,N_12388);
and U13342 (N_13342,N_12826,N_12330);
nand U13343 (N_13343,N_12845,N_12633);
xnor U13344 (N_13344,N_12111,N_12488);
xor U13345 (N_13345,N_12247,N_12034);
or U13346 (N_13346,N_12535,N_12611);
and U13347 (N_13347,N_12115,N_12272);
xnor U13348 (N_13348,N_12711,N_12642);
or U13349 (N_13349,N_12571,N_12169);
xnor U13350 (N_13350,N_12033,N_12786);
xnor U13351 (N_13351,N_12217,N_12063);
nor U13352 (N_13352,N_12857,N_12558);
and U13353 (N_13353,N_12982,N_12569);
xor U13354 (N_13354,N_12522,N_12072);
and U13355 (N_13355,N_12022,N_12553);
and U13356 (N_13356,N_12290,N_12363);
nand U13357 (N_13357,N_12429,N_12446);
and U13358 (N_13358,N_12347,N_12836);
nand U13359 (N_13359,N_12120,N_12842);
or U13360 (N_13360,N_12313,N_12190);
nand U13361 (N_13361,N_12135,N_12769);
nor U13362 (N_13362,N_12195,N_12218);
xnor U13363 (N_13363,N_12354,N_12211);
nand U13364 (N_13364,N_12696,N_12380);
nand U13365 (N_13365,N_12314,N_12419);
xnor U13366 (N_13366,N_12503,N_12596);
nor U13367 (N_13367,N_12645,N_12078);
nand U13368 (N_13368,N_12722,N_12567);
nor U13369 (N_13369,N_12554,N_12837);
and U13370 (N_13370,N_12248,N_12167);
or U13371 (N_13371,N_12699,N_12225);
xnor U13372 (N_13372,N_12895,N_12948);
or U13373 (N_13373,N_12138,N_12291);
xor U13374 (N_13374,N_12572,N_12674);
nor U13375 (N_13375,N_12840,N_12608);
xor U13376 (N_13376,N_12492,N_12004);
xor U13377 (N_13377,N_12089,N_12988);
and U13378 (N_13378,N_12318,N_12950);
nand U13379 (N_13379,N_12122,N_12610);
xor U13380 (N_13380,N_12454,N_12637);
nor U13381 (N_13381,N_12008,N_12032);
nor U13382 (N_13382,N_12096,N_12965);
and U13383 (N_13383,N_12518,N_12341);
nor U13384 (N_13384,N_12585,N_12482);
or U13385 (N_13385,N_12605,N_12728);
and U13386 (N_13386,N_12346,N_12300);
and U13387 (N_13387,N_12359,N_12867);
xor U13388 (N_13388,N_12798,N_12714);
or U13389 (N_13389,N_12245,N_12685);
nor U13390 (N_13390,N_12896,N_12444);
and U13391 (N_13391,N_12640,N_12053);
and U13392 (N_13392,N_12376,N_12698);
xor U13393 (N_13393,N_12933,N_12042);
xnor U13394 (N_13394,N_12426,N_12148);
nor U13395 (N_13395,N_12387,N_12413);
nor U13396 (N_13396,N_12055,N_12887);
nand U13397 (N_13397,N_12041,N_12882);
and U13398 (N_13398,N_12951,N_12788);
nor U13399 (N_13399,N_12231,N_12370);
xor U13400 (N_13400,N_12332,N_12304);
and U13401 (N_13401,N_12094,N_12793);
or U13402 (N_13402,N_12177,N_12393);
nor U13403 (N_13403,N_12533,N_12510);
and U13404 (N_13404,N_12733,N_12139);
nand U13405 (N_13405,N_12400,N_12486);
nor U13406 (N_13406,N_12467,N_12307);
nand U13407 (N_13407,N_12152,N_12773);
or U13408 (N_13408,N_12027,N_12923);
nand U13409 (N_13409,N_12995,N_12877);
or U13410 (N_13410,N_12500,N_12766);
or U13411 (N_13411,N_12324,N_12891);
xnor U13412 (N_13412,N_12244,N_12495);
or U13413 (N_13413,N_12265,N_12192);
or U13414 (N_13414,N_12118,N_12990);
xnor U13415 (N_13415,N_12539,N_12369);
or U13416 (N_13416,N_12687,N_12281);
or U13417 (N_13417,N_12013,N_12546);
nor U13418 (N_13418,N_12855,N_12514);
nand U13419 (N_13419,N_12869,N_12395);
nor U13420 (N_13420,N_12656,N_12526);
nor U13421 (N_13421,N_12958,N_12158);
and U13422 (N_13422,N_12070,N_12464);
xor U13423 (N_13423,N_12852,N_12944);
or U13424 (N_13424,N_12658,N_12161);
xnor U13425 (N_13425,N_12333,N_12663);
nand U13426 (N_13426,N_12595,N_12196);
or U13427 (N_13427,N_12938,N_12643);
or U13428 (N_13428,N_12056,N_12021);
nand U13429 (N_13429,N_12991,N_12871);
or U13430 (N_13430,N_12306,N_12654);
nand U13431 (N_13431,N_12331,N_12474);
nand U13432 (N_13432,N_12974,N_12438);
or U13433 (N_13433,N_12345,N_12079);
nor U13434 (N_13434,N_12978,N_12154);
xor U13435 (N_13435,N_12294,N_12521);
or U13436 (N_13436,N_12641,N_12402);
or U13437 (N_13437,N_12308,N_12912);
and U13438 (N_13438,N_12303,N_12997);
nor U13439 (N_13439,N_12417,N_12955);
nand U13440 (N_13440,N_12422,N_12075);
nand U13441 (N_13441,N_12415,N_12049);
xor U13442 (N_13442,N_12677,N_12582);
or U13443 (N_13443,N_12391,N_12494);
and U13444 (N_13444,N_12802,N_12787);
and U13445 (N_13445,N_12784,N_12451);
and U13446 (N_13446,N_12059,N_12548);
nand U13447 (N_13447,N_12006,N_12209);
xnor U13448 (N_13448,N_12747,N_12003);
or U13449 (N_13449,N_12664,N_12295);
and U13450 (N_13450,N_12412,N_12980);
nand U13451 (N_13451,N_12803,N_12668);
and U13452 (N_13452,N_12109,N_12183);
and U13453 (N_13453,N_12157,N_12434);
and U13454 (N_13454,N_12760,N_12918);
nand U13455 (N_13455,N_12445,N_12919);
and U13456 (N_13456,N_12329,N_12077);
nand U13457 (N_13457,N_12009,N_12326);
nor U13458 (N_13458,N_12179,N_12888);
nor U13459 (N_13459,N_12136,N_12025);
xnor U13460 (N_13460,N_12942,N_12141);
xor U13461 (N_13461,N_12527,N_12397);
nor U13462 (N_13462,N_12186,N_12481);
nor U13463 (N_13463,N_12288,N_12275);
or U13464 (N_13464,N_12545,N_12886);
or U13465 (N_13465,N_12531,N_12810);
nor U13466 (N_13466,N_12894,N_12203);
xnor U13467 (N_13467,N_12038,N_12576);
xnor U13468 (N_13468,N_12578,N_12660);
nand U13469 (N_13469,N_12067,N_12254);
and U13470 (N_13470,N_12448,N_12661);
nor U13471 (N_13471,N_12850,N_12017);
xor U13472 (N_13472,N_12208,N_12207);
nand U13473 (N_13473,N_12941,N_12998);
nand U13474 (N_13474,N_12889,N_12966);
nor U13475 (N_13475,N_12897,N_12352);
and U13476 (N_13476,N_12924,N_12993);
nand U13477 (N_13477,N_12859,N_12420);
or U13478 (N_13478,N_12512,N_12470);
nor U13479 (N_13479,N_12751,N_12466);
or U13480 (N_13480,N_12453,N_12385);
nor U13481 (N_13481,N_12754,N_12732);
nand U13482 (N_13482,N_12012,N_12761);
xor U13483 (N_13483,N_12251,N_12808);
and U13484 (N_13484,N_12418,N_12591);
or U13485 (N_13485,N_12830,N_12968);
and U13486 (N_13486,N_12822,N_12839);
nor U13487 (N_13487,N_12935,N_12772);
or U13488 (N_13488,N_12020,N_12178);
nand U13489 (N_13489,N_12544,N_12336);
or U13490 (N_13490,N_12112,N_12785);
or U13491 (N_13491,N_12173,N_12524);
and U13492 (N_13492,N_12727,N_12639);
xor U13493 (N_13493,N_12425,N_12015);
xnor U13494 (N_13494,N_12738,N_12405);
xnor U13495 (N_13495,N_12261,N_12911);
or U13496 (N_13496,N_12019,N_12469);
nand U13497 (N_13497,N_12198,N_12629);
or U13498 (N_13498,N_12796,N_12091);
and U13499 (N_13499,N_12283,N_12964);
and U13500 (N_13500,N_12289,N_12124);
xor U13501 (N_13501,N_12205,N_12142);
and U13502 (N_13502,N_12893,N_12813);
nand U13503 (N_13503,N_12154,N_12238);
nor U13504 (N_13504,N_12805,N_12495);
and U13505 (N_13505,N_12357,N_12592);
nand U13506 (N_13506,N_12644,N_12048);
or U13507 (N_13507,N_12241,N_12607);
nand U13508 (N_13508,N_12392,N_12483);
xor U13509 (N_13509,N_12922,N_12484);
xnor U13510 (N_13510,N_12177,N_12789);
and U13511 (N_13511,N_12847,N_12275);
nor U13512 (N_13512,N_12464,N_12437);
or U13513 (N_13513,N_12035,N_12756);
nand U13514 (N_13514,N_12242,N_12139);
and U13515 (N_13515,N_12479,N_12964);
nor U13516 (N_13516,N_12078,N_12402);
nand U13517 (N_13517,N_12084,N_12435);
and U13518 (N_13518,N_12969,N_12529);
and U13519 (N_13519,N_12890,N_12816);
and U13520 (N_13520,N_12552,N_12176);
nor U13521 (N_13521,N_12767,N_12458);
xnor U13522 (N_13522,N_12472,N_12205);
xor U13523 (N_13523,N_12506,N_12017);
or U13524 (N_13524,N_12446,N_12663);
or U13525 (N_13525,N_12890,N_12901);
and U13526 (N_13526,N_12849,N_12324);
xor U13527 (N_13527,N_12592,N_12319);
nor U13528 (N_13528,N_12619,N_12432);
or U13529 (N_13529,N_12467,N_12860);
nand U13530 (N_13530,N_12734,N_12323);
and U13531 (N_13531,N_12249,N_12178);
or U13532 (N_13532,N_12873,N_12245);
or U13533 (N_13533,N_12079,N_12019);
xnor U13534 (N_13534,N_12893,N_12205);
nor U13535 (N_13535,N_12133,N_12234);
nand U13536 (N_13536,N_12277,N_12631);
nor U13537 (N_13537,N_12134,N_12818);
nor U13538 (N_13538,N_12780,N_12864);
xnor U13539 (N_13539,N_12659,N_12393);
nor U13540 (N_13540,N_12490,N_12004);
or U13541 (N_13541,N_12019,N_12386);
nand U13542 (N_13542,N_12369,N_12940);
nand U13543 (N_13543,N_12585,N_12373);
and U13544 (N_13544,N_12071,N_12619);
nor U13545 (N_13545,N_12766,N_12835);
or U13546 (N_13546,N_12780,N_12846);
and U13547 (N_13547,N_12358,N_12953);
or U13548 (N_13548,N_12735,N_12297);
nand U13549 (N_13549,N_12666,N_12241);
xnor U13550 (N_13550,N_12629,N_12564);
nor U13551 (N_13551,N_12120,N_12466);
nand U13552 (N_13552,N_12727,N_12477);
or U13553 (N_13553,N_12351,N_12963);
nor U13554 (N_13554,N_12006,N_12448);
or U13555 (N_13555,N_12313,N_12252);
nor U13556 (N_13556,N_12462,N_12096);
nand U13557 (N_13557,N_12621,N_12963);
or U13558 (N_13558,N_12711,N_12508);
or U13559 (N_13559,N_12973,N_12178);
or U13560 (N_13560,N_12273,N_12344);
or U13561 (N_13561,N_12861,N_12897);
and U13562 (N_13562,N_12847,N_12990);
nand U13563 (N_13563,N_12965,N_12645);
or U13564 (N_13564,N_12029,N_12546);
nor U13565 (N_13565,N_12741,N_12166);
nand U13566 (N_13566,N_12334,N_12613);
nand U13567 (N_13567,N_12895,N_12646);
xor U13568 (N_13568,N_12828,N_12432);
nor U13569 (N_13569,N_12108,N_12521);
and U13570 (N_13570,N_12291,N_12372);
or U13571 (N_13571,N_12125,N_12694);
nor U13572 (N_13572,N_12951,N_12900);
or U13573 (N_13573,N_12838,N_12889);
nand U13574 (N_13574,N_12777,N_12378);
xnor U13575 (N_13575,N_12414,N_12411);
nor U13576 (N_13576,N_12564,N_12379);
nor U13577 (N_13577,N_12980,N_12063);
nand U13578 (N_13578,N_12745,N_12186);
or U13579 (N_13579,N_12915,N_12568);
xnor U13580 (N_13580,N_12177,N_12413);
and U13581 (N_13581,N_12965,N_12098);
nand U13582 (N_13582,N_12475,N_12453);
and U13583 (N_13583,N_12479,N_12892);
and U13584 (N_13584,N_12963,N_12237);
and U13585 (N_13585,N_12138,N_12062);
xor U13586 (N_13586,N_12586,N_12139);
xnor U13587 (N_13587,N_12947,N_12061);
and U13588 (N_13588,N_12856,N_12097);
nor U13589 (N_13589,N_12049,N_12796);
nand U13590 (N_13590,N_12521,N_12304);
xnor U13591 (N_13591,N_12114,N_12213);
nand U13592 (N_13592,N_12756,N_12079);
and U13593 (N_13593,N_12210,N_12577);
nand U13594 (N_13594,N_12405,N_12823);
or U13595 (N_13595,N_12912,N_12200);
xor U13596 (N_13596,N_12416,N_12683);
xnor U13597 (N_13597,N_12568,N_12874);
nand U13598 (N_13598,N_12302,N_12524);
xor U13599 (N_13599,N_12889,N_12750);
or U13600 (N_13600,N_12424,N_12010);
or U13601 (N_13601,N_12441,N_12422);
or U13602 (N_13602,N_12983,N_12819);
nor U13603 (N_13603,N_12740,N_12708);
or U13604 (N_13604,N_12515,N_12964);
xnor U13605 (N_13605,N_12073,N_12973);
or U13606 (N_13606,N_12363,N_12354);
nor U13607 (N_13607,N_12153,N_12956);
and U13608 (N_13608,N_12577,N_12166);
nand U13609 (N_13609,N_12166,N_12665);
and U13610 (N_13610,N_12692,N_12509);
and U13611 (N_13611,N_12434,N_12314);
nand U13612 (N_13612,N_12684,N_12561);
nor U13613 (N_13613,N_12144,N_12406);
xor U13614 (N_13614,N_12280,N_12935);
nand U13615 (N_13615,N_12587,N_12850);
or U13616 (N_13616,N_12272,N_12947);
and U13617 (N_13617,N_12830,N_12573);
xnor U13618 (N_13618,N_12064,N_12887);
nand U13619 (N_13619,N_12706,N_12231);
or U13620 (N_13620,N_12519,N_12587);
xor U13621 (N_13621,N_12701,N_12091);
xor U13622 (N_13622,N_12304,N_12046);
or U13623 (N_13623,N_12479,N_12286);
or U13624 (N_13624,N_12992,N_12254);
nor U13625 (N_13625,N_12711,N_12638);
and U13626 (N_13626,N_12519,N_12113);
and U13627 (N_13627,N_12299,N_12423);
and U13628 (N_13628,N_12525,N_12674);
nand U13629 (N_13629,N_12112,N_12248);
nor U13630 (N_13630,N_12124,N_12405);
nand U13631 (N_13631,N_12117,N_12922);
and U13632 (N_13632,N_12308,N_12116);
nand U13633 (N_13633,N_12181,N_12027);
nor U13634 (N_13634,N_12926,N_12487);
nor U13635 (N_13635,N_12179,N_12047);
or U13636 (N_13636,N_12014,N_12543);
and U13637 (N_13637,N_12966,N_12208);
and U13638 (N_13638,N_12236,N_12697);
or U13639 (N_13639,N_12738,N_12234);
xnor U13640 (N_13640,N_12579,N_12590);
xnor U13641 (N_13641,N_12424,N_12584);
nand U13642 (N_13642,N_12542,N_12454);
or U13643 (N_13643,N_12180,N_12743);
nand U13644 (N_13644,N_12170,N_12863);
nor U13645 (N_13645,N_12975,N_12136);
nand U13646 (N_13646,N_12669,N_12130);
or U13647 (N_13647,N_12245,N_12358);
nand U13648 (N_13648,N_12358,N_12653);
nand U13649 (N_13649,N_12483,N_12338);
xnor U13650 (N_13650,N_12516,N_12819);
and U13651 (N_13651,N_12450,N_12024);
xnor U13652 (N_13652,N_12794,N_12042);
nand U13653 (N_13653,N_12944,N_12868);
and U13654 (N_13654,N_12402,N_12565);
and U13655 (N_13655,N_12708,N_12964);
nor U13656 (N_13656,N_12532,N_12094);
nor U13657 (N_13657,N_12625,N_12945);
and U13658 (N_13658,N_12394,N_12359);
nor U13659 (N_13659,N_12634,N_12864);
xnor U13660 (N_13660,N_12801,N_12133);
or U13661 (N_13661,N_12046,N_12499);
and U13662 (N_13662,N_12726,N_12806);
or U13663 (N_13663,N_12127,N_12224);
xor U13664 (N_13664,N_12168,N_12532);
and U13665 (N_13665,N_12403,N_12474);
nand U13666 (N_13666,N_12344,N_12951);
nand U13667 (N_13667,N_12648,N_12426);
or U13668 (N_13668,N_12336,N_12194);
xnor U13669 (N_13669,N_12974,N_12609);
and U13670 (N_13670,N_12903,N_12099);
or U13671 (N_13671,N_12434,N_12771);
or U13672 (N_13672,N_12101,N_12463);
or U13673 (N_13673,N_12975,N_12813);
and U13674 (N_13674,N_12119,N_12570);
nor U13675 (N_13675,N_12762,N_12707);
nor U13676 (N_13676,N_12236,N_12596);
or U13677 (N_13677,N_12146,N_12250);
xor U13678 (N_13678,N_12274,N_12307);
or U13679 (N_13679,N_12146,N_12525);
and U13680 (N_13680,N_12178,N_12352);
nand U13681 (N_13681,N_12172,N_12355);
nand U13682 (N_13682,N_12055,N_12568);
and U13683 (N_13683,N_12020,N_12419);
nor U13684 (N_13684,N_12625,N_12757);
nor U13685 (N_13685,N_12907,N_12392);
nand U13686 (N_13686,N_12455,N_12236);
xor U13687 (N_13687,N_12604,N_12357);
or U13688 (N_13688,N_12245,N_12135);
or U13689 (N_13689,N_12316,N_12547);
xnor U13690 (N_13690,N_12278,N_12492);
or U13691 (N_13691,N_12225,N_12176);
xor U13692 (N_13692,N_12914,N_12997);
and U13693 (N_13693,N_12035,N_12339);
and U13694 (N_13694,N_12591,N_12022);
or U13695 (N_13695,N_12799,N_12514);
and U13696 (N_13696,N_12888,N_12344);
or U13697 (N_13697,N_12459,N_12659);
or U13698 (N_13698,N_12494,N_12549);
and U13699 (N_13699,N_12007,N_12537);
or U13700 (N_13700,N_12487,N_12343);
nand U13701 (N_13701,N_12529,N_12836);
xnor U13702 (N_13702,N_12188,N_12517);
nor U13703 (N_13703,N_12711,N_12955);
or U13704 (N_13704,N_12798,N_12029);
and U13705 (N_13705,N_12154,N_12410);
nor U13706 (N_13706,N_12111,N_12266);
nand U13707 (N_13707,N_12610,N_12921);
xor U13708 (N_13708,N_12617,N_12926);
and U13709 (N_13709,N_12841,N_12754);
nor U13710 (N_13710,N_12306,N_12814);
xnor U13711 (N_13711,N_12369,N_12635);
xnor U13712 (N_13712,N_12198,N_12904);
nor U13713 (N_13713,N_12322,N_12988);
and U13714 (N_13714,N_12797,N_12466);
nand U13715 (N_13715,N_12943,N_12487);
nor U13716 (N_13716,N_12120,N_12452);
xnor U13717 (N_13717,N_12146,N_12485);
xnor U13718 (N_13718,N_12191,N_12690);
nor U13719 (N_13719,N_12588,N_12039);
nand U13720 (N_13720,N_12937,N_12051);
nand U13721 (N_13721,N_12370,N_12034);
nor U13722 (N_13722,N_12492,N_12843);
nand U13723 (N_13723,N_12058,N_12390);
and U13724 (N_13724,N_12264,N_12991);
nor U13725 (N_13725,N_12295,N_12913);
nor U13726 (N_13726,N_12073,N_12157);
and U13727 (N_13727,N_12796,N_12729);
nand U13728 (N_13728,N_12547,N_12376);
xor U13729 (N_13729,N_12538,N_12375);
xor U13730 (N_13730,N_12101,N_12776);
and U13731 (N_13731,N_12300,N_12335);
or U13732 (N_13732,N_12475,N_12918);
nand U13733 (N_13733,N_12598,N_12267);
nand U13734 (N_13734,N_12109,N_12650);
and U13735 (N_13735,N_12408,N_12072);
and U13736 (N_13736,N_12431,N_12913);
nor U13737 (N_13737,N_12854,N_12685);
or U13738 (N_13738,N_12920,N_12954);
and U13739 (N_13739,N_12907,N_12627);
or U13740 (N_13740,N_12599,N_12416);
xnor U13741 (N_13741,N_12270,N_12868);
or U13742 (N_13742,N_12138,N_12159);
or U13743 (N_13743,N_12244,N_12660);
nor U13744 (N_13744,N_12360,N_12409);
or U13745 (N_13745,N_12593,N_12645);
or U13746 (N_13746,N_12171,N_12521);
or U13747 (N_13747,N_12173,N_12910);
xor U13748 (N_13748,N_12448,N_12380);
nand U13749 (N_13749,N_12960,N_12419);
and U13750 (N_13750,N_12960,N_12742);
and U13751 (N_13751,N_12541,N_12657);
nand U13752 (N_13752,N_12624,N_12941);
nor U13753 (N_13753,N_12472,N_12933);
nand U13754 (N_13754,N_12576,N_12740);
and U13755 (N_13755,N_12282,N_12118);
or U13756 (N_13756,N_12956,N_12150);
nor U13757 (N_13757,N_12463,N_12905);
and U13758 (N_13758,N_12572,N_12143);
xnor U13759 (N_13759,N_12527,N_12922);
nor U13760 (N_13760,N_12386,N_12722);
nor U13761 (N_13761,N_12446,N_12112);
nor U13762 (N_13762,N_12357,N_12369);
xnor U13763 (N_13763,N_12769,N_12363);
nand U13764 (N_13764,N_12238,N_12639);
and U13765 (N_13765,N_12027,N_12702);
and U13766 (N_13766,N_12180,N_12161);
xor U13767 (N_13767,N_12438,N_12026);
or U13768 (N_13768,N_12340,N_12398);
nor U13769 (N_13769,N_12450,N_12887);
and U13770 (N_13770,N_12909,N_12937);
nand U13771 (N_13771,N_12385,N_12340);
xnor U13772 (N_13772,N_12560,N_12205);
xor U13773 (N_13773,N_12914,N_12915);
nand U13774 (N_13774,N_12239,N_12350);
xor U13775 (N_13775,N_12853,N_12304);
and U13776 (N_13776,N_12408,N_12294);
nor U13777 (N_13777,N_12423,N_12901);
and U13778 (N_13778,N_12515,N_12083);
or U13779 (N_13779,N_12410,N_12752);
xnor U13780 (N_13780,N_12327,N_12889);
and U13781 (N_13781,N_12854,N_12954);
and U13782 (N_13782,N_12135,N_12019);
xor U13783 (N_13783,N_12418,N_12130);
nand U13784 (N_13784,N_12341,N_12706);
or U13785 (N_13785,N_12434,N_12879);
nand U13786 (N_13786,N_12811,N_12835);
nor U13787 (N_13787,N_12528,N_12500);
nand U13788 (N_13788,N_12388,N_12492);
nor U13789 (N_13789,N_12125,N_12520);
and U13790 (N_13790,N_12325,N_12092);
nand U13791 (N_13791,N_12624,N_12285);
xor U13792 (N_13792,N_12047,N_12963);
nand U13793 (N_13793,N_12387,N_12078);
and U13794 (N_13794,N_12648,N_12995);
or U13795 (N_13795,N_12341,N_12556);
or U13796 (N_13796,N_12018,N_12990);
or U13797 (N_13797,N_12917,N_12285);
or U13798 (N_13798,N_12736,N_12959);
nand U13799 (N_13799,N_12065,N_12506);
nand U13800 (N_13800,N_12427,N_12686);
and U13801 (N_13801,N_12730,N_12738);
or U13802 (N_13802,N_12800,N_12598);
xor U13803 (N_13803,N_12535,N_12599);
nand U13804 (N_13804,N_12544,N_12282);
or U13805 (N_13805,N_12811,N_12500);
nor U13806 (N_13806,N_12759,N_12095);
xor U13807 (N_13807,N_12725,N_12568);
or U13808 (N_13808,N_12567,N_12841);
xnor U13809 (N_13809,N_12264,N_12496);
nand U13810 (N_13810,N_12923,N_12828);
or U13811 (N_13811,N_12460,N_12034);
nor U13812 (N_13812,N_12409,N_12558);
nand U13813 (N_13813,N_12209,N_12318);
nor U13814 (N_13814,N_12828,N_12004);
and U13815 (N_13815,N_12528,N_12356);
or U13816 (N_13816,N_12394,N_12361);
nor U13817 (N_13817,N_12470,N_12460);
or U13818 (N_13818,N_12880,N_12092);
nand U13819 (N_13819,N_12452,N_12019);
nor U13820 (N_13820,N_12670,N_12116);
xnor U13821 (N_13821,N_12323,N_12524);
nor U13822 (N_13822,N_12002,N_12129);
nor U13823 (N_13823,N_12030,N_12453);
nor U13824 (N_13824,N_12980,N_12226);
and U13825 (N_13825,N_12825,N_12552);
and U13826 (N_13826,N_12414,N_12207);
or U13827 (N_13827,N_12602,N_12091);
nand U13828 (N_13828,N_12700,N_12777);
or U13829 (N_13829,N_12771,N_12581);
nand U13830 (N_13830,N_12674,N_12834);
or U13831 (N_13831,N_12542,N_12943);
nand U13832 (N_13832,N_12517,N_12668);
nor U13833 (N_13833,N_12825,N_12760);
xnor U13834 (N_13834,N_12893,N_12077);
nand U13835 (N_13835,N_12094,N_12572);
or U13836 (N_13836,N_12740,N_12028);
and U13837 (N_13837,N_12974,N_12729);
nand U13838 (N_13838,N_12414,N_12189);
nor U13839 (N_13839,N_12375,N_12751);
nor U13840 (N_13840,N_12966,N_12745);
and U13841 (N_13841,N_12528,N_12886);
or U13842 (N_13842,N_12699,N_12693);
nand U13843 (N_13843,N_12700,N_12431);
and U13844 (N_13844,N_12121,N_12128);
nand U13845 (N_13845,N_12420,N_12058);
nor U13846 (N_13846,N_12720,N_12603);
nand U13847 (N_13847,N_12849,N_12421);
nand U13848 (N_13848,N_12121,N_12954);
nor U13849 (N_13849,N_12376,N_12827);
and U13850 (N_13850,N_12290,N_12660);
nand U13851 (N_13851,N_12917,N_12682);
or U13852 (N_13852,N_12681,N_12293);
nand U13853 (N_13853,N_12711,N_12160);
and U13854 (N_13854,N_12465,N_12403);
xnor U13855 (N_13855,N_12341,N_12811);
xnor U13856 (N_13856,N_12983,N_12901);
or U13857 (N_13857,N_12505,N_12260);
or U13858 (N_13858,N_12552,N_12435);
nand U13859 (N_13859,N_12842,N_12756);
nor U13860 (N_13860,N_12907,N_12099);
and U13861 (N_13861,N_12789,N_12225);
and U13862 (N_13862,N_12953,N_12877);
xnor U13863 (N_13863,N_12587,N_12468);
and U13864 (N_13864,N_12184,N_12112);
xor U13865 (N_13865,N_12349,N_12854);
and U13866 (N_13866,N_12246,N_12001);
nor U13867 (N_13867,N_12633,N_12076);
xor U13868 (N_13868,N_12127,N_12077);
nand U13869 (N_13869,N_12973,N_12428);
nand U13870 (N_13870,N_12401,N_12857);
nand U13871 (N_13871,N_12896,N_12775);
nand U13872 (N_13872,N_12637,N_12262);
or U13873 (N_13873,N_12722,N_12009);
nand U13874 (N_13874,N_12234,N_12690);
or U13875 (N_13875,N_12631,N_12970);
xnor U13876 (N_13876,N_12892,N_12253);
nand U13877 (N_13877,N_12526,N_12912);
and U13878 (N_13878,N_12819,N_12820);
nor U13879 (N_13879,N_12335,N_12301);
nand U13880 (N_13880,N_12837,N_12570);
nand U13881 (N_13881,N_12924,N_12773);
nand U13882 (N_13882,N_12720,N_12343);
and U13883 (N_13883,N_12306,N_12614);
nor U13884 (N_13884,N_12142,N_12257);
and U13885 (N_13885,N_12316,N_12072);
nand U13886 (N_13886,N_12360,N_12811);
nor U13887 (N_13887,N_12893,N_12038);
xnor U13888 (N_13888,N_12722,N_12526);
or U13889 (N_13889,N_12640,N_12884);
nand U13890 (N_13890,N_12212,N_12220);
or U13891 (N_13891,N_12692,N_12701);
or U13892 (N_13892,N_12362,N_12001);
nor U13893 (N_13893,N_12363,N_12476);
or U13894 (N_13894,N_12816,N_12683);
or U13895 (N_13895,N_12159,N_12437);
xor U13896 (N_13896,N_12539,N_12845);
nor U13897 (N_13897,N_12497,N_12631);
and U13898 (N_13898,N_12849,N_12024);
nor U13899 (N_13899,N_12448,N_12557);
xnor U13900 (N_13900,N_12007,N_12501);
nor U13901 (N_13901,N_12192,N_12149);
or U13902 (N_13902,N_12967,N_12127);
or U13903 (N_13903,N_12829,N_12422);
or U13904 (N_13904,N_12420,N_12631);
nor U13905 (N_13905,N_12056,N_12061);
or U13906 (N_13906,N_12893,N_12928);
xnor U13907 (N_13907,N_12577,N_12548);
or U13908 (N_13908,N_12121,N_12932);
nor U13909 (N_13909,N_12018,N_12539);
xnor U13910 (N_13910,N_12149,N_12202);
nand U13911 (N_13911,N_12583,N_12749);
nor U13912 (N_13912,N_12784,N_12279);
nand U13913 (N_13913,N_12298,N_12961);
or U13914 (N_13914,N_12939,N_12993);
nand U13915 (N_13915,N_12007,N_12239);
and U13916 (N_13916,N_12961,N_12170);
or U13917 (N_13917,N_12734,N_12979);
nand U13918 (N_13918,N_12323,N_12038);
nand U13919 (N_13919,N_12379,N_12441);
nor U13920 (N_13920,N_12611,N_12149);
xnor U13921 (N_13921,N_12291,N_12249);
nor U13922 (N_13922,N_12026,N_12113);
xnor U13923 (N_13923,N_12574,N_12169);
or U13924 (N_13924,N_12221,N_12761);
xnor U13925 (N_13925,N_12441,N_12286);
xnor U13926 (N_13926,N_12045,N_12437);
xnor U13927 (N_13927,N_12090,N_12827);
nand U13928 (N_13928,N_12773,N_12738);
and U13929 (N_13929,N_12469,N_12422);
nor U13930 (N_13930,N_12654,N_12408);
xnor U13931 (N_13931,N_12116,N_12635);
or U13932 (N_13932,N_12235,N_12976);
and U13933 (N_13933,N_12292,N_12116);
xor U13934 (N_13934,N_12203,N_12218);
nand U13935 (N_13935,N_12316,N_12329);
nand U13936 (N_13936,N_12813,N_12208);
xnor U13937 (N_13937,N_12138,N_12111);
or U13938 (N_13938,N_12750,N_12125);
xnor U13939 (N_13939,N_12776,N_12745);
or U13940 (N_13940,N_12933,N_12529);
xnor U13941 (N_13941,N_12128,N_12728);
xor U13942 (N_13942,N_12168,N_12290);
xor U13943 (N_13943,N_12545,N_12113);
and U13944 (N_13944,N_12912,N_12077);
xnor U13945 (N_13945,N_12798,N_12459);
nand U13946 (N_13946,N_12731,N_12108);
and U13947 (N_13947,N_12587,N_12789);
or U13948 (N_13948,N_12336,N_12520);
nand U13949 (N_13949,N_12931,N_12612);
and U13950 (N_13950,N_12530,N_12741);
xnor U13951 (N_13951,N_12774,N_12079);
nor U13952 (N_13952,N_12380,N_12639);
or U13953 (N_13953,N_12453,N_12936);
xnor U13954 (N_13954,N_12218,N_12331);
or U13955 (N_13955,N_12137,N_12408);
nand U13956 (N_13956,N_12309,N_12985);
nor U13957 (N_13957,N_12054,N_12462);
and U13958 (N_13958,N_12651,N_12005);
and U13959 (N_13959,N_12698,N_12935);
or U13960 (N_13960,N_12889,N_12488);
and U13961 (N_13961,N_12809,N_12508);
and U13962 (N_13962,N_12896,N_12310);
nor U13963 (N_13963,N_12112,N_12996);
xor U13964 (N_13964,N_12269,N_12265);
xnor U13965 (N_13965,N_12640,N_12969);
nor U13966 (N_13966,N_12071,N_12742);
nand U13967 (N_13967,N_12307,N_12123);
nor U13968 (N_13968,N_12910,N_12765);
or U13969 (N_13969,N_12400,N_12385);
or U13970 (N_13970,N_12781,N_12928);
nand U13971 (N_13971,N_12990,N_12865);
and U13972 (N_13972,N_12170,N_12388);
and U13973 (N_13973,N_12490,N_12750);
nand U13974 (N_13974,N_12383,N_12636);
xor U13975 (N_13975,N_12277,N_12203);
xnor U13976 (N_13976,N_12521,N_12295);
and U13977 (N_13977,N_12218,N_12637);
or U13978 (N_13978,N_12462,N_12385);
nor U13979 (N_13979,N_12843,N_12494);
or U13980 (N_13980,N_12490,N_12379);
nor U13981 (N_13981,N_12934,N_12939);
or U13982 (N_13982,N_12797,N_12628);
nand U13983 (N_13983,N_12417,N_12212);
nor U13984 (N_13984,N_12932,N_12817);
nand U13985 (N_13985,N_12008,N_12960);
nand U13986 (N_13986,N_12950,N_12539);
xor U13987 (N_13987,N_12067,N_12078);
or U13988 (N_13988,N_12064,N_12531);
nor U13989 (N_13989,N_12310,N_12290);
nand U13990 (N_13990,N_12263,N_12034);
or U13991 (N_13991,N_12675,N_12796);
nand U13992 (N_13992,N_12119,N_12563);
xnor U13993 (N_13993,N_12049,N_12062);
nor U13994 (N_13994,N_12352,N_12560);
nor U13995 (N_13995,N_12507,N_12596);
nor U13996 (N_13996,N_12195,N_12907);
xor U13997 (N_13997,N_12852,N_12341);
or U13998 (N_13998,N_12450,N_12617);
xor U13999 (N_13999,N_12210,N_12523);
and U14000 (N_14000,N_13098,N_13903);
and U14001 (N_14001,N_13097,N_13899);
and U14002 (N_14002,N_13251,N_13748);
xnor U14003 (N_14003,N_13104,N_13528);
nand U14004 (N_14004,N_13729,N_13188);
nand U14005 (N_14005,N_13516,N_13341);
nand U14006 (N_14006,N_13226,N_13541);
and U14007 (N_14007,N_13487,N_13044);
or U14008 (N_14008,N_13025,N_13122);
nor U14009 (N_14009,N_13908,N_13453);
and U14010 (N_14010,N_13915,N_13235);
or U14011 (N_14011,N_13520,N_13625);
nand U14012 (N_14012,N_13547,N_13338);
nor U14013 (N_14013,N_13950,N_13054);
or U14014 (N_14014,N_13726,N_13126);
and U14015 (N_14015,N_13739,N_13928);
xnor U14016 (N_14016,N_13172,N_13198);
xor U14017 (N_14017,N_13135,N_13527);
and U14018 (N_14018,N_13461,N_13454);
and U14019 (N_14019,N_13942,N_13807);
or U14020 (N_14020,N_13584,N_13447);
or U14021 (N_14021,N_13138,N_13163);
and U14022 (N_14022,N_13103,N_13546);
xor U14023 (N_14023,N_13946,N_13678);
xor U14024 (N_14024,N_13810,N_13558);
and U14025 (N_14025,N_13094,N_13068);
nor U14026 (N_14026,N_13857,N_13995);
xor U14027 (N_14027,N_13909,N_13140);
nor U14028 (N_14028,N_13473,N_13051);
and U14029 (N_14029,N_13313,N_13202);
nor U14030 (N_14030,N_13399,N_13674);
nor U14031 (N_14031,N_13187,N_13060);
nand U14032 (N_14032,N_13328,N_13976);
nand U14033 (N_14033,N_13016,N_13334);
or U14034 (N_14034,N_13760,N_13885);
nand U14035 (N_14035,N_13715,N_13250);
nor U14036 (N_14036,N_13593,N_13600);
nor U14037 (N_14037,N_13771,N_13291);
xor U14038 (N_14038,N_13773,N_13981);
nor U14039 (N_14039,N_13323,N_13434);
or U14040 (N_14040,N_13299,N_13204);
xnor U14041 (N_14041,N_13883,N_13196);
nand U14042 (N_14042,N_13175,N_13468);
and U14043 (N_14043,N_13040,N_13021);
nor U14044 (N_14044,N_13502,N_13431);
nor U14045 (N_14045,N_13258,N_13296);
or U14046 (N_14046,N_13999,N_13550);
or U14047 (N_14047,N_13471,N_13295);
nor U14048 (N_14048,N_13630,N_13317);
or U14049 (N_14049,N_13798,N_13038);
or U14050 (N_14050,N_13503,N_13426);
xor U14051 (N_14051,N_13752,N_13953);
and U14052 (N_14052,N_13274,N_13083);
and U14053 (N_14053,N_13462,N_13114);
and U14054 (N_14054,N_13948,N_13701);
and U14055 (N_14055,N_13116,N_13939);
xnor U14056 (N_14056,N_13457,N_13256);
xor U14057 (N_14057,N_13894,N_13694);
nor U14058 (N_14058,N_13840,N_13848);
nand U14059 (N_14059,N_13713,N_13688);
and U14060 (N_14060,N_13003,N_13601);
xor U14061 (N_14061,N_13576,N_13452);
nor U14062 (N_14062,N_13190,N_13725);
nor U14063 (N_14063,N_13746,N_13563);
and U14064 (N_14064,N_13310,N_13469);
xor U14065 (N_14065,N_13160,N_13968);
and U14066 (N_14066,N_13566,N_13232);
or U14067 (N_14067,N_13061,N_13074);
or U14068 (N_14068,N_13936,N_13489);
xnor U14069 (N_14069,N_13648,N_13684);
nor U14070 (N_14070,N_13384,N_13002);
or U14071 (N_14071,N_13552,N_13286);
nand U14072 (N_14072,N_13392,N_13095);
xor U14073 (N_14073,N_13082,N_13785);
and U14074 (N_14074,N_13270,N_13853);
or U14075 (N_14075,N_13671,N_13424);
nor U14076 (N_14076,N_13194,N_13358);
xor U14077 (N_14077,N_13540,N_13951);
nand U14078 (N_14078,N_13134,N_13505);
xor U14079 (N_14079,N_13032,N_13904);
nor U14080 (N_14080,N_13120,N_13460);
xnor U14081 (N_14081,N_13749,N_13962);
xor U14082 (N_14082,N_13761,N_13930);
nand U14083 (N_14083,N_13022,N_13917);
xnor U14084 (N_14084,N_13011,N_13151);
nand U14085 (N_14085,N_13791,N_13534);
nor U14086 (N_14086,N_13978,N_13186);
nor U14087 (N_14087,N_13716,N_13657);
or U14088 (N_14088,N_13886,N_13211);
or U14089 (N_14089,N_13742,N_13153);
nor U14090 (N_14090,N_13944,N_13170);
or U14091 (N_14091,N_13348,N_13989);
xnor U14092 (N_14092,N_13796,N_13176);
nor U14093 (N_14093,N_13632,N_13435);
nand U14094 (N_14094,N_13689,N_13660);
or U14095 (N_14095,N_13283,N_13998);
nand U14096 (N_14096,N_13219,N_13272);
or U14097 (N_14097,N_13493,N_13914);
xor U14098 (N_14098,N_13931,N_13672);
and U14099 (N_14099,N_13402,N_13562);
and U14100 (N_14100,N_13182,N_13314);
xnor U14101 (N_14101,N_13586,N_13751);
or U14102 (N_14102,N_13730,N_13259);
xor U14103 (N_14103,N_13832,N_13269);
xor U14104 (N_14104,N_13561,N_13128);
or U14105 (N_14105,N_13375,N_13071);
nor U14106 (N_14106,N_13037,N_13257);
nand U14107 (N_14107,N_13922,N_13929);
and U14108 (N_14108,N_13934,N_13843);
nand U14109 (N_14109,N_13197,N_13124);
xnor U14110 (N_14110,N_13475,N_13847);
and U14111 (N_14111,N_13906,N_13486);
xor U14112 (N_14112,N_13620,N_13644);
xor U14113 (N_14113,N_13776,N_13597);
nand U14114 (N_14114,N_13254,N_13209);
nor U14115 (N_14115,N_13548,N_13611);
or U14116 (N_14116,N_13788,N_13279);
and U14117 (N_14117,N_13902,N_13261);
and U14118 (N_14118,N_13479,N_13582);
or U14119 (N_14119,N_13873,N_13432);
xnor U14120 (N_14120,N_13136,N_13718);
xnor U14121 (N_14121,N_13991,N_13941);
nand U14122 (N_14122,N_13084,N_13531);
nand U14123 (N_14123,N_13523,N_13265);
nor U14124 (N_14124,N_13979,N_13281);
and U14125 (N_14125,N_13380,N_13680);
nand U14126 (N_14126,N_13736,N_13240);
nor U14127 (N_14127,N_13482,N_13638);
and U14128 (N_14128,N_13855,N_13234);
and U14129 (N_14129,N_13223,N_13072);
or U14130 (N_14130,N_13093,N_13280);
nor U14131 (N_14131,N_13782,N_13096);
or U14132 (N_14132,N_13542,N_13229);
nand U14133 (N_14133,N_13667,N_13307);
and U14134 (N_14134,N_13410,N_13964);
and U14135 (N_14135,N_13288,N_13860);
nand U14136 (N_14136,N_13405,N_13019);
or U14137 (N_14137,N_13926,N_13819);
nand U14138 (N_14138,N_13518,N_13697);
xnor U14139 (N_14139,N_13987,N_13125);
nand U14140 (N_14140,N_13714,N_13318);
xor U14141 (N_14141,N_13193,N_13164);
and U14142 (N_14142,N_13682,N_13608);
xor U14143 (N_14143,N_13804,N_13501);
or U14144 (N_14144,N_13612,N_13101);
xor U14145 (N_14145,N_13794,N_13438);
and U14146 (N_14146,N_13661,N_13494);
and U14147 (N_14147,N_13877,N_13195);
xor U14148 (N_14148,N_13275,N_13543);
xor U14149 (N_14149,N_13969,N_13532);
xnor U14150 (N_14150,N_13161,N_13937);
xor U14151 (N_14151,N_13433,N_13439);
and U14152 (N_14152,N_13738,N_13861);
nand U14153 (N_14153,N_13631,N_13708);
or U14154 (N_14154,N_13789,N_13409);
or U14155 (N_14155,N_13845,N_13614);
xnor U14156 (N_14156,N_13227,N_13321);
and U14157 (N_14157,N_13677,N_13339);
xnor U14158 (N_14158,N_13703,N_13519);
and U14159 (N_14159,N_13342,N_13028);
and U14160 (N_14160,N_13833,N_13893);
or U14161 (N_14161,N_13900,N_13168);
and U14162 (N_14162,N_13757,N_13535);
or U14163 (N_14163,N_13685,N_13344);
xor U14164 (N_14164,N_13663,N_13376);
or U14165 (N_14165,N_13300,N_13615);
and U14166 (N_14166,N_13112,N_13755);
xnor U14167 (N_14167,N_13719,N_13485);
nand U14168 (N_14168,N_13735,N_13076);
nor U14169 (N_14169,N_13427,N_13192);
or U14170 (N_14170,N_13598,N_13242);
nand U14171 (N_14171,N_13717,N_13997);
xnor U14172 (N_14172,N_13759,N_13133);
or U14173 (N_14173,N_13337,N_13610);
nand U14174 (N_14174,N_13653,N_13692);
and U14175 (N_14175,N_13106,N_13572);
nand U14176 (N_14176,N_13619,N_13090);
nor U14177 (N_14177,N_13092,N_13580);
nand U14178 (N_14178,N_13705,N_13013);
nand U14179 (N_14179,N_13277,N_13822);
nand U14180 (N_14180,N_13975,N_13465);
and U14181 (N_14181,N_13208,N_13818);
nor U14182 (N_14182,N_13472,N_13216);
xor U14183 (N_14183,N_13595,N_13370);
or U14184 (N_14184,N_13721,N_13784);
xor U14185 (N_14185,N_13142,N_13005);
xor U14186 (N_14186,N_13217,N_13711);
or U14187 (N_14187,N_13152,N_13617);
nor U14188 (N_14188,N_13560,N_13816);
nand U14189 (N_14189,N_13252,N_13329);
or U14190 (N_14190,N_13581,N_13876);
and U14191 (N_14191,N_13429,N_13606);
xor U14192 (N_14192,N_13925,N_13312);
xnor U14193 (N_14193,N_13393,N_13722);
nand U14194 (N_14194,N_13449,N_13728);
nor U14195 (N_14195,N_13360,N_13799);
nor U14196 (N_14196,N_13316,N_13311);
nand U14197 (N_14197,N_13564,N_13345);
nand U14198 (N_14198,N_13043,N_13629);
xor U14199 (N_14199,N_13417,N_13635);
nand U14200 (N_14200,N_13215,N_13118);
xnor U14201 (N_14201,N_13779,N_13642);
xor U14202 (N_14202,N_13699,N_13511);
and U14203 (N_14203,N_13377,N_13102);
and U14204 (N_14204,N_13408,N_13298);
and U14205 (N_14205,N_13495,N_13734);
and U14206 (N_14206,N_13368,N_13545);
nor U14207 (N_14207,N_13292,N_13374);
and U14208 (N_14208,N_13686,N_13228);
and U14209 (N_14209,N_13897,N_13165);
or U14210 (N_14210,N_13079,N_13144);
nand U14211 (N_14211,N_13813,N_13693);
or U14212 (N_14212,N_13765,N_13797);
nand U14213 (N_14213,N_13591,N_13347);
xnor U14214 (N_14214,N_13207,N_13415);
nor U14215 (N_14215,N_13354,N_13145);
xnor U14216 (N_14216,N_13920,N_13696);
nand U14217 (N_14217,N_13826,N_13573);
and U14218 (N_14218,N_13089,N_13023);
nand U14219 (N_14219,N_13756,N_13325);
or U14220 (N_14220,N_13828,N_13067);
nand U14221 (N_14221,N_13080,N_13436);
and U14222 (N_14222,N_13363,N_13880);
and U14223 (N_14223,N_13842,N_13982);
nand U14224 (N_14224,N_13983,N_13960);
or U14225 (N_14225,N_13895,N_13958);
nor U14226 (N_14226,N_13220,N_13400);
nor U14227 (N_14227,N_13233,N_13515);
or U14228 (N_14228,N_13753,N_13859);
nor U14229 (N_14229,N_13727,N_13086);
nand U14230 (N_14230,N_13935,N_13639);
and U14231 (N_14231,N_13988,N_13009);
nand U14232 (N_14232,N_13646,N_13050);
or U14233 (N_14233,N_13008,N_13437);
and U14234 (N_14234,N_13015,N_13108);
and U14235 (N_14235,N_13687,N_13959);
nor U14236 (N_14236,N_13679,N_13733);
and U14237 (N_14237,N_13825,N_13309);
or U14238 (N_14238,N_13070,N_13210);
xnor U14239 (N_14239,N_13767,N_13156);
xnor U14240 (N_14240,N_13866,N_13780);
nor U14241 (N_14241,N_13655,N_13557);
and U14242 (N_14242,N_13398,N_13879);
and U14243 (N_14243,N_13792,N_13000);
or U14244 (N_14244,N_13297,N_13319);
nand U14245 (N_14245,N_13910,N_13884);
nor U14246 (N_14246,N_13121,N_13647);
nor U14247 (N_14247,N_13504,N_13356);
or U14248 (N_14248,N_13383,N_13184);
nand U14249 (N_14249,N_13744,N_13030);
nor U14250 (N_14250,N_13724,N_13521);
nor U14251 (N_14251,N_13622,N_13173);
and U14252 (N_14252,N_13916,N_13575);
or U14253 (N_14253,N_13676,N_13419);
nand U14254 (N_14254,N_13602,N_13373);
nand U14255 (N_14255,N_13039,N_13115);
xnor U14256 (N_14256,N_13260,N_13059);
nand U14257 (N_14257,N_13111,N_13484);
and U14258 (N_14258,N_13150,N_13568);
nor U14259 (N_14259,N_13241,N_13322);
nor U14260 (N_14260,N_13474,N_13222);
xor U14261 (N_14261,N_13177,N_13993);
or U14262 (N_14262,N_13887,N_13649);
and U14263 (N_14263,N_13651,N_13673);
nand U14264 (N_14264,N_13556,N_13938);
or U14265 (N_14265,N_13965,N_13616);
or U14266 (N_14266,N_13183,N_13056);
xnor U14267 (N_14267,N_13821,N_13483);
and U14268 (N_14268,N_13132,N_13466);
xnor U14269 (N_14269,N_13440,N_13180);
xnor U14270 (N_14270,N_13191,N_13411);
nor U14271 (N_14271,N_13470,N_13255);
or U14272 (N_14272,N_13167,N_13918);
xor U14273 (N_14273,N_13031,N_13872);
nor U14274 (N_14274,N_13605,N_13587);
xnor U14275 (N_14275,N_13123,N_13852);
and U14276 (N_14276,N_13130,N_13795);
xor U14277 (N_14277,N_13571,N_13057);
and U14278 (N_14278,N_13006,N_13603);
nor U14279 (N_14279,N_13413,N_13069);
nor U14280 (N_14280,N_13555,N_13882);
xor U14281 (N_14281,N_13662,N_13065);
and U14282 (N_14282,N_13446,N_13851);
or U14283 (N_14283,N_13805,N_13850);
xnor U14284 (N_14284,N_13559,N_13034);
and U14285 (N_14285,N_13898,N_13954);
or U14286 (N_14286,N_13787,N_13737);
nor U14287 (N_14287,N_13707,N_13837);
or U14288 (N_14288,N_13428,N_13357);
or U14289 (N_14289,N_13583,N_13509);
nor U14290 (N_14290,N_13589,N_13327);
and U14291 (N_14291,N_13670,N_13731);
xor U14292 (N_14292,N_13977,N_13814);
or U14293 (N_14293,N_13927,N_13248);
nand U14294 (N_14294,N_13522,N_13533);
nand U14295 (N_14295,N_13924,N_13970);
xnor U14296 (N_14296,N_13838,N_13513);
nor U14297 (N_14297,N_13154,N_13014);
and U14298 (N_14298,N_13225,N_13001);
or U14299 (N_14299,N_13129,N_13336);
or U14300 (N_14300,N_13350,N_13875);
or U14301 (N_14301,N_13458,N_13035);
nor U14302 (N_14302,N_13754,N_13407);
xor U14303 (N_14303,N_13803,N_13247);
and U14304 (N_14304,N_13359,N_13169);
or U14305 (N_14305,N_13430,N_13723);
or U14306 (N_14306,N_13675,N_13010);
nor U14307 (N_14307,N_13397,N_13517);
nand U14308 (N_14308,N_13656,N_13956);
and U14309 (N_14309,N_13236,N_13117);
and U14310 (N_14310,N_13913,N_13775);
nor U14311 (N_14311,N_13088,N_13075);
xnor U14312 (N_14312,N_13127,N_13854);
and U14313 (N_14313,N_13514,N_13783);
or U14314 (N_14314,N_13282,N_13634);
or U14315 (N_14315,N_13416,N_13626);
xnor U14316 (N_14316,N_13985,N_13865);
nor U14317 (N_14317,N_13574,N_13823);
and U14318 (N_14318,N_13500,N_13862);
nand U14319 (N_14319,N_13864,N_13890);
or U14320 (N_14320,N_13268,N_13324);
nand U14321 (N_14321,N_13806,N_13218);
or U14322 (N_14322,N_13996,N_13055);
xnor U14323 (N_14323,N_13740,N_13790);
nor U14324 (N_14324,N_13786,N_13802);
nor U14325 (N_14325,N_13621,N_13698);
xor U14326 (N_14326,N_13955,N_13294);
and U14327 (N_14327,N_13947,N_13800);
or U14328 (N_14328,N_13905,N_13669);
or U14329 (N_14329,N_13063,N_13366);
xnor U14330 (N_14330,N_13231,N_13459);
nor U14331 (N_14331,N_13867,N_13654);
nor U14332 (N_14332,N_13308,N_13476);
nand U14333 (N_14333,N_13637,N_13801);
xnor U14334 (N_14334,N_13107,N_13645);
and U14335 (N_14335,N_13881,N_13706);
nor U14336 (N_14336,N_13162,N_13414);
or U14337 (N_14337,N_13214,N_13200);
nand U14338 (N_14338,N_13418,N_13372);
nand U14339 (N_14339,N_13577,N_13596);
and U14340 (N_14340,N_13491,N_13896);
nand U14341 (N_14341,N_13369,N_13640);
or U14342 (N_14342,N_13143,N_13387);
nor U14343 (N_14343,N_13390,N_13808);
nor U14344 (N_14344,N_13599,N_13388);
and U14345 (N_14345,N_13224,N_13641);
xor U14346 (N_14346,N_13974,N_13213);
or U14347 (N_14347,N_13244,N_13036);
xor U14348 (N_14348,N_13665,N_13333);
nand U14349 (N_14349,N_13488,N_13538);
and U14350 (N_14350,N_13249,N_13178);
or U14351 (N_14351,N_13253,N_13421);
xnor U14352 (N_14352,N_13045,N_13874);
nand U14353 (N_14353,N_13058,N_13841);
or U14354 (N_14354,N_13441,N_13443);
nand U14355 (N_14355,N_13769,N_13844);
nor U14356 (N_14356,N_13967,N_13159);
nor U14357 (N_14357,N_13704,N_13066);
xor U14358 (N_14358,N_13588,N_13870);
or U14359 (N_14359,N_13994,N_13199);
nand U14360 (N_14360,N_13046,N_13778);
and U14361 (N_14361,N_13404,N_13456);
and U14362 (N_14362,N_13181,N_13592);
nand U14363 (N_14363,N_13078,N_13772);
nor U14364 (N_14364,N_13131,N_13012);
nor U14365 (N_14365,N_13238,N_13442);
or U14366 (N_14366,N_13110,N_13529);
xor U14367 (N_14367,N_13444,N_13892);
and U14368 (N_14368,N_13467,N_13349);
and U14369 (N_14369,N_13966,N_13174);
nand U14370 (N_14370,N_13099,N_13451);
or U14371 (N_14371,N_13971,N_13266);
xnor U14372 (N_14372,N_13980,N_13029);
xor U14373 (N_14373,N_13026,N_13607);
xnor U14374 (N_14374,N_13246,N_13712);
or U14375 (N_14375,N_13406,N_13945);
and U14376 (N_14376,N_13817,N_13047);
or U14377 (N_14377,N_13304,N_13835);
nor U14378 (N_14378,N_13284,N_13766);
and U14379 (N_14379,N_13664,N_13113);
xnor U14380 (N_14380,N_13839,N_13189);
or U14381 (N_14381,N_13027,N_13303);
nor U14382 (N_14382,N_13510,N_13412);
xnor U14383 (N_14383,N_13381,N_13496);
and U14384 (N_14384,N_13774,N_13379);
and U14385 (N_14385,N_13353,N_13149);
nor U14386 (N_14386,N_13957,N_13481);
or U14387 (N_14387,N_13691,N_13508);
nor U14388 (N_14388,N_13100,N_13477);
and U14389 (N_14389,N_13048,N_13633);
nor U14390 (N_14390,N_13394,N_13933);
xnor U14391 (N_14391,N_13391,N_13171);
nor U14392 (N_14392,N_13148,N_13385);
or U14393 (N_14393,N_13267,N_13973);
or U14394 (N_14394,N_13263,N_13963);
xnor U14395 (N_14395,N_13365,N_13590);
xnor U14396 (N_14396,N_13332,N_13554);
and U14397 (N_14397,N_13949,N_13681);
or U14398 (N_14398,N_13695,N_13203);
or U14399 (N_14399,N_13340,N_13371);
or U14400 (N_14400,N_13109,N_13290);
xor U14401 (N_14401,N_13758,N_13659);
nand U14402 (N_14402,N_13346,N_13450);
nand U14403 (N_14403,N_13330,N_13326);
xnor U14404 (N_14404,N_13585,N_13888);
or U14405 (N_14405,N_13793,N_13306);
xor U14406 (N_14406,N_13553,N_13352);
xor U14407 (N_14407,N_13445,N_13081);
nor U14408 (N_14408,N_13343,N_13565);
xor U14409 (N_14409,N_13666,N_13750);
or U14410 (N_14410,N_13829,N_13932);
xnor U14411 (N_14411,N_13157,N_13273);
nor U14412 (N_14412,N_13085,N_13239);
and U14413 (N_14413,N_13463,N_13869);
xnor U14414 (N_14414,N_13480,N_13062);
xnor U14415 (N_14415,N_13033,N_13020);
nand U14416 (N_14416,N_13745,N_13395);
nand U14417 (N_14417,N_13004,N_13389);
or U14418 (N_14418,N_13741,N_13525);
or U14419 (N_14419,N_13425,N_13650);
nor U14420 (N_14420,N_13492,N_13849);
xnor U14421 (N_14421,N_13567,N_13331);
nor U14422 (N_14422,N_13064,N_13907);
or U14423 (N_14423,N_13700,N_13315);
xnor U14424 (N_14424,N_13105,N_13185);
xnor U14425 (N_14425,N_13053,N_13815);
nand U14426 (N_14426,N_13831,N_13830);
or U14427 (N_14427,N_13961,N_13539);
xor U14428 (N_14428,N_13579,N_13448);
or U14429 (N_14429,N_13747,N_13042);
nand U14430 (N_14430,N_13278,N_13628);
nand U14431 (N_14431,N_13382,N_13570);
and U14432 (N_14432,N_13361,N_13041);
xnor U14433 (N_14433,N_13986,N_13179);
nand U14434 (N_14434,N_13243,N_13024);
xnor U14435 (N_14435,N_13627,N_13091);
nor U14436 (N_14436,N_13396,N_13720);
and U14437 (N_14437,N_13710,N_13658);
xor U14438 (N_14438,N_13139,N_13386);
and U14439 (N_14439,N_13604,N_13507);
xor U14440 (N_14440,N_13732,N_13537);
or U14441 (N_14441,N_13891,N_13351);
and U14442 (N_14442,N_13536,N_13245);
xor U14443 (N_14443,N_13919,N_13668);
nor U14444 (N_14444,N_13205,N_13578);
nor U14445 (N_14445,N_13293,N_13868);
and U14446 (N_14446,N_13320,N_13155);
xnor U14447 (N_14447,N_13403,N_13301);
nor U14448 (N_14448,N_13871,N_13305);
xor U14449 (N_14449,N_13827,N_13878);
nor U14450 (N_14450,N_13287,N_13940);
and U14451 (N_14451,N_13624,N_13478);
nand U14452 (N_14452,N_13856,N_13137);
and U14453 (N_14453,N_13623,N_13636);
or U14454 (N_14454,N_13990,N_13709);
and U14455 (N_14455,N_13569,N_13166);
nand U14456 (N_14456,N_13992,N_13367);
nor U14457 (N_14457,N_13212,N_13362);
xnor U14458 (N_14458,N_13355,N_13943);
and U14459 (N_14459,N_13764,N_13643);
or U14460 (N_14460,N_13812,N_13912);
xor U14461 (N_14461,N_13762,N_13498);
or U14462 (N_14462,N_13276,N_13763);
or U14463 (N_14463,N_13146,N_13007);
and U14464 (N_14464,N_13618,N_13952);
nand U14465 (N_14465,N_13455,N_13770);
nand U14466 (N_14466,N_13499,N_13530);
xor U14467 (N_14467,N_13834,N_13690);
xnor U14468 (N_14468,N_13018,N_13289);
nor U14469 (N_14469,N_13049,N_13364);
and U14470 (N_14470,N_13230,N_13464);
or U14471 (N_14471,N_13158,N_13262);
or U14472 (N_14472,N_13423,N_13087);
nor U14473 (N_14473,N_13077,N_13846);
nor U14474 (N_14474,N_13777,N_13921);
xnor U14475 (N_14475,N_13524,N_13335);
xnor U14476 (N_14476,N_13613,N_13141);
nor U14477 (N_14477,N_13512,N_13652);
or U14478 (N_14478,N_13052,N_13863);
and U14479 (N_14479,N_13683,N_13147);
xor U14480 (N_14480,N_13206,N_13811);
and U14481 (N_14481,N_13702,N_13221);
or U14482 (N_14482,N_13594,N_13984);
xor U14483 (N_14483,N_13858,N_13271);
nand U14484 (N_14484,N_13544,N_13285);
and U14485 (N_14485,N_13809,N_13073);
and U14486 (N_14486,N_13506,N_13923);
or U14487 (N_14487,N_13422,N_13824);
xor U14488 (N_14488,N_13526,N_13889);
nand U14489 (N_14489,N_13237,N_13119);
or U14490 (N_14490,N_13972,N_13017);
nor U14491 (N_14491,N_13911,N_13201);
or U14492 (N_14492,N_13901,N_13378);
or U14493 (N_14493,N_13836,N_13609);
xnor U14494 (N_14494,N_13401,N_13551);
nor U14495 (N_14495,N_13820,N_13781);
and U14496 (N_14496,N_13490,N_13768);
nand U14497 (N_14497,N_13302,N_13497);
or U14498 (N_14498,N_13420,N_13264);
xor U14499 (N_14499,N_13743,N_13549);
and U14500 (N_14500,N_13872,N_13099);
nor U14501 (N_14501,N_13086,N_13959);
xnor U14502 (N_14502,N_13517,N_13753);
nand U14503 (N_14503,N_13052,N_13227);
or U14504 (N_14504,N_13422,N_13076);
xor U14505 (N_14505,N_13441,N_13224);
xor U14506 (N_14506,N_13340,N_13039);
xor U14507 (N_14507,N_13456,N_13664);
nand U14508 (N_14508,N_13103,N_13918);
and U14509 (N_14509,N_13434,N_13965);
or U14510 (N_14510,N_13735,N_13827);
xor U14511 (N_14511,N_13582,N_13170);
nand U14512 (N_14512,N_13958,N_13777);
or U14513 (N_14513,N_13935,N_13670);
and U14514 (N_14514,N_13388,N_13073);
nand U14515 (N_14515,N_13322,N_13158);
and U14516 (N_14516,N_13516,N_13679);
nand U14517 (N_14517,N_13036,N_13661);
or U14518 (N_14518,N_13422,N_13899);
or U14519 (N_14519,N_13835,N_13662);
or U14520 (N_14520,N_13211,N_13970);
nor U14521 (N_14521,N_13004,N_13039);
nor U14522 (N_14522,N_13167,N_13973);
nand U14523 (N_14523,N_13023,N_13704);
nor U14524 (N_14524,N_13708,N_13935);
and U14525 (N_14525,N_13529,N_13810);
xor U14526 (N_14526,N_13176,N_13184);
xor U14527 (N_14527,N_13839,N_13498);
and U14528 (N_14528,N_13778,N_13760);
xor U14529 (N_14529,N_13748,N_13643);
or U14530 (N_14530,N_13711,N_13943);
xnor U14531 (N_14531,N_13132,N_13701);
and U14532 (N_14532,N_13208,N_13514);
nand U14533 (N_14533,N_13959,N_13725);
or U14534 (N_14534,N_13698,N_13135);
nor U14535 (N_14535,N_13692,N_13897);
nor U14536 (N_14536,N_13837,N_13186);
nand U14537 (N_14537,N_13527,N_13355);
xor U14538 (N_14538,N_13517,N_13817);
and U14539 (N_14539,N_13085,N_13836);
nor U14540 (N_14540,N_13468,N_13500);
nor U14541 (N_14541,N_13165,N_13550);
nor U14542 (N_14542,N_13394,N_13254);
xnor U14543 (N_14543,N_13582,N_13790);
or U14544 (N_14544,N_13038,N_13241);
or U14545 (N_14545,N_13346,N_13894);
and U14546 (N_14546,N_13385,N_13608);
xnor U14547 (N_14547,N_13586,N_13418);
nand U14548 (N_14548,N_13479,N_13938);
or U14549 (N_14549,N_13665,N_13324);
or U14550 (N_14550,N_13494,N_13350);
and U14551 (N_14551,N_13315,N_13961);
and U14552 (N_14552,N_13245,N_13153);
nand U14553 (N_14553,N_13885,N_13282);
or U14554 (N_14554,N_13890,N_13790);
nand U14555 (N_14555,N_13672,N_13940);
or U14556 (N_14556,N_13752,N_13260);
nand U14557 (N_14557,N_13554,N_13097);
xnor U14558 (N_14558,N_13673,N_13638);
nand U14559 (N_14559,N_13051,N_13244);
and U14560 (N_14560,N_13997,N_13160);
or U14561 (N_14561,N_13418,N_13434);
nand U14562 (N_14562,N_13029,N_13075);
nand U14563 (N_14563,N_13590,N_13914);
and U14564 (N_14564,N_13590,N_13184);
and U14565 (N_14565,N_13587,N_13782);
xor U14566 (N_14566,N_13337,N_13525);
xnor U14567 (N_14567,N_13570,N_13429);
nor U14568 (N_14568,N_13229,N_13901);
nor U14569 (N_14569,N_13861,N_13412);
or U14570 (N_14570,N_13926,N_13253);
nand U14571 (N_14571,N_13147,N_13059);
xor U14572 (N_14572,N_13466,N_13263);
nor U14573 (N_14573,N_13443,N_13462);
nand U14574 (N_14574,N_13407,N_13387);
and U14575 (N_14575,N_13600,N_13842);
nor U14576 (N_14576,N_13385,N_13273);
xor U14577 (N_14577,N_13286,N_13037);
or U14578 (N_14578,N_13173,N_13884);
and U14579 (N_14579,N_13587,N_13861);
nor U14580 (N_14580,N_13747,N_13028);
or U14581 (N_14581,N_13263,N_13881);
nand U14582 (N_14582,N_13172,N_13199);
nor U14583 (N_14583,N_13782,N_13972);
or U14584 (N_14584,N_13721,N_13255);
nor U14585 (N_14585,N_13170,N_13077);
xnor U14586 (N_14586,N_13286,N_13401);
or U14587 (N_14587,N_13121,N_13742);
nor U14588 (N_14588,N_13301,N_13615);
or U14589 (N_14589,N_13186,N_13249);
nor U14590 (N_14590,N_13231,N_13934);
nand U14591 (N_14591,N_13539,N_13020);
and U14592 (N_14592,N_13389,N_13756);
and U14593 (N_14593,N_13617,N_13419);
xor U14594 (N_14594,N_13769,N_13899);
xnor U14595 (N_14595,N_13229,N_13046);
nand U14596 (N_14596,N_13767,N_13390);
nand U14597 (N_14597,N_13520,N_13539);
xor U14598 (N_14598,N_13358,N_13040);
nand U14599 (N_14599,N_13376,N_13685);
nor U14600 (N_14600,N_13118,N_13388);
nand U14601 (N_14601,N_13805,N_13818);
and U14602 (N_14602,N_13783,N_13386);
nand U14603 (N_14603,N_13812,N_13412);
nor U14604 (N_14604,N_13645,N_13451);
xor U14605 (N_14605,N_13750,N_13724);
nand U14606 (N_14606,N_13033,N_13276);
nor U14607 (N_14607,N_13741,N_13147);
and U14608 (N_14608,N_13292,N_13065);
and U14609 (N_14609,N_13288,N_13117);
xnor U14610 (N_14610,N_13895,N_13703);
and U14611 (N_14611,N_13754,N_13460);
or U14612 (N_14612,N_13865,N_13732);
and U14613 (N_14613,N_13108,N_13503);
and U14614 (N_14614,N_13429,N_13684);
and U14615 (N_14615,N_13628,N_13143);
and U14616 (N_14616,N_13193,N_13656);
nor U14617 (N_14617,N_13301,N_13446);
nand U14618 (N_14618,N_13719,N_13402);
xor U14619 (N_14619,N_13105,N_13004);
or U14620 (N_14620,N_13909,N_13933);
xnor U14621 (N_14621,N_13445,N_13488);
or U14622 (N_14622,N_13247,N_13412);
and U14623 (N_14623,N_13156,N_13090);
and U14624 (N_14624,N_13548,N_13087);
xor U14625 (N_14625,N_13687,N_13420);
or U14626 (N_14626,N_13820,N_13756);
and U14627 (N_14627,N_13331,N_13498);
nand U14628 (N_14628,N_13816,N_13244);
and U14629 (N_14629,N_13593,N_13614);
or U14630 (N_14630,N_13449,N_13512);
or U14631 (N_14631,N_13206,N_13285);
nand U14632 (N_14632,N_13913,N_13791);
or U14633 (N_14633,N_13987,N_13046);
nor U14634 (N_14634,N_13601,N_13742);
nor U14635 (N_14635,N_13647,N_13346);
or U14636 (N_14636,N_13477,N_13988);
nand U14637 (N_14637,N_13836,N_13029);
nor U14638 (N_14638,N_13948,N_13831);
nand U14639 (N_14639,N_13320,N_13090);
and U14640 (N_14640,N_13296,N_13292);
nor U14641 (N_14641,N_13480,N_13459);
nand U14642 (N_14642,N_13372,N_13286);
xnor U14643 (N_14643,N_13248,N_13098);
xnor U14644 (N_14644,N_13259,N_13856);
nand U14645 (N_14645,N_13193,N_13397);
or U14646 (N_14646,N_13462,N_13414);
and U14647 (N_14647,N_13734,N_13921);
and U14648 (N_14648,N_13260,N_13868);
nand U14649 (N_14649,N_13596,N_13884);
xor U14650 (N_14650,N_13830,N_13700);
xor U14651 (N_14651,N_13817,N_13337);
nand U14652 (N_14652,N_13636,N_13774);
nand U14653 (N_14653,N_13463,N_13046);
and U14654 (N_14654,N_13147,N_13485);
nand U14655 (N_14655,N_13208,N_13022);
or U14656 (N_14656,N_13142,N_13267);
xor U14657 (N_14657,N_13033,N_13957);
or U14658 (N_14658,N_13592,N_13890);
nor U14659 (N_14659,N_13867,N_13799);
and U14660 (N_14660,N_13014,N_13117);
and U14661 (N_14661,N_13268,N_13704);
nor U14662 (N_14662,N_13445,N_13052);
and U14663 (N_14663,N_13674,N_13227);
and U14664 (N_14664,N_13447,N_13631);
nor U14665 (N_14665,N_13817,N_13417);
and U14666 (N_14666,N_13447,N_13304);
nand U14667 (N_14667,N_13863,N_13984);
nand U14668 (N_14668,N_13748,N_13220);
or U14669 (N_14669,N_13738,N_13406);
nand U14670 (N_14670,N_13432,N_13330);
nand U14671 (N_14671,N_13497,N_13618);
xnor U14672 (N_14672,N_13678,N_13176);
and U14673 (N_14673,N_13414,N_13952);
or U14674 (N_14674,N_13734,N_13081);
or U14675 (N_14675,N_13021,N_13508);
or U14676 (N_14676,N_13999,N_13823);
nor U14677 (N_14677,N_13680,N_13873);
xor U14678 (N_14678,N_13267,N_13187);
nor U14679 (N_14679,N_13955,N_13401);
xnor U14680 (N_14680,N_13143,N_13822);
and U14681 (N_14681,N_13202,N_13031);
nand U14682 (N_14682,N_13135,N_13045);
nor U14683 (N_14683,N_13463,N_13674);
and U14684 (N_14684,N_13257,N_13350);
nor U14685 (N_14685,N_13656,N_13604);
or U14686 (N_14686,N_13443,N_13942);
xor U14687 (N_14687,N_13234,N_13500);
nand U14688 (N_14688,N_13489,N_13231);
or U14689 (N_14689,N_13584,N_13849);
or U14690 (N_14690,N_13235,N_13674);
and U14691 (N_14691,N_13307,N_13149);
nand U14692 (N_14692,N_13049,N_13538);
and U14693 (N_14693,N_13633,N_13152);
nand U14694 (N_14694,N_13639,N_13702);
and U14695 (N_14695,N_13920,N_13321);
and U14696 (N_14696,N_13740,N_13632);
nor U14697 (N_14697,N_13330,N_13570);
xor U14698 (N_14698,N_13477,N_13505);
and U14699 (N_14699,N_13867,N_13001);
nand U14700 (N_14700,N_13496,N_13445);
or U14701 (N_14701,N_13364,N_13269);
nor U14702 (N_14702,N_13377,N_13957);
or U14703 (N_14703,N_13211,N_13410);
xnor U14704 (N_14704,N_13342,N_13672);
nand U14705 (N_14705,N_13109,N_13198);
and U14706 (N_14706,N_13473,N_13863);
or U14707 (N_14707,N_13086,N_13837);
or U14708 (N_14708,N_13162,N_13508);
nand U14709 (N_14709,N_13329,N_13135);
xor U14710 (N_14710,N_13748,N_13908);
nand U14711 (N_14711,N_13380,N_13054);
xnor U14712 (N_14712,N_13711,N_13506);
nor U14713 (N_14713,N_13430,N_13182);
or U14714 (N_14714,N_13651,N_13878);
or U14715 (N_14715,N_13028,N_13502);
nor U14716 (N_14716,N_13664,N_13815);
nand U14717 (N_14717,N_13370,N_13207);
nor U14718 (N_14718,N_13276,N_13456);
or U14719 (N_14719,N_13055,N_13168);
or U14720 (N_14720,N_13096,N_13277);
nor U14721 (N_14721,N_13713,N_13075);
nor U14722 (N_14722,N_13439,N_13342);
nor U14723 (N_14723,N_13197,N_13960);
nor U14724 (N_14724,N_13144,N_13339);
and U14725 (N_14725,N_13637,N_13143);
or U14726 (N_14726,N_13014,N_13360);
nand U14727 (N_14727,N_13407,N_13147);
xor U14728 (N_14728,N_13410,N_13068);
nor U14729 (N_14729,N_13311,N_13127);
nor U14730 (N_14730,N_13016,N_13080);
xnor U14731 (N_14731,N_13440,N_13474);
and U14732 (N_14732,N_13282,N_13417);
nand U14733 (N_14733,N_13998,N_13343);
xnor U14734 (N_14734,N_13849,N_13644);
or U14735 (N_14735,N_13024,N_13458);
or U14736 (N_14736,N_13153,N_13715);
nand U14737 (N_14737,N_13798,N_13713);
and U14738 (N_14738,N_13898,N_13977);
nand U14739 (N_14739,N_13042,N_13124);
xnor U14740 (N_14740,N_13708,N_13936);
nor U14741 (N_14741,N_13322,N_13732);
and U14742 (N_14742,N_13561,N_13442);
nor U14743 (N_14743,N_13157,N_13008);
and U14744 (N_14744,N_13291,N_13511);
xor U14745 (N_14745,N_13030,N_13753);
or U14746 (N_14746,N_13041,N_13777);
nor U14747 (N_14747,N_13852,N_13976);
xnor U14748 (N_14748,N_13343,N_13726);
nand U14749 (N_14749,N_13997,N_13209);
nand U14750 (N_14750,N_13852,N_13951);
nor U14751 (N_14751,N_13830,N_13750);
nand U14752 (N_14752,N_13305,N_13490);
and U14753 (N_14753,N_13276,N_13772);
nand U14754 (N_14754,N_13540,N_13195);
nor U14755 (N_14755,N_13635,N_13108);
nand U14756 (N_14756,N_13165,N_13126);
nor U14757 (N_14757,N_13007,N_13060);
or U14758 (N_14758,N_13592,N_13975);
nand U14759 (N_14759,N_13896,N_13336);
xnor U14760 (N_14760,N_13635,N_13222);
nor U14761 (N_14761,N_13608,N_13898);
or U14762 (N_14762,N_13064,N_13416);
xnor U14763 (N_14763,N_13621,N_13762);
xor U14764 (N_14764,N_13334,N_13146);
or U14765 (N_14765,N_13508,N_13861);
and U14766 (N_14766,N_13504,N_13682);
and U14767 (N_14767,N_13220,N_13559);
or U14768 (N_14768,N_13994,N_13741);
and U14769 (N_14769,N_13587,N_13678);
nand U14770 (N_14770,N_13367,N_13832);
and U14771 (N_14771,N_13488,N_13394);
nand U14772 (N_14772,N_13566,N_13373);
nand U14773 (N_14773,N_13208,N_13792);
nand U14774 (N_14774,N_13018,N_13610);
xnor U14775 (N_14775,N_13495,N_13435);
and U14776 (N_14776,N_13610,N_13232);
and U14777 (N_14777,N_13906,N_13749);
and U14778 (N_14778,N_13644,N_13750);
nor U14779 (N_14779,N_13580,N_13194);
and U14780 (N_14780,N_13409,N_13884);
or U14781 (N_14781,N_13444,N_13094);
nor U14782 (N_14782,N_13681,N_13749);
xor U14783 (N_14783,N_13537,N_13850);
nor U14784 (N_14784,N_13146,N_13679);
or U14785 (N_14785,N_13799,N_13062);
and U14786 (N_14786,N_13309,N_13733);
or U14787 (N_14787,N_13203,N_13902);
and U14788 (N_14788,N_13039,N_13088);
and U14789 (N_14789,N_13936,N_13540);
xor U14790 (N_14790,N_13119,N_13317);
and U14791 (N_14791,N_13159,N_13262);
or U14792 (N_14792,N_13787,N_13974);
or U14793 (N_14793,N_13983,N_13475);
nor U14794 (N_14794,N_13070,N_13677);
or U14795 (N_14795,N_13013,N_13408);
and U14796 (N_14796,N_13375,N_13470);
and U14797 (N_14797,N_13437,N_13915);
and U14798 (N_14798,N_13166,N_13787);
nor U14799 (N_14799,N_13846,N_13651);
and U14800 (N_14800,N_13996,N_13821);
nand U14801 (N_14801,N_13522,N_13134);
and U14802 (N_14802,N_13517,N_13220);
and U14803 (N_14803,N_13734,N_13828);
and U14804 (N_14804,N_13409,N_13781);
and U14805 (N_14805,N_13944,N_13295);
and U14806 (N_14806,N_13139,N_13062);
nand U14807 (N_14807,N_13807,N_13494);
nor U14808 (N_14808,N_13752,N_13748);
or U14809 (N_14809,N_13406,N_13817);
nor U14810 (N_14810,N_13665,N_13006);
xor U14811 (N_14811,N_13206,N_13850);
xnor U14812 (N_14812,N_13222,N_13931);
xor U14813 (N_14813,N_13554,N_13984);
or U14814 (N_14814,N_13369,N_13311);
or U14815 (N_14815,N_13405,N_13408);
and U14816 (N_14816,N_13666,N_13035);
and U14817 (N_14817,N_13372,N_13157);
nand U14818 (N_14818,N_13720,N_13637);
nor U14819 (N_14819,N_13509,N_13575);
and U14820 (N_14820,N_13738,N_13389);
xor U14821 (N_14821,N_13082,N_13366);
nand U14822 (N_14822,N_13071,N_13758);
xnor U14823 (N_14823,N_13591,N_13377);
xnor U14824 (N_14824,N_13946,N_13553);
and U14825 (N_14825,N_13492,N_13421);
nor U14826 (N_14826,N_13908,N_13505);
xnor U14827 (N_14827,N_13339,N_13717);
and U14828 (N_14828,N_13490,N_13268);
nor U14829 (N_14829,N_13176,N_13626);
nand U14830 (N_14830,N_13211,N_13560);
nand U14831 (N_14831,N_13986,N_13380);
xor U14832 (N_14832,N_13434,N_13343);
nor U14833 (N_14833,N_13622,N_13692);
nand U14834 (N_14834,N_13176,N_13078);
or U14835 (N_14835,N_13153,N_13336);
or U14836 (N_14836,N_13040,N_13693);
nor U14837 (N_14837,N_13835,N_13588);
nor U14838 (N_14838,N_13998,N_13048);
xnor U14839 (N_14839,N_13907,N_13258);
nor U14840 (N_14840,N_13957,N_13553);
nand U14841 (N_14841,N_13568,N_13535);
nor U14842 (N_14842,N_13299,N_13134);
and U14843 (N_14843,N_13994,N_13109);
or U14844 (N_14844,N_13018,N_13470);
xor U14845 (N_14845,N_13368,N_13229);
xor U14846 (N_14846,N_13258,N_13007);
xor U14847 (N_14847,N_13015,N_13310);
and U14848 (N_14848,N_13799,N_13778);
xor U14849 (N_14849,N_13174,N_13150);
nand U14850 (N_14850,N_13210,N_13152);
nor U14851 (N_14851,N_13953,N_13588);
nand U14852 (N_14852,N_13364,N_13133);
nor U14853 (N_14853,N_13724,N_13310);
or U14854 (N_14854,N_13751,N_13870);
or U14855 (N_14855,N_13418,N_13968);
nand U14856 (N_14856,N_13058,N_13303);
xor U14857 (N_14857,N_13997,N_13332);
nor U14858 (N_14858,N_13854,N_13125);
xor U14859 (N_14859,N_13437,N_13390);
nor U14860 (N_14860,N_13662,N_13092);
nor U14861 (N_14861,N_13926,N_13237);
nor U14862 (N_14862,N_13098,N_13867);
nor U14863 (N_14863,N_13504,N_13083);
nor U14864 (N_14864,N_13965,N_13139);
nor U14865 (N_14865,N_13051,N_13518);
nor U14866 (N_14866,N_13585,N_13414);
or U14867 (N_14867,N_13463,N_13280);
and U14868 (N_14868,N_13227,N_13890);
nand U14869 (N_14869,N_13164,N_13493);
nand U14870 (N_14870,N_13337,N_13485);
xor U14871 (N_14871,N_13658,N_13513);
xnor U14872 (N_14872,N_13147,N_13320);
or U14873 (N_14873,N_13693,N_13271);
and U14874 (N_14874,N_13818,N_13038);
and U14875 (N_14875,N_13971,N_13888);
or U14876 (N_14876,N_13989,N_13688);
nand U14877 (N_14877,N_13684,N_13511);
nand U14878 (N_14878,N_13693,N_13225);
nand U14879 (N_14879,N_13017,N_13016);
nand U14880 (N_14880,N_13982,N_13204);
xnor U14881 (N_14881,N_13436,N_13553);
and U14882 (N_14882,N_13997,N_13283);
or U14883 (N_14883,N_13796,N_13531);
or U14884 (N_14884,N_13544,N_13907);
or U14885 (N_14885,N_13144,N_13053);
xor U14886 (N_14886,N_13942,N_13549);
nor U14887 (N_14887,N_13337,N_13805);
nor U14888 (N_14888,N_13541,N_13523);
nand U14889 (N_14889,N_13957,N_13893);
xnor U14890 (N_14890,N_13399,N_13560);
nand U14891 (N_14891,N_13095,N_13824);
nand U14892 (N_14892,N_13349,N_13667);
xnor U14893 (N_14893,N_13270,N_13922);
nor U14894 (N_14894,N_13752,N_13440);
xor U14895 (N_14895,N_13531,N_13401);
nor U14896 (N_14896,N_13857,N_13358);
nand U14897 (N_14897,N_13817,N_13636);
nand U14898 (N_14898,N_13868,N_13204);
and U14899 (N_14899,N_13890,N_13187);
or U14900 (N_14900,N_13146,N_13276);
nor U14901 (N_14901,N_13431,N_13882);
xnor U14902 (N_14902,N_13580,N_13844);
or U14903 (N_14903,N_13497,N_13065);
xor U14904 (N_14904,N_13707,N_13458);
or U14905 (N_14905,N_13503,N_13760);
nor U14906 (N_14906,N_13435,N_13011);
and U14907 (N_14907,N_13668,N_13056);
nor U14908 (N_14908,N_13494,N_13203);
nand U14909 (N_14909,N_13501,N_13576);
nand U14910 (N_14910,N_13128,N_13762);
or U14911 (N_14911,N_13171,N_13862);
or U14912 (N_14912,N_13653,N_13858);
xor U14913 (N_14913,N_13920,N_13226);
nor U14914 (N_14914,N_13995,N_13257);
and U14915 (N_14915,N_13271,N_13159);
nand U14916 (N_14916,N_13966,N_13617);
nand U14917 (N_14917,N_13108,N_13268);
nor U14918 (N_14918,N_13926,N_13007);
or U14919 (N_14919,N_13342,N_13711);
xor U14920 (N_14920,N_13164,N_13469);
and U14921 (N_14921,N_13031,N_13661);
nor U14922 (N_14922,N_13669,N_13384);
and U14923 (N_14923,N_13475,N_13563);
or U14924 (N_14924,N_13786,N_13243);
nor U14925 (N_14925,N_13491,N_13819);
xnor U14926 (N_14926,N_13800,N_13608);
and U14927 (N_14927,N_13961,N_13356);
xor U14928 (N_14928,N_13447,N_13989);
nand U14929 (N_14929,N_13654,N_13605);
nor U14930 (N_14930,N_13261,N_13783);
or U14931 (N_14931,N_13903,N_13198);
nand U14932 (N_14932,N_13419,N_13260);
nand U14933 (N_14933,N_13768,N_13523);
or U14934 (N_14934,N_13274,N_13897);
or U14935 (N_14935,N_13343,N_13892);
and U14936 (N_14936,N_13071,N_13239);
and U14937 (N_14937,N_13423,N_13219);
xor U14938 (N_14938,N_13752,N_13877);
xnor U14939 (N_14939,N_13396,N_13162);
and U14940 (N_14940,N_13785,N_13579);
xor U14941 (N_14941,N_13006,N_13998);
and U14942 (N_14942,N_13046,N_13428);
nor U14943 (N_14943,N_13607,N_13395);
xor U14944 (N_14944,N_13087,N_13801);
and U14945 (N_14945,N_13244,N_13825);
nand U14946 (N_14946,N_13073,N_13277);
and U14947 (N_14947,N_13687,N_13129);
xor U14948 (N_14948,N_13698,N_13073);
and U14949 (N_14949,N_13556,N_13715);
or U14950 (N_14950,N_13309,N_13440);
nor U14951 (N_14951,N_13597,N_13442);
xnor U14952 (N_14952,N_13922,N_13000);
and U14953 (N_14953,N_13096,N_13356);
xnor U14954 (N_14954,N_13389,N_13447);
or U14955 (N_14955,N_13238,N_13329);
or U14956 (N_14956,N_13252,N_13110);
nor U14957 (N_14957,N_13598,N_13606);
nand U14958 (N_14958,N_13926,N_13119);
or U14959 (N_14959,N_13272,N_13650);
xnor U14960 (N_14960,N_13605,N_13306);
nor U14961 (N_14961,N_13249,N_13930);
or U14962 (N_14962,N_13856,N_13774);
and U14963 (N_14963,N_13275,N_13012);
or U14964 (N_14964,N_13758,N_13202);
and U14965 (N_14965,N_13550,N_13746);
or U14966 (N_14966,N_13931,N_13907);
and U14967 (N_14967,N_13269,N_13343);
nor U14968 (N_14968,N_13742,N_13788);
nor U14969 (N_14969,N_13823,N_13033);
or U14970 (N_14970,N_13318,N_13282);
nand U14971 (N_14971,N_13423,N_13810);
nor U14972 (N_14972,N_13976,N_13539);
nand U14973 (N_14973,N_13894,N_13850);
or U14974 (N_14974,N_13360,N_13580);
nand U14975 (N_14975,N_13815,N_13042);
and U14976 (N_14976,N_13477,N_13436);
nand U14977 (N_14977,N_13279,N_13732);
and U14978 (N_14978,N_13929,N_13276);
or U14979 (N_14979,N_13624,N_13824);
xnor U14980 (N_14980,N_13167,N_13217);
and U14981 (N_14981,N_13376,N_13413);
nor U14982 (N_14982,N_13823,N_13297);
nand U14983 (N_14983,N_13429,N_13515);
nor U14984 (N_14984,N_13861,N_13470);
and U14985 (N_14985,N_13232,N_13294);
xnor U14986 (N_14986,N_13418,N_13114);
xor U14987 (N_14987,N_13364,N_13062);
or U14988 (N_14988,N_13874,N_13695);
nand U14989 (N_14989,N_13775,N_13028);
or U14990 (N_14990,N_13092,N_13795);
and U14991 (N_14991,N_13220,N_13482);
nand U14992 (N_14992,N_13493,N_13335);
xor U14993 (N_14993,N_13944,N_13265);
nor U14994 (N_14994,N_13062,N_13231);
nor U14995 (N_14995,N_13508,N_13894);
nand U14996 (N_14996,N_13211,N_13259);
or U14997 (N_14997,N_13241,N_13471);
and U14998 (N_14998,N_13192,N_13625);
and U14999 (N_14999,N_13804,N_13047);
xor U15000 (N_15000,N_14156,N_14118);
and U15001 (N_15001,N_14354,N_14802);
or U15002 (N_15002,N_14426,N_14404);
or U15003 (N_15003,N_14159,N_14849);
and U15004 (N_15004,N_14615,N_14377);
nand U15005 (N_15005,N_14359,N_14391);
and U15006 (N_15006,N_14934,N_14878);
and U15007 (N_15007,N_14526,N_14991);
and U15008 (N_15008,N_14613,N_14385);
nand U15009 (N_15009,N_14548,N_14144);
or U15010 (N_15010,N_14501,N_14846);
nor U15011 (N_15011,N_14599,N_14503);
nor U15012 (N_15012,N_14357,N_14128);
xor U15013 (N_15013,N_14004,N_14082);
or U15014 (N_15014,N_14361,N_14198);
nor U15015 (N_15015,N_14561,N_14964);
nand U15016 (N_15016,N_14057,N_14940);
nor U15017 (N_15017,N_14433,N_14437);
or U15018 (N_15018,N_14746,N_14689);
xnor U15019 (N_15019,N_14957,N_14735);
nand U15020 (N_15020,N_14710,N_14738);
xnor U15021 (N_15021,N_14112,N_14324);
or U15022 (N_15022,N_14602,N_14372);
nor U15023 (N_15023,N_14865,N_14789);
xnor U15024 (N_15024,N_14092,N_14723);
and U15025 (N_15025,N_14739,N_14512);
nand U15026 (N_15026,N_14472,N_14708);
nor U15027 (N_15027,N_14392,N_14193);
xnor U15028 (N_15028,N_14380,N_14674);
xor U15029 (N_15029,N_14913,N_14384);
or U15030 (N_15030,N_14105,N_14477);
xnor U15031 (N_15031,N_14311,N_14416);
nor U15032 (N_15032,N_14199,N_14819);
or U15033 (N_15033,N_14217,N_14524);
nor U15034 (N_15034,N_14267,N_14342);
nand U15035 (N_15035,N_14375,N_14451);
and U15036 (N_15036,N_14314,N_14966);
nand U15037 (N_15037,N_14691,N_14232);
or U15038 (N_15038,N_14035,N_14097);
nor U15039 (N_15039,N_14812,N_14823);
or U15040 (N_15040,N_14133,N_14126);
nand U15041 (N_15041,N_14557,N_14420);
and U15042 (N_15042,N_14461,N_14149);
xor U15043 (N_15043,N_14320,N_14347);
or U15044 (N_15044,N_14645,N_14170);
xor U15045 (N_15045,N_14269,N_14210);
nor U15046 (N_15046,N_14047,N_14993);
nand U15047 (N_15047,N_14449,N_14188);
nor U15048 (N_15048,N_14363,N_14860);
and U15049 (N_15049,N_14173,N_14204);
nor U15050 (N_15050,N_14396,N_14318);
or U15051 (N_15051,N_14148,N_14132);
nor U15052 (N_15052,N_14284,N_14489);
and U15053 (N_15053,N_14953,N_14901);
nand U15054 (N_15054,N_14631,N_14587);
nor U15055 (N_15055,N_14495,N_14143);
nand U15056 (N_15056,N_14240,N_14916);
xor U15057 (N_15057,N_14397,N_14300);
xor U15058 (N_15058,N_14681,N_14340);
nand U15059 (N_15059,N_14720,N_14983);
and U15060 (N_15060,N_14381,N_14544);
nor U15061 (N_15061,N_14251,N_14053);
or U15062 (N_15062,N_14833,N_14555);
or U15063 (N_15063,N_14959,N_14002);
or U15064 (N_15064,N_14005,N_14996);
or U15065 (N_15065,N_14929,N_14260);
and U15066 (N_15066,N_14831,N_14475);
and U15067 (N_15067,N_14625,N_14013);
xnor U15068 (N_15068,N_14902,N_14030);
or U15069 (N_15069,N_14688,N_14017);
nor U15070 (N_15070,N_14247,N_14094);
and U15071 (N_15071,N_14768,N_14473);
or U15072 (N_15072,N_14067,N_14226);
nand U15073 (N_15073,N_14784,N_14339);
and U15074 (N_15074,N_14276,N_14265);
and U15075 (N_15075,N_14673,N_14761);
nor U15076 (N_15076,N_14223,N_14037);
and U15077 (N_15077,N_14535,N_14672);
or U15078 (N_15078,N_14273,N_14713);
or U15079 (N_15079,N_14791,N_14301);
or U15080 (N_15080,N_14614,N_14576);
xor U15081 (N_15081,N_14575,N_14671);
nor U15082 (N_15082,N_14182,N_14459);
and U15083 (N_15083,N_14146,N_14923);
nand U15084 (N_15084,N_14732,N_14452);
or U15085 (N_15085,N_14965,N_14487);
and U15086 (N_15086,N_14655,N_14421);
and U15087 (N_15087,N_14060,N_14448);
and U15088 (N_15088,N_14109,N_14563);
nand U15089 (N_15089,N_14491,N_14716);
and U15090 (N_15090,N_14306,N_14838);
or U15091 (N_15091,N_14282,N_14064);
nand U15092 (N_15092,N_14317,N_14656);
nor U15093 (N_15093,N_14443,N_14758);
nor U15094 (N_15094,N_14153,N_14606);
or U15095 (N_15095,N_14863,N_14619);
or U15096 (N_15096,N_14346,N_14830);
or U15097 (N_15097,N_14928,N_14853);
or U15098 (N_15098,N_14087,N_14176);
xnor U15099 (N_15099,N_14436,N_14794);
xor U15100 (N_15100,N_14580,N_14261);
and U15101 (N_15101,N_14400,N_14155);
and U15102 (N_15102,N_14970,N_14231);
and U15103 (N_15103,N_14626,N_14235);
xnor U15104 (N_15104,N_14025,N_14084);
nor U15105 (N_15105,N_14186,N_14291);
nand U15106 (N_15106,N_14683,N_14862);
and U15107 (N_15107,N_14889,N_14056);
xor U15108 (N_15108,N_14401,N_14679);
nand U15109 (N_15109,N_14795,N_14653);
and U15110 (N_15110,N_14597,N_14944);
or U15111 (N_15111,N_14299,N_14869);
nand U15112 (N_15112,N_14010,N_14936);
and U15113 (N_15113,N_14187,N_14102);
xnor U15114 (N_15114,N_14344,N_14727);
xnor U15115 (N_15115,N_14325,N_14113);
or U15116 (N_15116,N_14032,N_14570);
xor U15117 (N_15117,N_14780,N_14603);
and U15118 (N_15118,N_14556,N_14196);
nand U15119 (N_15119,N_14518,N_14814);
nand U15120 (N_15120,N_14158,N_14027);
and U15121 (N_15121,N_14590,N_14506);
nand U15122 (N_15122,N_14793,N_14984);
and U15123 (N_15123,N_14997,N_14922);
xor U15124 (N_15124,N_14079,N_14481);
nand U15125 (N_15125,N_14701,N_14697);
nor U15126 (N_15126,N_14721,N_14191);
xnor U15127 (N_15127,N_14522,N_14090);
and U15128 (N_15128,N_14667,N_14510);
and U15129 (N_15129,N_14546,N_14760);
and U15130 (N_15130,N_14043,N_14935);
and U15131 (N_15131,N_14254,N_14622);
nand U15132 (N_15132,N_14242,N_14729);
nor U15133 (N_15133,N_14020,N_14915);
xor U15134 (N_15134,N_14164,N_14661);
xor U15135 (N_15135,N_14638,N_14938);
or U15136 (N_15136,N_14086,N_14414);
or U15137 (N_15137,N_14909,N_14920);
and U15138 (N_15138,N_14586,N_14600);
or U15139 (N_15139,N_14428,N_14894);
xnor U15140 (N_15140,N_14341,N_14917);
nand U15141 (N_15141,N_14817,N_14755);
nand U15142 (N_15142,N_14685,N_14244);
nand U15143 (N_15143,N_14841,N_14558);
and U15144 (N_15144,N_14539,N_14596);
xnor U15145 (N_15145,N_14330,N_14933);
nand U15146 (N_15146,N_14624,N_14668);
or U15147 (N_15147,N_14537,N_14649);
and U15148 (N_15148,N_14302,N_14618);
or U15149 (N_15149,N_14429,N_14621);
or U15150 (N_15150,N_14435,N_14811);
nor U15151 (N_15151,N_14104,N_14022);
or U15152 (N_15152,N_14887,N_14852);
nor U15153 (N_15153,N_14634,N_14982);
or U15154 (N_15154,N_14771,N_14183);
and U15155 (N_15155,N_14808,N_14099);
and U15156 (N_15156,N_14055,N_14975);
nor U15157 (N_15157,N_14835,N_14338);
nand U15158 (N_15158,N_14085,N_14875);
nor U15159 (N_15159,N_14776,N_14332);
or U15160 (N_15160,N_14026,N_14943);
nand U15161 (N_15161,N_14545,N_14549);
and U15162 (N_15162,N_14932,N_14504);
xor U15163 (N_15163,N_14827,N_14167);
nand U15164 (N_15164,N_14927,N_14759);
nor U15165 (N_15165,N_14677,N_14924);
nor U15166 (N_15166,N_14682,N_14644);
nand U15167 (N_15167,N_14930,N_14999);
nor U15168 (N_15168,N_14772,N_14611);
or U15169 (N_15169,N_14464,N_14439);
or U15170 (N_15170,N_14230,N_14145);
nor U15171 (N_15171,N_14532,N_14093);
or U15172 (N_15172,N_14294,N_14177);
nor U15173 (N_15173,N_14507,N_14492);
and U15174 (N_15174,N_14581,N_14277);
xnor U15175 (N_15175,N_14015,N_14169);
or U15176 (N_15176,N_14029,N_14650);
nand U15177 (N_15177,N_14245,N_14750);
nor U15178 (N_15178,N_14648,N_14637);
and U15179 (N_15179,N_14088,N_14591);
nor U15180 (N_15180,N_14388,N_14463);
nand U15181 (N_15181,N_14947,N_14103);
or U15182 (N_15182,N_14218,N_14365);
or U15183 (N_15183,N_14698,N_14858);
nor U15184 (N_15184,N_14742,N_14528);
nand U15185 (N_15185,N_14327,N_14471);
and U15186 (N_15186,N_14304,N_14166);
and U15187 (N_15187,N_14562,N_14333);
xor U15188 (N_15188,N_14490,N_14257);
nor U15189 (N_15189,N_14309,N_14574);
nand U15190 (N_15190,N_14140,N_14468);
and U15191 (N_15191,N_14214,N_14425);
nor U15192 (N_15192,N_14151,N_14009);
xor U15193 (N_15193,N_14994,N_14350);
nor U15194 (N_15194,N_14237,N_14559);
and U15195 (N_15195,N_14598,N_14798);
or U15196 (N_15196,N_14584,N_14500);
and U15197 (N_15197,N_14807,N_14051);
xor U15198 (N_15198,N_14628,N_14289);
nand U15199 (N_15199,N_14937,N_14142);
nor U15200 (N_15200,N_14730,N_14568);
nand U15201 (N_15201,N_14271,N_14076);
xor U15202 (N_15202,N_14553,N_14121);
nor U15203 (N_15203,N_14221,N_14253);
nand U15204 (N_15204,N_14620,N_14702);
and U15205 (N_15205,N_14859,N_14162);
nor U15206 (N_15206,N_14297,N_14243);
or U15207 (N_15207,N_14378,N_14255);
xor U15208 (N_15208,N_14496,N_14527);
and U15209 (N_15209,N_14881,N_14470);
or U15210 (N_15210,N_14213,N_14680);
nand U15211 (N_15211,N_14855,N_14172);
nand U15212 (N_15212,N_14023,N_14872);
nand U15213 (N_15213,N_14441,N_14896);
xnor U15214 (N_15214,N_14058,N_14305);
nand U15215 (N_15215,N_14577,N_14321);
xor U15216 (N_15216,N_14949,N_14871);
or U15217 (N_15217,N_14456,N_14044);
xor U15218 (N_15218,N_14405,N_14059);
nor U15219 (N_15219,N_14951,N_14116);
or U15220 (N_15220,N_14290,N_14212);
xor U15221 (N_15221,N_14206,N_14345);
xor U15222 (N_15222,N_14762,N_14081);
nor U15223 (N_15223,N_14019,N_14505);
or U15224 (N_15224,N_14885,N_14788);
nor U15225 (N_15225,N_14379,N_14390);
xor U15226 (N_15226,N_14467,N_14786);
nand U15227 (N_15227,N_14856,N_14124);
and U15228 (N_15228,N_14279,N_14753);
and U15229 (N_15229,N_14733,N_14376);
nand U15230 (N_15230,N_14850,N_14248);
nor U15231 (N_15231,N_14709,N_14281);
xor U15232 (N_15232,N_14431,N_14062);
or U15233 (N_15233,N_14236,N_14407);
and U15234 (N_15234,N_14326,N_14669);
nor U15235 (N_15235,N_14063,N_14007);
or U15236 (N_15236,N_14529,N_14373);
and U15237 (N_15237,N_14045,N_14484);
xor U15238 (N_15238,N_14851,N_14643);
nand U15239 (N_15239,N_14465,N_14870);
nor U15240 (N_15240,N_14985,N_14152);
nand U15241 (N_15241,N_14147,N_14815);
xor U15242 (N_15242,N_14402,N_14604);
and U15243 (N_15243,N_14509,N_14482);
nor U15244 (N_15244,N_14640,N_14696);
xor U15245 (N_15245,N_14120,N_14785);
nor U15246 (N_15246,N_14612,N_14411);
nor U15247 (N_15247,N_14160,N_14246);
nand U15248 (N_15248,N_14898,N_14201);
nor U15249 (N_15249,N_14919,N_14741);
nand U15250 (N_15250,N_14796,N_14866);
nand U15251 (N_15251,N_14348,N_14117);
nor U15252 (N_15252,N_14303,N_14962);
nor U15253 (N_15253,N_14781,N_14497);
or U15254 (N_15254,N_14216,N_14816);
nand U15255 (N_15255,N_14387,N_14905);
and U15256 (N_15256,N_14080,N_14038);
xor U15257 (N_15257,N_14419,N_14770);
nand U15258 (N_15258,N_14829,N_14498);
xor U15259 (N_15259,N_14207,N_14971);
nor U15260 (N_15260,N_14534,N_14605);
nor U15261 (N_15261,N_14123,N_14594);
nand U15262 (N_15262,N_14399,N_14891);
and U15263 (N_15263,N_14783,N_14179);
nand U15264 (N_15264,N_14538,N_14515);
or U15265 (N_15265,N_14782,N_14728);
nand U15266 (N_15266,N_14973,N_14046);
or U15267 (N_15267,N_14111,N_14945);
nand U15268 (N_15268,N_14234,N_14367);
nand U15269 (N_15269,N_14266,N_14961);
nand U15270 (N_15270,N_14749,N_14694);
and U15271 (N_15271,N_14189,N_14393);
nand U15272 (N_15272,N_14184,N_14968);
xor U15273 (N_15273,N_14194,N_14593);
xor U15274 (N_15274,N_14130,N_14219);
and U15275 (N_15275,N_14434,N_14692);
or U15276 (N_15276,N_14228,N_14748);
nand U15277 (N_15277,N_14826,N_14034);
and U15278 (N_15278,N_14369,N_14886);
or U15279 (N_15279,N_14647,N_14601);
nand U15280 (N_15280,N_14180,N_14907);
and U15281 (N_15281,N_14288,N_14800);
or U15282 (N_15282,N_14980,N_14664);
and U15283 (N_15283,N_14890,N_14520);
nand U15284 (N_15284,N_14211,N_14939);
nand U15285 (N_15285,N_14734,N_14633);
nor U15286 (N_15286,N_14892,N_14777);
nand U15287 (N_15287,N_14114,N_14368);
nand U15288 (N_15288,N_14089,N_14845);
xor U15289 (N_15289,N_14163,N_14494);
or U15290 (N_15290,N_14722,N_14233);
and U15291 (N_15291,N_14926,N_14810);
or U15292 (N_15292,N_14447,N_14867);
and U15293 (N_15293,N_14293,N_14629);
xnor U15294 (N_15294,N_14003,N_14285);
xor U15295 (N_15295,N_14048,N_14565);
and U15296 (N_15296,N_14806,N_14747);
nor U15297 (N_15297,N_14115,N_14229);
and U15298 (N_15298,N_14705,N_14769);
or U15299 (N_15299,N_14925,N_14715);
nand U15300 (N_15300,N_14918,N_14660);
or U15301 (N_15301,N_14403,N_14541);
nand U15302 (N_15302,N_14767,N_14566);
xor U15303 (N_15303,N_14882,N_14262);
nor U15304 (N_15304,N_14988,N_14220);
xor U15305 (N_15305,N_14567,N_14323);
nor U15306 (N_15306,N_14954,N_14275);
nand U15307 (N_15307,N_14595,N_14824);
xnor U15308 (N_15308,N_14825,N_14848);
xor U15309 (N_15309,N_14479,N_14844);
xnor U15310 (N_15310,N_14676,N_14197);
xnor U15311 (N_15311,N_14171,N_14989);
nor U15312 (N_15312,N_14805,N_14139);
xor U15313 (N_15313,N_14445,N_14942);
nand U15314 (N_15314,N_14249,N_14724);
xor U15315 (N_15315,N_14745,N_14790);
or U15316 (N_15316,N_14427,N_14474);
xnor U15317 (N_15317,N_14582,N_14502);
nor U15318 (N_15318,N_14836,N_14021);
xnor U15319 (N_15319,N_14774,N_14238);
or U15320 (N_15320,N_14134,N_14879);
nor U15321 (N_15321,N_14684,N_14315);
xnor U15322 (N_15322,N_14083,N_14740);
nor U15323 (N_15323,N_14349,N_14054);
and U15324 (N_15324,N_14259,N_14398);
nand U15325 (N_15325,N_14061,N_14642);
xor U15326 (N_15326,N_14884,N_14704);
xnor U15327 (N_15327,N_14900,N_14412);
and U15328 (N_15328,N_14066,N_14039);
xor U15329 (N_15329,N_14658,N_14707);
and U15330 (N_15330,N_14091,N_14070);
nor U15331 (N_15331,N_14921,N_14799);
xor U15332 (N_15332,N_14178,N_14543);
or U15333 (N_15333,N_14787,N_14700);
or U15334 (N_15334,N_14639,N_14876);
nor U15335 (N_15335,N_14334,N_14014);
nand U15336 (N_15336,N_14395,N_14573);
xnor U15337 (N_15337,N_14979,N_14822);
nor U15338 (N_15338,N_14880,N_14508);
and U15339 (N_15339,N_14071,N_14736);
or U15340 (N_15340,N_14157,N_14636);
nor U15341 (N_15341,N_14287,N_14554);
xor U15342 (N_15342,N_14239,N_14313);
nand U15343 (N_15343,N_14356,N_14296);
nor U15344 (N_15344,N_14442,N_14222);
xor U15345 (N_15345,N_14589,N_14531);
and U15346 (N_15346,N_14828,N_14803);
and U15347 (N_15347,N_14352,N_14072);
and U15348 (N_15348,N_14609,N_14731);
xnor U15349 (N_15349,N_14737,N_14024);
nand U15350 (N_15350,N_14389,N_14406);
nand U15351 (N_15351,N_14270,N_14857);
and U15352 (N_15352,N_14224,N_14726);
nor U15353 (N_15353,N_14560,N_14422);
nand U15354 (N_15354,N_14711,N_14394);
xnor U15355 (N_15355,N_14756,N_14610);
xor U15356 (N_15356,N_14174,N_14635);
and U15357 (N_15357,N_14202,N_14847);
xor U15358 (N_15358,N_14329,N_14280);
nand U15359 (N_15359,N_14948,N_14252);
and U15360 (N_15360,N_14154,N_14763);
nor U15361 (N_15361,N_14779,N_14241);
nor U15362 (N_15362,N_14227,N_14525);
xor U15363 (N_15363,N_14670,N_14382);
nor U15364 (N_15364,N_14131,N_14873);
and U15365 (N_15365,N_14675,N_14078);
nand U15366 (N_15366,N_14579,N_14536);
nor U15367 (N_15367,N_14754,N_14564);
xor U15368 (N_15368,N_14818,N_14699);
xor U15369 (N_15369,N_14883,N_14488);
or U15370 (N_15370,N_14200,N_14617);
xor U15371 (N_15371,N_14190,N_14572);
nor U15372 (N_15372,N_14264,N_14274);
nor U15373 (N_15373,N_14351,N_14813);
or U15374 (N_15374,N_14757,N_14513);
xnor U15375 (N_15375,N_14977,N_14050);
and U15376 (N_15376,N_14272,N_14328);
and U15377 (N_15377,N_14129,N_14832);
xnor U15378 (N_15378,N_14141,N_14998);
or U15379 (N_15379,N_14941,N_14308);
and U15380 (N_15380,N_14417,N_14161);
nor U15381 (N_15381,N_14001,N_14652);
xnor U15382 (N_15382,N_14225,N_14460);
nand U15383 (N_15383,N_14583,N_14018);
xor U15384 (N_15384,N_14840,N_14992);
and U15385 (N_15385,N_14911,N_14455);
nor U15386 (N_15386,N_14410,N_14972);
nand U15387 (N_15387,N_14530,N_14974);
xnor U15388 (N_15388,N_14842,N_14519);
and U15389 (N_15389,N_14665,N_14904);
nor U15390 (N_15390,N_14310,N_14874);
nand U15391 (N_15391,N_14343,N_14792);
and U15392 (N_15392,N_14585,N_14523);
nor U15393 (N_15393,N_14976,N_14215);
or U15394 (N_15394,N_14136,N_14374);
xnor U15395 (N_15395,N_14627,N_14571);
or U15396 (N_15396,N_14820,N_14335);
nor U15397 (N_15397,N_14371,N_14666);
or U15398 (N_15398,N_14250,N_14719);
nand U15399 (N_15399,N_14485,N_14963);
nor U15400 (N_15400,N_14322,N_14775);
or U15401 (N_15401,N_14821,N_14843);
xor U15402 (N_15402,N_14712,N_14175);
nor U15403 (N_15403,N_14370,N_14469);
and U15404 (N_15404,N_14108,N_14077);
xor U15405 (N_15405,N_14517,N_14074);
and U15406 (N_15406,N_14483,N_14877);
nand U15407 (N_15407,N_14868,N_14444);
nand U15408 (N_15408,N_14542,N_14854);
and U15409 (N_15409,N_14906,N_14990);
nand U15410 (N_15410,N_14286,N_14967);
nor U15411 (N_15411,N_14458,N_14861);
or U15412 (N_15412,N_14511,N_14106);
xnor U15413 (N_15413,N_14457,N_14068);
and U15414 (N_15414,N_14307,N_14016);
xor U15415 (N_15415,N_14098,N_14119);
or U15416 (N_15416,N_14337,N_14897);
nand U15417 (N_15417,N_14192,N_14478);
nand U15418 (N_15418,N_14778,N_14075);
and U15419 (N_15419,N_14150,N_14298);
nand U15420 (N_15420,N_14205,N_14764);
nand U15421 (N_15421,N_14413,N_14987);
nor U15422 (N_15422,N_14041,N_14899);
nor U15423 (N_15423,N_14839,N_14283);
nand U15424 (N_15424,N_14608,N_14662);
and U15425 (N_15425,N_14446,N_14008);
xnor U15426 (N_15426,N_14895,N_14706);
xor U15427 (N_15427,N_14765,N_14258);
xor U15428 (N_15428,N_14100,N_14552);
or U15429 (N_15429,N_14168,N_14012);
and U15430 (N_15430,N_14903,N_14550);
nor U15431 (N_15431,N_14547,N_14033);
and U15432 (N_15432,N_14383,N_14096);
nand U15433 (N_15433,N_14744,N_14127);
nor U15434 (N_15434,N_14981,N_14203);
nor U15435 (N_15435,N_14908,N_14743);
nor U15436 (N_15436,N_14521,N_14837);
xor U15437 (N_15437,N_14956,N_14000);
and U15438 (N_15438,N_14362,N_14268);
xor U15439 (N_15439,N_14540,N_14773);
or U15440 (N_15440,N_14569,N_14718);
or U15441 (N_15441,N_14687,N_14424);
or U15442 (N_15442,N_14138,N_14185);
or U15443 (N_15443,N_14693,N_14809);
and U15444 (N_15444,N_14678,N_14137);
nand U15445 (N_15445,N_14031,N_14052);
nand U15446 (N_15446,N_14946,N_14319);
nand U15447 (N_15447,N_14292,N_14028);
xor U15448 (N_15448,N_14011,N_14751);
and U15449 (N_15449,N_14125,N_14766);
or U15450 (N_15450,N_14423,N_14657);
and U15451 (N_15451,N_14366,N_14432);
nor U15452 (N_15452,N_14358,N_14752);
and U15453 (N_15453,N_14960,N_14466);
nand U15454 (N_15454,N_14654,N_14592);
or U15455 (N_15455,N_14036,N_14632);
xnor U15456 (N_15456,N_14408,N_14360);
nand U15457 (N_15457,N_14295,N_14893);
xor U15458 (N_15458,N_14797,N_14516);
and U15459 (N_15459,N_14006,N_14914);
or U15460 (N_15460,N_14195,N_14430);
or U15461 (N_15461,N_14952,N_14486);
or U15462 (N_15462,N_14493,N_14386);
xnor U15463 (N_15463,N_14065,N_14514);
xnor U15464 (N_15464,N_14480,N_14256);
nor U15465 (N_15465,N_14073,N_14355);
nand U15466 (N_15466,N_14616,N_14101);
xor U15467 (N_15467,N_14418,N_14588);
or U15468 (N_15468,N_14208,N_14476);
xor U15469 (N_15469,N_14438,N_14331);
nor U15470 (N_15470,N_14110,N_14263);
nor U15471 (N_15471,N_14415,N_14703);
and U15472 (N_15472,N_14978,N_14040);
and U15473 (N_15473,N_14533,N_14107);
nand U15474 (N_15474,N_14095,N_14440);
nor U15475 (N_15475,N_14714,N_14641);
xor U15476 (N_15476,N_14955,N_14630);
or U15477 (N_15477,N_14364,N_14165);
xnor U15478 (N_15478,N_14686,N_14042);
nand U15479 (N_15479,N_14578,N_14607);
nand U15480 (N_15480,N_14834,N_14801);
xor U15481 (N_15481,N_14659,N_14986);
nand U15482 (N_15482,N_14181,N_14353);
or U15483 (N_15483,N_14049,N_14912);
nand U15484 (N_15484,N_14312,N_14695);
nand U15485 (N_15485,N_14336,N_14910);
nor U15486 (N_15486,N_14462,N_14209);
and U15487 (N_15487,N_14725,N_14278);
xor U15488 (N_15488,N_14969,N_14995);
nor U15489 (N_15489,N_14454,N_14646);
nor U15490 (N_15490,N_14453,N_14888);
xnor U15491 (N_15491,N_14450,N_14651);
or U15492 (N_15492,N_14717,N_14135);
xor U15493 (N_15493,N_14950,N_14499);
or U15494 (N_15494,N_14663,N_14931);
or U15495 (N_15495,N_14122,N_14864);
xnor U15496 (N_15496,N_14551,N_14958);
nor U15497 (N_15497,N_14690,N_14409);
xnor U15498 (N_15498,N_14069,N_14804);
nand U15499 (N_15499,N_14623,N_14316);
xor U15500 (N_15500,N_14320,N_14022);
nand U15501 (N_15501,N_14090,N_14624);
and U15502 (N_15502,N_14489,N_14721);
xor U15503 (N_15503,N_14315,N_14917);
nand U15504 (N_15504,N_14882,N_14625);
nand U15505 (N_15505,N_14104,N_14313);
nor U15506 (N_15506,N_14351,N_14279);
nor U15507 (N_15507,N_14428,N_14877);
nor U15508 (N_15508,N_14223,N_14293);
and U15509 (N_15509,N_14464,N_14592);
nor U15510 (N_15510,N_14531,N_14739);
nand U15511 (N_15511,N_14317,N_14242);
and U15512 (N_15512,N_14705,N_14198);
xnor U15513 (N_15513,N_14527,N_14034);
nand U15514 (N_15514,N_14663,N_14413);
nor U15515 (N_15515,N_14808,N_14943);
or U15516 (N_15516,N_14347,N_14273);
and U15517 (N_15517,N_14357,N_14188);
or U15518 (N_15518,N_14227,N_14753);
nor U15519 (N_15519,N_14151,N_14215);
or U15520 (N_15520,N_14247,N_14294);
or U15521 (N_15521,N_14855,N_14631);
or U15522 (N_15522,N_14069,N_14682);
nand U15523 (N_15523,N_14327,N_14629);
and U15524 (N_15524,N_14991,N_14842);
nor U15525 (N_15525,N_14409,N_14726);
or U15526 (N_15526,N_14355,N_14642);
or U15527 (N_15527,N_14574,N_14072);
and U15528 (N_15528,N_14030,N_14130);
or U15529 (N_15529,N_14746,N_14634);
xor U15530 (N_15530,N_14804,N_14542);
and U15531 (N_15531,N_14835,N_14992);
nand U15532 (N_15532,N_14672,N_14750);
nand U15533 (N_15533,N_14183,N_14626);
xor U15534 (N_15534,N_14726,N_14533);
and U15535 (N_15535,N_14549,N_14176);
or U15536 (N_15536,N_14037,N_14679);
nor U15537 (N_15537,N_14552,N_14159);
xnor U15538 (N_15538,N_14533,N_14547);
nand U15539 (N_15539,N_14761,N_14967);
xor U15540 (N_15540,N_14299,N_14333);
nand U15541 (N_15541,N_14476,N_14831);
nor U15542 (N_15542,N_14189,N_14728);
or U15543 (N_15543,N_14389,N_14231);
nor U15544 (N_15544,N_14043,N_14889);
and U15545 (N_15545,N_14762,N_14303);
xnor U15546 (N_15546,N_14746,N_14977);
and U15547 (N_15547,N_14512,N_14352);
and U15548 (N_15548,N_14404,N_14707);
nand U15549 (N_15549,N_14002,N_14061);
nor U15550 (N_15550,N_14857,N_14576);
xor U15551 (N_15551,N_14889,N_14371);
nand U15552 (N_15552,N_14439,N_14725);
or U15553 (N_15553,N_14967,N_14614);
and U15554 (N_15554,N_14952,N_14115);
nor U15555 (N_15555,N_14979,N_14157);
nor U15556 (N_15556,N_14332,N_14945);
nand U15557 (N_15557,N_14650,N_14797);
xor U15558 (N_15558,N_14863,N_14795);
and U15559 (N_15559,N_14714,N_14669);
xnor U15560 (N_15560,N_14983,N_14480);
and U15561 (N_15561,N_14781,N_14923);
and U15562 (N_15562,N_14215,N_14766);
nor U15563 (N_15563,N_14331,N_14821);
and U15564 (N_15564,N_14263,N_14058);
xor U15565 (N_15565,N_14919,N_14602);
nand U15566 (N_15566,N_14279,N_14192);
nand U15567 (N_15567,N_14938,N_14846);
nand U15568 (N_15568,N_14877,N_14941);
xor U15569 (N_15569,N_14514,N_14479);
or U15570 (N_15570,N_14507,N_14880);
and U15571 (N_15571,N_14260,N_14785);
or U15572 (N_15572,N_14864,N_14517);
nor U15573 (N_15573,N_14162,N_14683);
xnor U15574 (N_15574,N_14656,N_14525);
or U15575 (N_15575,N_14136,N_14954);
or U15576 (N_15576,N_14599,N_14935);
nor U15577 (N_15577,N_14772,N_14678);
nand U15578 (N_15578,N_14608,N_14494);
nor U15579 (N_15579,N_14702,N_14442);
nand U15580 (N_15580,N_14844,N_14297);
nor U15581 (N_15581,N_14258,N_14069);
and U15582 (N_15582,N_14747,N_14940);
nor U15583 (N_15583,N_14819,N_14240);
xor U15584 (N_15584,N_14697,N_14533);
nand U15585 (N_15585,N_14527,N_14384);
xnor U15586 (N_15586,N_14995,N_14784);
or U15587 (N_15587,N_14655,N_14886);
and U15588 (N_15588,N_14275,N_14606);
xor U15589 (N_15589,N_14507,N_14678);
or U15590 (N_15590,N_14874,N_14230);
xnor U15591 (N_15591,N_14155,N_14892);
and U15592 (N_15592,N_14109,N_14657);
nand U15593 (N_15593,N_14596,N_14880);
nand U15594 (N_15594,N_14574,N_14048);
xnor U15595 (N_15595,N_14519,N_14464);
or U15596 (N_15596,N_14552,N_14704);
nand U15597 (N_15597,N_14714,N_14755);
or U15598 (N_15598,N_14959,N_14651);
and U15599 (N_15599,N_14567,N_14821);
and U15600 (N_15600,N_14819,N_14150);
nor U15601 (N_15601,N_14593,N_14762);
nor U15602 (N_15602,N_14085,N_14332);
nand U15603 (N_15603,N_14878,N_14931);
xnor U15604 (N_15604,N_14477,N_14547);
nor U15605 (N_15605,N_14744,N_14178);
and U15606 (N_15606,N_14740,N_14990);
xnor U15607 (N_15607,N_14804,N_14225);
and U15608 (N_15608,N_14264,N_14935);
or U15609 (N_15609,N_14644,N_14394);
nor U15610 (N_15610,N_14019,N_14842);
nor U15611 (N_15611,N_14629,N_14918);
and U15612 (N_15612,N_14853,N_14919);
nor U15613 (N_15613,N_14053,N_14199);
and U15614 (N_15614,N_14558,N_14620);
nand U15615 (N_15615,N_14371,N_14723);
nor U15616 (N_15616,N_14926,N_14637);
nor U15617 (N_15617,N_14928,N_14494);
or U15618 (N_15618,N_14707,N_14454);
nor U15619 (N_15619,N_14764,N_14632);
or U15620 (N_15620,N_14871,N_14457);
and U15621 (N_15621,N_14686,N_14170);
nand U15622 (N_15622,N_14580,N_14740);
nand U15623 (N_15623,N_14634,N_14124);
xnor U15624 (N_15624,N_14840,N_14750);
xnor U15625 (N_15625,N_14324,N_14387);
nand U15626 (N_15626,N_14351,N_14814);
nor U15627 (N_15627,N_14216,N_14925);
nor U15628 (N_15628,N_14036,N_14340);
nand U15629 (N_15629,N_14409,N_14800);
nand U15630 (N_15630,N_14619,N_14688);
or U15631 (N_15631,N_14449,N_14574);
nand U15632 (N_15632,N_14856,N_14165);
and U15633 (N_15633,N_14033,N_14353);
xor U15634 (N_15634,N_14470,N_14448);
nor U15635 (N_15635,N_14977,N_14713);
or U15636 (N_15636,N_14860,N_14685);
and U15637 (N_15637,N_14005,N_14429);
and U15638 (N_15638,N_14165,N_14029);
and U15639 (N_15639,N_14022,N_14298);
nor U15640 (N_15640,N_14890,N_14304);
nand U15641 (N_15641,N_14675,N_14856);
or U15642 (N_15642,N_14672,N_14419);
xor U15643 (N_15643,N_14096,N_14967);
nor U15644 (N_15644,N_14441,N_14256);
or U15645 (N_15645,N_14142,N_14115);
nand U15646 (N_15646,N_14013,N_14220);
nand U15647 (N_15647,N_14535,N_14838);
nand U15648 (N_15648,N_14533,N_14172);
xnor U15649 (N_15649,N_14897,N_14329);
or U15650 (N_15650,N_14289,N_14208);
or U15651 (N_15651,N_14249,N_14827);
xnor U15652 (N_15652,N_14633,N_14186);
nor U15653 (N_15653,N_14492,N_14566);
or U15654 (N_15654,N_14321,N_14367);
nand U15655 (N_15655,N_14065,N_14927);
nor U15656 (N_15656,N_14704,N_14266);
nand U15657 (N_15657,N_14831,N_14249);
and U15658 (N_15658,N_14316,N_14289);
and U15659 (N_15659,N_14696,N_14743);
and U15660 (N_15660,N_14368,N_14216);
or U15661 (N_15661,N_14968,N_14481);
and U15662 (N_15662,N_14210,N_14577);
xor U15663 (N_15663,N_14406,N_14847);
or U15664 (N_15664,N_14739,N_14317);
and U15665 (N_15665,N_14566,N_14156);
and U15666 (N_15666,N_14629,N_14999);
xor U15667 (N_15667,N_14549,N_14842);
or U15668 (N_15668,N_14497,N_14329);
xnor U15669 (N_15669,N_14869,N_14906);
nor U15670 (N_15670,N_14147,N_14645);
and U15671 (N_15671,N_14144,N_14920);
xor U15672 (N_15672,N_14358,N_14087);
nor U15673 (N_15673,N_14548,N_14890);
xor U15674 (N_15674,N_14794,N_14883);
nor U15675 (N_15675,N_14256,N_14808);
nor U15676 (N_15676,N_14969,N_14315);
xnor U15677 (N_15677,N_14517,N_14229);
and U15678 (N_15678,N_14218,N_14389);
nand U15679 (N_15679,N_14216,N_14980);
or U15680 (N_15680,N_14208,N_14686);
nand U15681 (N_15681,N_14535,N_14106);
and U15682 (N_15682,N_14178,N_14445);
or U15683 (N_15683,N_14249,N_14207);
nand U15684 (N_15684,N_14523,N_14535);
or U15685 (N_15685,N_14474,N_14810);
nand U15686 (N_15686,N_14900,N_14749);
and U15687 (N_15687,N_14774,N_14381);
and U15688 (N_15688,N_14147,N_14728);
and U15689 (N_15689,N_14057,N_14010);
and U15690 (N_15690,N_14554,N_14902);
or U15691 (N_15691,N_14888,N_14156);
and U15692 (N_15692,N_14344,N_14462);
xor U15693 (N_15693,N_14219,N_14599);
xor U15694 (N_15694,N_14161,N_14285);
nor U15695 (N_15695,N_14128,N_14312);
nand U15696 (N_15696,N_14938,N_14976);
nor U15697 (N_15697,N_14834,N_14276);
nand U15698 (N_15698,N_14752,N_14134);
or U15699 (N_15699,N_14408,N_14277);
nand U15700 (N_15700,N_14574,N_14264);
or U15701 (N_15701,N_14998,N_14112);
and U15702 (N_15702,N_14226,N_14512);
nand U15703 (N_15703,N_14477,N_14968);
nand U15704 (N_15704,N_14151,N_14524);
or U15705 (N_15705,N_14819,N_14827);
nand U15706 (N_15706,N_14117,N_14821);
or U15707 (N_15707,N_14641,N_14707);
nand U15708 (N_15708,N_14241,N_14162);
nand U15709 (N_15709,N_14310,N_14408);
xor U15710 (N_15710,N_14235,N_14923);
xor U15711 (N_15711,N_14536,N_14531);
or U15712 (N_15712,N_14555,N_14525);
xor U15713 (N_15713,N_14211,N_14598);
or U15714 (N_15714,N_14519,N_14063);
nand U15715 (N_15715,N_14262,N_14953);
nand U15716 (N_15716,N_14365,N_14888);
and U15717 (N_15717,N_14901,N_14101);
nor U15718 (N_15718,N_14445,N_14010);
nor U15719 (N_15719,N_14586,N_14838);
and U15720 (N_15720,N_14701,N_14361);
or U15721 (N_15721,N_14572,N_14973);
or U15722 (N_15722,N_14562,N_14786);
nor U15723 (N_15723,N_14237,N_14764);
nor U15724 (N_15724,N_14588,N_14546);
and U15725 (N_15725,N_14196,N_14181);
or U15726 (N_15726,N_14281,N_14712);
nand U15727 (N_15727,N_14665,N_14174);
nand U15728 (N_15728,N_14469,N_14280);
or U15729 (N_15729,N_14516,N_14126);
and U15730 (N_15730,N_14253,N_14293);
xor U15731 (N_15731,N_14980,N_14954);
xnor U15732 (N_15732,N_14326,N_14313);
nand U15733 (N_15733,N_14922,N_14193);
nand U15734 (N_15734,N_14486,N_14877);
xnor U15735 (N_15735,N_14345,N_14297);
nor U15736 (N_15736,N_14520,N_14775);
nand U15737 (N_15737,N_14627,N_14520);
or U15738 (N_15738,N_14610,N_14879);
nor U15739 (N_15739,N_14002,N_14145);
xnor U15740 (N_15740,N_14026,N_14685);
and U15741 (N_15741,N_14565,N_14273);
nand U15742 (N_15742,N_14116,N_14213);
xor U15743 (N_15743,N_14792,N_14897);
nand U15744 (N_15744,N_14827,N_14265);
and U15745 (N_15745,N_14270,N_14078);
and U15746 (N_15746,N_14567,N_14186);
nand U15747 (N_15747,N_14606,N_14392);
nor U15748 (N_15748,N_14052,N_14980);
xor U15749 (N_15749,N_14878,N_14702);
xnor U15750 (N_15750,N_14319,N_14060);
nor U15751 (N_15751,N_14649,N_14429);
and U15752 (N_15752,N_14376,N_14445);
and U15753 (N_15753,N_14041,N_14414);
xor U15754 (N_15754,N_14289,N_14759);
xor U15755 (N_15755,N_14791,N_14777);
xnor U15756 (N_15756,N_14475,N_14015);
and U15757 (N_15757,N_14922,N_14905);
and U15758 (N_15758,N_14565,N_14098);
xor U15759 (N_15759,N_14196,N_14735);
nand U15760 (N_15760,N_14588,N_14166);
and U15761 (N_15761,N_14630,N_14735);
nand U15762 (N_15762,N_14098,N_14650);
nor U15763 (N_15763,N_14899,N_14827);
xor U15764 (N_15764,N_14193,N_14153);
or U15765 (N_15765,N_14606,N_14795);
nor U15766 (N_15766,N_14837,N_14610);
nand U15767 (N_15767,N_14528,N_14676);
nor U15768 (N_15768,N_14078,N_14165);
and U15769 (N_15769,N_14166,N_14139);
nor U15770 (N_15770,N_14919,N_14343);
and U15771 (N_15771,N_14063,N_14891);
xor U15772 (N_15772,N_14596,N_14521);
nand U15773 (N_15773,N_14561,N_14091);
nor U15774 (N_15774,N_14292,N_14737);
nor U15775 (N_15775,N_14994,N_14193);
nand U15776 (N_15776,N_14878,N_14335);
nor U15777 (N_15777,N_14823,N_14093);
nand U15778 (N_15778,N_14248,N_14280);
or U15779 (N_15779,N_14618,N_14751);
and U15780 (N_15780,N_14957,N_14632);
or U15781 (N_15781,N_14043,N_14667);
xnor U15782 (N_15782,N_14990,N_14586);
xnor U15783 (N_15783,N_14434,N_14255);
nor U15784 (N_15784,N_14358,N_14894);
nand U15785 (N_15785,N_14445,N_14409);
nor U15786 (N_15786,N_14398,N_14901);
nand U15787 (N_15787,N_14182,N_14039);
and U15788 (N_15788,N_14826,N_14119);
and U15789 (N_15789,N_14219,N_14636);
or U15790 (N_15790,N_14498,N_14200);
or U15791 (N_15791,N_14346,N_14804);
nand U15792 (N_15792,N_14537,N_14016);
nor U15793 (N_15793,N_14990,N_14235);
nor U15794 (N_15794,N_14359,N_14450);
xnor U15795 (N_15795,N_14430,N_14815);
or U15796 (N_15796,N_14522,N_14606);
nand U15797 (N_15797,N_14196,N_14353);
xnor U15798 (N_15798,N_14243,N_14768);
xor U15799 (N_15799,N_14217,N_14739);
nand U15800 (N_15800,N_14208,N_14116);
nand U15801 (N_15801,N_14815,N_14878);
nand U15802 (N_15802,N_14888,N_14261);
nor U15803 (N_15803,N_14545,N_14758);
and U15804 (N_15804,N_14968,N_14040);
or U15805 (N_15805,N_14459,N_14048);
or U15806 (N_15806,N_14384,N_14535);
or U15807 (N_15807,N_14783,N_14120);
nand U15808 (N_15808,N_14612,N_14637);
or U15809 (N_15809,N_14822,N_14892);
and U15810 (N_15810,N_14459,N_14561);
nand U15811 (N_15811,N_14150,N_14122);
nor U15812 (N_15812,N_14271,N_14560);
nand U15813 (N_15813,N_14561,N_14348);
xnor U15814 (N_15814,N_14734,N_14298);
nand U15815 (N_15815,N_14370,N_14823);
or U15816 (N_15816,N_14642,N_14450);
xnor U15817 (N_15817,N_14250,N_14524);
or U15818 (N_15818,N_14878,N_14944);
nand U15819 (N_15819,N_14099,N_14406);
xnor U15820 (N_15820,N_14722,N_14719);
nand U15821 (N_15821,N_14621,N_14823);
xnor U15822 (N_15822,N_14426,N_14504);
and U15823 (N_15823,N_14603,N_14128);
nand U15824 (N_15824,N_14364,N_14739);
nand U15825 (N_15825,N_14279,N_14779);
and U15826 (N_15826,N_14728,N_14166);
and U15827 (N_15827,N_14680,N_14631);
nor U15828 (N_15828,N_14095,N_14406);
nor U15829 (N_15829,N_14790,N_14515);
and U15830 (N_15830,N_14505,N_14280);
nor U15831 (N_15831,N_14029,N_14312);
nor U15832 (N_15832,N_14529,N_14595);
or U15833 (N_15833,N_14494,N_14262);
nand U15834 (N_15834,N_14146,N_14525);
and U15835 (N_15835,N_14148,N_14916);
xor U15836 (N_15836,N_14062,N_14677);
and U15837 (N_15837,N_14510,N_14947);
nor U15838 (N_15838,N_14710,N_14801);
nor U15839 (N_15839,N_14530,N_14479);
nor U15840 (N_15840,N_14900,N_14010);
xnor U15841 (N_15841,N_14410,N_14578);
xnor U15842 (N_15842,N_14187,N_14834);
and U15843 (N_15843,N_14734,N_14338);
or U15844 (N_15844,N_14766,N_14043);
nor U15845 (N_15845,N_14928,N_14187);
and U15846 (N_15846,N_14008,N_14516);
xor U15847 (N_15847,N_14879,N_14035);
nor U15848 (N_15848,N_14263,N_14428);
nor U15849 (N_15849,N_14356,N_14708);
nor U15850 (N_15850,N_14321,N_14876);
or U15851 (N_15851,N_14328,N_14452);
xor U15852 (N_15852,N_14918,N_14939);
nand U15853 (N_15853,N_14631,N_14448);
xnor U15854 (N_15854,N_14246,N_14289);
or U15855 (N_15855,N_14054,N_14153);
nor U15856 (N_15856,N_14065,N_14811);
and U15857 (N_15857,N_14336,N_14084);
and U15858 (N_15858,N_14678,N_14496);
xnor U15859 (N_15859,N_14797,N_14929);
and U15860 (N_15860,N_14839,N_14439);
xor U15861 (N_15861,N_14750,N_14580);
nand U15862 (N_15862,N_14745,N_14833);
or U15863 (N_15863,N_14558,N_14743);
nor U15864 (N_15864,N_14585,N_14224);
xor U15865 (N_15865,N_14814,N_14523);
nor U15866 (N_15866,N_14222,N_14175);
nor U15867 (N_15867,N_14564,N_14222);
xnor U15868 (N_15868,N_14290,N_14968);
xnor U15869 (N_15869,N_14542,N_14304);
nor U15870 (N_15870,N_14701,N_14516);
nor U15871 (N_15871,N_14643,N_14482);
nand U15872 (N_15872,N_14542,N_14930);
or U15873 (N_15873,N_14311,N_14422);
and U15874 (N_15874,N_14529,N_14649);
nor U15875 (N_15875,N_14745,N_14565);
or U15876 (N_15876,N_14691,N_14546);
and U15877 (N_15877,N_14766,N_14926);
nand U15878 (N_15878,N_14919,N_14463);
or U15879 (N_15879,N_14221,N_14626);
xor U15880 (N_15880,N_14057,N_14453);
nand U15881 (N_15881,N_14129,N_14634);
nand U15882 (N_15882,N_14490,N_14912);
or U15883 (N_15883,N_14105,N_14896);
and U15884 (N_15884,N_14456,N_14022);
nand U15885 (N_15885,N_14171,N_14079);
nor U15886 (N_15886,N_14049,N_14954);
nand U15887 (N_15887,N_14691,N_14079);
or U15888 (N_15888,N_14691,N_14349);
nor U15889 (N_15889,N_14817,N_14525);
and U15890 (N_15890,N_14664,N_14266);
xor U15891 (N_15891,N_14631,N_14220);
or U15892 (N_15892,N_14249,N_14052);
nand U15893 (N_15893,N_14310,N_14761);
and U15894 (N_15894,N_14325,N_14012);
nand U15895 (N_15895,N_14228,N_14843);
nor U15896 (N_15896,N_14192,N_14087);
nor U15897 (N_15897,N_14315,N_14072);
xnor U15898 (N_15898,N_14766,N_14361);
and U15899 (N_15899,N_14447,N_14217);
nand U15900 (N_15900,N_14374,N_14936);
or U15901 (N_15901,N_14736,N_14974);
nor U15902 (N_15902,N_14097,N_14908);
and U15903 (N_15903,N_14622,N_14377);
nand U15904 (N_15904,N_14013,N_14187);
or U15905 (N_15905,N_14136,N_14224);
nand U15906 (N_15906,N_14915,N_14030);
or U15907 (N_15907,N_14194,N_14317);
and U15908 (N_15908,N_14726,N_14776);
nand U15909 (N_15909,N_14714,N_14214);
nor U15910 (N_15910,N_14493,N_14511);
and U15911 (N_15911,N_14915,N_14873);
nor U15912 (N_15912,N_14855,N_14405);
nand U15913 (N_15913,N_14471,N_14433);
nor U15914 (N_15914,N_14834,N_14435);
xor U15915 (N_15915,N_14038,N_14828);
or U15916 (N_15916,N_14020,N_14927);
nand U15917 (N_15917,N_14926,N_14501);
nor U15918 (N_15918,N_14383,N_14262);
or U15919 (N_15919,N_14212,N_14541);
xor U15920 (N_15920,N_14218,N_14418);
nor U15921 (N_15921,N_14071,N_14487);
nor U15922 (N_15922,N_14269,N_14915);
or U15923 (N_15923,N_14596,N_14592);
or U15924 (N_15924,N_14495,N_14128);
nand U15925 (N_15925,N_14454,N_14511);
xor U15926 (N_15926,N_14475,N_14546);
nor U15927 (N_15927,N_14417,N_14980);
nor U15928 (N_15928,N_14371,N_14854);
nor U15929 (N_15929,N_14024,N_14449);
nor U15930 (N_15930,N_14400,N_14088);
nor U15931 (N_15931,N_14181,N_14476);
and U15932 (N_15932,N_14115,N_14491);
or U15933 (N_15933,N_14701,N_14686);
nor U15934 (N_15934,N_14063,N_14593);
and U15935 (N_15935,N_14749,N_14286);
or U15936 (N_15936,N_14763,N_14262);
nand U15937 (N_15937,N_14712,N_14033);
xor U15938 (N_15938,N_14150,N_14834);
nor U15939 (N_15939,N_14953,N_14370);
xor U15940 (N_15940,N_14623,N_14890);
xor U15941 (N_15941,N_14852,N_14627);
or U15942 (N_15942,N_14057,N_14609);
and U15943 (N_15943,N_14721,N_14245);
nand U15944 (N_15944,N_14729,N_14555);
nor U15945 (N_15945,N_14988,N_14236);
and U15946 (N_15946,N_14387,N_14336);
or U15947 (N_15947,N_14884,N_14010);
xnor U15948 (N_15948,N_14593,N_14870);
and U15949 (N_15949,N_14385,N_14078);
and U15950 (N_15950,N_14960,N_14526);
nand U15951 (N_15951,N_14455,N_14818);
and U15952 (N_15952,N_14430,N_14153);
xnor U15953 (N_15953,N_14358,N_14524);
xor U15954 (N_15954,N_14824,N_14280);
nor U15955 (N_15955,N_14916,N_14693);
nor U15956 (N_15956,N_14357,N_14649);
nor U15957 (N_15957,N_14744,N_14476);
or U15958 (N_15958,N_14341,N_14350);
xor U15959 (N_15959,N_14136,N_14468);
or U15960 (N_15960,N_14684,N_14313);
nor U15961 (N_15961,N_14320,N_14413);
or U15962 (N_15962,N_14013,N_14114);
or U15963 (N_15963,N_14648,N_14135);
nor U15964 (N_15964,N_14313,N_14766);
or U15965 (N_15965,N_14917,N_14560);
or U15966 (N_15966,N_14232,N_14944);
xor U15967 (N_15967,N_14542,N_14402);
xor U15968 (N_15968,N_14257,N_14122);
nand U15969 (N_15969,N_14208,N_14888);
xnor U15970 (N_15970,N_14895,N_14846);
or U15971 (N_15971,N_14477,N_14165);
and U15972 (N_15972,N_14637,N_14224);
xnor U15973 (N_15973,N_14103,N_14701);
nor U15974 (N_15974,N_14238,N_14762);
nand U15975 (N_15975,N_14717,N_14007);
nor U15976 (N_15976,N_14693,N_14301);
nor U15977 (N_15977,N_14684,N_14718);
or U15978 (N_15978,N_14592,N_14262);
nor U15979 (N_15979,N_14516,N_14269);
nor U15980 (N_15980,N_14577,N_14909);
and U15981 (N_15981,N_14673,N_14498);
nand U15982 (N_15982,N_14452,N_14174);
nand U15983 (N_15983,N_14698,N_14857);
nor U15984 (N_15984,N_14051,N_14659);
and U15985 (N_15985,N_14113,N_14147);
xnor U15986 (N_15986,N_14835,N_14360);
nor U15987 (N_15987,N_14923,N_14191);
xor U15988 (N_15988,N_14917,N_14294);
nand U15989 (N_15989,N_14071,N_14587);
nand U15990 (N_15990,N_14792,N_14790);
nand U15991 (N_15991,N_14371,N_14197);
nor U15992 (N_15992,N_14785,N_14459);
nand U15993 (N_15993,N_14075,N_14261);
nor U15994 (N_15994,N_14313,N_14764);
nand U15995 (N_15995,N_14165,N_14091);
or U15996 (N_15996,N_14589,N_14392);
xnor U15997 (N_15997,N_14976,N_14296);
xnor U15998 (N_15998,N_14713,N_14216);
or U15999 (N_15999,N_14617,N_14553);
nor U16000 (N_16000,N_15750,N_15865);
xnor U16001 (N_16001,N_15243,N_15478);
xnor U16002 (N_16002,N_15950,N_15852);
and U16003 (N_16003,N_15521,N_15647);
nand U16004 (N_16004,N_15678,N_15605);
nand U16005 (N_16005,N_15897,N_15926);
nor U16006 (N_16006,N_15386,N_15325);
xnor U16007 (N_16007,N_15819,N_15525);
xnor U16008 (N_16008,N_15848,N_15223);
xnor U16009 (N_16009,N_15473,N_15481);
and U16010 (N_16010,N_15810,N_15145);
nor U16011 (N_16011,N_15299,N_15660);
and U16012 (N_16012,N_15611,N_15390);
and U16013 (N_16013,N_15416,N_15528);
xor U16014 (N_16014,N_15377,N_15707);
or U16015 (N_16015,N_15382,N_15796);
xor U16016 (N_16016,N_15064,N_15503);
nor U16017 (N_16017,N_15895,N_15373);
or U16018 (N_16018,N_15091,N_15984);
nor U16019 (N_16019,N_15332,N_15162);
nand U16020 (N_16020,N_15550,N_15081);
nand U16021 (N_16021,N_15639,N_15253);
and U16022 (N_16022,N_15094,N_15705);
nor U16023 (N_16023,N_15049,N_15055);
nand U16024 (N_16024,N_15847,N_15589);
nor U16025 (N_16025,N_15306,N_15463);
nand U16026 (N_16026,N_15420,N_15490);
nor U16027 (N_16027,N_15684,N_15524);
xnor U16028 (N_16028,N_15997,N_15493);
xnor U16029 (N_16029,N_15307,N_15009);
nor U16030 (N_16030,N_15472,N_15352);
and U16031 (N_16031,N_15188,N_15276);
nand U16032 (N_16032,N_15551,N_15393);
xor U16033 (N_16033,N_15242,N_15457);
nor U16034 (N_16034,N_15155,N_15185);
or U16035 (N_16035,N_15534,N_15830);
and U16036 (N_16036,N_15047,N_15782);
nor U16037 (N_16037,N_15902,N_15686);
nor U16038 (N_16038,N_15154,N_15728);
nor U16039 (N_16039,N_15281,N_15807);
or U16040 (N_16040,N_15339,N_15877);
xor U16041 (N_16041,N_15289,N_15908);
and U16042 (N_16042,N_15446,N_15288);
xnor U16043 (N_16043,N_15492,N_15506);
nor U16044 (N_16044,N_15685,N_15361);
xnor U16045 (N_16045,N_15236,N_15788);
xor U16046 (N_16046,N_15137,N_15957);
or U16047 (N_16047,N_15201,N_15709);
and U16048 (N_16048,N_15499,N_15884);
nor U16049 (N_16049,N_15056,N_15101);
or U16050 (N_16050,N_15290,N_15209);
nor U16051 (N_16051,N_15619,N_15026);
nor U16052 (N_16052,N_15922,N_15933);
nand U16053 (N_16053,N_15115,N_15072);
nand U16054 (N_16054,N_15644,N_15590);
or U16055 (N_16055,N_15418,N_15917);
nor U16056 (N_16056,N_15756,N_15649);
nor U16057 (N_16057,N_15417,N_15261);
nand U16058 (N_16058,N_15850,N_15641);
and U16059 (N_16059,N_15934,N_15718);
xnor U16060 (N_16060,N_15568,N_15683);
xnor U16061 (N_16061,N_15400,N_15855);
nor U16062 (N_16062,N_15798,N_15227);
or U16063 (N_16063,N_15766,N_15980);
xor U16064 (N_16064,N_15826,N_15286);
nor U16065 (N_16065,N_15458,N_15929);
nand U16066 (N_16066,N_15633,N_15015);
nand U16067 (N_16067,N_15392,N_15033);
nor U16068 (N_16068,N_15821,N_15962);
or U16069 (N_16069,N_15184,N_15772);
nand U16070 (N_16070,N_15229,N_15904);
nand U16071 (N_16071,N_15273,N_15967);
or U16072 (N_16072,N_15832,N_15448);
or U16073 (N_16073,N_15964,N_15876);
or U16074 (N_16074,N_15000,N_15177);
and U16075 (N_16075,N_15120,N_15182);
nor U16076 (N_16076,N_15424,N_15735);
xnor U16077 (N_16077,N_15058,N_15439);
and U16078 (N_16078,N_15447,N_15125);
or U16079 (N_16079,N_15511,N_15956);
nand U16080 (N_16080,N_15300,N_15747);
and U16081 (N_16081,N_15381,N_15912);
nand U16082 (N_16082,N_15618,N_15096);
xor U16083 (N_16083,N_15725,N_15313);
nor U16084 (N_16084,N_15498,N_15631);
or U16085 (N_16085,N_15349,N_15219);
xor U16086 (N_16086,N_15305,N_15779);
nand U16087 (N_16087,N_15794,N_15138);
and U16088 (N_16088,N_15991,N_15801);
and U16089 (N_16089,N_15333,N_15191);
or U16090 (N_16090,N_15742,N_15022);
and U16091 (N_16091,N_15336,N_15006);
nand U16092 (N_16092,N_15330,N_15398);
and U16093 (N_16093,N_15347,N_15932);
xnor U16094 (N_16094,N_15536,N_15052);
or U16095 (N_16095,N_15566,N_15475);
xnor U16096 (N_16096,N_15909,N_15806);
nor U16097 (N_16097,N_15749,N_15609);
or U16098 (N_16098,N_15573,N_15990);
xnor U16099 (N_16099,N_15411,N_15724);
and U16100 (N_16100,N_15993,N_15346);
or U16101 (N_16101,N_15438,N_15892);
nand U16102 (N_16102,N_15719,N_15245);
and U16103 (N_16103,N_15161,N_15041);
nand U16104 (N_16104,N_15319,N_15889);
or U16105 (N_16105,N_15051,N_15989);
or U16106 (N_16106,N_15940,N_15858);
and U16107 (N_16107,N_15190,N_15250);
nor U16108 (N_16108,N_15399,N_15602);
nand U16109 (N_16109,N_15743,N_15837);
nor U16110 (N_16110,N_15960,N_15773);
nor U16111 (N_16111,N_15264,N_15415);
or U16112 (N_16112,N_15112,N_15936);
and U16113 (N_16113,N_15547,N_15353);
xor U16114 (N_16114,N_15710,N_15959);
or U16115 (N_16115,N_15843,N_15700);
and U16116 (N_16116,N_15459,N_15105);
nand U16117 (N_16117,N_15217,N_15070);
nand U16118 (N_16118,N_15553,N_15999);
nor U16119 (N_16119,N_15218,N_15764);
xor U16120 (N_16120,N_15230,N_15966);
nor U16121 (N_16121,N_15340,N_15040);
nand U16122 (N_16122,N_15900,N_15642);
and U16123 (N_16123,N_15467,N_15513);
and U16124 (N_16124,N_15808,N_15523);
and U16125 (N_16125,N_15476,N_15401);
xor U16126 (N_16126,N_15938,N_15651);
and U16127 (N_16127,N_15696,N_15968);
xor U16128 (N_16128,N_15215,N_15180);
xor U16129 (N_16129,N_15574,N_15638);
or U16130 (N_16130,N_15714,N_15042);
and U16131 (N_16131,N_15898,N_15527);
xor U16132 (N_16132,N_15158,N_15387);
nor U16133 (N_16133,N_15531,N_15495);
nand U16134 (N_16134,N_15505,N_15578);
nor U16135 (N_16135,N_15862,N_15163);
and U16136 (N_16136,N_15488,N_15587);
nor U16137 (N_16137,N_15664,N_15486);
nand U16138 (N_16138,N_15159,N_15681);
xnor U16139 (N_16139,N_15376,N_15857);
and U16140 (N_16140,N_15269,N_15147);
nand U16141 (N_16141,N_15221,N_15903);
nor U16142 (N_16142,N_15024,N_15228);
nand U16143 (N_16143,N_15925,N_15485);
or U16144 (N_16144,N_15713,N_15791);
and U16145 (N_16145,N_15595,N_15767);
nor U16146 (N_16146,N_15383,N_15468);
xnor U16147 (N_16147,N_15045,N_15114);
nor U16148 (N_16148,N_15150,N_15635);
and U16149 (N_16149,N_15192,N_15890);
xor U16150 (N_16150,N_15133,N_15711);
or U16151 (N_16151,N_15835,N_15745);
nor U16152 (N_16152,N_15751,N_15414);
nand U16153 (N_16153,N_15057,N_15507);
and U16154 (N_16154,N_15315,N_15753);
xor U16155 (N_16155,N_15156,N_15872);
and U16156 (N_16156,N_15437,N_15792);
xor U16157 (N_16157,N_15804,N_15500);
and U16158 (N_16158,N_15755,N_15085);
nor U16159 (N_16159,N_15822,N_15126);
nand U16160 (N_16160,N_15691,N_15405);
and U16161 (N_16161,N_15617,N_15456);
xor U16162 (N_16162,N_15028,N_15128);
or U16163 (N_16163,N_15093,N_15246);
or U16164 (N_16164,N_15825,N_15483);
xor U16165 (N_16165,N_15206,N_15296);
and U16166 (N_16166,N_15443,N_15292);
nor U16167 (N_16167,N_15634,N_15918);
nand U16168 (N_16168,N_15734,N_15121);
nand U16169 (N_16169,N_15021,N_15196);
xnor U16170 (N_16170,N_15883,N_15484);
and U16171 (N_16171,N_15765,N_15001);
and U16172 (N_16172,N_15673,N_15576);
or U16173 (N_16173,N_15043,N_15628);
or U16174 (N_16174,N_15019,N_15391);
or U16175 (N_16175,N_15087,N_15202);
and U16176 (N_16176,N_15563,N_15099);
and U16177 (N_16177,N_15092,N_15477);
nor U16178 (N_16178,N_15915,N_15258);
xnor U16179 (N_16179,N_15280,N_15329);
or U16180 (N_16180,N_15863,N_15655);
nor U16181 (N_16181,N_15951,N_15777);
and U16182 (N_16182,N_15715,N_15232);
and U16183 (N_16183,N_15682,N_15135);
nand U16184 (N_16184,N_15435,N_15839);
or U16185 (N_16185,N_15981,N_15924);
or U16186 (N_16186,N_15856,N_15294);
xor U16187 (N_16187,N_15372,N_15688);
nor U16188 (N_16188,N_15178,N_15355);
or U16189 (N_16189,N_15032,N_15471);
nand U16190 (N_16190,N_15031,N_15901);
nand U16191 (N_16191,N_15899,N_15762);
and U16192 (N_16192,N_15455,N_15431);
nand U16193 (N_16193,N_15833,N_15529);
or U16194 (N_16194,N_15433,N_15518);
nor U16195 (N_16195,N_15680,N_15697);
nor U16196 (N_16196,N_15263,N_15712);
or U16197 (N_16197,N_15954,N_15259);
xnor U16198 (N_16198,N_15648,N_15846);
or U16199 (N_16199,N_15775,N_15367);
nor U16200 (N_16200,N_15348,N_15097);
or U16201 (N_16201,N_15010,N_15591);
xor U16202 (N_16202,N_15763,N_15036);
and U16203 (N_16203,N_15656,N_15271);
nor U16204 (N_16204,N_15975,N_15882);
nor U16205 (N_16205,N_15255,N_15017);
or U16206 (N_16206,N_15310,N_15131);
xor U16207 (N_16207,N_15733,N_15987);
xnor U16208 (N_16208,N_15816,N_15914);
or U16209 (N_16209,N_15632,N_15942);
nand U16210 (N_16210,N_15864,N_15759);
xor U16211 (N_16211,N_15295,N_15226);
nand U16212 (N_16212,N_15265,N_15474);
nand U16213 (N_16213,N_15974,N_15335);
and U16214 (N_16214,N_15434,N_15768);
nor U16215 (N_16215,N_15593,N_15197);
xor U16216 (N_16216,N_15564,N_15164);
and U16217 (N_16217,N_15103,N_15025);
xor U16218 (N_16218,N_15166,N_15893);
xor U16219 (N_16219,N_15314,N_15107);
nor U16220 (N_16220,N_15614,N_15887);
or U16221 (N_16221,N_15692,N_15110);
or U16222 (N_16222,N_15410,N_15778);
xor U16223 (N_16223,N_15020,N_15624);
nand U16224 (N_16224,N_15018,N_15504);
xor U16225 (N_16225,N_15879,N_15341);
or U16226 (N_16226,N_15216,N_15011);
xnor U16227 (N_16227,N_15034,N_15548);
xor U16228 (N_16228,N_15327,N_15667);
xor U16229 (N_16229,N_15854,N_15491);
nand U16230 (N_16230,N_15257,N_15181);
xnor U16231 (N_16231,N_15193,N_15913);
xor U16232 (N_16232,N_15211,N_15165);
xor U16233 (N_16233,N_15666,N_15570);
xor U16234 (N_16234,N_15996,N_15646);
xnor U16235 (N_16235,N_15213,N_15650);
and U16236 (N_16236,N_15630,N_15127);
nand U16237 (N_16237,N_15169,N_15144);
nor U16238 (N_16238,N_15172,N_15117);
nand U16239 (N_16239,N_15059,N_15986);
or U16240 (N_16240,N_15640,N_15874);
nor U16241 (N_16241,N_15428,N_15809);
nand U16242 (N_16242,N_15384,N_15780);
and U16243 (N_16243,N_15703,N_15971);
and U16244 (N_16244,N_15343,N_15911);
and U16245 (N_16245,N_15797,N_15061);
or U16246 (N_16246,N_15248,N_15291);
or U16247 (N_16247,N_15783,N_15748);
nand U16248 (N_16248,N_15077,N_15321);
and U16249 (N_16249,N_15254,N_15124);
nand U16250 (N_16250,N_15441,N_15425);
or U16251 (N_16251,N_15469,N_15198);
and U16252 (N_16252,N_15016,N_15316);
nand U16253 (N_16253,N_15298,N_15823);
and U16254 (N_16254,N_15979,N_15075);
nor U16255 (N_16255,N_15027,N_15878);
and U16256 (N_16256,N_15946,N_15311);
nand U16257 (N_16257,N_15937,N_15394);
or U16258 (N_16258,N_15413,N_15304);
or U16259 (N_16259,N_15442,N_15958);
and U16260 (N_16260,N_15342,N_15111);
or U16261 (N_16261,N_15881,N_15706);
nor U16262 (N_16262,N_15970,N_15931);
xor U16263 (N_16263,N_15616,N_15985);
or U16264 (N_16264,N_15338,N_15214);
or U16265 (N_16265,N_15921,N_15366);
and U16266 (N_16266,N_15123,N_15407);
xnor U16267 (N_16267,N_15482,N_15030);
nand U16268 (N_16268,N_15406,N_15351);
nor U16269 (N_16269,N_15039,N_15541);
nor U16270 (N_16270,N_15562,N_15168);
xnor U16271 (N_16271,N_15820,N_15556);
nand U16272 (N_16272,N_15008,N_15063);
nand U16273 (N_16273,N_15585,N_15580);
and U16274 (N_16274,N_15690,N_15653);
or U16275 (N_16275,N_15535,N_15194);
or U16276 (N_16276,N_15817,N_15995);
nand U16277 (N_16277,N_15761,N_15322);
xor U16278 (N_16278,N_15676,N_15982);
and U16279 (N_16279,N_15453,N_15544);
xor U16280 (N_16280,N_15861,N_15282);
nand U16281 (N_16281,N_15238,N_15873);
or U16282 (N_16282,N_15053,N_15770);
or U16283 (N_16283,N_15359,N_15251);
and U16284 (N_16284,N_15082,N_15470);
nor U16285 (N_16285,N_15663,N_15941);
nand U16286 (N_16286,N_15445,N_15203);
and U16287 (N_16287,N_15179,N_15757);
xor U16288 (N_16288,N_15905,N_15139);
xor U16289 (N_16289,N_15549,N_15466);
and U16290 (N_16290,N_15350,N_15429);
and U16291 (N_16291,N_15657,N_15831);
nor U16292 (N_16292,N_15244,N_15565);
xnor U16293 (N_16293,N_15037,N_15514);
nand U16294 (N_16294,N_15868,N_15601);
and U16295 (N_16295,N_15012,N_15038);
and U16296 (N_16296,N_15814,N_15677);
xnor U16297 (N_16297,N_15939,N_15005);
and U16298 (N_16298,N_15241,N_15395);
nand U16299 (N_16299,N_15774,N_15388);
xnor U16300 (N_16300,N_15795,N_15919);
nor U16301 (N_16301,N_15317,N_15326);
xor U16302 (N_16302,N_15818,N_15113);
and U16303 (N_16303,N_15187,N_15787);
xnor U16304 (N_16304,N_15916,N_15369);
nor U16305 (N_16305,N_15119,N_15068);
nand U16306 (N_16306,N_15205,N_15284);
nand U16307 (N_16307,N_15859,N_15622);
xnor U16308 (N_16308,N_15983,N_15247);
nand U16309 (N_16309,N_15594,N_15771);
nand U16310 (N_16310,N_15277,N_15427);
xnor U16311 (N_16311,N_15278,N_15436);
and U16312 (N_16312,N_15212,N_15907);
or U16313 (N_16313,N_15270,N_15220);
nand U16314 (N_16314,N_15567,N_15645);
or U16315 (N_16315,N_15378,N_15397);
or U16316 (N_16316,N_15303,N_15841);
nor U16317 (N_16317,N_15621,N_15698);
and U16318 (N_16318,N_15404,N_15331);
or U16319 (N_16319,N_15952,N_15323);
nand U16320 (N_16320,N_15722,N_15363);
or U16321 (N_16321,N_15084,N_15575);
nand U16322 (N_16322,N_15130,N_15606);
or U16323 (N_16323,N_15994,N_15955);
xor U16324 (N_16324,N_15176,N_15256);
or U16325 (N_16325,N_15360,N_15412);
xor U16326 (N_16326,N_15204,N_15963);
or U16327 (N_16327,N_15146,N_15149);
xnor U16328 (N_16328,N_15231,N_15118);
or U16329 (N_16329,N_15610,N_15658);
xnor U16330 (N_16330,N_15561,N_15554);
nor U16331 (N_16331,N_15953,N_15625);
or U16332 (N_16332,N_15972,N_15167);
nor U16333 (N_16333,N_15208,N_15786);
xnor U16334 (N_16334,N_15636,N_15785);
or U16335 (N_16335,N_15389,N_15210);
nor U16336 (N_16336,N_15637,N_15572);
or U16337 (N_16337,N_15744,N_15927);
or U16338 (N_16338,N_15007,N_15569);
nand U16339 (N_16339,N_15935,N_15626);
nor U16340 (N_16340,N_15334,N_15324);
nor U16341 (N_16341,N_15409,N_15449);
nand U16342 (N_16342,N_15522,N_15344);
nand U16343 (N_16343,N_15888,N_15370);
xnor U16344 (N_16344,N_15802,N_15860);
nor U16345 (N_16345,N_15662,N_15444);
and U16346 (N_16346,N_15558,N_15252);
xnor U16347 (N_16347,N_15815,N_15354);
and U16348 (N_16348,N_15297,N_15838);
or U16349 (N_16349,N_15702,N_15048);
nor U16350 (N_16350,N_15828,N_15827);
or U16351 (N_16351,N_15704,N_15803);
nand U16352 (N_16352,N_15517,N_15516);
nand U16353 (N_16353,N_15152,N_15740);
or U16354 (N_16354,N_15419,N_15533);
xnor U16355 (N_16355,N_15992,N_15600);
and U16356 (N_16356,N_15375,N_15539);
nand U16357 (N_16357,N_15422,N_15003);
xnor U16358 (N_16358,N_15875,N_15089);
nand U16359 (N_16359,N_15845,N_15362);
or U16360 (N_16360,N_15451,N_15699);
nand U16361 (N_16361,N_15612,N_15423);
and U16362 (N_16362,N_15496,N_15896);
nor U16363 (N_16363,N_15440,N_15701);
nor U16364 (N_16364,N_15054,N_15141);
or U16365 (N_16365,N_15060,N_15538);
nand U16366 (N_16366,N_15674,N_15170);
nand U16367 (N_16367,N_15973,N_15171);
and U16368 (N_16368,N_15100,N_15153);
nor U16369 (N_16369,N_15080,N_15174);
or U16370 (N_16370,N_15928,N_15268);
or U16371 (N_16371,N_15450,N_15186);
or U16372 (N_16372,N_15301,N_15739);
nand U16373 (N_16373,N_15623,N_15283);
or U16374 (N_16374,N_15643,N_15867);
nor U16375 (N_16375,N_15894,N_15559);
xnor U16376 (N_16376,N_15824,N_15998);
and U16377 (N_16377,N_15368,N_15721);
xor U16378 (N_16378,N_15235,N_15526);
nor U16379 (N_16379,N_15930,N_15988);
or U16380 (N_16380,N_15560,N_15949);
and U16381 (N_16381,N_15035,N_15509);
or U16382 (N_16382,N_15737,N_15224);
nand U16383 (N_16383,N_15597,N_15813);
xnor U16384 (N_16384,N_15195,N_15104);
nand U16385 (N_16385,N_15122,N_15279);
xor U16386 (N_16386,N_15151,N_15920);
or U16387 (N_16387,N_15604,N_15479);
or U16388 (N_16388,N_15659,N_15044);
or U16389 (N_16389,N_15769,N_15784);
or U16390 (N_16390,N_15046,N_15754);
and U16391 (N_16391,N_15976,N_15866);
nand U16392 (N_16392,N_15542,N_15840);
nor U16393 (N_16393,N_15800,N_15066);
nor U16394 (N_16394,N_15947,N_15462);
and U16395 (N_16395,N_15002,N_15309);
and U16396 (N_16396,N_15134,N_15615);
nand U16397 (N_16397,N_15098,N_15870);
xor U16398 (N_16398,N_15736,N_15487);
nor U16399 (N_16399,N_15379,N_15079);
or U16400 (N_16400,N_15727,N_15083);
or U16401 (N_16401,N_15760,N_15207);
nor U16402 (N_16402,N_15004,N_15708);
nor U16403 (N_16403,N_15374,N_15078);
or U16404 (N_16404,N_15851,N_15948);
nor U16405 (N_16405,N_15222,N_15789);
nand U16406 (N_16406,N_15106,N_15189);
nor U16407 (N_16407,N_15603,N_15586);
and U16408 (N_16408,N_15050,N_15013);
xor U16409 (N_16409,N_15944,N_15074);
nand U16410 (N_16410,N_15726,N_15853);
nor U16411 (N_16411,N_15588,N_15086);
nor U16412 (N_16412,N_15140,N_15287);
nand U16413 (N_16413,N_15421,N_15834);
nor U16414 (N_16414,N_15654,N_15582);
xor U16415 (N_16415,N_15285,N_15512);
and U16416 (N_16416,N_15460,N_15687);
and U16417 (N_16417,N_15129,N_15571);
and U16418 (N_16418,N_15272,N_15365);
nor U16419 (N_16419,N_15842,N_15508);
and U16420 (N_16420,N_15665,N_15869);
and U16421 (N_16421,N_15579,N_15260);
xor U16422 (N_16422,N_15545,N_15746);
xnor U16423 (N_16423,N_15577,N_15670);
nor U16424 (N_16424,N_15175,N_15396);
xnor U16425 (N_16425,N_15065,N_15200);
and U16426 (N_16426,N_15607,N_15694);
nor U16427 (N_16427,N_15454,N_15108);
xor U16428 (N_16428,N_15720,N_15627);
nand U16429 (N_16429,N_15402,N_15109);
nor U16430 (N_16430,N_15318,N_15675);
nor U16431 (N_16431,N_15225,N_15965);
or U16432 (N_16432,N_15520,N_15143);
nand U16433 (N_16433,N_15717,N_15584);
and U16434 (N_16434,N_15275,N_15961);
or U16435 (N_16435,N_15132,N_15844);
nor U16436 (N_16436,N_15608,N_15738);
nand U16437 (N_16437,N_15886,N_15945);
xor U16438 (N_16438,N_15943,N_15308);
and U16439 (N_16439,N_15519,N_15599);
nor U16440 (N_16440,N_15502,N_15811);
or U16441 (N_16441,N_15237,N_15157);
nand U16442 (N_16442,N_15652,N_15546);
or U16443 (N_16443,N_15752,N_15978);
nor U16444 (N_16444,N_15581,N_15661);
nor U16445 (N_16445,N_15408,N_15532);
xor U16446 (N_16446,N_15358,N_15328);
or U16447 (N_16447,N_15812,N_15076);
or U16448 (N_16448,N_15380,N_15781);
nor U16449 (N_16449,N_15183,N_15793);
nand U16450 (N_16450,N_15403,N_15302);
nand U16451 (N_16451,N_15239,N_15062);
xnor U16452 (N_16452,N_15758,N_15977);
nor U16453 (N_16453,N_15148,N_15530);
nor U16454 (N_16454,N_15116,N_15267);
or U16455 (N_16455,N_15432,N_15262);
nand U16456 (N_16456,N_15356,N_15014);
nand U16457 (N_16457,N_15836,N_15693);
and U16458 (N_16458,N_15629,N_15452);
nand U16459 (N_16459,N_15266,N_15880);
nand U16460 (N_16460,N_15088,N_15293);
or U16461 (N_16461,N_15776,N_15029);
nand U16462 (N_16462,N_15073,N_15312);
nand U16463 (N_16463,N_15805,N_15969);
xor U16464 (N_16464,N_15849,N_15464);
xor U16465 (N_16465,N_15199,N_15501);
nand U16466 (N_16466,N_15515,N_15669);
nor U16467 (N_16467,N_15552,N_15337);
or U16468 (N_16468,N_15385,N_15741);
xnor U16469 (N_16469,N_15480,N_15136);
nor U16470 (N_16470,N_15557,N_15071);
or U16471 (N_16471,N_15672,N_15142);
and U16472 (N_16472,N_15274,N_15465);
nor U16473 (N_16473,N_15489,N_15731);
nor U16474 (N_16474,N_15497,N_15730);
xnor U16475 (N_16475,N_15923,N_15689);
and U16476 (N_16476,N_15829,N_15371);
or U16477 (N_16477,N_15537,N_15430);
and U16478 (N_16478,N_15364,N_15716);
nand U16479 (N_16479,N_15906,N_15885);
and U16480 (N_16480,N_15668,N_15679);
nor U16481 (N_16481,N_15357,N_15160);
or U16482 (N_16482,N_15426,N_15598);
and U16483 (N_16483,N_15732,N_15173);
nor U16484 (N_16484,N_15596,N_15320);
xnor U16485 (N_16485,N_15102,N_15799);
and U16486 (N_16486,N_15067,N_15345);
or U16487 (N_16487,N_15729,N_15090);
nand U16488 (N_16488,N_15790,N_15540);
nand U16489 (N_16489,N_15069,N_15910);
xor U16490 (N_16490,N_15671,N_15494);
nor U16491 (N_16491,N_15510,N_15240);
and U16492 (N_16492,N_15891,N_15583);
xnor U16493 (N_16493,N_15695,N_15592);
or U16494 (N_16494,N_15613,N_15023);
nand U16495 (N_16495,N_15233,N_15249);
or U16496 (N_16496,N_15871,N_15095);
and U16497 (N_16497,N_15555,N_15234);
and U16498 (N_16498,N_15620,N_15543);
and U16499 (N_16499,N_15461,N_15723);
and U16500 (N_16500,N_15942,N_15937);
nor U16501 (N_16501,N_15804,N_15376);
xor U16502 (N_16502,N_15940,N_15272);
nor U16503 (N_16503,N_15431,N_15619);
or U16504 (N_16504,N_15144,N_15652);
nand U16505 (N_16505,N_15337,N_15708);
and U16506 (N_16506,N_15272,N_15454);
and U16507 (N_16507,N_15735,N_15581);
xnor U16508 (N_16508,N_15645,N_15162);
or U16509 (N_16509,N_15682,N_15756);
xnor U16510 (N_16510,N_15489,N_15282);
or U16511 (N_16511,N_15211,N_15000);
nor U16512 (N_16512,N_15864,N_15919);
nand U16513 (N_16513,N_15398,N_15391);
nand U16514 (N_16514,N_15983,N_15127);
nand U16515 (N_16515,N_15427,N_15301);
xnor U16516 (N_16516,N_15341,N_15469);
nand U16517 (N_16517,N_15053,N_15124);
nor U16518 (N_16518,N_15857,N_15811);
xor U16519 (N_16519,N_15085,N_15414);
nor U16520 (N_16520,N_15653,N_15285);
xnor U16521 (N_16521,N_15820,N_15562);
nand U16522 (N_16522,N_15574,N_15509);
xnor U16523 (N_16523,N_15120,N_15341);
nor U16524 (N_16524,N_15702,N_15370);
nand U16525 (N_16525,N_15451,N_15452);
nand U16526 (N_16526,N_15590,N_15771);
or U16527 (N_16527,N_15805,N_15387);
and U16528 (N_16528,N_15875,N_15463);
nor U16529 (N_16529,N_15130,N_15280);
xor U16530 (N_16530,N_15929,N_15916);
or U16531 (N_16531,N_15950,N_15608);
or U16532 (N_16532,N_15932,N_15793);
and U16533 (N_16533,N_15427,N_15663);
xor U16534 (N_16534,N_15214,N_15989);
nand U16535 (N_16535,N_15677,N_15461);
xnor U16536 (N_16536,N_15462,N_15340);
and U16537 (N_16537,N_15017,N_15549);
nand U16538 (N_16538,N_15393,N_15818);
nand U16539 (N_16539,N_15111,N_15244);
and U16540 (N_16540,N_15982,N_15204);
nor U16541 (N_16541,N_15860,N_15286);
nand U16542 (N_16542,N_15598,N_15876);
and U16543 (N_16543,N_15229,N_15965);
nor U16544 (N_16544,N_15918,N_15258);
xor U16545 (N_16545,N_15850,N_15216);
nand U16546 (N_16546,N_15852,N_15519);
and U16547 (N_16547,N_15757,N_15237);
nand U16548 (N_16548,N_15373,N_15449);
xnor U16549 (N_16549,N_15814,N_15605);
xor U16550 (N_16550,N_15770,N_15967);
or U16551 (N_16551,N_15746,N_15851);
or U16552 (N_16552,N_15834,N_15052);
xor U16553 (N_16553,N_15098,N_15460);
and U16554 (N_16554,N_15749,N_15255);
nor U16555 (N_16555,N_15173,N_15607);
and U16556 (N_16556,N_15529,N_15625);
xnor U16557 (N_16557,N_15583,N_15910);
and U16558 (N_16558,N_15672,N_15466);
xor U16559 (N_16559,N_15205,N_15131);
and U16560 (N_16560,N_15540,N_15499);
xnor U16561 (N_16561,N_15558,N_15388);
nand U16562 (N_16562,N_15919,N_15118);
or U16563 (N_16563,N_15669,N_15363);
and U16564 (N_16564,N_15915,N_15450);
nor U16565 (N_16565,N_15890,N_15119);
xor U16566 (N_16566,N_15071,N_15188);
or U16567 (N_16567,N_15310,N_15740);
nand U16568 (N_16568,N_15807,N_15176);
or U16569 (N_16569,N_15916,N_15747);
or U16570 (N_16570,N_15089,N_15171);
and U16571 (N_16571,N_15522,N_15529);
xnor U16572 (N_16572,N_15142,N_15483);
and U16573 (N_16573,N_15897,N_15345);
or U16574 (N_16574,N_15134,N_15942);
xnor U16575 (N_16575,N_15455,N_15895);
or U16576 (N_16576,N_15481,N_15332);
nor U16577 (N_16577,N_15705,N_15602);
and U16578 (N_16578,N_15276,N_15555);
xnor U16579 (N_16579,N_15522,N_15361);
nand U16580 (N_16580,N_15150,N_15816);
or U16581 (N_16581,N_15865,N_15615);
or U16582 (N_16582,N_15754,N_15816);
nand U16583 (N_16583,N_15170,N_15655);
or U16584 (N_16584,N_15719,N_15945);
nand U16585 (N_16585,N_15536,N_15288);
or U16586 (N_16586,N_15602,N_15335);
nand U16587 (N_16587,N_15746,N_15733);
xor U16588 (N_16588,N_15991,N_15296);
or U16589 (N_16589,N_15154,N_15185);
nor U16590 (N_16590,N_15188,N_15954);
xnor U16591 (N_16591,N_15587,N_15578);
nor U16592 (N_16592,N_15108,N_15085);
nand U16593 (N_16593,N_15849,N_15670);
nor U16594 (N_16594,N_15913,N_15313);
and U16595 (N_16595,N_15211,N_15905);
and U16596 (N_16596,N_15588,N_15525);
nand U16597 (N_16597,N_15146,N_15242);
nand U16598 (N_16598,N_15647,N_15473);
nand U16599 (N_16599,N_15577,N_15744);
xnor U16600 (N_16600,N_15294,N_15439);
and U16601 (N_16601,N_15650,N_15046);
and U16602 (N_16602,N_15990,N_15110);
or U16603 (N_16603,N_15030,N_15014);
xor U16604 (N_16604,N_15199,N_15884);
and U16605 (N_16605,N_15135,N_15765);
nor U16606 (N_16606,N_15583,N_15920);
nor U16607 (N_16607,N_15659,N_15984);
xor U16608 (N_16608,N_15945,N_15152);
nand U16609 (N_16609,N_15111,N_15291);
or U16610 (N_16610,N_15502,N_15829);
or U16611 (N_16611,N_15923,N_15291);
and U16612 (N_16612,N_15886,N_15649);
xor U16613 (N_16613,N_15034,N_15057);
or U16614 (N_16614,N_15777,N_15445);
nand U16615 (N_16615,N_15244,N_15955);
xnor U16616 (N_16616,N_15389,N_15496);
or U16617 (N_16617,N_15885,N_15099);
xor U16618 (N_16618,N_15408,N_15883);
xnor U16619 (N_16619,N_15686,N_15270);
nor U16620 (N_16620,N_15927,N_15502);
nand U16621 (N_16621,N_15332,N_15516);
nor U16622 (N_16622,N_15558,N_15387);
nand U16623 (N_16623,N_15219,N_15802);
nand U16624 (N_16624,N_15056,N_15599);
or U16625 (N_16625,N_15247,N_15356);
nand U16626 (N_16626,N_15302,N_15158);
nor U16627 (N_16627,N_15617,N_15417);
nand U16628 (N_16628,N_15739,N_15073);
nor U16629 (N_16629,N_15662,N_15086);
nand U16630 (N_16630,N_15731,N_15164);
xor U16631 (N_16631,N_15134,N_15466);
and U16632 (N_16632,N_15386,N_15309);
nand U16633 (N_16633,N_15231,N_15078);
nand U16634 (N_16634,N_15050,N_15291);
nor U16635 (N_16635,N_15522,N_15887);
or U16636 (N_16636,N_15807,N_15566);
or U16637 (N_16637,N_15976,N_15679);
xor U16638 (N_16638,N_15512,N_15982);
nor U16639 (N_16639,N_15657,N_15817);
xor U16640 (N_16640,N_15240,N_15768);
nor U16641 (N_16641,N_15874,N_15524);
and U16642 (N_16642,N_15509,N_15263);
xor U16643 (N_16643,N_15751,N_15818);
or U16644 (N_16644,N_15724,N_15407);
nand U16645 (N_16645,N_15559,N_15040);
nor U16646 (N_16646,N_15559,N_15214);
xnor U16647 (N_16647,N_15481,N_15355);
nor U16648 (N_16648,N_15514,N_15342);
nand U16649 (N_16649,N_15575,N_15975);
and U16650 (N_16650,N_15843,N_15905);
nor U16651 (N_16651,N_15781,N_15536);
or U16652 (N_16652,N_15694,N_15381);
xor U16653 (N_16653,N_15564,N_15090);
xnor U16654 (N_16654,N_15636,N_15144);
or U16655 (N_16655,N_15734,N_15275);
nand U16656 (N_16656,N_15477,N_15882);
nand U16657 (N_16657,N_15301,N_15116);
or U16658 (N_16658,N_15940,N_15664);
and U16659 (N_16659,N_15118,N_15962);
and U16660 (N_16660,N_15687,N_15413);
xnor U16661 (N_16661,N_15989,N_15918);
nor U16662 (N_16662,N_15777,N_15995);
nand U16663 (N_16663,N_15738,N_15378);
nand U16664 (N_16664,N_15872,N_15884);
and U16665 (N_16665,N_15821,N_15124);
or U16666 (N_16666,N_15468,N_15845);
nor U16667 (N_16667,N_15065,N_15539);
nor U16668 (N_16668,N_15680,N_15113);
and U16669 (N_16669,N_15841,N_15211);
and U16670 (N_16670,N_15971,N_15473);
nor U16671 (N_16671,N_15204,N_15039);
nand U16672 (N_16672,N_15687,N_15929);
nor U16673 (N_16673,N_15424,N_15052);
nand U16674 (N_16674,N_15964,N_15385);
xnor U16675 (N_16675,N_15273,N_15880);
nand U16676 (N_16676,N_15484,N_15392);
or U16677 (N_16677,N_15107,N_15973);
and U16678 (N_16678,N_15940,N_15951);
xor U16679 (N_16679,N_15763,N_15068);
nor U16680 (N_16680,N_15782,N_15340);
and U16681 (N_16681,N_15031,N_15106);
and U16682 (N_16682,N_15381,N_15553);
xor U16683 (N_16683,N_15345,N_15390);
and U16684 (N_16684,N_15434,N_15247);
or U16685 (N_16685,N_15122,N_15641);
and U16686 (N_16686,N_15825,N_15591);
and U16687 (N_16687,N_15960,N_15573);
and U16688 (N_16688,N_15763,N_15477);
or U16689 (N_16689,N_15300,N_15140);
and U16690 (N_16690,N_15259,N_15850);
xor U16691 (N_16691,N_15365,N_15226);
nor U16692 (N_16692,N_15684,N_15902);
nor U16693 (N_16693,N_15955,N_15641);
nor U16694 (N_16694,N_15888,N_15671);
nand U16695 (N_16695,N_15207,N_15183);
and U16696 (N_16696,N_15767,N_15768);
and U16697 (N_16697,N_15752,N_15561);
nor U16698 (N_16698,N_15451,N_15549);
nor U16699 (N_16699,N_15817,N_15457);
and U16700 (N_16700,N_15106,N_15774);
nor U16701 (N_16701,N_15123,N_15881);
and U16702 (N_16702,N_15742,N_15347);
xnor U16703 (N_16703,N_15934,N_15782);
nor U16704 (N_16704,N_15450,N_15249);
xor U16705 (N_16705,N_15860,N_15477);
or U16706 (N_16706,N_15053,N_15409);
xnor U16707 (N_16707,N_15708,N_15650);
or U16708 (N_16708,N_15687,N_15948);
and U16709 (N_16709,N_15209,N_15624);
or U16710 (N_16710,N_15602,N_15242);
and U16711 (N_16711,N_15505,N_15616);
nand U16712 (N_16712,N_15101,N_15560);
nand U16713 (N_16713,N_15440,N_15398);
nor U16714 (N_16714,N_15471,N_15687);
nand U16715 (N_16715,N_15151,N_15694);
nand U16716 (N_16716,N_15485,N_15356);
nor U16717 (N_16717,N_15598,N_15798);
nand U16718 (N_16718,N_15320,N_15217);
nor U16719 (N_16719,N_15771,N_15469);
nor U16720 (N_16720,N_15570,N_15931);
nor U16721 (N_16721,N_15080,N_15796);
or U16722 (N_16722,N_15361,N_15487);
nand U16723 (N_16723,N_15899,N_15181);
xor U16724 (N_16724,N_15750,N_15063);
nand U16725 (N_16725,N_15058,N_15491);
nand U16726 (N_16726,N_15892,N_15217);
xnor U16727 (N_16727,N_15441,N_15107);
nor U16728 (N_16728,N_15865,N_15029);
nand U16729 (N_16729,N_15839,N_15888);
or U16730 (N_16730,N_15164,N_15949);
or U16731 (N_16731,N_15314,N_15516);
nor U16732 (N_16732,N_15544,N_15993);
nor U16733 (N_16733,N_15923,N_15510);
nand U16734 (N_16734,N_15419,N_15976);
nor U16735 (N_16735,N_15816,N_15373);
nor U16736 (N_16736,N_15957,N_15557);
and U16737 (N_16737,N_15028,N_15377);
xnor U16738 (N_16738,N_15601,N_15086);
xor U16739 (N_16739,N_15628,N_15888);
nor U16740 (N_16740,N_15144,N_15429);
and U16741 (N_16741,N_15756,N_15033);
nand U16742 (N_16742,N_15970,N_15167);
and U16743 (N_16743,N_15401,N_15995);
nor U16744 (N_16744,N_15252,N_15853);
xnor U16745 (N_16745,N_15352,N_15773);
or U16746 (N_16746,N_15258,N_15870);
and U16747 (N_16747,N_15398,N_15061);
nor U16748 (N_16748,N_15287,N_15507);
and U16749 (N_16749,N_15818,N_15870);
xor U16750 (N_16750,N_15892,N_15219);
nor U16751 (N_16751,N_15867,N_15411);
nand U16752 (N_16752,N_15960,N_15471);
xor U16753 (N_16753,N_15773,N_15937);
and U16754 (N_16754,N_15340,N_15564);
and U16755 (N_16755,N_15207,N_15659);
nor U16756 (N_16756,N_15890,N_15735);
xor U16757 (N_16757,N_15972,N_15274);
or U16758 (N_16758,N_15300,N_15310);
nor U16759 (N_16759,N_15814,N_15738);
nand U16760 (N_16760,N_15970,N_15756);
xnor U16761 (N_16761,N_15663,N_15724);
or U16762 (N_16762,N_15670,N_15279);
xnor U16763 (N_16763,N_15100,N_15119);
or U16764 (N_16764,N_15924,N_15237);
and U16765 (N_16765,N_15446,N_15296);
or U16766 (N_16766,N_15962,N_15237);
xor U16767 (N_16767,N_15903,N_15948);
or U16768 (N_16768,N_15596,N_15739);
nor U16769 (N_16769,N_15094,N_15837);
nand U16770 (N_16770,N_15593,N_15130);
xor U16771 (N_16771,N_15591,N_15680);
xor U16772 (N_16772,N_15055,N_15413);
xnor U16773 (N_16773,N_15486,N_15654);
nor U16774 (N_16774,N_15932,N_15917);
nor U16775 (N_16775,N_15786,N_15713);
nor U16776 (N_16776,N_15881,N_15842);
nor U16777 (N_16777,N_15423,N_15203);
nor U16778 (N_16778,N_15382,N_15053);
or U16779 (N_16779,N_15657,N_15616);
or U16780 (N_16780,N_15120,N_15574);
nor U16781 (N_16781,N_15873,N_15272);
or U16782 (N_16782,N_15749,N_15820);
nor U16783 (N_16783,N_15126,N_15250);
or U16784 (N_16784,N_15457,N_15839);
xor U16785 (N_16785,N_15675,N_15788);
and U16786 (N_16786,N_15074,N_15546);
and U16787 (N_16787,N_15478,N_15282);
and U16788 (N_16788,N_15495,N_15955);
nor U16789 (N_16789,N_15005,N_15511);
nor U16790 (N_16790,N_15881,N_15527);
and U16791 (N_16791,N_15030,N_15937);
and U16792 (N_16792,N_15387,N_15959);
nand U16793 (N_16793,N_15844,N_15368);
nand U16794 (N_16794,N_15594,N_15322);
or U16795 (N_16795,N_15828,N_15888);
or U16796 (N_16796,N_15384,N_15155);
nand U16797 (N_16797,N_15553,N_15874);
xnor U16798 (N_16798,N_15133,N_15152);
nor U16799 (N_16799,N_15891,N_15705);
nor U16800 (N_16800,N_15673,N_15335);
or U16801 (N_16801,N_15301,N_15944);
and U16802 (N_16802,N_15959,N_15369);
nor U16803 (N_16803,N_15573,N_15941);
nor U16804 (N_16804,N_15273,N_15475);
xor U16805 (N_16805,N_15684,N_15512);
or U16806 (N_16806,N_15917,N_15020);
or U16807 (N_16807,N_15115,N_15620);
or U16808 (N_16808,N_15195,N_15759);
nand U16809 (N_16809,N_15651,N_15762);
nand U16810 (N_16810,N_15245,N_15671);
xnor U16811 (N_16811,N_15579,N_15315);
nand U16812 (N_16812,N_15883,N_15301);
xnor U16813 (N_16813,N_15591,N_15585);
nor U16814 (N_16814,N_15414,N_15493);
or U16815 (N_16815,N_15076,N_15134);
nor U16816 (N_16816,N_15559,N_15036);
xnor U16817 (N_16817,N_15659,N_15774);
nand U16818 (N_16818,N_15200,N_15730);
and U16819 (N_16819,N_15412,N_15399);
and U16820 (N_16820,N_15121,N_15615);
nor U16821 (N_16821,N_15508,N_15802);
nor U16822 (N_16822,N_15158,N_15726);
xor U16823 (N_16823,N_15692,N_15563);
and U16824 (N_16824,N_15507,N_15958);
xnor U16825 (N_16825,N_15542,N_15475);
xnor U16826 (N_16826,N_15055,N_15734);
xor U16827 (N_16827,N_15265,N_15828);
nor U16828 (N_16828,N_15430,N_15077);
nand U16829 (N_16829,N_15782,N_15372);
and U16830 (N_16830,N_15159,N_15994);
and U16831 (N_16831,N_15035,N_15991);
xnor U16832 (N_16832,N_15810,N_15640);
and U16833 (N_16833,N_15767,N_15020);
nor U16834 (N_16834,N_15328,N_15149);
xnor U16835 (N_16835,N_15775,N_15267);
nor U16836 (N_16836,N_15335,N_15145);
nand U16837 (N_16837,N_15558,N_15428);
and U16838 (N_16838,N_15144,N_15452);
nand U16839 (N_16839,N_15045,N_15205);
or U16840 (N_16840,N_15486,N_15546);
nand U16841 (N_16841,N_15654,N_15595);
nor U16842 (N_16842,N_15636,N_15589);
nand U16843 (N_16843,N_15961,N_15324);
nor U16844 (N_16844,N_15566,N_15789);
nand U16845 (N_16845,N_15956,N_15054);
or U16846 (N_16846,N_15639,N_15996);
or U16847 (N_16847,N_15279,N_15254);
nor U16848 (N_16848,N_15420,N_15556);
nor U16849 (N_16849,N_15836,N_15309);
and U16850 (N_16850,N_15466,N_15145);
xor U16851 (N_16851,N_15953,N_15818);
nand U16852 (N_16852,N_15938,N_15206);
xnor U16853 (N_16853,N_15935,N_15753);
and U16854 (N_16854,N_15426,N_15865);
nor U16855 (N_16855,N_15660,N_15460);
and U16856 (N_16856,N_15790,N_15282);
and U16857 (N_16857,N_15605,N_15303);
nand U16858 (N_16858,N_15040,N_15373);
or U16859 (N_16859,N_15337,N_15525);
nor U16860 (N_16860,N_15246,N_15747);
xor U16861 (N_16861,N_15456,N_15717);
and U16862 (N_16862,N_15039,N_15623);
xor U16863 (N_16863,N_15193,N_15745);
xnor U16864 (N_16864,N_15471,N_15484);
and U16865 (N_16865,N_15876,N_15033);
xnor U16866 (N_16866,N_15546,N_15713);
xor U16867 (N_16867,N_15238,N_15700);
or U16868 (N_16868,N_15685,N_15294);
and U16869 (N_16869,N_15965,N_15660);
xor U16870 (N_16870,N_15037,N_15945);
nand U16871 (N_16871,N_15966,N_15341);
nor U16872 (N_16872,N_15955,N_15150);
or U16873 (N_16873,N_15173,N_15325);
xnor U16874 (N_16874,N_15381,N_15215);
nand U16875 (N_16875,N_15538,N_15830);
and U16876 (N_16876,N_15720,N_15076);
nand U16877 (N_16877,N_15012,N_15644);
or U16878 (N_16878,N_15290,N_15538);
xnor U16879 (N_16879,N_15250,N_15617);
or U16880 (N_16880,N_15328,N_15771);
nor U16881 (N_16881,N_15334,N_15435);
nor U16882 (N_16882,N_15952,N_15594);
or U16883 (N_16883,N_15748,N_15143);
or U16884 (N_16884,N_15901,N_15693);
nand U16885 (N_16885,N_15064,N_15621);
xor U16886 (N_16886,N_15631,N_15241);
nand U16887 (N_16887,N_15487,N_15260);
xnor U16888 (N_16888,N_15372,N_15972);
nand U16889 (N_16889,N_15206,N_15157);
or U16890 (N_16890,N_15921,N_15874);
xnor U16891 (N_16891,N_15758,N_15248);
or U16892 (N_16892,N_15411,N_15273);
xor U16893 (N_16893,N_15254,N_15657);
nor U16894 (N_16894,N_15718,N_15841);
xnor U16895 (N_16895,N_15558,N_15507);
nor U16896 (N_16896,N_15369,N_15331);
nor U16897 (N_16897,N_15458,N_15984);
or U16898 (N_16898,N_15825,N_15785);
xnor U16899 (N_16899,N_15030,N_15187);
nand U16900 (N_16900,N_15925,N_15806);
and U16901 (N_16901,N_15978,N_15646);
nor U16902 (N_16902,N_15077,N_15510);
or U16903 (N_16903,N_15061,N_15916);
nand U16904 (N_16904,N_15668,N_15568);
nand U16905 (N_16905,N_15960,N_15026);
xor U16906 (N_16906,N_15165,N_15408);
and U16907 (N_16907,N_15914,N_15639);
nand U16908 (N_16908,N_15115,N_15205);
or U16909 (N_16909,N_15954,N_15341);
nor U16910 (N_16910,N_15317,N_15761);
or U16911 (N_16911,N_15135,N_15197);
or U16912 (N_16912,N_15470,N_15269);
nor U16913 (N_16913,N_15991,N_15470);
and U16914 (N_16914,N_15774,N_15551);
nor U16915 (N_16915,N_15066,N_15289);
or U16916 (N_16916,N_15427,N_15751);
nand U16917 (N_16917,N_15019,N_15396);
or U16918 (N_16918,N_15242,N_15254);
nor U16919 (N_16919,N_15195,N_15689);
nor U16920 (N_16920,N_15522,N_15550);
or U16921 (N_16921,N_15097,N_15121);
and U16922 (N_16922,N_15645,N_15716);
nand U16923 (N_16923,N_15149,N_15544);
nor U16924 (N_16924,N_15560,N_15672);
and U16925 (N_16925,N_15912,N_15854);
xor U16926 (N_16926,N_15090,N_15766);
nor U16927 (N_16927,N_15583,N_15570);
nand U16928 (N_16928,N_15970,N_15264);
and U16929 (N_16929,N_15275,N_15309);
and U16930 (N_16930,N_15089,N_15372);
or U16931 (N_16931,N_15989,N_15813);
nor U16932 (N_16932,N_15642,N_15368);
and U16933 (N_16933,N_15097,N_15796);
and U16934 (N_16934,N_15288,N_15722);
xor U16935 (N_16935,N_15948,N_15739);
or U16936 (N_16936,N_15479,N_15286);
or U16937 (N_16937,N_15531,N_15119);
xor U16938 (N_16938,N_15708,N_15112);
and U16939 (N_16939,N_15226,N_15847);
and U16940 (N_16940,N_15189,N_15488);
and U16941 (N_16941,N_15753,N_15295);
nor U16942 (N_16942,N_15219,N_15388);
and U16943 (N_16943,N_15358,N_15988);
and U16944 (N_16944,N_15842,N_15565);
nor U16945 (N_16945,N_15383,N_15116);
nand U16946 (N_16946,N_15233,N_15438);
nor U16947 (N_16947,N_15975,N_15722);
nand U16948 (N_16948,N_15201,N_15156);
nand U16949 (N_16949,N_15854,N_15100);
and U16950 (N_16950,N_15522,N_15455);
nand U16951 (N_16951,N_15755,N_15603);
nand U16952 (N_16952,N_15836,N_15809);
nor U16953 (N_16953,N_15336,N_15554);
and U16954 (N_16954,N_15302,N_15447);
and U16955 (N_16955,N_15581,N_15454);
nor U16956 (N_16956,N_15609,N_15877);
nand U16957 (N_16957,N_15937,N_15326);
and U16958 (N_16958,N_15300,N_15597);
xor U16959 (N_16959,N_15725,N_15084);
nor U16960 (N_16960,N_15594,N_15705);
xnor U16961 (N_16961,N_15372,N_15948);
or U16962 (N_16962,N_15331,N_15726);
or U16963 (N_16963,N_15299,N_15927);
or U16964 (N_16964,N_15663,N_15080);
xnor U16965 (N_16965,N_15327,N_15143);
and U16966 (N_16966,N_15837,N_15426);
and U16967 (N_16967,N_15934,N_15498);
xor U16968 (N_16968,N_15330,N_15661);
and U16969 (N_16969,N_15700,N_15411);
nand U16970 (N_16970,N_15025,N_15905);
nand U16971 (N_16971,N_15634,N_15155);
or U16972 (N_16972,N_15907,N_15363);
nand U16973 (N_16973,N_15755,N_15934);
nand U16974 (N_16974,N_15741,N_15100);
nand U16975 (N_16975,N_15680,N_15080);
and U16976 (N_16976,N_15774,N_15003);
or U16977 (N_16977,N_15077,N_15701);
xnor U16978 (N_16978,N_15781,N_15403);
xnor U16979 (N_16979,N_15013,N_15229);
and U16980 (N_16980,N_15489,N_15852);
or U16981 (N_16981,N_15669,N_15779);
and U16982 (N_16982,N_15344,N_15253);
xor U16983 (N_16983,N_15335,N_15477);
and U16984 (N_16984,N_15877,N_15927);
and U16985 (N_16985,N_15869,N_15527);
or U16986 (N_16986,N_15782,N_15427);
nand U16987 (N_16987,N_15394,N_15842);
and U16988 (N_16988,N_15211,N_15890);
nor U16989 (N_16989,N_15090,N_15651);
nand U16990 (N_16990,N_15744,N_15540);
xor U16991 (N_16991,N_15868,N_15746);
and U16992 (N_16992,N_15082,N_15300);
nor U16993 (N_16993,N_15804,N_15816);
and U16994 (N_16994,N_15514,N_15234);
or U16995 (N_16995,N_15715,N_15583);
nand U16996 (N_16996,N_15113,N_15514);
xnor U16997 (N_16997,N_15572,N_15393);
xor U16998 (N_16998,N_15788,N_15199);
and U16999 (N_16999,N_15855,N_15539);
nand U17000 (N_17000,N_16183,N_16685);
or U17001 (N_17001,N_16781,N_16537);
or U17002 (N_17002,N_16069,N_16786);
nor U17003 (N_17003,N_16611,N_16332);
xor U17004 (N_17004,N_16251,N_16408);
nor U17005 (N_17005,N_16006,N_16617);
xnor U17006 (N_17006,N_16501,N_16861);
or U17007 (N_17007,N_16126,N_16149);
nor U17008 (N_17008,N_16499,N_16842);
nor U17009 (N_17009,N_16736,N_16667);
nor U17010 (N_17010,N_16462,N_16592);
and U17011 (N_17011,N_16797,N_16366);
or U17012 (N_17012,N_16027,N_16487);
and U17013 (N_17013,N_16282,N_16729);
nand U17014 (N_17014,N_16692,N_16690);
xor U17015 (N_17015,N_16572,N_16148);
or U17016 (N_17016,N_16376,N_16803);
xor U17017 (N_17017,N_16991,N_16377);
xor U17018 (N_17018,N_16684,N_16841);
and U17019 (N_17019,N_16065,N_16862);
nor U17020 (N_17020,N_16832,N_16243);
nor U17021 (N_17021,N_16210,N_16494);
xor U17022 (N_17022,N_16099,N_16691);
and U17023 (N_17023,N_16722,N_16478);
or U17024 (N_17024,N_16364,N_16988);
and U17025 (N_17025,N_16312,N_16048);
nor U17026 (N_17026,N_16155,N_16383);
or U17027 (N_17027,N_16698,N_16926);
nand U17028 (N_17028,N_16008,N_16568);
and U17029 (N_17029,N_16876,N_16616);
or U17030 (N_17030,N_16902,N_16680);
and U17031 (N_17031,N_16378,N_16262);
nor U17032 (N_17032,N_16012,N_16195);
and U17033 (N_17033,N_16821,N_16629);
or U17034 (N_17034,N_16475,N_16819);
nand U17035 (N_17035,N_16504,N_16765);
or U17036 (N_17036,N_16283,N_16101);
and U17037 (N_17037,N_16163,N_16066);
and U17038 (N_17038,N_16359,N_16843);
nand U17039 (N_17039,N_16347,N_16314);
or U17040 (N_17040,N_16423,N_16836);
nor U17041 (N_17041,N_16563,N_16479);
and U17042 (N_17042,N_16165,N_16724);
or U17043 (N_17043,N_16433,N_16256);
nand U17044 (N_17044,N_16938,N_16705);
or U17045 (N_17045,N_16587,N_16986);
and U17046 (N_17046,N_16707,N_16770);
xor U17047 (N_17047,N_16947,N_16513);
and U17048 (N_17048,N_16872,N_16193);
and U17049 (N_17049,N_16473,N_16522);
xor U17050 (N_17050,N_16429,N_16823);
nand U17051 (N_17051,N_16141,N_16581);
nor U17052 (N_17052,N_16084,N_16734);
nor U17053 (N_17053,N_16854,N_16606);
xnor U17054 (N_17054,N_16943,N_16791);
nor U17055 (N_17055,N_16090,N_16010);
xnor U17056 (N_17056,N_16888,N_16583);
or U17057 (N_17057,N_16093,N_16655);
xor U17058 (N_17058,N_16554,N_16915);
or U17059 (N_17059,N_16735,N_16425);
nor U17060 (N_17060,N_16981,N_16026);
or U17061 (N_17061,N_16485,N_16622);
or U17062 (N_17062,N_16397,N_16457);
and U17063 (N_17063,N_16777,N_16815);
or U17064 (N_17064,N_16236,N_16247);
nand U17065 (N_17065,N_16345,N_16086);
or U17066 (N_17066,N_16711,N_16644);
and U17067 (N_17067,N_16933,N_16410);
or U17068 (N_17068,N_16758,N_16204);
and U17069 (N_17069,N_16388,N_16496);
nand U17070 (N_17070,N_16580,N_16182);
xnor U17071 (N_17071,N_16545,N_16444);
xor U17072 (N_17072,N_16398,N_16437);
or U17073 (N_17073,N_16367,N_16699);
nand U17074 (N_17074,N_16952,N_16325);
nand U17075 (N_17075,N_16212,N_16826);
nand U17076 (N_17076,N_16929,N_16845);
or U17077 (N_17077,N_16994,N_16795);
nand U17078 (N_17078,N_16802,N_16194);
nor U17079 (N_17079,N_16111,N_16414);
xor U17080 (N_17080,N_16743,N_16600);
nand U17081 (N_17081,N_16466,N_16497);
xnor U17082 (N_17082,N_16351,N_16411);
or U17083 (N_17083,N_16089,N_16328);
nand U17084 (N_17084,N_16272,N_16471);
nor U17085 (N_17085,N_16483,N_16740);
and U17086 (N_17086,N_16597,N_16811);
nor U17087 (N_17087,N_16331,N_16258);
or U17088 (N_17088,N_16674,N_16436);
xnor U17089 (N_17089,N_16894,N_16002);
xor U17090 (N_17090,N_16558,N_16983);
or U17091 (N_17091,N_16748,N_16123);
xnor U17092 (N_17092,N_16028,N_16418);
xor U17093 (N_17093,N_16589,N_16118);
nor U17094 (N_17094,N_16595,N_16989);
nor U17095 (N_17095,N_16827,N_16159);
nand U17096 (N_17096,N_16224,N_16532);
xnor U17097 (N_17097,N_16395,N_16682);
nor U17098 (N_17098,N_16396,N_16403);
xnor U17099 (N_17099,N_16630,N_16225);
and U17100 (N_17100,N_16556,N_16879);
nand U17101 (N_17101,N_16577,N_16753);
or U17102 (N_17102,N_16199,N_16566);
nor U17103 (N_17103,N_16930,N_16604);
xnor U17104 (N_17104,N_16533,N_16480);
and U17105 (N_17105,N_16144,N_16439);
xnor U17106 (N_17106,N_16454,N_16688);
nor U17107 (N_17107,N_16263,N_16078);
xnor U17108 (N_17108,N_16279,N_16432);
nand U17109 (N_17109,N_16030,N_16979);
nand U17110 (N_17110,N_16571,N_16387);
or U17111 (N_17111,N_16920,N_16640);
and U17112 (N_17112,N_16723,N_16130);
xnor U17113 (N_17113,N_16421,N_16461);
and U17114 (N_17114,N_16612,N_16113);
nand U17115 (N_17115,N_16467,N_16664);
nor U17116 (N_17116,N_16694,N_16759);
xor U17117 (N_17117,N_16881,N_16095);
nor U17118 (N_17118,N_16072,N_16883);
nor U17119 (N_17119,N_16603,N_16767);
or U17120 (N_17120,N_16763,N_16591);
and U17121 (N_17121,N_16202,N_16878);
and U17122 (N_17122,N_16162,N_16553);
nor U17123 (N_17123,N_16908,N_16018);
nand U17124 (N_17124,N_16151,N_16135);
xnor U17125 (N_17125,N_16169,N_16393);
and U17126 (N_17126,N_16493,N_16207);
xor U17127 (N_17127,N_16642,N_16284);
nor U17128 (N_17128,N_16338,N_16799);
or U17129 (N_17129,N_16870,N_16904);
nand U17130 (N_17130,N_16211,N_16570);
xnor U17131 (N_17131,N_16448,N_16489);
nand U17132 (N_17132,N_16768,N_16999);
and U17133 (N_17133,N_16818,N_16059);
xor U17134 (N_17134,N_16713,N_16716);
nand U17135 (N_17135,N_16961,N_16068);
or U17136 (N_17136,N_16939,N_16209);
nand U17137 (N_17137,N_16588,N_16316);
and U17138 (N_17138,N_16678,N_16001);
xnor U17139 (N_17139,N_16661,N_16333);
or U17140 (N_17140,N_16228,N_16932);
or U17141 (N_17141,N_16775,N_16728);
and U17142 (N_17142,N_16732,N_16715);
nand U17143 (N_17143,N_16341,N_16040);
or U17144 (N_17144,N_16222,N_16746);
nor U17145 (N_17145,N_16017,N_16356);
nor U17146 (N_17146,N_16276,N_16181);
nor U17147 (N_17147,N_16773,N_16557);
and U17148 (N_17148,N_16146,N_16175);
nor U17149 (N_17149,N_16108,N_16274);
xor U17150 (N_17150,N_16598,N_16428);
or U17151 (N_17151,N_16087,N_16374);
or U17152 (N_17152,N_16621,N_16669);
and U17153 (N_17153,N_16838,N_16180);
and U17154 (N_17154,N_16186,N_16188);
xor U17155 (N_17155,N_16683,N_16252);
nand U17156 (N_17156,N_16131,N_16754);
nand U17157 (N_17157,N_16830,N_16191);
xor U17158 (N_17158,N_16071,N_16668);
or U17159 (N_17159,N_16197,N_16492);
xor U17160 (N_17160,N_16599,N_16745);
nor U17161 (N_17161,N_16968,N_16807);
or U17162 (N_17162,N_16885,N_16127);
nand U17163 (N_17163,N_16280,N_16384);
nor U17164 (N_17164,N_16415,N_16465);
xnor U17165 (N_17165,N_16995,N_16585);
and U17166 (N_17166,N_16275,N_16452);
or U17167 (N_17167,N_16360,N_16992);
xnor U17168 (N_17168,N_16075,N_16547);
nand U17169 (N_17169,N_16520,N_16652);
and U17170 (N_17170,N_16132,N_16663);
or U17171 (N_17171,N_16601,N_16829);
nor U17172 (N_17172,N_16925,N_16311);
and U17173 (N_17173,N_16246,N_16404);
xor U17174 (N_17174,N_16326,N_16910);
xor U17175 (N_17175,N_16476,N_16718);
nor U17176 (N_17176,N_16498,N_16831);
nand U17177 (N_17177,N_16302,N_16851);
or U17178 (N_17178,N_16613,N_16079);
xor U17179 (N_17179,N_16747,N_16117);
and U17180 (N_17180,N_16731,N_16633);
nand U17181 (N_17181,N_16297,N_16164);
nor U17182 (N_17182,N_16092,N_16295);
nand U17183 (N_17183,N_16844,N_16950);
and U17184 (N_17184,N_16919,N_16420);
nand U17185 (N_17185,N_16561,N_16525);
nor U17186 (N_17186,N_16771,N_16172);
nand U17187 (N_17187,N_16864,N_16317);
nand U17188 (N_17188,N_16218,N_16975);
or U17189 (N_17189,N_16637,N_16049);
and U17190 (N_17190,N_16594,N_16299);
nand U17191 (N_17191,N_16430,N_16413);
nor U17192 (N_17192,N_16103,N_16120);
nor U17193 (N_17193,N_16638,N_16177);
nor U17194 (N_17194,N_16179,N_16798);
nor U17195 (N_17195,N_16329,N_16858);
or U17196 (N_17196,N_16353,N_16835);
or U17197 (N_17197,N_16456,N_16080);
and U17198 (N_17198,N_16004,N_16375);
xor U17199 (N_17199,N_16038,N_16041);
xor U17200 (N_17200,N_16447,N_16714);
and U17201 (N_17201,N_16305,N_16890);
nor U17202 (N_17202,N_16727,N_16273);
nand U17203 (N_17203,N_16145,N_16521);
and U17204 (N_17204,N_16552,N_16906);
nor U17205 (N_17205,N_16646,N_16506);
xor U17206 (N_17206,N_16515,N_16647);
nand U17207 (N_17207,N_16837,N_16708);
and U17208 (N_17208,N_16666,N_16227);
or U17209 (N_17209,N_16726,N_16201);
or U17210 (N_17210,N_16871,N_16023);
or U17211 (N_17211,N_16076,N_16689);
and U17212 (N_17212,N_16945,N_16507);
and U17213 (N_17213,N_16468,N_16056);
nor U17214 (N_17214,N_16266,N_16278);
and U17215 (N_17215,N_16917,N_16636);
nor U17216 (N_17216,N_16639,N_16189);
nand U17217 (N_17217,N_16741,N_16531);
or U17218 (N_17218,N_16060,N_16565);
nand U17219 (N_17219,N_16336,N_16451);
or U17220 (N_17220,N_16882,N_16789);
xnor U17221 (N_17221,N_16527,N_16957);
or U17222 (N_17222,N_16912,N_16379);
xnor U17223 (N_17223,N_16907,N_16422);
or U17224 (N_17224,N_16304,N_16675);
nand U17225 (N_17225,N_16058,N_16490);
and U17226 (N_17226,N_16972,N_16441);
nor U17227 (N_17227,N_16769,N_16486);
nand U17228 (N_17228,N_16013,N_16369);
and U17229 (N_17229,N_16956,N_16955);
nand U17230 (N_17230,N_16213,N_16516);
or U17231 (N_17231,N_16687,N_16648);
nand U17232 (N_17232,N_16112,N_16863);
or U17233 (N_17233,N_16511,N_16443);
xor U17234 (N_17234,N_16147,N_16916);
and U17235 (N_17235,N_16372,N_16880);
xnor U17236 (N_17236,N_16055,N_16154);
xnor U17237 (N_17237,N_16898,N_16509);
xnor U17238 (N_17238,N_16405,N_16381);
xnor U17239 (N_17239,N_16964,N_16899);
and U17240 (N_17240,N_16321,N_16564);
xnor U17241 (N_17241,N_16751,N_16082);
nand U17242 (N_17242,N_16470,N_16229);
and U17243 (N_17243,N_16039,N_16801);
or U17244 (N_17244,N_16971,N_16105);
nand U17245 (N_17245,N_16551,N_16942);
nand U17246 (N_17246,N_16518,N_16267);
nor U17247 (N_17247,N_16869,N_16709);
nand U17248 (N_17248,N_16535,N_16217);
nand U17249 (N_17249,N_16253,N_16744);
and U17250 (N_17250,N_16053,N_16109);
and U17251 (N_17251,N_16867,N_16996);
xor U17252 (N_17252,N_16185,N_16043);
xnor U17253 (N_17253,N_16969,N_16074);
nand U17254 (N_17254,N_16339,N_16820);
nor U17255 (N_17255,N_16755,N_16787);
nand U17256 (N_17256,N_16503,N_16584);
and U17257 (N_17257,N_16987,N_16085);
xor U17258 (N_17258,N_16358,N_16800);
xor U17259 (N_17259,N_16665,N_16635);
or U17260 (N_17260,N_16788,N_16241);
nand U17261 (N_17261,N_16081,N_16104);
or U17262 (N_17262,N_16346,N_16340);
nand U17263 (N_17263,N_16784,N_16070);
nor U17264 (N_17264,N_16774,N_16052);
nor U17265 (N_17265,N_16555,N_16719);
xor U17266 (N_17266,N_16575,N_16324);
nor U17267 (N_17267,N_16142,N_16519);
and U17268 (N_17268,N_16481,N_16416);
and U17269 (N_17269,N_16913,N_16125);
nand U17270 (N_17270,N_16538,N_16288);
xor U17271 (N_17271,N_16290,N_16510);
xnor U17272 (N_17272,N_16849,N_16064);
nand U17273 (N_17273,N_16319,N_16946);
xor U17274 (N_17274,N_16050,N_16805);
or U17275 (N_17275,N_16828,N_16344);
nand U17276 (N_17276,N_16671,N_16242);
or U17277 (N_17277,N_16540,N_16446);
nor U17278 (N_17278,N_16037,N_16891);
or U17279 (N_17279,N_16419,N_16286);
nor U17280 (N_17280,N_16931,N_16610);
nor U17281 (N_17281,N_16921,N_16122);
xnor U17282 (N_17282,N_16614,N_16063);
or U17283 (N_17283,N_16624,N_16119);
or U17284 (N_17284,N_16237,N_16459);
nand U17285 (N_17285,N_16641,N_16400);
nor U17286 (N_17286,N_16918,N_16619);
xnor U17287 (N_17287,N_16173,N_16960);
xnor U17288 (N_17288,N_16752,N_16783);
and U17289 (N_17289,N_16015,N_16717);
and U17290 (N_17290,N_16327,N_16281);
or U17291 (N_17291,N_16382,N_16500);
or U17292 (N_17292,N_16067,N_16596);
and U17293 (N_17293,N_16261,N_16772);
nand U17294 (N_17294,N_16143,N_16895);
nand U17295 (N_17295,N_16541,N_16025);
and U17296 (N_17296,N_16623,N_16865);
xor U17297 (N_17297,N_16285,N_16115);
nand U17298 (N_17298,N_16927,N_16137);
or U17299 (N_17299,N_16576,N_16649);
nand U17300 (N_17300,N_16350,N_16114);
nand U17301 (N_17301,N_16094,N_16593);
nor U17302 (N_17302,N_16007,N_16679);
nand U17303 (N_17303,N_16733,N_16116);
nor U17304 (N_17304,N_16196,N_16477);
nand U17305 (N_17305,N_16928,N_16003);
xor U17306 (N_17306,N_16270,N_16550);
or U17307 (N_17307,N_16233,N_16737);
xor U17308 (N_17308,N_16293,N_16238);
nand U17309 (N_17309,N_16965,N_16847);
nand U17310 (N_17310,N_16349,N_16255);
or U17311 (N_17311,N_16192,N_16984);
xor U17312 (N_17312,N_16721,N_16824);
nor U17313 (N_17313,N_16098,N_16982);
and U17314 (N_17314,N_16259,N_16216);
xor U17315 (N_17315,N_16287,N_16993);
and U17316 (N_17316,N_16368,N_16062);
nand U17317 (N_17317,N_16582,N_16045);
nor U17318 (N_17318,N_16019,N_16232);
xnor U17319 (N_17319,N_16677,N_16884);
nand U17320 (N_17320,N_16488,N_16778);
nand U17321 (N_17321,N_16846,N_16277);
or U17322 (N_17322,N_16296,N_16785);
nor U17323 (N_17323,N_16790,N_16703);
nand U17324 (N_17324,N_16330,N_16036);
nor U17325 (N_17325,N_16412,N_16502);
nor U17326 (N_17326,N_16107,N_16586);
nor U17327 (N_17327,N_16817,N_16607);
and U17328 (N_17328,N_16720,N_16442);
xnor U17329 (N_17329,N_16234,N_16549);
nor U17330 (N_17330,N_16460,N_16491);
or U17331 (N_17331,N_16569,N_16438);
nand U17332 (N_17332,N_16529,N_16187);
xor U17333 (N_17333,N_16054,N_16974);
nor U17334 (N_17334,N_16934,N_16046);
xnor U17335 (N_17335,N_16980,N_16463);
and U17336 (N_17336,N_16365,N_16424);
nor U17337 (N_17337,N_16985,N_16348);
and U17338 (N_17338,N_16219,N_16014);
or U17339 (N_17339,N_16294,N_16660);
or U17340 (N_17340,N_16264,N_16352);
or U17341 (N_17341,N_16306,N_16402);
nor U17342 (N_17342,N_16361,N_16833);
and U17343 (N_17343,N_16035,N_16291);
nand U17344 (N_17344,N_16335,N_16176);
and U17345 (N_17345,N_16031,N_16962);
and U17346 (N_17346,N_16651,N_16909);
xnor U17347 (N_17347,N_16091,N_16248);
or U17348 (N_17348,N_16860,N_16696);
xnor U17349 (N_17349,N_16453,N_16954);
nor U17350 (N_17350,N_16464,N_16710);
xnor U17351 (N_17351,N_16536,N_16385);
and U17352 (N_17352,N_16150,N_16897);
nand U17353 (N_17353,N_16997,N_16271);
nor U17354 (N_17354,N_16548,N_16407);
and U17355 (N_17355,N_16203,N_16840);
nor U17356 (N_17356,N_16579,N_16399);
nor U17357 (N_17357,N_16578,N_16124);
and U17358 (N_17358,N_16215,N_16848);
nor U17359 (N_17359,N_16922,N_16370);
and U17360 (N_17360,N_16362,N_16469);
xnor U17361 (N_17361,N_16776,N_16605);
nor U17362 (N_17362,N_16033,N_16005);
and U17363 (N_17363,N_16978,N_16935);
or U17364 (N_17364,N_16235,N_16307);
and U17365 (N_17365,N_16334,N_16310);
nand U17366 (N_17366,N_16426,N_16450);
nand U17367 (N_17367,N_16766,N_16656);
and U17368 (N_17368,N_16941,N_16022);
nor U17369 (N_17369,N_16153,N_16102);
xnor U17370 (N_17370,N_16673,N_16260);
or U17371 (N_17371,N_16896,N_16289);
nand U17372 (N_17372,N_16544,N_16914);
nor U17373 (N_17373,N_16292,N_16427);
and U17374 (N_17374,N_16738,N_16940);
or U17375 (N_17375,N_16615,N_16160);
nor U17376 (N_17376,N_16905,N_16354);
xor U17377 (N_17377,N_16371,N_16546);
and U17378 (N_17378,N_16524,N_16810);
nor U17379 (N_17379,N_16574,N_16355);
nor U17380 (N_17380,N_16138,N_16514);
nor U17381 (N_17381,N_16530,N_16839);
or U17382 (N_17382,N_16812,N_16873);
and U17383 (N_17383,N_16061,N_16000);
nand U17384 (N_17384,N_16024,N_16313);
nand U17385 (N_17385,N_16875,N_16166);
nor U17386 (N_17386,N_16814,N_16756);
or U17387 (N_17387,N_16866,N_16976);
nand U17388 (N_17388,N_16449,N_16445);
or U17389 (N_17389,N_16517,N_16363);
or U17390 (N_17390,N_16032,N_16226);
nand U17391 (N_17391,N_16662,N_16936);
or U17392 (N_17392,N_16152,N_16484);
xnor U17393 (N_17393,N_16857,N_16813);
nor U17394 (N_17394,N_16750,N_16170);
or U17395 (N_17395,N_16590,N_16762);
xor U17396 (N_17396,N_16602,N_16850);
xor U17397 (N_17397,N_16171,N_16967);
nand U17398 (N_17398,N_16676,N_16609);
and U17399 (N_17399,N_16077,N_16816);
nand U17400 (N_17400,N_16392,N_16409);
or U17401 (N_17401,N_16659,N_16323);
nand U17402 (N_17402,N_16508,N_16200);
or U17403 (N_17403,N_16792,N_16534);
nand U17404 (N_17404,N_16106,N_16998);
nor U17405 (N_17405,N_16889,N_16697);
nand U17406 (N_17406,N_16834,N_16300);
or U17407 (N_17407,N_16859,N_16764);
nor U17408 (N_17408,N_16139,N_16780);
nand U17409 (N_17409,N_16309,N_16240);
xnor U17410 (N_17410,N_16900,N_16949);
nor U17411 (N_17411,N_16220,N_16244);
nand U17412 (N_17412,N_16097,N_16853);
nor U17413 (N_17413,N_16631,N_16704);
nor U17414 (N_17414,N_16560,N_16632);
or U17415 (N_17415,N_16214,N_16269);
or U17416 (N_17416,N_16318,N_16695);
or U17417 (N_17417,N_16455,N_16342);
and U17418 (N_17418,N_16406,N_16208);
and U17419 (N_17419,N_16653,N_16953);
nor U17420 (N_17420,N_16794,N_16742);
and U17421 (N_17421,N_16057,N_16245);
nor U17422 (N_17422,N_16990,N_16923);
nand U17423 (N_17423,N_16944,N_16657);
nor U17424 (N_17424,N_16482,N_16051);
xnor U17425 (N_17425,N_16128,N_16793);
xor U17426 (N_17426,N_16110,N_16526);
xor U17427 (N_17427,N_16136,N_16205);
and U17428 (N_17428,N_16250,N_16417);
nor U17429 (N_17429,N_16239,N_16628);
or U17430 (N_17430,N_16730,N_16198);
xnor U17431 (N_17431,N_16693,N_16320);
and U17432 (N_17432,N_16658,N_16825);
nand U17433 (N_17433,N_16431,N_16959);
or U17434 (N_17434,N_16394,N_16343);
nand U17435 (N_17435,N_16528,N_16523);
nor U17436 (N_17436,N_16073,N_16458);
xor U17437 (N_17437,N_16626,N_16706);
or U17438 (N_17438,N_16887,N_16702);
or U17439 (N_17439,N_16686,N_16391);
xnor U17440 (N_17440,N_16654,N_16643);
nand U17441 (N_17441,N_16380,N_16701);
nand U17442 (N_17442,N_16474,N_16133);
or U17443 (N_17443,N_16440,N_16167);
or U17444 (N_17444,N_16782,N_16357);
nand U17445 (N_17445,N_16505,N_16650);
nand U17446 (N_17446,N_16096,N_16559);
or U17447 (N_17447,N_16620,N_16373);
nand U17448 (N_17448,N_16042,N_16796);
or U17449 (N_17449,N_16562,N_16963);
xnor U17450 (N_17450,N_16308,N_16977);
nor U17451 (N_17451,N_16011,N_16009);
or U17452 (N_17452,N_16855,N_16121);
xor U17453 (N_17453,N_16924,N_16761);
xor U17454 (N_17454,N_16168,N_16757);
and U17455 (N_17455,N_16966,N_16044);
and U17456 (N_17456,N_16970,N_16749);
nor U17457 (N_17457,N_16911,N_16760);
xor U17458 (N_17458,N_16495,N_16034);
or U17459 (N_17459,N_16948,N_16856);
and U17460 (N_17460,N_16809,N_16618);
and U17461 (N_17461,N_16184,N_16221);
or U17462 (N_17462,N_16901,N_16020);
nand U17463 (N_17463,N_16301,N_16223);
nand U17464 (N_17464,N_16021,N_16337);
or U17465 (N_17465,N_16088,N_16973);
and U17466 (N_17466,N_16190,N_16512);
nand U17467 (N_17467,N_16134,N_16157);
xnor U17468 (N_17468,N_16877,N_16886);
nor U17469 (N_17469,N_16543,N_16230);
nor U17470 (N_17470,N_16156,N_16958);
xnor U17471 (N_17471,N_16100,N_16083);
nor U17472 (N_17472,N_16401,N_16852);
xnor U17473 (N_17473,N_16472,N_16634);
nor U17474 (N_17474,N_16892,N_16322);
xor U17475 (N_17475,N_16542,N_16206);
nor U17476 (N_17476,N_16303,N_16567);
or U17477 (N_17477,N_16386,N_16231);
and U17478 (N_17478,N_16268,N_16047);
nand U17479 (N_17479,N_16645,N_16315);
nor U17480 (N_17480,N_16903,N_16389);
xor U17481 (N_17481,N_16739,N_16937);
or U17482 (N_17482,N_16178,N_16804);
nand U17483 (N_17483,N_16029,N_16779);
nand U17484 (N_17484,N_16874,N_16808);
or U17485 (N_17485,N_16681,N_16700);
xnor U17486 (N_17486,N_16608,N_16806);
or U17487 (N_17487,N_16712,N_16822);
nand U17488 (N_17488,N_16868,N_16265);
nand U17489 (N_17489,N_16298,N_16435);
and U17490 (N_17490,N_16174,N_16670);
nand U17491 (N_17491,N_16539,N_16016);
xor U17492 (N_17492,N_16390,N_16257);
xor U17493 (N_17493,N_16254,N_16725);
nand U17494 (N_17494,N_16434,N_16161);
or U17495 (N_17495,N_16573,N_16129);
nand U17496 (N_17496,N_16140,N_16625);
and U17497 (N_17497,N_16672,N_16627);
xnor U17498 (N_17498,N_16158,N_16951);
nand U17499 (N_17499,N_16249,N_16893);
xor U17500 (N_17500,N_16037,N_16944);
xor U17501 (N_17501,N_16115,N_16046);
nor U17502 (N_17502,N_16184,N_16896);
and U17503 (N_17503,N_16978,N_16147);
or U17504 (N_17504,N_16456,N_16192);
nand U17505 (N_17505,N_16657,N_16746);
and U17506 (N_17506,N_16620,N_16301);
xnor U17507 (N_17507,N_16671,N_16426);
and U17508 (N_17508,N_16519,N_16313);
and U17509 (N_17509,N_16776,N_16545);
nor U17510 (N_17510,N_16900,N_16586);
nand U17511 (N_17511,N_16151,N_16988);
xor U17512 (N_17512,N_16141,N_16629);
nor U17513 (N_17513,N_16373,N_16296);
nor U17514 (N_17514,N_16051,N_16864);
or U17515 (N_17515,N_16401,N_16199);
xnor U17516 (N_17516,N_16453,N_16380);
and U17517 (N_17517,N_16976,N_16679);
or U17518 (N_17518,N_16998,N_16242);
or U17519 (N_17519,N_16559,N_16037);
and U17520 (N_17520,N_16527,N_16826);
or U17521 (N_17521,N_16223,N_16349);
nor U17522 (N_17522,N_16601,N_16043);
nor U17523 (N_17523,N_16685,N_16988);
and U17524 (N_17524,N_16655,N_16866);
xor U17525 (N_17525,N_16865,N_16695);
and U17526 (N_17526,N_16862,N_16008);
nor U17527 (N_17527,N_16410,N_16924);
nand U17528 (N_17528,N_16077,N_16064);
and U17529 (N_17529,N_16798,N_16300);
or U17530 (N_17530,N_16068,N_16511);
nand U17531 (N_17531,N_16742,N_16110);
xnor U17532 (N_17532,N_16410,N_16990);
xnor U17533 (N_17533,N_16411,N_16616);
nor U17534 (N_17534,N_16561,N_16912);
or U17535 (N_17535,N_16259,N_16391);
nor U17536 (N_17536,N_16887,N_16901);
xor U17537 (N_17537,N_16134,N_16844);
and U17538 (N_17538,N_16516,N_16973);
or U17539 (N_17539,N_16246,N_16471);
or U17540 (N_17540,N_16989,N_16349);
nor U17541 (N_17541,N_16037,N_16634);
and U17542 (N_17542,N_16303,N_16417);
nor U17543 (N_17543,N_16647,N_16514);
xor U17544 (N_17544,N_16721,N_16782);
or U17545 (N_17545,N_16269,N_16487);
nand U17546 (N_17546,N_16798,N_16604);
or U17547 (N_17547,N_16044,N_16914);
nor U17548 (N_17548,N_16680,N_16325);
xor U17549 (N_17549,N_16176,N_16561);
and U17550 (N_17550,N_16710,N_16741);
nand U17551 (N_17551,N_16263,N_16077);
nor U17552 (N_17552,N_16565,N_16576);
and U17553 (N_17553,N_16701,N_16012);
xor U17554 (N_17554,N_16078,N_16053);
xor U17555 (N_17555,N_16574,N_16201);
or U17556 (N_17556,N_16864,N_16526);
or U17557 (N_17557,N_16667,N_16434);
nand U17558 (N_17558,N_16423,N_16115);
nor U17559 (N_17559,N_16295,N_16442);
nand U17560 (N_17560,N_16440,N_16609);
xnor U17561 (N_17561,N_16316,N_16696);
nor U17562 (N_17562,N_16272,N_16172);
nor U17563 (N_17563,N_16076,N_16524);
nor U17564 (N_17564,N_16594,N_16688);
and U17565 (N_17565,N_16281,N_16334);
xnor U17566 (N_17566,N_16439,N_16497);
nand U17567 (N_17567,N_16274,N_16915);
nand U17568 (N_17568,N_16110,N_16178);
and U17569 (N_17569,N_16536,N_16856);
or U17570 (N_17570,N_16694,N_16218);
nand U17571 (N_17571,N_16981,N_16190);
nand U17572 (N_17572,N_16004,N_16313);
xnor U17573 (N_17573,N_16035,N_16020);
xor U17574 (N_17574,N_16888,N_16293);
nand U17575 (N_17575,N_16628,N_16959);
nor U17576 (N_17576,N_16603,N_16275);
nand U17577 (N_17577,N_16670,N_16815);
and U17578 (N_17578,N_16394,N_16095);
and U17579 (N_17579,N_16805,N_16304);
nor U17580 (N_17580,N_16964,N_16129);
and U17581 (N_17581,N_16694,N_16086);
or U17582 (N_17582,N_16020,N_16717);
nand U17583 (N_17583,N_16672,N_16336);
and U17584 (N_17584,N_16696,N_16629);
or U17585 (N_17585,N_16164,N_16818);
nor U17586 (N_17586,N_16068,N_16747);
nor U17587 (N_17587,N_16707,N_16547);
and U17588 (N_17588,N_16024,N_16762);
nand U17589 (N_17589,N_16015,N_16512);
nor U17590 (N_17590,N_16713,N_16730);
nor U17591 (N_17591,N_16462,N_16464);
xor U17592 (N_17592,N_16148,N_16423);
nor U17593 (N_17593,N_16409,N_16722);
nor U17594 (N_17594,N_16707,N_16480);
nand U17595 (N_17595,N_16716,N_16699);
nor U17596 (N_17596,N_16603,N_16641);
nor U17597 (N_17597,N_16875,N_16828);
xnor U17598 (N_17598,N_16349,N_16516);
nor U17599 (N_17599,N_16038,N_16061);
xnor U17600 (N_17600,N_16995,N_16151);
xnor U17601 (N_17601,N_16191,N_16565);
nor U17602 (N_17602,N_16237,N_16317);
and U17603 (N_17603,N_16397,N_16499);
nand U17604 (N_17604,N_16560,N_16238);
and U17605 (N_17605,N_16170,N_16386);
nor U17606 (N_17606,N_16476,N_16922);
and U17607 (N_17607,N_16585,N_16306);
or U17608 (N_17608,N_16041,N_16272);
nor U17609 (N_17609,N_16289,N_16209);
and U17610 (N_17610,N_16020,N_16116);
or U17611 (N_17611,N_16752,N_16673);
nor U17612 (N_17612,N_16600,N_16648);
nor U17613 (N_17613,N_16467,N_16702);
nand U17614 (N_17614,N_16161,N_16694);
or U17615 (N_17615,N_16821,N_16088);
xor U17616 (N_17616,N_16393,N_16472);
nor U17617 (N_17617,N_16016,N_16619);
or U17618 (N_17618,N_16475,N_16199);
and U17619 (N_17619,N_16786,N_16490);
and U17620 (N_17620,N_16426,N_16032);
nor U17621 (N_17621,N_16254,N_16214);
nor U17622 (N_17622,N_16338,N_16028);
nor U17623 (N_17623,N_16911,N_16334);
and U17624 (N_17624,N_16758,N_16623);
or U17625 (N_17625,N_16079,N_16574);
nand U17626 (N_17626,N_16637,N_16339);
xor U17627 (N_17627,N_16037,N_16576);
xor U17628 (N_17628,N_16801,N_16792);
nor U17629 (N_17629,N_16551,N_16866);
nand U17630 (N_17630,N_16559,N_16064);
nor U17631 (N_17631,N_16524,N_16555);
nor U17632 (N_17632,N_16810,N_16700);
xnor U17633 (N_17633,N_16529,N_16108);
xor U17634 (N_17634,N_16071,N_16270);
and U17635 (N_17635,N_16705,N_16412);
and U17636 (N_17636,N_16408,N_16489);
xor U17637 (N_17637,N_16767,N_16636);
nand U17638 (N_17638,N_16383,N_16933);
and U17639 (N_17639,N_16654,N_16163);
or U17640 (N_17640,N_16113,N_16151);
nand U17641 (N_17641,N_16870,N_16209);
and U17642 (N_17642,N_16102,N_16065);
xor U17643 (N_17643,N_16769,N_16006);
nand U17644 (N_17644,N_16493,N_16165);
nor U17645 (N_17645,N_16063,N_16692);
or U17646 (N_17646,N_16536,N_16464);
nor U17647 (N_17647,N_16276,N_16699);
nor U17648 (N_17648,N_16850,N_16405);
or U17649 (N_17649,N_16431,N_16341);
xnor U17650 (N_17650,N_16821,N_16971);
xnor U17651 (N_17651,N_16353,N_16752);
xnor U17652 (N_17652,N_16647,N_16354);
nor U17653 (N_17653,N_16424,N_16915);
or U17654 (N_17654,N_16899,N_16641);
nand U17655 (N_17655,N_16649,N_16816);
nor U17656 (N_17656,N_16659,N_16812);
and U17657 (N_17657,N_16464,N_16759);
or U17658 (N_17658,N_16726,N_16270);
xnor U17659 (N_17659,N_16964,N_16486);
xor U17660 (N_17660,N_16044,N_16378);
and U17661 (N_17661,N_16025,N_16619);
nand U17662 (N_17662,N_16618,N_16894);
or U17663 (N_17663,N_16126,N_16963);
or U17664 (N_17664,N_16107,N_16042);
nand U17665 (N_17665,N_16285,N_16430);
and U17666 (N_17666,N_16250,N_16061);
nand U17667 (N_17667,N_16166,N_16421);
and U17668 (N_17668,N_16348,N_16908);
nor U17669 (N_17669,N_16281,N_16010);
or U17670 (N_17670,N_16567,N_16960);
or U17671 (N_17671,N_16144,N_16232);
and U17672 (N_17672,N_16949,N_16443);
nand U17673 (N_17673,N_16422,N_16730);
nor U17674 (N_17674,N_16922,N_16589);
nand U17675 (N_17675,N_16607,N_16804);
nor U17676 (N_17676,N_16547,N_16647);
nor U17677 (N_17677,N_16436,N_16764);
nand U17678 (N_17678,N_16026,N_16558);
nand U17679 (N_17679,N_16494,N_16361);
nand U17680 (N_17680,N_16800,N_16577);
nor U17681 (N_17681,N_16584,N_16481);
and U17682 (N_17682,N_16106,N_16874);
xnor U17683 (N_17683,N_16101,N_16687);
xnor U17684 (N_17684,N_16882,N_16957);
nand U17685 (N_17685,N_16516,N_16825);
xnor U17686 (N_17686,N_16215,N_16875);
or U17687 (N_17687,N_16024,N_16721);
and U17688 (N_17688,N_16620,N_16513);
and U17689 (N_17689,N_16514,N_16785);
nor U17690 (N_17690,N_16561,N_16885);
or U17691 (N_17691,N_16632,N_16272);
or U17692 (N_17692,N_16769,N_16714);
nor U17693 (N_17693,N_16528,N_16989);
nand U17694 (N_17694,N_16704,N_16040);
and U17695 (N_17695,N_16440,N_16313);
nor U17696 (N_17696,N_16169,N_16974);
xnor U17697 (N_17697,N_16658,N_16069);
nor U17698 (N_17698,N_16468,N_16185);
xnor U17699 (N_17699,N_16835,N_16760);
and U17700 (N_17700,N_16255,N_16859);
or U17701 (N_17701,N_16208,N_16478);
and U17702 (N_17702,N_16259,N_16428);
xnor U17703 (N_17703,N_16644,N_16122);
nand U17704 (N_17704,N_16029,N_16865);
xnor U17705 (N_17705,N_16980,N_16892);
or U17706 (N_17706,N_16512,N_16443);
xor U17707 (N_17707,N_16732,N_16380);
or U17708 (N_17708,N_16697,N_16200);
and U17709 (N_17709,N_16472,N_16591);
nor U17710 (N_17710,N_16263,N_16800);
nand U17711 (N_17711,N_16529,N_16666);
xor U17712 (N_17712,N_16441,N_16255);
and U17713 (N_17713,N_16344,N_16947);
and U17714 (N_17714,N_16132,N_16726);
or U17715 (N_17715,N_16415,N_16821);
nor U17716 (N_17716,N_16956,N_16756);
xor U17717 (N_17717,N_16445,N_16444);
and U17718 (N_17718,N_16860,N_16814);
and U17719 (N_17719,N_16382,N_16024);
or U17720 (N_17720,N_16054,N_16356);
nand U17721 (N_17721,N_16879,N_16428);
or U17722 (N_17722,N_16463,N_16106);
nand U17723 (N_17723,N_16333,N_16191);
and U17724 (N_17724,N_16977,N_16705);
nand U17725 (N_17725,N_16419,N_16845);
nor U17726 (N_17726,N_16882,N_16172);
and U17727 (N_17727,N_16855,N_16183);
nor U17728 (N_17728,N_16635,N_16308);
xor U17729 (N_17729,N_16197,N_16577);
nand U17730 (N_17730,N_16447,N_16682);
nand U17731 (N_17731,N_16247,N_16906);
xnor U17732 (N_17732,N_16783,N_16214);
and U17733 (N_17733,N_16613,N_16802);
nor U17734 (N_17734,N_16635,N_16646);
nand U17735 (N_17735,N_16075,N_16694);
nand U17736 (N_17736,N_16526,N_16844);
xnor U17737 (N_17737,N_16605,N_16381);
xnor U17738 (N_17738,N_16303,N_16570);
nand U17739 (N_17739,N_16925,N_16394);
xnor U17740 (N_17740,N_16731,N_16766);
nor U17741 (N_17741,N_16067,N_16192);
or U17742 (N_17742,N_16086,N_16872);
and U17743 (N_17743,N_16761,N_16577);
and U17744 (N_17744,N_16662,N_16569);
and U17745 (N_17745,N_16781,N_16695);
nor U17746 (N_17746,N_16679,N_16736);
and U17747 (N_17747,N_16286,N_16833);
nor U17748 (N_17748,N_16317,N_16488);
and U17749 (N_17749,N_16884,N_16074);
or U17750 (N_17750,N_16075,N_16754);
nor U17751 (N_17751,N_16018,N_16574);
or U17752 (N_17752,N_16526,N_16388);
xor U17753 (N_17753,N_16958,N_16031);
nor U17754 (N_17754,N_16259,N_16513);
nor U17755 (N_17755,N_16412,N_16981);
or U17756 (N_17756,N_16838,N_16634);
nor U17757 (N_17757,N_16833,N_16377);
nor U17758 (N_17758,N_16857,N_16516);
nor U17759 (N_17759,N_16969,N_16938);
nor U17760 (N_17760,N_16218,N_16559);
and U17761 (N_17761,N_16706,N_16030);
xor U17762 (N_17762,N_16714,N_16301);
xnor U17763 (N_17763,N_16035,N_16233);
nor U17764 (N_17764,N_16542,N_16021);
or U17765 (N_17765,N_16396,N_16945);
nor U17766 (N_17766,N_16481,N_16804);
nand U17767 (N_17767,N_16323,N_16533);
nand U17768 (N_17768,N_16272,N_16942);
xor U17769 (N_17769,N_16148,N_16496);
xnor U17770 (N_17770,N_16238,N_16463);
or U17771 (N_17771,N_16828,N_16140);
xnor U17772 (N_17772,N_16405,N_16205);
nand U17773 (N_17773,N_16430,N_16783);
nand U17774 (N_17774,N_16527,N_16333);
nor U17775 (N_17775,N_16646,N_16601);
or U17776 (N_17776,N_16560,N_16056);
xor U17777 (N_17777,N_16837,N_16570);
nor U17778 (N_17778,N_16812,N_16992);
nand U17779 (N_17779,N_16131,N_16344);
or U17780 (N_17780,N_16173,N_16930);
xor U17781 (N_17781,N_16347,N_16397);
nand U17782 (N_17782,N_16385,N_16477);
nor U17783 (N_17783,N_16977,N_16230);
or U17784 (N_17784,N_16178,N_16992);
nor U17785 (N_17785,N_16117,N_16731);
or U17786 (N_17786,N_16052,N_16394);
nand U17787 (N_17787,N_16142,N_16136);
and U17788 (N_17788,N_16865,N_16468);
nor U17789 (N_17789,N_16089,N_16243);
xnor U17790 (N_17790,N_16774,N_16733);
nor U17791 (N_17791,N_16261,N_16726);
nor U17792 (N_17792,N_16533,N_16347);
and U17793 (N_17793,N_16793,N_16310);
nand U17794 (N_17794,N_16647,N_16877);
nand U17795 (N_17795,N_16386,N_16609);
xnor U17796 (N_17796,N_16175,N_16730);
xnor U17797 (N_17797,N_16150,N_16030);
and U17798 (N_17798,N_16243,N_16732);
nand U17799 (N_17799,N_16506,N_16993);
or U17800 (N_17800,N_16638,N_16613);
nand U17801 (N_17801,N_16779,N_16535);
or U17802 (N_17802,N_16412,N_16393);
xnor U17803 (N_17803,N_16362,N_16358);
or U17804 (N_17804,N_16427,N_16563);
nor U17805 (N_17805,N_16655,N_16115);
or U17806 (N_17806,N_16134,N_16875);
or U17807 (N_17807,N_16992,N_16259);
xor U17808 (N_17808,N_16283,N_16083);
or U17809 (N_17809,N_16584,N_16439);
nor U17810 (N_17810,N_16513,N_16374);
nor U17811 (N_17811,N_16725,N_16186);
xor U17812 (N_17812,N_16807,N_16771);
and U17813 (N_17813,N_16387,N_16052);
nand U17814 (N_17814,N_16088,N_16751);
nor U17815 (N_17815,N_16273,N_16078);
nor U17816 (N_17816,N_16142,N_16449);
nand U17817 (N_17817,N_16692,N_16228);
nor U17818 (N_17818,N_16282,N_16538);
nor U17819 (N_17819,N_16519,N_16597);
xor U17820 (N_17820,N_16332,N_16107);
or U17821 (N_17821,N_16760,N_16108);
nand U17822 (N_17822,N_16221,N_16798);
nor U17823 (N_17823,N_16299,N_16314);
nor U17824 (N_17824,N_16941,N_16991);
nor U17825 (N_17825,N_16388,N_16927);
and U17826 (N_17826,N_16789,N_16456);
nand U17827 (N_17827,N_16523,N_16237);
nand U17828 (N_17828,N_16973,N_16744);
xnor U17829 (N_17829,N_16031,N_16298);
and U17830 (N_17830,N_16529,N_16832);
or U17831 (N_17831,N_16006,N_16796);
or U17832 (N_17832,N_16596,N_16319);
nand U17833 (N_17833,N_16458,N_16856);
xor U17834 (N_17834,N_16921,N_16884);
nand U17835 (N_17835,N_16735,N_16739);
xor U17836 (N_17836,N_16309,N_16184);
xor U17837 (N_17837,N_16551,N_16696);
nor U17838 (N_17838,N_16142,N_16731);
nor U17839 (N_17839,N_16613,N_16273);
or U17840 (N_17840,N_16531,N_16142);
nor U17841 (N_17841,N_16754,N_16935);
nor U17842 (N_17842,N_16690,N_16686);
xor U17843 (N_17843,N_16988,N_16226);
or U17844 (N_17844,N_16577,N_16802);
nand U17845 (N_17845,N_16070,N_16405);
or U17846 (N_17846,N_16430,N_16903);
xnor U17847 (N_17847,N_16053,N_16973);
or U17848 (N_17848,N_16288,N_16321);
nor U17849 (N_17849,N_16863,N_16337);
or U17850 (N_17850,N_16151,N_16824);
xor U17851 (N_17851,N_16021,N_16793);
or U17852 (N_17852,N_16245,N_16196);
and U17853 (N_17853,N_16640,N_16885);
nand U17854 (N_17854,N_16752,N_16523);
xnor U17855 (N_17855,N_16759,N_16647);
nand U17856 (N_17856,N_16666,N_16573);
nand U17857 (N_17857,N_16436,N_16661);
xor U17858 (N_17858,N_16310,N_16629);
nand U17859 (N_17859,N_16347,N_16853);
nor U17860 (N_17860,N_16421,N_16095);
nand U17861 (N_17861,N_16914,N_16956);
or U17862 (N_17862,N_16526,N_16206);
or U17863 (N_17863,N_16561,N_16490);
nand U17864 (N_17864,N_16184,N_16925);
xnor U17865 (N_17865,N_16444,N_16857);
xnor U17866 (N_17866,N_16336,N_16924);
nand U17867 (N_17867,N_16660,N_16216);
or U17868 (N_17868,N_16772,N_16499);
nand U17869 (N_17869,N_16367,N_16238);
or U17870 (N_17870,N_16374,N_16508);
nor U17871 (N_17871,N_16540,N_16408);
or U17872 (N_17872,N_16968,N_16747);
or U17873 (N_17873,N_16681,N_16264);
nand U17874 (N_17874,N_16167,N_16528);
or U17875 (N_17875,N_16719,N_16944);
nand U17876 (N_17876,N_16670,N_16718);
xnor U17877 (N_17877,N_16597,N_16237);
and U17878 (N_17878,N_16205,N_16309);
nor U17879 (N_17879,N_16586,N_16830);
or U17880 (N_17880,N_16284,N_16682);
or U17881 (N_17881,N_16595,N_16755);
or U17882 (N_17882,N_16219,N_16524);
xor U17883 (N_17883,N_16262,N_16992);
or U17884 (N_17884,N_16109,N_16505);
or U17885 (N_17885,N_16198,N_16577);
nand U17886 (N_17886,N_16186,N_16885);
nor U17887 (N_17887,N_16556,N_16564);
nand U17888 (N_17888,N_16432,N_16916);
nor U17889 (N_17889,N_16382,N_16874);
and U17890 (N_17890,N_16964,N_16356);
or U17891 (N_17891,N_16658,N_16402);
xnor U17892 (N_17892,N_16278,N_16414);
nor U17893 (N_17893,N_16499,N_16605);
or U17894 (N_17894,N_16013,N_16232);
nand U17895 (N_17895,N_16009,N_16283);
or U17896 (N_17896,N_16303,N_16840);
or U17897 (N_17897,N_16423,N_16595);
nand U17898 (N_17898,N_16616,N_16198);
and U17899 (N_17899,N_16447,N_16945);
xnor U17900 (N_17900,N_16020,N_16323);
nor U17901 (N_17901,N_16636,N_16276);
and U17902 (N_17902,N_16604,N_16881);
and U17903 (N_17903,N_16254,N_16206);
nand U17904 (N_17904,N_16601,N_16991);
xnor U17905 (N_17905,N_16434,N_16646);
or U17906 (N_17906,N_16633,N_16504);
xor U17907 (N_17907,N_16458,N_16450);
xnor U17908 (N_17908,N_16964,N_16839);
or U17909 (N_17909,N_16117,N_16131);
nand U17910 (N_17910,N_16037,N_16194);
and U17911 (N_17911,N_16737,N_16511);
nor U17912 (N_17912,N_16169,N_16306);
xnor U17913 (N_17913,N_16548,N_16247);
or U17914 (N_17914,N_16943,N_16862);
nor U17915 (N_17915,N_16989,N_16775);
xor U17916 (N_17916,N_16734,N_16590);
and U17917 (N_17917,N_16843,N_16740);
and U17918 (N_17918,N_16208,N_16355);
or U17919 (N_17919,N_16541,N_16464);
and U17920 (N_17920,N_16114,N_16702);
nor U17921 (N_17921,N_16234,N_16146);
or U17922 (N_17922,N_16469,N_16497);
xor U17923 (N_17923,N_16306,N_16133);
xor U17924 (N_17924,N_16127,N_16492);
and U17925 (N_17925,N_16215,N_16006);
xor U17926 (N_17926,N_16882,N_16267);
nor U17927 (N_17927,N_16755,N_16865);
or U17928 (N_17928,N_16299,N_16395);
xnor U17929 (N_17929,N_16284,N_16707);
nor U17930 (N_17930,N_16822,N_16296);
or U17931 (N_17931,N_16752,N_16535);
and U17932 (N_17932,N_16145,N_16575);
nand U17933 (N_17933,N_16730,N_16819);
or U17934 (N_17934,N_16958,N_16369);
nand U17935 (N_17935,N_16430,N_16876);
or U17936 (N_17936,N_16655,N_16668);
xor U17937 (N_17937,N_16580,N_16382);
or U17938 (N_17938,N_16959,N_16733);
nand U17939 (N_17939,N_16669,N_16160);
or U17940 (N_17940,N_16891,N_16781);
or U17941 (N_17941,N_16368,N_16375);
or U17942 (N_17942,N_16568,N_16527);
and U17943 (N_17943,N_16906,N_16606);
nor U17944 (N_17944,N_16640,N_16979);
nor U17945 (N_17945,N_16711,N_16759);
nand U17946 (N_17946,N_16729,N_16021);
nand U17947 (N_17947,N_16495,N_16879);
and U17948 (N_17948,N_16892,N_16917);
xnor U17949 (N_17949,N_16193,N_16495);
xnor U17950 (N_17950,N_16838,N_16546);
xnor U17951 (N_17951,N_16400,N_16697);
or U17952 (N_17952,N_16536,N_16809);
xnor U17953 (N_17953,N_16853,N_16507);
nand U17954 (N_17954,N_16288,N_16700);
nand U17955 (N_17955,N_16694,N_16178);
nand U17956 (N_17956,N_16232,N_16917);
xnor U17957 (N_17957,N_16097,N_16123);
xnor U17958 (N_17958,N_16960,N_16288);
nor U17959 (N_17959,N_16205,N_16657);
xor U17960 (N_17960,N_16302,N_16418);
xor U17961 (N_17961,N_16246,N_16490);
nand U17962 (N_17962,N_16797,N_16468);
xor U17963 (N_17963,N_16911,N_16451);
nand U17964 (N_17964,N_16162,N_16429);
and U17965 (N_17965,N_16341,N_16966);
or U17966 (N_17966,N_16611,N_16139);
or U17967 (N_17967,N_16292,N_16093);
and U17968 (N_17968,N_16287,N_16571);
nor U17969 (N_17969,N_16818,N_16418);
nor U17970 (N_17970,N_16241,N_16554);
xor U17971 (N_17971,N_16384,N_16837);
and U17972 (N_17972,N_16971,N_16588);
nand U17973 (N_17973,N_16500,N_16668);
xor U17974 (N_17974,N_16343,N_16379);
xor U17975 (N_17975,N_16938,N_16841);
nand U17976 (N_17976,N_16567,N_16696);
and U17977 (N_17977,N_16220,N_16198);
or U17978 (N_17978,N_16286,N_16443);
nand U17979 (N_17979,N_16736,N_16059);
and U17980 (N_17980,N_16447,N_16974);
nor U17981 (N_17981,N_16309,N_16241);
or U17982 (N_17982,N_16695,N_16677);
and U17983 (N_17983,N_16935,N_16769);
nor U17984 (N_17984,N_16161,N_16889);
xor U17985 (N_17985,N_16838,N_16059);
xnor U17986 (N_17986,N_16354,N_16057);
xnor U17987 (N_17987,N_16681,N_16575);
or U17988 (N_17988,N_16635,N_16418);
xnor U17989 (N_17989,N_16419,N_16203);
and U17990 (N_17990,N_16671,N_16175);
and U17991 (N_17991,N_16241,N_16624);
and U17992 (N_17992,N_16486,N_16866);
xnor U17993 (N_17993,N_16624,N_16705);
and U17994 (N_17994,N_16691,N_16843);
nor U17995 (N_17995,N_16493,N_16537);
nand U17996 (N_17996,N_16922,N_16138);
nor U17997 (N_17997,N_16970,N_16922);
and U17998 (N_17998,N_16588,N_16394);
and U17999 (N_17999,N_16632,N_16124);
and U18000 (N_18000,N_17887,N_17736);
nor U18001 (N_18001,N_17821,N_17065);
and U18002 (N_18002,N_17341,N_17290);
or U18003 (N_18003,N_17277,N_17741);
and U18004 (N_18004,N_17940,N_17322);
nand U18005 (N_18005,N_17832,N_17441);
nor U18006 (N_18006,N_17607,N_17566);
and U18007 (N_18007,N_17299,N_17579);
or U18008 (N_18008,N_17924,N_17937);
or U18009 (N_18009,N_17011,N_17306);
or U18010 (N_18010,N_17409,N_17108);
and U18011 (N_18011,N_17119,N_17723);
nor U18012 (N_18012,N_17898,N_17684);
nor U18013 (N_18013,N_17549,N_17681);
nand U18014 (N_18014,N_17808,N_17249);
and U18015 (N_18015,N_17205,N_17484);
or U18016 (N_18016,N_17383,N_17444);
xnor U18017 (N_18017,N_17342,N_17452);
and U18018 (N_18018,N_17365,N_17507);
or U18019 (N_18019,N_17642,N_17235);
xnor U18020 (N_18020,N_17548,N_17401);
nor U18021 (N_18021,N_17818,N_17885);
and U18022 (N_18022,N_17155,N_17686);
xor U18023 (N_18023,N_17067,N_17649);
nor U18024 (N_18024,N_17653,N_17530);
nand U18025 (N_18025,N_17150,N_17433);
or U18026 (N_18026,N_17115,N_17387);
xor U18027 (N_18027,N_17586,N_17469);
and U18028 (N_18028,N_17269,N_17578);
or U18029 (N_18029,N_17671,N_17225);
xnor U18030 (N_18030,N_17001,N_17170);
or U18031 (N_18031,N_17542,N_17817);
and U18032 (N_18032,N_17377,N_17582);
or U18033 (N_18033,N_17921,N_17123);
nand U18034 (N_18034,N_17532,N_17279);
or U18035 (N_18035,N_17938,N_17431);
nor U18036 (N_18036,N_17983,N_17396);
and U18037 (N_18037,N_17997,N_17258);
nand U18038 (N_18038,N_17035,N_17192);
and U18039 (N_18039,N_17724,N_17386);
or U18040 (N_18040,N_17630,N_17312);
nand U18041 (N_18041,N_17545,N_17000);
and U18042 (N_18042,N_17491,N_17238);
or U18043 (N_18043,N_17526,N_17019);
and U18044 (N_18044,N_17841,N_17591);
or U18045 (N_18045,N_17795,N_17149);
and U18046 (N_18046,N_17091,N_17104);
nand U18047 (N_18047,N_17250,N_17971);
xnor U18048 (N_18048,N_17540,N_17505);
or U18049 (N_18049,N_17423,N_17927);
or U18050 (N_18050,N_17136,N_17959);
and U18051 (N_18051,N_17758,N_17512);
or U18052 (N_18052,N_17086,N_17862);
nor U18053 (N_18053,N_17884,N_17581);
or U18054 (N_18054,N_17730,N_17802);
and U18055 (N_18055,N_17234,N_17738);
nand U18056 (N_18056,N_17535,N_17767);
nor U18057 (N_18057,N_17111,N_17561);
nor U18058 (N_18058,N_17658,N_17044);
xor U18059 (N_18059,N_17445,N_17371);
or U18060 (N_18060,N_17287,N_17904);
or U18061 (N_18061,N_17114,N_17391);
and U18062 (N_18062,N_17351,N_17198);
or U18063 (N_18063,N_17156,N_17994);
xnor U18064 (N_18064,N_17641,N_17665);
nor U18065 (N_18065,N_17664,N_17644);
or U18066 (N_18066,N_17077,N_17326);
or U18067 (N_18067,N_17964,N_17853);
and U18068 (N_18068,N_17627,N_17575);
and U18069 (N_18069,N_17487,N_17837);
xor U18070 (N_18070,N_17403,N_17872);
nor U18071 (N_18071,N_17259,N_17295);
nand U18072 (N_18072,N_17868,N_17133);
nor U18073 (N_18073,N_17493,N_17027);
xor U18074 (N_18074,N_17138,N_17110);
xor U18075 (N_18075,N_17131,N_17834);
nand U18076 (N_18076,N_17023,N_17304);
or U18077 (N_18077,N_17359,N_17462);
nand U18078 (N_18078,N_17236,N_17333);
and U18079 (N_18079,N_17437,N_17856);
nand U18080 (N_18080,N_17038,N_17463);
and U18081 (N_18081,N_17789,N_17122);
nor U18082 (N_18082,N_17314,N_17558);
nand U18083 (N_18083,N_17323,N_17621);
nand U18084 (N_18084,N_17729,N_17501);
nand U18085 (N_18085,N_17405,N_17555);
nand U18086 (N_18086,N_17211,N_17912);
xnor U18087 (N_18087,N_17254,N_17256);
and U18088 (N_18088,N_17251,N_17537);
or U18089 (N_18089,N_17842,N_17890);
nor U18090 (N_18090,N_17950,N_17804);
xor U18091 (N_18091,N_17895,N_17367);
xor U18092 (N_18092,N_17151,N_17682);
and U18093 (N_18093,N_17756,N_17228);
and U18094 (N_18094,N_17113,N_17404);
nor U18095 (N_18095,N_17517,N_17846);
xnor U18096 (N_18096,N_17800,N_17244);
xnor U18097 (N_18097,N_17922,N_17661);
and U18098 (N_18098,N_17416,N_17739);
xor U18099 (N_18099,N_17593,N_17137);
xnor U18100 (N_18100,N_17373,N_17508);
xor U18101 (N_18101,N_17353,N_17216);
nor U18102 (N_18102,N_17900,N_17363);
and U18103 (N_18103,N_17089,N_17048);
nand U18104 (N_18104,N_17705,N_17985);
xnor U18105 (N_18105,N_17278,N_17810);
and U18106 (N_18106,N_17654,N_17204);
xor U18107 (N_18107,N_17446,N_17081);
xnor U18108 (N_18108,N_17509,N_17390);
xnor U18109 (N_18109,N_17179,N_17161);
or U18110 (N_18110,N_17024,N_17475);
xor U18111 (N_18111,N_17100,N_17613);
xnor U18112 (N_18112,N_17087,N_17374);
xnor U18113 (N_18113,N_17241,N_17305);
or U18114 (N_18114,N_17899,N_17597);
nand U18115 (N_18115,N_17564,N_17783);
nand U18116 (N_18116,N_17061,N_17090);
nand U18117 (N_18117,N_17500,N_17757);
xnor U18118 (N_18118,N_17918,N_17527);
xnor U18119 (N_18119,N_17267,N_17199);
nor U18120 (N_18120,N_17215,N_17124);
and U18121 (N_18121,N_17768,N_17703);
nand U18122 (N_18122,N_17667,N_17521);
xnor U18123 (N_18123,N_17970,N_17625);
nand U18124 (N_18124,N_17273,N_17690);
xnor U18125 (N_18125,N_17563,N_17955);
and U18126 (N_18126,N_17084,N_17458);
xnor U18127 (N_18127,N_17932,N_17078);
and U18128 (N_18128,N_17335,N_17980);
xor U18129 (N_18129,N_17714,N_17949);
nor U18130 (N_18130,N_17849,N_17280);
and U18131 (N_18131,N_17375,N_17550);
nor U18132 (N_18132,N_17186,N_17343);
or U18133 (N_18133,N_17042,N_17608);
xor U18134 (N_18134,N_17788,N_17047);
or U18135 (N_18135,N_17942,N_17812);
nor U18136 (N_18136,N_17126,N_17928);
xor U18137 (N_18137,N_17447,N_17300);
nor U18138 (N_18138,N_17953,N_17693);
nand U18139 (N_18139,N_17709,N_17666);
xnor U18140 (N_18140,N_17825,N_17276);
or U18141 (N_18141,N_17439,N_17088);
nor U18142 (N_18142,N_17622,N_17141);
nand U18143 (N_18143,N_17878,N_17606);
and U18144 (N_18144,N_17984,N_17822);
and U18145 (N_18145,N_17683,N_17197);
xor U18146 (N_18146,N_17961,N_17497);
nor U18147 (N_18147,N_17407,N_17903);
xnor U18148 (N_18148,N_17847,N_17428);
nand U18149 (N_18149,N_17412,N_17232);
or U18150 (N_18150,N_17292,N_17960);
xor U18151 (N_18151,N_17525,N_17454);
nand U18152 (N_18152,N_17321,N_17720);
or U18153 (N_18153,N_17003,N_17626);
and U18154 (N_18154,N_17784,N_17346);
xnor U18155 (N_18155,N_17162,N_17601);
or U18156 (N_18156,N_17806,N_17520);
nand U18157 (N_18157,N_17307,N_17262);
nor U18158 (N_18158,N_17726,N_17761);
nor U18159 (N_18159,N_17408,N_17702);
xnor U18160 (N_18160,N_17422,N_17995);
xnor U18161 (N_18161,N_17132,N_17368);
xor U18162 (N_18162,N_17930,N_17399);
or U18163 (N_18163,N_17184,N_17330);
or U18164 (N_18164,N_17093,N_17191);
and U18165 (N_18165,N_17740,N_17175);
xnor U18166 (N_18166,N_17461,N_17313);
nor U18167 (N_18167,N_17117,N_17118);
nor U18168 (N_18168,N_17202,N_17209);
or U18169 (N_18169,N_17163,N_17587);
or U18170 (N_18170,N_17687,N_17999);
xor U18171 (N_18171,N_17006,N_17778);
nand U18172 (N_18172,N_17239,N_17261);
and U18173 (N_18173,N_17397,N_17018);
nand U18174 (N_18174,N_17460,N_17157);
nor U18175 (N_18175,N_17640,N_17317);
and U18176 (N_18176,N_17680,N_17531);
and U18177 (N_18177,N_17638,N_17602);
or U18178 (N_18178,N_17325,N_17424);
or U18179 (N_18179,N_17701,N_17340);
nor U18180 (N_18180,N_17908,N_17263);
nor U18181 (N_18181,N_17518,N_17334);
nand U18182 (N_18182,N_17577,N_17190);
or U18183 (N_18183,N_17410,N_17376);
or U18184 (N_18184,N_17320,N_17712);
nor U18185 (N_18185,N_17870,N_17886);
nand U18186 (N_18186,N_17554,N_17893);
nor U18187 (N_18187,N_17229,N_17839);
and U18188 (N_18188,N_17245,N_17448);
xnor U18189 (N_18189,N_17674,N_17356);
or U18190 (N_18190,N_17324,N_17901);
or U18191 (N_18191,N_17384,N_17533);
nand U18192 (N_18192,N_17698,N_17871);
or U18193 (N_18193,N_17880,N_17694);
or U18194 (N_18194,N_17989,N_17008);
nand U18195 (N_18195,N_17844,N_17296);
xnor U18196 (N_18196,N_17430,N_17515);
and U18197 (N_18197,N_17056,N_17127);
or U18198 (N_18198,N_17028,N_17544);
or U18199 (N_18199,N_17939,N_17105);
or U18200 (N_18200,N_17897,N_17635);
nor U18201 (N_18201,N_17025,N_17836);
or U18202 (N_18202,N_17426,N_17467);
and U18203 (N_18203,N_17583,N_17851);
and U18204 (N_18204,N_17392,N_17243);
xnor U18205 (N_18205,N_17957,N_17786);
or U18206 (N_18206,N_17470,N_17145);
or U18207 (N_18207,N_17748,N_17297);
xor U18208 (N_18208,N_17629,N_17831);
or U18209 (N_18209,N_17121,N_17095);
or U18210 (N_18210,N_17233,N_17109);
and U18211 (N_18211,N_17843,N_17920);
and U18212 (N_18212,N_17417,N_17315);
and U18213 (N_18213,N_17616,N_17183);
nand U18214 (N_18214,N_17045,N_17991);
nor U18215 (N_18215,N_17845,N_17776);
and U18216 (N_18216,N_17814,N_17473);
and U18217 (N_18217,N_17755,N_17639);
nor U18218 (N_18218,N_17576,N_17620);
nand U18219 (N_18219,N_17743,N_17455);
and U18220 (N_18220,N_17840,N_17826);
xnor U18221 (N_18221,N_17919,N_17859);
and U18222 (N_18222,N_17348,N_17394);
or U18223 (N_18223,N_17442,N_17492);
xor U18224 (N_18224,N_17506,N_17079);
or U18225 (N_18225,N_17609,N_17436);
and U18226 (N_18226,N_17742,N_17972);
or U18227 (N_18227,N_17043,N_17434);
xor U18228 (N_18228,N_17062,N_17504);
and U18229 (N_18229,N_17350,N_17538);
xor U18230 (N_18230,N_17754,N_17264);
nor U18231 (N_18231,N_17354,N_17026);
xor U18232 (N_18232,N_17553,N_17708);
or U18233 (N_18233,N_17503,N_17598);
or U18234 (N_18234,N_17242,N_17231);
nor U18235 (N_18235,N_17944,N_17283);
nor U18236 (N_18236,N_17827,N_17207);
nand U18237 (N_18237,N_17612,N_17913);
or U18238 (N_18238,N_17567,N_17771);
xnor U18239 (N_18239,N_17050,N_17072);
nor U18240 (N_18240,N_17173,N_17811);
nand U18241 (N_18241,N_17803,N_17107);
nand U18242 (N_18242,N_17302,N_17060);
and U18243 (N_18243,N_17160,N_17438);
nor U18244 (N_18244,N_17716,N_17007);
xnor U18245 (N_18245,N_17772,N_17660);
nand U18246 (N_18246,N_17857,N_17332);
xor U18247 (N_18247,N_17338,N_17096);
or U18248 (N_18248,N_17339,N_17753);
and U18249 (N_18249,N_17744,N_17707);
nand U18250 (N_18250,N_17522,N_17166);
or U18251 (N_18251,N_17352,N_17221);
nand U18252 (N_18252,N_17479,N_17294);
nand U18253 (N_18253,N_17910,N_17185);
nor U18254 (N_18254,N_17572,N_17935);
or U18255 (N_18255,N_17734,N_17398);
nor U18256 (N_18256,N_17167,N_17059);
xnor U18257 (N_18257,N_17990,N_17240);
xnor U18258 (N_18258,N_17465,N_17632);
or U18259 (N_18259,N_17485,N_17976);
or U18260 (N_18260,N_17429,N_17615);
or U18261 (N_18261,N_17456,N_17415);
nor U18262 (N_18262,N_17152,N_17936);
nand U18263 (N_18263,N_17728,N_17568);
or U18264 (N_18264,N_17551,N_17931);
and U18265 (N_18265,N_17057,N_17435);
and U18266 (N_18266,N_17865,N_17481);
nor U18267 (N_18267,N_17528,N_17765);
nor U18268 (N_18268,N_17692,N_17604);
nor U18269 (N_18269,N_17891,N_17719);
nand U18270 (N_18270,N_17271,N_17592);
nor U18271 (N_18271,N_17361,N_17382);
xor U18272 (N_18272,N_17345,N_17174);
nand U18273 (N_18273,N_17083,N_17792);
and U18274 (N_18274,N_17926,N_17766);
xor U18275 (N_18275,N_17070,N_17385);
and U18276 (N_18276,N_17303,N_17466);
or U18277 (N_18277,N_17097,N_17732);
and U18278 (N_18278,N_17066,N_17663);
xnor U18279 (N_18279,N_17459,N_17219);
or U18280 (N_18280,N_17925,N_17293);
xnor U18281 (N_18281,N_17206,N_17055);
nor U18282 (N_18282,N_17982,N_17002);
and U18283 (N_18283,N_17902,N_17787);
or U18284 (N_18284,N_17427,N_17881);
nand U18285 (N_18285,N_17963,N_17706);
xnor U18286 (N_18286,N_17889,N_17074);
and U18287 (N_18287,N_17696,N_17112);
xnor U18288 (N_18288,N_17679,N_17850);
nand U18289 (N_18289,N_17943,N_17907);
nand U18290 (N_18290,N_17967,N_17443);
nand U18291 (N_18291,N_17634,N_17611);
nor U18292 (N_18292,N_17071,N_17180);
or U18293 (N_18293,N_17879,N_17051);
or U18294 (N_18294,N_17678,N_17432);
nand U18295 (N_18295,N_17248,N_17020);
or U18296 (N_18296,N_17565,N_17717);
or U18297 (N_18297,N_17182,N_17569);
xnor U18298 (N_18298,N_17673,N_17349);
and U18299 (N_18299,N_17861,N_17364);
nand U18300 (N_18300,N_17981,N_17883);
nand U18301 (N_18301,N_17973,N_17134);
nor U18302 (N_18302,N_17780,N_17951);
xnor U18303 (N_18303,N_17733,N_17449);
and U18304 (N_18304,N_17536,N_17624);
nor U18305 (N_18305,N_17829,N_17556);
nand U18306 (N_18306,N_17158,N_17165);
nand U18307 (N_18307,N_17237,N_17725);
nand U18308 (N_18308,N_17511,N_17782);
nor U18309 (N_18309,N_17494,N_17181);
and U18310 (N_18310,N_17268,N_17146);
or U18311 (N_18311,N_17617,N_17979);
nor U18312 (N_18312,N_17476,N_17519);
nand U18313 (N_18313,N_17274,N_17213);
nor U18314 (N_18314,N_17662,N_17013);
and U18315 (N_18315,N_17774,N_17402);
nor U18316 (N_18316,N_17370,N_17381);
nor U18317 (N_18317,N_17058,N_17425);
or U18318 (N_18318,N_17488,N_17017);
xnor U18319 (N_18319,N_17646,N_17882);
or U18320 (N_18320,N_17128,N_17453);
and U18321 (N_18321,N_17194,N_17781);
nor U18322 (N_18322,N_17418,N_17393);
nand U18323 (N_18323,N_17762,N_17866);
nand U18324 (N_18324,N_17965,N_17220);
and U18325 (N_18325,N_17805,N_17669);
nand U18326 (N_18326,N_17212,N_17790);
and U18327 (N_18327,N_17539,N_17021);
nor U18328 (N_18328,N_17763,N_17308);
and U18329 (N_18329,N_17421,N_17594);
nand U18330 (N_18330,N_17218,N_17691);
and U18331 (N_18331,N_17824,N_17760);
and U18332 (N_18332,N_17956,N_17828);
and U18333 (N_18333,N_17208,N_17380);
and U18334 (N_18334,N_17543,N_17954);
xnor U18335 (N_18335,N_17775,N_17929);
and U18336 (N_18336,N_17801,N_17791);
or U18337 (N_18337,N_17695,N_17914);
nand U18338 (N_18338,N_17715,N_17977);
xor U18339 (N_18339,N_17478,N_17288);
nor U18340 (N_18340,N_17941,N_17721);
xor U18341 (N_18341,N_17049,N_17144);
or U18342 (N_18342,N_17773,N_17195);
xor U18343 (N_18343,N_17033,N_17281);
and U18344 (N_18344,N_17210,N_17934);
or U18345 (N_18345,N_17286,N_17012);
or U18346 (N_18346,N_17498,N_17863);
nand U18347 (N_18347,N_17796,N_17636);
nand U18348 (N_18348,N_17360,N_17188);
xnor U18349 (N_18349,N_17759,N_17962);
and U18350 (N_18350,N_17489,N_17030);
nand U18351 (N_18351,N_17987,N_17187);
and U18352 (N_18352,N_17499,N_17894);
and U18353 (N_18353,N_17852,N_17189);
nor U18354 (N_18354,N_17655,N_17154);
and U18355 (N_18355,N_17820,N_17203);
xor U18356 (N_18356,N_17214,N_17041);
nor U18357 (N_18357,N_17004,N_17514);
nor U18358 (N_18358,N_17833,N_17659);
nor U18359 (N_18359,N_17073,N_17988);
xor U18360 (N_18360,N_17600,N_17978);
and U18361 (N_18361,N_17672,N_17336);
nor U18362 (N_18362,N_17737,N_17406);
xor U18363 (N_18363,N_17486,N_17272);
nor U18364 (N_18364,N_17395,N_17474);
nand U18365 (N_18365,N_17596,N_17400);
or U18366 (N_18366,N_17546,N_17923);
nor U18367 (N_18367,N_17357,N_17319);
nand U18368 (N_18368,N_17275,N_17477);
xor U18369 (N_18369,N_17177,N_17316);
and U18370 (N_18370,N_17676,N_17223);
nor U18371 (N_18371,N_17911,N_17589);
nand U18372 (N_18372,N_17524,N_17605);
nor U18373 (N_18373,N_17888,N_17585);
nand U18374 (N_18374,N_17142,N_17046);
or U18375 (N_18375,N_17201,N_17054);
or U18376 (N_18376,N_17329,N_17657);
xor U18377 (N_18377,N_17064,N_17647);
nand U18378 (N_18378,N_17656,N_17670);
xnor U18379 (N_18379,N_17362,N_17917);
nor U18380 (N_18380,N_17750,N_17289);
and U18381 (N_18381,N_17366,N_17063);
xnor U18382 (N_18382,N_17651,N_17298);
xnor U18383 (N_18383,N_17747,N_17076);
xnor U18384 (N_18384,N_17603,N_17085);
or U18385 (N_18385,N_17103,N_17713);
or U18386 (N_18386,N_17129,N_17147);
xnor U18387 (N_18387,N_17413,N_17628);
nand U18388 (N_18388,N_17619,N_17140);
xnor U18389 (N_18389,N_17623,N_17411);
or U18390 (N_18390,N_17252,N_17875);
or U18391 (N_18391,N_17143,N_17779);
or U18392 (N_18392,N_17529,N_17016);
and U18393 (N_18393,N_17794,N_17584);
nor U18394 (N_18394,N_17253,N_17178);
nor U18395 (N_18395,N_17574,N_17069);
and U18396 (N_18396,N_17785,N_17668);
or U18397 (N_18397,N_17222,N_17358);
nor U18398 (N_18398,N_17958,N_17120);
nand U18399 (N_18399,N_17699,N_17440);
nand U18400 (N_18400,N_17637,N_17948);
nand U18401 (N_18401,N_17685,N_17052);
and U18402 (N_18402,N_17916,N_17945);
xor U18403 (N_18403,N_17075,N_17727);
nor U18404 (N_18404,N_17704,N_17135);
nor U18405 (N_18405,N_17284,N_17710);
or U18406 (N_18406,N_17388,N_17793);
nor U18407 (N_18407,N_17688,N_17807);
nor U18408 (N_18408,N_17102,N_17819);
or U18409 (N_18409,N_17159,N_17010);
nand U18410 (N_18410,N_17260,N_17590);
xor U18411 (N_18411,N_17547,N_17139);
nand U18412 (N_18412,N_17631,N_17854);
or U18413 (N_18413,N_17311,N_17310);
nand U18414 (N_18414,N_17968,N_17813);
nand U18415 (N_18415,N_17344,N_17777);
or U18416 (N_18416,N_17595,N_17552);
nand U18417 (N_18417,N_17675,N_17838);
xnor U18418 (N_18418,N_17764,N_17414);
nand U18419 (N_18419,N_17082,N_17337);
nand U18420 (N_18420,N_17643,N_17257);
or U18421 (N_18421,N_17495,N_17892);
nand U18422 (N_18422,N_17169,N_17633);
xor U18423 (N_18423,N_17039,N_17573);
nand U18424 (N_18424,N_17974,N_17282);
nand U18425 (N_18425,N_17472,N_17718);
nand U18426 (N_18426,N_17513,N_17450);
xnor U18427 (N_18427,N_17798,N_17464);
xnor U18428 (N_18428,N_17722,N_17992);
nor U18429 (N_18429,N_17580,N_17947);
or U18430 (N_18430,N_17752,N_17516);
nand U18431 (N_18431,N_17031,N_17099);
and U18432 (N_18432,N_17022,N_17098);
nand U18433 (N_18433,N_17372,N_17815);
xor U18434 (N_18434,N_17092,N_17379);
nor U18435 (N_18435,N_17318,N_17614);
nor U18436 (N_18436,N_17876,N_17224);
nor U18437 (N_18437,N_17700,N_17559);
or U18438 (N_18438,N_17193,N_17797);
xnor U18439 (N_18439,N_17933,N_17285);
nor U18440 (N_18440,N_17172,N_17749);
nand U18441 (N_18441,N_17745,N_17015);
nor U18442 (N_18442,N_17034,N_17130);
xnor U18443 (N_18443,N_17153,N_17906);
and U18444 (N_18444,N_17451,N_17711);
or U18445 (N_18445,N_17420,N_17909);
or U18446 (N_18446,N_17226,N_17246);
xnor U18447 (N_18447,N_17419,N_17998);
nand U18448 (N_18448,N_17993,N_17848);
and U18449 (N_18449,N_17094,N_17480);
or U18450 (N_18450,N_17247,N_17053);
and U18451 (N_18451,N_17227,N_17830);
xnor U18452 (N_18452,N_17080,N_17331);
xor U18453 (N_18453,N_17523,N_17648);
or U18454 (N_18454,N_17562,N_17217);
or U18455 (N_18455,N_17869,N_17106);
xor U18456 (N_18456,N_17176,N_17689);
xor U18457 (N_18457,N_17867,N_17541);
or U18458 (N_18458,N_17490,N_17471);
and U18459 (N_18459,N_17255,N_17915);
and U18460 (N_18460,N_17036,N_17571);
and U18461 (N_18461,N_17037,N_17969);
nor U18462 (N_18462,N_17291,N_17483);
xor U18463 (N_18463,N_17645,N_17230);
nand U18464 (N_18464,N_17389,N_17873);
nor U18465 (N_18465,N_17196,N_17327);
nor U18466 (N_18466,N_17966,N_17534);
nor U18467 (N_18467,N_17618,N_17560);
and U18468 (N_18468,N_17116,N_17816);
nand U18469 (N_18469,N_17877,N_17029);
nand U18470 (N_18470,N_17168,N_17005);
nor U18471 (N_18471,N_17009,N_17457);
nor U18472 (N_18472,N_17650,N_17874);
xor U18473 (N_18473,N_17952,N_17986);
nor U18474 (N_18474,N_17496,N_17164);
xnor U18475 (N_18475,N_17858,N_17468);
and U18476 (N_18476,N_17040,N_17355);
nor U18477 (N_18477,N_17265,N_17996);
and U18478 (N_18478,N_17677,N_17502);
xnor U18479 (N_18479,N_17769,N_17014);
or U18480 (N_18480,N_17266,N_17946);
nor U18481 (N_18481,N_17746,N_17482);
or U18482 (N_18482,N_17347,N_17557);
nor U18483 (N_18483,N_17905,N_17855);
or U18484 (N_18484,N_17378,N_17860);
nor U18485 (N_18485,N_17735,N_17570);
nor U18486 (N_18486,N_17975,N_17809);
or U18487 (N_18487,N_17599,N_17171);
or U18488 (N_18488,N_17200,N_17835);
xor U18489 (N_18489,N_17369,N_17697);
and U18490 (N_18490,N_17301,N_17770);
or U18491 (N_18491,N_17823,N_17101);
nor U18492 (N_18492,N_17588,N_17148);
or U18493 (N_18493,N_17652,N_17610);
or U18494 (N_18494,N_17068,N_17799);
nand U18495 (N_18495,N_17751,N_17896);
or U18496 (N_18496,N_17270,N_17510);
nand U18497 (N_18497,N_17864,N_17731);
and U18498 (N_18498,N_17309,N_17328);
nand U18499 (N_18499,N_17125,N_17032);
and U18500 (N_18500,N_17327,N_17186);
or U18501 (N_18501,N_17062,N_17933);
and U18502 (N_18502,N_17207,N_17798);
nor U18503 (N_18503,N_17568,N_17553);
xnor U18504 (N_18504,N_17639,N_17515);
and U18505 (N_18505,N_17989,N_17524);
xor U18506 (N_18506,N_17690,N_17183);
nand U18507 (N_18507,N_17963,N_17364);
and U18508 (N_18508,N_17553,N_17567);
and U18509 (N_18509,N_17465,N_17844);
xor U18510 (N_18510,N_17366,N_17305);
or U18511 (N_18511,N_17303,N_17618);
nor U18512 (N_18512,N_17715,N_17180);
nor U18513 (N_18513,N_17031,N_17597);
nand U18514 (N_18514,N_17497,N_17551);
or U18515 (N_18515,N_17163,N_17517);
nand U18516 (N_18516,N_17917,N_17343);
nand U18517 (N_18517,N_17242,N_17971);
or U18518 (N_18518,N_17281,N_17515);
xnor U18519 (N_18519,N_17464,N_17724);
or U18520 (N_18520,N_17604,N_17886);
nand U18521 (N_18521,N_17237,N_17290);
and U18522 (N_18522,N_17062,N_17555);
xnor U18523 (N_18523,N_17650,N_17269);
or U18524 (N_18524,N_17481,N_17846);
and U18525 (N_18525,N_17693,N_17128);
nand U18526 (N_18526,N_17923,N_17696);
nand U18527 (N_18527,N_17949,N_17106);
nand U18528 (N_18528,N_17555,N_17778);
or U18529 (N_18529,N_17287,N_17733);
nor U18530 (N_18530,N_17174,N_17826);
nand U18531 (N_18531,N_17019,N_17543);
and U18532 (N_18532,N_17306,N_17934);
xnor U18533 (N_18533,N_17324,N_17018);
nor U18534 (N_18534,N_17790,N_17881);
or U18535 (N_18535,N_17423,N_17320);
xnor U18536 (N_18536,N_17742,N_17272);
xnor U18537 (N_18537,N_17149,N_17121);
nor U18538 (N_18538,N_17271,N_17549);
nor U18539 (N_18539,N_17313,N_17783);
nand U18540 (N_18540,N_17497,N_17236);
nor U18541 (N_18541,N_17171,N_17456);
and U18542 (N_18542,N_17690,N_17299);
or U18543 (N_18543,N_17496,N_17610);
xor U18544 (N_18544,N_17255,N_17392);
and U18545 (N_18545,N_17633,N_17486);
nor U18546 (N_18546,N_17316,N_17481);
nor U18547 (N_18547,N_17502,N_17192);
nor U18548 (N_18548,N_17661,N_17156);
xnor U18549 (N_18549,N_17385,N_17601);
and U18550 (N_18550,N_17299,N_17334);
or U18551 (N_18551,N_17763,N_17362);
or U18552 (N_18552,N_17244,N_17735);
nor U18553 (N_18553,N_17440,N_17023);
or U18554 (N_18554,N_17859,N_17598);
and U18555 (N_18555,N_17359,N_17585);
xor U18556 (N_18556,N_17156,N_17514);
xor U18557 (N_18557,N_17826,N_17441);
nand U18558 (N_18558,N_17524,N_17688);
xor U18559 (N_18559,N_17619,N_17057);
xnor U18560 (N_18560,N_17144,N_17991);
and U18561 (N_18561,N_17621,N_17652);
or U18562 (N_18562,N_17177,N_17365);
and U18563 (N_18563,N_17296,N_17072);
xnor U18564 (N_18564,N_17514,N_17554);
and U18565 (N_18565,N_17620,N_17211);
nor U18566 (N_18566,N_17326,N_17342);
and U18567 (N_18567,N_17737,N_17869);
and U18568 (N_18568,N_17434,N_17763);
xnor U18569 (N_18569,N_17886,N_17268);
nand U18570 (N_18570,N_17639,N_17546);
xnor U18571 (N_18571,N_17063,N_17722);
and U18572 (N_18572,N_17126,N_17163);
nand U18573 (N_18573,N_17017,N_17918);
nor U18574 (N_18574,N_17432,N_17058);
or U18575 (N_18575,N_17095,N_17524);
nand U18576 (N_18576,N_17737,N_17175);
xnor U18577 (N_18577,N_17959,N_17625);
and U18578 (N_18578,N_17524,N_17284);
nand U18579 (N_18579,N_17493,N_17803);
and U18580 (N_18580,N_17669,N_17923);
nand U18581 (N_18581,N_17699,N_17651);
and U18582 (N_18582,N_17528,N_17227);
nand U18583 (N_18583,N_17598,N_17225);
nand U18584 (N_18584,N_17479,N_17771);
nand U18585 (N_18585,N_17830,N_17782);
and U18586 (N_18586,N_17326,N_17266);
and U18587 (N_18587,N_17809,N_17120);
nand U18588 (N_18588,N_17454,N_17244);
or U18589 (N_18589,N_17739,N_17893);
xor U18590 (N_18590,N_17534,N_17844);
or U18591 (N_18591,N_17343,N_17612);
xnor U18592 (N_18592,N_17450,N_17408);
or U18593 (N_18593,N_17919,N_17982);
nor U18594 (N_18594,N_17765,N_17354);
nor U18595 (N_18595,N_17954,N_17524);
and U18596 (N_18596,N_17124,N_17569);
or U18597 (N_18597,N_17951,N_17587);
nand U18598 (N_18598,N_17814,N_17646);
nor U18599 (N_18599,N_17946,N_17243);
or U18600 (N_18600,N_17683,N_17048);
and U18601 (N_18601,N_17235,N_17331);
nand U18602 (N_18602,N_17505,N_17832);
nor U18603 (N_18603,N_17044,N_17349);
nand U18604 (N_18604,N_17487,N_17767);
xor U18605 (N_18605,N_17121,N_17300);
nor U18606 (N_18606,N_17218,N_17672);
xor U18607 (N_18607,N_17807,N_17583);
nand U18608 (N_18608,N_17683,N_17423);
xor U18609 (N_18609,N_17078,N_17148);
nand U18610 (N_18610,N_17033,N_17742);
xnor U18611 (N_18611,N_17184,N_17714);
xnor U18612 (N_18612,N_17324,N_17626);
xor U18613 (N_18613,N_17290,N_17738);
or U18614 (N_18614,N_17586,N_17926);
nand U18615 (N_18615,N_17045,N_17193);
or U18616 (N_18616,N_17644,N_17208);
nor U18617 (N_18617,N_17709,N_17365);
or U18618 (N_18618,N_17821,N_17786);
nor U18619 (N_18619,N_17982,N_17235);
and U18620 (N_18620,N_17900,N_17494);
and U18621 (N_18621,N_17792,N_17768);
nor U18622 (N_18622,N_17782,N_17764);
or U18623 (N_18623,N_17150,N_17095);
nor U18624 (N_18624,N_17019,N_17280);
or U18625 (N_18625,N_17598,N_17120);
xor U18626 (N_18626,N_17384,N_17315);
nand U18627 (N_18627,N_17221,N_17813);
nand U18628 (N_18628,N_17954,N_17544);
nand U18629 (N_18629,N_17044,N_17176);
and U18630 (N_18630,N_17963,N_17877);
and U18631 (N_18631,N_17566,N_17759);
and U18632 (N_18632,N_17656,N_17116);
nand U18633 (N_18633,N_17073,N_17839);
or U18634 (N_18634,N_17265,N_17428);
xor U18635 (N_18635,N_17726,N_17989);
nor U18636 (N_18636,N_17441,N_17171);
nor U18637 (N_18637,N_17708,N_17737);
and U18638 (N_18638,N_17421,N_17850);
nor U18639 (N_18639,N_17334,N_17600);
nand U18640 (N_18640,N_17132,N_17197);
and U18641 (N_18641,N_17651,N_17852);
or U18642 (N_18642,N_17834,N_17683);
xnor U18643 (N_18643,N_17986,N_17570);
or U18644 (N_18644,N_17188,N_17452);
nand U18645 (N_18645,N_17259,N_17870);
and U18646 (N_18646,N_17656,N_17642);
and U18647 (N_18647,N_17783,N_17222);
or U18648 (N_18648,N_17977,N_17142);
or U18649 (N_18649,N_17327,N_17382);
or U18650 (N_18650,N_17908,N_17481);
nand U18651 (N_18651,N_17320,N_17240);
nor U18652 (N_18652,N_17233,N_17485);
xnor U18653 (N_18653,N_17880,N_17279);
nand U18654 (N_18654,N_17474,N_17741);
and U18655 (N_18655,N_17248,N_17581);
and U18656 (N_18656,N_17048,N_17652);
or U18657 (N_18657,N_17992,N_17765);
xor U18658 (N_18658,N_17053,N_17324);
nand U18659 (N_18659,N_17735,N_17968);
nor U18660 (N_18660,N_17625,N_17415);
xnor U18661 (N_18661,N_17944,N_17818);
or U18662 (N_18662,N_17155,N_17312);
nand U18663 (N_18663,N_17655,N_17232);
xnor U18664 (N_18664,N_17927,N_17938);
nand U18665 (N_18665,N_17966,N_17976);
nor U18666 (N_18666,N_17145,N_17187);
and U18667 (N_18667,N_17302,N_17820);
xnor U18668 (N_18668,N_17721,N_17923);
xor U18669 (N_18669,N_17821,N_17888);
and U18670 (N_18670,N_17499,N_17200);
and U18671 (N_18671,N_17120,N_17647);
nor U18672 (N_18672,N_17017,N_17855);
nor U18673 (N_18673,N_17849,N_17510);
nand U18674 (N_18674,N_17228,N_17225);
or U18675 (N_18675,N_17119,N_17817);
xnor U18676 (N_18676,N_17435,N_17741);
or U18677 (N_18677,N_17769,N_17551);
nand U18678 (N_18678,N_17096,N_17747);
or U18679 (N_18679,N_17939,N_17921);
nor U18680 (N_18680,N_17805,N_17360);
nor U18681 (N_18681,N_17005,N_17629);
or U18682 (N_18682,N_17960,N_17434);
nand U18683 (N_18683,N_17144,N_17579);
nand U18684 (N_18684,N_17632,N_17035);
and U18685 (N_18685,N_17706,N_17727);
nor U18686 (N_18686,N_17320,N_17257);
nor U18687 (N_18687,N_17476,N_17758);
or U18688 (N_18688,N_17028,N_17640);
and U18689 (N_18689,N_17937,N_17566);
nand U18690 (N_18690,N_17589,N_17213);
nand U18691 (N_18691,N_17689,N_17112);
nor U18692 (N_18692,N_17683,N_17626);
nor U18693 (N_18693,N_17316,N_17279);
nor U18694 (N_18694,N_17579,N_17065);
and U18695 (N_18695,N_17501,N_17823);
or U18696 (N_18696,N_17118,N_17450);
or U18697 (N_18697,N_17959,N_17536);
or U18698 (N_18698,N_17501,N_17106);
and U18699 (N_18699,N_17898,N_17315);
or U18700 (N_18700,N_17413,N_17465);
nor U18701 (N_18701,N_17755,N_17291);
nand U18702 (N_18702,N_17457,N_17941);
nor U18703 (N_18703,N_17450,N_17718);
nand U18704 (N_18704,N_17346,N_17886);
nor U18705 (N_18705,N_17410,N_17190);
nor U18706 (N_18706,N_17458,N_17013);
xnor U18707 (N_18707,N_17316,N_17766);
nand U18708 (N_18708,N_17657,N_17331);
nand U18709 (N_18709,N_17853,N_17194);
nand U18710 (N_18710,N_17178,N_17565);
or U18711 (N_18711,N_17413,N_17132);
or U18712 (N_18712,N_17603,N_17333);
or U18713 (N_18713,N_17572,N_17975);
and U18714 (N_18714,N_17080,N_17328);
nand U18715 (N_18715,N_17704,N_17915);
nand U18716 (N_18716,N_17956,N_17550);
and U18717 (N_18717,N_17894,N_17405);
xnor U18718 (N_18718,N_17109,N_17958);
and U18719 (N_18719,N_17725,N_17972);
nand U18720 (N_18720,N_17776,N_17913);
and U18721 (N_18721,N_17432,N_17433);
xor U18722 (N_18722,N_17179,N_17805);
nor U18723 (N_18723,N_17211,N_17703);
nor U18724 (N_18724,N_17236,N_17766);
xnor U18725 (N_18725,N_17364,N_17687);
xnor U18726 (N_18726,N_17165,N_17253);
or U18727 (N_18727,N_17601,N_17012);
nand U18728 (N_18728,N_17617,N_17694);
nand U18729 (N_18729,N_17577,N_17015);
xor U18730 (N_18730,N_17134,N_17777);
xnor U18731 (N_18731,N_17563,N_17598);
xnor U18732 (N_18732,N_17978,N_17949);
and U18733 (N_18733,N_17072,N_17728);
and U18734 (N_18734,N_17757,N_17633);
xor U18735 (N_18735,N_17054,N_17402);
nand U18736 (N_18736,N_17518,N_17899);
and U18737 (N_18737,N_17102,N_17292);
and U18738 (N_18738,N_17123,N_17412);
nand U18739 (N_18739,N_17857,N_17402);
nand U18740 (N_18740,N_17512,N_17116);
nand U18741 (N_18741,N_17361,N_17521);
nand U18742 (N_18742,N_17789,N_17852);
nor U18743 (N_18743,N_17932,N_17978);
xor U18744 (N_18744,N_17758,N_17376);
xnor U18745 (N_18745,N_17295,N_17041);
xor U18746 (N_18746,N_17809,N_17617);
nor U18747 (N_18747,N_17029,N_17009);
and U18748 (N_18748,N_17956,N_17778);
xor U18749 (N_18749,N_17534,N_17360);
xor U18750 (N_18750,N_17449,N_17804);
nor U18751 (N_18751,N_17675,N_17159);
xor U18752 (N_18752,N_17967,N_17497);
nand U18753 (N_18753,N_17100,N_17826);
nand U18754 (N_18754,N_17877,N_17159);
nand U18755 (N_18755,N_17956,N_17271);
nor U18756 (N_18756,N_17369,N_17419);
xor U18757 (N_18757,N_17896,N_17174);
nand U18758 (N_18758,N_17616,N_17263);
and U18759 (N_18759,N_17855,N_17133);
or U18760 (N_18760,N_17789,N_17027);
nor U18761 (N_18761,N_17762,N_17227);
or U18762 (N_18762,N_17908,N_17975);
xor U18763 (N_18763,N_17869,N_17657);
xor U18764 (N_18764,N_17476,N_17901);
nand U18765 (N_18765,N_17354,N_17890);
nor U18766 (N_18766,N_17585,N_17136);
or U18767 (N_18767,N_17284,N_17532);
xnor U18768 (N_18768,N_17527,N_17004);
xor U18769 (N_18769,N_17515,N_17895);
and U18770 (N_18770,N_17384,N_17367);
and U18771 (N_18771,N_17407,N_17869);
nor U18772 (N_18772,N_17349,N_17129);
nand U18773 (N_18773,N_17944,N_17773);
xor U18774 (N_18774,N_17617,N_17504);
or U18775 (N_18775,N_17789,N_17386);
xnor U18776 (N_18776,N_17601,N_17605);
xor U18777 (N_18777,N_17526,N_17633);
nand U18778 (N_18778,N_17880,N_17962);
nand U18779 (N_18779,N_17431,N_17646);
nand U18780 (N_18780,N_17095,N_17117);
or U18781 (N_18781,N_17393,N_17375);
or U18782 (N_18782,N_17496,N_17604);
nand U18783 (N_18783,N_17750,N_17825);
nand U18784 (N_18784,N_17861,N_17028);
xnor U18785 (N_18785,N_17176,N_17976);
xnor U18786 (N_18786,N_17086,N_17318);
or U18787 (N_18787,N_17899,N_17305);
nor U18788 (N_18788,N_17187,N_17489);
and U18789 (N_18789,N_17849,N_17471);
and U18790 (N_18790,N_17179,N_17299);
nand U18791 (N_18791,N_17610,N_17616);
or U18792 (N_18792,N_17601,N_17559);
and U18793 (N_18793,N_17310,N_17323);
or U18794 (N_18794,N_17307,N_17806);
and U18795 (N_18795,N_17424,N_17861);
nand U18796 (N_18796,N_17166,N_17457);
or U18797 (N_18797,N_17553,N_17182);
or U18798 (N_18798,N_17491,N_17542);
or U18799 (N_18799,N_17665,N_17253);
and U18800 (N_18800,N_17390,N_17480);
nand U18801 (N_18801,N_17957,N_17881);
or U18802 (N_18802,N_17026,N_17972);
or U18803 (N_18803,N_17822,N_17343);
and U18804 (N_18804,N_17340,N_17197);
nor U18805 (N_18805,N_17606,N_17197);
xor U18806 (N_18806,N_17243,N_17447);
or U18807 (N_18807,N_17411,N_17662);
nand U18808 (N_18808,N_17251,N_17174);
nand U18809 (N_18809,N_17713,N_17017);
nand U18810 (N_18810,N_17852,N_17439);
nor U18811 (N_18811,N_17120,N_17753);
nor U18812 (N_18812,N_17178,N_17662);
xnor U18813 (N_18813,N_17098,N_17469);
xor U18814 (N_18814,N_17696,N_17864);
nand U18815 (N_18815,N_17412,N_17031);
nor U18816 (N_18816,N_17301,N_17992);
xor U18817 (N_18817,N_17452,N_17095);
xnor U18818 (N_18818,N_17980,N_17807);
nor U18819 (N_18819,N_17977,N_17570);
nor U18820 (N_18820,N_17170,N_17830);
nand U18821 (N_18821,N_17392,N_17561);
and U18822 (N_18822,N_17034,N_17828);
and U18823 (N_18823,N_17686,N_17671);
or U18824 (N_18824,N_17135,N_17582);
nor U18825 (N_18825,N_17141,N_17799);
nand U18826 (N_18826,N_17966,N_17075);
and U18827 (N_18827,N_17650,N_17129);
xnor U18828 (N_18828,N_17770,N_17852);
nand U18829 (N_18829,N_17426,N_17093);
nor U18830 (N_18830,N_17908,N_17024);
and U18831 (N_18831,N_17628,N_17721);
xnor U18832 (N_18832,N_17740,N_17531);
nand U18833 (N_18833,N_17718,N_17764);
or U18834 (N_18834,N_17922,N_17027);
or U18835 (N_18835,N_17433,N_17541);
and U18836 (N_18836,N_17532,N_17818);
nor U18837 (N_18837,N_17896,N_17755);
or U18838 (N_18838,N_17631,N_17937);
xnor U18839 (N_18839,N_17743,N_17009);
nand U18840 (N_18840,N_17613,N_17334);
nand U18841 (N_18841,N_17708,N_17421);
or U18842 (N_18842,N_17618,N_17986);
or U18843 (N_18843,N_17960,N_17778);
and U18844 (N_18844,N_17952,N_17348);
and U18845 (N_18845,N_17961,N_17673);
xnor U18846 (N_18846,N_17237,N_17315);
or U18847 (N_18847,N_17572,N_17873);
or U18848 (N_18848,N_17750,N_17474);
xnor U18849 (N_18849,N_17654,N_17731);
nand U18850 (N_18850,N_17003,N_17745);
or U18851 (N_18851,N_17229,N_17141);
and U18852 (N_18852,N_17804,N_17367);
nor U18853 (N_18853,N_17144,N_17406);
xor U18854 (N_18854,N_17318,N_17909);
and U18855 (N_18855,N_17754,N_17184);
and U18856 (N_18856,N_17989,N_17423);
nor U18857 (N_18857,N_17635,N_17087);
xnor U18858 (N_18858,N_17552,N_17849);
nor U18859 (N_18859,N_17035,N_17796);
xor U18860 (N_18860,N_17253,N_17818);
xor U18861 (N_18861,N_17873,N_17133);
or U18862 (N_18862,N_17142,N_17300);
xor U18863 (N_18863,N_17307,N_17015);
nand U18864 (N_18864,N_17499,N_17705);
or U18865 (N_18865,N_17866,N_17074);
nand U18866 (N_18866,N_17468,N_17788);
nand U18867 (N_18867,N_17388,N_17771);
xor U18868 (N_18868,N_17202,N_17547);
xnor U18869 (N_18869,N_17210,N_17477);
nor U18870 (N_18870,N_17414,N_17286);
nor U18871 (N_18871,N_17767,N_17500);
nand U18872 (N_18872,N_17982,N_17634);
nand U18873 (N_18873,N_17015,N_17687);
nor U18874 (N_18874,N_17624,N_17750);
nor U18875 (N_18875,N_17174,N_17675);
or U18876 (N_18876,N_17480,N_17724);
or U18877 (N_18877,N_17905,N_17102);
nor U18878 (N_18878,N_17064,N_17410);
nor U18879 (N_18879,N_17520,N_17002);
xor U18880 (N_18880,N_17999,N_17253);
and U18881 (N_18881,N_17591,N_17561);
xor U18882 (N_18882,N_17360,N_17745);
xor U18883 (N_18883,N_17751,N_17959);
nor U18884 (N_18884,N_17914,N_17245);
nand U18885 (N_18885,N_17700,N_17637);
or U18886 (N_18886,N_17777,N_17636);
and U18887 (N_18887,N_17963,N_17404);
or U18888 (N_18888,N_17547,N_17901);
nand U18889 (N_18889,N_17831,N_17975);
nor U18890 (N_18890,N_17299,N_17262);
and U18891 (N_18891,N_17840,N_17102);
and U18892 (N_18892,N_17793,N_17216);
nand U18893 (N_18893,N_17734,N_17240);
xnor U18894 (N_18894,N_17241,N_17539);
or U18895 (N_18895,N_17114,N_17537);
or U18896 (N_18896,N_17560,N_17600);
nand U18897 (N_18897,N_17832,N_17254);
xnor U18898 (N_18898,N_17784,N_17979);
and U18899 (N_18899,N_17831,N_17596);
xor U18900 (N_18900,N_17180,N_17827);
xor U18901 (N_18901,N_17780,N_17101);
or U18902 (N_18902,N_17847,N_17590);
or U18903 (N_18903,N_17085,N_17999);
xor U18904 (N_18904,N_17043,N_17585);
or U18905 (N_18905,N_17674,N_17847);
and U18906 (N_18906,N_17137,N_17404);
and U18907 (N_18907,N_17478,N_17467);
xnor U18908 (N_18908,N_17478,N_17816);
and U18909 (N_18909,N_17735,N_17838);
nor U18910 (N_18910,N_17171,N_17934);
nor U18911 (N_18911,N_17257,N_17107);
or U18912 (N_18912,N_17412,N_17325);
or U18913 (N_18913,N_17914,N_17517);
nand U18914 (N_18914,N_17095,N_17780);
nor U18915 (N_18915,N_17446,N_17285);
or U18916 (N_18916,N_17717,N_17185);
xor U18917 (N_18917,N_17804,N_17507);
nand U18918 (N_18918,N_17942,N_17577);
and U18919 (N_18919,N_17561,N_17060);
and U18920 (N_18920,N_17225,N_17661);
nand U18921 (N_18921,N_17391,N_17771);
nor U18922 (N_18922,N_17035,N_17991);
nor U18923 (N_18923,N_17113,N_17122);
nor U18924 (N_18924,N_17784,N_17536);
and U18925 (N_18925,N_17459,N_17802);
nand U18926 (N_18926,N_17981,N_17870);
nand U18927 (N_18927,N_17536,N_17193);
or U18928 (N_18928,N_17467,N_17835);
or U18929 (N_18929,N_17174,N_17383);
or U18930 (N_18930,N_17738,N_17441);
or U18931 (N_18931,N_17555,N_17922);
nand U18932 (N_18932,N_17918,N_17781);
nor U18933 (N_18933,N_17918,N_17272);
nand U18934 (N_18934,N_17871,N_17766);
or U18935 (N_18935,N_17230,N_17390);
and U18936 (N_18936,N_17940,N_17247);
and U18937 (N_18937,N_17409,N_17886);
nand U18938 (N_18938,N_17380,N_17100);
or U18939 (N_18939,N_17566,N_17793);
nand U18940 (N_18940,N_17453,N_17173);
xor U18941 (N_18941,N_17486,N_17916);
xnor U18942 (N_18942,N_17945,N_17600);
and U18943 (N_18943,N_17297,N_17551);
or U18944 (N_18944,N_17322,N_17975);
nor U18945 (N_18945,N_17240,N_17322);
or U18946 (N_18946,N_17712,N_17478);
xnor U18947 (N_18947,N_17588,N_17655);
nand U18948 (N_18948,N_17750,N_17662);
nand U18949 (N_18949,N_17948,N_17666);
nand U18950 (N_18950,N_17532,N_17727);
nor U18951 (N_18951,N_17920,N_17757);
or U18952 (N_18952,N_17533,N_17569);
xnor U18953 (N_18953,N_17196,N_17304);
nand U18954 (N_18954,N_17882,N_17638);
and U18955 (N_18955,N_17447,N_17644);
xnor U18956 (N_18956,N_17859,N_17696);
or U18957 (N_18957,N_17999,N_17236);
nor U18958 (N_18958,N_17660,N_17471);
and U18959 (N_18959,N_17236,N_17747);
nand U18960 (N_18960,N_17855,N_17620);
and U18961 (N_18961,N_17240,N_17495);
nand U18962 (N_18962,N_17421,N_17671);
or U18963 (N_18963,N_17075,N_17498);
and U18964 (N_18964,N_17701,N_17797);
xnor U18965 (N_18965,N_17576,N_17402);
or U18966 (N_18966,N_17490,N_17187);
or U18967 (N_18967,N_17548,N_17567);
and U18968 (N_18968,N_17474,N_17770);
xor U18969 (N_18969,N_17983,N_17845);
xnor U18970 (N_18970,N_17754,N_17358);
xnor U18971 (N_18971,N_17373,N_17701);
or U18972 (N_18972,N_17865,N_17518);
nand U18973 (N_18973,N_17163,N_17788);
nor U18974 (N_18974,N_17255,N_17469);
xor U18975 (N_18975,N_17160,N_17654);
or U18976 (N_18976,N_17722,N_17298);
nor U18977 (N_18977,N_17482,N_17854);
nand U18978 (N_18978,N_17029,N_17163);
or U18979 (N_18979,N_17770,N_17980);
xor U18980 (N_18980,N_17382,N_17270);
nor U18981 (N_18981,N_17718,N_17251);
nor U18982 (N_18982,N_17547,N_17244);
and U18983 (N_18983,N_17766,N_17158);
nor U18984 (N_18984,N_17107,N_17519);
and U18985 (N_18985,N_17774,N_17695);
nand U18986 (N_18986,N_17427,N_17166);
or U18987 (N_18987,N_17645,N_17188);
and U18988 (N_18988,N_17220,N_17962);
and U18989 (N_18989,N_17791,N_17152);
xnor U18990 (N_18990,N_17802,N_17030);
and U18991 (N_18991,N_17396,N_17788);
nand U18992 (N_18992,N_17928,N_17308);
nor U18993 (N_18993,N_17890,N_17869);
nand U18994 (N_18994,N_17246,N_17208);
nand U18995 (N_18995,N_17553,N_17414);
or U18996 (N_18996,N_17772,N_17990);
and U18997 (N_18997,N_17689,N_17770);
or U18998 (N_18998,N_17647,N_17327);
nor U18999 (N_18999,N_17040,N_17835);
or U19000 (N_19000,N_18185,N_18971);
nand U19001 (N_19001,N_18866,N_18047);
nand U19002 (N_19002,N_18074,N_18594);
nand U19003 (N_19003,N_18063,N_18716);
and U19004 (N_19004,N_18588,N_18407);
or U19005 (N_19005,N_18555,N_18893);
and U19006 (N_19006,N_18933,N_18108);
xnor U19007 (N_19007,N_18448,N_18714);
nand U19008 (N_19008,N_18348,N_18245);
or U19009 (N_19009,N_18042,N_18119);
nor U19010 (N_19010,N_18599,N_18331);
nor U19011 (N_19011,N_18600,N_18068);
nand U19012 (N_19012,N_18030,N_18373);
or U19013 (N_19013,N_18269,N_18831);
and U19014 (N_19014,N_18703,N_18051);
and U19015 (N_19015,N_18015,N_18697);
xnor U19016 (N_19016,N_18680,N_18718);
and U19017 (N_19017,N_18424,N_18295);
or U19018 (N_19018,N_18707,N_18136);
and U19019 (N_19019,N_18862,N_18694);
nand U19020 (N_19020,N_18853,N_18940);
nand U19021 (N_19021,N_18651,N_18539);
nor U19022 (N_19022,N_18398,N_18195);
nand U19023 (N_19023,N_18580,N_18918);
nand U19024 (N_19024,N_18548,N_18649);
xor U19025 (N_19025,N_18330,N_18067);
nand U19026 (N_19026,N_18957,N_18705);
nand U19027 (N_19027,N_18490,N_18762);
nand U19028 (N_19028,N_18550,N_18142);
or U19029 (N_19029,N_18568,N_18809);
or U19030 (N_19030,N_18652,N_18432);
nand U19031 (N_19031,N_18208,N_18537);
nand U19032 (N_19032,N_18477,N_18304);
and U19033 (N_19033,N_18668,N_18368);
xor U19034 (N_19034,N_18681,N_18271);
nand U19035 (N_19035,N_18754,N_18732);
or U19036 (N_19036,N_18571,N_18779);
or U19037 (N_19037,N_18184,N_18221);
xor U19038 (N_19038,N_18494,N_18527);
nand U19039 (N_19039,N_18766,N_18876);
xnor U19040 (N_19040,N_18531,N_18917);
nor U19041 (N_19041,N_18219,N_18929);
nor U19042 (N_19042,N_18370,N_18767);
nand U19043 (N_19043,N_18881,N_18238);
and U19044 (N_19044,N_18394,N_18510);
nor U19045 (N_19045,N_18518,N_18974);
xnor U19046 (N_19046,N_18909,N_18721);
nor U19047 (N_19047,N_18228,N_18105);
nand U19048 (N_19048,N_18521,N_18639);
nor U19049 (N_19049,N_18114,N_18196);
nand U19050 (N_19050,N_18376,N_18444);
nor U19051 (N_19051,N_18728,N_18653);
and U19052 (N_19052,N_18775,N_18073);
nor U19053 (N_19053,N_18798,N_18402);
nand U19054 (N_19054,N_18229,N_18225);
and U19055 (N_19055,N_18473,N_18043);
nand U19056 (N_19056,N_18606,N_18735);
nor U19057 (N_19057,N_18856,N_18936);
nand U19058 (N_19058,N_18272,N_18730);
and U19059 (N_19059,N_18204,N_18702);
xnor U19060 (N_19060,N_18602,N_18771);
nand U19061 (N_19061,N_18621,N_18144);
or U19062 (N_19062,N_18520,N_18834);
nor U19063 (N_19063,N_18815,N_18797);
and U19064 (N_19064,N_18495,N_18223);
nand U19065 (N_19065,N_18019,N_18146);
nand U19066 (N_19066,N_18554,N_18637);
nor U19067 (N_19067,N_18454,N_18158);
nand U19068 (N_19068,N_18317,N_18822);
and U19069 (N_19069,N_18266,N_18711);
or U19070 (N_19070,N_18596,N_18173);
xor U19071 (N_19071,N_18006,N_18143);
nand U19072 (N_19072,N_18032,N_18871);
and U19073 (N_19073,N_18590,N_18084);
and U19074 (N_19074,N_18787,N_18191);
nor U19075 (N_19075,N_18188,N_18870);
and U19076 (N_19076,N_18018,N_18608);
xnor U19077 (N_19077,N_18844,N_18041);
xnor U19078 (N_19078,N_18695,N_18461);
xor U19079 (N_19079,N_18906,N_18823);
and U19080 (N_19080,N_18827,N_18337);
and U19081 (N_19081,N_18632,N_18889);
or U19082 (N_19082,N_18855,N_18717);
and U19083 (N_19083,N_18701,N_18682);
nand U19084 (N_19084,N_18841,N_18115);
nor U19085 (N_19085,N_18215,N_18811);
nor U19086 (N_19086,N_18045,N_18462);
nand U19087 (N_19087,N_18489,N_18253);
xor U19088 (N_19088,N_18307,N_18848);
nor U19089 (N_19089,N_18300,N_18130);
nand U19090 (N_19090,N_18380,N_18562);
and U19091 (N_19091,N_18665,N_18077);
nand U19092 (N_19092,N_18891,N_18615);
and U19093 (N_19093,N_18127,N_18742);
nand U19094 (N_19094,N_18347,N_18968);
xnor U19095 (N_19095,N_18138,N_18340);
or U19096 (N_19096,N_18658,N_18626);
xor U19097 (N_19097,N_18022,N_18297);
and U19098 (N_19098,N_18670,N_18365);
nor U19099 (N_19099,N_18839,N_18913);
or U19100 (N_19100,N_18560,N_18507);
xnor U19101 (N_19101,N_18724,N_18328);
nand U19102 (N_19102,N_18515,N_18828);
nand U19103 (N_19103,N_18218,N_18401);
nand U19104 (N_19104,N_18178,N_18264);
nor U19105 (N_19105,N_18303,N_18847);
nand U19106 (N_19106,N_18542,N_18627);
nor U19107 (N_19107,N_18411,N_18984);
xnor U19108 (N_19108,N_18897,N_18120);
xor U19109 (N_19109,N_18796,N_18381);
xor U19110 (N_19110,N_18650,N_18291);
and U19111 (N_19111,N_18217,N_18082);
or U19112 (N_19112,N_18151,N_18288);
nand U19113 (N_19113,N_18430,N_18964);
nor U19114 (N_19114,N_18751,N_18688);
and U19115 (N_19115,N_18403,N_18799);
xnor U19116 (N_19116,N_18565,N_18321);
nor U19117 (N_19117,N_18165,N_18298);
xnor U19118 (N_19118,N_18546,N_18850);
xnor U19119 (N_19119,N_18311,N_18698);
xor U19120 (N_19120,N_18353,N_18131);
or U19121 (N_19121,N_18479,N_18433);
or U19122 (N_19122,N_18247,N_18982);
or U19123 (N_19123,N_18336,N_18469);
nor U19124 (N_19124,N_18122,N_18205);
and U19125 (N_19125,N_18179,N_18660);
nand U19126 (N_19126,N_18919,N_18176);
and U19127 (N_19127,N_18584,N_18960);
xnor U19128 (N_19128,N_18912,N_18369);
nor U19129 (N_19129,N_18020,N_18329);
and U19130 (N_19130,N_18991,N_18260);
and U19131 (N_19131,N_18686,N_18171);
nor U19132 (N_19132,N_18593,N_18493);
and U19133 (N_19133,N_18558,N_18687);
nand U19134 (N_19134,N_18039,N_18523);
xor U19135 (N_19135,N_18564,N_18814);
nand U19136 (N_19136,N_18782,N_18884);
or U19137 (N_19137,N_18121,N_18163);
and U19138 (N_19138,N_18172,N_18065);
nand U19139 (N_19139,N_18945,N_18090);
or U19140 (N_19140,N_18154,N_18877);
and U19141 (N_19141,N_18306,N_18609);
or U19142 (N_19142,N_18509,N_18858);
nand U19143 (N_19143,N_18922,N_18690);
or U19144 (N_19144,N_18296,N_18880);
xnor U19145 (N_19145,N_18374,N_18784);
xnor U19146 (N_19146,N_18943,N_18149);
nand U19147 (N_19147,N_18854,N_18315);
nor U19148 (N_19148,N_18046,N_18362);
or U19149 (N_19149,N_18852,N_18139);
nor U19150 (N_19150,N_18333,N_18569);
and U19151 (N_19151,N_18604,N_18955);
nand U19152 (N_19152,N_18801,N_18156);
and U19153 (N_19153,N_18794,N_18441);
nor U19154 (N_19154,N_18692,N_18976);
nor U19155 (N_19155,N_18375,N_18747);
xor U19156 (N_19156,N_18058,N_18464);
or U19157 (N_19157,N_18453,N_18617);
nor U19158 (N_19158,N_18780,N_18764);
nor U19159 (N_19159,N_18415,N_18693);
nand U19160 (N_19160,N_18981,N_18085);
or U19161 (N_19161,N_18646,N_18123);
nor U19162 (N_19162,N_18998,N_18174);
or U19163 (N_19163,N_18585,N_18110);
nor U19164 (N_19164,N_18807,N_18613);
xnor U19165 (N_19165,N_18384,N_18731);
nand U19166 (N_19166,N_18969,N_18706);
and U19167 (N_19167,N_18332,N_18426);
xor U19168 (N_19168,N_18544,N_18399);
and U19169 (N_19169,N_18416,N_18440);
and U19170 (N_19170,N_18258,N_18497);
or U19171 (N_19171,N_18220,N_18486);
xor U19172 (N_19172,N_18959,N_18704);
xor U19173 (N_19173,N_18610,N_18699);
and U19174 (N_19174,N_18805,N_18256);
xnor U19175 (N_19175,N_18713,N_18434);
nor U19176 (N_19176,N_18587,N_18285);
or U19177 (N_19177,N_18145,N_18001);
or U19178 (N_19178,N_18683,N_18791);
nand U19179 (N_19179,N_18476,N_18346);
or U19180 (N_19180,N_18124,N_18267);
and U19181 (N_19181,N_18289,N_18352);
and U19182 (N_19182,N_18201,N_18248);
xor U19183 (N_19183,N_18227,N_18182);
xnor U19184 (N_19184,N_18232,N_18935);
nand U19185 (N_19185,N_18339,N_18678);
or U19186 (N_19186,N_18103,N_18761);
nand U19187 (N_19187,N_18106,N_18508);
and U19188 (N_19188,N_18437,N_18563);
or U19189 (N_19189,N_18422,N_18206);
nor U19190 (N_19190,N_18979,N_18934);
or U19191 (N_19191,N_18010,N_18069);
or U19192 (N_19192,N_18236,N_18180);
nor U19193 (N_19193,N_18614,N_18710);
nand U19194 (N_19194,N_18098,N_18741);
nand U19195 (N_19195,N_18377,N_18886);
xor U19196 (N_19196,N_18684,N_18199);
nor U19197 (N_19197,N_18282,N_18418);
and U19198 (N_19198,N_18474,N_18349);
xnor U19199 (N_19199,N_18134,N_18391);
and U19200 (N_19200,N_18029,N_18159);
and U19201 (N_19201,N_18641,N_18715);
nand U19202 (N_19202,N_18107,N_18630);
and U19203 (N_19203,N_18985,N_18458);
nor U19204 (N_19204,N_18488,N_18958);
nand U19205 (N_19205,N_18659,N_18292);
xor U19206 (N_19206,N_18435,N_18900);
and U19207 (N_19207,N_18007,N_18233);
xor U19208 (N_19208,N_18412,N_18756);
xor U19209 (N_19209,N_18284,N_18150);
xor U19210 (N_19210,N_18733,N_18170);
or U19211 (N_19211,N_18186,N_18857);
and U19212 (N_19212,N_18746,N_18556);
xnor U19213 (N_19213,N_18427,N_18790);
and U19214 (N_19214,N_18089,N_18883);
nand U19215 (N_19215,N_18978,N_18005);
nand U19216 (N_19216,N_18002,N_18447);
or U19217 (N_19217,N_18419,N_18193);
nor U19218 (N_19218,N_18152,N_18091);
nand U19219 (N_19219,N_18483,N_18845);
and U19220 (N_19220,N_18319,N_18096);
or U19221 (N_19221,N_18765,N_18071);
and U19222 (N_19222,N_18318,N_18648);
nor U19223 (N_19223,N_18551,N_18977);
and U19224 (N_19224,N_18720,N_18663);
or U19225 (N_19225,N_18250,N_18946);
or U19226 (N_19226,N_18552,N_18950);
xnor U19227 (N_19227,N_18901,N_18343);
nand U19228 (N_19228,N_18803,N_18409);
or U19229 (N_19229,N_18287,N_18079);
nor U19230 (N_19230,N_18111,N_18334);
xor U19231 (N_19231,N_18363,N_18431);
and U19232 (N_19232,N_18017,N_18824);
and U19233 (N_19233,N_18719,N_18487);
xnor U19234 (N_19234,N_18953,N_18101);
or U19235 (N_19235,N_18070,N_18770);
xnor U19236 (N_19236,N_18522,N_18472);
xor U19237 (N_19237,N_18467,N_18470);
nor U19238 (N_19238,N_18169,N_18538);
or U19239 (N_19239,N_18664,N_18456);
nand U19240 (N_19240,N_18443,N_18025);
nor U19241 (N_19241,N_18438,N_18161);
nand U19242 (N_19242,N_18261,N_18983);
xnor U19243 (N_19243,N_18423,N_18601);
nand U19244 (N_19244,N_18400,N_18885);
nor U19245 (N_19245,N_18578,N_18168);
nor U19246 (N_19246,N_18502,N_18364);
or U19247 (N_19247,N_18988,N_18093);
nand U19248 (N_19248,N_18436,N_18956);
nand U19249 (N_19249,N_18605,N_18753);
nor U19250 (N_19250,N_18102,N_18278);
or U19251 (N_19251,N_18778,N_18576);
or U19252 (N_19252,N_18457,N_18194);
nor U19253 (N_19253,N_18583,N_18439);
nand U19254 (N_19254,N_18833,N_18887);
and U19255 (N_19255,N_18442,N_18942);
or U19256 (N_19256,N_18836,N_18361);
or U19257 (N_19257,N_18989,N_18760);
or U19258 (N_19258,N_18481,N_18994);
xnor U19259 (N_19259,N_18305,N_18390);
and U19260 (N_19260,N_18873,N_18410);
xnor U19261 (N_19261,N_18175,N_18057);
and U19262 (N_19262,N_18924,N_18244);
nand U19263 (N_19263,N_18446,N_18776);
nand U19264 (N_19264,N_18009,N_18820);
xnor U19265 (N_19265,N_18132,N_18449);
or U19266 (N_19266,N_18777,N_18072);
or U19267 (N_19267,N_18393,N_18000);
nand U19268 (N_19268,N_18125,N_18459);
nor U19269 (N_19269,N_18414,N_18624);
xnor U19270 (N_19270,N_18386,N_18890);
nand U19271 (N_19271,N_18997,N_18644);
nor U19272 (N_19272,N_18725,N_18902);
xor U19273 (N_19273,N_18092,N_18354);
nand U19274 (N_19274,N_18226,N_18314);
nand U19275 (N_19275,N_18620,N_18817);
and U19276 (N_19276,N_18758,N_18262);
nand U19277 (N_19277,N_18054,N_18972);
nor U19278 (N_19278,N_18903,N_18975);
and U19279 (N_19279,N_18948,N_18342);
and U19280 (N_19280,N_18781,N_18892);
nor U19281 (N_19281,N_18938,N_18635);
nor U19282 (N_19282,N_18265,N_18603);
nor U19283 (N_19283,N_18246,N_18597);
or U19284 (N_19284,N_18212,N_18530);
and U19285 (N_19285,N_18575,N_18743);
nand U19286 (N_19286,N_18094,N_18395);
or U19287 (N_19287,N_18869,N_18944);
nor U19288 (N_19288,N_18643,N_18155);
or U19289 (N_19289,N_18910,N_18750);
nand U19290 (N_19290,N_18048,N_18567);
xnor U19291 (N_19291,N_18053,N_18335);
nor U19292 (N_19292,N_18829,N_18358);
nand U19293 (N_19293,N_18177,N_18691);
or U19294 (N_19294,N_18749,N_18468);
nor U19295 (N_19295,N_18224,N_18534);
xor U19296 (N_19296,N_18579,N_18524);
nor U19297 (N_19297,N_18581,N_18372);
or U19298 (N_19298,N_18512,N_18478);
nand U19299 (N_19299,N_18928,N_18034);
nor U19300 (N_19300,N_18793,N_18612);
nand U19301 (N_19301,N_18216,N_18513);
or U19302 (N_19302,N_18939,N_18638);
nand U19303 (N_19303,N_18973,N_18965);
nor U19304 (N_19304,N_18677,N_18460);
and U19305 (N_19305,N_18506,N_18533);
nor U19306 (N_19306,N_18086,N_18843);
xnor U19307 (N_19307,N_18947,N_18345);
or U19308 (N_19308,N_18745,N_18417);
and U19309 (N_19309,N_18655,N_18726);
xnor U19310 (N_19310,N_18322,N_18408);
xor U19311 (N_19311,N_18813,N_18326);
and U19312 (N_19312,N_18842,N_18276);
nor U19313 (N_19313,N_18021,N_18389);
nor U19314 (N_19314,N_18341,N_18392);
xor U19315 (N_19315,N_18211,N_18657);
xnor U19316 (N_19316,N_18455,N_18190);
and U19317 (N_19317,N_18927,N_18385);
or U19318 (N_19318,N_18097,N_18806);
or U19319 (N_19319,N_18141,N_18181);
nand U19320 (N_19320,N_18421,N_18826);
nor U19321 (N_19321,N_18789,N_18859);
and U19322 (N_19322,N_18727,N_18148);
nor U19323 (N_19323,N_18214,N_18825);
and U19324 (N_19324,N_18874,N_18708);
or U19325 (N_19325,N_18081,N_18004);
xor U19326 (N_19326,N_18299,N_18656);
or U19327 (N_19327,N_18095,N_18905);
xor U19328 (N_19328,N_18553,N_18970);
or U19329 (N_19329,N_18954,N_18633);
xor U19330 (N_19330,N_18294,N_18485);
or U19331 (N_19331,N_18209,N_18252);
nor U19332 (N_19332,N_18273,N_18712);
nor U19333 (N_19333,N_18207,N_18323);
nor U19334 (N_19334,N_18259,N_18894);
and U19335 (N_19335,N_18290,N_18075);
and U19336 (N_19336,N_18709,N_18837);
nor U19337 (N_19337,N_18532,N_18033);
nor U19338 (N_19338,N_18768,N_18312);
xor U19339 (N_19339,N_18896,N_18672);
and U19340 (N_19340,N_18616,N_18044);
nor U19341 (N_19341,N_18099,N_18160);
nor U19342 (N_19342,N_18308,N_18310);
nand U19343 (N_19343,N_18202,N_18147);
nand U19344 (N_19344,N_18113,N_18203);
nor U19345 (N_19345,N_18952,N_18013);
and U19346 (N_19346,N_18722,N_18595);
nand U19347 (N_19347,N_18872,N_18541);
nor U19348 (N_19348,N_18559,N_18642);
or U19349 (N_19349,N_18925,N_18213);
xnor U19350 (N_19350,N_18367,N_18350);
xnor U19351 (N_19351,N_18235,N_18078);
xnor U19352 (N_19352,N_18838,N_18023);
or U19353 (N_19353,N_18230,N_18661);
nand U19354 (N_19354,N_18561,N_18519);
and U19355 (N_19355,N_18183,N_18028);
and U19356 (N_19356,N_18425,N_18325);
nand U19357 (N_19357,N_18254,N_18234);
and U19358 (N_19358,N_18008,N_18451);
xor U19359 (N_19359,N_18810,N_18257);
and U19360 (N_19360,N_18619,N_18625);
nor U19361 (N_19361,N_18198,N_18816);
xnor U19362 (N_19362,N_18937,N_18309);
and U19363 (N_19363,N_18623,N_18492);
or U19364 (N_19364,N_18066,N_18505);
nor U19365 (N_19365,N_18882,N_18355);
xor U19366 (N_19366,N_18274,N_18812);
and U19367 (N_19367,N_18986,N_18654);
nor U19368 (N_19368,N_18769,N_18240);
nand U19369 (N_19369,N_18062,N_18967);
or U19370 (N_19370,N_18821,N_18499);
nand U19371 (N_19371,N_18543,N_18878);
nor U19372 (N_19372,N_18237,N_18573);
nand U19373 (N_19373,N_18832,N_18961);
and U19374 (N_19374,N_18557,N_18445);
or U19375 (N_19375,N_18413,N_18526);
nor U19376 (N_19376,N_18126,N_18359);
nor U19377 (N_19377,N_18286,N_18050);
xnor U19378 (N_19378,N_18673,N_18669);
xor U19379 (N_19379,N_18491,N_18772);
nand U19380 (N_19380,N_18868,N_18049);
nand U19381 (N_19381,N_18420,N_18808);
and U19382 (N_19382,N_18990,N_18549);
xnor U19383 (N_19383,N_18923,N_18404);
xor U19384 (N_19384,N_18966,N_18275);
xor U19385 (N_19385,N_18031,N_18640);
or U19386 (N_19386,N_18327,N_18999);
nor U19387 (N_19387,N_18040,N_18366);
xor U19388 (N_19388,N_18572,N_18591);
nand U19389 (N_19389,N_18993,N_18995);
nor U19390 (N_19390,N_18429,N_18128);
nand U19391 (N_19391,N_18729,N_18773);
nor U19392 (N_19392,N_18759,N_18851);
nand U19393 (N_19393,N_18788,N_18503);
nand U19394 (N_19394,N_18496,N_18210);
nand U19395 (N_19395,N_18689,N_18428);
nand U19396 (N_19396,N_18525,N_18200);
nand U19397 (N_19397,N_18570,N_18344);
xnor U19398 (N_19398,N_18243,N_18574);
and U19399 (N_19399,N_18840,N_18739);
or U19400 (N_19400,N_18916,N_18511);
nand U19401 (N_19401,N_18313,N_18700);
nand U19402 (N_19402,N_18397,N_18338);
nor U19403 (N_19403,N_18647,N_18405);
and U19404 (N_19404,N_18498,N_18270);
nand U19405 (N_19405,N_18088,N_18675);
xnor U19406 (N_19406,N_18387,N_18501);
nand U19407 (N_19407,N_18802,N_18109);
nor U19408 (N_19408,N_18059,N_18586);
or U19409 (N_19409,N_18895,N_18915);
or U19410 (N_19410,N_18012,N_18582);
or U19411 (N_19411,N_18388,N_18117);
xor U19412 (N_19412,N_18835,N_18757);
or U19413 (N_19413,N_18011,N_18504);
xnor U19414 (N_19414,N_18536,N_18666);
or U19415 (N_19415,N_18083,N_18187);
xor U19416 (N_19416,N_18450,N_18949);
nand U19417 (N_19417,N_18293,N_18622);
and U19418 (N_19418,N_18135,N_18737);
nor U19419 (N_19419,N_18100,N_18951);
nand U19420 (N_19420,N_18819,N_18360);
or U19421 (N_19421,N_18056,N_18268);
or U19422 (N_19422,N_18566,N_18875);
and U19423 (N_19423,N_18133,N_18301);
and U19424 (N_19424,N_18904,N_18888);
or U19425 (N_19425,N_18351,N_18849);
nand U19426 (N_19426,N_18996,N_18785);
xnor U19427 (N_19427,N_18383,N_18104);
and U19428 (N_19428,N_18357,N_18679);
nor U19429 (N_19429,N_18898,N_18774);
nor U19430 (N_19430,N_18516,N_18723);
xnor U19431 (N_19431,N_18241,N_18861);
nor U19432 (N_19432,N_18752,N_18545);
nand U19433 (N_19433,N_18540,N_18197);
or U19434 (N_19434,N_18239,N_18899);
nand U19435 (N_19435,N_18060,N_18026);
and U19436 (N_19436,N_18055,N_18598);
or U19437 (N_19437,N_18645,N_18140);
xnor U19438 (N_19438,N_18744,N_18577);
or U19439 (N_19439,N_18396,N_18992);
or U19440 (N_19440,N_18003,N_18482);
nand U19441 (N_19441,N_18736,N_18980);
nor U19442 (N_19442,N_18676,N_18879);
xor U19443 (N_19443,N_18631,N_18763);
or U19444 (N_19444,N_18795,N_18281);
and U19445 (N_19445,N_18027,N_18076);
nand U19446 (N_19446,N_18465,N_18863);
nor U19447 (N_19447,N_18378,N_18471);
nor U19448 (N_19448,N_18356,N_18255);
or U19449 (N_19449,N_18517,N_18167);
xnor U19450 (N_19450,N_18911,N_18475);
and U19451 (N_19451,N_18222,N_18528);
nand U19452 (N_19452,N_18112,N_18607);
xnor U19453 (N_19453,N_18302,N_18907);
nand U19454 (N_19454,N_18251,N_18371);
xnor U19455 (N_19455,N_18037,N_18052);
nor U19456 (N_19456,N_18783,N_18864);
nor U19457 (N_19457,N_18466,N_18932);
or U19458 (N_19458,N_18786,N_18738);
nor U19459 (N_19459,N_18589,N_18036);
nor U19460 (N_19460,N_18634,N_18860);
nand U19461 (N_19461,N_18930,N_18189);
nor U19462 (N_19462,N_18324,N_18792);
or U19463 (N_19463,N_18164,N_18611);
nor U19464 (N_19464,N_18231,N_18463);
or U19465 (N_19465,N_18628,N_18064);
and U19466 (N_19466,N_18320,N_18667);
or U19467 (N_19467,N_18024,N_18116);
nand U19468 (N_19468,N_18500,N_18263);
xor U19469 (N_19469,N_18242,N_18192);
or U19470 (N_19470,N_18618,N_18908);
xnor U19471 (N_19471,N_18671,N_18316);
nand U19472 (N_19472,N_18035,N_18480);
xor U19473 (N_19473,N_18529,N_18283);
nand U19474 (N_19474,N_18734,N_18830);
nand U19475 (N_19475,N_18137,N_18514);
and U19476 (N_19476,N_18921,N_18129);
and U19477 (N_19477,N_18038,N_18685);
nor U19478 (N_19478,N_18941,N_18535);
or U19479 (N_19479,N_18061,N_18800);
xor U19480 (N_19480,N_18748,N_18740);
or U19481 (N_19481,N_18846,N_18920);
nor U19482 (N_19482,N_18484,N_18804);
nand U19483 (N_19483,N_18016,N_18629);
xnor U19484 (N_19484,N_18674,N_18926);
xnor U19485 (N_19485,N_18987,N_18867);
xnor U19486 (N_19486,N_18162,N_18865);
and U19487 (N_19487,N_18379,N_18962);
nand U19488 (N_19488,N_18452,N_18166);
nor U19489 (N_19489,N_18592,N_18636);
and U19490 (N_19490,N_18662,N_18157);
and U19491 (N_19491,N_18279,N_18931);
or U19492 (N_19492,N_18118,N_18382);
and U19493 (N_19493,N_18963,N_18014);
and U19494 (N_19494,N_18277,N_18406);
nand U19495 (N_19495,N_18249,N_18755);
and U19496 (N_19496,N_18696,N_18818);
nor U19497 (N_19497,N_18547,N_18087);
nand U19498 (N_19498,N_18153,N_18080);
nor U19499 (N_19499,N_18280,N_18914);
nand U19500 (N_19500,N_18301,N_18308);
xnor U19501 (N_19501,N_18053,N_18879);
nand U19502 (N_19502,N_18941,N_18612);
nand U19503 (N_19503,N_18841,N_18336);
nand U19504 (N_19504,N_18491,N_18174);
nor U19505 (N_19505,N_18145,N_18833);
xnor U19506 (N_19506,N_18606,N_18269);
nor U19507 (N_19507,N_18215,N_18708);
nor U19508 (N_19508,N_18539,N_18565);
xnor U19509 (N_19509,N_18549,N_18076);
nor U19510 (N_19510,N_18964,N_18867);
xnor U19511 (N_19511,N_18263,N_18446);
and U19512 (N_19512,N_18690,N_18400);
and U19513 (N_19513,N_18075,N_18246);
and U19514 (N_19514,N_18033,N_18686);
nor U19515 (N_19515,N_18590,N_18825);
nand U19516 (N_19516,N_18148,N_18424);
or U19517 (N_19517,N_18271,N_18228);
nand U19518 (N_19518,N_18101,N_18731);
xnor U19519 (N_19519,N_18402,N_18363);
nor U19520 (N_19520,N_18225,N_18823);
or U19521 (N_19521,N_18716,N_18181);
or U19522 (N_19522,N_18205,N_18438);
or U19523 (N_19523,N_18196,N_18235);
nor U19524 (N_19524,N_18484,N_18046);
xnor U19525 (N_19525,N_18887,N_18366);
or U19526 (N_19526,N_18625,N_18252);
xor U19527 (N_19527,N_18488,N_18239);
xnor U19528 (N_19528,N_18035,N_18825);
nand U19529 (N_19529,N_18259,N_18701);
xor U19530 (N_19530,N_18617,N_18534);
xnor U19531 (N_19531,N_18587,N_18119);
xor U19532 (N_19532,N_18695,N_18006);
xnor U19533 (N_19533,N_18208,N_18865);
or U19534 (N_19534,N_18110,N_18997);
nand U19535 (N_19535,N_18464,N_18328);
nand U19536 (N_19536,N_18001,N_18130);
and U19537 (N_19537,N_18859,N_18143);
and U19538 (N_19538,N_18743,N_18972);
nor U19539 (N_19539,N_18081,N_18845);
xor U19540 (N_19540,N_18788,N_18082);
xnor U19541 (N_19541,N_18051,N_18169);
or U19542 (N_19542,N_18863,N_18071);
nand U19543 (N_19543,N_18189,N_18571);
xnor U19544 (N_19544,N_18134,N_18841);
xor U19545 (N_19545,N_18865,N_18125);
and U19546 (N_19546,N_18463,N_18230);
nor U19547 (N_19547,N_18359,N_18793);
nand U19548 (N_19548,N_18090,N_18240);
nand U19549 (N_19549,N_18269,N_18825);
xnor U19550 (N_19550,N_18886,N_18908);
or U19551 (N_19551,N_18422,N_18402);
nor U19552 (N_19552,N_18300,N_18873);
xnor U19553 (N_19553,N_18733,N_18221);
nor U19554 (N_19554,N_18164,N_18301);
xor U19555 (N_19555,N_18180,N_18333);
xor U19556 (N_19556,N_18625,N_18079);
xnor U19557 (N_19557,N_18981,N_18396);
xnor U19558 (N_19558,N_18156,N_18947);
nand U19559 (N_19559,N_18793,N_18546);
and U19560 (N_19560,N_18215,N_18285);
and U19561 (N_19561,N_18768,N_18215);
nand U19562 (N_19562,N_18939,N_18682);
xor U19563 (N_19563,N_18123,N_18752);
or U19564 (N_19564,N_18091,N_18564);
and U19565 (N_19565,N_18934,N_18413);
or U19566 (N_19566,N_18026,N_18411);
xor U19567 (N_19567,N_18739,N_18492);
nand U19568 (N_19568,N_18587,N_18461);
nand U19569 (N_19569,N_18481,N_18949);
or U19570 (N_19570,N_18753,N_18689);
or U19571 (N_19571,N_18758,N_18187);
xor U19572 (N_19572,N_18206,N_18135);
and U19573 (N_19573,N_18393,N_18193);
nand U19574 (N_19574,N_18766,N_18900);
nor U19575 (N_19575,N_18285,N_18652);
xnor U19576 (N_19576,N_18040,N_18304);
and U19577 (N_19577,N_18444,N_18180);
nor U19578 (N_19578,N_18683,N_18962);
and U19579 (N_19579,N_18420,N_18635);
and U19580 (N_19580,N_18511,N_18977);
nand U19581 (N_19581,N_18452,N_18467);
xnor U19582 (N_19582,N_18627,N_18984);
xor U19583 (N_19583,N_18179,N_18324);
nand U19584 (N_19584,N_18225,N_18674);
nor U19585 (N_19585,N_18934,N_18412);
nand U19586 (N_19586,N_18783,N_18194);
or U19587 (N_19587,N_18326,N_18632);
xor U19588 (N_19588,N_18458,N_18087);
or U19589 (N_19589,N_18741,N_18931);
or U19590 (N_19590,N_18425,N_18871);
and U19591 (N_19591,N_18606,N_18088);
xnor U19592 (N_19592,N_18632,N_18123);
and U19593 (N_19593,N_18387,N_18313);
nand U19594 (N_19594,N_18894,N_18339);
nor U19595 (N_19595,N_18151,N_18939);
nor U19596 (N_19596,N_18326,N_18294);
nor U19597 (N_19597,N_18977,N_18515);
and U19598 (N_19598,N_18781,N_18111);
nand U19599 (N_19599,N_18917,N_18286);
nor U19600 (N_19600,N_18683,N_18919);
nor U19601 (N_19601,N_18833,N_18625);
nand U19602 (N_19602,N_18210,N_18520);
nor U19603 (N_19603,N_18615,N_18317);
or U19604 (N_19604,N_18035,N_18452);
xnor U19605 (N_19605,N_18078,N_18790);
or U19606 (N_19606,N_18129,N_18076);
or U19607 (N_19607,N_18724,N_18808);
and U19608 (N_19608,N_18474,N_18219);
and U19609 (N_19609,N_18880,N_18142);
nor U19610 (N_19610,N_18100,N_18144);
xnor U19611 (N_19611,N_18568,N_18529);
or U19612 (N_19612,N_18173,N_18913);
or U19613 (N_19613,N_18935,N_18394);
and U19614 (N_19614,N_18983,N_18100);
nor U19615 (N_19615,N_18432,N_18066);
xor U19616 (N_19616,N_18395,N_18624);
nand U19617 (N_19617,N_18162,N_18433);
or U19618 (N_19618,N_18976,N_18739);
nand U19619 (N_19619,N_18892,N_18443);
xor U19620 (N_19620,N_18413,N_18222);
or U19621 (N_19621,N_18931,N_18098);
xnor U19622 (N_19622,N_18601,N_18511);
nand U19623 (N_19623,N_18424,N_18970);
and U19624 (N_19624,N_18190,N_18688);
or U19625 (N_19625,N_18536,N_18817);
and U19626 (N_19626,N_18469,N_18684);
nor U19627 (N_19627,N_18526,N_18244);
nand U19628 (N_19628,N_18696,N_18842);
xor U19629 (N_19629,N_18060,N_18423);
nor U19630 (N_19630,N_18638,N_18983);
nor U19631 (N_19631,N_18637,N_18534);
or U19632 (N_19632,N_18438,N_18002);
or U19633 (N_19633,N_18747,N_18689);
xor U19634 (N_19634,N_18760,N_18235);
and U19635 (N_19635,N_18824,N_18574);
or U19636 (N_19636,N_18262,N_18955);
nor U19637 (N_19637,N_18376,N_18308);
xnor U19638 (N_19638,N_18039,N_18072);
and U19639 (N_19639,N_18837,N_18926);
nand U19640 (N_19640,N_18905,N_18491);
xnor U19641 (N_19641,N_18945,N_18893);
or U19642 (N_19642,N_18221,N_18565);
xor U19643 (N_19643,N_18909,N_18219);
or U19644 (N_19644,N_18850,N_18854);
xor U19645 (N_19645,N_18078,N_18172);
nand U19646 (N_19646,N_18432,N_18753);
nor U19647 (N_19647,N_18920,N_18278);
nand U19648 (N_19648,N_18531,N_18090);
or U19649 (N_19649,N_18500,N_18439);
and U19650 (N_19650,N_18517,N_18449);
xnor U19651 (N_19651,N_18752,N_18189);
nand U19652 (N_19652,N_18140,N_18915);
xor U19653 (N_19653,N_18600,N_18941);
or U19654 (N_19654,N_18594,N_18010);
nand U19655 (N_19655,N_18484,N_18890);
or U19656 (N_19656,N_18345,N_18856);
xor U19657 (N_19657,N_18678,N_18739);
nor U19658 (N_19658,N_18170,N_18756);
or U19659 (N_19659,N_18915,N_18684);
or U19660 (N_19660,N_18278,N_18057);
xnor U19661 (N_19661,N_18971,N_18047);
or U19662 (N_19662,N_18010,N_18083);
xor U19663 (N_19663,N_18054,N_18980);
or U19664 (N_19664,N_18857,N_18070);
or U19665 (N_19665,N_18086,N_18767);
nand U19666 (N_19666,N_18756,N_18916);
xor U19667 (N_19667,N_18625,N_18152);
nand U19668 (N_19668,N_18560,N_18649);
or U19669 (N_19669,N_18957,N_18258);
or U19670 (N_19670,N_18628,N_18631);
or U19671 (N_19671,N_18807,N_18365);
xnor U19672 (N_19672,N_18468,N_18130);
or U19673 (N_19673,N_18417,N_18049);
nand U19674 (N_19674,N_18137,N_18398);
or U19675 (N_19675,N_18667,N_18627);
and U19676 (N_19676,N_18647,N_18887);
and U19677 (N_19677,N_18467,N_18208);
and U19678 (N_19678,N_18742,N_18844);
and U19679 (N_19679,N_18715,N_18306);
xnor U19680 (N_19680,N_18328,N_18460);
or U19681 (N_19681,N_18098,N_18893);
nor U19682 (N_19682,N_18315,N_18439);
and U19683 (N_19683,N_18951,N_18386);
nor U19684 (N_19684,N_18112,N_18858);
and U19685 (N_19685,N_18710,N_18316);
and U19686 (N_19686,N_18762,N_18578);
or U19687 (N_19687,N_18558,N_18628);
nand U19688 (N_19688,N_18703,N_18132);
nor U19689 (N_19689,N_18781,N_18929);
xnor U19690 (N_19690,N_18569,N_18419);
and U19691 (N_19691,N_18243,N_18115);
nor U19692 (N_19692,N_18123,N_18262);
and U19693 (N_19693,N_18088,N_18886);
nor U19694 (N_19694,N_18968,N_18385);
and U19695 (N_19695,N_18900,N_18376);
xnor U19696 (N_19696,N_18830,N_18593);
xor U19697 (N_19697,N_18148,N_18335);
and U19698 (N_19698,N_18251,N_18834);
xor U19699 (N_19699,N_18432,N_18130);
nor U19700 (N_19700,N_18140,N_18458);
nor U19701 (N_19701,N_18532,N_18784);
nand U19702 (N_19702,N_18425,N_18185);
or U19703 (N_19703,N_18931,N_18102);
or U19704 (N_19704,N_18442,N_18290);
xnor U19705 (N_19705,N_18314,N_18634);
xnor U19706 (N_19706,N_18504,N_18557);
and U19707 (N_19707,N_18203,N_18831);
xnor U19708 (N_19708,N_18354,N_18886);
or U19709 (N_19709,N_18744,N_18035);
and U19710 (N_19710,N_18377,N_18117);
or U19711 (N_19711,N_18087,N_18222);
xor U19712 (N_19712,N_18851,N_18724);
xor U19713 (N_19713,N_18121,N_18507);
nor U19714 (N_19714,N_18881,N_18683);
or U19715 (N_19715,N_18451,N_18578);
and U19716 (N_19716,N_18994,N_18839);
or U19717 (N_19717,N_18092,N_18405);
nor U19718 (N_19718,N_18494,N_18388);
xor U19719 (N_19719,N_18044,N_18641);
nand U19720 (N_19720,N_18312,N_18204);
or U19721 (N_19721,N_18925,N_18179);
and U19722 (N_19722,N_18962,N_18744);
nand U19723 (N_19723,N_18256,N_18568);
nand U19724 (N_19724,N_18709,N_18773);
nor U19725 (N_19725,N_18938,N_18305);
xor U19726 (N_19726,N_18480,N_18709);
or U19727 (N_19727,N_18118,N_18832);
xnor U19728 (N_19728,N_18451,N_18959);
nand U19729 (N_19729,N_18212,N_18601);
or U19730 (N_19730,N_18538,N_18148);
xor U19731 (N_19731,N_18771,N_18649);
and U19732 (N_19732,N_18612,N_18263);
nand U19733 (N_19733,N_18252,N_18604);
or U19734 (N_19734,N_18776,N_18364);
nand U19735 (N_19735,N_18005,N_18823);
xnor U19736 (N_19736,N_18222,N_18762);
or U19737 (N_19737,N_18744,N_18271);
nand U19738 (N_19738,N_18065,N_18151);
nand U19739 (N_19739,N_18718,N_18466);
nand U19740 (N_19740,N_18567,N_18480);
or U19741 (N_19741,N_18985,N_18632);
or U19742 (N_19742,N_18925,N_18369);
and U19743 (N_19743,N_18928,N_18133);
and U19744 (N_19744,N_18552,N_18030);
or U19745 (N_19745,N_18762,N_18153);
nand U19746 (N_19746,N_18831,N_18240);
or U19747 (N_19747,N_18429,N_18386);
nor U19748 (N_19748,N_18656,N_18794);
nand U19749 (N_19749,N_18937,N_18356);
or U19750 (N_19750,N_18695,N_18884);
or U19751 (N_19751,N_18759,N_18504);
or U19752 (N_19752,N_18376,N_18595);
nor U19753 (N_19753,N_18873,N_18026);
nand U19754 (N_19754,N_18850,N_18055);
nor U19755 (N_19755,N_18296,N_18898);
nand U19756 (N_19756,N_18205,N_18108);
xor U19757 (N_19757,N_18467,N_18528);
and U19758 (N_19758,N_18662,N_18351);
nand U19759 (N_19759,N_18308,N_18625);
and U19760 (N_19760,N_18541,N_18927);
nand U19761 (N_19761,N_18837,N_18983);
and U19762 (N_19762,N_18161,N_18500);
nor U19763 (N_19763,N_18664,N_18247);
or U19764 (N_19764,N_18419,N_18071);
nor U19765 (N_19765,N_18264,N_18130);
nand U19766 (N_19766,N_18905,N_18601);
nand U19767 (N_19767,N_18581,N_18010);
and U19768 (N_19768,N_18019,N_18499);
nand U19769 (N_19769,N_18057,N_18859);
xnor U19770 (N_19770,N_18928,N_18787);
xnor U19771 (N_19771,N_18277,N_18303);
and U19772 (N_19772,N_18685,N_18030);
or U19773 (N_19773,N_18601,N_18718);
and U19774 (N_19774,N_18523,N_18136);
or U19775 (N_19775,N_18433,N_18520);
xnor U19776 (N_19776,N_18162,N_18692);
and U19777 (N_19777,N_18919,N_18319);
or U19778 (N_19778,N_18131,N_18498);
nor U19779 (N_19779,N_18919,N_18765);
nand U19780 (N_19780,N_18833,N_18853);
nand U19781 (N_19781,N_18493,N_18566);
nor U19782 (N_19782,N_18105,N_18505);
or U19783 (N_19783,N_18869,N_18768);
nor U19784 (N_19784,N_18611,N_18919);
or U19785 (N_19785,N_18863,N_18471);
xnor U19786 (N_19786,N_18016,N_18966);
or U19787 (N_19787,N_18021,N_18690);
nor U19788 (N_19788,N_18688,N_18371);
and U19789 (N_19789,N_18179,N_18016);
nand U19790 (N_19790,N_18308,N_18383);
xor U19791 (N_19791,N_18706,N_18331);
or U19792 (N_19792,N_18872,N_18134);
nand U19793 (N_19793,N_18782,N_18152);
or U19794 (N_19794,N_18790,N_18548);
xnor U19795 (N_19795,N_18747,N_18999);
nor U19796 (N_19796,N_18341,N_18000);
or U19797 (N_19797,N_18361,N_18043);
xor U19798 (N_19798,N_18896,N_18354);
nor U19799 (N_19799,N_18970,N_18718);
nand U19800 (N_19800,N_18055,N_18431);
nand U19801 (N_19801,N_18147,N_18036);
nor U19802 (N_19802,N_18760,N_18136);
nand U19803 (N_19803,N_18290,N_18920);
xor U19804 (N_19804,N_18748,N_18373);
and U19805 (N_19805,N_18234,N_18620);
nand U19806 (N_19806,N_18598,N_18007);
xnor U19807 (N_19807,N_18452,N_18615);
and U19808 (N_19808,N_18851,N_18220);
nor U19809 (N_19809,N_18170,N_18229);
and U19810 (N_19810,N_18787,N_18476);
or U19811 (N_19811,N_18717,N_18847);
nand U19812 (N_19812,N_18589,N_18694);
nand U19813 (N_19813,N_18814,N_18915);
xnor U19814 (N_19814,N_18739,N_18980);
nand U19815 (N_19815,N_18027,N_18902);
nor U19816 (N_19816,N_18556,N_18083);
nor U19817 (N_19817,N_18278,N_18520);
xor U19818 (N_19818,N_18757,N_18911);
and U19819 (N_19819,N_18023,N_18118);
xnor U19820 (N_19820,N_18214,N_18057);
nor U19821 (N_19821,N_18785,N_18751);
xnor U19822 (N_19822,N_18837,N_18886);
and U19823 (N_19823,N_18719,N_18256);
nand U19824 (N_19824,N_18917,N_18871);
xor U19825 (N_19825,N_18587,N_18690);
nand U19826 (N_19826,N_18245,N_18914);
and U19827 (N_19827,N_18736,N_18187);
nor U19828 (N_19828,N_18756,N_18806);
and U19829 (N_19829,N_18928,N_18456);
nand U19830 (N_19830,N_18774,N_18794);
xnor U19831 (N_19831,N_18743,N_18460);
nor U19832 (N_19832,N_18068,N_18948);
xnor U19833 (N_19833,N_18661,N_18491);
nor U19834 (N_19834,N_18932,N_18491);
nor U19835 (N_19835,N_18385,N_18041);
and U19836 (N_19836,N_18931,N_18732);
and U19837 (N_19837,N_18914,N_18674);
and U19838 (N_19838,N_18452,N_18029);
nor U19839 (N_19839,N_18362,N_18104);
xor U19840 (N_19840,N_18232,N_18259);
or U19841 (N_19841,N_18158,N_18104);
xor U19842 (N_19842,N_18945,N_18207);
or U19843 (N_19843,N_18849,N_18829);
nand U19844 (N_19844,N_18430,N_18057);
and U19845 (N_19845,N_18194,N_18703);
nand U19846 (N_19846,N_18254,N_18189);
nand U19847 (N_19847,N_18964,N_18869);
nand U19848 (N_19848,N_18224,N_18535);
or U19849 (N_19849,N_18449,N_18623);
nor U19850 (N_19850,N_18707,N_18292);
or U19851 (N_19851,N_18851,N_18820);
xnor U19852 (N_19852,N_18131,N_18985);
nor U19853 (N_19853,N_18541,N_18291);
xor U19854 (N_19854,N_18461,N_18436);
and U19855 (N_19855,N_18891,N_18433);
xor U19856 (N_19856,N_18489,N_18833);
nor U19857 (N_19857,N_18765,N_18317);
or U19858 (N_19858,N_18027,N_18261);
or U19859 (N_19859,N_18529,N_18848);
or U19860 (N_19860,N_18273,N_18838);
nand U19861 (N_19861,N_18868,N_18836);
and U19862 (N_19862,N_18396,N_18334);
and U19863 (N_19863,N_18488,N_18050);
nor U19864 (N_19864,N_18176,N_18928);
nor U19865 (N_19865,N_18387,N_18877);
nor U19866 (N_19866,N_18860,N_18696);
and U19867 (N_19867,N_18222,N_18404);
nand U19868 (N_19868,N_18096,N_18248);
nor U19869 (N_19869,N_18683,N_18488);
nor U19870 (N_19870,N_18328,N_18563);
nand U19871 (N_19871,N_18989,N_18822);
and U19872 (N_19872,N_18522,N_18758);
and U19873 (N_19873,N_18259,N_18631);
or U19874 (N_19874,N_18663,N_18935);
or U19875 (N_19875,N_18889,N_18716);
xor U19876 (N_19876,N_18927,N_18623);
nand U19877 (N_19877,N_18068,N_18259);
and U19878 (N_19878,N_18861,N_18842);
nand U19879 (N_19879,N_18629,N_18964);
nand U19880 (N_19880,N_18790,N_18200);
xnor U19881 (N_19881,N_18203,N_18817);
or U19882 (N_19882,N_18453,N_18070);
or U19883 (N_19883,N_18971,N_18653);
and U19884 (N_19884,N_18061,N_18174);
nand U19885 (N_19885,N_18432,N_18403);
nand U19886 (N_19886,N_18488,N_18070);
or U19887 (N_19887,N_18580,N_18602);
or U19888 (N_19888,N_18662,N_18963);
and U19889 (N_19889,N_18224,N_18267);
nor U19890 (N_19890,N_18963,N_18177);
xor U19891 (N_19891,N_18590,N_18528);
and U19892 (N_19892,N_18655,N_18697);
nor U19893 (N_19893,N_18934,N_18357);
xor U19894 (N_19894,N_18989,N_18882);
or U19895 (N_19895,N_18769,N_18667);
or U19896 (N_19896,N_18920,N_18481);
nand U19897 (N_19897,N_18036,N_18171);
nor U19898 (N_19898,N_18595,N_18430);
or U19899 (N_19899,N_18652,N_18634);
nor U19900 (N_19900,N_18356,N_18538);
nor U19901 (N_19901,N_18375,N_18441);
and U19902 (N_19902,N_18095,N_18355);
and U19903 (N_19903,N_18839,N_18569);
nor U19904 (N_19904,N_18399,N_18696);
or U19905 (N_19905,N_18102,N_18505);
xnor U19906 (N_19906,N_18457,N_18528);
nor U19907 (N_19907,N_18985,N_18103);
nand U19908 (N_19908,N_18107,N_18775);
and U19909 (N_19909,N_18823,N_18275);
nand U19910 (N_19910,N_18022,N_18423);
or U19911 (N_19911,N_18889,N_18520);
nand U19912 (N_19912,N_18513,N_18753);
nand U19913 (N_19913,N_18300,N_18036);
and U19914 (N_19914,N_18099,N_18984);
and U19915 (N_19915,N_18723,N_18419);
nand U19916 (N_19916,N_18210,N_18132);
or U19917 (N_19917,N_18822,N_18357);
nand U19918 (N_19918,N_18073,N_18367);
nand U19919 (N_19919,N_18172,N_18892);
or U19920 (N_19920,N_18778,N_18953);
and U19921 (N_19921,N_18962,N_18619);
and U19922 (N_19922,N_18147,N_18173);
xnor U19923 (N_19923,N_18302,N_18624);
xor U19924 (N_19924,N_18125,N_18299);
and U19925 (N_19925,N_18958,N_18557);
xor U19926 (N_19926,N_18341,N_18464);
or U19927 (N_19927,N_18534,N_18410);
nor U19928 (N_19928,N_18228,N_18450);
nor U19929 (N_19929,N_18605,N_18234);
or U19930 (N_19930,N_18446,N_18267);
or U19931 (N_19931,N_18845,N_18562);
nand U19932 (N_19932,N_18634,N_18865);
nor U19933 (N_19933,N_18829,N_18071);
xor U19934 (N_19934,N_18822,N_18671);
nand U19935 (N_19935,N_18923,N_18558);
nor U19936 (N_19936,N_18223,N_18355);
and U19937 (N_19937,N_18795,N_18135);
and U19938 (N_19938,N_18902,N_18712);
nor U19939 (N_19939,N_18174,N_18603);
xnor U19940 (N_19940,N_18421,N_18105);
xor U19941 (N_19941,N_18020,N_18388);
nand U19942 (N_19942,N_18759,N_18465);
or U19943 (N_19943,N_18890,N_18057);
or U19944 (N_19944,N_18510,N_18293);
nor U19945 (N_19945,N_18975,N_18381);
nor U19946 (N_19946,N_18992,N_18231);
or U19947 (N_19947,N_18816,N_18465);
nand U19948 (N_19948,N_18722,N_18936);
nand U19949 (N_19949,N_18275,N_18609);
nor U19950 (N_19950,N_18032,N_18814);
and U19951 (N_19951,N_18157,N_18685);
or U19952 (N_19952,N_18807,N_18888);
nor U19953 (N_19953,N_18926,N_18049);
xor U19954 (N_19954,N_18455,N_18661);
xnor U19955 (N_19955,N_18062,N_18994);
and U19956 (N_19956,N_18596,N_18570);
xnor U19957 (N_19957,N_18686,N_18621);
nand U19958 (N_19958,N_18361,N_18286);
nand U19959 (N_19959,N_18158,N_18738);
nor U19960 (N_19960,N_18919,N_18968);
and U19961 (N_19961,N_18190,N_18792);
xor U19962 (N_19962,N_18272,N_18611);
xnor U19963 (N_19963,N_18034,N_18853);
and U19964 (N_19964,N_18821,N_18542);
nor U19965 (N_19965,N_18527,N_18227);
nor U19966 (N_19966,N_18623,N_18974);
or U19967 (N_19967,N_18682,N_18428);
or U19968 (N_19968,N_18841,N_18539);
xor U19969 (N_19969,N_18055,N_18775);
nor U19970 (N_19970,N_18179,N_18985);
nand U19971 (N_19971,N_18749,N_18569);
nor U19972 (N_19972,N_18812,N_18288);
and U19973 (N_19973,N_18922,N_18138);
and U19974 (N_19974,N_18460,N_18812);
nand U19975 (N_19975,N_18497,N_18567);
and U19976 (N_19976,N_18567,N_18280);
nand U19977 (N_19977,N_18847,N_18747);
nor U19978 (N_19978,N_18564,N_18206);
nand U19979 (N_19979,N_18057,N_18748);
nor U19980 (N_19980,N_18648,N_18698);
xnor U19981 (N_19981,N_18871,N_18313);
nor U19982 (N_19982,N_18729,N_18357);
nor U19983 (N_19983,N_18428,N_18980);
xnor U19984 (N_19984,N_18009,N_18072);
and U19985 (N_19985,N_18055,N_18331);
and U19986 (N_19986,N_18184,N_18804);
and U19987 (N_19987,N_18140,N_18398);
xor U19988 (N_19988,N_18445,N_18578);
nand U19989 (N_19989,N_18374,N_18460);
xnor U19990 (N_19990,N_18141,N_18194);
xnor U19991 (N_19991,N_18452,N_18732);
or U19992 (N_19992,N_18222,N_18500);
nor U19993 (N_19993,N_18646,N_18280);
and U19994 (N_19994,N_18353,N_18130);
or U19995 (N_19995,N_18698,N_18155);
xnor U19996 (N_19996,N_18086,N_18771);
nor U19997 (N_19997,N_18622,N_18415);
nand U19998 (N_19998,N_18436,N_18453);
nand U19999 (N_19999,N_18181,N_18537);
nand U20000 (N_20000,N_19018,N_19476);
nand U20001 (N_20001,N_19742,N_19947);
and U20002 (N_20002,N_19532,N_19284);
xor U20003 (N_20003,N_19114,N_19340);
nor U20004 (N_20004,N_19332,N_19734);
and U20005 (N_20005,N_19876,N_19237);
nor U20006 (N_20006,N_19050,N_19273);
nand U20007 (N_20007,N_19611,N_19472);
nor U20008 (N_20008,N_19017,N_19227);
xor U20009 (N_20009,N_19987,N_19820);
or U20010 (N_20010,N_19622,N_19246);
and U20011 (N_20011,N_19475,N_19562);
nor U20012 (N_20012,N_19564,N_19295);
nand U20013 (N_20013,N_19244,N_19449);
and U20014 (N_20014,N_19037,N_19026);
and U20015 (N_20015,N_19899,N_19552);
or U20016 (N_20016,N_19910,N_19197);
and U20017 (N_20017,N_19623,N_19720);
nor U20018 (N_20018,N_19436,N_19047);
xor U20019 (N_20019,N_19470,N_19399);
nor U20020 (N_20020,N_19956,N_19378);
xnor U20021 (N_20021,N_19211,N_19132);
xnor U20022 (N_20022,N_19610,N_19941);
nor U20023 (N_20023,N_19333,N_19639);
nand U20024 (N_20024,N_19774,N_19542);
nor U20025 (N_20025,N_19831,N_19558);
nand U20026 (N_20026,N_19784,N_19369);
and U20027 (N_20027,N_19609,N_19903);
and U20028 (N_20028,N_19940,N_19543);
nand U20029 (N_20029,N_19514,N_19446);
xor U20030 (N_20030,N_19042,N_19595);
or U20031 (N_20031,N_19326,N_19215);
xnor U20032 (N_20032,N_19366,N_19465);
nor U20033 (N_20033,N_19041,N_19346);
xor U20034 (N_20034,N_19756,N_19459);
nand U20035 (N_20035,N_19683,N_19559);
or U20036 (N_20036,N_19663,N_19766);
or U20037 (N_20037,N_19155,N_19557);
or U20038 (N_20038,N_19833,N_19196);
or U20039 (N_20039,N_19396,N_19515);
nor U20040 (N_20040,N_19953,N_19823);
xnor U20041 (N_20041,N_19177,N_19904);
nor U20042 (N_20042,N_19240,N_19834);
nor U20043 (N_20043,N_19590,N_19394);
and U20044 (N_20044,N_19123,N_19529);
xor U20045 (N_20045,N_19567,N_19137);
or U20046 (N_20046,N_19250,N_19403);
nand U20047 (N_20047,N_19839,N_19430);
nand U20048 (N_20048,N_19835,N_19624);
xor U20049 (N_20049,N_19738,N_19750);
nand U20050 (N_20050,N_19686,N_19889);
nor U20051 (N_20051,N_19646,N_19619);
xnor U20052 (N_20052,N_19317,N_19805);
or U20053 (N_20053,N_19108,N_19966);
nand U20054 (N_20054,N_19670,N_19799);
nand U20055 (N_20055,N_19874,N_19431);
xnor U20056 (N_20056,N_19395,N_19585);
nand U20057 (N_20057,N_19019,N_19676);
xnor U20058 (N_20058,N_19583,N_19969);
or U20059 (N_20059,N_19822,N_19357);
and U20060 (N_20060,N_19363,N_19763);
and U20061 (N_20061,N_19687,N_19827);
or U20062 (N_20062,N_19570,N_19199);
and U20063 (N_20063,N_19933,N_19679);
nand U20064 (N_20064,N_19934,N_19817);
xnor U20065 (N_20065,N_19844,N_19882);
or U20066 (N_20066,N_19927,N_19209);
nand U20067 (N_20067,N_19741,N_19471);
or U20068 (N_20068,N_19483,N_19792);
nand U20069 (N_20069,N_19528,N_19451);
nor U20070 (N_20070,N_19918,N_19325);
nand U20071 (N_20071,N_19468,N_19860);
nor U20072 (N_20072,N_19389,N_19535);
and U20073 (N_20073,N_19189,N_19490);
xor U20074 (N_20074,N_19186,N_19656);
nor U20075 (N_20075,N_19764,N_19975);
and U20076 (N_20076,N_19594,N_19090);
xnor U20077 (N_20077,N_19531,N_19522);
or U20078 (N_20078,N_19992,N_19185);
xor U20079 (N_20079,N_19702,N_19599);
or U20080 (N_20080,N_19616,N_19011);
nand U20081 (N_20081,N_19296,N_19384);
nor U20082 (N_20082,N_19020,N_19418);
xor U20083 (N_20083,N_19963,N_19689);
or U20084 (N_20084,N_19809,N_19501);
nor U20085 (N_20085,N_19849,N_19103);
xor U20086 (N_20086,N_19724,N_19003);
and U20087 (N_20087,N_19086,N_19651);
nor U20088 (N_20088,N_19694,N_19761);
and U20089 (N_20089,N_19748,N_19524);
nand U20090 (N_20090,N_19314,N_19193);
or U20091 (N_20091,N_19053,N_19510);
nor U20092 (N_20092,N_19950,N_19888);
xor U20093 (N_20093,N_19278,N_19156);
and U20094 (N_20094,N_19589,N_19055);
or U20095 (N_20095,N_19322,N_19051);
and U20096 (N_20096,N_19582,N_19007);
or U20097 (N_20097,N_19659,N_19856);
or U20098 (N_20098,N_19723,N_19015);
nand U20099 (N_20099,N_19715,N_19069);
and U20100 (N_20100,N_19083,N_19424);
or U20101 (N_20101,N_19421,N_19790);
xor U20102 (N_20102,N_19016,N_19235);
xnor U20103 (N_20103,N_19440,N_19548);
xnor U20104 (N_20104,N_19283,N_19508);
xor U20105 (N_20105,N_19085,N_19710);
nor U20106 (N_20106,N_19310,N_19920);
nor U20107 (N_20107,N_19124,N_19749);
nand U20108 (N_20108,N_19349,N_19913);
xnor U20109 (N_20109,N_19816,N_19150);
xor U20110 (N_20110,N_19388,N_19350);
xnor U20111 (N_20111,N_19785,N_19168);
or U20112 (N_20112,N_19243,N_19365);
xor U20113 (N_20113,N_19668,N_19182);
nand U20114 (N_20114,N_19719,N_19348);
and U20115 (N_20115,N_19484,N_19635);
and U20116 (N_20116,N_19536,N_19793);
nand U20117 (N_20117,N_19461,N_19167);
nand U20118 (N_20118,N_19187,N_19245);
and U20119 (N_20119,N_19022,N_19667);
and U20120 (N_20120,N_19525,N_19276);
or U20121 (N_20121,N_19226,N_19126);
xnor U20122 (N_20122,N_19337,N_19690);
or U20123 (N_20123,N_19464,N_19566);
and U20124 (N_20124,N_19824,N_19607);
nand U20125 (N_20125,N_19873,N_19173);
or U20126 (N_20126,N_19640,N_19408);
xnor U20127 (N_20127,N_19454,N_19338);
and U20128 (N_20128,N_19819,N_19780);
nand U20129 (N_20129,N_19485,N_19821);
or U20130 (N_20130,N_19642,N_19212);
nand U20131 (N_20131,N_19135,N_19077);
xnor U20132 (N_20132,N_19239,N_19968);
or U20133 (N_20133,N_19142,N_19358);
nand U20134 (N_20134,N_19703,N_19068);
xor U20135 (N_20135,N_19154,N_19166);
nor U20136 (N_20136,N_19178,N_19000);
or U20137 (N_20137,N_19079,N_19251);
and U20138 (N_20138,N_19084,N_19813);
xnor U20139 (N_20139,N_19519,N_19708);
nand U20140 (N_20140,N_19818,N_19134);
nor U20141 (N_20141,N_19443,N_19989);
xor U20142 (N_20142,N_19262,N_19621);
nand U20143 (N_20143,N_19955,N_19588);
or U20144 (N_20144,N_19788,N_19576);
nor U20145 (N_20145,N_19843,N_19417);
xor U20146 (N_20146,N_19188,N_19803);
nor U20147 (N_20147,N_19480,N_19422);
and U20148 (N_20148,N_19939,N_19184);
and U20149 (N_20149,N_19046,N_19441);
or U20150 (N_20150,N_19974,N_19321);
xnor U20151 (N_20151,N_19192,N_19098);
xor U20152 (N_20152,N_19125,N_19405);
nand U20153 (N_20153,N_19347,N_19481);
and U20154 (N_20154,N_19049,N_19315);
or U20155 (N_20155,N_19128,N_19665);
or U20156 (N_20156,N_19620,N_19078);
and U20157 (N_20157,N_19540,N_19554);
and U20158 (N_20158,N_19630,N_19592);
nor U20159 (N_20159,N_19469,N_19213);
nand U20160 (N_20160,N_19311,N_19252);
nand U20161 (N_20161,N_19980,N_19129);
and U20162 (N_20162,N_19368,N_19765);
nor U20163 (N_20163,N_19677,N_19351);
xnor U20164 (N_20164,N_19911,N_19027);
and U20165 (N_20165,N_19247,N_19059);
nand U20166 (N_20166,N_19058,N_19754);
nor U20167 (N_20167,N_19716,N_19662);
xnor U20168 (N_20168,N_19398,N_19930);
nand U20169 (N_20169,N_19204,N_19136);
nand U20170 (N_20170,N_19367,N_19444);
or U20171 (N_20171,N_19201,N_19162);
and U20172 (N_20172,N_19241,N_19807);
or U20173 (N_20173,N_19830,N_19488);
nand U20174 (N_20174,N_19804,N_19385);
or U20175 (N_20175,N_19778,N_19313);
and U20176 (N_20176,N_19248,N_19320);
and U20177 (N_20177,N_19163,N_19513);
xor U20178 (N_20178,N_19442,N_19221);
nand U20179 (N_20179,N_19413,N_19717);
and U20180 (N_20180,N_19060,N_19419);
xor U20181 (N_20181,N_19695,N_19954);
xor U20182 (N_20182,N_19293,N_19923);
or U20183 (N_20183,N_19133,N_19905);
nand U20184 (N_20184,N_19074,N_19033);
xor U20185 (N_20185,N_19721,N_19447);
xnor U20186 (N_20186,N_19467,N_19257);
and U20187 (N_20187,N_19301,N_19837);
nand U20188 (N_20188,N_19373,N_19025);
or U20189 (N_20189,N_19897,N_19757);
nand U20190 (N_20190,N_19509,N_19104);
or U20191 (N_20191,N_19100,N_19001);
nand U20192 (N_20192,N_19743,N_19238);
nor U20193 (N_20193,N_19127,N_19190);
or U20194 (N_20194,N_19815,N_19453);
or U20195 (N_20195,N_19770,N_19195);
nor U20196 (N_20196,N_19907,N_19885);
or U20197 (N_20197,N_19316,N_19675);
nand U20198 (N_20198,N_19099,N_19021);
xor U20199 (N_20199,N_19236,N_19220);
nand U20200 (N_20200,N_19896,N_19744);
nor U20201 (N_20201,N_19795,N_19879);
or U20202 (N_20202,N_19404,N_19674);
and U20203 (N_20203,N_19655,N_19569);
or U20204 (N_20204,N_19353,N_19426);
nand U20205 (N_20205,N_19502,N_19961);
nand U20206 (N_20206,N_19280,N_19706);
nand U20207 (N_20207,N_19063,N_19288);
or U20208 (N_20208,N_19629,N_19714);
nand U20209 (N_20209,N_19306,N_19959);
and U20210 (N_20210,N_19832,N_19729);
and U20211 (N_20211,N_19080,N_19153);
or U20212 (N_20212,N_19908,N_19962);
and U20213 (N_20213,N_19632,N_19254);
xnor U20214 (N_20214,N_19160,N_19932);
nand U20215 (N_20215,N_19685,N_19682);
nand U20216 (N_20216,N_19596,N_19300);
nor U20217 (N_20217,N_19777,N_19265);
and U20218 (N_20218,N_19797,N_19507);
nor U20219 (N_20219,N_19354,N_19909);
xor U20220 (N_20220,N_19650,N_19870);
nor U20221 (N_20221,N_19157,N_19994);
xor U20222 (N_20222,N_19216,N_19092);
or U20223 (N_20223,N_19376,N_19194);
xor U20224 (N_20224,N_19070,N_19038);
xnor U20225 (N_20225,N_19291,N_19214);
xor U20226 (N_20226,N_19277,N_19842);
or U20227 (N_20227,N_19584,N_19746);
xor U20228 (N_20228,N_19854,N_19298);
or U20229 (N_20229,N_19409,N_19556);
nand U20230 (N_20230,N_19180,N_19638);
or U20231 (N_20231,N_19740,N_19942);
nor U20232 (N_20232,N_19004,N_19372);
nand U20233 (N_20233,N_19474,N_19304);
xor U20234 (N_20234,N_19169,N_19960);
and U20235 (N_20235,N_19944,N_19993);
xnor U20236 (N_20236,N_19445,N_19981);
or U20237 (N_20237,N_19534,N_19122);
and U20238 (N_20238,N_19645,N_19782);
xor U20239 (N_20239,N_19081,N_19499);
and U20240 (N_20240,N_19794,N_19530);
nand U20241 (N_20241,N_19005,N_19343);
or U20242 (N_20242,N_19627,N_19275);
nand U20243 (N_20243,N_19572,N_19512);
nor U20244 (N_20244,N_19506,N_19867);
or U20245 (N_20245,N_19952,N_19497);
xor U20246 (N_20246,N_19853,N_19149);
and U20247 (N_20247,N_19318,N_19684);
nor U20248 (N_20248,N_19951,N_19840);
nand U20249 (N_20249,N_19931,N_19551);
nand U20250 (N_20250,N_19730,N_19270);
nand U20251 (N_20251,N_19170,N_19680);
nor U20252 (N_20252,N_19460,N_19852);
and U20253 (N_20253,N_19605,N_19926);
nor U20254 (N_20254,N_19767,N_19877);
nor U20255 (N_20255,N_19202,N_19052);
nor U20256 (N_20256,N_19733,N_19511);
nand U20257 (N_20257,N_19228,N_19139);
nand U20258 (N_20258,N_19979,N_19117);
or U20259 (N_20259,N_19625,N_19075);
or U20260 (N_20260,N_19056,N_19073);
or U20261 (N_20261,N_19224,N_19158);
nand U20262 (N_20262,N_19586,N_19455);
nand U20263 (N_20263,N_19571,N_19102);
nor U20264 (N_20264,N_19242,N_19577);
and U20265 (N_20265,N_19323,N_19341);
nor U20266 (N_20266,N_19486,N_19152);
nand U20267 (N_20267,N_19089,N_19798);
nand U20268 (N_20268,N_19014,N_19118);
nor U20269 (N_20269,N_19891,N_19678);
and U20270 (N_20270,N_19545,N_19845);
or U20271 (N_20271,N_19407,N_19527);
or U20272 (N_20272,N_19279,N_19549);
nor U20273 (N_20273,N_19705,N_19713);
xor U20274 (N_20274,N_19660,N_19072);
xor U20275 (N_20275,N_19290,N_19045);
or U20276 (N_20276,N_19009,N_19985);
nand U20277 (N_20277,N_19802,N_19673);
and U20278 (N_20278,N_19339,N_19364);
and U20279 (N_20279,N_19786,N_19324);
or U20280 (N_20280,N_19429,N_19151);
and U20281 (N_20281,N_19500,N_19159);
xor U20282 (N_20282,N_19161,N_19334);
nand U20283 (N_20283,N_19995,N_19412);
nor U20284 (N_20284,N_19144,N_19495);
xnor U20285 (N_20285,N_19023,N_19165);
xor U20286 (N_20286,N_19671,N_19119);
and U20287 (N_20287,N_19064,N_19915);
xor U20288 (N_20288,N_19810,N_19071);
or U20289 (N_20289,N_19600,N_19681);
or U20290 (N_20290,N_19967,N_19760);
nand U20291 (N_20291,N_19416,N_19574);
or U20292 (N_20292,N_19303,N_19390);
xnor U20293 (N_20293,N_19336,N_19294);
or U20294 (N_20294,N_19111,N_19539);
nor U20295 (N_20295,N_19652,N_19614);
xnor U20296 (N_20296,N_19223,N_19482);
and U20297 (N_20297,N_19986,N_19550);
and U20298 (N_20298,N_19400,N_19203);
and U20299 (N_20299,N_19983,N_19762);
xnor U20300 (N_20300,N_19565,N_19957);
nor U20301 (N_20301,N_19858,N_19411);
nor U20302 (N_20302,N_19919,N_19308);
and U20303 (N_20303,N_19973,N_19737);
or U20304 (N_20304,N_19697,N_19886);
and U20305 (N_20305,N_19759,N_19379);
nor U20306 (N_20306,N_19800,N_19601);
and U20307 (N_20307,N_19851,N_19386);
and U20308 (N_20308,N_19634,N_19829);
xor U20309 (N_20309,N_19861,N_19002);
nor U20310 (N_20310,N_19207,N_19253);
nor U20311 (N_20311,N_19965,N_19887);
nand U20312 (N_20312,N_19289,N_19863);
nor U20313 (N_20313,N_19937,N_19666);
nand U20314 (N_20314,N_19012,N_19146);
xor U20315 (N_20315,N_19044,N_19330);
xnor U20316 (N_20316,N_19437,N_19608);
or U20317 (N_20317,N_19106,N_19894);
and U20318 (N_20318,N_19722,N_19631);
nand U20319 (N_20319,N_19029,N_19493);
nand U20320 (N_20320,N_19617,N_19260);
or U20321 (N_20321,N_19949,N_19101);
nand U20322 (N_20322,N_19272,N_19925);
nand U20323 (N_20323,N_19375,N_19219);
or U20324 (N_20324,N_19520,N_19263);
nand U20325 (N_20325,N_19884,N_19718);
xnor U20326 (N_20326,N_19107,N_19751);
nor U20327 (N_20327,N_19848,N_19649);
or U20328 (N_20328,N_19898,N_19043);
xor U20329 (N_20329,N_19233,N_19274);
and U20330 (N_20330,N_19113,N_19523);
nand U20331 (N_20331,N_19477,N_19095);
and U20332 (N_20332,N_19948,N_19864);
or U20333 (N_20333,N_19647,N_19626);
or U20334 (N_20334,N_19563,N_19024);
nand U20335 (N_20335,N_19922,N_19603);
and U20336 (N_20336,N_19381,N_19964);
and U20337 (N_20337,N_19172,N_19587);
xor U20338 (N_20338,N_19836,N_19342);
nand U20339 (N_20339,N_19521,N_19067);
and U20340 (N_20340,N_19654,N_19657);
nor U20341 (N_20341,N_19115,N_19555);
nor U20342 (N_20342,N_19148,N_19838);
and U20343 (N_20343,N_19517,N_19597);
and U20344 (N_20344,N_19061,N_19880);
and U20345 (N_20345,N_19008,N_19120);
and U20346 (N_20346,N_19560,N_19496);
and U20347 (N_20347,N_19281,N_19054);
nor U20348 (N_20348,N_19039,N_19175);
or U20349 (N_20349,N_19847,N_19808);
nand U20350 (N_20350,N_19494,N_19999);
and U20351 (N_20351,N_19425,N_19344);
and U20352 (N_20352,N_19711,N_19269);
or U20353 (N_20353,N_19602,N_19487);
nor U20354 (N_20354,N_19504,N_19264);
nand U20355 (N_20355,N_19789,N_19091);
and U20356 (N_20356,N_19814,N_19773);
nor U20357 (N_20357,N_19065,N_19735);
or U20358 (N_20358,N_19147,N_19928);
xor U20359 (N_20359,N_19096,N_19463);
or U20360 (N_20360,N_19618,N_19781);
nor U20361 (N_20361,N_19648,N_19094);
nand U20362 (N_20362,N_19997,N_19544);
xor U20363 (N_20363,N_19812,N_19062);
and U20364 (N_20364,N_19006,N_19892);
nor U20365 (N_20365,N_19093,N_19359);
nand U20366 (N_20366,N_19971,N_19935);
and U20367 (N_20367,N_19698,N_19653);
or U20368 (N_20368,N_19361,N_19450);
or U20369 (N_20369,N_19034,N_19796);
or U20370 (N_20370,N_19143,N_19533);
nand U20371 (N_20371,N_19747,N_19598);
and U20372 (N_20372,N_19181,N_19636);
and U20373 (N_20373,N_19806,N_19538);
or U20374 (N_20374,N_19725,N_19200);
and U20375 (N_20375,N_19218,N_19701);
and U20376 (N_20376,N_19772,N_19669);
and U20377 (N_20377,N_19414,N_19140);
or U20378 (N_20378,N_19391,N_19319);
xor U20379 (N_20379,N_19259,N_19526);
nand U20380 (N_20380,N_19036,N_19580);
nand U20381 (N_20381,N_19109,N_19518);
or U20382 (N_20382,N_19739,N_19374);
xnor U20383 (N_20383,N_19901,N_19914);
xor U20384 (N_20384,N_19991,N_19727);
nand U20385 (N_20385,N_19745,N_19872);
nand U20386 (N_20386,N_19230,N_19553);
and U20387 (N_20387,N_19097,N_19292);
xnor U20388 (N_20388,N_19057,N_19664);
or U20389 (N_20389,N_19356,N_19312);
nand U20390 (N_20390,N_19256,N_19775);
and U20391 (N_20391,N_19401,N_19633);
and U20392 (N_20392,N_19862,N_19452);
nand U20393 (N_20393,N_19672,N_19906);
or U20394 (N_20394,N_19268,N_19732);
or U20395 (N_20395,N_19434,N_19176);
nor U20396 (N_20396,N_19731,N_19392);
nand U20397 (N_20397,N_19779,N_19699);
nand U20398 (N_20398,N_19846,N_19998);
xor U20399 (N_20399,N_19433,N_19088);
nand U20400 (N_20400,N_19435,N_19641);
xor U20401 (N_20401,N_19866,N_19547);
and U20402 (N_20402,N_19771,N_19383);
xor U20403 (N_20403,N_19371,N_19145);
nand U20404 (N_20404,N_19415,N_19438);
xnor U20405 (N_20405,N_19758,N_19871);
or U20406 (N_20406,N_19406,N_19769);
and U20407 (N_20407,N_19828,N_19752);
and U20408 (N_20408,N_19225,N_19217);
or U20409 (N_20409,N_19945,N_19783);
xnor U20410 (N_20410,N_19335,N_19164);
and U20411 (N_20411,N_19691,N_19801);
or U20412 (N_20412,N_19516,N_19458);
xor U20413 (N_20413,N_19473,N_19255);
and U20414 (N_20414,N_19958,N_19287);
xnor U20415 (N_20415,N_19984,N_19138);
nor U20416 (N_20416,N_19561,N_19787);
xor U20417 (N_20417,N_19893,N_19229);
and U20418 (N_20418,N_19491,N_19028);
nand U20419 (N_20419,N_19420,N_19210);
xor U20420 (N_20420,N_19568,N_19615);
and U20421 (N_20421,N_19205,N_19988);
or U20422 (N_20422,N_19883,N_19970);
or U20423 (N_20423,N_19261,N_19208);
and U20424 (N_20424,N_19895,N_19282);
nand U20425 (N_20425,N_19696,N_19466);
nand U20426 (N_20426,N_19581,N_19031);
or U20427 (N_20427,N_19393,N_19360);
and U20428 (N_20428,N_19105,N_19032);
nand U20429 (N_20429,N_19087,N_19286);
nor U20430 (N_20430,N_19841,N_19936);
nand U20431 (N_20431,N_19130,N_19643);
or U20432 (N_20432,N_19776,N_19258);
nand U20433 (N_20433,N_19387,N_19753);
and U20434 (N_20434,N_19370,N_19355);
nor U20435 (N_20435,N_19040,N_19693);
nand U20436 (N_20436,N_19110,N_19878);
nor U20437 (N_20437,N_19362,N_19612);
and U20438 (N_20438,N_19305,N_19943);
nor U20439 (N_20439,N_19076,N_19112);
xor U20440 (N_20440,N_19726,N_19875);
nor U20441 (N_20441,N_19902,N_19505);
nand U20442 (N_20442,N_19977,N_19035);
nand U20443 (N_20443,N_19912,N_19066);
or U20444 (N_20444,N_19121,N_19428);
nand U20445 (N_20445,N_19857,N_19191);
xor U20446 (N_20446,N_19791,N_19397);
xnor U20447 (N_20447,N_19946,N_19116);
xnor U20448 (N_20448,N_19990,N_19859);
and U20449 (N_20449,N_19704,N_19498);
and U20450 (N_20450,N_19141,N_19171);
or U20451 (N_20451,N_19266,N_19658);
xnor U20452 (N_20452,N_19768,N_19329);
and U20453 (N_20453,N_19503,N_19345);
and U20454 (N_20454,N_19996,N_19377);
or U20455 (N_20455,N_19712,N_19688);
nor U20456 (N_20456,N_19613,N_19606);
nor U20457 (N_20457,N_19082,N_19234);
or U20458 (N_20458,N_19546,N_19881);
nor U20459 (N_20459,N_19728,N_19232);
and U20460 (N_20460,N_19736,N_19231);
and U20461 (N_20461,N_19978,N_19307);
or U20462 (N_20462,N_19579,N_19709);
and U20463 (N_20463,N_19380,N_19328);
nor U20464 (N_20464,N_19825,N_19198);
nor U20465 (N_20465,N_19013,N_19222);
or U20466 (N_20466,N_19976,N_19479);
or U20467 (N_20467,N_19299,N_19929);
xnor U20468 (N_20468,N_19423,N_19637);
or U20469 (N_20469,N_19179,N_19448);
nor U20470 (N_20470,N_19972,N_19309);
nor U20471 (N_20471,N_19593,N_19302);
and U20472 (N_20472,N_19541,N_19537);
nor U20473 (N_20473,N_19700,N_19489);
or U20474 (N_20474,N_19327,N_19573);
xor U20475 (N_20475,N_19462,N_19048);
or U20476 (N_20476,N_19644,N_19850);
nor U20477 (N_20477,N_19826,N_19492);
xnor U20478 (N_20478,N_19604,N_19938);
xor U20479 (N_20479,N_19578,N_19575);
nand U20480 (N_20480,N_19811,N_19628);
nor U20481 (N_20481,N_19900,N_19457);
and U20482 (N_20482,N_19855,N_19410);
nand U20483 (N_20483,N_19271,N_19030);
nand U20484 (N_20484,N_19868,N_19206);
xnor U20485 (N_20485,N_19924,N_19249);
nor U20486 (N_20486,N_19010,N_19456);
nand U20487 (N_20487,N_19707,N_19755);
and U20488 (N_20488,N_19331,N_19890);
nand U20489 (N_20489,N_19916,N_19174);
nor U20490 (N_20490,N_19865,N_19297);
xor U20491 (N_20491,N_19478,N_19591);
or U20492 (N_20492,N_19917,N_19131);
or U20493 (N_20493,N_19285,N_19427);
nand U20494 (N_20494,N_19183,N_19921);
or U20495 (N_20495,N_19267,N_19382);
or U20496 (N_20496,N_19661,N_19402);
xor U20497 (N_20497,N_19869,N_19432);
xnor U20498 (N_20498,N_19982,N_19352);
or U20499 (N_20499,N_19439,N_19692);
and U20500 (N_20500,N_19690,N_19123);
xor U20501 (N_20501,N_19348,N_19566);
nand U20502 (N_20502,N_19387,N_19417);
nand U20503 (N_20503,N_19771,N_19991);
and U20504 (N_20504,N_19671,N_19036);
and U20505 (N_20505,N_19521,N_19864);
xnor U20506 (N_20506,N_19853,N_19244);
or U20507 (N_20507,N_19671,N_19605);
or U20508 (N_20508,N_19936,N_19881);
or U20509 (N_20509,N_19480,N_19541);
nor U20510 (N_20510,N_19598,N_19878);
and U20511 (N_20511,N_19464,N_19991);
and U20512 (N_20512,N_19180,N_19562);
xnor U20513 (N_20513,N_19680,N_19318);
nand U20514 (N_20514,N_19894,N_19347);
and U20515 (N_20515,N_19038,N_19084);
and U20516 (N_20516,N_19569,N_19669);
or U20517 (N_20517,N_19901,N_19075);
or U20518 (N_20518,N_19062,N_19805);
and U20519 (N_20519,N_19569,N_19399);
or U20520 (N_20520,N_19406,N_19602);
nor U20521 (N_20521,N_19722,N_19344);
and U20522 (N_20522,N_19775,N_19530);
nor U20523 (N_20523,N_19113,N_19075);
xor U20524 (N_20524,N_19534,N_19052);
and U20525 (N_20525,N_19906,N_19075);
and U20526 (N_20526,N_19642,N_19247);
and U20527 (N_20527,N_19345,N_19296);
or U20528 (N_20528,N_19880,N_19433);
nand U20529 (N_20529,N_19550,N_19125);
xor U20530 (N_20530,N_19932,N_19487);
xnor U20531 (N_20531,N_19556,N_19381);
and U20532 (N_20532,N_19039,N_19404);
nor U20533 (N_20533,N_19404,N_19233);
nand U20534 (N_20534,N_19923,N_19297);
nand U20535 (N_20535,N_19358,N_19060);
xnor U20536 (N_20536,N_19242,N_19422);
nor U20537 (N_20537,N_19180,N_19048);
and U20538 (N_20538,N_19809,N_19775);
nand U20539 (N_20539,N_19938,N_19103);
xnor U20540 (N_20540,N_19201,N_19602);
nand U20541 (N_20541,N_19142,N_19868);
and U20542 (N_20542,N_19116,N_19885);
and U20543 (N_20543,N_19605,N_19929);
or U20544 (N_20544,N_19537,N_19793);
or U20545 (N_20545,N_19354,N_19763);
or U20546 (N_20546,N_19945,N_19509);
xnor U20547 (N_20547,N_19722,N_19112);
and U20548 (N_20548,N_19599,N_19283);
or U20549 (N_20549,N_19450,N_19580);
or U20550 (N_20550,N_19287,N_19435);
xnor U20551 (N_20551,N_19632,N_19269);
nand U20552 (N_20552,N_19386,N_19115);
or U20553 (N_20553,N_19193,N_19749);
nand U20554 (N_20554,N_19400,N_19063);
xor U20555 (N_20555,N_19171,N_19689);
nor U20556 (N_20556,N_19930,N_19705);
or U20557 (N_20557,N_19212,N_19737);
and U20558 (N_20558,N_19708,N_19776);
or U20559 (N_20559,N_19173,N_19608);
or U20560 (N_20560,N_19652,N_19022);
nand U20561 (N_20561,N_19679,N_19179);
and U20562 (N_20562,N_19355,N_19175);
xor U20563 (N_20563,N_19139,N_19362);
nor U20564 (N_20564,N_19785,N_19830);
xor U20565 (N_20565,N_19013,N_19012);
nand U20566 (N_20566,N_19932,N_19812);
xor U20567 (N_20567,N_19146,N_19682);
or U20568 (N_20568,N_19560,N_19015);
nor U20569 (N_20569,N_19640,N_19626);
nand U20570 (N_20570,N_19498,N_19728);
xnor U20571 (N_20571,N_19129,N_19559);
nor U20572 (N_20572,N_19972,N_19315);
and U20573 (N_20573,N_19872,N_19058);
xnor U20574 (N_20574,N_19779,N_19465);
or U20575 (N_20575,N_19394,N_19388);
and U20576 (N_20576,N_19364,N_19647);
and U20577 (N_20577,N_19322,N_19897);
or U20578 (N_20578,N_19707,N_19248);
or U20579 (N_20579,N_19162,N_19717);
xnor U20580 (N_20580,N_19521,N_19249);
nor U20581 (N_20581,N_19336,N_19717);
nor U20582 (N_20582,N_19774,N_19882);
xor U20583 (N_20583,N_19315,N_19765);
and U20584 (N_20584,N_19960,N_19343);
xor U20585 (N_20585,N_19749,N_19177);
nor U20586 (N_20586,N_19502,N_19366);
or U20587 (N_20587,N_19566,N_19016);
or U20588 (N_20588,N_19516,N_19832);
nor U20589 (N_20589,N_19763,N_19930);
xnor U20590 (N_20590,N_19661,N_19510);
nor U20591 (N_20591,N_19314,N_19326);
and U20592 (N_20592,N_19350,N_19636);
or U20593 (N_20593,N_19097,N_19820);
or U20594 (N_20594,N_19200,N_19442);
xor U20595 (N_20595,N_19261,N_19000);
nand U20596 (N_20596,N_19392,N_19895);
xor U20597 (N_20597,N_19203,N_19957);
xnor U20598 (N_20598,N_19104,N_19507);
xnor U20599 (N_20599,N_19170,N_19273);
or U20600 (N_20600,N_19259,N_19669);
xnor U20601 (N_20601,N_19212,N_19954);
xnor U20602 (N_20602,N_19584,N_19830);
nand U20603 (N_20603,N_19762,N_19778);
or U20604 (N_20604,N_19499,N_19026);
or U20605 (N_20605,N_19586,N_19140);
xnor U20606 (N_20606,N_19948,N_19170);
and U20607 (N_20607,N_19131,N_19883);
nand U20608 (N_20608,N_19230,N_19090);
nand U20609 (N_20609,N_19047,N_19064);
and U20610 (N_20610,N_19452,N_19508);
and U20611 (N_20611,N_19924,N_19677);
nand U20612 (N_20612,N_19417,N_19512);
or U20613 (N_20613,N_19615,N_19524);
or U20614 (N_20614,N_19504,N_19690);
and U20615 (N_20615,N_19472,N_19048);
nor U20616 (N_20616,N_19105,N_19338);
nor U20617 (N_20617,N_19349,N_19804);
or U20618 (N_20618,N_19099,N_19907);
nand U20619 (N_20619,N_19618,N_19979);
nand U20620 (N_20620,N_19060,N_19150);
and U20621 (N_20621,N_19359,N_19711);
or U20622 (N_20622,N_19435,N_19475);
nor U20623 (N_20623,N_19985,N_19741);
or U20624 (N_20624,N_19012,N_19988);
xor U20625 (N_20625,N_19156,N_19733);
nand U20626 (N_20626,N_19460,N_19188);
and U20627 (N_20627,N_19495,N_19629);
nor U20628 (N_20628,N_19848,N_19268);
xor U20629 (N_20629,N_19682,N_19161);
xor U20630 (N_20630,N_19914,N_19155);
nor U20631 (N_20631,N_19398,N_19141);
nor U20632 (N_20632,N_19312,N_19353);
nor U20633 (N_20633,N_19842,N_19320);
and U20634 (N_20634,N_19541,N_19936);
xnor U20635 (N_20635,N_19070,N_19122);
and U20636 (N_20636,N_19244,N_19769);
nor U20637 (N_20637,N_19698,N_19115);
and U20638 (N_20638,N_19751,N_19281);
and U20639 (N_20639,N_19215,N_19495);
xnor U20640 (N_20640,N_19462,N_19091);
and U20641 (N_20641,N_19668,N_19739);
nand U20642 (N_20642,N_19221,N_19890);
and U20643 (N_20643,N_19257,N_19513);
or U20644 (N_20644,N_19504,N_19932);
nor U20645 (N_20645,N_19943,N_19123);
and U20646 (N_20646,N_19040,N_19745);
and U20647 (N_20647,N_19191,N_19291);
xor U20648 (N_20648,N_19958,N_19546);
nor U20649 (N_20649,N_19137,N_19869);
xor U20650 (N_20650,N_19261,N_19136);
and U20651 (N_20651,N_19643,N_19437);
or U20652 (N_20652,N_19372,N_19931);
nor U20653 (N_20653,N_19651,N_19825);
and U20654 (N_20654,N_19258,N_19066);
nor U20655 (N_20655,N_19533,N_19269);
or U20656 (N_20656,N_19328,N_19921);
and U20657 (N_20657,N_19834,N_19095);
or U20658 (N_20658,N_19100,N_19019);
xnor U20659 (N_20659,N_19229,N_19710);
nand U20660 (N_20660,N_19615,N_19323);
xor U20661 (N_20661,N_19437,N_19333);
xor U20662 (N_20662,N_19490,N_19645);
nor U20663 (N_20663,N_19132,N_19199);
nor U20664 (N_20664,N_19782,N_19023);
xnor U20665 (N_20665,N_19612,N_19189);
nor U20666 (N_20666,N_19026,N_19273);
nor U20667 (N_20667,N_19212,N_19983);
and U20668 (N_20668,N_19933,N_19620);
nand U20669 (N_20669,N_19012,N_19512);
xnor U20670 (N_20670,N_19778,N_19546);
nor U20671 (N_20671,N_19581,N_19945);
or U20672 (N_20672,N_19013,N_19611);
or U20673 (N_20673,N_19796,N_19592);
nor U20674 (N_20674,N_19091,N_19724);
nor U20675 (N_20675,N_19051,N_19104);
nor U20676 (N_20676,N_19338,N_19013);
or U20677 (N_20677,N_19637,N_19117);
xor U20678 (N_20678,N_19966,N_19145);
or U20679 (N_20679,N_19142,N_19359);
nor U20680 (N_20680,N_19366,N_19734);
nand U20681 (N_20681,N_19886,N_19117);
or U20682 (N_20682,N_19370,N_19729);
or U20683 (N_20683,N_19466,N_19368);
or U20684 (N_20684,N_19275,N_19044);
nand U20685 (N_20685,N_19995,N_19536);
nor U20686 (N_20686,N_19852,N_19669);
or U20687 (N_20687,N_19522,N_19788);
or U20688 (N_20688,N_19043,N_19300);
xnor U20689 (N_20689,N_19792,N_19127);
nor U20690 (N_20690,N_19578,N_19974);
or U20691 (N_20691,N_19599,N_19396);
nand U20692 (N_20692,N_19593,N_19140);
nor U20693 (N_20693,N_19984,N_19378);
and U20694 (N_20694,N_19822,N_19364);
or U20695 (N_20695,N_19899,N_19777);
nor U20696 (N_20696,N_19596,N_19338);
xnor U20697 (N_20697,N_19235,N_19418);
nor U20698 (N_20698,N_19140,N_19953);
xor U20699 (N_20699,N_19681,N_19496);
nor U20700 (N_20700,N_19982,N_19948);
or U20701 (N_20701,N_19546,N_19791);
nand U20702 (N_20702,N_19102,N_19143);
and U20703 (N_20703,N_19620,N_19547);
nor U20704 (N_20704,N_19490,N_19341);
nor U20705 (N_20705,N_19456,N_19038);
and U20706 (N_20706,N_19348,N_19564);
nor U20707 (N_20707,N_19214,N_19518);
nand U20708 (N_20708,N_19232,N_19794);
xor U20709 (N_20709,N_19231,N_19017);
nor U20710 (N_20710,N_19378,N_19368);
nor U20711 (N_20711,N_19383,N_19571);
and U20712 (N_20712,N_19132,N_19861);
or U20713 (N_20713,N_19811,N_19839);
and U20714 (N_20714,N_19246,N_19303);
or U20715 (N_20715,N_19506,N_19090);
and U20716 (N_20716,N_19871,N_19181);
and U20717 (N_20717,N_19488,N_19952);
or U20718 (N_20718,N_19955,N_19217);
and U20719 (N_20719,N_19887,N_19902);
or U20720 (N_20720,N_19554,N_19017);
xor U20721 (N_20721,N_19899,N_19016);
xnor U20722 (N_20722,N_19674,N_19379);
nor U20723 (N_20723,N_19246,N_19347);
xnor U20724 (N_20724,N_19501,N_19566);
or U20725 (N_20725,N_19635,N_19192);
xor U20726 (N_20726,N_19326,N_19850);
nand U20727 (N_20727,N_19996,N_19525);
nor U20728 (N_20728,N_19451,N_19745);
and U20729 (N_20729,N_19639,N_19105);
or U20730 (N_20730,N_19532,N_19485);
nand U20731 (N_20731,N_19310,N_19036);
nor U20732 (N_20732,N_19128,N_19188);
or U20733 (N_20733,N_19789,N_19289);
nand U20734 (N_20734,N_19093,N_19434);
xnor U20735 (N_20735,N_19353,N_19177);
nor U20736 (N_20736,N_19799,N_19968);
and U20737 (N_20737,N_19453,N_19206);
xor U20738 (N_20738,N_19243,N_19468);
or U20739 (N_20739,N_19093,N_19667);
nor U20740 (N_20740,N_19307,N_19360);
and U20741 (N_20741,N_19946,N_19529);
or U20742 (N_20742,N_19990,N_19213);
xnor U20743 (N_20743,N_19773,N_19653);
or U20744 (N_20744,N_19003,N_19112);
or U20745 (N_20745,N_19481,N_19341);
or U20746 (N_20746,N_19061,N_19002);
nand U20747 (N_20747,N_19987,N_19379);
nand U20748 (N_20748,N_19457,N_19154);
nor U20749 (N_20749,N_19742,N_19504);
xnor U20750 (N_20750,N_19678,N_19055);
or U20751 (N_20751,N_19387,N_19964);
or U20752 (N_20752,N_19651,N_19377);
and U20753 (N_20753,N_19626,N_19173);
nand U20754 (N_20754,N_19950,N_19681);
and U20755 (N_20755,N_19372,N_19378);
nand U20756 (N_20756,N_19487,N_19805);
nand U20757 (N_20757,N_19598,N_19815);
and U20758 (N_20758,N_19241,N_19644);
nand U20759 (N_20759,N_19307,N_19672);
or U20760 (N_20760,N_19785,N_19791);
or U20761 (N_20761,N_19592,N_19975);
or U20762 (N_20762,N_19098,N_19789);
or U20763 (N_20763,N_19857,N_19427);
nor U20764 (N_20764,N_19186,N_19955);
nor U20765 (N_20765,N_19173,N_19597);
nand U20766 (N_20766,N_19438,N_19156);
and U20767 (N_20767,N_19160,N_19573);
nand U20768 (N_20768,N_19491,N_19106);
and U20769 (N_20769,N_19033,N_19116);
nand U20770 (N_20770,N_19372,N_19433);
and U20771 (N_20771,N_19737,N_19352);
xnor U20772 (N_20772,N_19988,N_19317);
nand U20773 (N_20773,N_19482,N_19625);
nand U20774 (N_20774,N_19842,N_19972);
xnor U20775 (N_20775,N_19275,N_19181);
nand U20776 (N_20776,N_19807,N_19194);
or U20777 (N_20777,N_19388,N_19449);
and U20778 (N_20778,N_19684,N_19276);
and U20779 (N_20779,N_19873,N_19169);
or U20780 (N_20780,N_19273,N_19659);
or U20781 (N_20781,N_19492,N_19066);
xnor U20782 (N_20782,N_19939,N_19887);
or U20783 (N_20783,N_19584,N_19854);
nor U20784 (N_20784,N_19353,N_19449);
or U20785 (N_20785,N_19503,N_19322);
nand U20786 (N_20786,N_19123,N_19645);
xnor U20787 (N_20787,N_19368,N_19440);
and U20788 (N_20788,N_19602,N_19149);
nand U20789 (N_20789,N_19377,N_19419);
nand U20790 (N_20790,N_19965,N_19340);
and U20791 (N_20791,N_19725,N_19523);
and U20792 (N_20792,N_19436,N_19773);
nor U20793 (N_20793,N_19815,N_19845);
or U20794 (N_20794,N_19115,N_19101);
nand U20795 (N_20795,N_19005,N_19028);
nand U20796 (N_20796,N_19815,N_19138);
or U20797 (N_20797,N_19227,N_19411);
xor U20798 (N_20798,N_19426,N_19442);
nand U20799 (N_20799,N_19998,N_19333);
nand U20800 (N_20800,N_19177,N_19112);
nor U20801 (N_20801,N_19133,N_19394);
nand U20802 (N_20802,N_19134,N_19367);
and U20803 (N_20803,N_19424,N_19583);
xnor U20804 (N_20804,N_19511,N_19485);
xor U20805 (N_20805,N_19744,N_19681);
xor U20806 (N_20806,N_19278,N_19412);
and U20807 (N_20807,N_19914,N_19291);
xnor U20808 (N_20808,N_19626,N_19162);
nand U20809 (N_20809,N_19105,N_19783);
or U20810 (N_20810,N_19207,N_19105);
nor U20811 (N_20811,N_19167,N_19760);
or U20812 (N_20812,N_19978,N_19092);
and U20813 (N_20813,N_19577,N_19045);
nor U20814 (N_20814,N_19508,N_19281);
and U20815 (N_20815,N_19584,N_19836);
and U20816 (N_20816,N_19012,N_19381);
xnor U20817 (N_20817,N_19277,N_19455);
nand U20818 (N_20818,N_19957,N_19732);
nor U20819 (N_20819,N_19899,N_19953);
nand U20820 (N_20820,N_19322,N_19402);
nor U20821 (N_20821,N_19768,N_19316);
and U20822 (N_20822,N_19271,N_19235);
or U20823 (N_20823,N_19500,N_19686);
or U20824 (N_20824,N_19174,N_19121);
nand U20825 (N_20825,N_19473,N_19082);
xnor U20826 (N_20826,N_19365,N_19984);
or U20827 (N_20827,N_19185,N_19908);
and U20828 (N_20828,N_19182,N_19396);
or U20829 (N_20829,N_19198,N_19401);
xor U20830 (N_20830,N_19060,N_19200);
xnor U20831 (N_20831,N_19799,N_19925);
and U20832 (N_20832,N_19429,N_19560);
nor U20833 (N_20833,N_19445,N_19090);
xor U20834 (N_20834,N_19450,N_19197);
or U20835 (N_20835,N_19506,N_19150);
nand U20836 (N_20836,N_19981,N_19025);
nor U20837 (N_20837,N_19486,N_19719);
xnor U20838 (N_20838,N_19927,N_19827);
or U20839 (N_20839,N_19464,N_19929);
or U20840 (N_20840,N_19564,N_19478);
and U20841 (N_20841,N_19463,N_19285);
xor U20842 (N_20842,N_19783,N_19156);
nand U20843 (N_20843,N_19069,N_19917);
and U20844 (N_20844,N_19148,N_19776);
and U20845 (N_20845,N_19069,N_19823);
and U20846 (N_20846,N_19722,N_19264);
nor U20847 (N_20847,N_19455,N_19050);
nor U20848 (N_20848,N_19033,N_19244);
xor U20849 (N_20849,N_19537,N_19258);
xor U20850 (N_20850,N_19591,N_19167);
nor U20851 (N_20851,N_19680,N_19171);
and U20852 (N_20852,N_19843,N_19176);
or U20853 (N_20853,N_19700,N_19784);
nand U20854 (N_20854,N_19544,N_19280);
and U20855 (N_20855,N_19355,N_19464);
nand U20856 (N_20856,N_19571,N_19068);
and U20857 (N_20857,N_19672,N_19748);
or U20858 (N_20858,N_19588,N_19035);
nor U20859 (N_20859,N_19879,N_19268);
or U20860 (N_20860,N_19937,N_19385);
nand U20861 (N_20861,N_19157,N_19022);
xnor U20862 (N_20862,N_19404,N_19298);
xor U20863 (N_20863,N_19926,N_19047);
and U20864 (N_20864,N_19679,N_19924);
nand U20865 (N_20865,N_19587,N_19417);
and U20866 (N_20866,N_19277,N_19200);
nor U20867 (N_20867,N_19915,N_19060);
nand U20868 (N_20868,N_19178,N_19142);
xor U20869 (N_20869,N_19487,N_19917);
or U20870 (N_20870,N_19888,N_19414);
and U20871 (N_20871,N_19659,N_19043);
xnor U20872 (N_20872,N_19458,N_19237);
nor U20873 (N_20873,N_19453,N_19258);
or U20874 (N_20874,N_19760,N_19570);
and U20875 (N_20875,N_19172,N_19467);
nand U20876 (N_20876,N_19063,N_19520);
nor U20877 (N_20877,N_19839,N_19022);
or U20878 (N_20878,N_19550,N_19849);
and U20879 (N_20879,N_19249,N_19278);
xor U20880 (N_20880,N_19975,N_19991);
nand U20881 (N_20881,N_19307,N_19570);
nor U20882 (N_20882,N_19276,N_19694);
nand U20883 (N_20883,N_19673,N_19713);
and U20884 (N_20884,N_19753,N_19126);
or U20885 (N_20885,N_19068,N_19041);
xor U20886 (N_20886,N_19135,N_19425);
nand U20887 (N_20887,N_19408,N_19827);
xnor U20888 (N_20888,N_19844,N_19445);
xor U20889 (N_20889,N_19692,N_19870);
xor U20890 (N_20890,N_19057,N_19762);
nor U20891 (N_20891,N_19666,N_19916);
xor U20892 (N_20892,N_19868,N_19723);
nand U20893 (N_20893,N_19237,N_19267);
nor U20894 (N_20894,N_19061,N_19351);
nand U20895 (N_20895,N_19081,N_19855);
nand U20896 (N_20896,N_19421,N_19746);
nor U20897 (N_20897,N_19293,N_19420);
or U20898 (N_20898,N_19801,N_19347);
nor U20899 (N_20899,N_19524,N_19710);
nor U20900 (N_20900,N_19868,N_19302);
nand U20901 (N_20901,N_19879,N_19238);
nand U20902 (N_20902,N_19145,N_19959);
and U20903 (N_20903,N_19700,N_19862);
nand U20904 (N_20904,N_19716,N_19036);
nand U20905 (N_20905,N_19678,N_19418);
nand U20906 (N_20906,N_19394,N_19627);
nand U20907 (N_20907,N_19515,N_19993);
xor U20908 (N_20908,N_19892,N_19338);
nand U20909 (N_20909,N_19714,N_19282);
nor U20910 (N_20910,N_19617,N_19819);
nor U20911 (N_20911,N_19749,N_19759);
and U20912 (N_20912,N_19214,N_19681);
xor U20913 (N_20913,N_19363,N_19159);
nor U20914 (N_20914,N_19644,N_19263);
and U20915 (N_20915,N_19719,N_19735);
nor U20916 (N_20916,N_19125,N_19751);
or U20917 (N_20917,N_19991,N_19788);
or U20918 (N_20918,N_19274,N_19163);
xnor U20919 (N_20919,N_19551,N_19168);
nand U20920 (N_20920,N_19202,N_19899);
nor U20921 (N_20921,N_19126,N_19113);
nor U20922 (N_20922,N_19470,N_19573);
and U20923 (N_20923,N_19096,N_19167);
nor U20924 (N_20924,N_19076,N_19282);
and U20925 (N_20925,N_19210,N_19100);
or U20926 (N_20926,N_19119,N_19716);
nor U20927 (N_20927,N_19387,N_19534);
nand U20928 (N_20928,N_19599,N_19864);
or U20929 (N_20929,N_19209,N_19317);
or U20930 (N_20930,N_19009,N_19519);
or U20931 (N_20931,N_19237,N_19651);
nand U20932 (N_20932,N_19607,N_19493);
or U20933 (N_20933,N_19061,N_19804);
and U20934 (N_20934,N_19147,N_19187);
or U20935 (N_20935,N_19644,N_19859);
nand U20936 (N_20936,N_19170,N_19581);
and U20937 (N_20937,N_19426,N_19885);
nand U20938 (N_20938,N_19284,N_19079);
or U20939 (N_20939,N_19045,N_19846);
and U20940 (N_20940,N_19710,N_19449);
nand U20941 (N_20941,N_19089,N_19088);
nor U20942 (N_20942,N_19446,N_19627);
xnor U20943 (N_20943,N_19764,N_19337);
nor U20944 (N_20944,N_19193,N_19966);
and U20945 (N_20945,N_19685,N_19248);
xnor U20946 (N_20946,N_19552,N_19282);
and U20947 (N_20947,N_19380,N_19430);
and U20948 (N_20948,N_19921,N_19340);
xnor U20949 (N_20949,N_19591,N_19622);
nand U20950 (N_20950,N_19947,N_19611);
or U20951 (N_20951,N_19569,N_19247);
nand U20952 (N_20952,N_19399,N_19139);
nand U20953 (N_20953,N_19460,N_19072);
xnor U20954 (N_20954,N_19634,N_19937);
and U20955 (N_20955,N_19416,N_19677);
or U20956 (N_20956,N_19983,N_19332);
and U20957 (N_20957,N_19768,N_19047);
nand U20958 (N_20958,N_19700,N_19407);
nor U20959 (N_20959,N_19734,N_19422);
xor U20960 (N_20960,N_19408,N_19678);
nand U20961 (N_20961,N_19094,N_19282);
xnor U20962 (N_20962,N_19912,N_19103);
and U20963 (N_20963,N_19157,N_19075);
nand U20964 (N_20964,N_19826,N_19873);
and U20965 (N_20965,N_19092,N_19862);
and U20966 (N_20966,N_19182,N_19139);
or U20967 (N_20967,N_19646,N_19647);
nand U20968 (N_20968,N_19876,N_19872);
and U20969 (N_20969,N_19444,N_19951);
or U20970 (N_20970,N_19930,N_19291);
and U20971 (N_20971,N_19089,N_19459);
or U20972 (N_20972,N_19168,N_19947);
and U20973 (N_20973,N_19766,N_19485);
and U20974 (N_20974,N_19445,N_19653);
or U20975 (N_20975,N_19281,N_19855);
nand U20976 (N_20976,N_19497,N_19624);
and U20977 (N_20977,N_19764,N_19974);
nor U20978 (N_20978,N_19833,N_19882);
nand U20979 (N_20979,N_19660,N_19938);
nor U20980 (N_20980,N_19163,N_19073);
nand U20981 (N_20981,N_19998,N_19455);
nand U20982 (N_20982,N_19546,N_19705);
or U20983 (N_20983,N_19506,N_19351);
nor U20984 (N_20984,N_19852,N_19510);
and U20985 (N_20985,N_19014,N_19153);
nand U20986 (N_20986,N_19012,N_19932);
or U20987 (N_20987,N_19451,N_19431);
nor U20988 (N_20988,N_19153,N_19969);
xor U20989 (N_20989,N_19863,N_19549);
nand U20990 (N_20990,N_19159,N_19681);
nand U20991 (N_20991,N_19875,N_19761);
xor U20992 (N_20992,N_19093,N_19223);
and U20993 (N_20993,N_19284,N_19353);
nor U20994 (N_20994,N_19721,N_19843);
nor U20995 (N_20995,N_19621,N_19975);
nor U20996 (N_20996,N_19147,N_19226);
nand U20997 (N_20997,N_19940,N_19295);
nand U20998 (N_20998,N_19486,N_19253);
and U20999 (N_20999,N_19767,N_19157);
xnor U21000 (N_21000,N_20246,N_20073);
nor U21001 (N_21001,N_20485,N_20807);
and U21002 (N_21002,N_20334,N_20927);
or U21003 (N_21003,N_20100,N_20935);
and U21004 (N_21004,N_20337,N_20095);
or U21005 (N_21005,N_20620,N_20721);
nor U21006 (N_21006,N_20134,N_20933);
xnor U21007 (N_21007,N_20143,N_20871);
xnor U21008 (N_21008,N_20266,N_20087);
nand U21009 (N_21009,N_20712,N_20790);
or U21010 (N_21010,N_20922,N_20780);
nor U21011 (N_21011,N_20473,N_20245);
xnor U21012 (N_21012,N_20235,N_20763);
nand U21013 (N_21013,N_20255,N_20068);
nand U21014 (N_21014,N_20888,N_20045);
xor U21015 (N_21015,N_20432,N_20634);
nand U21016 (N_21016,N_20328,N_20355);
nor U21017 (N_21017,N_20614,N_20331);
nand U21018 (N_21018,N_20274,N_20942);
nor U21019 (N_21019,N_20020,N_20227);
or U21020 (N_21020,N_20399,N_20768);
and U21021 (N_21021,N_20532,N_20693);
xnor U21022 (N_21022,N_20716,N_20081);
and U21023 (N_21023,N_20105,N_20875);
or U21024 (N_21024,N_20259,N_20299);
nand U21025 (N_21025,N_20155,N_20909);
xnor U21026 (N_21026,N_20581,N_20315);
nand U21027 (N_21027,N_20397,N_20044);
nand U21028 (N_21028,N_20225,N_20347);
and U21029 (N_21029,N_20421,N_20574);
or U21030 (N_21030,N_20270,N_20643);
or U21031 (N_21031,N_20603,N_20164);
and U21032 (N_21032,N_20769,N_20496);
or U21033 (N_21033,N_20236,N_20286);
or U21034 (N_21034,N_20111,N_20744);
and U21035 (N_21035,N_20356,N_20253);
nor U21036 (N_21036,N_20514,N_20625);
and U21037 (N_21037,N_20759,N_20216);
and U21038 (N_21038,N_20772,N_20316);
and U21039 (N_21039,N_20985,N_20403);
and U21040 (N_21040,N_20173,N_20362);
nor U21041 (N_21041,N_20925,N_20152);
or U21042 (N_21042,N_20953,N_20549);
and U21043 (N_21043,N_20661,N_20254);
xnor U21044 (N_21044,N_20703,N_20314);
or U21045 (N_21045,N_20615,N_20418);
xor U21046 (N_21046,N_20907,N_20836);
and U21047 (N_21047,N_20525,N_20520);
and U21048 (N_21048,N_20926,N_20709);
nand U21049 (N_21049,N_20477,N_20491);
nor U21050 (N_21050,N_20011,N_20671);
or U21051 (N_21051,N_20683,N_20470);
nor U21052 (N_21052,N_20672,N_20382);
or U21053 (N_21053,N_20506,N_20823);
xnor U21054 (N_21054,N_20770,N_20480);
and U21055 (N_21055,N_20147,N_20472);
nand U21056 (N_21056,N_20417,N_20946);
or U21057 (N_21057,N_20917,N_20032);
nand U21058 (N_21058,N_20536,N_20969);
nor U21059 (N_21059,N_20656,N_20024);
xor U21060 (N_21060,N_20552,N_20419);
nand U21061 (N_21061,N_20967,N_20080);
and U21062 (N_21062,N_20723,N_20298);
nor U21063 (N_21063,N_20320,N_20635);
or U21064 (N_21064,N_20988,N_20345);
and U21065 (N_21065,N_20715,N_20488);
or U21066 (N_21066,N_20296,N_20159);
or U21067 (N_21067,N_20700,N_20519);
xnor U21068 (N_21068,N_20069,N_20944);
or U21069 (N_21069,N_20966,N_20810);
and U21070 (N_21070,N_20384,N_20630);
and U21071 (N_21071,N_20001,N_20279);
nor U21072 (N_21072,N_20776,N_20426);
and U21073 (N_21073,N_20055,N_20596);
and U21074 (N_21074,N_20762,N_20013);
xnor U21075 (N_21075,N_20998,N_20117);
nor U21076 (N_21076,N_20075,N_20895);
or U21077 (N_21077,N_20208,N_20741);
xor U21078 (N_21078,N_20722,N_20806);
or U21079 (N_21079,N_20636,N_20214);
nor U21080 (N_21080,N_20207,N_20481);
or U21081 (N_21081,N_20198,N_20128);
nor U21082 (N_21082,N_20792,N_20711);
nor U21083 (N_21083,N_20802,N_20420);
xnor U21084 (N_21084,N_20934,N_20766);
nand U21085 (N_21085,N_20058,N_20748);
nand U21086 (N_21086,N_20775,N_20735);
nand U21087 (N_21087,N_20333,N_20789);
or U21088 (N_21088,N_20957,N_20076);
nand U21089 (N_21089,N_20017,N_20241);
or U21090 (N_21090,N_20194,N_20754);
and U21091 (N_21091,N_20510,N_20771);
nor U21092 (N_21092,N_20996,N_20070);
nor U21093 (N_21093,N_20978,N_20847);
and U21094 (N_21094,N_20023,N_20653);
or U21095 (N_21095,N_20975,N_20739);
or U21096 (N_21096,N_20457,N_20950);
xor U21097 (N_21097,N_20912,N_20434);
xnor U21098 (N_21098,N_20688,N_20446);
and U21099 (N_21099,N_20610,N_20714);
xnor U21100 (N_21100,N_20862,N_20959);
nand U21101 (N_21101,N_20827,N_20821);
or U21102 (N_21102,N_20553,N_20752);
xor U21103 (N_21103,N_20439,N_20843);
or U21104 (N_21104,N_20077,N_20006);
nor U21105 (N_21105,N_20850,N_20452);
and U21106 (N_21106,N_20025,N_20260);
or U21107 (N_21107,N_20228,N_20012);
nand U21108 (N_21108,N_20606,N_20640);
xor U21109 (N_21109,N_20995,N_20613);
nor U21110 (N_21110,N_20649,N_20889);
nor U21111 (N_21111,N_20518,N_20326);
xor U21112 (N_21112,N_20300,N_20226);
nand U21113 (N_21113,N_20000,N_20166);
xor U21114 (N_21114,N_20571,N_20358);
or U21115 (N_21115,N_20002,N_20468);
or U21116 (N_21116,N_20604,N_20018);
nor U21117 (N_21117,N_20327,N_20601);
xnor U21118 (N_21118,N_20951,N_20324);
nand U21119 (N_21119,N_20153,N_20056);
or U21120 (N_21120,N_20687,N_20037);
and U21121 (N_21121,N_20088,N_20185);
xnor U21122 (N_21122,N_20960,N_20484);
xnor U21123 (N_21123,N_20729,N_20605);
and U21124 (N_21124,N_20497,N_20199);
and U21125 (N_21125,N_20220,N_20611);
nor U21126 (N_21126,N_20212,N_20706);
and U21127 (N_21127,N_20923,N_20448);
and U21128 (N_21128,N_20513,N_20276);
or U21129 (N_21129,N_20727,N_20303);
or U21130 (N_21130,N_20047,N_20264);
nor U21131 (N_21131,N_20569,N_20961);
nor U21132 (N_21132,N_20145,N_20206);
nand U21133 (N_21133,N_20968,N_20804);
nor U21134 (N_21134,N_20502,N_20049);
or U21135 (N_21135,N_20638,N_20921);
nor U21136 (N_21136,N_20007,N_20668);
nand U21137 (N_21137,N_20425,N_20662);
and U21138 (N_21138,N_20460,N_20547);
xor U21139 (N_21139,N_20414,N_20312);
xnor U21140 (N_21140,N_20783,N_20554);
or U21141 (N_21141,N_20641,N_20781);
nor U21142 (N_21142,N_20292,N_20093);
xnor U21143 (N_21143,N_20422,N_20539);
or U21144 (N_21144,N_20224,N_20980);
or U21145 (N_21145,N_20652,N_20952);
xor U21146 (N_21146,N_20537,N_20247);
nand U21147 (N_21147,N_20118,N_20550);
and U21148 (N_21148,N_20365,N_20408);
and U21149 (N_21149,N_20778,N_20283);
nand U21150 (N_21150,N_20902,N_20677);
and U21151 (N_21151,N_20751,N_20785);
xnor U21152 (N_21152,N_20387,N_20126);
nor U21153 (N_21153,N_20191,N_20336);
and U21154 (N_21154,N_20116,N_20026);
nand U21155 (N_21155,N_20142,N_20034);
xor U21156 (N_21156,N_20915,N_20577);
xor U21157 (N_21157,N_20137,N_20738);
nor U21158 (N_21158,N_20107,N_20992);
or U21159 (N_21159,N_20555,N_20174);
and U21160 (N_21160,N_20494,N_20708);
nor U21161 (N_21161,N_20449,N_20846);
or U21162 (N_21162,N_20072,N_20628);
or U21163 (N_21163,N_20936,N_20637);
nor U21164 (N_21164,N_20830,N_20745);
nand U21165 (N_21165,N_20787,N_20750);
and U21166 (N_21166,N_20565,N_20568);
nor U21167 (N_21167,N_20021,N_20534);
nand U21168 (N_21168,N_20444,N_20913);
xor U21169 (N_21169,N_20190,N_20035);
xor U21170 (N_21170,N_20469,N_20930);
nand U21171 (N_21171,N_20788,N_20033);
or U21172 (N_21172,N_20841,N_20837);
xor U21173 (N_21173,N_20172,N_20386);
or U21174 (N_21174,N_20309,N_20083);
xor U21175 (N_21175,N_20891,N_20091);
xnor U21176 (N_21176,N_20500,N_20140);
nand U21177 (N_21177,N_20812,N_20873);
nor U21178 (N_21178,N_20391,N_20658);
xor U21179 (N_21179,N_20455,N_20808);
nand U21180 (N_21180,N_20219,N_20139);
and U21181 (N_21181,N_20991,N_20962);
xnor U21182 (N_21182,N_20433,N_20592);
nand U21183 (N_21183,N_20311,N_20607);
xnor U21184 (N_21184,N_20395,N_20517);
or U21185 (N_21185,N_20445,N_20036);
xor U21186 (N_21186,N_20119,N_20881);
nor U21187 (N_21187,N_20796,N_20731);
xor U21188 (N_21188,N_20029,N_20820);
and U21189 (N_21189,N_20949,N_20618);
and U21190 (N_21190,N_20048,N_20475);
nand U21191 (N_21191,N_20389,N_20579);
nand U21192 (N_21192,N_20878,N_20233);
nand U21193 (N_21193,N_20705,N_20619);
nand U21194 (N_21194,N_20240,N_20608);
or U21195 (N_21195,N_20645,N_20057);
nor U21196 (N_21196,N_20278,N_20101);
and U21197 (N_21197,N_20857,N_20284);
nand U21198 (N_21198,N_20261,N_20461);
nor U21199 (N_21199,N_20244,N_20740);
or U21200 (N_21200,N_20060,N_20867);
nand U21201 (N_21201,N_20123,N_20773);
nand U21202 (N_21202,N_20149,N_20492);
xor U21203 (N_21203,N_20795,N_20512);
xnor U21204 (N_21204,N_20487,N_20388);
or U21205 (N_21205,N_20318,N_20924);
or U21206 (N_21206,N_20663,N_20914);
nor U21207 (N_21207,N_20825,N_20162);
or U21208 (N_21208,N_20690,N_20970);
or U21209 (N_21209,N_20238,N_20108);
and U21210 (N_21210,N_20495,N_20993);
xor U21211 (N_21211,N_20466,N_20256);
and U21212 (N_21212,N_20374,N_20136);
nor U21213 (N_21213,N_20680,N_20218);
and U21214 (N_21214,N_20937,N_20015);
nand U21215 (N_21215,N_20815,N_20313);
and U21216 (N_21216,N_20725,N_20633);
and U21217 (N_21217,N_20588,N_20193);
xnor U21218 (N_21218,N_20416,N_20456);
xnor U21219 (N_21219,N_20590,N_20543);
and U21220 (N_21220,N_20252,N_20761);
xor U21221 (N_21221,N_20901,N_20209);
nor U21222 (N_21222,N_20258,N_20086);
xor U21223 (N_21223,N_20573,N_20732);
or U21224 (N_21224,N_20046,N_20591);
nor U21225 (N_21225,N_20660,N_20476);
nand U21226 (N_21226,N_20885,N_20308);
nor U21227 (N_21227,N_20533,N_20098);
and U21228 (N_21228,N_20053,N_20431);
or U21229 (N_21229,N_20443,N_20564);
nor U21230 (N_21230,N_20178,N_20289);
xnor U21231 (N_21231,N_20409,N_20724);
or U21232 (N_21232,N_20522,N_20490);
nand U21233 (N_21233,N_20793,N_20129);
nand U21234 (N_21234,N_20682,N_20765);
and U21235 (N_21235,N_20666,N_20281);
and U21236 (N_21236,N_20361,N_20824);
or U21237 (N_21237,N_20801,N_20749);
or U21238 (N_21238,N_20424,N_20063);
nor U21239 (N_21239,N_20064,N_20956);
and U21240 (N_21240,N_20364,N_20989);
xnor U21241 (N_21241,N_20438,N_20170);
nor U21242 (N_21242,N_20816,N_20335);
nand U21243 (N_21243,N_20521,N_20165);
and U21244 (N_21244,N_20676,N_20498);
xor U21245 (N_21245,N_20197,N_20401);
nor U21246 (N_21246,N_20883,N_20528);
and U21247 (N_21247,N_20437,N_20505);
nor U21248 (N_21248,N_20357,N_20798);
or U21249 (N_21249,N_20595,N_20965);
or U21250 (N_21250,N_20861,N_20188);
nand U21251 (N_21251,N_20657,N_20459);
or U21252 (N_21252,N_20858,N_20065);
xor U21253 (N_21253,N_20544,N_20974);
or U21254 (N_21254,N_20650,N_20042);
nand U21255 (N_21255,N_20451,N_20144);
nor U21256 (N_21256,N_20398,N_20535);
xnor U21257 (N_21257,N_20955,N_20478);
and U21258 (N_21258,N_20629,N_20849);
or U21259 (N_21259,N_20854,N_20367);
and U21260 (N_21260,N_20008,N_20231);
nand U21261 (N_21261,N_20856,N_20287);
xnor U21262 (N_21262,N_20329,N_20515);
nand U21263 (N_21263,N_20125,N_20994);
nor U21264 (N_21264,N_20039,N_20330);
nor U21265 (N_21265,N_20647,N_20339);
or U21266 (N_21266,N_20894,N_20141);
xor U21267 (N_21267,N_20538,N_20103);
nand U21268 (N_21268,N_20094,N_20866);
nand U21269 (N_21269,N_20121,N_20631);
or U21270 (N_21270,N_20919,N_20844);
and U21271 (N_21271,N_20890,N_20400);
xnor U21272 (N_21272,N_20864,N_20654);
nor U21273 (N_21273,N_20710,N_20435);
or U21274 (N_21274,N_20175,N_20192);
and U21275 (N_21275,N_20833,N_20832);
and U21276 (N_21276,N_20265,N_20644);
and U21277 (N_21277,N_20148,N_20599);
xnor U21278 (N_21278,N_20028,N_20757);
xnor U21279 (N_21279,N_20385,N_20393);
and U21280 (N_21280,N_20120,N_20349);
xnor U21281 (N_21281,N_20493,N_20523);
nor U21282 (N_21282,N_20343,N_20842);
nor U21283 (N_21283,N_20341,N_20217);
and U21284 (N_21284,N_20911,N_20089);
xor U21285 (N_21285,N_20079,N_20558);
and U21286 (N_21286,N_20288,N_20559);
or U21287 (N_21287,N_20102,N_20066);
and U21288 (N_21288,N_20051,N_20131);
or U21289 (N_21289,N_20078,N_20370);
or U21290 (N_21290,N_20753,N_20720);
nand U21291 (N_21291,N_20351,N_20378);
or U21292 (N_21292,N_20239,N_20084);
nor U21293 (N_21293,N_20737,N_20879);
nand U21294 (N_21294,N_20642,N_20784);
nand U21295 (N_21295,N_20779,N_20639);
or U21296 (N_21296,N_20582,N_20646);
nand U21297 (N_21297,N_20758,N_20003);
or U21298 (N_21298,N_20561,N_20813);
xor U21299 (N_21299,N_20305,N_20019);
and U21300 (N_21300,N_20074,N_20760);
or U21301 (N_21301,N_20267,N_20667);
xor U21302 (N_21302,N_20809,N_20584);
and U21303 (N_21303,N_20352,N_20454);
and U21304 (N_21304,N_20189,N_20504);
nor U21305 (N_21305,N_20377,N_20838);
nand U21306 (N_21306,N_20691,N_20453);
nor U21307 (N_21307,N_20109,N_20730);
and U21308 (N_21308,N_20860,N_20811);
and U21309 (N_21309,N_20171,N_20892);
nor U21310 (N_21310,N_20195,N_20943);
and U21311 (N_21311,N_20929,N_20905);
or U21312 (N_21312,N_20747,N_20132);
nor U21313 (N_21313,N_20085,N_20718);
nand U21314 (N_21314,N_20585,N_20767);
nor U21315 (N_21315,N_20229,N_20479);
xor U21316 (N_21316,N_20350,N_20627);
and U21317 (N_21317,N_20376,N_20511);
xnor U21318 (N_21318,N_20402,N_20508);
nand U21319 (N_21319,N_20407,N_20685);
or U21320 (N_21320,N_20567,N_20575);
nand U21321 (N_21321,N_20187,N_20560);
and U21322 (N_21322,N_20290,N_20791);
or U21323 (N_21323,N_20412,N_20462);
or U21324 (N_21324,N_20697,N_20692);
or U21325 (N_21325,N_20999,N_20576);
or U21326 (N_21326,N_20368,N_20133);
xnor U21327 (N_21327,N_20373,N_20509);
and U21328 (N_21328,N_20593,N_20948);
nor U21329 (N_21329,N_20851,N_20659);
and U21330 (N_21330,N_20736,N_20963);
xnor U21331 (N_21331,N_20186,N_20898);
or U21332 (N_21332,N_20797,N_20939);
or U21333 (N_21333,N_20176,N_20282);
nor U21334 (N_21334,N_20104,N_20344);
or U21335 (N_21335,N_20363,N_20160);
nor U21336 (N_21336,N_20215,N_20594);
nor U21337 (N_21337,N_20733,N_20756);
and U21338 (N_21338,N_20180,N_20516);
xnor U21339 (N_21339,N_20669,N_20548);
xnor U21340 (N_21340,N_20562,N_20423);
and U21341 (N_21341,N_20920,N_20545);
xnor U21342 (N_21342,N_20158,N_20285);
nor U21343 (N_21343,N_20410,N_20884);
nand U21344 (N_21344,N_20156,N_20067);
or U21345 (N_21345,N_20904,N_20893);
and U21346 (N_21346,N_20578,N_20230);
nand U21347 (N_21347,N_20670,N_20157);
nand U21348 (N_21348,N_20127,N_20940);
or U21349 (N_21349,N_20853,N_20719);
or U21350 (N_21350,N_20726,N_20598);
nand U21351 (N_21351,N_20200,N_20232);
nor U21352 (N_21352,N_20262,N_20202);
nor U21353 (N_21353,N_20221,N_20794);
nor U21354 (N_21354,N_20958,N_20870);
xor U21355 (N_21355,N_20698,N_20203);
xor U21356 (N_21356,N_20291,N_20876);
nor U21357 (N_21357,N_20906,N_20396);
nor U21358 (N_21358,N_20413,N_20556);
nand U21359 (N_21359,N_20293,N_20237);
nand U21360 (N_21360,N_20415,N_20673);
and U21361 (N_21361,N_20566,N_20168);
xor U21362 (N_21362,N_20899,N_20728);
nand U21363 (N_21363,N_20984,N_20301);
xnor U21364 (N_21364,N_20865,N_20005);
nor U21365 (N_21365,N_20524,N_20746);
nand U21366 (N_21366,N_20845,N_20383);
nand U21367 (N_21367,N_20234,N_20546);
and U21368 (N_21368,N_20819,N_20482);
nand U21369 (N_21369,N_20257,N_20800);
nor U21370 (N_21370,N_20931,N_20163);
xor U21371 (N_21371,N_20332,N_20271);
or U21372 (N_21372,N_20059,N_20110);
nand U21373 (N_21373,N_20348,N_20112);
nor U21374 (N_21374,N_20394,N_20831);
nor U21375 (N_21375,N_20938,N_20242);
and U21376 (N_21376,N_20755,N_20817);
and U21377 (N_21377,N_20294,N_20277);
nor U21378 (N_21378,N_20474,N_20622);
and U21379 (N_21379,N_20050,N_20828);
nor U21380 (N_21380,N_20822,N_20205);
or U21381 (N_21381,N_20135,N_20211);
and U21382 (N_21382,N_20503,N_20983);
and U21383 (N_21383,N_20406,N_20932);
nor U21384 (N_21384,N_20689,N_20447);
nor U21385 (N_21385,N_20030,N_20359);
nor U21386 (N_21386,N_20014,N_20799);
and U21387 (N_21387,N_20805,N_20179);
xnor U21388 (N_21388,N_20375,N_20243);
nor U21389 (N_21389,N_20213,N_20465);
xnor U21390 (N_21390,N_20918,N_20223);
or U21391 (N_21391,N_20609,N_20529);
xor U21392 (N_21392,N_20621,N_20874);
and U21393 (N_21393,N_20092,N_20429);
nor U21394 (N_21394,N_20530,N_20295);
and U21395 (N_21395,N_20655,N_20686);
and U21396 (N_21396,N_20353,N_20371);
nand U21397 (N_21397,N_20115,N_20675);
or U21398 (N_21398,N_20997,N_20707);
and U21399 (N_21399,N_20979,N_20346);
and U21400 (N_21400,N_20082,N_20557);
nor U21401 (N_21401,N_20713,N_20430);
and U21402 (N_21402,N_20090,N_20436);
or U21403 (N_21403,N_20183,N_20201);
or U21404 (N_21404,N_20704,N_20977);
nor U21405 (N_21405,N_20097,N_20863);
xor U21406 (N_21406,N_20269,N_20695);
xnor U21407 (N_21407,N_20304,N_20321);
nand U21408 (N_21408,N_20440,N_20678);
or U21409 (N_21409,N_20380,N_20903);
or U21410 (N_21410,N_20411,N_20222);
nand U21411 (N_21411,N_20626,N_20651);
nor U21412 (N_21412,N_20829,N_20840);
xor U21413 (N_21413,N_20004,N_20022);
or U21414 (N_21414,N_20580,N_20541);
xor U21415 (N_21415,N_20273,N_20826);
and U21416 (N_21416,N_20181,N_20325);
nor U21417 (N_21417,N_20182,N_20124);
and U21418 (N_21418,N_20501,N_20859);
nor U21419 (N_21419,N_20427,N_20317);
xnor U21420 (N_21420,N_20855,N_20319);
or U21421 (N_21421,N_20563,N_20664);
nand U21422 (N_21422,N_20322,N_20196);
or U21423 (N_21423,N_20031,N_20428);
nor U21424 (N_21424,N_20982,N_20272);
nand U21425 (N_21425,N_20210,N_20251);
nand U21426 (N_21426,N_20717,N_20010);
nand U21427 (N_21427,N_20602,N_20877);
or U21428 (N_21428,N_20062,N_20372);
nand U21429 (N_21429,N_20130,N_20947);
nor U21430 (N_21430,N_20540,N_20872);
nor U21431 (N_21431,N_20441,N_20354);
or U21432 (N_21432,N_20852,N_20586);
or U21433 (N_21433,N_20674,N_20679);
nor U21434 (N_21434,N_20150,N_20467);
nor U21435 (N_21435,N_20458,N_20551);
nor U21436 (N_21436,N_20471,N_20009);
nor U21437 (N_21437,N_20250,N_20971);
and U21438 (N_21438,N_20096,N_20887);
nor U21439 (N_21439,N_20527,N_20868);
nand U21440 (N_21440,N_20848,N_20616);
xnor U21441 (N_21441,N_20987,N_20263);
nor U21442 (N_21442,N_20138,N_20597);
and U21443 (N_21443,N_20280,N_20764);
nor U21444 (N_21444,N_20379,N_20910);
xnor U21445 (N_21445,N_20338,N_20973);
xor U21446 (N_21446,N_20169,N_20880);
nor U21447 (N_21447,N_20310,N_20834);
and U21448 (N_21448,N_20106,N_20507);
nor U21449 (N_21449,N_20099,N_20570);
xor U21450 (N_21450,N_20486,N_20990);
and U21451 (N_21451,N_20177,N_20161);
nand U21452 (N_21452,N_20648,N_20694);
nor U21453 (N_21453,N_20531,N_20945);
or U21454 (N_21454,N_20307,N_20390);
nand U21455 (N_21455,N_20743,N_20869);
xnor U21456 (N_21456,N_20572,N_20268);
and U21457 (N_21457,N_20442,N_20803);
nand U21458 (N_21458,N_20450,N_20976);
nand U21459 (N_21459,N_20151,N_20040);
nor U21460 (N_21460,N_20302,N_20665);
nor U21461 (N_21461,N_20814,N_20297);
xnor U21462 (N_21462,N_20941,N_20835);
and U21463 (N_21463,N_20886,N_20734);
nor U21464 (N_21464,N_20964,N_20323);
xor U21465 (N_21465,N_20600,N_20632);
and U21466 (N_21466,N_20340,N_20954);
and U21467 (N_21467,N_20146,N_20041);
xnor U21468 (N_21468,N_20392,N_20054);
nor U21469 (N_21469,N_20897,N_20908);
nor U21470 (N_21470,N_20916,N_20369);
xor U21471 (N_21471,N_20786,N_20617);
nand U21472 (N_21472,N_20154,N_20542);
nor U21473 (N_21473,N_20587,N_20167);
nand U21474 (N_21474,N_20612,N_20702);
xor U21475 (N_21475,N_20249,N_20061);
nand U21476 (N_21476,N_20405,N_20742);
nand U21477 (N_21477,N_20818,N_20113);
nand U21478 (N_21478,N_20366,N_20027);
xor U21479 (N_21479,N_20275,N_20464);
and U21480 (N_21480,N_20071,N_20782);
and U21481 (N_21481,N_20489,N_20204);
and U21482 (N_21482,N_20699,N_20981);
nand U21483 (N_21483,N_20928,N_20583);
or U21484 (N_21484,N_20701,N_20114);
xnor U21485 (N_21485,N_20882,N_20681);
or U21486 (N_21486,N_20184,N_20306);
or U21487 (N_21487,N_20499,N_20624);
and U21488 (N_21488,N_20777,N_20900);
and U21489 (N_21489,N_20360,N_20342);
and U21490 (N_21490,N_20381,N_20839);
or U21491 (N_21491,N_20696,N_20896);
or U21492 (N_21492,N_20684,N_20589);
xor U21493 (N_21493,N_20122,N_20463);
nand U21494 (N_21494,N_20043,N_20483);
and U21495 (N_21495,N_20774,N_20404);
xnor U21496 (N_21496,N_20052,N_20972);
nor U21497 (N_21497,N_20248,N_20986);
or U21498 (N_21498,N_20016,N_20623);
nand U21499 (N_21499,N_20526,N_20038);
or U21500 (N_21500,N_20370,N_20896);
nand U21501 (N_21501,N_20488,N_20784);
xnor U21502 (N_21502,N_20595,N_20467);
xnor U21503 (N_21503,N_20182,N_20289);
nand U21504 (N_21504,N_20835,N_20240);
nand U21505 (N_21505,N_20426,N_20769);
xnor U21506 (N_21506,N_20693,N_20155);
and U21507 (N_21507,N_20929,N_20510);
xor U21508 (N_21508,N_20034,N_20017);
xnor U21509 (N_21509,N_20166,N_20462);
nor U21510 (N_21510,N_20641,N_20083);
xor U21511 (N_21511,N_20621,N_20051);
or U21512 (N_21512,N_20380,N_20523);
nand U21513 (N_21513,N_20411,N_20010);
or U21514 (N_21514,N_20722,N_20754);
nor U21515 (N_21515,N_20397,N_20740);
or U21516 (N_21516,N_20328,N_20092);
and U21517 (N_21517,N_20840,N_20736);
xnor U21518 (N_21518,N_20833,N_20230);
or U21519 (N_21519,N_20697,N_20967);
nor U21520 (N_21520,N_20680,N_20076);
nand U21521 (N_21521,N_20568,N_20232);
and U21522 (N_21522,N_20666,N_20246);
nor U21523 (N_21523,N_20365,N_20293);
or U21524 (N_21524,N_20194,N_20917);
xnor U21525 (N_21525,N_20061,N_20866);
and U21526 (N_21526,N_20752,N_20759);
or U21527 (N_21527,N_20349,N_20501);
nand U21528 (N_21528,N_20998,N_20249);
nand U21529 (N_21529,N_20285,N_20238);
and U21530 (N_21530,N_20673,N_20373);
or U21531 (N_21531,N_20915,N_20103);
or U21532 (N_21532,N_20242,N_20510);
and U21533 (N_21533,N_20242,N_20073);
xor U21534 (N_21534,N_20824,N_20083);
nor U21535 (N_21535,N_20756,N_20827);
xnor U21536 (N_21536,N_20144,N_20386);
or U21537 (N_21537,N_20789,N_20991);
or U21538 (N_21538,N_20690,N_20476);
xnor U21539 (N_21539,N_20412,N_20840);
nor U21540 (N_21540,N_20340,N_20425);
nand U21541 (N_21541,N_20869,N_20669);
xnor U21542 (N_21542,N_20580,N_20209);
and U21543 (N_21543,N_20841,N_20947);
nor U21544 (N_21544,N_20573,N_20441);
xnor U21545 (N_21545,N_20533,N_20807);
nand U21546 (N_21546,N_20902,N_20222);
xnor U21547 (N_21547,N_20852,N_20654);
nor U21548 (N_21548,N_20398,N_20980);
nand U21549 (N_21549,N_20122,N_20004);
and U21550 (N_21550,N_20809,N_20044);
nand U21551 (N_21551,N_20530,N_20706);
or U21552 (N_21552,N_20459,N_20261);
or U21553 (N_21553,N_20820,N_20522);
and U21554 (N_21554,N_20370,N_20500);
or U21555 (N_21555,N_20709,N_20849);
nand U21556 (N_21556,N_20767,N_20307);
xnor U21557 (N_21557,N_20111,N_20882);
xnor U21558 (N_21558,N_20673,N_20687);
nor U21559 (N_21559,N_20449,N_20218);
and U21560 (N_21560,N_20123,N_20342);
nand U21561 (N_21561,N_20144,N_20429);
xor U21562 (N_21562,N_20000,N_20247);
and U21563 (N_21563,N_20324,N_20049);
xnor U21564 (N_21564,N_20220,N_20114);
or U21565 (N_21565,N_20345,N_20288);
or U21566 (N_21566,N_20603,N_20902);
or U21567 (N_21567,N_20945,N_20291);
nand U21568 (N_21568,N_20804,N_20832);
xnor U21569 (N_21569,N_20161,N_20282);
xor U21570 (N_21570,N_20719,N_20372);
or U21571 (N_21571,N_20357,N_20155);
nand U21572 (N_21572,N_20824,N_20775);
nand U21573 (N_21573,N_20288,N_20099);
and U21574 (N_21574,N_20207,N_20864);
nand U21575 (N_21575,N_20657,N_20988);
xnor U21576 (N_21576,N_20802,N_20946);
nor U21577 (N_21577,N_20079,N_20252);
xnor U21578 (N_21578,N_20324,N_20668);
nand U21579 (N_21579,N_20446,N_20786);
and U21580 (N_21580,N_20395,N_20659);
nand U21581 (N_21581,N_20845,N_20156);
and U21582 (N_21582,N_20735,N_20996);
and U21583 (N_21583,N_20236,N_20694);
xor U21584 (N_21584,N_20192,N_20440);
nand U21585 (N_21585,N_20403,N_20630);
nand U21586 (N_21586,N_20578,N_20113);
and U21587 (N_21587,N_20143,N_20641);
nand U21588 (N_21588,N_20154,N_20408);
or U21589 (N_21589,N_20312,N_20199);
nor U21590 (N_21590,N_20645,N_20437);
xor U21591 (N_21591,N_20882,N_20902);
xor U21592 (N_21592,N_20293,N_20646);
and U21593 (N_21593,N_20407,N_20938);
xnor U21594 (N_21594,N_20169,N_20685);
xnor U21595 (N_21595,N_20511,N_20444);
and U21596 (N_21596,N_20650,N_20916);
nor U21597 (N_21597,N_20925,N_20679);
and U21598 (N_21598,N_20785,N_20610);
and U21599 (N_21599,N_20945,N_20334);
or U21600 (N_21600,N_20988,N_20955);
and U21601 (N_21601,N_20283,N_20723);
xnor U21602 (N_21602,N_20188,N_20865);
nand U21603 (N_21603,N_20733,N_20523);
or U21604 (N_21604,N_20904,N_20432);
and U21605 (N_21605,N_20018,N_20620);
and U21606 (N_21606,N_20304,N_20541);
or U21607 (N_21607,N_20507,N_20121);
xor U21608 (N_21608,N_20962,N_20803);
nand U21609 (N_21609,N_20737,N_20097);
and U21610 (N_21610,N_20249,N_20777);
or U21611 (N_21611,N_20819,N_20910);
or U21612 (N_21612,N_20332,N_20375);
nand U21613 (N_21613,N_20330,N_20218);
xnor U21614 (N_21614,N_20897,N_20368);
nor U21615 (N_21615,N_20200,N_20850);
xor U21616 (N_21616,N_20520,N_20413);
xor U21617 (N_21617,N_20441,N_20140);
nor U21618 (N_21618,N_20032,N_20595);
nor U21619 (N_21619,N_20640,N_20524);
nor U21620 (N_21620,N_20601,N_20550);
xnor U21621 (N_21621,N_20309,N_20555);
nor U21622 (N_21622,N_20619,N_20986);
nor U21623 (N_21623,N_20898,N_20411);
and U21624 (N_21624,N_20451,N_20980);
nor U21625 (N_21625,N_20806,N_20178);
and U21626 (N_21626,N_20652,N_20444);
nand U21627 (N_21627,N_20357,N_20690);
nand U21628 (N_21628,N_20493,N_20980);
or U21629 (N_21629,N_20047,N_20336);
and U21630 (N_21630,N_20780,N_20626);
or U21631 (N_21631,N_20506,N_20608);
nor U21632 (N_21632,N_20961,N_20500);
xor U21633 (N_21633,N_20937,N_20516);
and U21634 (N_21634,N_20333,N_20259);
nand U21635 (N_21635,N_20357,N_20538);
or U21636 (N_21636,N_20044,N_20668);
and U21637 (N_21637,N_20095,N_20549);
or U21638 (N_21638,N_20672,N_20522);
xnor U21639 (N_21639,N_20648,N_20972);
xnor U21640 (N_21640,N_20493,N_20020);
xor U21641 (N_21641,N_20346,N_20614);
xnor U21642 (N_21642,N_20075,N_20149);
and U21643 (N_21643,N_20518,N_20403);
xnor U21644 (N_21644,N_20867,N_20049);
nand U21645 (N_21645,N_20893,N_20090);
nand U21646 (N_21646,N_20714,N_20320);
xnor U21647 (N_21647,N_20726,N_20781);
or U21648 (N_21648,N_20084,N_20649);
nor U21649 (N_21649,N_20792,N_20642);
xor U21650 (N_21650,N_20021,N_20935);
nor U21651 (N_21651,N_20661,N_20061);
nand U21652 (N_21652,N_20467,N_20178);
nor U21653 (N_21653,N_20917,N_20207);
nand U21654 (N_21654,N_20496,N_20382);
or U21655 (N_21655,N_20032,N_20839);
or U21656 (N_21656,N_20004,N_20726);
or U21657 (N_21657,N_20639,N_20468);
or U21658 (N_21658,N_20310,N_20885);
nor U21659 (N_21659,N_20075,N_20232);
xnor U21660 (N_21660,N_20631,N_20723);
and U21661 (N_21661,N_20976,N_20950);
nor U21662 (N_21662,N_20426,N_20888);
and U21663 (N_21663,N_20598,N_20669);
nand U21664 (N_21664,N_20423,N_20520);
nand U21665 (N_21665,N_20369,N_20448);
or U21666 (N_21666,N_20159,N_20072);
and U21667 (N_21667,N_20983,N_20484);
or U21668 (N_21668,N_20651,N_20901);
xor U21669 (N_21669,N_20601,N_20195);
nor U21670 (N_21670,N_20318,N_20488);
nand U21671 (N_21671,N_20004,N_20637);
and U21672 (N_21672,N_20446,N_20080);
or U21673 (N_21673,N_20727,N_20366);
xnor U21674 (N_21674,N_20038,N_20988);
and U21675 (N_21675,N_20425,N_20300);
xor U21676 (N_21676,N_20920,N_20967);
nand U21677 (N_21677,N_20470,N_20187);
or U21678 (N_21678,N_20373,N_20526);
nand U21679 (N_21679,N_20928,N_20977);
xnor U21680 (N_21680,N_20687,N_20653);
or U21681 (N_21681,N_20622,N_20833);
or U21682 (N_21682,N_20346,N_20829);
and U21683 (N_21683,N_20313,N_20912);
and U21684 (N_21684,N_20758,N_20789);
nand U21685 (N_21685,N_20769,N_20578);
nand U21686 (N_21686,N_20966,N_20943);
or U21687 (N_21687,N_20872,N_20096);
nor U21688 (N_21688,N_20576,N_20127);
nor U21689 (N_21689,N_20867,N_20891);
xor U21690 (N_21690,N_20125,N_20674);
and U21691 (N_21691,N_20302,N_20760);
nand U21692 (N_21692,N_20548,N_20499);
and U21693 (N_21693,N_20441,N_20743);
and U21694 (N_21694,N_20080,N_20416);
nand U21695 (N_21695,N_20942,N_20306);
nand U21696 (N_21696,N_20722,N_20618);
nand U21697 (N_21697,N_20920,N_20127);
xnor U21698 (N_21698,N_20192,N_20243);
and U21699 (N_21699,N_20775,N_20216);
xor U21700 (N_21700,N_20636,N_20528);
nand U21701 (N_21701,N_20439,N_20115);
nand U21702 (N_21702,N_20678,N_20364);
nor U21703 (N_21703,N_20442,N_20573);
xor U21704 (N_21704,N_20967,N_20040);
nand U21705 (N_21705,N_20265,N_20990);
xnor U21706 (N_21706,N_20485,N_20871);
xor U21707 (N_21707,N_20369,N_20719);
and U21708 (N_21708,N_20415,N_20958);
or U21709 (N_21709,N_20104,N_20826);
xnor U21710 (N_21710,N_20199,N_20022);
nor U21711 (N_21711,N_20561,N_20112);
nor U21712 (N_21712,N_20744,N_20742);
or U21713 (N_21713,N_20909,N_20353);
nand U21714 (N_21714,N_20128,N_20464);
xnor U21715 (N_21715,N_20470,N_20706);
xor U21716 (N_21716,N_20615,N_20867);
nor U21717 (N_21717,N_20113,N_20434);
and U21718 (N_21718,N_20684,N_20061);
nor U21719 (N_21719,N_20492,N_20926);
nor U21720 (N_21720,N_20007,N_20901);
nor U21721 (N_21721,N_20809,N_20764);
nor U21722 (N_21722,N_20872,N_20293);
nand U21723 (N_21723,N_20205,N_20443);
nand U21724 (N_21724,N_20239,N_20703);
and U21725 (N_21725,N_20802,N_20059);
or U21726 (N_21726,N_20033,N_20205);
xor U21727 (N_21727,N_20908,N_20162);
xor U21728 (N_21728,N_20920,N_20690);
and U21729 (N_21729,N_20318,N_20996);
and U21730 (N_21730,N_20877,N_20090);
nor U21731 (N_21731,N_20364,N_20066);
and U21732 (N_21732,N_20407,N_20219);
nor U21733 (N_21733,N_20052,N_20937);
or U21734 (N_21734,N_20760,N_20277);
nand U21735 (N_21735,N_20143,N_20893);
or U21736 (N_21736,N_20499,N_20780);
nor U21737 (N_21737,N_20216,N_20683);
nand U21738 (N_21738,N_20514,N_20380);
and U21739 (N_21739,N_20618,N_20244);
and U21740 (N_21740,N_20417,N_20542);
or U21741 (N_21741,N_20846,N_20792);
or U21742 (N_21742,N_20274,N_20266);
nand U21743 (N_21743,N_20552,N_20151);
nand U21744 (N_21744,N_20721,N_20532);
xor U21745 (N_21745,N_20681,N_20511);
and U21746 (N_21746,N_20469,N_20796);
and U21747 (N_21747,N_20860,N_20985);
and U21748 (N_21748,N_20644,N_20885);
xor U21749 (N_21749,N_20468,N_20359);
and U21750 (N_21750,N_20964,N_20130);
or U21751 (N_21751,N_20776,N_20385);
or U21752 (N_21752,N_20107,N_20117);
or U21753 (N_21753,N_20202,N_20621);
nand U21754 (N_21754,N_20493,N_20950);
nand U21755 (N_21755,N_20130,N_20321);
xor U21756 (N_21756,N_20482,N_20633);
xnor U21757 (N_21757,N_20656,N_20689);
nor U21758 (N_21758,N_20150,N_20719);
or U21759 (N_21759,N_20733,N_20968);
and U21760 (N_21760,N_20339,N_20596);
xor U21761 (N_21761,N_20467,N_20121);
nand U21762 (N_21762,N_20758,N_20537);
or U21763 (N_21763,N_20684,N_20607);
nor U21764 (N_21764,N_20037,N_20299);
nand U21765 (N_21765,N_20669,N_20081);
or U21766 (N_21766,N_20366,N_20446);
or U21767 (N_21767,N_20372,N_20209);
nand U21768 (N_21768,N_20679,N_20455);
nor U21769 (N_21769,N_20940,N_20158);
and U21770 (N_21770,N_20472,N_20646);
or U21771 (N_21771,N_20505,N_20741);
and U21772 (N_21772,N_20942,N_20421);
nor U21773 (N_21773,N_20762,N_20590);
xnor U21774 (N_21774,N_20159,N_20018);
xor U21775 (N_21775,N_20460,N_20806);
or U21776 (N_21776,N_20577,N_20191);
or U21777 (N_21777,N_20807,N_20875);
nor U21778 (N_21778,N_20934,N_20676);
or U21779 (N_21779,N_20617,N_20744);
xnor U21780 (N_21780,N_20473,N_20021);
nand U21781 (N_21781,N_20232,N_20526);
nand U21782 (N_21782,N_20836,N_20430);
nand U21783 (N_21783,N_20191,N_20087);
or U21784 (N_21784,N_20368,N_20231);
and U21785 (N_21785,N_20387,N_20432);
xor U21786 (N_21786,N_20078,N_20423);
xnor U21787 (N_21787,N_20171,N_20753);
and U21788 (N_21788,N_20711,N_20769);
and U21789 (N_21789,N_20849,N_20660);
and U21790 (N_21790,N_20193,N_20475);
nand U21791 (N_21791,N_20110,N_20382);
or U21792 (N_21792,N_20795,N_20022);
xnor U21793 (N_21793,N_20604,N_20190);
and U21794 (N_21794,N_20934,N_20829);
xor U21795 (N_21795,N_20882,N_20247);
and U21796 (N_21796,N_20916,N_20829);
xor U21797 (N_21797,N_20318,N_20759);
or U21798 (N_21798,N_20866,N_20194);
nor U21799 (N_21799,N_20100,N_20397);
or U21800 (N_21800,N_20206,N_20461);
or U21801 (N_21801,N_20019,N_20551);
xnor U21802 (N_21802,N_20887,N_20760);
and U21803 (N_21803,N_20038,N_20009);
or U21804 (N_21804,N_20960,N_20517);
nor U21805 (N_21805,N_20191,N_20830);
and U21806 (N_21806,N_20099,N_20497);
xor U21807 (N_21807,N_20307,N_20715);
or U21808 (N_21808,N_20421,N_20933);
nor U21809 (N_21809,N_20937,N_20002);
and U21810 (N_21810,N_20618,N_20582);
or U21811 (N_21811,N_20075,N_20908);
nand U21812 (N_21812,N_20554,N_20522);
xor U21813 (N_21813,N_20980,N_20301);
nand U21814 (N_21814,N_20792,N_20450);
xor U21815 (N_21815,N_20038,N_20869);
or U21816 (N_21816,N_20775,N_20033);
xor U21817 (N_21817,N_20516,N_20278);
and U21818 (N_21818,N_20262,N_20038);
nand U21819 (N_21819,N_20631,N_20717);
or U21820 (N_21820,N_20961,N_20488);
nand U21821 (N_21821,N_20089,N_20045);
nor U21822 (N_21822,N_20142,N_20721);
nor U21823 (N_21823,N_20781,N_20985);
or U21824 (N_21824,N_20975,N_20486);
nand U21825 (N_21825,N_20154,N_20911);
nor U21826 (N_21826,N_20773,N_20131);
or U21827 (N_21827,N_20765,N_20113);
and U21828 (N_21828,N_20042,N_20213);
nand U21829 (N_21829,N_20971,N_20754);
or U21830 (N_21830,N_20010,N_20354);
or U21831 (N_21831,N_20474,N_20565);
nor U21832 (N_21832,N_20057,N_20476);
or U21833 (N_21833,N_20462,N_20361);
xor U21834 (N_21834,N_20272,N_20837);
xnor U21835 (N_21835,N_20829,N_20110);
or U21836 (N_21836,N_20031,N_20431);
nand U21837 (N_21837,N_20683,N_20886);
nor U21838 (N_21838,N_20742,N_20658);
and U21839 (N_21839,N_20966,N_20020);
xnor U21840 (N_21840,N_20352,N_20944);
and U21841 (N_21841,N_20626,N_20258);
and U21842 (N_21842,N_20326,N_20078);
and U21843 (N_21843,N_20853,N_20175);
or U21844 (N_21844,N_20952,N_20053);
xor U21845 (N_21845,N_20705,N_20059);
nor U21846 (N_21846,N_20378,N_20754);
xnor U21847 (N_21847,N_20801,N_20169);
xor U21848 (N_21848,N_20153,N_20594);
xnor U21849 (N_21849,N_20017,N_20799);
or U21850 (N_21850,N_20448,N_20190);
or U21851 (N_21851,N_20386,N_20747);
nand U21852 (N_21852,N_20915,N_20022);
nand U21853 (N_21853,N_20762,N_20560);
xor U21854 (N_21854,N_20579,N_20185);
nor U21855 (N_21855,N_20216,N_20283);
nand U21856 (N_21856,N_20096,N_20763);
xnor U21857 (N_21857,N_20134,N_20994);
nand U21858 (N_21858,N_20494,N_20681);
or U21859 (N_21859,N_20278,N_20876);
nand U21860 (N_21860,N_20677,N_20422);
nor U21861 (N_21861,N_20756,N_20520);
nand U21862 (N_21862,N_20244,N_20692);
xor U21863 (N_21863,N_20363,N_20197);
and U21864 (N_21864,N_20379,N_20841);
and U21865 (N_21865,N_20110,N_20340);
nand U21866 (N_21866,N_20925,N_20295);
xor U21867 (N_21867,N_20735,N_20130);
nor U21868 (N_21868,N_20549,N_20011);
nand U21869 (N_21869,N_20740,N_20777);
and U21870 (N_21870,N_20691,N_20410);
nor U21871 (N_21871,N_20871,N_20236);
nor U21872 (N_21872,N_20042,N_20147);
and U21873 (N_21873,N_20551,N_20452);
nor U21874 (N_21874,N_20143,N_20839);
or U21875 (N_21875,N_20975,N_20618);
xnor U21876 (N_21876,N_20568,N_20199);
nand U21877 (N_21877,N_20814,N_20684);
or U21878 (N_21878,N_20385,N_20387);
nand U21879 (N_21879,N_20172,N_20516);
nor U21880 (N_21880,N_20038,N_20041);
or U21881 (N_21881,N_20338,N_20866);
xor U21882 (N_21882,N_20523,N_20060);
and U21883 (N_21883,N_20271,N_20311);
xor U21884 (N_21884,N_20063,N_20811);
and U21885 (N_21885,N_20398,N_20246);
and U21886 (N_21886,N_20681,N_20939);
nand U21887 (N_21887,N_20341,N_20907);
nand U21888 (N_21888,N_20729,N_20191);
nand U21889 (N_21889,N_20132,N_20460);
or U21890 (N_21890,N_20851,N_20222);
nand U21891 (N_21891,N_20670,N_20907);
nand U21892 (N_21892,N_20616,N_20511);
nor U21893 (N_21893,N_20676,N_20249);
xor U21894 (N_21894,N_20311,N_20603);
nor U21895 (N_21895,N_20221,N_20701);
nor U21896 (N_21896,N_20642,N_20173);
xor U21897 (N_21897,N_20920,N_20534);
nor U21898 (N_21898,N_20864,N_20418);
xnor U21899 (N_21899,N_20501,N_20374);
and U21900 (N_21900,N_20343,N_20669);
xnor U21901 (N_21901,N_20290,N_20526);
nor U21902 (N_21902,N_20750,N_20267);
nor U21903 (N_21903,N_20925,N_20359);
xnor U21904 (N_21904,N_20456,N_20194);
nor U21905 (N_21905,N_20701,N_20542);
nor U21906 (N_21906,N_20028,N_20842);
and U21907 (N_21907,N_20723,N_20514);
xnor U21908 (N_21908,N_20520,N_20054);
and U21909 (N_21909,N_20298,N_20935);
nor U21910 (N_21910,N_20726,N_20943);
nor U21911 (N_21911,N_20143,N_20097);
nand U21912 (N_21912,N_20019,N_20529);
nand U21913 (N_21913,N_20103,N_20764);
nand U21914 (N_21914,N_20278,N_20588);
nor U21915 (N_21915,N_20508,N_20226);
and U21916 (N_21916,N_20804,N_20579);
nor U21917 (N_21917,N_20829,N_20215);
or U21918 (N_21918,N_20995,N_20740);
xor U21919 (N_21919,N_20354,N_20173);
xnor U21920 (N_21920,N_20432,N_20978);
or U21921 (N_21921,N_20154,N_20682);
nor U21922 (N_21922,N_20618,N_20187);
nand U21923 (N_21923,N_20127,N_20098);
or U21924 (N_21924,N_20610,N_20589);
and U21925 (N_21925,N_20360,N_20819);
nand U21926 (N_21926,N_20439,N_20186);
and U21927 (N_21927,N_20874,N_20122);
nor U21928 (N_21928,N_20208,N_20081);
and U21929 (N_21929,N_20675,N_20908);
or U21930 (N_21930,N_20069,N_20666);
nor U21931 (N_21931,N_20200,N_20171);
or U21932 (N_21932,N_20470,N_20223);
and U21933 (N_21933,N_20041,N_20483);
or U21934 (N_21934,N_20727,N_20866);
and U21935 (N_21935,N_20330,N_20255);
nand U21936 (N_21936,N_20729,N_20808);
nor U21937 (N_21937,N_20620,N_20962);
nand U21938 (N_21938,N_20472,N_20164);
nand U21939 (N_21939,N_20857,N_20803);
and U21940 (N_21940,N_20126,N_20169);
nor U21941 (N_21941,N_20427,N_20858);
nor U21942 (N_21942,N_20031,N_20479);
nor U21943 (N_21943,N_20059,N_20221);
and U21944 (N_21944,N_20177,N_20609);
and U21945 (N_21945,N_20885,N_20068);
nand U21946 (N_21946,N_20858,N_20401);
nor U21947 (N_21947,N_20962,N_20451);
and U21948 (N_21948,N_20632,N_20900);
nor U21949 (N_21949,N_20787,N_20591);
xor U21950 (N_21950,N_20494,N_20095);
or U21951 (N_21951,N_20107,N_20816);
nor U21952 (N_21952,N_20896,N_20886);
nand U21953 (N_21953,N_20192,N_20314);
xor U21954 (N_21954,N_20686,N_20233);
nand U21955 (N_21955,N_20721,N_20374);
nand U21956 (N_21956,N_20573,N_20075);
nand U21957 (N_21957,N_20433,N_20419);
nand U21958 (N_21958,N_20032,N_20921);
nor U21959 (N_21959,N_20687,N_20586);
or U21960 (N_21960,N_20045,N_20412);
or U21961 (N_21961,N_20930,N_20129);
xor U21962 (N_21962,N_20398,N_20539);
or U21963 (N_21963,N_20856,N_20245);
nor U21964 (N_21964,N_20767,N_20923);
or U21965 (N_21965,N_20287,N_20076);
nand U21966 (N_21966,N_20919,N_20782);
or U21967 (N_21967,N_20809,N_20052);
and U21968 (N_21968,N_20644,N_20784);
or U21969 (N_21969,N_20348,N_20748);
nand U21970 (N_21970,N_20900,N_20145);
or U21971 (N_21971,N_20275,N_20910);
nand U21972 (N_21972,N_20778,N_20169);
or U21973 (N_21973,N_20916,N_20889);
nand U21974 (N_21974,N_20635,N_20136);
xnor U21975 (N_21975,N_20526,N_20939);
and U21976 (N_21976,N_20085,N_20136);
nor U21977 (N_21977,N_20813,N_20264);
xnor U21978 (N_21978,N_20512,N_20432);
or U21979 (N_21979,N_20672,N_20317);
nand U21980 (N_21980,N_20797,N_20145);
nand U21981 (N_21981,N_20710,N_20652);
nor U21982 (N_21982,N_20295,N_20929);
or U21983 (N_21983,N_20128,N_20158);
nor U21984 (N_21984,N_20959,N_20065);
nand U21985 (N_21985,N_20532,N_20190);
xnor U21986 (N_21986,N_20651,N_20274);
nand U21987 (N_21987,N_20239,N_20675);
xnor U21988 (N_21988,N_20046,N_20066);
nand U21989 (N_21989,N_20483,N_20447);
or U21990 (N_21990,N_20384,N_20946);
and U21991 (N_21991,N_20889,N_20920);
nor U21992 (N_21992,N_20366,N_20751);
nand U21993 (N_21993,N_20275,N_20069);
and U21994 (N_21994,N_20642,N_20811);
nand U21995 (N_21995,N_20576,N_20366);
nand U21996 (N_21996,N_20154,N_20575);
nor U21997 (N_21997,N_20055,N_20608);
or U21998 (N_21998,N_20257,N_20350);
nand U21999 (N_21999,N_20840,N_20664);
nand U22000 (N_22000,N_21853,N_21829);
and U22001 (N_22001,N_21336,N_21975);
and U22002 (N_22002,N_21688,N_21894);
and U22003 (N_22003,N_21966,N_21800);
nor U22004 (N_22004,N_21370,N_21376);
and U22005 (N_22005,N_21458,N_21302);
or U22006 (N_22006,N_21816,N_21416);
xor U22007 (N_22007,N_21731,N_21826);
or U22008 (N_22008,N_21264,N_21553);
xor U22009 (N_22009,N_21864,N_21722);
nand U22010 (N_22010,N_21385,N_21533);
and U22011 (N_22011,N_21981,N_21954);
xnor U22012 (N_22012,N_21228,N_21283);
nor U22013 (N_22013,N_21477,N_21292);
nor U22014 (N_22014,N_21271,N_21601);
nor U22015 (N_22015,N_21665,N_21298);
nor U22016 (N_22016,N_21166,N_21708);
or U22017 (N_22017,N_21782,N_21639);
xor U22018 (N_22018,N_21532,N_21592);
xor U22019 (N_22019,N_21783,N_21739);
nand U22020 (N_22020,N_21487,N_21658);
and U22021 (N_22021,N_21801,N_21990);
xnor U22022 (N_22022,N_21939,N_21721);
nor U22023 (N_22023,N_21220,N_21326);
nand U22024 (N_22024,N_21539,N_21199);
nand U22025 (N_22025,N_21439,N_21677);
or U22026 (N_22026,N_21243,N_21896);
and U22027 (N_22027,N_21834,N_21471);
or U22028 (N_22028,N_21707,N_21420);
nor U22029 (N_22029,N_21261,N_21647);
or U22030 (N_22030,N_21158,N_21673);
and U22031 (N_22031,N_21219,N_21106);
and U22032 (N_22032,N_21361,N_21053);
and U22033 (N_22033,N_21769,N_21702);
xnor U22034 (N_22034,N_21167,N_21478);
xor U22035 (N_22035,N_21656,N_21317);
or U22036 (N_22036,N_21107,N_21987);
and U22037 (N_22037,N_21935,N_21664);
or U22038 (N_22038,N_21996,N_21484);
xor U22039 (N_22039,N_21295,N_21010);
xnor U22040 (N_22040,N_21367,N_21549);
xnor U22041 (N_22041,N_21171,N_21156);
xnor U22042 (N_22042,N_21511,N_21129);
nand U22043 (N_22043,N_21610,N_21852);
and U22044 (N_22044,N_21431,N_21470);
or U22045 (N_22045,N_21191,N_21644);
nor U22046 (N_22046,N_21615,N_21718);
nor U22047 (N_22047,N_21895,N_21161);
or U22048 (N_22048,N_21402,N_21753);
xor U22049 (N_22049,N_21081,N_21200);
nor U22050 (N_22050,N_21841,N_21071);
and U22051 (N_22051,N_21960,N_21066);
or U22052 (N_22052,N_21537,N_21133);
nor U22053 (N_22053,N_21555,N_21248);
xor U22054 (N_22054,N_21510,N_21744);
nor U22055 (N_22055,N_21837,N_21629);
or U22056 (N_22056,N_21775,N_21715);
and U22057 (N_22057,N_21189,N_21284);
or U22058 (N_22058,N_21903,N_21092);
nand U22059 (N_22059,N_21922,N_21565);
and U22060 (N_22060,N_21872,N_21597);
and U22061 (N_22061,N_21230,N_21029);
or U22062 (N_22062,N_21719,N_21277);
or U22063 (N_22063,N_21031,N_21689);
or U22064 (N_22064,N_21022,N_21464);
and U22065 (N_22065,N_21595,N_21232);
nand U22066 (N_22066,N_21598,N_21341);
or U22067 (N_22067,N_21324,N_21860);
xor U22068 (N_22068,N_21803,N_21737);
xor U22069 (N_22069,N_21596,N_21907);
and U22070 (N_22070,N_21999,N_21176);
or U22071 (N_22071,N_21509,N_21818);
and U22072 (N_22072,N_21440,N_21628);
or U22073 (N_22073,N_21157,N_21560);
and U22074 (N_22074,N_21934,N_21641);
and U22075 (N_22075,N_21006,N_21869);
xor U22076 (N_22076,N_21705,N_21774);
nor U22077 (N_22077,N_21172,N_21884);
or U22078 (N_22078,N_21337,N_21952);
nand U22079 (N_22079,N_21983,N_21997);
and U22080 (N_22080,N_21246,N_21923);
nand U22081 (N_22081,N_21086,N_21977);
or U22082 (N_22082,N_21388,N_21300);
and U22083 (N_22083,N_21461,N_21181);
xnor U22084 (N_22084,N_21384,N_21058);
and U22085 (N_22085,N_21048,N_21141);
nor U22086 (N_22086,N_21512,N_21459);
nand U22087 (N_22087,N_21968,N_21832);
xnor U22088 (N_22088,N_21185,N_21674);
and U22089 (N_22089,N_21480,N_21550);
xnor U22090 (N_22090,N_21498,N_21584);
nand U22091 (N_22091,N_21383,N_21415);
and U22092 (N_22092,N_21606,N_21957);
or U22093 (N_22093,N_21055,N_21469);
xor U22094 (N_22094,N_21237,N_21716);
nor U22095 (N_22095,N_21779,N_21563);
nor U22096 (N_22096,N_21661,N_21136);
or U22097 (N_22097,N_21362,N_21492);
and U22098 (N_22098,N_21519,N_21898);
or U22099 (N_22099,N_21871,N_21706);
xor U22100 (N_22100,N_21881,N_21720);
nand U22101 (N_22101,N_21486,N_21211);
or U22102 (N_22102,N_21877,N_21238);
xor U22103 (N_22103,N_21016,N_21789);
nand U22104 (N_22104,N_21426,N_21148);
xor U22105 (N_22105,N_21710,N_21137);
xnor U22106 (N_22106,N_21224,N_21638);
or U22107 (N_22107,N_21807,N_21585);
or U22108 (N_22108,N_21620,N_21698);
and U22109 (N_22109,N_21085,N_21114);
or U22110 (N_22110,N_21034,N_21989);
and U22111 (N_22111,N_21493,N_21712);
and U22112 (N_22112,N_21495,N_21462);
or U22113 (N_22113,N_21540,N_21182);
nor U22114 (N_22114,N_21848,N_21036);
xor U22115 (N_22115,N_21235,N_21334);
or U22116 (N_22116,N_21032,N_21150);
nand U22117 (N_22117,N_21355,N_21963);
or U22118 (N_22118,N_21578,N_21339);
xnor U22119 (N_22119,N_21475,N_21918);
xnor U22120 (N_22120,N_21733,N_21736);
or U22121 (N_22121,N_21692,N_21504);
or U22122 (N_22122,N_21076,N_21748);
and U22123 (N_22123,N_21303,N_21310);
xor U22124 (N_22124,N_21075,N_21763);
xor U22125 (N_22125,N_21056,N_21988);
and U22126 (N_22126,N_21602,N_21915);
and U22127 (N_22127,N_21955,N_21932);
and U22128 (N_22128,N_21521,N_21589);
and U22129 (N_22129,N_21855,N_21645);
and U22130 (N_22130,N_21472,N_21522);
and U22131 (N_22131,N_21695,N_21242);
nand U22132 (N_22132,N_21924,N_21659);
or U22133 (N_22133,N_21322,N_21282);
nand U22134 (N_22134,N_21704,N_21179);
nand U22135 (N_22135,N_21164,N_21587);
and U22136 (N_22136,N_21770,N_21364);
or U22137 (N_22137,N_21314,N_21691);
xnor U22138 (N_22138,N_21212,N_21494);
nor U22139 (N_22139,N_21503,N_21218);
and U22140 (N_22140,N_21173,N_21759);
nor U22141 (N_22141,N_21274,N_21613);
nand U22142 (N_22142,N_21128,N_21350);
xor U22143 (N_22143,N_21079,N_21815);
xnor U22144 (N_22144,N_21103,N_21417);
or U22145 (N_22145,N_21208,N_21541);
and U22146 (N_22146,N_21299,N_21259);
nand U22147 (N_22147,N_21247,N_21657);
nand U22148 (N_22148,N_21023,N_21139);
nand U22149 (N_22149,N_21389,N_21594);
and U22150 (N_22150,N_21378,N_21073);
nand U22151 (N_22151,N_21184,N_21045);
xnor U22152 (N_22152,N_21885,N_21979);
xor U22153 (N_22153,N_21944,N_21352);
nor U22154 (N_22154,N_21743,N_21140);
or U22155 (N_22155,N_21751,N_21011);
or U22156 (N_22156,N_21328,N_21080);
and U22157 (N_22157,N_21529,N_21660);
xor U22158 (N_22158,N_21279,N_21059);
or U22159 (N_22159,N_21198,N_21926);
or U22160 (N_22160,N_21791,N_21348);
nor U22161 (N_22161,N_21395,N_21091);
xor U22162 (N_22162,N_21887,N_21570);
nor U22163 (N_22163,N_21687,N_21856);
or U22164 (N_22164,N_21608,N_21531);
nand U22165 (N_22165,N_21125,N_21343);
nand U22166 (N_22166,N_21929,N_21973);
nand U22167 (N_22167,N_21202,N_21667);
nor U22168 (N_22168,N_21857,N_21094);
xor U22169 (N_22169,N_21342,N_21825);
or U22170 (N_22170,N_21307,N_21183);
nor U22171 (N_22171,N_21456,N_21497);
nand U22172 (N_22172,N_21393,N_21870);
xnor U22173 (N_22173,N_21646,N_21758);
xor U22174 (N_22174,N_21001,N_21483);
nor U22175 (N_22175,N_21703,N_21412);
nand U22176 (N_22176,N_21113,N_21254);
and U22177 (N_22177,N_21734,N_21377);
nand U22178 (N_22178,N_21285,N_21488);
and U22179 (N_22179,N_21382,N_21481);
nand U22180 (N_22180,N_21095,N_21294);
and U22181 (N_22181,N_21245,N_21580);
or U22182 (N_22182,N_21306,N_21672);
nand U22183 (N_22183,N_21528,N_21162);
or U22184 (N_22184,N_21003,N_21234);
nand U22185 (N_22185,N_21479,N_21649);
or U22186 (N_22186,N_21700,N_21399);
or U22187 (N_22187,N_21270,N_21757);
xor U22188 (N_22188,N_21018,N_21159);
and U22189 (N_22189,N_21305,N_21077);
and U22190 (N_22190,N_21177,N_21227);
xnor U22191 (N_22191,N_21397,N_21313);
and U22192 (N_22192,N_21709,N_21724);
nand U22193 (N_22193,N_21950,N_21210);
xor U22194 (N_22194,N_21226,N_21956);
nor U22195 (N_22195,N_21363,N_21526);
xnor U22196 (N_22196,N_21216,N_21192);
nor U22197 (N_22197,N_21214,N_21090);
nor U22198 (N_22198,N_21831,N_21976);
nor U22199 (N_22199,N_21680,N_21463);
and U22200 (N_22200,N_21400,N_21040);
xor U22201 (N_22201,N_21043,N_21222);
nand U22202 (N_22202,N_21686,N_21605);
xor U22203 (N_22203,N_21804,N_21122);
and U22204 (N_22204,N_21061,N_21905);
nor U22205 (N_22205,N_21108,N_21930);
or U22206 (N_22206,N_21046,N_21749);
xor U22207 (N_22207,N_21438,N_21675);
or U22208 (N_22208,N_21648,N_21862);
nor U22209 (N_22209,N_21845,N_21728);
nor U22210 (N_22210,N_21943,N_21683);
or U22211 (N_22211,N_21787,N_21972);
and U22212 (N_22212,N_21111,N_21369);
nand U22213 (N_22213,N_21784,N_21165);
nand U22214 (N_22214,N_21250,N_21145);
xor U22215 (N_22215,N_21696,N_21941);
nand U22216 (N_22216,N_21600,N_21586);
or U22217 (N_22217,N_21229,N_21714);
nand U22218 (N_22218,N_21699,N_21514);
xor U22219 (N_22219,N_21795,N_21747);
xor U22220 (N_22220,N_21265,N_21231);
nand U22221 (N_22221,N_21876,N_21269);
or U22222 (N_22222,N_21499,N_21899);
and U22223 (N_22223,N_21293,N_21882);
nor U22224 (N_22224,N_21636,N_21655);
nor U22225 (N_22225,N_21886,N_21335);
xor U22226 (N_22226,N_21599,N_21102);
nand U22227 (N_22227,N_21682,N_21117);
or U22228 (N_22228,N_21255,N_21788);
or U22229 (N_22229,N_21315,N_21275);
xor U22230 (N_22230,N_21785,N_21132);
nand U22231 (N_22231,N_21823,N_21821);
nand U22232 (N_22232,N_21154,N_21917);
xor U22233 (N_22233,N_21945,N_21515);
nand U22234 (N_22234,N_21505,N_21604);
and U22235 (N_22235,N_21065,N_21062);
xor U22236 (N_22236,N_21304,N_21513);
and U22237 (N_22237,N_21365,N_21217);
and U22238 (N_22238,N_21017,N_21266);
xnor U22239 (N_22239,N_21776,N_21101);
and U22240 (N_22240,N_21349,N_21379);
and U22241 (N_22241,N_21865,N_21033);
nand U22242 (N_22242,N_21225,N_21742);
nor U22243 (N_22243,N_21735,N_21603);
xnor U22244 (N_22244,N_21811,N_21021);
nor U22245 (N_22245,N_21233,N_21418);
xnor U22246 (N_22246,N_21067,N_21196);
nand U22247 (N_22247,N_21962,N_21965);
xor U22248 (N_22248,N_21491,N_21442);
nand U22249 (N_22249,N_21617,N_21750);
or U22250 (N_22250,N_21760,N_21490);
xnor U22251 (N_22251,N_21407,N_21567);
or U22252 (N_22252,N_21566,N_21425);
and U22253 (N_22253,N_21391,N_21288);
xor U22254 (N_22254,N_21878,N_21556);
xnor U22255 (N_22255,N_21007,N_21449);
nand U22256 (N_22256,N_21590,N_21452);
nor U22257 (N_22257,N_21790,N_21741);
nor U22258 (N_22258,N_21901,N_21465);
or U22259 (N_22259,N_21916,N_21340);
nand U22260 (N_22260,N_21851,N_21518);
nor U22261 (N_22261,N_21197,N_21174);
nand U22262 (N_22262,N_21535,N_21195);
nor U22263 (N_22263,N_21263,N_21398);
xnor U22264 (N_22264,N_21879,N_21588);
and U22265 (N_22265,N_21296,N_21621);
and U22266 (N_22266,N_21039,N_21701);
nand U22267 (N_22267,N_21347,N_21612);
xnor U22268 (N_22268,N_21726,N_21429);
nand U22269 (N_22269,N_21571,N_21890);
and U22270 (N_22270,N_21051,N_21467);
xnor U22271 (N_22271,N_21893,N_21839);
and U22272 (N_22272,N_21037,N_21558);
and U22273 (N_22273,N_21764,N_21013);
nand U22274 (N_22274,N_21631,N_21931);
nand U22275 (N_22275,N_21244,N_21386);
or U22276 (N_22276,N_21793,N_21151);
or U22277 (N_22277,N_21445,N_21074);
nor U22278 (N_22278,N_21951,N_21408);
xnor U22279 (N_22279,N_21551,N_21523);
nor U22280 (N_22280,N_21543,N_21502);
and U22281 (N_22281,N_21969,N_21614);
nor U22282 (N_22282,N_21685,N_21766);
or U22283 (N_22283,N_21097,N_21024);
nor U22284 (N_22284,N_21506,N_21912);
or U22285 (N_22285,N_21607,N_21520);
xnor U22286 (N_22286,N_21451,N_21180);
xnor U22287 (N_22287,N_21557,N_21489);
nor U22288 (N_22288,N_21914,N_21538);
nor U22289 (N_22289,N_21536,N_21327);
nor U22290 (N_22290,N_21260,N_21149);
nor U22291 (N_22291,N_21160,N_21118);
nor U22292 (N_22292,N_21297,N_21119);
and U22293 (N_22293,N_21762,N_21325);
nor U22294 (N_22294,N_21863,N_21640);
xor U22295 (N_22295,N_21994,N_21444);
and U22296 (N_22296,N_21135,N_21875);
nand U22297 (N_22297,N_21430,N_21880);
or U22298 (N_22298,N_21373,N_21690);
xnor U22299 (N_22299,N_21933,N_21980);
or U22300 (N_22300,N_21666,N_21581);
nor U22301 (N_22301,N_21205,N_21711);
or U22302 (N_22302,N_21047,N_21593);
and U22303 (N_22303,N_21725,N_21846);
and U22304 (N_22304,N_21971,N_21679);
and U22305 (N_22305,N_21781,N_21552);
xor U22306 (N_22306,N_21651,N_21168);
xnor U22307 (N_22307,N_21730,N_21146);
nor U22308 (N_22308,N_21240,N_21262);
nand U22309 (N_22309,N_21188,N_21088);
xnor U22310 (N_22310,N_21542,N_21100);
and U22311 (N_22311,N_21946,N_21115);
nand U22312 (N_22312,N_21874,N_21850);
nor U22313 (N_22313,N_21561,N_21170);
nor U22314 (N_22314,N_21249,N_21959);
and U22315 (N_22315,N_21669,N_21568);
xor U22316 (N_22316,N_21153,N_21267);
and U22317 (N_22317,N_21802,N_21681);
nor U22318 (N_22318,N_21403,N_21792);
and U22319 (N_22319,N_21995,N_21799);
nand U22320 (N_22320,N_21911,N_21050);
nand U22321 (N_22321,N_21241,N_21359);
or U22322 (N_22322,N_21970,N_21019);
or U22323 (N_22323,N_21671,N_21676);
or U22324 (N_22324,N_21193,N_21654);
nand U22325 (N_22325,N_21009,N_21072);
nor U22326 (N_22326,N_21508,N_21138);
nor U22327 (N_22327,N_21842,N_21986);
xor U22328 (N_22328,N_21413,N_21474);
or U22329 (N_22329,N_21866,N_21330);
nand U22330 (N_22330,N_21252,N_21213);
xor U22331 (N_22331,N_21311,N_21632);
nand U22332 (N_22332,N_21745,N_21353);
and U22333 (N_22333,N_21559,N_21308);
and U22334 (N_22334,N_21668,N_21372);
nor U22335 (N_22335,N_21466,N_21134);
and U22336 (N_22336,N_21754,N_21419);
nand U22337 (N_22337,N_21187,N_21358);
nor U22338 (N_22338,N_21859,N_21404);
xor U22339 (N_22339,N_21796,N_21028);
xor U22340 (N_22340,N_21717,N_21063);
or U22341 (N_22341,N_21321,N_21152);
nor U22342 (N_22342,N_21756,N_21268);
nand U22343 (N_22343,N_21190,N_21947);
and U22344 (N_22344,N_21889,N_21847);
xor U22345 (N_22345,N_21083,N_21366);
xnor U22346 (N_22346,N_21333,N_21752);
xor U22347 (N_22347,N_21131,N_21354);
or U22348 (N_22348,N_21958,N_21390);
nand U22349 (N_22349,N_21096,N_21993);
and U22350 (N_22350,N_21124,N_21435);
or U22351 (N_22351,N_21000,N_21982);
nor U22352 (N_22352,N_21064,N_21808);
or U22353 (N_22353,N_21178,N_21287);
nor U22354 (N_22354,N_21814,N_21583);
nand U22355 (N_22355,N_21794,N_21253);
xnor U22356 (N_22356,N_21500,N_21099);
xnor U22357 (N_22357,N_21574,N_21964);
nor U22358 (N_22358,N_21309,N_21127);
or U22359 (N_22359,N_21272,N_21052);
nand U22360 (N_22360,N_21175,N_21098);
or U22361 (N_22361,N_21371,N_21109);
nand U22362 (N_22362,N_21454,N_21446);
xor U22363 (N_22363,N_21809,N_21992);
xor U22364 (N_22364,N_21937,N_21069);
xnor U22365 (N_22365,N_21961,N_21761);
xor U22366 (N_22366,N_21280,N_21624);
nand U22367 (N_22367,N_21819,N_21949);
or U22368 (N_22368,N_21653,N_21286);
xor U22369 (N_22369,N_21394,N_21093);
or U22370 (N_22370,N_21281,N_21836);
xnor U22371 (N_22371,N_21374,N_21693);
or U22372 (N_22372,N_21273,N_21025);
nand U22373 (N_22373,N_21057,N_21723);
or U22374 (N_22374,N_21729,N_21546);
nand U22375 (N_22375,N_21323,N_21356);
and U22376 (N_22376,N_21833,N_21611);
or U22377 (N_22377,N_21545,N_21078);
nor U22378 (N_22378,N_21562,N_21392);
and U22379 (N_22379,N_21437,N_21633);
nor U22380 (N_22380,N_21577,N_21768);
and U22381 (N_22381,N_21824,N_21888);
and U22382 (N_22382,N_21038,N_21974);
or U22383 (N_22383,N_21547,N_21998);
or U22384 (N_22384,N_21517,N_21978);
nor U22385 (N_22385,N_21116,N_21643);
nor U22386 (N_22386,N_21256,N_21854);
or U22387 (N_22387,N_21591,N_21953);
nand U22388 (N_22388,N_21068,N_21920);
or U22389 (N_22389,N_21530,N_21110);
xnor U22390 (N_22390,N_21448,N_21817);
or U22391 (N_22391,N_21991,N_21421);
xor U22392 (N_22392,N_21873,N_21121);
and U22393 (N_22393,N_21209,N_21634);
or U22394 (N_22394,N_21527,N_21312);
and U22395 (N_22395,N_21004,N_21460);
nand U22396 (N_22396,N_21401,N_21618);
nor U22397 (N_22397,N_21123,N_21927);
xor U22398 (N_22398,N_21380,N_21027);
xnor U22399 (N_22399,N_21858,N_21206);
nor U22400 (N_22400,N_21482,N_21221);
xnor U22401 (N_22401,N_21396,N_21316);
nor U22402 (N_22402,N_21130,N_21433);
xnor U22403 (N_22403,N_21332,N_21186);
xor U22404 (N_22404,N_21575,N_21967);
or U22405 (N_22405,N_21650,N_21485);
xor U22406 (N_22406,N_21453,N_21375);
or U22407 (N_22407,N_21070,N_21126);
and U22408 (N_22408,N_21773,N_21891);
xnor U22409 (N_22409,N_21236,N_21662);
xnor U22410 (N_22410,N_21910,N_21544);
or U22411 (N_22411,N_21900,N_21319);
and U22412 (N_22412,N_21622,N_21838);
nand U22413 (N_22413,N_21331,N_21169);
nor U22414 (N_22414,N_21525,N_21548);
xor U22415 (N_22415,N_21642,N_21805);
and U22416 (N_22416,N_21904,N_21105);
nand U22417 (N_22417,N_21663,N_21201);
and U22418 (N_22418,N_21940,N_21501);
nor U22419 (N_22419,N_21534,N_21777);
nor U22420 (N_22420,N_21861,N_21427);
and U22421 (N_22421,N_21616,N_21827);
nand U22422 (N_22422,N_21868,N_21928);
nand U22423 (N_22423,N_21713,N_21849);
or U22424 (N_22424,N_21345,N_21609);
and U22425 (N_22425,N_21434,N_21089);
and U22426 (N_22426,N_21694,N_21360);
nand U22427 (N_22427,N_21812,N_21573);
and U22428 (N_22428,N_21806,N_21797);
nand U22429 (N_22429,N_21516,N_21147);
xor U22430 (N_22430,N_21780,N_21697);
nor U22431 (N_22431,N_21044,N_21258);
nor U22432 (N_22432,N_21767,N_21630);
or U22433 (N_22433,N_21625,N_21441);
xnor U22434 (N_22434,N_21087,N_21740);
xor U22435 (N_22435,N_21450,N_21828);
xor U22436 (N_22436,N_21985,N_21251);
nand U22437 (N_22437,N_21572,N_21443);
nand U22438 (N_22438,N_21042,N_21919);
and U22439 (N_22439,N_21942,N_21938);
nor U22440 (N_22440,N_21948,N_21030);
xor U22441 (N_22441,N_21346,N_21468);
or U22442 (N_22442,N_21289,N_21223);
xnor U22443 (N_22443,N_21344,N_21627);
or U22444 (N_22444,N_21897,N_21778);
or U22445 (N_22445,N_21652,N_21329);
or U22446 (N_22446,N_21002,N_21084);
and U22447 (N_22447,N_21772,N_21867);
xor U22448 (N_22448,N_21432,N_21422);
and U22449 (N_22449,N_21921,N_21005);
or U22450 (N_22450,N_21423,N_21883);
or U22451 (N_22451,N_21357,N_21755);
and U22452 (N_22452,N_21060,N_21844);
and U22453 (N_22453,N_21194,N_21635);
nand U22454 (N_22454,N_21405,N_21409);
or U22455 (N_22455,N_21381,N_21155);
or U22456 (N_22456,N_21020,N_21623);
nand U22457 (N_22457,N_21015,N_21727);
or U22458 (N_22458,N_21320,N_21524);
nor U22459 (N_22459,N_21239,N_21902);
xor U22460 (N_22460,N_21843,N_21582);
or U22461 (N_22461,N_21908,N_21626);
xor U22462 (N_22462,N_21008,N_21082);
or U22463 (N_22463,N_21142,N_21351);
nor U22464 (N_22464,N_21746,N_21207);
xor U22465 (N_22465,N_21112,N_21765);
and U22466 (N_22466,N_21455,N_21054);
nand U22467 (N_22467,N_21906,N_21012);
nand U22468 (N_22468,N_21318,N_21840);
or U22469 (N_22469,N_21569,N_21496);
xnor U22470 (N_22470,N_21041,N_21411);
xnor U22471 (N_22471,N_21406,N_21909);
nor U22472 (N_22472,N_21203,N_21771);
xnor U22473 (N_22473,N_21936,N_21368);
xor U22474 (N_22474,N_21798,N_21338);
nand U22475 (N_22475,N_21301,N_21822);
nor U22476 (N_22476,N_21447,N_21424);
nand U22477 (N_22477,N_21144,N_21564);
or U22478 (N_22478,N_21143,N_21436);
and U22479 (N_22479,N_21120,N_21913);
nand U22480 (N_22480,N_21554,N_21835);
xnor U22481 (N_22481,N_21257,N_21278);
xnor U22482 (N_22482,N_21507,N_21414);
nor U22483 (N_22483,N_21457,N_21035);
nand U22484 (N_22484,N_21290,N_21984);
and U22485 (N_22485,N_21892,N_21276);
and U22486 (N_22486,N_21291,N_21684);
or U22487 (N_22487,N_21738,N_21473);
xnor U22488 (N_22488,N_21619,N_21163);
nand U22489 (N_22489,N_21925,N_21670);
nand U22490 (N_22490,N_21813,N_21428);
or U22491 (N_22491,N_21830,N_21810);
or U22492 (N_22492,N_21387,N_21678);
xnor U22493 (N_22493,N_21637,N_21820);
and U22494 (N_22494,N_21204,N_21026);
xnor U22495 (N_22495,N_21579,N_21786);
nand U22496 (N_22496,N_21476,N_21104);
nor U22497 (N_22497,N_21732,N_21215);
and U22498 (N_22498,N_21049,N_21576);
nand U22499 (N_22499,N_21014,N_21410);
xnor U22500 (N_22500,N_21283,N_21976);
and U22501 (N_22501,N_21542,N_21287);
nand U22502 (N_22502,N_21713,N_21064);
nor U22503 (N_22503,N_21313,N_21902);
and U22504 (N_22504,N_21433,N_21921);
and U22505 (N_22505,N_21615,N_21548);
or U22506 (N_22506,N_21978,N_21311);
xor U22507 (N_22507,N_21697,N_21935);
nand U22508 (N_22508,N_21838,N_21683);
xnor U22509 (N_22509,N_21682,N_21055);
xor U22510 (N_22510,N_21427,N_21588);
or U22511 (N_22511,N_21483,N_21655);
or U22512 (N_22512,N_21052,N_21502);
nand U22513 (N_22513,N_21900,N_21234);
or U22514 (N_22514,N_21262,N_21621);
nand U22515 (N_22515,N_21548,N_21090);
xnor U22516 (N_22516,N_21670,N_21780);
xnor U22517 (N_22517,N_21170,N_21823);
and U22518 (N_22518,N_21703,N_21671);
or U22519 (N_22519,N_21846,N_21131);
nand U22520 (N_22520,N_21622,N_21307);
and U22521 (N_22521,N_21312,N_21191);
and U22522 (N_22522,N_21635,N_21530);
nand U22523 (N_22523,N_21314,N_21999);
or U22524 (N_22524,N_21211,N_21973);
xnor U22525 (N_22525,N_21355,N_21797);
or U22526 (N_22526,N_21219,N_21788);
nor U22527 (N_22527,N_21849,N_21336);
nand U22528 (N_22528,N_21530,N_21440);
nand U22529 (N_22529,N_21312,N_21814);
or U22530 (N_22530,N_21523,N_21861);
and U22531 (N_22531,N_21890,N_21064);
xor U22532 (N_22532,N_21446,N_21303);
or U22533 (N_22533,N_21310,N_21198);
or U22534 (N_22534,N_21981,N_21415);
xnor U22535 (N_22535,N_21285,N_21310);
nand U22536 (N_22536,N_21020,N_21927);
xor U22537 (N_22537,N_21194,N_21362);
nand U22538 (N_22538,N_21993,N_21258);
and U22539 (N_22539,N_21065,N_21685);
nor U22540 (N_22540,N_21645,N_21228);
and U22541 (N_22541,N_21576,N_21235);
xnor U22542 (N_22542,N_21403,N_21463);
and U22543 (N_22543,N_21355,N_21947);
nor U22544 (N_22544,N_21079,N_21449);
xnor U22545 (N_22545,N_21146,N_21856);
xor U22546 (N_22546,N_21297,N_21686);
or U22547 (N_22547,N_21641,N_21727);
xor U22548 (N_22548,N_21488,N_21646);
or U22549 (N_22549,N_21156,N_21386);
and U22550 (N_22550,N_21388,N_21810);
nor U22551 (N_22551,N_21537,N_21034);
and U22552 (N_22552,N_21295,N_21646);
or U22553 (N_22553,N_21375,N_21173);
nand U22554 (N_22554,N_21281,N_21230);
nand U22555 (N_22555,N_21077,N_21335);
xor U22556 (N_22556,N_21716,N_21862);
nor U22557 (N_22557,N_21899,N_21440);
nand U22558 (N_22558,N_21009,N_21342);
xor U22559 (N_22559,N_21131,N_21682);
and U22560 (N_22560,N_21223,N_21115);
and U22561 (N_22561,N_21414,N_21778);
nand U22562 (N_22562,N_21991,N_21473);
nand U22563 (N_22563,N_21264,N_21254);
nand U22564 (N_22564,N_21466,N_21003);
or U22565 (N_22565,N_21136,N_21889);
or U22566 (N_22566,N_21245,N_21778);
xor U22567 (N_22567,N_21585,N_21678);
nand U22568 (N_22568,N_21825,N_21589);
and U22569 (N_22569,N_21755,N_21970);
xnor U22570 (N_22570,N_21486,N_21440);
and U22571 (N_22571,N_21677,N_21210);
nor U22572 (N_22572,N_21773,N_21593);
or U22573 (N_22573,N_21353,N_21597);
and U22574 (N_22574,N_21982,N_21999);
nand U22575 (N_22575,N_21878,N_21672);
xnor U22576 (N_22576,N_21418,N_21764);
nor U22577 (N_22577,N_21006,N_21984);
and U22578 (N_22578,N_21592,N_21106);
or U22579 (N_22579,N_21718,N_21688);
nor U22580 (N_22580,N_21296,N_21669);
nor U22581 (N_22581,N_21875,N_21296);
and U22582 (N_22582,N_21534,N_21270);
xnor U22583 (N_22583,N_21092,N_21897);
or U22584 (N_22584,N_21244,N_21880);
and U22585 (N_22585,N_21626,N_21984);
nor U22586 (N_22586,N_21920,N_21493);
xnor U22587 (N_22587,N_21929,N_21327);
nand U22588 (N_22588,N_21339,N_21267);
nor U22589 (N_22589,N_21369,N_21597);
or U22590 (N_22590,N_21709,N_21881);
xor U22591 (N_22591,N_21485,N_21514);
xor U22592 (N_22592,N_21303,N_21817);
and U22593 (N_22593,N_21264,N_21029);
nor U22594 (N_22594,N_21764,N_21519);
or U22595 (N_22595,N_21803,N_21576);
nand U22596 (N_22596,N_21236,N_21360);
or U22597 (N_22597,N_21355,N_21408);
xor U22598 (N_22598,N_21336,N_21322);
nor U22599 (N_22599,N_21505,N_21764);
nand U22600 (N_22600,N_21067,N_21901);
xor U22601 (N_22601,N_21459,N_21602);
xnor U22602 (N_22602,N_21868,N_21000);
and U22603 (N_22603,N_21863,N_21655);
or U22604 (N_22604,N_21431,N_21364);
xnor U22605 (N_22605,N_21240,N_21736);
or U22606 (N_22606,N_21091,N_21925);
or U22607 (N_22607,N_21827,N_21437);
xor U22608 (N_22608,N_21297,N_21698);
xnor U22609 (N_22609,N_21013,N_21515);
nor U22610 (N_22610,N_21073,N_21652);
nand U22611 (N_22611,N_21766,N_21425);
and U22612 (N_22612,N_21701,N_21817);
or U22613 (N_22613,N_21910,N_21986);
xnor U22614 (N_22614,N_21228,N_21830);
nand U22615 (N_22615,N_21962,N_21185);
xor U22616 (N_22616,N_21149,N_21543);
and U22617 (N_22617,N_21469,N_21077);
and U22618 (N_22618,N_21082,N_21507);
or U22619 (N_22619,N_21474,N_21960);
or U22620 (N_22620,N_21238,N_21922);
and U22621 (N_22621,N_21616,N_21586);
or U22622 (N_22622,N_21642,N_21471);
nand U22623 (N_22623,N_21119,N_21549);
or U22624 (N_22624,N_21829,N_21505);
or U22625 (N_22625,N_21706,N_21838);
nand U22626 (N_22626,N_21597,N_21199);
xor U22627 (N_22627,N_21370,N_21864);
or U22628 (N_22628,N_21653,N_21841);
nand U22629 (N_22629,N_21526,N_21688);
nand U22630 (N_22630,N_21207,N_21379);
or U22631 (N_22631,N_21200,N_21297);
nor U22632 (N_22632,N_21301,N_21864);
or U22633 (N_22633,N_21790,N_21592);
nor U22634 (N_22634,N_21851,N_21007);
xnor U22635 (N_22635,N_21761,N_21269);
and U22636 (N_22636,N_21701,N_21808);
nor U22637 (N_22637,N_21830,N_21332);
xor U22638 (N_22638,N_21711,N_21856);
xor U22639 (N_22639,N_21530,N_21660);
or U22640 (N_22640,N_21990,N_21339);
nor U22641 (N_22641,N_21727,N_21653);
nor U22642 (N_22642,N_21143,N_21791);
or U22643 (N_22643,N_21790,N_21457);
xnor U22644 (N_22644,N_21056,N_21763);
nand U22645 (N_22645,N_21527,N_21032);
and U22646 (N_22646,N_21425,N_21225);
nor U22647 (N_22647,N_21705,N_21725);
nor U22648 (N_22648,N_21087,N_21809);
xnor U22649 (N_22649,N_21896,N_21448);
and U22650 (N_22650,N_21267,N_21475);
nand U22651 (N_22651,N_21436,N_21927);
nor U22652 (N_22652,N_21393,N_21986);
and U22653 (N_22653,N_21025,N_21811);
and U22654 (N_22654,N_21755,N_21577);
nand U22655 (N_22655,N_21271,N_21290);
or U22656 (N_22656,N_21593,N_21807);
and U22657 (N_22657,N_21593,N_21390);
nor U22658 (N_22658,N_21813,N_21039);
xnor U22659 (N_22659,N_21691,N_21557);
or U22660 (N_22660,N_21976,N_21408);
or U22661 (N_22661,N_21033,N_21762);
nor U22662 (N_22662,N_21589,N_21209);
nand U22663 (N_22663,N_21413,N_21332);
nand U22664 (N_22664,N_21174,N_21000);
nand U22665 (N_22665,N_21880,N_21781);
nand U22666 (N_22666,N_21677,N_21652);
nor U22667 (N_22667,N_21732,N_21667);
nand U22668 (N_22668,N_21418,N_21845);
and U22669 (N_22669,N_21032,N_21874);
xor U22670 (N_22670,N_21068,N_21984);
nor U22671 (N_22671,N_21276,N_21495);
nand U22672 (N_22672,N_21262,N_21859);
xor U22673 (N_22673,N_21026,N_21429);
or U22674 (N_22674,N_21995,N_21521);
nor U22675 (N_22675,N_21320,N_21952);
xor U22676 (N_22676,N_21785,N_21731);
xor U22677 (N_22677,N_21748,N_21422);
nand U22678 (N_22678,N_21746,N_21949);
nor U22679 (N_22679,N_21894,N_21405);
nor U22680 (N_22680,N_21506,N_21575);
or U22681 (N_22681,N_21384,N_21479);
xor U22682 (N_22682,N_21237,N_21758);
xor U22683 (N_22683,N_21931,N_21887);
and U22684 (N_22684,N_21214,N_21577);
and U22685 (N_22685,N_21013,N_21128);
and U22686 (N_22686,N_21957,N_21455);
xor U22687 (N_22687,N_21867,N_21278);
nor U22688 (N_22688,N_21593,N_21186);
nand U22689 (N_22689,N_21470,N_21114);
xor U22690 (N_22690,N_21925,N_21858);
or U22691 (N_22691,N_21279,N_21900);
or U22692 (N_22692,N_21328,N_21800);
nand U22693 (N_22693,N_21763,N_21000);
xor U22694 (N_22694,N_21862,N_21045);
and U22695 (N_22695,N_21590,N_21588);
nor U22696 (N_22696,N_21299,N_21821);
nor U22697 (N_22697,N_21153,N_21832);
nor U22698 (N_22698,N_21441,N_21298);
nand U22699 (N_22699,N_21515,N_21351);
xnor U22700 (N_22700,N_21999,N_21041);
or U22701 (N_22701,N_21241,N_21280);
and U22702 (N_22702,N_21521,N_21081);
xnor U22703 (N_22703,N_21180,N_21473);
nor U22704 (N_22704,N_21641,N_21517);
and U22705 (N_22705,N_21167,N_21809);
xnor U22706 (N_22706,N_21923,N_21266);
xor U22707 (N_22707,N_21468,N_21000);
and U22708 (N_22708,N_21975,N_21030);
xnor U22709 (N_22709,N_21182,N_21495);
or U22710 (N_22710,N_21987,N_21399);
or U22711 (N_22711,N_21373,N_21935);
or U22712 (N_22712,N_21578,N_21953);
or U22713 (N_22713,N_21454,N_21580);
nor U22714 (N_22714,N_21537,N_21891);
nand U22715 (N_22715,N_21827,N_21347);
xnor U22716 (N_22716,N_21243,N_21786);
and U22717 (N_22717,N_21003,N_21944);
nor U22718 (N_22718,N_21463,N_21362);
nand U22719 (N_22719,N_21071,N_21309);
and U22720 (N_22720,N_21046,N_21178);
or U22721 (N_22721,N_21275,N_21940);
xnor U22722 (N_22722,N_21780,N_21125);
or U22723 (N_22723,N_21986,N_21509);
and U22724 (N_22724,N_21993,N_21420);
and U22725 (N_22725,N_21907,N_21715);
xor U22726 (N_22726,N_21763,N_21749);
or U22727 (N_22727,N_21713,N_21331);
nand U22728 (N_22728,N_21347,N_21937);
or U22729 (N_22729,N_21616,N_21261);
xor U22730 (N_22730,N_21132,N_21749);
nor U22731 (N_22731,N_21900,N_21020);
or U22732 (N_22732,N_21151,N_21847);
and U22733 (N_22733,N_21907,N_21292);
xor U22734 (N_22734,N_21179,N_21454);
and U22735 (N_22735,N_21348,N_21678);
nor U22736 (N_22736,N_21901,N_21763);
xor U22737 (N_22737,N_21712,N_21412);
nor U22738 (N_22738,N_21245,N_21990);
xnor U22739 (N_22739,N_21414,N_21707);
or U22740 (N_22740,N_21459,N_21770);
nor U22741 (N_22741,N_21886,N_21260);
nand U22742 (N_22742,N_21083,N_21602);
nor U22743 (N_22743,N_21851,N_21460);
or U22744 (N_22744,N_21924,N_21559);
nand U22745 (N_22745,N_21579,N_21342);
and U22746 (N_22746,N_21716,N_21759);
nand U22747 (N_22747,N_21906,N_21266);
xnor U22748 (N_22748,N_21651,N_21645);
and U22749 (N_22749,N_21479,N_21381);
or U22750 (N_22750,N_21366,N_21426);
xnor U22751 (N_22751,N_21637,N_21265);
or U22752 (N_22752,N_21995,N_21825);
xor U22753 (N_22753,N_21100,N_21426);
and U22754 (N_22754,N_21483,N_21059);
or U22755 (N_22755,N_21670,N_21744);
and U22756 (N_22756,N_21005,N_21390);
or U22757 (N_22757,N_21261,N_21255);
nor U22758 (N_22758,N_21661,N_21298);
nand U22759 (N_22759,N_21638,N_21437);
nor U22760 (N_22760,N_21309,N_21278);
nor U22761 (N_22761,N_21493,N_21129);
and U22762 (N_22762,N_21650,N_21040);
nor U22763 (N_22763,N_21463,N_21305);
xor U22764 (N_22764,N_21260,N_21525);
xnor U22765 (N_22765,N_21102,N_21824);
nor U22766 (N_22766,N_21222,N_21723);
and U22767 (N_22767,N_21915,N_21683);
nand U22768 (N_22768,N_21924,N_21577);
nand U22769 (N_22769,N_21077,N_21212);
nand U22770 (N_22770,N_21932,N_21814);
and U22771 (N_22771,N_21334,N_21707);
nor U22772 (N_22772,N_21154,N_21651);
nand U22773 (N_22773,N_21916,N_21704);
and U22774 (N_22774,N_21669,N_21037);
nor U22775 (N_22775,N_21308,N_21938);
xor U22776 (N_22776,N_21196,N_21256);
nand U22777 (N_22777,N_21829,N_21692);
nor U22778 (N_22778,N_21486,N_21127);
xnor U22779 (N_22779,N_21728,N_21021);
and U22780 (N_22780,N_21037,N_21348);
nand U22781 (N_22781,N_21636,N_21791);
or U22782 (N_22782,N_21301,N_21555);
xor U22783 (N_22783,N_21150,N_21633);
xnor U22784 (N_22784,N_21556,N_21469);
and U22785 (N_22785,N_21797,N_21381);
and U22786 (N_22786,N_21803,N_21978);
xor U22787 (N_22787,N_21491,N_21828);
nor U22788 (N_22788,N_21139,N_21459);
xnor U22789 (N_22789,N_21660,N_21693);
or U22790 (N_22790,N_21265,N_21464);
or U22791 (N_22791,N_21645,N_21451);
or U22792 (N_22792,N_21034,N_21703);
xor U22793 (N_22793,N_21582,N_21230);
xnor U22794 (N_22794,N_21998,N_21076);
xnor U22795 (N_22795,N_21124,N_21508);
or U22796 (N_22796,N_21182,N_21659);
nor U22797 (N_22797,N_21880,N_21748);
xnor U22798 (N_22798,N_21164,N_21202);
xor U22799 (N_22799,N_21328,N_21330);
nand U22800 (N_22800,N_21549,N_21471);
and U22801 (N_22801,N_21313,N_21185);
or U22802 (N_22802,N_21605,N_21108);
and U22803 (N_22803,N_21368,N_21383);
and U22804 (N_22804,N_21572,N_21246);
nor U22805 (N_22805,N_21685,N_21507);
or U22806 (N_22806,N_21194,N_21460);
xnor U22807 (N_22807,N_21022,N_21766);
and U22808 (N_22808,N_21531,N_21930);
xnor U22809 (N_22809,N_21592,N_21389);
nor U22810 (N_22810,N_21632,N_21346);
nand U22811 (N_22811,N_21997,N_21207);
and U22812 (N_22812,N_21362,N_21092);
nor U22813 (N_22813,N_21936,N_21085);
and U22814 (N_22814,N_21307,N_21582);
xnor U22815 (N_22815,N_21134,N_21893);
or U22816 (N_22816,N_21333,N_21338);
and U22817 (N_22817,N_21229,N_21967);
xor U22818 (N_22818,N_21113,N_21028);
nand U22819 (N_22819,N_21416,N_21717);
and U22820 (N_22820,N_21302,N_21689);
and U22821 (N_22821,N_21434,N_21734);
xor U22822 (N_22822,N_21607,N_21761);
and U22823 (N_22823,N_21182,N_21290);
nand U22824 (N_22824,N_21820,N_21007);
and U22825 (N_22825,N_21435,N_21094);
and U22826 (N_22826,N_21427,N_21755);
xor U22827 (N_22827,N_21857,N_21290);
xnor U22828 (N_22828,N_21208,N_21754);
or U22829 (N_22829,N_21921,N_21414);
nor U22830 (N_22830,N_21303,N_21775);
nor U22831 (N_22831,N_21966,N_21255);
and U22832 (N_22832,N_21473,N_21981);
nand U22833 (N_22833,N_21473,N_21466);
nand U22834 (N_22834,N_21004,N_21791);
and U22835 (N_22835,N_21692,N_21908);
xnor U22836 (N_22836,N_21844,N_21717);
xor U22837 (N_22837,N_21956,N_21184);
nand U22838 (N_22838,N_21531,N_21475);
nand U22839 (N_22839,N_21046,N_21008);
and U22840 (N_22840,N_21631,N_21325);
nor U22841 (N_22841,N_21490,N_21728);
or U22842 (N_22842,N_21068,N_21962);
or U22843 (N_22843,N_21365,N_21769);
nand U22844 (N_22844,N_21623,N_21226);
and U22845 (N_22845,N_21363,N_21899);
and U22846 (N_22846,N_21504,N_21222);
xnor U22847 (N_22847,N_21685,N_21650);
and U22848 (N_22848,N_21165,N_21654);
nor U22849 (N_22849,N_21487,N_21831);
xnor U22850 (N_22850,N_21232,N_21915);
nand U22851 (N_22851,N_21714,N_21196);
and U22852 (N_22852,N_21704,N_21550);
or U22853 (N_22853,N_21005,N_21887);
or U22854 (N_22854,N_21221,N_21433);
nand U22855 (N_22855,N_21741,N_21254);
or U22856 (N_22856,N_21006,N_21461);
and U22857 (N_22857,N_21277,N_21556);
and U22858 (N_22858,N_21975,N_21468);
nand U22859 (N_22859,N_21632,N_21733);
xnor U22860 (N_22860,N_21654,N_21639);
nand U22861 (N_22861,N_21315,N_21153);
nand U22862 (N_22862,N_21524,N_21401);
and U22863 (N_22863,N_21869,N_21176);
nor U22864 (N_22864,N_21211,N_21970);
or U22865 (N_22865,N_21427,N_21827);
or U22866 (N_22866,N_21187,N_21147);
nor U22867 (N_22867,N_21871,N_21043);
xnor U22868 (N_22868,N_21022,N_21950);
nand U22869 (N_22869,N_21497,N_21404);
or U22870 (N_22870,N_21330,N_21084);
xor U22871 (N_22871,N_21770,N_21358);
nand U22872 (N_22872,N_21369,N_21758);
or U22873 (N_22873,N_21072,N_21490);
or U22874 (N_22874,N_21326,N_21755);
or U22875 (N_22875,N_21115,N_21005);
nor U22876 (N_22876,N_21678,N_21550);
nand U22877 (N_22877,N_21158,N_21199);
nor U22878 (N_22878,N_21367,N_21012);
and U22879 (N_22879,N_21496,N_21060);
or U22880 (N_22880,N_21859,N_21501);
or U22881 (N_22881,N_21065,N_21567);
or U22882 (N_22882,N_21461,N_21775);
or U22883 (N_22883,N_21211,N_21458);
nor U22884 (N_22884,N_21067,N_21599);
nand U22885 (N_22885,N_21278,N_21759);
and U22886 (N_22886,N_21519,N_21967);
xor U22887 (N_22887,N_21454,N_21165);
xnor U22888 (N_22888,N_21379,N_21226);
nand U22889 (N_22889,N_21488,N_21202);
or U22890 (N_22890,N_21444,N_21588);
or U22891 (N_22891,N_21289,N_21024);
and U22892 (N_22892,N_21167,N_21049);
nor U22893 (N_22893,N_21425,N_21931);
and U22894 (N_22894,N_21785,N_21263);
or U22895 (N_22895,N_21370,N_21025);
nand U22896 (N_22896,N_21108,N_21163);
or U22897 (N_22897,N_21754,N_21998);
nand U22898 (N_22898,N_21872,N_21417);
nor U22899 (N_22899,N_21155,N_21545);
and U22900 (N_22900,N_21630,N_21214);
or U22901 (N_22901,N_21713,N_21447);
nand U22902 (N_22902,N_21563,N_21742);
nand U22903 (N_22903,N_21154,N_21099);
xor U22904 (N_22904,N_21499,N_21224);
xor U22905 (N_22905,N_21603,N_21960);
or U22906 (N_22906,N_21790,N_21942);
nand U22907 (N_22907,N_21881,N_21882);
nand U22908 (N_22908,N_21798,N_21997);
and U22909 (N_22909,N_21491,N_21276);
nand U22910 (N_22910,N_21915,N_21025);
or U22911 (N_22911,N_21070,N_21499);
xnor U22912 (N_22912,N_21536,N_21609);
nand U22913 (N_22913,N_21880,N_21103);
and U22914 (N_22914,N_21006,N_21172);
and U22915 (N_22915,N_21541,N_21469);
xor U22916 (N_22916,N_21018,N_21181);
nor U22917 (N_22917,N_21324,N_21410);
xor U22918 (N_22918,N_21805,N_21119);
xnor U22919 (N_22919,N_21855,N_21373);
xor U22920 (N_22920,N_21783,N_21857);
nor U22921 (N_22921,N_21185,N_21293);
and U22922 (N_22922,N_21845,N_21315);
or U22923 (N_22923,N_21153,N_21937);
or U22924 (N_22924,N_21663,N_21069);
and U22925 (N_22925,N_21305,N_21114);
nor U22926 (N_22926,N_21174,N_21707);
xnor U22927 (N_22927,N_21510,N_21908);
xor U22928 (N_22928,N_21087,N_21690);
and U22929 (N_22929,N_21015,N_21532);
xnor U22930 (N_22930,N_21372,N_21075);
nand U22931 (N_22931,N_21530,N_21942);
nor U22932 (N_22932,N_21688,N_21852);
nor U22933 (N_22933,N_21722,N_21779);
or U22934 (N_22934,N_21508,N_21553);
xnor U22935 (N_22935,N_21825,N_21464);
nand U22936 (N_22936,N_21009,N_21023);
nand U22937 (N_22937,N_21994,N_21261);
xor U22938 (N_22938,N_21237,N_21770);
nand U22939 (N_22939,N_21246,N_21479);
xnor U22940 (N_22940,N_21011,N_21601);
nand U22941 (N_22941,N_21854,N_21552);
nand U22942 (N_22942,N_21942,N_21999);
nand U22943 (N_22943,N_21055,N_21283);
xor U22944 (N_22944,N_21261,N_21522);
or U22945 (N_22945,N_21388,N_21039);
nand U22946 (N_22946,N_21168,N_21797);
nand U22947 (N_22947,N_21632,N_21097);
nand U22948 (N_22948,N_21399,N_21922);
nor U22949 (N_22949,N_21488,N_21267);
and U22950 (N_22950,N_21040,N_21607);
xor U22951 (N_22951,N_21000,N_21293);
nor U22952 (N_22952,N_21720,N_21109);
or U22953 (N_22953,N_21111,N_21492);
and U22954 (N_22954,N_21696,N_21175);
nand U22955 (N_22955,N_21689,N_21453);
xor U22956 (N_22956,N_21020,N_21847);
or U22957 (N_22957,N_21993,N_21255);
and U22958 (N_22958,N_21855,N_21996);
nand U22959 (N_22959,N_21012,N_21960);
nor U22960 (N_22960,N_21963,N_21563);
nand U22961 (N_22961,N_21565,N_21227);
nor U22962 (N_22962,N_21500,N_21991);
or U22963 (N_22963,N_21250,N_21354);
or U22964 (N_22964,N_21918,N_21931);
xor U22965 (N_22965,N_21114,N_21693);
nor U22966 (N_22966,N_21827,N_21074);
nand U22967 (N_22967,N_21202,N_21261);
and U22968 (N_22968,N_21965,N_21422);
nor U22969 (N_22969,N_21610,N_21867);
xor U22970 (N_22970,N_21348,N_21240);
xnor U22971 (N_22971,N_21806,N_21003);
nor U22972 (N_22972,N_21427,N_21031);
nand U22973 (N_22973,N_21212,N_21609);
xor U22974 (N_22974,N_21334,N_21808);
xor U22975 (N_22975,N_21314,N_21624);
nor U22976 (N_22976,N_21125,N_21462);
or U22977 (N_22977,N_21959,N_21087);
xor U22978 (N_22978,N_21228,N_21234);
nand U22979 (N_22979,N_21724,N_21911);
xor U22980 (N_22980,N_21374,N_21874);
xnor U22981 (N_22981,N_21081,N_21973);
and U22982 (N_22982,N_21255,N_21283);
xnor U22983 (N_22983,N_21334,N_21783);
nand U22984 (N_22984,N_21471,N_21074);
nand U22985 (N_22985,N_21415,N_21835);
and U22986 (N_22986,N_21892,N_21081);
and U22987 (N_22987,N_21208,N_21450);
nor U22988 (N_22988,N_21470,N_21875);
or U22989 (N_22989,N_21079,N_21412);
and U22990 (N_22990,N_21720,N_21129);
and U22991 (N_22991,N_21098,N_21998);
or U22992 (N_22992,N_21917,N_21363);
nand U22993 (N_22993,N_21270,N_21828);
or U22994 (N_22994,N_21370,N_21127);
nand U22995 (N_22995,N_21749,N_21438);
and U22996 (N_22996,N_21738,N_21448);
and U22997 (N_22997,N_21605,N_21571);
nor U22998 (N_22998,N_21439,N_21788);
nor U22999 (N_22999,N_21305,N_21065);
nand U23000 (N_23000,N_22033,N_22288);
xnor U23001 (N_23001,N_22811,N_22788);
or U23002 (N_23002,N_22947,N_22827);
nor U23003 (N_23003,N_22525,N_22317);
xnor U23004 (N_23004,N_22904,N_22804);
or U23005 (N_23005,N_22863,N_22550);
nor U23006 (N_23006,N_22920,N_22865);
or U23007 (N_23007,N_22361,N_22564);
nor U23008 (N_23008,N_22056,N_22612);
xor U23009 (N_23009,N_22501,N_22994);
nand U23010 (N_23010,N_22896,N_22700);
and U23011 (N_23011,N_22184,N_22977);
xnor U23012 (N_23012,N_22793,N_22653);
xnor U23013 (N_23013,N_22413,N_22208);
xor U23014 (N_23014,N_22967,N_22672);
and U23015 (N_23015,N_22402,N_22576);
or U23016 (N_23016,N_22440,N_22602);
nand U23017 (N_23017,N_22030,N_22284);
or U23018 (N_23018,N_22183,N_22095);
xor U23019 (N_23019,N_22332,N_22328);
nand U23020 (N_23020,N_22324,N_22177);
nor U23021 (N_23021,N_22489,N_22560);
xor U23022 (N_23022,N_22379,N_22728);
and U23023 (N_23023,N_22151,N_22983);
xnor U23024 (N_23024,N_22296,N_22460);
and U23025 (N_23025,N_22817,N_22104);
xnor U23026 (N_23026,N_22866,N_22207);
nand U23027 (N_23027,N_22805,N_22764);
nand U23028 (N_23028,N_22452,N_22676);
xor U23029 (N_23029,N_22267,N_22956);
and U23030 (N_23030,N_22495,N_22506);
and U23031 (N_23031,N_22380,N_22225);
and U23032 (N_23032,N_22523,N_22373);
and U23033 (N_23033,N_22575,N_22893);
nand U23034 (N_23034,N_22099,N_22930);
nor U23035 (N_23035,N_22935,N_22340);
xor U23036 (N_23036,N_22618,N_22200);
or U23037 (N_23037,N_22769,N_22483);
nor U23038 (N_23038,N_22129,N_22914);
xnor U23039 (N_23039,N_22195,N_22339);
or U23040 (N_23040,N_22305,N_22203);
or U23041 (N_23041,N_22012,N_22980);
xor U23042 (N_23042,N_22437,N_22021);
nor U23043 (N_23043,N_22610,N_22916);
xor U23044 (N_23044,N_22997,N_22958);
xor U23045 (N_23045,N_22657,N_22868);
xor U23046 (N_23046,N_22076,N_22051);
nand U23047 (N_23047,N_22392,N_22266);
nor U23048 (N_23048,N_22140,N_22156);
and U23049 (N_23049,N_22924,N_22526);
and U23050 (N_23050,N_22342,N_22420);
and U23051 (N_23051,N_22633,N_22659);
or U23052 (N_23052,N_22219,N_22019);
nor U23053 (N_23053,N_22972,N_22372);
xor U23054 (N_23054,N_22290,N_22889);
and U23055 (N_23055,N_22799,N_22418);
nand U23056 (N_23056,N_22157,N_22120);
or U23057 (N_23057,N_22170,N_22806);
nor U23058 (N_23058,N_22708,N_22790);
nand U23059 (N_23059,N_22243,N_22253);
nor U23060 (N_23060,N_22858,N_22443);
or U23061 (N_23061,N_22285,N_22730);
or U23062 (N_23062,N_22695,N_22687);
nand U23063 (N_23063,N_22415,N_22301);
nand U23064 (N_23064,N_22583,N_22394);
and U23065 (N_23065,N_22240,N_22458);
xnor U23066 (N_23066,N_22666,N_22322);
xnor U23067 (N_23067,N_22250,N_22173);
nor U23068 (N_23068,N_22636,N_22386);
nand U23069 (N_23069,N_22941,N_22142);
or U23070 (N_23070,N_22066,N_22566);
and U23071 (N_23071,N_22106,N_22473);
xor U23072 (N_23072,N_22193,N_22993);
nor U23073 (N_23073,N_22098,N_22595);
and U23074 (N_23074,N_22900,N_22292);
nor U23075 (N_23075,N_22356,N_22204);
and U23076 (N_23076,N_22622,N_22410);
nand U23077 (N_23077,N_22505,N_22289);
xor U23078 (N_23078,N_22234,N_22894);
nand U23079 (N_23079,N_22025,N_22946);
xnor U23080 (N_23080,N_22824,N_22553);
or U23081 (N_23081,N_22009,N_22963);
nand U23082 (N_23082,N_22599,N_22527);
nor U23083 (N_23083,N_22870,N_22760);
or U23084 (N_23084,N_22821,N_22351);
xor U23085 (N_23085,N_22875,N_22513);
nor U23086 (N_23086,N_22918,N_22067);
nand U23087 (N_23087,N_22884,N_22965);
xnor U23088 (N_23088,N_22022,N_22024);
and U23089 (N_23089,N_22381,N_22375);
or U23090 (N_23090,N_22744,N_22973);
xnor U23091 (N_23091,N_22925,N_22346);
and U23092 (N_23092,N_22275,N_22217);
and U23093 (N_23093,N_22913,N_22449);
and U23094 (N_23094,N_22349,N_22154);
xor U23095 (N_23095,N_22403,N_22953);
or U23096 (N_23096,N_22807,N_22548);
and U23097 (N_23097,N_22959,N_22942);
nand U23098 (N_23098,N_22196,N_22368);
and U23099 (N_23099,N_22160,N_22694);
nor U23100 (N_23100,N_22391,N_22216);
or U23101 (N_23101,N_22163,N_22699);
xor U23102 (N_23102,N_22431,N_22629);
nand U23103 (N_23103,N_22014,N_22632);
nand U23104 (N_23104,N_22951,N_22646);
and U23105 (N_23105,N_22678,N_22178);
nor U23106 (N_23106,N_22291,N_22737);
nor U23107 (N_23107,N_22887,N_22181);
xor U23108 (N_23108,N_22830,N_22114);
or U23109 (N_23109,N_22631,N_22003);
nor U23110 (N_23110,N_22626,N_22890);
or U23111 (N_23111,N_22283,N_22544);
and U23112 (N_23112,N_22318,N_22258);
and U23113 (N_23113,N_22222,N_22600);
or U23114 (N_23114,N_22310,N_22681);
xnor U23115 (N_23115,N_22406,N_22774);
nand U23116 (N_23116,N_22046,N_22689);
or U23117 (N_23117,N_22647,N_22319);
xor U23118 (N_23118,N_22693,N_22126);
and U23119 (N_23119,N_22643,N_22090);
nor U23120 (N_23120,N_22214,N_22607);
and U23121 (N_23121,N_22882,N_22143);
nand U23122 (N_23122,N_22069,N_22434);
nand U23123 (N_23123,N_22976,N_22175);
or U23124 (N_23124,N_22574,N_22054);
xnor U23125 (N_23125,N_22109,N_22615);
xnor U23126 (N_23126,N_22209,N_22344);
and U23127 (N_23127,N_22902,N_22795);
or U23128 (N_23128,N_22844,N_22781);
xnor U23129 (N_23129,N_22740,N_22748);
nand U23130 (N_23130,N_22915,N_22869);
and U23131 (N_23131,N_22210,N_22725);
or U23132 (N_23132,N_22899,N_22419);
and U23133 (N_23133,N_22389,N_22171);
or U23134 (N_23134,N_22087,N_22385);
nor U23135 (N_23135,N_22064,N_22702);
and U23136 (N_23136,N_22039,N_22187);
xor U23137 (N_23137,N_22004,N_22573);
and U23138 (N_23138,N_22227,N_22848);
or U23139 (N_23139,N_22684,N_22464);
or U23140 (N_23140,N_22100,N_22966);
or U23141 (N_23141,N_22818,N_22701);
and U23142 (N_23142,N_22759,N_22442);
nor U23143 (N_23143,N_22749,N_22743);
and U23144 (N_23144,N_22042,N_22286);
xor U23145 (N_23145,N_22864,N_22815);
nor U23146 (N_23146,N_22427,N_22911);
xor U23147 (N_23147,N_22282,N_22132);
or U23148 (N_23148,N_22457,N_22704);
xnor U23149 (N_23149,N_22493,N_22975);
nor U23150 (N_23150,N_22934,N_22484);
nor U23151 (N_23151,N_22362,N_22147);
xnor U23152 (N_23152,N_22639,N_22561);
nand U23153 (N_23153,N_22080,N_22088);
nand U23154 (N_23154,N_22119,N_22426);
xor U23155 (N_23155,N_22465,N_22376);
nand U23156 (N_23156,N_22589,N_22241);
nor U23157 (N_23157,N_22948,N_22587);
nor U23158 (N_23158,N_22245,N_22238);
nand U23159 (N_23159,N_22488,N_22127);
nand U23160 (N_23160,N_22136,N_22885);
and U23161 (N_23161,N_22118,N_22813);
nor U23162 (N_23162,N_22360,N_22335);
and U23163 (N_23163,N_22532,N_22365);
or U23164 (N_23164,N_22679,N_22331);
nand U23165 (N_23165,N_22476,N_22783);
nor U23166 (N_23166,N_22761,N_22763);
nand U23167 (N_23167,N_22060,N_22228);
or U23168 (N_23168,N_22537,N_22979);
nor U23169 (N_23169,N_22078,N_22558);
or U23170 (N_23170,N_22623,N_22981);
and U23171 (N_23171,N_22026,N_22037);
nand U23172 (N_23172,N_22919,N_22874);
nand U23173 (N_23173,N_22557,N_22206);
nor U23174 (N_23174,N_22727,N_22881);
nor U23175 (N_23175,N_22131,N_22496);
nor U23176 (N_23176,N_22665,N_22825);
or U23177 (N_23177,N_22441,N_22792);
nor U23178 (N_23178,N_22753,N_22150);
nand U23179 (N_23179,N_22731,N_22279);
or U23180 (N_23180,N_22964,N_22563);
or U23181 (N_23181,N_22668,N_22928);
or U23182 (N_23182,N_22779,N_22358);
xnor U23183 (N_23183,N_22614,N_22117);
and U23184 (N_23184,N_22188,N_22800);
or U23185 (N_23185,N_22252,N_22524);
or U23186 (N_23186,N_22459,N_22316);
and U23187 (N_23187,N_22852,N_22667);
nand U23188 (N_23188,N_22153,N_22438);
and U23189 (N_23189,N_22061,N_22311);
nand U23190 (N_23190,N_22604,N_22498);
nor U23191 (N_23191,N_22303,N_22507);
nand U23192 (N_23192,N_22399,N_22313);
and U23193 (N_23193,N_22338,N_22264);
xor U23194 (N_23194,N_22326,N_22398);
or U23195 (N_23195,N_22627,N_22194);
xor U23196 (N_23196,N_22397,N_22901);
xnor U23197 (N_23197,N_22096,N_22685);
nand U23198 (N_23198,N_22439,N_22097);
xor U23199 (N_23199,N_22363,N_22407);
nand U23200 (N_23200,N_22211,N_22172);
xor U23201 (N_23201,N_22122,N_22485);
or U23202 (N_23202,N_22933,N_22536);
xnor U23203 (N_23203,N_22638,N_22535);
xor U23204 (N_23204,N_22733,N_22735);
or U23205 (N_23205,N_22226,N_22213);
and U23206 (N_23206,N_22487,N_22314);
and U23207 (N_23207,N_22027,N_22932);
or U23208 (N_23208,N_22642,N_22071);
nand U23209 (N_23209,N_22816,N_22005);
nor U23210 (N_23210,N_22931,N_22530);
nor U23211 (N_23211,N_22182,N_22628);
xnor U23212 (N_23212,N_22814,N_22113);
nand U23213 (N_23213,N_22405,N_22220);
nand U23214 (N_23214,N_22533,N_22531);
xor U23215 (N_23215,N_22327,N_22224);
nand U23216 (N_23216,N_22174,N_22218);
and U23217 (N_23217,N_22989,N_22384);
nand U23218 (N_23218,N_22242,N_22886);
nor U23219 (N_23219,N_22011,N_22121);
and U23220 (N_23220,N_22768,N_22509);
nor U23221 (N_23221,N_22709,N_22660);
and U23222 (N_23222,N_22231,N_22084);
nand U23223 (N_23223,N_22717,N_22957);
xor U23224 (N_23224,N_22630,N_22357);
nor U23225 (N_23225,N_22579,N_22149);
or U23226 (N_23226,N_22123,N_22337);
nand U23227 (N_23227,N_22998,N_22256);
xnor U23228 (N_23228,N_22393,N_22594);
xnor U23229 (N_23229,N_22855,N_22169);
xor U23230 (N_23230,N_22680,N_22294);
and U23231 (N_23231,N_22857,N_22738);
or U23232 (N_23232,N_22773,N_22850);
or U23233 (N_23233,N_22081,N_22479);
xor U23234 (N_23234,N_22671,N_22697);
and U23235 (N_23235,N_22649,N_22777);
or U23236 (N_23236,N_22751,N_22837);
xor U23237 (N_23237,N_22370,N_22089);
and U23238 (N_23238,N_22260,N_22674);
nor U23239 (N_23239,N_22762,N_22180);
nand U23240 (N_23240,N_22782,N_22581);
nor U23241 (N_23241,N_22766,N_22995);
nand U23242 (N_23242,N_22378,N_22261);
or U23243 (N_23243,N_22237,N_22045);
or U23244 (N_23244,N_22750,N_22955);
xnor U23245 (N_23245,N_22770,N_22820);
nor U23246 (N_23246,N_22201,N_22785);
or U23247 (N_23247,N_22000,N_22545);
nor U23248 (N_23248,N_22396,N_22107);
and U23249 (N_23249,N_22463,N_22233);
and U23250 (N_23250,N_22836,N_22739);
nor U23251 (N_23251,N_22703,N_22897);
or U23252 (N_23252,N_22306,N_22462);
or U23253 (N_23253,N_22323,N_22036);
nor U23254 (N_23254,N_22984,N_22616);
or U23255 (N_23255,N_22115,N_22822);
and U23256 (N_23256,N_22843,N_22650);
xor U23257 (N_23257,N_22255,N_22705);
and U23258 (N_23258,N_22269,N_22878);
and U23259 (N_23259,N_22974,N_22374);
xor U23260 (N_23260,N_22624,N_22982);
and U23261 (N_23261,N_22845,N_22791);
xor U23262 (N_23262,N_22448,N_22582);
xor U23263 (N_23263,N_22377,N_22569);
xnor U23264 (N_23264,N_22585,N_22521);
xor U23265 (N_23265,N_22189,N_22741);
or U23266 (N_23266,N_22670,N_22721);
or U23267 (N_23267,N_22609,N_22789);
and U23268 (N_23268,N_22608,N_22823);
and U23269 (N_23269,N_22819,N_22613);
and U23270 (N_23270,N_22246,N_22148);
and U23271 (N_23271,N_22390,N_22778);
xnor U23272 (N_23272,N_22943,N_22455);
xnor U23273 (N_23273,N_22508,N_22839);
nor U23274 (N_23274,N_22249,N_22161);
xor U23275 (N_23275,N_22146,N_22929);
nand U23276 (N_23276,N_22765,N_22077);
nor U23277 (N_23277,N_22223,N_22414);
xnor U23278 (N_23278,N_22265,N_22041);
or U23279 (N_23279,N_22645,N_22343);
xor U23280 (N_23280,N_22796,N_22451);
nor U23281 (N_23281,N_22949,N_22565);
or U23282 (N_23282,N_22514,N_22519);
nor U23283 (N_23283,N_22002,N_22141);
xor U23284 (N_23284,N_22517,N_22802);
and U23285 (N_23285,N_22345,N_22467);
xor U23286 (N_23286,N_22571,N_22510);
or U23287 (N_23287,N_22103,N_22101);
nor U23288 (N_23288,N_22747,N_22682);
nor U23289 (N_23289,N_22723,N_22499);
or U23290 (N_23290,N_22347,N_22404);
nor U23291 (N_23291,N_22450,N_22917);
or U23292 (N_23292,N_22539,N_22910);
xor U23293 (N_23293,N_22734,N_22826);
and U23294 (N_23294,N_22176,N_22834);
nand U23295 (N_23295,N_22528,N_22771);
nand U23296 (N_23296,N_22471,N_22350);
or U23297 (N_23297,N_22133,N_22468);
xor U23298 (N_23298,N_22554,N_22675);
nand U23299 (N_23299,N_22683,N_22474);
or U23300 (N_23300,N_22718,N_22031);
xor U23301 (N_23301,N_22883,N_22297);
nand U23302 (N_23302,N_22593,N_22480);
nor U23303 (N_23303,N_22167,N_22546);
nor U23304 (N_23304,N_22722,N_22619);
nor U23305 (N_23305,N_22927,N_22062);
and U23306 (N_23306,N_22754,N_22273);
and U23307 (N_23307,N_22658,N_22477);
xor U23308 (N_23308,N_22590,N_22732);
or U23309 (N_23309,N_22716,N_22656);
and U23310 (N_23310,N_22567,N_22945);
xor U23311 (N_23311,N_22831,N_22726);
xnor U23312 (N_23312,N_22411,N_22634);
nor U23313 (N_23313,N_22274,N_22192);
nand U23314 (N_23314,N_22075,N_22198);
nand U23315 (N_23315,N_22833,N_22862);
nand U23316 (N_23316,N_22259,N_22308);
nand U23317 (N_23317,N_22986,N_22230);
xor U23318 (N_23318,N_22861,N_22348);
nor U23319 (N_23319,N_22110,N_22742);
and U23320 (N_23320,N_22854,N_22416);
xor U23321 (N_23321,N_22293,N_22125);
and U23322 (N_23322,N_22591,N_22707);
xnor U23323 (N_23323,N_22641,N_22159);
nand U23324 (N_23324,N_22417,N_22808);
xnor U23325 (N_23325,N_22073,N_22300);
and U23326 (N_23326,N_22102,N_22637);
nand U23327 (N_23327,N_22355,N_22034);
xnor U23328 (N_23328,N_22454,N_22755);
xor U23329 (N_23329,N_22944,N_22094);
and U23330 (N_23330,N_22272,N_22736);
nor U23331 (N_23331,N_22775,N_22325);
xor U23332 (N_23332,N_22152,N_22877);
nand U23333 (N_23333,N_22185,N_22664);
xor U23334 (N_23334,N_22138,N_22020);
nand U23335 (N_23335,N_22706,N_22715);
or U23336 (N_23336,N_22052,N_22063);
xnor U23337 (N_23337,N_22369,N_22444);
or U23338 (N_23338,N_22661,N_22729);
nor U23339 (N_23339,N_22652,N_22212);
nand U23340 (N_23340,N_22922,N_22654);
xnor U23341 (N_23341,N_22085,N_22516);
or U23342 (N_23342,N_22787,N_22842);
xor U23343 (N_23343,N_22598,N_22570);
nand U23344 (N_23344,N_22239,N_22908);
or U23345 (N_23345,N_22606,N_22853);
nand U23346 (N_23346,N_22466,N_22784);
or U23347 (N_23347,N_22307,N_22926);
and U23348 (N_23348,N_22511,N_22710);
nand U23349 (N_23349,N_22401,N_22801);
nor U23350 (N_23350,N_22746,N_22053);
nor U23351 (N_23351,N_22412,N_22835);
and U23352 (N_23352,N_22662,N_22475);
nor U23353 (N_23353,N_22696,N_22724);
nand U23354 (N_23354,N_22478,N_22597);
and U23355 (N_23355,N_22522,N_22559);
and U23356 (N_23356,N_22540,N_22482);
xor U23357 (N_23357,N_22006,N_22518);
nor U23358 (N_23358,N_22035,N_22542);
or U23359 (N_23359,N_22023,N_22992);
or U23360 (N_23360,N_22058,N_22938);
xor U23361 (N_23361,N_22068,N_22408);
nor U23362 (N_23362,N_22333,N_22280);
xor U23363 (N_23363,N_22111,N_22688);
and U23364 (N_23364,N_22903,N_22798);
nor U23365 (N_23365,N_22860,N_22872);
nor U23366 (N_23366,N_22832,N_22072);
nor U23367 (N_23367,N_22829,N_22047);
nor U23368 (N_23368,N_22436,N_22856);
and U23369 (N_23369,N_22712,N_22898);
nand U23370 (N_23370,N_22555,N_22999);
and U23371 (N_23371,N_22312,N_22341);
nand U23372 (N_23372,N_22572,N_22082);
xor U23373 (N_23373,N_22644,N_22371);
or U23374 (N_23374,N_22888,N_22010);
and U23375 (N_23375,N_22070,N_22758);
and U23376 (N_23376,N_22205,N_22382);
and U23377 (N_23377,N_22083,N_22359);
xnor U23378 (N_23378,N_22329,N_22429);
and U23379 (N_23379,N_22008,N_22655);
and U23380 (N_23380,N_22015,N_22470);
nor U23381 (N_23381,N_22277,N_22032);
xor U23382 (N_23382,N_22491,N_22907);
xnor U23383 (N_23383,N_22446,N_22162);
or U23384 (N_23384,N_22302,N_22968);
or U23385 (N_23385,N_22987,N_22422);
nor U23386 (N_23386,N_22871,N_22481);
nand U23387 (N_23387,N_22295,N_22846);
and U23388 (N_23388,N_22486,N_22445);
or U23389 (N_23389,N_22691,N_22309);
nand U23390 (N_23390,N_22952,N_22909);
or U23391 (N_23391,N_22797,N_22472);
nand U23392 (N_23392,N_22752,N_22937);
xor U23393 (N_23393,N_22625,N_22108);
nor U23394 (N_23394,N_22124,N_22425);
nor U23395 (N_23395,N_22092,N_22601);
nor U23396 (N_23396,N_22503,N_22847);
or U23397 (N_23397,N_22534,N_22859);
and U23398 (N_23398,N_22139,N_22692);
or U23399 (N_23399,N_22936,N_22838);
nor U23400 (N_23400,N_22134,N_22424);
nor U23401 (N_23401,N_22040,N_22892);
xnor U23402 (N_23402,N_22320,N_22669);
nor U23403 (N_23403,N_22512,N_22215);
nand U23404 (N_23404,N_22248,N_22592);
or U23405 (N_23405,N_22043,N_22954);
nand U23406 (N_23406,N_22840,N_22428);
nand U23407 (N_23407,N_22961,N_22996);
nand U23408 (N_23408,N_22018,N_22586);
nor U23409 (N_23409,N_22383,N_22158);
and U23410 (N_23410,N_22016,N_22017);
nand U23411 (N_23411,N_22044,N_22520);
nor U23412 (N_23412,N_22577,N_22812);
or U23413 (N_23413,N_22304,N_22757);
or U23414 (N_23414,N_22809,N_22074);
or U23415 (N_23415,N_22584,N_22130);
and U23416 (N_23416,N_22492,N_22851);
xor U23417 (N_23417,N_22556,N_22876);
nor U23418 (N_23418,N_22112,N_22611);
nand U23419 (N_23419,N_22190,N_22617);
xnor U23420 (N_23420,N_22299,N_22352);
nand U23421 (N_23421,N_22767,N_22271);
and U23422 (N_23422,N_22270,N_22698);
or U23423 (N_23423,N_22780,N_22247);
and U23424 (N_23424,N_22543,N_22409);
nand U23425 (N_23425,N_22596,N_22873);
or U23426 (N_23426,N_22321,N_22315);
nand U23427 (N_23427,N_22199,N_22906);
nand U23428 (N_23428,N_22435,N_22278);
and U23429 (N_23429,N_22251,N_22810);
and U23430 (N_23430,N_22776,N_22235);
nor U23431 (N_23431,N_22867,N_22552);
xnor U23432 (N_23432,N_22686,N_22794);
or U23433 (N_23433,N_22202,N_22690);
or U23434 (N_23434,N_22912,N_22353);
nor U23435 (N_23435,N_22713,N_22461);
nor U23436 (N_23436,N_22990,N_22988);
or U23437 (N_23437,N_22165,N_22456);
nand U23438 (N_23438,N_22116,N_22497);
and U23439 (N_23439,N_22921,N_22529);
nand U23440 (N_23440,N_22950,N_22504);
and U23441 (N_23441,N_22354,N_22786);
nand U23442 (N_23442,N_22547,N_22939);
nand U23443 (N_23443,N_22940,N_22421);
nor U23444 (N_23444,N_22849,N_22186);
nor U23445 (N_23445,N_22756,N_22050);
xor U23446 (N_23446,N_22254,N_22145);
nor U23447 (N_23447,N_22276,N_22879);
and U23448 (N_23448,N_22221,N_22960);
nor U23449 (N_23449,N_22091,N_22978);
xor U23450 (N_23450,N_22962,N_22055);
and U23451 (N_23451,N_22079,N_22364);
nor U23452 (N_23452,N_22330,N_22168);
xnor U23453 (N_23453,N_22494,N_22164);
nand U23454 (N_23454,N_22970,N_22578);
or U23455 (N_23455,N_22433,N_22155);
xor U23456 (N_23456,N_22719,N_22605);
nor U23457 (N_23457,N_22621,N_22257);
xor U23458 (N_23458,N_22387,N_22828);
and U23459 (N_23459,N_22880,N_22191);
and U23460 (N_23460,N_22541,N_22001);
nand U23461 (N_23461,N_22336,N_22395);
nor U23462 (N_23462,N_22086,N_22137);
nand U23463 (N_23463,N_22007,N_22469);
nor U23464 (N_23464,N_22745,N_22551);
nor U23465 (N_23465,N_22603,N_22366);
nor U23466 (N_23466,N_22065,N_22772);
xor U23467 (N_23467,N_22588,N_22244);
nand U23468 (N_23468,N_22490,N_22057);
nor U23469 (N_23469,N_22648,N_22549);
xnor U23470 (N_23470,N_22803,N_22028);
nand U23471 (N_23471,N_22711,N_22515);
xnor U23472 (N_23472,N_22673,N_22502);
nand U23473 (N_23473,N_22423,N_22236);
and U23474 (N_23474,N_22268,N_22640);
xor U23475 (N_23475,N_22197,N_22367);
and U23476 (N_23476,N_22388,N_22049);
or U23477 (N_23477,N_22538,N_22500);
nand U23478 (N_23478,N_22895,N_22232);
nor U23479 (N_23479,N_22059,N_22430);
or U23480 (N_23480,N_22105,N_22562);
nor U23481 (N_23481,N_22038,N_22166);
nand U23482 (N_23482,N_22298,N_22334);
nand U23483 (N_23483,N_22969,N_22144);
and U23484 (N_23484,N_22093,N_22432);
and U23485 (N_23485,N_22923,N_22635);
or U23486 (N_23486,N_22287,N_22013);
nand U23487 (N_23487,N_22400,N_22841);
nor U23488 (N_23488,N_22677,N_22453);
nand U23489 (N_23489,N_22651,N_22229);
or U23490 (N_23490,N_22135,N_22262);
or U23491 (N_23491,N_22048,N_22029);
xnor U23492 (N_23492,N_22263,N_22714);
or U23493 (N_23493,N_22281,N_22128);
and U23494 (N_23494,N_22179,N_22663);
nor U23495 (N_23495,N_22905,N_22891);
nand U23496 (N_23496,N_22985,N_22620);
xor U23497 (N_23497,N_22580,N_22568);
or U23498 (N_23498,N_22991,N_22971);
nand U23499 (N_23499,N_22720,N_22447);
or U23500 (N_23500,N_22050,N_22870);
xor U23501 (N_23501,N_22788,N_22991);
and U23502 (N_23502,N_22143,N_22255);
and U23503 (N_23503,N_22051,N_22976);
or U23504 (N_23504,N_22459,N_22418);
or U23505 (N_23505,N_22446,N_22120);
nand U23506 (N_23506,N_22959,N_22591);
and U23507 (N_23507,N_22681,N_22915);
xor U23508 (N_23508,N_22773,N_22353);
xnor U23509 (N_23509,N_22246,N_22970);
and U23510 (N_23510,N_22884,N_22995);
nor U23511 (N_23511,N_22012,N_22516);
nor U23512 (N_23512,N_22311,N_22436);
and U23513 (N_23513,N_22659,N_22491);
nand U23514 (N_23514,N_22319,N_22036);
nand U23515 (N_23515,N_22273,N_22450);
xnor U23516 (N_23516,N_22019,N_22798);
and U23517 (N_23517,N_22276,N_22383);
nand U23518 (N_23518,N_22334,N_22989);
or U23519 (N_23519,N_22866,N_22117);
nand U23520 (N_23520,N_22083,N_22080);
or U23521 (N_23521,N_22295,N_22428);
or U23522 (N_23522,N_22663,N_22634);
nor U23523 (N_23523,N_22637,N_22665);
xnor U23524 (N_23524,N_22052,N_22248);
nor U23525 (N_23525,N_22549,N_22849);
nand U23526 (N_23526,N_22904,N_22067);
nand U23527 (N_23527,N_22769,N_22758);
or U23528 (N_23528,N_22032,N_22301);
xnor U23529 (N_23529,N_22654,N_22235);
or U23530 (N_23530,N_22724,N_22373);
nand U23531 (N_23531,N_22201,N_22323);
xnor U23532 (N_23532,N_22285,N_22799);
or U23533 (N_23533,N_22835,N_22882);
nand U23534 (N_23534,N_22103,N_22989);
nand U23535 (N_23535,N_22670,N_22848);
xor U23536 (N_23536,N_22020,N_22523);
and U23537 (N_23537,N_22040,N_22870);
or U23538 (N_23538,N_22163,N_22620);
nor U23539 (N_23539,N_22424,N_22234);
xor U23540 (N_23540,N_22362,N_22339);
nand U23541 (N_23541,N_22633,N_22945);
or U23542 (N_23542,N_22436,N_22569);
or U23543 (N_23543,N_22283,N_22869);
nand U23544 (N_23544,N_22642,N_22940);
and U23545 (N_23545,N_22541,N_22460);
xnor U23546 (N_23546,N_22594,N_22652);
xnor U23547 (N_23547,N_22560,N_22125);
and U23548 (N_23548,N_22794,N_22647);
nand U23549 (N_23549,N_22929,N_22952);
nand U23550 (N_23550,N_22679,N_22635);
or U23551 (N_23551,N_22105,N_22440);
or U23552 (N_23552,N_22504,N_22924);
or U23553 (N_23553,N_22070,N_22550);
xor U23554 (N_23554,N_22346,N_22877);
xnor U23555 (N_23555,N_22189,N_22697);
nor U23556 (N_23556,N_22811,N_22552);
nor U23557 (N_23557,N_22197,N_22707);
xor U23558 (N_23558,N_22430,N_22701);
and U23559 (N_23559,N_22659,N_22756);
xnor U23560 (N_23560,N_22463,N_22010);
or U23561 (N_23561,N_22804,N_22077);
or U23562 (N_23562,N_22834,N_22063);
or U23563 (N_23563,N_22039,N_22469);
nor U23564 (N_23564,N_22886,N_22712);
xor U23565 (N_23565,N_22107,N_22170);
nand U23566 (N_23566,N_22943,N_22371);
and U23567 (N_23567,N_22113,N_22841);
or U23568 (N_23568,N_22222,N_22838);
nor U23569 (N_23569,N_22934,N_22000);
and U23570 (N_23570,N_22193,N_22632);
xor U23571 (N_23571,N_22450,N_22275);
xor U23572 (N_23572,N_22216,N_22414);
xor U23573 (N_23573,N_22716,N_22488);
or U23574 (N_23574,N_22666,N_22764);
nor U23575 (N_23575,N_22364,N_22410);
or U23576 (N_23576,N_22574,N_22400);
or U23577 (N_23577,N_22336,N_22685);
nor U23578 (N_23578,N_22969,N_22831);
and U23579 (N_23579,N_22901,N_22584);
xor U23580 (N_23580,N_22339,N_22565);
nor U23581 (N_23581,N_22288,N_22572);
or U23582 (N_23582,N_22217,N_22637);
nor U23583 (N_23583,N_22346,N_22585);
nand U23584 (N_23584,N_22788,N_22783);
nor U23585 (N_23585,N_22030,N_22625);
xor U23586 (N_23586,N_22618,N_22547);
nor U23587 (N_23587,N_22977,N_22877);
nor U23588 (N_23588,N_22990,N_22681);
xor U23589 (N_23589,N_22609,N_22314);
nand U23590 (N_23590,N_22183,N_22343);
or U23591 (N_23591,N_22629,N_22368);
xor U23592 (N_23592,N_22673,N_22821);
xnor U23593 (N_23593,N_22789,N_22524);
and U23594 (N_23594,N_22838,N_22006);
nor U23595 (N_23595,N_22101,N_22011);
or U23596 (N_23596,N_22578,N_22007);
nor U23597 (N_23597,N_22630,N_22482);
nand U23598 (N_23598,N_22961,N_22765);
xor U23599 (N_23599,N_22509,N_22194);
or U23600 (N_23600,N_22690,N_22072);
or U23601 (N_23601,N_22041,N_22395);
and U23602 (N_23602,N_22948,N_22480);
nand U23603 (N_23603,N_22207,N_22598);
nand U23604 (N_23604,N_22680,N_22610);
xnor U23605 (N_23605,N_22242,N_22556);
nand U23606 (N_23606,N_22176,N_22651);
xnor U23607 (N_23607,N_22399,N_22110);
or U23608 (N_23608,N_22143,N_22794);
nand U23609 (N_23609,N_22265,N_22941);
nand U23610 (N_23610,N_22403,N_22249);
nor U23611 (N_23611,N_22697,N_22729);
xnor U23612 (N_23612,N_22401,N_22080);
or U23613 (N_23613,N_22405,N_22410);
or U23614 (N_23614,N_22752,N_22071);
or U23615 (N_23615,N_22411,N_22296);
nand U23616 (N_23616,N_22777,N_22629);
nand U23617 (N_23617,N_22061,N_22607);
nand U23618 (N_23618,N_22153,N_22530);
nor U23619 (N_23619,N_22772,N_22682);
nor U23620 (N_23620,N_22197,N_22452);
nand U23621 (N_23621,N_22575,N_22847);
and U23622 (N_23622,N_22340,N_22567);
nor U23623 (N_23623,N_22688,N_22619);
xnor U23624 (N_23624,N_22979,N_22834);
xnor U23625 (N_23625,N_22709,N_22566);
and U23626 (N_23626,N_22708,N_22662);
or U23627 (N_23627,N_22957,N_22687);
nor U23628 (N_23628,N_22785,N_22516);
or U23629 (N_23629,N_22046,N_22605);
nand U23630 (N_23630,N_22544,N_22570);
and U23631 (N_23631,N_22430,N_22739);
xnor U23632 (N_23632,N_22350,N_22283);
or U23633 (N_23633,N_22313,N_22661);
nor U23634 (N_23634,N_22687,N_22211);
nand U23635 (N_23635,N_22125,N_22495);
nand U23636 (N_23636,N_22243,N_22329);
nand U23637 (N_23637,N_22365,N_22553);
nor U23638 (N_23638,N_22276,N_22852);
xor U23639 (N_23639,N_22708,N_22563);
and U23640 (N_23640,N_22733,N_22197);
nand U23641 (N_23641,N_22888,N_22803);
xor U23642 (N_23642,N_22045,N_22876);
and U23643 (N_23643,N_22626,N_22759);
and U23644 (N_23644,N_22362,N_22497);
and U23645 (N_23645,N_22638,N_22272);
nand U23646 (N_23646,N_22470,N_22884);
nand U23647 (N_23647,N_22993,N_22325);
nor U23648 (N_23648,N_22990,N_22941);
nand U23649 (N_23649,N_22668,N_22247);
nor U23650 (N_23650,N_22854,N_22400);
xnor U23651 (N_23651,N_22972,N_22279);
and U23652 (N_23652,N_22321,N_22394);
or U23653 (N_23653,N_22515,N_22748);
and U23654 (N_23654,N_22098,N_22113);
or U23655 (N_23655,N_22523,N_22475);
nor U23656 (N_23656,N_22563,N_22833);
nor U23657 (N_23657,N_22654,N_22229);
or U23658 (N_23658,N_22075,N_22616);
nand U23659 (N_23659,N_22885,N_22150);
and U23660 (N_23660,N_22730,N_22457);
nand U23661 (N_23661,N_22596,N_22243);
or U23662 (N_23662,N_22464,N_22731);
and U23663 (N_23663,N_22932,N_22976);
xor U23664 (N_23664,N_22812,N_22571);
xnor U23665 (N_23665,N_22415,N_22565);
xnor U23666 (N_23666,N_22655,N_22115);
nor U23667 (N_23667,N_22435,N_22649);
and U23668 (N_23668,N_22957,N_22947);
nor U23669 (N_23669,N_22270,N_22854);
xor U23670 (N_23670,N_22595,N_22134);
and U23671 (N_23671,N_22988,N_22914);
nor U23672 (N_23672,N_22975,N_22264);
or U23673 (N_23673,N_22757,N_22744);
xnor U23674 (N_23674,N_22883,N_22619);
nand U23675 (N_23675,N_22287,N_22788);
xnor U23676 (N_23676,N_22794,N_22290);
nor U23677 (N_23677,N_22848,N_22190);
xnor U23678 (N_23678,N_22605,N_22256);
nand U23679 (N_23679,N_22456,N_22974);
or U23680 (N_23680,N_22553,N_22772);
and U23681 (N_23681,N_22044,N_22923);
or U23682 (N_23682,N_22772,N_22365);
nand U23683 (N_23683,N_22956,N_22349);
and U23684 (N_23684,N_22952,N_22856);
xnor U23685 (N_23685,N_22438,N_22525);
nor U23686 (N_23686,N_22744,N_22770);
or U23687 (N_23687,N_22097,N_22565);
xnor U23688 (N_23688,N_22200,N_22837);
nand U23689 (N_23689,N_22912,N_22770);
and U23690 (N_23690,N_22703,N_22872);
nand U23691 (N_23691,N_22110,N_22509);
xnor U23692 (N_23692,N_22127,N_22280);
nor U23693 (N_23693,N_22868,N_22924);
or U23694 (N_23694,N_22640,N_22975);
xnor U23695 (N_23695,N_22406,N_22728);
and U23696 (N_23696,N_22263,N_22153);
or U23697 (N_23697,N_22325,N_22987);
or U23698 (N_23698,N_22710,N_22384);
xnor U23699 (N_23699,N_22165,N_22560);
xnor U23700 (N_23700,N_22825,N_22113);
nand U23701 (N_23701,N_22858,N_22405);
nand U23702 (N_23702,N_22524,N_22394);
and U23703 (N_23703,N_22555,N_22788);
and U23704 (N_23704,N_22363,N_22725);
xor U23705 (N_23705,N_22538,N_22100);
xor U23706 (N_23706,N_22711,N_22033);
and U23707 (N_23707,N_22279,N_22573);
xnor U23708 (N_23708,N_22101,N_22609);
or U23709 (N_23709,N_22204,N_22577);
nor U23710 (N_23710,N_22934,N_22632);
or U23711 (N_23711,N_22368,N_22425);
xnor U23712 (N_23712,N_22501,N_22256);
nand U23713 (N_23713,N_22320,N_22312);
xnor U23714 (N_23714,N_22071,N_22366);
nor U23715 (N_23715,N_22230,N_22846);
and U23716 (N_23716,N_22154,N_22514);
nor U23717 (N_23717,N_22870,N_22125);
or U23718 (N_23718,N_22789,N_22545);
or U23719 (N_23719,N_22162,N_22445);
or U23720 (N_23720,N_22354,N_22091);
xor U23721 (N_23721,N_22447,N_22396);
or U23722 (N_23722,N_22664,N_22525);
xor U23723 (N_23723,N_22736,N_22152);
xor U23724 (N_23724,N_22623,N_22809);
nand U23725 (N_23725,N_22621,N_22805);
or U23726 (N_23726,N_22382,N_22841);
nor U23727 (N_23727,N_22833,N_22965);
nand U23728 (N_23728,N_22340,N_22791);
or U23729 (N_23729,N_22068,N_22432);
nand U23730 (N_23730,N_22886,N_22362);
nand U23731 (N_23731,N_22963,N_22880);
or U23732 (N_23732,N_22130,N_22407);
nor U23733 (N_23733,N_22590,N_22114);
nor U23734 (N_23734,N_22606,N_22533);
xnor U23735 (N_23735,N_22028,N_22378);
or U23736 (N_23736,N_22648,N_22058);
or U23737 (N_23737,N_22644,N_22267);
or U23738 (N_23738,N_22793,N_22316);
or U23739 (N_23739,N_22548,N_22808);
and U23740 (N_23740,N_22830,N_22567);
nor U23741 (N_23741,N_22306,N_22078);
nor U23742 (N_23742,N_22822,N_22437);
and U23743 (N_23743,N_22974,N_22991);
or U23744 (N_23744,N_22035,N_22426);
xor U23745 (N_23745,N_22214,N_22346);
xor U23746 (N_23746,N_22674,N_22571);
nor U23747 (N_23747,N_22492,N_22954);
and U23748 (N_23748,N_22579,N_22390);
nor U23749 (N_23749,N_22357,N_22807);
or U23750 (N_23750,N_22632,N_22175);
nor U23751 (N_23751,N_22638,N_22603);
or U23752 (N_23752,N_22659,N_22531);
or U23753 (N_23753,N_22683,N_22522);
nand U23754 (N_23754,N_22821,N_22402);
xor U23755 (N_23755,N_22361,N_22260);
nand U23756 (N_23756,N_22261,N_22301);
nor U23757 (N_23757,N_22484,N_22415);
nand U23758 (N_23758,N_22003,N_22115);
or U23759 (N_23759,N_22449,N_22279);
nor U23760 (N_23760,N_22589,N_22075);
nor U23761 (N_23761,N_22920,N_22693);
xor U23762 (N_23762,N_22562,N_22271);
nor U23763 (N_23763,N_22167,N_22478);
nor U23764 (N_23764,N_22400,N_22879);
and U23765 (N_23765,N_22418,N_22023);
nand U23766 (N_23766,N_22673,N_22968);
nand U23767 (N_23767,N_22773,N_22297);
nand U23768 (N_23768,N_22428,N_22231);
xor U23769 (N_23769,N_22481,N_22385);
xor U23770 (N_23770,N_22600,N_22206);
nor U23771 (N_23771,N_22831,N_22389);
and U23772 (N_23772,N_22226,N_22310);
or U23773 (N_23773,N_22302,N_22156);
nor U23774 (N_23774,N_22308,N_22108);
nor U23775 (N_23775,N_22103,N_22147);
nor U23776 (N_23776,N_22502,N_22367);
and U23777 (N_23777,N_22616,N_22047);
and U23778 (N_23778,N_22270,N_22358);
xor U23779 (N_23779,N_22934,N_22252);
nand U23780 (N_23780,N_22394,N_22191);
or U23781 (N_23781,N_22925,N_22420);
nor U23782 (N_23782,N_22880,N_22903);
nand U23783 (N_23783,N_22178,N_22829);
or U23784 (N_23784,N_22409,N_22885);
nand U23785 (N_23785,N_22066,N_22647);
and U23786 (N_23786,N_22981,N_22080);
nor U23787 (N_23787,N_22937,N_22284);
xor U23788 (N_23788,N_22731,N_22065);
or U23789 (N_23789,N_22798,N_22746);
and U23790 (N_23790,N_22863,N_22742);
and U23791 (N_23791,N_22459,N_22789);
and U23792 (N_23792,N_22022,N_22019);
nor U23793 (N_23793,N_22013,N_22926);
xor U23794 (N_23794,N_22887,N_22200);
or U23795 (N_23795,N_22115,N_22430);
nand U23796 (N_23796,N_22436,N_22163);
or U23797 (N_23797,N_22771,N_22288);
or U23798 (N_23798,N_22751,N_22499);
nor U23799 (N_23799,N_22412,N_22625);
nand U23800 (N_23800,N_22596,N_22615);
xnor U23801 (N_23801,N_22705,N_22813);
and U23802 (N_23802,N_22599,N_22400);
nand U23803 (N_23803,N_22431,N_22178);
or U23804 (N_23804,N_22751,N_22867);
and U23805 (N_23805,N_22843,N_22354);
nor U23806 (N_23806,N_22084,N_22365);
and U23807 (N_23807,N_22682,N_22132);
nand U23808 (N_23808,N_22524,N_22458);
nor U23809 (N_23809,N_22487,N_22101);
and U23810 (N_23810,N_22057,N_22477);
and U23811 (N_23811,N_22292,N_22824);
xor U23812 (N_23812,N_22491,N_22209);
and U23813 (N_23813,N_22734,N_22340);
or U23814 (N_23814,N_22288,N_22769);
xor U23815 (N_23815,N_22788,N_22399);
nor U23816 (N_23816,N_22604,N_22741);
nand U23817 (N_23817,N_22908,N_22283);
nand U23818 (N_23818,N_22494,N_22620);
and U23819 (N_23819,N_22208,N_22867);
or U23820 (N_23820,N_22431,N_22666);
nor U23821 (N_23821,N_22787,N_22226);
nand U23822 (N_23822,N_22923,N_22496);
nand U23823 (N_23823,N_22413,N_22738);
xor U23824 (N_23824,N_22668,N_22755);
nand U23825 (N_23825,N_22061,N_22772);
nand U23826 (N_23826,N_22270,N_22021);
and U23827 (N_23827,N_22203,N_22399);
nand U23828 (N_23828,N_22162,N_22609);
xor U23829 (N_23829,N_22472,N_22282);
nand U23830 (N_23830,N_22128,N_22911);
nor U23831 (N_23831,N_22475,N_22988);
nor U23832 (N_23832,N_22590,N_22060);
nand U23833 (N_23833,N_22962,N_22164);
nor U23834 (N_23834,N_22286,N_22058);
nand U23835 (N_23835,N_22880,N_22905);
xnor U23836 (N_23836,N_22664,N_22556);
and U23837 (N_23837,N_22243,N_22496);
or U23838 (N_23838,N_22593,N_22101);
nand U23839 (N_23839,N_22831,N_22115);
and U23840 (N_23840,N_22094,N_22112);
or U23841 (N_23841,N_22408,N_22464);
and U23842 (N_23842,N_22297,N_22775);
xnor U23843 (N_23843,N_22554,N_22269);
xor U23844 (N_23844,N_22721,N_22119);
nand U23845 (N_23845,N_22357,N_22574);
nor U23846 (N_23846,N_22997,N_22928);
xor U23847 (N_23847,N_22115,N_22458);
nand U23848 (N_23848,N_22554,N_22178);
and U23849 (N_23849,N_22818,N_22643);
xor U23850 (N_23850,N_22677,N_22164);
nand U23851 (N_23851,N_22478,N_22733);
and U23852 (N_23852,N_22409,N_22154);
nand U23853 (N_23853,N_22602,N_22899);
nor U23854 (N_23854,N_22100,N_22769);
nor U23855 (N_23855,N_22954,N_22668);
nand U23856 (N_23856,N_22459,N_22417);
xor U23857 (N_23857,N_22020,N_22511);
nor U23858 (N_23858,N_22292,N_22301);
and U23859 (N_23859,N_22962,N_22359);
nand U23860 (N_23860,N_22174,N_22573);
nand U23861 (N_23861,N_22386,N_22810);
nor U23862 (N_23862,N_22270,N_22991);
nor U23863 (N_23863,N_22244,N_22734);
nor U23864 (N_23864,N_22242,N_22830);
nor U23865 (N_23865,N_22694,N_22758);
nor U23866 (N_23866,N_22572,N_22001);
and U23867 (N_23867,N_22539,N_22797);
and U23868 (N_23868,N_22376,N_22073);
nand U23869 (N_23869,N_22380,N_22715);
or U23870 (N_23870,N_22666,N_22845);
xnor U23871 (N_23871,N_22805,N_22553);
or U23872 (N_23872,N_22387,N_22464);
xor U23873 (N_23873,N_22821,N_22670);
nor U23874 (N_23874,N_22945,N_22289);
nor U23875 (N_23875,N_22297,N_22275);
and U23876 (N_23876,N_22386,N_22785);
nor U23877 (N_23877,N_22068,N_22314);
nand U23878 (N_23878,N_22302,N_22834);
or U23879 (N_23879,N_22353,N_22576);
nand U23880 (N_23880,N_22990,N_22580);
xor U23881 (N_23881,N_22008,N_22047);
and U23882 (N_23882,N_22346,N_22115);
nand U23883 (N_23883,N_22654,N_22261);
nor U23884 (N_23884,N_22985,N_22605);
xor U23885 (N_23885,N_22490,N_22118);
or U23886 (N_23886,N_22072,N_22544);
nand U23887 (N_23887,N_22478,N_22045);
and U23888 (N_23888,N_22571,N_22773);
and U23889 (N_23889,N_22246,N_22168);
nor U23890 (N_23890,N_22466,N_22571);
and U23891 (N_23891,N_22904,N_22254);
or U23892 (N_23892,N_22217,N_22644);
nor U23893 (N_23893,N_22132,N_22245);
nand U23894 (N_23894,N_22807,N_22645);
and U23895 (N_23895,N_22951,N_22453);
nor U23896 (N_23896,N_22489,N_22927);
xnor U23897 (N_23897,N_22395,N_22891);
nor U23898 (N_23898,N_22479,N_22549);
nor U23899 (N_23899,N_22918,N_22219);
nand U23900 (N_23900,N_22139,N_22738);
xnor U23901 (N_23901,N_22242,N_22008);
or U23902 (N_23902,N_22362,N_22521);
nand U23903 (N_23903,N_22561,N_22960);
and U23904 (N_23904,N_22776,N_22364);
nand U23905 (N_23905,N_22193,N_22081);
xor U23906 (N_23906,N_22996,N_22340);
xnor U23907 (N_23907,N_22979,N_22815);
nor U23908 (N_23908,N_22072,N_22391);
nor U23909 (N_23909,N_22019,N_22197);
xnor U23910 (N_23910,N_22724,N_22577);
xor U23911 (N_23911,N_22785,N_22404);
xor U23912 (N_23912,N_22532,N_22632);
or U23913 (N_23913,N_22942,N_22170);
and U23914 (N_23914,N_22883,N_22332);
xor U23915 (N_23915,N_22713,N_22568);
xnor U23916 (N_23916,N_22873,N_22085);
nor U23917 (N_23917,N_22988,N_22953);
nand U23918 (N_23918,N_22659,N_22318);
or U23919 (N_23919,N_22953,N_22763);
nand U23920 (N_23920,N_22728,N_22527);
and U23921 (N_23921,N_22263,N_22136);
nor U23922 (N_23922,N_22170,N_22543);
xnor U23923 (N_23923,N_22747,N_22547);
nor U23924 (N_23924,N_22082,N_22520);
nand U23925 (N_23925,N_22982,N_22200);
and U23926 (N_23926,N_22608,N_22840);
nor U23927 (N_23927,N_22800,N_22434);
or U23928 (N_23928,N_22762,N_22536);
and U23929 (N_23929,N_22357,N_22694);
and U23930 (N_23930,N_22806,N_22146);
xnor U23931 (N_23931,N_22458,N_22060);
or U23932 (N_23932,N_22367,N_22442);
nand U23933 (N_23933,N_22486,N_22597);
xor U23934 (N_23934,N_22081,N_22222);
nand U23935 (N_23935,N_22495,N_22727);
nand U23936 (N_23936,N_22148,N_22676);
nand U23937 (N_23937,N_22628,N_22086);
nor U23938 (N_23938,N_22329,N_22279);
nor U23939 (N_23939,N_22742,N_22868);
xnor U23940 (N_23940,N_22412,N_22486);
xor U23941 (N_23941,N_22672,N_22709);
xnor U23942 (N_23942,N_22344,N_22662);
and U23943 (N_23943,N_22232,N_22040);
and U23944 (N_23944,N_22383,N_22975);
or U23945 (N_23945,N_22015,N_22989);
nor U23946 (N_23946,N_22785,N_22686);
or U23947 (N_23947,N_22520,N_22633);
xnor U23948 (N_23948,N_22879,N_22725);
nand U23949 (N_23949,N_22358,N_22176);
or U23950 (N_23950,N_22427,N_22748);
nor U23951 (N_23951,N_22207,N_22877);
and U23952 (N_23952,N_22158,N_22922);
xnor U23953 (N_23953,N_22303,N_22825);
nand U23954 (N_23954,N_22146,N_22382);
and U23955 (N_23955,N_22661,N_22851);
or U23956 (N_23956,N_22875,N_22417);
or U23957 (N_23957,N_22046,N_22816);
xor U23958 (N_23958,N_22782,N_22055);
or U23959 (N_23959,N_22602,N_22210);
nand U23960 (N_23960,N_22023,N_22161);
and U23961 (N_23961,N_22216,N_22453);
nand U23962 (N_23962,N_22856,N_22836);
xor U23963 (N_23963,N_22434,N_22272);
and U23964 (N_23964,N_22066,N_22240);
or U23965 (N_23965,N_22835,N_22109);
nand U23966 (N_23966,N_22616,N_22548);
nand U23967 (N_23967,N_22212,N_22610);
nand U23968 (N_23968,N_22357,N_22504);
nor U23969 (N_23969,N_22576,N_22542);
xor U23970 (N_23970,N_22688,N_22360);
xnor U23971 (N_23971,N_22619,N_22258);
xnor U23972 (N_23972,N_22384,N_22628);
nand U23973 (N_23973,N_22453,N_22329);
nand U23974 (N_23974,N_22670,N_22677);
nand U23975 (N_23975,N_22204,N_22592);
nor U23976 (N_23976,N_22784,N_22660);
and U23977 (N_23977,N_22834,N_22337);
nor U23978 (N_23978,N_22750,N_22488);
xnor U23979 (N_23979,N_22127,N_22337);
and U23980 (N_23980,N_22268,N_22634);
nand U23981 (N_23981,N_22251,N_22901);
and U23982 (N_23982,N_22112,N_22828);
xnor U23983 (N_23983,N_22635,N_22386);
nand U23984 (N_23984,N_22450,N_22676);
xor U23985 (N_23985,N_22356,N_22268);
or U23986 (N_23986,N_22876,N_22383);
nor U23987 (N_23987,N_22252,N_22828);
nor U23988 (N_23988,N_22513,N_22913);
or U23989 (N_23989,N_22729,N_22213);
nor U23990 (N_23990,N_22990,N_22883);
and U23991 (N_23991,N_22749,N_22387);
nand U23992 (N_23992,N_22748,N_22762);
or U23993 (N_23993,N_22017,N_22130);
and U23994 (N_23994,N_22012,N_22434);
nor U23995 (N_23995,N_22157,N_22736);
or U23996 (N_23996,N_22988,N_22372);
xor U23997 (N_23997,N_22552,N_22909);
and U23998 (N_23998,N_22460,N_22437);
or U23999 (N_23999,N_22503,N_22293);
nor U24000 (N_24000,N_23909,N_23249);
xor U24001 (N_24001,N_23683,N_23261);
and U24002 (N_24002,N_23213,N_23963);
nor U24003 (N_24003,N_23485,N_23778);
nor U24004 (N_24004,N_23855,N_23137);
or U24005 (N_24005,N_23423,N_23748);
and U24006 (N_24006,N_23527,N_23230);
nand U24007 (N_24007,N_23179,N_23545);
and U24008 (N_24008,N_23845,N_23952);
or U24009 (N_24009,N_23890,N_23223);
or U24010 (N_24010,N_23838,N_23517);
xor U24011 (N_24011,N_23734,N_23309);
nor U24012 (N_24012,N_23481,N_23823);
xnor U24013 (N_24013,N_23056,N_23035);
nor U24014 (N_24014,N_23062,N_23843);
or U24015 (N_24015,N_23661,N_23727);
or U24016 (N_24016,N_23819,N_23987);
or U24017 (N_24017,N_23132,N_23708);
xnor U24018 (N_24018,N_23717,N_23725);
or U24019 (N_24019,N_23977,N_23453);
nand U24020 (N_24020,N_23447,N_23216);
nand U24021 (N_24021,N_23617,N_23189);
xor U24022 (N_24022,N_23707,N_23271);
or U24023 (N_24023,N_23245,N_23197);
xnor U24024 (N_24024,N_23492,N_23573);
and U24025 (N_24025,N_23943,N_23070);
or U24026 (N_24026,N_23215,N_23495);
and U24027 (N_24027,N_23418,N_23972);
nor U24028 (N_24028,N_23822,N_23983);
xor U24029 (N_24029,N_23883,N_23367);
nor U24030 (N_24030,N_23012,N_23970);
nor U24031 (N_24031,N_23145,N_23746);
and U24032 (N_24032,N_23089,N_23994);
xnor U24033 (N_24033,N_23633,N_23523);
nor U24034 (N_24034,N_23281,N_23072);
and U24035 (N_24035,N_23700,N_23280);
nor U24036 (N_24036,N_23731,N_23858);
or U24037 (N_24037,N_23368,N_23775);
nor U24038 (N_24038,N_23627,N_23552);
and U24039 (N_24039,N_23854,N_23896);
or U24040 (N_24040,N_23759,N_23059);
and U24041 (N_24041,N_23672,N_23766);
nand U24042 (N_24042,N_23018,N_23780);
or U24043 (N_24043,N_23124,N_23566);
nand U24044 (N_24044,N_23160,N_23014);
xor U24045 (N_24045,N_23004,N_23509);
nor U24046 (N_24046,N_23798,N_23642);
nor U24047 (N_24047,N_23944,N_23763);
nor U24048 (N_24048,N_23171,N_23345);
or U24049 (N_24049,N_23872,N_23114);
or U24050 (N_24050,N_23220,N_23113);
or U24051 (N_24051,N_23088,N_23363);
nand U24052 (N_24052,N_23928,N_23126);
and U24053 (N_24053,N_23643,N_23242);
or U24054 (N_24054,N_23602,N_23597);
and U24055 (N_24055,N_23128,N_23592);
and U24056 (N_24056,N_23096,N_23108);
xnor U24057 (N_24057,N_23715,N_23730);
or U24058 (N_24058,N_23741,N_23955);
and U24059 (N_24059,N_23448,N_23739);
or U24060 (N_24060,N_23724,N_23155);
or U24061 (N_24061,N_23637,N_23461);
nor U24062 (N_24062,N_23873,N_23596);
or U24063 (N_24063,N_23678,N_23080);
nand U24064 (N_24064,N_23939,N_23657);
nor U24065 (N_24065,N_23805,N_23282);
nor U24066 (N_24066,N_23359,N_23920);
nor U24067 (N_24067,N_23962,N_23227);
xnor U24068 (N_24068,N_23037,N_23360);
xnor U24069 (N_24069,N_23081,N_23516);
nor U24070 (N_24070,N_23310,N_23737);
or U24071 (N_24071,N_23621,N_23346);
and U24072 (N_24072,N_23269,N_23229);
nor U24073 (N_24073,N_23842,N_23589);
or U24074 (N_24074,N_23050,N_23630);
nand U24075 (N_24075,N_23380,N_23288);
xnor U24076 (N_24076,N_23325,N_23320);
xnor U24077 (N_24077,N_23903,N_23378);
and U24078 (N_24078,N_23090,N_23290);
nand U24079 (N_24079,N_23046,N_23184);
nand U24080 (N_24080,N_23513,N_23567);
and U24081 (N_24081,N_23697,N_23996);
or U24082 (N_24082,N_23499,N_23951);
or U24083 (N_24083,N_23364,N_23802);
nor U24084 (N_24084,N_23752,N_23277);
nor U24085 (N_24085,N_23942,N_23973);
nor U24086 (N_24086,N_23878,N_23777);
and U24087 (N_24087,N_23480,N_23395);
or U24088 (N_24088,N_23714,N_23236);
nor U24089 (N_24089,N_23584,N_23579);
xor U24090 (N_24090,N_23680,N_23486);
nand U24091 (N_24091,N_23922,N_23631);
xnor U24092 (N_24092,N_23040,N_23311);
and U24093 (N_24093,N_23995,N_23696);
nor U24094 (N_24094,N_23097,N_23287);
nor U24095 (N_24095,N_23074,N_23392);
and U24096 (N_24096,N_23001,N_23740);
and U24097 (N_24097,N_23853,N_23474);
xnor U24098 (N_24098,N_23576,N_23235);
or U24099 (N_24099,N_23029,N_23426);
and U24100 (N_24100,N_23259,N_23990);
and U24101 (N_24101,N_23300,N_23723);
or U24102 (N_24102,N_23443,N_23301);
and U24103 (N_24103,N_23340,N_23162);
nor U24104 (N_24104,N_23221,N_23782);
or U24105 (N_24105,N_23403,N_23302);
and U24106 (N_24106,N_23256,N_23025);
nor U24107 (N_24107,N_23837,N_23887);
nand U24108 (N_24108,N_23554,N_23571);
nand U24109 (N_24109,N_23253,N_23626);
and U24110 (N_24110,N_23002,N_23828);
nand U24111 (N_24111,N_23871,N_23634);
xnor U24112 (N_24112,N_23953,N_23515);
xnor U24113 (N_24113,N_23795,N_23112);
or U24114 (N_24114,N_23937,N_23398);
and U24115 (N_24115,N_23479,N_23975);
and U24116 (N_24116,N_23787,N_23670);
xor U24117 (N_24117,N_23514,N_23548);
nor U24118 (N_24118,N_23948,N_23611);
nand U24119 (N_24119,N_23747,N_23488);
nor U24120 (N_24120,N_23275,N_23956);
nor U24121 (N_24121,N_23885,N_23919);
nor U24122 (N_24122,N_23421,N_23228);
xnor U24123 (N_24123,N_23859,N_23652);
nand U24124 (N_24124,N_23231,N_23985);
and U24125 (N_24125,N_23671,N_23976);
xor U24126 (N_24126,N_23568,N_23107);
and U24127 (N_24127,N_23159,N_23744);
nor U24128 (N_24128,N_23565,N_23402);
or U24129 (N_24129,N_23319,N_23255);
xor U24130 (N_24130,N_23237,N_23415);
and U24131 (N_24131,N_23191,N_23372);
or U24132 (N_24132,N_23478,N_23613);
xor U24133 (N_24133,N_23452,N_23457);
nor U24134 (N_24134,N_23459,N_23882);
nor U24135 (N_24135,N_23668,N_23083);
xor U24136 (N_24136,N_23679,N_23243);
nor U24137 (N_24137,N_23122,N_23758);
or U24138 (N_24138,N_23846,N_23390);
nor U24139 (N_24139,N_23620,N_23265);
xor U24140 (N_24140,N_23291,N_23121);
nor U24141 (N_24141,N_23860,N_23503);
and U24142 (N_24142,N_23464,N_23923);
nand U24143 (N_24143,N_23793,N_23535);
or U24144 (N_24144,N_23017,N_23825);
xor U24145 (N_24145,N_23847,N_23988);
nand U24146 (N_24146,N_23590,N_23055);
nor U24147 (N_24147,N_23824,N_23416);
xor U24148 (N_24148,N_23911,N_23247);
nor U24149 (N_24149,N_23966,N_23130);
nand U24150 (N_24150,N_23466,N_23069);
nand U24151 (N_24151,N_23967,N_23019);
or U24152 (N_24152,N_23749,N_23343);
xnor U24153 (N_24153,N_23483,N_23536);
or U24154 (N_24154,N_23907,N_23323);
and U24155 (N_24155,N_23045,N_23157);
or U24156 (N_24156,N_23195,N_23831);
xor U24157 (N_24157,N_23574,N_23789);
or U24158 (N_24158,N_23303,N_23487);
and U24159 (N_24159,N_23519,N_23165);
xor U24160 (N_24160,N_23318,N_23224);
and U24161 (N_24161,N_23347,N_23511);
nor U24162 (N_24162,N_23353,N_23832);
or U24163 (N_24163,N_23469,N_23033);
xor U24164 (N_24164,N_23930,N_23098);
or U24165 (N_24165,N_23940,N_23272);
xor U24166 (N_24166,N_23609,N_23207);
or U24167 (N_24167,N_23028,N_23164);
nor U24168 (N_24168,N_23298,N_23935);
xnor U24169 (N_24169,N_23187,N_23582);
nand U24170 (N_24170,N_23989,N_23826);
nand U24171 (N_24171,N_23404,N_23964);
nor U24172 (N_24172,N_23965,N_23580);
xor U24173 (N_24173,N_23393,N_23530);
and U24174 (N_24174,N_23635,N_23583);
nor U24175 (N_24175,N_23719,N_23034);
and U24176 (N_24176,N_23413,N_23010);
nand U24177 (N_24177,N_23335,N_23677);
and U24178 (N_24178,N_23507,N_23772);
or U24179 (N_24179,N_23933,N_23148);
nand U24180 (N_24180,N_23119,N_23344);
xnor U24181 (N_24181,N_23695,N_23099);
xnor U24182 (N_24182,N_23877,N_23036);
nand U24183 (N_24183,N_23337,N_23118);
nor U24184 (N_24184,N_23640,N_23924);
nand U24185 (N_24185,N_23214,N_23278);
nand U24186 (N_24186,N_23106,N_23833);
nor U24187 (N_24187,N_23208,N_23341);
or U24188 (N_24188,N_23292,N_23039);
and U24189 (N_24189,N_23476,N_23917);
nor U24190 (N_24190,N_23077,N_23910);
nor U24191 (N_24191,N_23125,N_23891);
and U24192 (N_24192,N_23774,N_23501);
nor U24193 (N_24193,N_23295,N_23244);
and U24194 (N_24194,N_23586,N_23958);
xnor U24195 (N_24195,N_23628,N_23827);
nand U24196 (N_24196,N_23103,N_23500);
nor U24197 (N_24197,N_23257,N_23961);
and U24198 (N_24198,N_23960,N_23030);
xnor U24199 (N_24199,N_23424,N_23115);
xor U24200 (N_24200,N_23564,N_23716);
nand U24201 (N_24201,N_23386,N_23803);
nand U24202 (N_24202,N_23437,N_23941);
nor U24203 (N_24203,N_23146,N_23142);
and U24204 (N_24204,N_23477,N_23422);
and U24205 (N_24205,N_23065,N_23232);
and U24206 (N_24206,N_23218,N_23687);
and U24207 (N_24207,N_23117,N_23391);
nand U24208 (N_24208,N_23385,N_23225);
and U24209 (N_24209,N_23894,N_23068);
xnor U24210 (N_24210,N_23949,N_23784);
nand U24211 (N_24211,N_23524,N_23959);
and U24212 (N_24212,N_23296,N_23375);
nand U24213 (N_24213,N_23260,N_23434);
nand U24214 (N_24214,N_23502,N_23086);
nand U24215 (N_24215,N_23026,N_23100);
nand U24216 (N_24216,N_23765,N_23521);
xnor U24217 (N_24217,N_23783,N_23562);
or U24218 (N_24218,N_23166,N_23653);
nor U24219 (N_24219,N_23849,N_23508);
nand U24220 (N_24220,N_23095,N_23427);
nor U24221 (N_24221,N_23102,N_23312);
nand U24222 (N_24222,N_23879,N_23895);
nor U24223 (N_24223,N_23297,N_23123);
xor U24224 (N_24224,N_23092,N_23109);
or U24225 (N_24225,N_23969,N_23745);
nand U24226 (N_24226,N_23176,N_23968);
and U24227 (N_24227,N_23331,N_23264);
nand U24228 (N_24228,N_23556,N_23060);
nand U24229 (N_24229,N_23892,N_23591);
xor U24230 (N_24230,N_23713,N_23632);
xor U24231 (N_24231,N_23594,N_23192);
nand U24232 (N_24232,N_23681,N_23009);
nor U24233 (N_24233,N_23650,N_23250);
or U24234 (N_24234,N_23546,N_23647);
nor U24235 (N_24235,N_23870,N_23711);
nand U24236 (N_24236,N_23052,N_23091);
and U24237 (N_24237,N_23445,N_23755);
nand U24238 (N_24238,N_23601,N_23648);
xnor U24239 (N_24239,N_23575,N_23284);
nor U24240 (N_24240,N_23950,N_23305);
and U24241 (N_24241,N_23581,N_23471);
nor U24242 (N_24242,N_23742,N_23639);
nor U24243 (N_24243,N_23024,N_23354);
or U24244 (N_24244,N_23577,N_23274);
nor U24245 (N_24245,N_23936,N_23429);
nand U24246 (N_24246,N_23701,N_23432);
nor U24247 (N_24247,N_23369,N_23210);
or U24248 (N_24248,N_23902,N_23138);
nor U24249 (N_24249,N_23497,N_23205);
xor U24250 (N_24250,N_23665,N_23254);
or U24251 (N_24251,N_23356,N_23866);
xor U24252 (N_24252,N_23185,N_23408);
and U24253 (N_24253,N_23604,N_23266);
nand U24254 (N_24254,N_23931,N_23954);
or U24255 (N_24255,N_23776,N_23804);
nor U24256 (N_24256,N_23808,N_23921);
and U24257 (N_24257,N_23761,N_23867);
or U24258 (N_24258,N_23414,N_23856);
nand U24259 (N_24259,N_23134,N_23120);
xnor U24260 (N_24260,N_23135,N_23351);
and U24261 (N_24261,N_23893,N_23889);
nor U24262 (N_24262,N_23702,N_23217);
or U24263 (N_24263,N_23233,N_23041);
xor U24264 (N_24264,N_23876,N_23450);
nor U24265 (N_24265,N_23664,N_23797);
xnor U24266 (N_24266,N_23905,N_23992);
nand U24267 (N_24267,N_23182,N_23435);
xnor U24268 (N_24268,N_23504,N_23522);
nand U24269 (N_24269,N_23694,N_23439);
nand U24270 (N_24270,N_23624,N_23087);
xor U24271 (N_24271,N_23079,N_23051);
nor U24272 (N_24272,N_23649,N_23085);
and U24273 (N_24273,N_23490,N_23150);
and U24274 (N_24274,N_23181,N_23561);
or U24275 (N_24275,N_23178,N_23570);
nor U24276 (N_24276,N_23149,N_23689);
or U24277 (N_24277,N_23555,N_23547);
nor U24278 (N_24278,N_23455,N_23201);
and U24279 (N_24279,N_23406,N_23779);
nor U24280 (N_24280,N_23512,N_23463);
nor U24281 (N_24281,N_23934,N_23712);
nor U24282 (N_24282,N_23327,N_23467);
xnor U24283 (N_24283,N_23998,N_23685);
nor U24284 (N_24284,N_23811,N_23836);
xor U24285 (N_24285,N_23927,N_23127);
and U24286 (N_24286,N_23482,N_23686);
xor U24287 (N_24287,N_23984,N_23222);
or U24288 (N_24288,N_23153,N_23465);
xnor U24289 (N_24289,N_23007,N_23350);
and U24290 (N_24290,N_23874,N_23690);
xor U24291 (N_24291,N_23563,N_23316);
and U24292 (N_24292,N_23506,N_23807);
nor U24293 (N_24293,N_23194,N_23991);
or U24294 (N_24294,N_23067,N_23061);
xor U24295 (N_24295,N_23926,N_23349);
or U24296 (N_24296,N_23660,N_23918);
nand U24297 (N_24297,N_23361,N_23021);
nand U24298 (N_24298,N_23286,N_23143);
nor U24299 (N_24299,N_23252,N_23916);
nor U24300 (N_24300,N_23289,N_23412);
or U24301 (N_24301,N_23003,N_23908);
nand U24302 (N_24302,N_23704,N_23334);
xor U24303 (N_24303,N_23865,N_23411);
and U24304 (N_24304,N_23869,N_23559);
xnor U24305 (N_24305,N_23199,N_23321);
or U24306 (N_24306,N_23082,N_23794);
nor U24307 (N_24307,N_23262,N_23757);
nand U24308 (N_24308,N_23673,N_23800);
or U24309 (N_24309,N_23540,N_23382);
nand U24310 (N_24310,N_23336,N_23993);
xnor U24311 (N_24311,N_23806,N_23913);
xnor U24312 (N_24312,N_23440,N_23270);
nand U24313 (N_24313,N_23348,N_23809);
and U24314 (N_24314,N_23206,N_23156);
nand U24315 (N_24315,N_23371,N_23314);
nand U24316 (N_24316,N_23202,N_23644);
xor U24317 (N_24317,N_23615,N_23116);
xor U24318 (N_24318,N_23834,N_23821);
nand U24319 (N_24319,N_23979,N_23684);
nor U24320 (N_24320,N_23528,N_23456);
nand U24321 (N_24321,N_23330,N_23608);
nand U24322 (N_24322,N_23307,N_23888);
xnor U24323 (N_24323,N_23451,N_23267);
xnor U24324 (N_24324,N_23971,N_23365);
or U24325 (N_24325,N_23430,N_23792);
nor U24326 (N_24326,N_23006,N_23815);
xor U24327 (N_24327,N_23449,N_23655);
xnor U24328 (N_24328,N_23785,N_23675);
nor U24329 (N_24329,N_23258,N_23396);
or U24330 (N_24330,N_23158,N_23196);
nand U24331 (N_24331,N_23328,N_23433);
xnor U24332 (N_24332,N_23691,N_23801);
or U24333 (N_24333,N_23394,N_23706);
and U24334 (N_24334,N_23389,N_23729);
xor U24335 (N_24335,N_23728,N_23484);
nor U24336 (N_24336,N_23669,N_23606);
nor U24337 (N_24337,N_23332,N_23193);
or U24338 (N_24338,N_23234,N_23496);
xnor U24339 (N_24339,N_23073,N_23857);
nor U24340 (N_24340,N_23636,N_23897);
nor U24341 (N_24341,N_23428,N_23525);
xnor U24342 (N_24342,N_23549,N_23163);
xor U24343 (N_24343,N_23139,N_23770);
and U24344 (N_24344,N_23538,N_23829);
and U24345 (N_24345,N_23180,N_23063);
nor U24346 (N_24346,N_23442,N_23436);
xor U24347 (N_24347,N_23186,N_23978);
xor U24348 (N_24348,N_23900,N_23110);
and U24349 (N_24349,N_23101,N_23676);
nor U24350 (N_24350,N_23246,N_23498);
nor U24351 (N_24351,N_23384,N_23104);
xor U24352 (N_24352,N_23400,N_23470);
nor U24353 (N_24353,N_23638,N_23796);
nand U24354 (N_24354,N_23339,N_23692);
nor U24355 (N_24355,N_23397,N_23212);
nand U24356 (N_24356,N_23315,N_23454);
nand U24357 (N_24357,N_23674,N_23588);
and U24358 (N_24358,N_23151,N_23355);
or U24359 (N_24359,N_23835,N_23174);
or U24360 (N_24360,N_23446,N_23881);
or U24361 (N_24361,N_23285,N_23659);
and U24362 (N_24362,N_23534,N_23458);
xor U24363 (N_24363,N_23044,N_23557);
nand U24364 (N_24364,N_23377,N_23251);
nor U24365 (N_24365,N_23352,N_23058);
and U24366 (N_24366,N_23000,N_23342);
or U24367 (N_24367,N_23379,N_23722);
xnor U24368 (N_24368,N_23329,N_23767);
nand U24369 (N_24369,N_23263,N_23544);
or U24370 (N_24370,N_23015,N_23699);
or U24371 (N_24371,N_23313,N_23362);
or U24372 (N_24372,N_23338,N_23005);
nor U24373 (N_24373,N_23420,N_23733);
and U24374 (N_24374,N_23764,N_23738);
xnor U24375 (N_24375,N_23317,N_23839);
nor U24376 (N_24376,N_23884,N_23543);
nand U24377 (N_24377,N_23239,N_23152);
and U24378 (N_24378,N_23947,N_23333);
xnor U24379 (N_24379,N_23510,N_23023);
nand U24380 (N_24380,N_23306,N_23374);
or U24381 (N_24381,N_23226,N_23875);
nor U24382 (N_24382,N_23925,N_23013);
nor U24383 (N_24383,N_23868,N_23131);
xor U24384 (N_24384,N_23658,N_23175);
nand U24385 (N_24385,N_23771,N_23726);
or U24386 (N_24386,N_23376,N_23047);
nor U24387 (N_24387,N_23864,N_23852);
or U24388 (N_24388,N_23862,N_23629);
xor U24389 (N_24389,N_23732,N_23425);
xor U24390 (N_24390,N_23814,N_23326);
or U24391 (N_24391,N_23211,N_23473);
nor U24392 (N_24392,N_23760,N_23444);
nand U24393 (N_24393,N_23494,N_23204);
or U24394 (N_24394,N_23472,N_23986);
nand U24395 (N_24395,N_23999,N_23703);
nor U24396 (N_24396,N_23610,N_23539);
xnor U24397 (N_24397,N_23066,N_23324);
xnor U24398 (N_24398,N_23817,N_23753);
xor U24399 (N_24399,N_23754,N_23619);
or U24400 (N_24400,N_23721,N_23786);
nand U24401 (N_24401,N_23788,N_23308);
xor U24402 (N_24402,N_23645,N_23294);
and U24403 (N_24403,N_23848,N_23016);
nor U24404 (N_24404,N_23915,N_23144);
nor U24405 (N_24405,N_23084,N_23736);
xor U24406 (N_24406,N_23593,N_23932);
nor U24407 (N_24407,N_23898,N_23945);
and U24408 (N_24408,N_23491,N_23190);
xor U24409 (N_24409,N_23625,N_23054);
nor U24410 (N_24410,N_23622,N_23541);
nor U24411 (N_24411,N_23840,N_23997);
nor U24412 (N_24412,N_23974,N_23188);
nand U24413 (N_24413,N_23441,N_23399);
and U24414 (N_24414,N_23688,N_23520);
nor U24415 (N_24415,N_23929,N_23791);
and U24416 (N_24416,N_23183,N_23057);
nor U24417 (N_24417,N_23147,N_23946);
and U24418 (N_24418,N_23383,N_23718);
and U24419 (N_24419,N_23769,N_23572);
xnor U24420 (N_24420,N_23078,N_23076);
nor U24421 (N_24421,N_23667,N_23409);
xor U24422 (N_24422,N_23248,N_23167);
or U24423 (N_24423,N_23518,N_23553);
nor U24424 (N_24424,N_23200,N_23273);
and U24425 (N_24425,N_23407,N_23646);
xor U24426 (N_24426,N_23899,N_23008);
and U24427 (N_24427,N_23283,N_23799);
nand U24428 (N_24428,N_23022,N_23111);
or U24429 (N_24429,N_23585,N_23720);
xnor U24430 (N_24430,N_23980,N_23268);
nor U24431 (N_24431,N_23598,N_23462);
or U24432 (N_24432,N_23042,N_23388);
and U24433 (N_24433,N_23818,N_23542);
or U24434 (N_24434,N_23136,N_23735);
nand U24435 (N_24435,N_23914,N_23781);
and U24436 (N_24436,N_23533,N_23529);
xnor U24437 (N_24437,N_23616,N_23168);
nand U24438 (N_24438,N_23612,N_23219);
or U24439 (N_24439,N_23381,N_23299);
and U24440 (N_24440,N_23773,N_23094);
xnor U24441 (N_24441,N_23049,N_23161);
xor U24442 (N_24442,N_23276,N_23032);
xor U24443 (N_24443,N_23129,N_23537);
nand U24444 (N_24444,N_23651,N_23366);
nand U24445 (N_24445,N_23173,N_23603);
nand U24446 (N_24446,N_23607,N_23410);
xor U24447 (N_24447,N_23431,N_23880);
nand U24448 (N_24448,N_23031,N_23662);
or U24449 (N_24449,N_23666,N_23904);
or U24450 (N_24450,N_23209,N_23071);
or U24451 (N_24451,N_23750,N_23768);
nor U24452 (N_24452,N_23020,N_23460);
nor U24453 (N_24453,N_23813,N_23614);
or U24454 (N_24454,N_23475,N_23863);
xor U24455 (N_24455,N_23663,N_23938);
or U24456 (N_24456,N_23240,N_23560);
and U24457 (N_24457,N_23105,N_23532);
and U24458 (N_24458,N_23654,N_23698);
or U24459 (N_24459,N_23912,N_23526);
or U24460 (N_24460,N_23401,N_23605);
and U24461 (N_24461,N_23851,N_23293);
xor U24462 (N_24462,N_23844,N_23322);
nor U24463 (N_24463,N_23850,N_23762);
nor U24464 (N_24464,N_23505,N_23693);
nand U24465 (N_24465,N_23154,N_23438);
or U24466 (N_24466,N_23064,N_23841);
or U24467 (N_24467,N_23558,N_23493);
nand U24468 (N_24468,N_23038,N_23682);
and U24469 (N_24469,N_23756,N_23623);
nor U24470 (N_24470,N_23569,N_23551);
or U24471 (N_24471,N_23981,N_23531);
nand U24472 (N_24472,N_23358,N_23405);
or U24473 (N_24473,N_23790,N_23468);
nand U24474 (N_24474,N_23169,N_23133);
or U24475 (N_24475,N_23304,N_23140);
or U24476 (N_24476,N_23241,N_23820);
or U24477 (N_24477,N_23816,N_23641);
nand U24478 (N_24478,N_23075,N_23906);
or U24479 (N_24479,N_23177,N_23578);
xnor U24480 (N_24480,N_23743,N_23886);
xnor U24481 (N_24481,N_23810,N_23419);
nand U24482 (N_24482,N_23901,N_23861);
nand U24483 (N_24483,N_23587,N_23357);
or U24484 (N_24484,N_23417,N_23618);
or U24485 (N_24485,N_23053,N_23599);
or U24486 (N_24486,N_23595,N_23705);
nand U24487 (N_24487,N_23957,N_23982);
or U24488 (N_24488,N_23812,N_23203);
and U24489 (N_24489,N_23027,N_23093);
nand U24490 (N_24490,N_23600,N_23279);
xor U24491 (N_24491,N_23048,N_23656);
or U24492 (N_24492,N_23830,N_23489);
or U24493 (N_24493,N_23550,N_23172);
and U24494 (N_24494,N_23370,N_23710);
nor U24495 (N_24495,N_23387,N_23709);
and U24496 (N_24496,N_23751,N_23011);
nor U24497 (N_24497,N_23238,N_23170);
and U24498 (N_24498,N_23373,N_23141);
or U24499 (N_24499,N_23043,N_23198);
nand U24500 (N_24500,N_23765,N_23472);
xor U24501 (N_24501,N_23025,N_23716);
and U24502 (N_24502,N_23654,N_23874);
or U24503 (N_24503,N_23776,N_23374);
nor U24504 (N_24504,N_23394,N_23383);
or U24505 (N_24505,N_23922,N_23349);
or U24506 (N_24506,N_23035,N_23571);
or U24507 (N_24507,N_23494,N_23645);
or U24508 (N_24508,N_23362,N_23401);
xor U24509 (N_24509,N_23066,N_23388);
nand U24510 (N_24510,N_23278,N_23717);
or U24511 (N_24511,N_23340,N_23032);
or U24512 (N_24512,N_23578,N_23298);
or U24513 (N_24513,N_23126,N_23160);
or U24514 (N_24514,N_23506,N_23140);
xor U24515 (N_24515,N_23074,N_23619);
and U24516 (N_24516,N_23126,N_23384);
nor U24517 (N_24517,N_23373,N_23907);
xnor U24518 (N_24518,N_23011,N_23754);
or U24519 (N_24519,N_23890,N_23383);
xnor U24520 (N_24520,N_23153,N_23944);
or U24521 (N_24521,N_23722,N_23631);
or U24522 (N_24522,N_23677,N_23030);
or U24523 (N_24523,N_23642,N_23596);
and U24524 (N_24524,N_23384,N_23073);
xor U24525 (N_24525,N_23804,N_23436);
xor U24526 (N_24526,N_23249,N_23600);
or U24527 (N_24527,N_23642,N_23398);
or U24528 (N_24528,N_23930,N_23053);
nand U24529 (N_24529,N_23009,N_23362);
xnor U24530 (N_24530,N_23404,N_23570);
nor U24531 (N_24531,N_23876,N_23343);
and U24532 (N_24532,N_23406,N_23848);
and U24533 (N_24533,N_23481,N_23762);
xnor U24534 (N_24534,N_23817,N_23032);
nor U24535 (N_24535,N_23547,N_23924);
and U24536 (N_24536,N_23358,N_23172);
nand U24537 (N_24537,N_23596,N_23127);
nand U24538 (N_24538,N_23872,N_23165);
nor U24539 (N_24539,N_23665,N_23985);
and U24540 (N_24540,N_23530,N_23382);
xor U24541 (N_24541,N_23469,N_23904);
xnor U24542 (N_24542,N_23395,N_23170);
xor U24543 (N_24543,N_23139,N_23638);
and U24544 (N_24544,N_23822,N_23530);
and U24545 (N_24545,N_23193,N_23127);
nor U24546 (N_24546,N_23267,N_23436);
nand U24547 (N_24547,N_23699,N_23641);
nor U24548 (N_24548,N_23431,N_23480);
nand U24549 (N_24549,N_23083,N_23858);
or U24550 (N_24550,N_23750,N_23266);
nand U24551 (N_24551,N_23183,N_23083);
or U24552 (N_24552,N_23538,N_23465);
xnor U24553 (N_24553,N_23204,N_23261);
nor U24554 (N_24554,N_23229,N_23905);
nor U24555 (N_24555,N_23743,N_23765);
xor U24556 (N_24556,N_23426,N_23101);
xnor U24557 (N_24557,N_23486,N_23785);
xor U24558 (N_24558,N_23045,N_23120);
nor U24559 (N_24559,N_23880,N_23720);
and U24560 (N_24560,N_23652,N_23493);
nor U24561 (N_24561,N_23335,N_23554);
nand U24562 (N_24562,N_23550,N_23367);
nor U24563 (N_24563,N_23924,N_23245);
nor U24564 (N_24564,N_23576,N_23956);
and U24565 (N_24565,N_23040,N_23401);
and U24566 (N_24566,N_23739,N_23737);
and U24567 (N_24567,N_23029,N_23052);
and U24568 (N_24568,N_23136,N_23008);
nor U24569 (N_24569,N_23188,N_23443);
xnor U24570 (N_24570,N_23130,N_23937);
or U24571 (N_24571,N_23643,N_23862);
nor U24572 (N_24572,N_23363,N_23051);
nor U24573 (N_24573,N_23158,N_23663);
and U24574 (N_24574,N_23095,N_23028);
or U24575 (N_24575,N_23752,N_23327);
nor U24576 (N_24576,N_23424,N_23178);
or U24577 (N_24577,N_23373,N_23464);
xnor U24578 (N_24578,N_23842,N_23232);
nand U24579 (N_24579,N_23723,N_23342);
and U24580 (N_24580,N_23376,N_23914);
and U24581 (N_24581,N_23262,N_23390);
xor U24582 (N_24582,N_23329,N_23326);
or U24583 (N_24583,N_23421,N_23042);
xor U24584 (N_24584,N_23561,N_23096);
or U24585 (N_24585,N_23721,N_23900);
and U24586 (N_24586,N_23509,N_23221);
xor U24587 (N_24587,N_23321,N_23758);
and U24588 (N_24588,N_23433,N_23202);
xor U24589 (N_24589,N_23343,N_23566);
xnor U24590 (N_24590,N_23449,N_23379);
or U24591 (N_24591,N_23177,N_23269);
or U24592 (N_24592,N_23041,N_23875);
nor U24593 (N_24593,N_23429,N_23251);
nand U24594 (N_24594,N_23214,N_23235);
nor U24595 (N_24595,N_23304,N_23883);
xnor U24596 (N_24596,N_23128,N_23340);
nand U24597 (N_24597,N_23566,N_23116);
nor U24598 (N_24598,N_23821,N_23640);
xnor U24599 (N_24599,N_23391,N_23609);
or U24600 (N_24600,N_23975,N_23016);
nand U24601 (N_24601,N_23450,N_23227);
or U24602 (N_24602,N_23910,N_23471);
nor U24603 (N_24603,N_23461,N_23296);
nor U24604 (N_24604,N_23527,N_23500);
nand U24605 (N_24605,N_23066,N_23004);
and U24606 (N_24606,N_23730,N_23613);
nor U24607 (N_24607,N_23748,N_23207);
nor U24608 (N_24608,N_23486,N_23621);
nand U24609 (N_24609,N_23419,N_23245);
xor U24610 (N_24610,N_23066,N_23106);
or U24611 (N_24611,N_23278,N_23586);
nand U24612 (N_24612,N_23943,N_23970);
nor U24613 (N_24613,N_23817,N_23800);
or U24614 (N_24614,N_23464,N_23942);
or U24615 (N_24615,N_23046,N_23961);
and U24616 (N_24616,N_23794,N_23547);
or U24617 (N_24617,N_23364,N_23563);
nor U24618 (N_24618,N_23653,N_23508);
xor U24619 (N_24619,N_23880,N_23153);
and U24620 (N_24620,N_23196,N_23803);
xor U24621 (N_24621,N_23163,N_23045);
or U24622 (N_24622,N_23565,N_23789);
or U24623 (N_24623,N_23144,N_23271);
nand U24624 (N_24624,N_23787,N_23115);
xnor U24625 (N_24625,N_23278,N_23484);
nand U24626 (N_24626,N_23680,N_23242);
xor U24627 (N_24627,N_23148,N_23562);
nor U24628 (N_24628,N_23132,N_23287);
nor U24629 (N_24629,N_23920,N_23795);
nand U24630 (N_24630,N_23704,N_23143);
xor U24631 (N_24631,N_23679,N_23514);
xnor U24632 (N_24632,N_23536,N_23724);
nand U24633 (N_24633,N_23671,N_23943);
nand U24634 (N_24634,N_23905,N_23125);
and U24635 (N_24635,N_23034,N_23411);
nand U24636 (N_24636,N_23730,N_23065);
nand U24637 (N_24637,N_23762,N_23694);
nand U24638 (N_24638,N_23580,N_23168);
nand U24639 (N_24639,N_23542,N_23665);
nand U24640 (N_24640,N_23436,N_23300);
nand U24641 (N_24641,N_23543,N_23079);
and U24642 (N_24642,N_23702,N_23113);
and U24643 (N_24643,N_23994,N_23256);
nor U24644 (N_24644,N_23065,N_23912);
nor U24645 (N_24645,N_23937,N_23109);
nor U24646 (N_24646,N_23400,N_23999);
and U24647 (N_24647,N_23812,N_23246);
nor U24648 (N_24648,N_23894,N_23216);
nand U24649 (N_24649,N_23362,N_23549);
or U24650 (N_24650,N_23737,N_23593);
nand U24651 (N_24651,N_23320,N_23201);
or U24652 (N_24652,N_23335,N_23516);
and U24653 (N_24653,N_23583,N_23924);
nor U24654 (N_24654,N_23220,N_23165);
and U24655 (N_24655,N_23007,N_23069);
xnor U24656 (N_24656,N_23834,N_23884);
nor U24657 (N_24657,N_23399,N_23222);
xnor U24658 (N_24658,N_23557,N_23188);
or U24659 (N_24659,N_23046,N_23040);
nor U24660 (N_24660,N_23926,N_23627);
nor U24661 (N_24661,N_23994,N_23107);
nand U24662 (N_24662,N_23764,N_23702);
xor U24663 (N_24663,N_23320,N_23826);
nor U24664 (N_24664,N_23532,N_23934);
or U24665 (N_24665,N_23475,N_23563);
or U24666 (N_24666,N_23090,N_23402);
or U24667 (N_24667,N_23462,N_23834);
xor U24668 (N_24668,N_23950,N_23030);
or U24669 (N_24669,N_23848,N_23543);
xnor U24670 (N_24670,N_23543,N_23164);
xnor U24671 (N_24671,N_23256,N_23524);
xor U24672 (N_24672,N_23759,N_23162);
nor U24673 (N_24673,N_23811,N_23525);
nand U24674 (N_24674,N_23090,N_23188);
xnor U24675 (N_24675,N_23096,N_23675);
xnor U24676 (N_24676,N_23139,N_23548);
and U24677 (N_24677,N_23777,N_23814);
nor U24678 (N_24678,N_23407,N_23978);
or U24679 (N_24679,N_23972,N_23813);
nand U24680 (N_24680,N_23961,N_23579);
nand U24681 (N_24681,N_23608,N_23398);
or U24682 (N_24682,N_23497,N_23245);
nand U24683 (N_24683,N_23472,N_23846);
or U24684 (N_24684,N_23584,N_23697);
and U24685 (N_24685,N_23213,N_23404);
and U24686 (N_24686,N_23890,N_23423);
nor U24687 (N_24687,N_23383,N_23354);
or U24688 (N_24688,N_23217,N_23900);
nor U24689 (N_24689,N_23324,N_23620);
xnor U24690 (N_24690,N_23899,N_23887);
nand U24691 (N_24691,N_23521,N_23877);
xnor U24692 (N_24692,N_23852,N_23978);
and U24693 (N_24693,N_23875,N_23869);
nand U24694 (N_24694,N_23759,N_23150);
and U24695 (N_24695,N_23363,N_23156);
nor U24696 (N_24696,N_23272,N_23664);
nand U24697 (N_24697,N_23016,N_23824);
nand U24698 (N_24698,N_23436,N_23454);
nor U24699 (N_24699,N_23913,N_23186);
nand U24700 (N_24700,N_23014,N_23423);
or U24701 (N_24701,N_23707,N_23527);
or U24702 (N_24702,N_23592,N_23269);
nor U24703 (N_24703,N_23826,N_23215);
xnor U24704 (N_24704,N_23642,N_23534);
or U24705 (N_24705,N_23165,N_23617);
and U24706 (N_24706,N_23450,N_23985);
xnor U24707 (N_24707,N_23138,N_23497);
xor U24708 (N_24708,N_23627,N_23867);
xnor U24709 (N_24709,N_23285,N_23601);
nor U24710 (N_24710,N_23664,N_23178);
nor U24711 (N_24711,N_23522,N_23521);
or U24712 (N_24712,N_23668,N_23525);
and U24713 (N_24713,N_23155,N_23248);
and U24714 (N_24714,N_23928,N_23247);
or U24715 (N_24715,N_23822,N_23922);
or U24716 (N_24716,N_23446,N_23722);
nand U24717 (N_24717,N_23202,N_23063);
xor U24718 (N_24718,N_23873,N_23066);
nor U24719 (N_24719,N_23348,N_23777);
or U24720 (N_24720,N_23751,N_23962);
nor U24721 (N_24721,N_23001,N_23031);
and U24722 (N_24722,N_23060,N_23631);
or U24723 (N_24723,N_23626,N_23766);
and U24724 (N_24724,N_23588,N_23289);
xnor U24725 (N_24725,N_23264,N_23608);
nor U24726 (N_24726,N_23465,N_23531);
xor U24727 (N_24727,N_23972,N_23655);
and U24728 (N_24728,N_23211,N_23284);
nor U24729 (N_24729,N_23086,N_23220);
nand U24730 (N_24730,N_23568,N_23691);
nand U24731 (N_24731,N_23628,N_23363);
nand U24732 (N_24732,N_23497,N_23687);
or U24733 (N_24733,N_23710,N_23417);
xor U24734 (N_24734,N_23496,N_23043);
xnor U24735 (N_24735,N_23729,N_23252);
or U24736 (N_24736,N_23037,N_23934);
and U24737 (N_24737,N_23608,N_23412);
or U24738 (N_24738,N_23871,N_23331);
xnor U24739 (N_24739,N_23857,N_23449);
nor U24740 (N_24740,N_23074,N_23372);
or U24741 (N_24741,N_23713,N_23483);
nand U24742 (N_24742,N_23926,N_23550);
xnor U24743 (N_24743,N_23623,N_23195);
nand U24744 (N_24744,N_23229,N_23416);
or U24745 (N_24745,N_23196,N_23779);
xor U24746 (N_24746,N_23991,N_23369);
and U24747 (N_24747,N_23084,N_23398);
nor U24748 (N_24748,N_23258,N_23420);
and U24749 (N_24749,N_23210,N_23543);
nor U24750 (N_24750,N_23599,N_23479);
nor U24751 (N_24751,N_23782,N_23557);
nand U24752 (N_24752,N_23336,N_23362);
xor U24753 (N_24753,N_23288,N_23539);
and U24754 (N_24754,N_23595,N_23151);
xnor U24755 (N_24755,N_23074,N_23019);
xnor U24756 (N_24756,N_23207,N_23636);
nor U24757 (N_24757,N_23891,N_23399);
or U24758 (N_24758,N_23508,N_23570);
xor U24759 (N_24759,N_23104,N_23693);
xnor U24760 (N_24760,N_23489,N_23292);
nand U24761 (N_24761,N_23828,N_23696);
nand U24762 (N_24762,N_23699,N_23069);
nor U24763 (N_24763,N_23602,N_23835);
xnor U24764 (N_24764,N_23078,N_23798);
nor U24765 (N_24765,N_23712,N_23011);
xor U24766 (N_24766,N_23977,N_23959);
or U24767 (N_24767,N_23983,N_23750);
xnor U24768 (N_24768,N_23143,N_23457);
and U24769 (N_24769,N_23481,N_23160);
xor U24770 (N_24770,N_23292,N_23383);
and U24771 (N_24771,N_23800,N_23017);
and U24772 (N_24772,N_23659,N_23456);
or U24773 (N_24773,N_23503,N_23705);
nand U24774 (N_24774,N_23471,N_23338);
or U24775 (N_24775,N_23718,N_23106);
nand U24776 (N_24776,N_23992,N_23224);
nand U24777 (N_24777,N_23999,N_23129);
nand U24778 (N_24778,N_23231,N_23312);
or U24779 (N_24779,N_23109,N_23380);
nor U24780 (N_24780,N_23803,N_23792);
or U24781 (N_24781,N_23637,N_23373);
xnor U24782 (N_24782,N_23241,N_23739);
or U24783 (N_24783,N_23378,N_23383);
and U24784 (N_24784,N_23822,N_23605);
and U24785 (N_24785,N_23388,N_23393);
xor U24786 (N_24786,N_23637,N_23869);
or U24787 (N_24787,N_23082,N_23689);
nand U24788 (N_24788,N_23448,N_23329);
xnor U24789 (N_24789,N_23992,N_23711);
nand U24790 (N_24790,N_23558,N_23625);
and U24791 (N_24791,N_23359,N_23079);
and U24792 (N_24792,N_23277,N_23408);
nand U24793 (N_24793,N_23196,N_23519);
nand U24794 (N_24794,N_23878,N_23983);
nand U24795 (N_24795,N_23433,N_23677);
nor U24796 (N_24796,N_23503,N_23373);
nor U24797 (N_24797,N_23837,N_23311);
nand U24798 (N_24798,N_23646,N_23309);
nand U24799 (N_24799,N_23468,N_23037);
nand U24800 (N_24800,N_23421,N_23145);
or U24801 (N_24801,N_23608,N_23745);
nor U24802 (N_24802,N_23958,N_23566);
nand U24803 (N_24803,N_23805,N_23978);
or U24804 (N_24804,N_23016,N_23887);
or U24805 (N_24805,N_23515,N_23016);
and U24806 (N_24806,N_23969,N_23512);
or U24807 (N_24807,N_23102,N_23101);
and U24808 (N_24808,N_23840,N_23266);
xor U24809 (N_24809,N_23620,N_23624);
nor U24810 (N_24810,N_23933,N_23691);
nand U24811 (N_24811,N_23980,N_23400);
nand U24812 (N_24812,N_23821,N_23266);
or U24813 (N_24813,N_23429,N_23784);
nor U24814 (N_24814,N_23034,N_23683);
nand U24815 (N_24815,N_23070,N_23256);
nor U24816 (N_24816,N_23450,N_23987);
or U24817 (N_24817,N_23147,N_23108);
nand U24818 (N_24818,N_23057,N_23127);
xnor U24819 (N_24819,N_23111,N_23915);
nand U24820 (N_24820,N_23067,N_23807);
and U24821 (N_24821,N_23551,N_23031);
nand U24822 (N_24822,N_23335,N_23888);
xor U24823 (N_24823,N_23719,N_23441);
nor U24824 (N_24824,N_23263,N_23445);
and U24825 (N_24825,N_23151,N_23423);
or U24826 (N_24826,N_23937,N_23318);
xnor U24827 (N_24827,N_23401,N_23608);
nand U24828 (N_24828,N_23417,N_23040);
or U24829 (N_24829,N_23280,N_23826);
nand U24830 (N_24830,N_23371,N_23743);
nor U24831 (N_24831,N_23193,N_23620);
nand U24832 (N_24832,N_23576,N_23899);
or U24833 (N_24833,N_23112,N_23492);
nand U24834 (N_24834,N_23053,N_23610);
xnor U24835 (N_24835,N_23701,N_23256);
xnor U24836 (N_24836,N_23364,N_23755);
and U24837 (N_24837,N_23544,N_23839);
nor U24838 (N_24838,N_23160,N_23188);
and U24839 (N_24839,N_23978,N_23329);
and U24840 (N_24840,N_23422,N_23661);
or U24841 (N_24841,N_23353,N_23144);
and U24842 (N_24842,N_23494,N_23471);
xnor U24843 (N_24843,N_23192,N_23576);
or U24844 (N_24844,N_23454,N_23919);
xnor U24845 (N_24845,N_23222,N_23675);
nor U24846 (N_24846,N_23867,N_23065);
or U24847 (N_24847,N_23501,N_23406);
or U24848 (N_24848,N_23537,N_23362);
or U24849 (N_24849,N_23061,N_23249);
nand U24850 (N_24850,N_23259,N_23318);
or U24851 (N_24851,N_23519,N_23300);
nor U24852 (N_24852,N_23056,N_23795);
or U24853 (N_24853,N_23719,N_23049);
nand U24854 (N_24854,N_23261,N_23338);
xor U24855 (N_24855,N_23044,N_23324);
or U24856 (N_24856,N_23016,N_23693);
or U24857 (N_24857,N_23208,N_23014);
nand U24858 (N_24858,N_23350,N_23289);
and U24859 (N_24859,N_23909,N_23040);
or U24860 (N_24860,N_23733,N_23038);
nand U24861 (N_24861,N_23672,N_23784);
and U24862 (N_24862,N_23915,N_23492);
or U24863 (N_24863,N_23705,N_23650);
xnor U24864 (N_24864,N_23293,N_23057);
nor U24865 (N_24865,N_23376,N_23125);
nor U24866 (N_24866,N_23526,N_23646);
nand U24867 (N_24867,N_23694,N_23279);
or U24868 (N_24868,N_23605,N_23705);
or U24869 (N_24869,N_23997,N_23417);
or U24870 (N_24870,N_23129,N_23481);
and U24871 (N_24871,N_23633,N_23787);
and U24872 (N_24872,N_23097,N_23009);
xnor U24873 (N_24873,N_23248,N_23731);
or U24874 (N_24874,N_23273,N_23586);
xor U24875 (N_24875,N_23915,N_23531);
or U24876 (N_24876,N_23508,N_23483);
or U24877 (N_24877,N_23306,N_23201);
nor U24878 (N_24878,N_23443,N_23487);
nand U24879 (N_24879,N_23336,N_23119);
and U24880 (N_24880,N_23591,N_23874);
nor U24881 (N_24881,N_23588,N_23074);
or U24882 (N_24882,N_23824,N_23604);
nor U24883 (N_24883,N_23639,N_23796);
or U24884 (N_24884,N_23266,N_23882);
xnor U24885 (N_24885,N_23262,N_23110);
nand U24886 (N_24886,N_23938,N_23784);
nor U24887 (N_24887,N_23893,N_23376);
or U24888 (N_24888,N_23942,N_23855);
xor U24889 (N_24889,N_23044,N_23551);
or U24890 (N_24890,N_23406,N_23276);
nor U24891 (N_24891,N_23648,N_23238);
nor U24892 (N_24892,N_23926,N_23427);
nand U24893 (N_24893,N_23495,N_23506);
xor U24894 (N_24894,N_23018,N_23289);
or U24895 (N_24895,N_23061,N_23666);
nand U24896 (N_24896,N_23385,N_23025);
nand U24897 (N_24897,N_23267,N_23236);
or U24898 (N_24898,N_23192,N_23605);
or U24899 (N_24899,N_23001,N_23379);
or U24900 (N_24900,N_23496,N_23444);
xor U24901 (N_24901,N_23152,N_23195);
and U24902 (N_24902,N_23861,N_23539);
and U24903 (N_24903,N_23349,N_23354);
or U24904 (N_24904,N_23009,N_23058);
and U24905 (N_24905,N_23376,N_23071);
nand U24906 (N_24906,N_23887,N_23965);
nand U24907 (N_24907,N_23803,N_23781);
nand U24908 (N_24908,N_23402,N_23840);
or U24909 (N_24909,N_23248,N_23996);
nand U24910 (N_24910,N_23171,N_23575);
nand U24911 (N_24911,N_23374,N_23798);
xor U24912 (N_24912,N_23022,N_23306);
nor U24913 (N_24913,N_23317,N_23387);
or U24914 (N_24914,N_23900,N_23509);
and U24915 (N_24915,N_23142,N_23955);
nor U24916 (N_24916,N_23293,N_23505);
xnor U24917 (N_24917,N_23565,N_23962);
xor U24918 (N_24918,N_23720,N_23082);
nand U24919 (N_24919,N_23623,N_23420);
nand U24920 (N_24920,N_23702,N_23248);
xor U24921 (N_24921,N_23468,N_23363);
and U24922 (N_24922,N_23609,N_23028);
xnor U24923 (N_24923,N_23982,N_23812);
nand U24924 (N_24924,N_23475,N_23573);
or U24925 (N_24925,N_23624,N_23519);
xor U24926 (N_24926,N_23809,N_23180);
and U24927 (N_24927,N_23272,N_23121);
and U24928 (N_24928,N_23686,N_23875);
nand U24929 (N_24929,N_23341,N_23135);
or U24930 (N_24930,N_23776,N_23223);
nor U24931 (N_24931,N_23893,N_23610);
nand U24932 (N_24932,N_23311,N_23301);
or U24933 (N_24933,N_23073,N_23268);
or U24934 (N_24934,N_23895,N_23300);
nand U24935 (N_24935,N_23780,N_23855);
nor U24936 (N_24936,N_23089,N_23730);
nor U24937 (N_24937,N_23395,N_23912);
nor U24938 (N_24938,N_23411,N_23180);
xnor U24939 (N_24939,N_23728,N_23142);
or U24940 (N_24940,N_23002,N_23138);
nor U24941 (N_24941,N_23418,N_23653);
or U24942 (N_24942,N_23819,N_23292);
or U24943 (N_24943,N_23097,N_23124);
xor U24944 (N_24944,N_23342,N_23194);
xnor U24945 (N_24945,N_23946,N_23344);
xnor U24946 (N_24946,N_23886,N_23825);
and U24947 (N_24947,N_23227,N_23847);
xor U24948 (N_24948,N_23392,N_23080);
xor U24949 (N_24949,N_23997,N_23479);
xor U24950 (N_24950,N_23979,N_23934);
nand U24951 (N_24951,N_23764,N_23064);
nor U24952 (N_24952,N_23786,N_23411);
or U24953 (N_24953,N_23051,N_23686);
and U24954 (N_24954,N_23537,N_23369);
or U24955 (N_24955,N_23997,N_23079);
nor U24956 (N_24956,N_23884,N_23140);
and U24957 (N_24957,N_23901,N_23928);
and U24958 (N_24958,N_23320,N_23421);
and U24959 (N_24959,N_23761,N_23604);
or U24960 (N_24960,N_23222,N_23736);
nor U24961 (N_24961,N_23064,N_23147);
or U24962 (N_24962,N_23933,N_23381);
xor U24963 (N_24963,N_23434,N_23334);
nor U24964 (N_24964,N_23216,N_23557);
xnor U24965 (N_24965,N_23010,N_23783);
and U24966 (N_24966,N_23681,N_23179);
or U24967 (N_24967,N_23593,N_23046);
and U24968 (N_24968,N_23915,N_23194);
nor U24969 (N_24969,N_23962,N_23626);
and U24970 (N_24970,N_23492,N_23336);
and U24971 (N_24971,N_23567,N_23738);
and U24972 (N_24972,N_23109,N_23897);
or U24973 (N_24973,N_23755,N_23910);
and U24974 (N_24974,N_23592,N_23169);
or U24975 (N_24975,N_23979,N_23959);
nor U24976 (N_24976,N_23932,N_23359);
and U24977 (N_24977,N_23807,N_23187);
xnor U24978 (N_24978,N_23215,N_23936);
xor U24979 (N_24979,N_23175,N_23994);
xor U24980 (N_24980,N_23144,N_23586);
or U24981 (N_24981,N_23804,N_23331);
and U24982 (N_24982,N_23837,N_23125);
nand U24983 (N_24983,N_23358,N_23186);
or U24984 (N_24984,N_23118,N_23680);
nand U24985 (N_24985,N_23023,N_23975);
nor U24986 (N_24986,N_23459,N_23510);
and U24987 (N_24987,N_23654,N_23595);
xor U24988 (N_24988,N_23742,N_23051);
nand U24989 (N_24989,N_23398,N_23812);
xor U24990 (N_24990,N_23578,N_23461);
and U24991 (N_24991,N_23069,N_23588);
and U24992 (N_24992,N_23867,N_23915);
nor U24993 (N_24993,N_23562,N_23682);
and U24994 (N_24994,N_23457,N_23244);
nand U24995 (N_24995,N_23240,N_23232);
nand U24996 (N_24996,N_23034,N_23594);
nor U24997 (N_24997,N_23405,N_23280);
nor U24998 (N_24998,N_23147,N_23150);
and U24999 (N_24999,N_23337,N_23866);
xor UO_0 (O_0,N_24752,N_24829);
and UO_1 (O_1,N_24265,N_24890);
nand UO_2 (O_2,N_24973,N_24836);
nand UO_3 (O_3,N_24669,N_24127);
and UO_4 (O_4,N_24364,N_24059);
nor UO_5 (O_5,N_24738,N_24828);
and UO_6 (O_6,N_24697,N_24012);
xor UO_7 (O_7,N_24916,N_24299);
and UO_8 (O_8,N_24856,N_24156);
and UO_9 (O_9,N_24923,N_24827);
nand UO_10 (O_10,N_24121,N_24011);
nor UO_11 (O_11,N_24833,N_24564);
or UO_12 (O_12,N_24720,N_24897);
or UO_13 (O_13,N_24850,N_24427);
xor UO_14 (O_14,N_24096,N_24302);
xnor UO_15 (O_15,N_24081,N_24583);
nand UO_16 (O_16,N_24612,N_24538);
nor UO_17 (O_17,N_24470,N_24045);
or UO_18 (O_18,N_24180,N_24591);
or UO_19 (O_19,N_24805,N_24970);
nand UO_20 (O_20,N_24404,N_24608);
nor UO_21 (O_21,N_24135,N_24319);
xor UO_22 (O_22,N_24210,N_24702);
and UO_23 (O_23,N_24922,N_24606);
nor UO_24 (O_24,N_24871,N_24467);
or UO_25 (O_25,N_24323,N_24230);
nor UO_26 (O_26,N_24595,N_24682);
nor UO_27 (O_27,N_24434,N_24285);
or UO_28 (O_28,N_24561,N_24069);
nor UO_29 (O_29,N_24061,N_24109);
nand UO_30 (O_30,N_24423,N_24863);
nand UO_31 (O_31,N_24887,N_24052);
and UO_32 (O_32,N_24477,N_24563);
xor UO_33 (O_33,N_24892,N_24504);
xor UO_34 (O_34,N_24645,N_24592);
nor UO_35 (O_35,N_24830,N_24308);
and UO_36 (O_36,N_24484,N_24318);
or UO_37 (O_37,N_24353,N_24841);
xnor UO_38 (O_38,N_24558,N_24773);
nand UO_39 (O_39,N_24200,N_24220);
or UO_40 (O_40,N_24853,N_24243);
nand UO_41 (O_41,N_24118,N_24776);
or UO_42 (O_42,N_24932,N_24018);
and UO_43 (O_43,N_24029,N_24236);
nand UO_44 (O_44,N_24361,N_24491);
or UO_45 (O_45,N_24153,N_24198);
or UO_46 (O_46,N_24092,N_24646);
or UO_47 (O_47,N_24630,N_24884);
nor UO_48 (O_48,N_24136,N_24786);
or UO_49 (O_49,N_24722,N_24940);
or UO_50 (O_50,N_24909,N_24005);
and UO_51 (O_51,N_24448,N_24677);
or UO_52 (O_52,N_24024,N_24389);
or UO_53 (O_53,N_24769,N_24750);
nor UO_54 (O_54,N_24142,N_24600);
or UO_55 (O_55,N_24295,N_24416);
nand UO_56 (O_56,N_24380,N_24577);
or UO_57 (O_57,N_24067,N_24370);
and UO_58 (O_58,N_24189,N_24687);
or UO_59 (O_59,N_24958,N_24398);
nand UO_60 (O_60,N_24329,N_24823);
and UO_61 (O_61,N_24988,N_24694);
and UO_62 (O_62,N_24026,N_24399);
nor UO_63 (O_63,N_24528,N_24882);
xor UO_64 (O_64,N_24306,N_24986);
nand UO_65 (O_65,N_24290,N_24886);
nand UO_66 (O_66,N_24521,N_24326);
nor UO_67 (O_67,N_24551,N_24084);
and UO_68 (O_68,N_24861,N_24032);
nor UO_69 (O_69,N_24078,N_24145);
xnor UO_70 (O_70,N_24411,N_24334);
or UO_71 (O_71,N_24758,N_24281);
nand UO_72 (O_72,N_24545,N_24849);
or UO_73 (O_73,N_24679,N_24048);
nor UO_74 (O_74,N_24880,N_24794);
or UO_75 (O_75,N_24971,N_24692);
and UO_76 (O_76,N_24475,N_24409);
xor UO_77 (O_77,N_24859,N_24186);
nand UO_78 (O_78,N_24071,N_24928);
xor UO_79 (O_79,N_24944,N_24060);
nand UO_80 (O_80,N_24384,N_24190);
nor UO_81 (O_81,N_24267,N_24251);
and UO_82 (O_82,N_24047,N_24675);
nor UO_83 (O_83,N_24622,N_24670);
and UO_84 (O_84,N_24253,N_24063);
xnor UO_85 (O_85,N_24599,N_24442);
xnor UO_86 (O_86,N_24690,N_24161);
nor UO_87 (O_87,N_24468,N_24004);
and UO_88 (O_88,N_24627,N_24057);
xnor UO_89 (O_89,N_24676,N_24607);
xor UO_90 (O_90,N_24644,N_24369);
and UO_91 (O_91,N_24357,N_24378);
and UO_92 (O_92,N_24996,N_24201);
or UO_93 (O_93,N_24987,N_24065);
xor UO_94 (O_94,N_24574,N_24068);
nand UO_95 (O_95,N_24403,N_24050);
nor UO_96 (O_96,N_24616,N_24260);
xnor UO_97 (O_97,N_24426,N_24725);
or UO_98 (O_98,N_24402,N_24937);
nand UO_99 (O_99,N_24549,N_24994);
and UO_100 (O_100,N_24870,N_24862);
nor UO_101 (O_101,N_24680,N_24934);
xor UO_102 (O_102,N_24513,N_24514);
and UO_103 (O_103,N_24779,N_24215);
xor UO_104 (O_104,N_24383,N_24406);
and UO_105 (O_105,N_24494,N_24228);
or UO_106 (O_106,N_24959,N_24553);
or UO_107 (O_107,N_24347,N_24424);
xnor UO_108 (O_108,N_24258,N_24157);
nand UO_109 (O_109,N_24536,N_24554);
nor UO_110 (O_110,N_24245,N_24927);
or UO_111 (O_111,N_24386,N_24395);
nand UO_112 (O_112,N_24798,N_24183);
and UO_113 (O_113,N_24101,N_24232);
or UO_114 (O_114,N_24981,N_24704);
nor UO_115 (O_115,N_24873,N_24410);
xnor UO_116 (O_116,N_24723,N_24962);
xnor UO_117 (O_117,N_24175,N_24789);
and UO_118 (O_118,N_24901,N_24147);
xor UO_119 (O_119,N_24575,N_24103);
and UO_120 (O_120,N_24246,N_24053);
or UO_121 (O_121,N_24846,N_24414);
or UO_122 (O_122,N_24191,N_24605);
nor UO_123 (O_123,N_24681,N_24801);
xnor UO_124 (O_124,N_24977,N_24782);
xor UO_125 (O_125,N_24594,N_24234);
and UO_126 (O_126,N_24469,N_24982);
or UO_127 (O_127,N_24471,N_24479);
or UO_128 (O_128,N_24743,N_24685);
or UO_129 (O_129,N_24073,N_24998);
and UO_130 (O_130,N_24822,N_24523);
and UO_131 (O_131,N_24194,N_24847);
and UO_132 (O_132,N_24464,N_24272);
nand UO_133 (O_133,N_24167,N_24811);
and UO_134 (O_134,N_24223,N_24524);
or UO_135 (O_135,N_24008,N_24054);
nand UO_136 (O_136,N_24095,N_24356);
nand UO_137 (O_137,N_24613,N_24902);
xnor UO_138 (O_138,N_24333,N_24345);
or UO_139 (O_139,N_24120,N_24899);
and UO_140 (O_140,N_24585,N_24804);
and UO_141 (O_141,N_24858,N_24244);
and UO_142 (O_142,N_24891,N_24535);
and UO_143 (O_143,N_24555,N_24799);
or UO_144 (O_144,N_24039,N_24074);
and UO_145 (O_145,N_24221,N_24287);
and UO_146 (O_146,N_24114,N_24313);
xor UO_147 (O_147,N_24653,N_24527);
or UO_148 (O_148,N_24289,N_24310);
or UO_149 (O_149,N_24286,N_24755);
xnor UO_150 (O_150,N_24044,N_24911);
xnor UO_151 (O_151,N_24502,N_24956);
nor UO_152 (O_152,N_24541,N_24777);
nor UO_153 (O_153,N_24122,N_24275);
nor UO_154 (O_154,N_24297,N_24560);
xnor UO_155 (O_155,N_24741,N_24311);
and UO_156 (O_156,N_24445,N_24633);
and UO_157 (O_157,N_24879,N_24898);
and UO_158 (O_158,N_24664,N_24842);
xnor UO_159 (O_159,N_24990,N_24543);
or UO_160 (O_160,N_24385,N_24444);
nor UO_161 (O_161,N_24531,N_24184);
and UO_162 (O_162,N_24452,N_24581);
xor UO_163 (O_163,N_24337,N_24446);
nand UO_164 (O_164,N_24611,N_24056);
or UO_165 (O_165,N_24893,N_24497);
or UO_166 (O_166,N_24785,N_24344);
and UO_167 (O_167,N_24178,N_24261);
and UO_168 (O_168,N_24710,N_24817);
xnor UO_169 (O_169,N_24678,N_24952);
nor UO_170 (O_170,N_24010,N_24131);
nor UO_171 (O_171,N_24819,N_24740);
and UO_172 (O_172,N_24701,N_24854);
and UO_173 (O_173,N_24572,N_24516);
nand UO_174 (O_174,N_24413,N_24803);
nor UO_175 (O_175,N_24980,N_24134);
and UO_176 (O_176,N_24498,N_24300);
nand UO_177 (O_177,N_24759,N_24844);
nand UO_178 (O_178,N_24576,N_24624);
nand UO_179 (O_179,N_24366,N_24001);
or UO_180 (O_180,N_24511,N_24150);
nand UO_181 (O_181,N_24584,N_24152);
and UO_182 (O_182,N_24800,N_24992);
or UO_183 (O_183,N_24983,N_24542);
nand UO_184 (O_184,N_24518,N_24788);
xnor UO_185 (O_185,N_24734,N_24492);
and UO_186 (O_186,N_24111,N_24270);
xor UO_187 (O_187,N_24818,N_24271);
xnor UO_188 (O_188,N_24195,N_24124);
nor UO_189 (O_189,N_24003,N_24371);
nand UO_190 (O_190,N_24359,N_24128);
xnor UO_191 (O_191,N_24058,N_24415);
xnor UO_192 (O_192,N_24375,N_24877);
nor UO_193 (O_193,N_24835,N_24192);
and UO_194 (O_194,N_24064,N_24708);
or UO_195 (O_195,N_24137,N_24255);
or UO_196 (O_196,N_24571,N_24288);
nand UO_197 (O_197,N_24354,N_24099);
nand UO_198 (O_198,N_24961,N_24166);
xnor UO_199 (O_199,N_24187,N_24489);
and UO_200 (O_200,N_24957,N_24941);
and UO_201 (O_201,N_24515,N_24509);
or UO_202 (O_202,N_24763,N_24618);
xor UO_203 (O_203,N_24802,N_24568);
or UO_204 (O_204,N_24089,N_24193);
xor UO_205 (O_205,N_24066,N_24778);
nand UO_206 (O_206,N_24904,N_24642);
nor UO_207 (O_207,N_24433,N_24082);
and UO_208 (O_208,N_24628,N_24666);
nor UO_209 (O_209,N_24632,N_24430);
or UO_210 (O_210,N_24014,N_24865);
and UO_211 (O_211,N_24231,N_24726);
or UO_212 (O_212,N_24519,N_24869);
or UO_213 (O_213,N_24108,N_24159);
nor UO_214 (O_214,N_24698,N_24205);
or UO_215 (O_215,N_24390,N_24007);
xnor UO_216 (O_216,N_24761,N_24894);
or UO_217 (O_217,N_24325,N_24247);
nand UO_218 (O_218,N_24506,N_24783);
nor UO_219 (O_219,N_24459,N_24368);
and UO_220 (O_220,N_24090,N_24428);
nor UO_221 (O_221,N_24674,N_24874);
or UO_222 (O_222,N_24718,N_24550);
nand UO_223 (O_223,N_24917,N_24663);
nand UO_224 (O_224,N_24753,N_24105);
xnor UO_225 (O_225,N_24924,N_24578);
nor UO_226 (O_226,N_24895,N_24787);
nor UO_227 (O_227,N_24626,N_24635);
or UO_228 (O_228,N_24340,N_24587);
nor UO_229 (O_229,N_24652,N_24305);
xor UO_230 (O_230,N_24582,N_24490);
nand UO_231 (O_231,N_24714,N_24388);
and UO_232 (O_232,N_24387,N_24206);
nand UO_233 (O_233,N_24651,N_24684);
and UO_234 (O_234,N_24338,N_24921);
nand UO_235 (O_235,N_24840,N_24765);
or UO_236 (O_236,N_24526,N_24408);
nand UO_237 (O_237,N_24107,N_24482);
xor UO_238 (O_238,N_24950,N_24900);
or UO_239 (O_239,N_24707,N_24915);
xnor UO_240 (O_240,N_24177,N_24216);
and UO_241 (O_241,N_24252,N_24170);
or UO_242 (O_242,N_24693,N_24512);
nand UO_243 (O_243,N_24224,N_24327);
nand UO_244 (O_244,N_24620,N_24453);
or UO_245 (O_245,N_24144,N_24440);
nor UO_246 (O_246,N_24042,N_24372);
xor UO_247 (O_247,N_24838,N_24314);
and UO_248 (O_248,N_24839,N_24637);
nor UO_249 (O_249,N_24461,N_24396);
or UO_250 (O_250,N_24165,N_24552);
nand UO_251 (O_251,N_24181,N_24997);
nor UO_252 (O_252,N_24748,N_24631);
and UO_253 (O_253,N_24226,N_24619);
nor UO_254 (O_254,N_24093,N_24363);
xnor UO_255 (O_255,N_24196,N_24610);
nor UO_256 (O_256,N_24049,N_24905);
and UO_257 (O_257,N_24713,N_24559);
nand UO_258 (O_258,N_24907,N_24481);
xor UO_259 (O_259,N_24984,N_24328);
or UO_260 (O_260,N_24331,N_24925);
xnor UO_261 (O_261,N_24780,N_24496);
nor UO_262 (O_262,N_24155,N_24179);
or UO_263 (O_263,N_24355,N_24382);
xnor UO_264 (O_264,N_24022,N_24037);
or UO_265 (O_265,N_24813,N_24379);
nand UO_266 (O_266,N_24881,N_24432);
and UO_267 (O_267,N_24562,N_24168);
xor UO_268 (O_268,N_24070,N_24235);
and UO_269 (O_269,N_24154,N_24254);
or UO_270 (O_270,N_24762,N_24140);
nand UO_271 (O_271,N_24149,N_24636);
xor UO_272 (O_272,N_24995,N_24087);
nand UO_273 (O_273,N_24298,N_24505);
or UO_274 (O_274,N_24797,N_24548);
nand UO_275 (O_275,N_24671,N_24487);
or UO_276 (O_276,N_24367,N_24274);
and UO_277 (O_277,N_24656,N_24742);
nand UO_278 (O_278,N_24377,N_24604);
nor UO_279 (O_279,N_24754,N_24781);
and UO_280 (O_280,N_24162,N_24991);
or UO_281 (O_281,N_24943,N_24673);
nor UO_282 (O_282,N_24113,N_24979);
nor UO_283 (O_283,N_24381,N_24421);
nor UO_284 (O_284,N_24848,N_24534);
nor UO_285 (O_285,N_24972,N_24086);
and UO_286 (O_286,N_24598,N_24951);
nand UO_287 (O_287,N_24277,N_24662);
xor UO_288 (O_288,N_24532,N_24503);
nor UO_289 (O_289,N_24625,N_24213);
and UO_290 (O_290,N_24451,N_24936);
and UO_291 (O_291,N_24807,N_24463);
or UO_292 (O_292,N_24906,N_24772);
and UO_293 (O_293,N_24346,N_24160);
xnor UO_294 (O_294,N_24106,N_24358);
and UO_295 (O_295,N_24641,N_24974);
nor UO_296 (O_296,N_24292,N_24164);
nand UO_297 (O_297,N_24278,N_24659);
and UO_298 (O_298,N_24197,N_24621);
and UO_299 (O_299,N_24094,N_24110);
or UO_300 (O_300,N_24117,N_24914);
or UO_301 (O_301,N_24420,N_24696);
or UO_302 (O_302,N_24953,N_24309);
nand UO_303 (O_303,N_24209,N_24472);
xor UO_304 (O_304,N_24138,N_24699);
nor UO_305 (O_305,N_24268,N_24365);
nand UO_306 (O_306,N_24603,N_24654);
nand UO_307 (O_307,N_24163,N_24046);
xnor UO_308 (O_308,N_24257,N_24510);
and UO_309 (O_309,N_24174,N_24352);
nand UO_310 (O_310,N_24435,N_24954);
xor UO_311 (O_311,N_24454,N_24775);
nand UO_312 (O_312,N_24806,N_24668);
and UO_313 (O_313,N_24968,N_24263);
nor UO_314 (O_314,N_24883,N_24458);
and UO_315 (O_315,N_24264,N_24650);
and UO_316 (O_316,N_24332,N_24493);
or UO_317 (O_317,N_24965,N_24872);
nor UO_318 (O_318,N_24586,N_24691);
nand UO_319 (O_319,N_24960,N_24784);
and UO_320 (O_320,N_24262,N_24985);
nor UO_321 (O_321,N_24062,N_24028);
nand UO_322 (O_322,N_24700,N_24544);
xnor UO_323 (O_323,N_24296,N_24975);
nor UO_324 (O_324,N_24072,N_24273);
xnor UO_325 (O_325,N_24918,N_24649);
xnor UO_326 (O_326,N_24567,N_24412);
nor UO_327 (O_327,N_24425,N_24589);
or UO_328 (O_328,N_24455,N_24225);
nand UO_329 (O_329,N_24141,N_24341);
or UO_330 (O_330,N_24303,N_24351);
nand UO_331 (O_331,N_24736,N_24279);
xor UO_332 (O_332,N_24746,N_24580);
or UO_333 (O_333,N_24908,N_24967);
xnor UO_334 (O_334,N_24422,N_24115);
and UO_335 (O_335,N_24537,N_24768);
xnor UO_336 (O_336,N_24085,N_24033);
or UO_337 (O_337,N_24728,N_24031);
nand UO_338 (O_338,N_24293,N_24143);
nor UO_339 (O_339,N_24040,N_24130);
nand UO_340 (O_340,N_24266,N_24876);
and UO_341 (O_341,N_24926,N_24000);
xor UO_342 (O_342,N_24912,N_24450);
xnor UO_343 (O_343,N_24233,N_24376);
nor UO_344 (O_344,N_24397,N_24051);
nor UO_345 (O_345,N_24792,N_24570);
or UO_346 (O_346,N_24030,N_24816);
and UO_347 (O_347,N_24188,N_24832);
nor UO_348 (O_348,N_24724,N_24756);
nor UO_349 (O_349,N_24688,N_24217);
xor UO_350 (O_350,N_24500,N_24417);
or UO_351 (O_351,N_24540,N_24208);
nand UO_352 (O_352,N_24851,N_24431);
nand UO_353 (O_353,N_24878,N_24204);
xnor UO_354 (O_354,N_24336,N_24350);
nor UO_355 (O_355,N_24931,N_24182);
nor UO_356 (O_356,N_24933,N_24569);
or UO_357 (O_357,N_24533,N_24439);
and UO_358 (O_358,N_24767,N_24240);
xor UO_359 (O_359,N_24034,N_24989);
or UO_360 (O_360,N_24837,N_24812);
or UO_361 (O_361,N_24449,N_24834);
nor UO_362 (O_362,N_24035,N_24711);
nor UO_363 (O_363,N_24885,N_24719);
xor UO_364 (O_364,N_24655,N_24036);
or UO_365 (O_365,N_24815,N_24176);
xor UO_366 (O_366,N_24362,N_24083);
and UO_367 (O_367,N_24316,N_24112);
or UO_368 (O_368,N_24660,N_24405);
nand UO_369 (O_369,N_24732,N_24517);
xnor UO_370 (O_370,N_24485,N_24460);
or UO_371 (O_371,N_24025,N_24831);
nor UO_372 (O_372,N_24712,N_24969);
or UO_373 (O_373,N_24733,N_24947);
xnor UO_374 (O_374,N_24826,N_24639);
nand UO_375 (O_375,N_24942,N_24283);
nor UO_376 (O_376,N_24966,N_24602);
xnor UO_377 (O_377,N_24629,N_24237);
or UO_378 (O_378,N_24443,N_24465);
and UO_379 (O_379,N_24407,N_24749);
and UO_380 (O_380,N_24038,N_24955);
and UO_381 (O_381,N_24825,N_24557);
and UO_382 (O_382,N_24438,N_24250);
xor UO_383 (O_383,N_24593,N_24116);
and UO_384 (O_384,N_24091,N_24343);
xor UO_385 (O_385,N_24614,N_24665);
xnor UO_386 (O_386,N_24875,N_24808);
nor UO_387 (O_387,N_24330,N_24868);
xnor UO_388 (O_388,N_24020,N_24457);
or UO_389 (O_389,N_24796,N_24658);
nor UO_390 (O_390,N_24843,N_24478);
nor UO_391 (O_391,N_24978,N_24055);
and UO_392 (O_392,N_24565,N_24339);
nor UO_393 (O_393,N_24946,N_24320);
nor UO_394 (O_394,N_24400,N_24256);
xor UO_395 (O_395,N_24889,N_24342);
nand UO_396 (O_396,N_24214,N_24219);
xnor UO_397 (O_397,N_24790,N_24689);
nor UO_398 (O_398,N_24348,N_24896);
nor UO_399 (O_399,N_24123,N_24315);
xnor UO_400 (O_400,N_24716,N_24771);
xnor UO_401 (O_401,N_24102,N_24418);
nand UO_402 (O_402,N_24335,N_24867);
nor UO_403 (O_403,N_24860,N_24737);
xnor UO_404 (O_404,N_24088,N_24705);
and UO_405 (O_405,N_24019,N_24855);
nor UO_406 (O_406,N_24488,N_24211);
nor UO_407 (O_407,N_24016,N_24764);
or UO_408 (O_408,N_24770,N_24317);
or UO_409 (O_409,N_24814,N_24703);
nor UO_410 (O_410,N_24791,N_24321);
xnor UO_411 (O_411,N_24667,N_24312);
nand UO_412 (O_412,N_24239,N_24027);
xor UO_413 (O_413,N_24280,N_24766);
nand UO_414 (O_414,N_24579,N_24647);
nand UO_415 (O_415,N_24683,N_24075);
or UO_416 (O_416,N_24623,N_24546);
and UO_417 (O_417,N_24269,N_24419);
and UO_418 (O_418,N_24935,N_24999);
nor UO_419 (O_419,N_24360,N_24119);
and UO_420 (O_420,N_24507,N_24810);
and UO_421 (O_421,N_24919,N_24930);
nor UO_422 (O_422,N_24002,N_24238);
nor UO_423 (O_423,N_24203,N_24373);
nor UO_424 (O_424,N_24474,N_24171);
xnor UO_425 (O_425,N_24132,N_24638);
nor UO_426 (O_426,N_24158,N_24076);
nor UO_427 (O_427,N_24597,N_24199);
and UO_428 (O_428,N_24501,N_24888);
nor UO_429 (O_429,N_24709,N_24148);
nor UO_430 (O_430,N_24715,N_24249);
or UO_431 (O_431,N_24522,N_24207);
or UO_432 (O_432,N_24735,N_24282);
xnor UO_433 (O_433,N_24672,N_24126);
or UO_434 (O_434,N_24686,N_24437);
xnor UO_435 (O_435,N_24080,N_24222);
nor UO_436 (O_436,N_24456,N_24248);
nor UO_437 (O_437,N_24539,N_24009);
nand UO_438 (O_438,N_24401,N_24948);
and UO_439 (O_439,N_24747,N_24596);
or UO_440 (O_440,N_24774,N_24634);
nand UO_441 (O_441,N_24169,N_24441);
nand UO_442 (O_442,N_24436,N_24307);
nor UO_443 (O_443,N_24098,N_24721);
xnor UO_444 (O_444,N_24304,N_24483);
or UO_445 (O_445,N_24508,N_24963);
and UO_446 (O_446,N_24964,N_24617);
nand UO_447 (O_447,N_24609,N_24100);
xnor UO_448 (O_448,N_24525,N_24125);
nand UO_449 (O_449,N_24648,N_24473);
nand UO_450 (O_450,N_24601,N_24104);
nor UO_451 (O_451,N_24391,N_24015);
nor UO_452 (O_452,N_24910,N_24173);
nor UO_453 (O_453,N_24976,N_24041);
or UO_454 (O_454,N_24129,N_24023);
nand UO_455 (O_455,N_24938,N_24097);
or UO_456 (O_456,N_24706,N_24202);
nor UO_457 (O_457,N_24151,N_24229);
xor UO_458 (O_458,N_24845,N_24920);
nor UO_459 (O_459,N_24729,N_24824);
xor UO_460 (O_460,N_24556,N_24727);
nand UO_461 (O_461,N_24520,N_24745);
nand UO_462 (O_462,N_24429,N_24913);
or UO_463 (O_463,N_24573,N_24466);
xor UO_464 (O_464,N_24476,N_24043);
or UO_465 (O_465,N_24751,N_24394);
and UO_466 (O_466,N_24480,N_24757);
nand UO_467 (O_467,N_24857,N_24218);
nor UO_468 (O_468,N_24259,N_24486);
xnor UO_469 (O_469,N_24013,N_24566);
or UO_470 (O_470,N_24730,N_24939);
nand UO_471 (O_471,N_24657,N_24462);
nand UO_472 (O_472,N_24284,N_24447);
nand UO_473 (O_473,N_24006,N_24017);
or UO_474 (O_474,N_24294,N_24241);
xor UO_475 (O_475,N_24077,N_24276);
nand UO_476 (O_476,N_24793,N_24301);
nor UO_477 (O_477,N_24821,N_24392);
nor UO_478 (O_478,N_24530,N_24949);
nand UO_479 (O_479,N_24588,N_24795);
or UO_480 (O_480,N_24615,N_24744);
and UO_481 (O_481,N_24852,N_24393);
nand UO_482 (O_482,N_24324,N_24864);
nor UO_483 (O_483,N_24322,N_24499);
nand UO_484 (O_484,N_24809,N_24227);
nand UO_485 (O_485,N_24640,N_24139);
nand UO_486 (O_486,N_24717,N_24212);
and UO_487 (O_487,N_24661,N_24242);
nand UO_488 (O_488,N_24945,N_24993);
nand UO_489 (O_489,N_24760,N_24133);
nand UO_490 (O_490,N_24291,N_24820);
nor UO_491 (O_491,N_24695,N_24547);
nand UO_492 (O_492,N_24146,N_24021);
nor UO_493 (O_493,N_24929,N_24643);
nand UO_494 (O_494,N_24739,N_24731);
and UO_495 (O_495,N_24529,N_24866);
nor UO_496 (O_496,N_24495,N_24374);
nand UO_497 (O_497,N_24185,N_24590);
nand UO_498 (O_498,N_24349,N_24079);
or UO_499 (O_499,N_24903,N_24172);
nor UO_500 (O_500,N_24379,N_24734);
xor UO_501 (O_501,N_24225,N_24907);
or UO_502 (O_502,N_24185,N_24460);
nor UO_503 (O_503,N_24251,N_24592);
or UO_504 (O_504,N_24144,N_24723);
xnor UO_505 (O_505,N_24166,N_24171);
nand UO_506 (O_506,N_24396,N_24976);
nand UO_507 (O_507,N_24964,N_24737);
xnor UO_508 (O_508,N_24596,N_24257);
or UO_509 (O_509,N_24409,N_24807);
xor UO_510 (O_510,N_24088,N_24026);
nor UO_511 (O_511,N_24470,N_24372);
and UO_512 (O_512,N_24409,N_24191);
or UO_513 (O_513,N_24554,N_24131);
xnor UO_514 (O_514,N_24496,N_24985);
nand UO_515 (O_515,N_24317,N_24559);
nand UO_516 (O_516,N_24805,N_24224);
and UO_517 (O_517,N_24303,N_24214);
nor UO_518 (O_518,N_24254,N_24363);
nor UO_519 (O_519,N_24379,N_24610);
xor UO_520 (O_520,N_24273,N_24489);
nor UO_521 (O_521,N_24178,N_24950);
nand UO_522 (O_522,N_24854,N_24793);
nand UO_523 (O_523,N_24329,N_24237);
and UO_524 (O_524,N_24638,N_24807);
nor UO_525 (O_525,N_24848,N_24938);
nor UO_526 (O_526,N_24821,N_24976);
nor UO_527 (O_527,N_24315,N_24263);
or UO_528 (O_528,N_24067,N_24736);
or UO_529 (O_529,N_24594,N_24579);
or UO_530 (O_530,N_24447,N_24184);
nand UO_531 (O_531,N_24150,N_24400);
or UO_532 (O_532,N_24310,N_24211);
xor UO_533 (O_533,N_24426,N_24390);
and UO_534 (O_534,N_24073,N_24348);
or UO_535 (O_535,N_24447,N_24245);
nand UO_536 (O_536,N_24802,N_24368);
nand UO_537 (O_537,N_24703,N_24487);
nand UO_538 (O_538,N_24210,N_24600);
nor UO_539 (O_539,N_24342,N_24657);
xor UO_540 (O_540,N_24805,N_24649);
nor UO_541 (O_541,N_24555,N_24913);
xor UO_542 (O_542,N_24196,N_24455);
and UO_543 (O_543,N_24682,N_24208);
nor UO_544 (O_544,N_24388,N_24688);
and UO_545 (O_545,N_24118,N_24581);
or UO_546 (O_546,N_24325,N_24122);
or UO_547 (O_547,N_24556,N_24819);
and UO_548 (O_548,N_24554,N_24101);
xor UO_549 (O_549,N_24619,N_24198);
and UO_550 (O_550,N_24367,N_24781);
nand UO_551 (O_551,N_24135,N_24250);
or UO_552 (O_552,N_24688,N_24210);
and UO_553 (O_553,N_24983,N_24225);
nor UO_554 (O_554,N_24866,N_24896);
and UO_555 (O_555,N_24176,N_24109);
or UO_556 (O_556,N_24929,N_24528);
or UO_557 (O_557,N_24956,N_24673);
and UO_558 (O_558,N_24644,N_24354);
nor UO_559 (O_559,N_24981,N_24001);
and UO_560 (O_560,N_24425,N_24549);
xor UO_561 (O_561,N_24749,N_24747);
nand UO_562 (O_562,N_24536,N_24093);
and UO_563 (O_563,N_24495,N_24848);
nand UO_564 (O_564,N_24175,N_24208);
nand UO_565 (O_565,N_24595,N_24765);
or UO_566 (O_566,N_24037,N_24979);
and UO_567 (O_567,N_24830,N_24186);
xnor UO_568 (O_568,N_24865,N_24921);
nor UO_569 (O_569,N_24063,N_24122);
nor UO_570 (O_570,N_24611,N_24980);
nand UO_571 (O_571,N_24943,N_24061);
nor UO_572 (O_572,N_24703,N_24245);
nand UO_573 (O_573,N_24109,N_24653);
or UO_574 (O_574,N_24635,N_24399);
and UO_575 (O_575,N_24011,N_24659);
nor UO_576 (O_576,N_24567,N_24646);
and UO_577 (O_577,N_24110,N_24585);
nor UO_578 (O_578,N_24944,N_24566);
and UO_579 (O_579,N_24573,N_24062);
or UO_580 (O_580,N_24809,N_24368);
and UO_581 (O_581,N_24896,N_24135);
nor UO_582 (O_582,N_24563,N_24250);
xnor UO_583 (O_583,N_24040,N_24653);
xor UO_584 (O_584,N_24181,N_24226);
nand UO_585 (O_585,N_24429,N_24226);
nor UO_586 (O_586,N_24629,N_24711);
xnor UO_587 (O_587,N_24130,N_24568);
and UO_588 (O_588,N_24539,N_24553);
nor UO_589 (O_589,N_24587,N_24304);
or UO_590 (O_590,N_24117,N_24832);
nor UO_591 (O_591,N_24323,N_24179);
or UO_592 (O_592,N_24331,N_24735);
nand UO_593 (O_593,N_24589,N_24917);
or UO_594 (O_594,N_24996,N_24080);
nand UO_595 (O_595,N_24897,N_24226);
or UO_596 (O_596,N_24941,N_24744);
xor UO_597 (O_597,N_24393,N_24080);
or UO_598 (O_598,N_24528,N_24751);
nand UO_599 (O_599,N_24451,N_24679);
nand UO_600 (O_600,N_24982,N_24663);
or UO_601 (O_601,N_24912,N_24293);
and UO_602 (O_602,N_24261,N_24119);
and UO_603 (O_603,N_24522,N_24600);
nor UO_604 (O_604,N_24391,N_24308);
nor UO_605 (O_605,N_24358,N_24565);
nor UO_606 (O_606,N_24372,N_24514);
and UO_607 (O_607,N_24466,N_24990);
and UO_608 (O_608,N_24061,N_24718);
nor UO_609 (O_609,N_24419,N_24223);
nand UO_610 (O_610,N_24484,N_24730);
nor UO_611 (O_611,N_24700,N_24639);
nor UO_612 (O_612,N_24171,N_24504);
xor UO_613 (O_613,N_24344,N_24788);
nor UO_614 (O_614,N_24989,N_24298);
and UO_615 (O_615,N_24906,N_24932);
nor UO_616 (O_616,N_24079,N_24064);
nor UO_617 (O_617,N_24402,N_24595);
xnor UO_618 (O_618,N_24109,N_24005);
or UO_619 (O_619,N_24708,N_24028);
and UO_620 (O_620,N_24308,N_24300);
or UO_621 (O_621,N_24892,N_24894);
xnor UO_622 (O_622,N_24098,N_24934);
nand UO_623 (O_623,N_24594,N_24463);
or UO_624 (O_624,N_24659,N_24904);
nand UO_625 (O_625,N_24887,N_24081);
and UO_626 (O_626,N_24182,N_24912);
xor UO_627 (O_627,N_24912,N_24475);
or UO_628 (O_628,N_24076,N_24377);
or UO_629 (O_629,N_24788,N_24617);
or UO_630 (O_630,N_24614,N_24337);
or UO_631 (O_631,N_24990,N_24290);
xor UO_632 (O_632,N_24979,N_24027);
and UO_633 (O_633,N_24056,N_24656);
xor UO_634 (O_634,N_24355,N_24070);
nand UO_635 (O_635,N_24171,N_24025);
nor UO_636 (O_636,N_24423,N_24252);
and UO_637 (O_637,N_24049,N_24633);
or UO_638 (O_638,N_24857,N_24972);
and UO_639 (O_639,N_24315,N_24045);
xnor UO_640 (O_640,N_24529,N_24675);
nand UO_641 (O_641,N_24453,N_24352);
xnor UO_642 (O_642,N_24879,N_24069);
or UO_643 (O_643,N_24200,N_24533);
nand UO_644 (O_644,N_24424,N_24814);
xnor UO_645 (O_645,N_24566,N_24108);
nand UO_646 (O_646,N_24852,N_24030);
nand UO_647 (O_647,N_24098,N_24574);
and UO_648 (O_648,N_24845,N_24188);
and UO_649 (O_649,N_24378,N_24773);
and UO_650 (O_650,N_24559,N_24095);
nand UO_651 (O_651,N_24072,N_24417);
xnor UO_652 (O_652,N_24077,N_24237);
and UO_653 (O_653,N_24751,N_24189);
and UO_654 (O_654,N_24442,N_24405);
nor UO_655 (O_655,N_24550,N_24473);
nor UO_656 (O_656,N_24219,N_24629);
xor UO_657 (O_657,N_24870,N_24732);
xor UO_658 (O_658,N_24026,N_24306);
and UO_659 (O_659,N_24902,N_24184);
xor UO_660 (O_660,N_24305,N_24522);
nor UO_661 (O_661,N_24472,N_24659);
or UO_662 (O_662,N_24650,N_24474);
nor UO_663 (O_663,N_24528,N_24416);
xor UO_664 (O_664,N_24221,N_24306);
and UO_665 (O_665,N_24808,N_24756);
and UO_666 (O_666,N_24529,N_24587);
nand UO_667 (O_667,N_24613,N_24932);
or UO_668 (O_668,N_24373,N_24640);
nor UO_669 (O_669,N_24033,N_24100);
or UO_670 (O_670,N_24956,N_24147);
nand UO_671 (O_671,N_24779,N_24478);
and UO_672 (O_672,N_24448,N_24026);
nand UO_673 (O_673,N_24048,N_24576);
nand UO_674 (O_674,N_24423,N_24766);
or UO_675 (O_675,N_24619,N_24803);
and UO_676 (O_676,N_24617,N_24875);
xnor UO_677 (O_677,N_24733,N_24246);
xor UO_678 (O_678,N_24381,N_24270);
xor UO_679 (O_679,N_24180,N_24437);
nor UO_680 (O_680,N_24129,N_24610);
and UO_681 (O_681,N_24299,N_24933);
and UO_682 (O_682,N_24253,N_24298);
or UO_683 (O_683,N_24306,N_24970);
and UO_684 (O_684,N_24791,N_24188);
nor UO_685 (O_685,N_24564,N_24227);
or UO_686 (O_686,N_24213,N_24030);
and UO_687 (O_687,N_24081,N_24776);
or UO_688 (O_688,N_24501,N_24366);
nor UO_689 (O_689,N_24212,N_24348);
or UO_690 (O_690,N_24360,N_24335);
or UO_691 (O_691,N_24526,N_24974);
and UO_692 (O_692,N_24960,N_24516);
xor UO_693 (O_693,N_24165,N_24629);
xnor UO_694 (O_694,N_24107,N_24492);
or UO_695 (O_695,N_24915,N_24429);
or UO_696 (O_696,N_24648,N_24588);
or UO_697 (O_697,N_24405,N_24147);
and UO_698 (O_698,N_24720,N_24112);
nand UO_699 (O_699,N_24905,N_24232);
nand UO_700 (O_700,N_24740,N_24054);
or UO_701 (O_701,N_24279,N_24636);
xor UO_702 (O_702,N_24763,N_24114);
xnor UO_703 (O_703,N_24966,N_24159);
nand UO_704 (O_704,N_24469,N_24015);
xor UO_705 (O_705,N_24494,N_24762);
nand UO_706 (O_706,N_24674,N_24854);
xnor UO_707 (O_707,N_24510,N_24031);
or UO_708 (O_708,N_24983,N_24944);
nand UO_709 (O_709,N_24412,N_24900);
or UO_710 (O_710,N_24185,N_24083);
nor UO_711 (O_711,N_24042,N_24723);
and UO_712 (O_712,N_24408,N_24795);
and UO_713 (O_713,N_24566,N_24833);
nor UO_714 (O_714,N_24307,N_24234);
or UO_715 (O_715,N_24879,N_24771);
and UO_716 (O_716,N_24339,N_24179);
nor UO_717 (O_717,N_24144,N_24509);
or UO_718 (O_718,N_24736,N_24830);
nor UO_719 (O_719,N_24391,N_24071);
and UO_720 (O_720,N_24603,N_24174);
nand UO_721 (O_721,N_24273,N_24042);
or UO_722 (O_722,N_24917,N_24340);
or UO_723 (O_723,N_24720,N_24702);
nand UO_724 (O_724,N_24587,N_24639);
or UO_725 (O_725,N_24249,N_24145);
nor UO_726 (O_726,N_24439,N_24893);
and UO_727 (O_727,N_24740,N_24525);
or UO_728 (O_728,N_24202,N_24668);
nand UO_729 (O_729,N_24708,N_24336);
nand UO_730 (O_730,N_24875,N_24429);
or UO_731 (O_731,N_24517,N_24928);
xor UO_732 (O_732,N_24790,N_24571);
and UO_733 (O_733,N_24925,N_24689);
and UO_734 (O_734,N_24248,N_24729);
or UO_735 (O_735,N_24065,N_24158);
nand UO_736 (O_736,N_24231,N_24016);
nor UO_737 (O_737,N_24106,N_24884);
nand UO_738 (O_738,N_24232,N_24062);
xor UO_739 (O_739,N_24608,N_24870);
nor UO_740 (O_740,N_24585,N_24508);
nor UO_741 (O_741,N_24604,N_24865);
nand UO_742 (O_742,N_24398,N_24771);
and UO_743 (O_743,N_24993,N_24229);
nand UO_744 (O_744,N_24728,N_24953);
and UO_745 (O_745,N_24522,N_24750);
or UO_746 (O_746,N_24908,N_24588);
and UO_747 (O_747,N_24337,N_24325);
and UO_748 (O_748,N_24983,N_24592);
nor UO_749 (O_749,N_24974,N_24470);
or UO_750 (O_750,N_24750,N_24501);
and UO_751 (O_751,N_24912,N_24596);
or UO_752 (O_752,N_24567,N_24351);
and UO_753 (O_753,N_24137,N_24097);
or UO_754 (O_754,N_24305,N_24253);
nand UO_755 (O_755,N_24841,N_24526);
or UO_756 (O_756,N_24884,N_24869);
nor UO_757 (O_757,N_24383,N_24139);
nor UO_758 (O_758,N_24949,N_24917);
nor UO_759 (O_759,N_24247,N_24665);
or UO_760 (O_760,N_24119,N_24485);
nand UO_761 (O_761,N_24094,N_24866);
or UO_762 (O_762,N_24356,N_24861);
and UO_763 (O_763,N_24887,N_24566);
nor UO_764 (O_764,N_24799,N_24599);
nand UO_765 (O_765,N_24201,N_24076);
or UO_766 (O_766,N_24585,N_24309);
nand UO_767 (O_767,N_24202,N_24309);
xor UO_768 (O_768,N_24706,N_24886);
xor UO_769 (O_769,N_24328,N_24693);
and UO_770 (O_770,N_24245,N_24096);
xor UO_771 (O_771,N_24003,N_24956);
nor UO_772 (O_772,N_24103,N_24358);
nor UO_773 (O_773,N_24867,N_24908);
nor UO_774 (O_774,N_24485,N_24754);
xor UO_775 (O_775,N_24828,N_24903);
nand UO_776 (O_776,N_24127,N_24024);
and UO_777 (O_777,N_24203,N_24782);
nor UO_778 (O_778,N_24906,N_24045);
xor UO_779 (O_779,N_24406,N_24244);
xor UO_780 (O_780,N_24920,N_24469);
nor UO_781 (O_781,N_24194,N_24325);
nand UO_782 (O_782,N_24392,N_24136);
nand UO_783 (O_783,N_24911,N_24171);
nor UO_784 (O_784,N_24026,N_24139);
xor UO_785 (O_785,N_24396,N_24640);
or UO_786 (O_786,N_24992,N_24221);
nand UO_787 (O_787,N_24633,N_24593);
and UO_788 (O_788,N_24061,N_24249);
nand UO_789 (O_789,N_24856,N_24066);
nand UO_790 (O_790,N_24237,N_24106);
or UO_791 (O_791,N_24866,N_24760);
xnor UO_792 (O_792,N_24341,N_24346);
and UO_793 (O_793,N_24767,N_24511);
and UO_794 (O_794,N_24204,N_24217);
and UO_795 (O_795,N_24177,N_24051);
nand UO_796 (O_796,N_24991,N_24464);
or UO_797 (O_797,N_24467,N_24006);
xnor UO_798 (O_798,N_24400,N_24406);
or UO_799 (O_799,N_24941,N_24478);
and UO_800 (O_800,N_24156,N_24426);
xor UO_801 (O_801,N_24868,N_24603);
or UO_802 (O_802,N_24418,N_24334);
or UO_803 (O_803,N_24042,N_24096);
xor UO_804 (O_804,N_24261,N_24175);
nand UO_805 (O_805,N_24151,N_24856);
or UO_806 (O_806,N_24959,N_24679);
or UO_807 (O_807,N_24989,N_24157);
nand UO_808 (O_808,N_24455,N_24303);
xor UO_809 (O_809,N_24351,N_24198);
nand UO_810 (O_810,N_24354,N_24496);
or UO_811 (O_811,N_24975,N_24777);
and UO_812 (O_812,N_24281,N_24532);
nor UO_813 (O_813,N_24225,N_24744);
or UO_814 (O_814,N_24319,N_24592);
and UO_815 (O_815,N_24370,N_24907);
xor UO_816 (O_816,N_24494,N_24630);
xor UO_817 (O_817,N_24302,N_24523);
xnor UO_818 (O_818,N_24955,N_24623);
xnor UO_819 (O_819,N_24299,N_24190);
and UO_820 (O_820,N_24151,N_24658);
nor UO_821 (O_821,N_24276,N_24438);
xnor UO_822 (O_822,N_24099,N_24835);
nand UO_823 (O_823,N_24808,N_24496);
or UO_824 (O_824,N_24545,N_24123);
nor UO_825 (O_825,N_24132,N_24778);
xnor UO_826 (O_826,N_24921,N_24108);
xor UO_827 (O_827,N_24758,N_24948);
nor UO_828 (O_828,N_24698,N_24489);
and UO_829 (O_829,N_24078,N_24416);
xnor UO_830 (O_830,N_24084,N_24909);
and UO_831 (O_831,N_24566,N_24410);
or UO_832 (O_832,N_24521,N_24691);
nand UO_833 (O_833,N_24188,N_24878);
nand UO_834 (O_834,N_24634,N_24487);
nor UO_835 (O_835,N_24078,N_24442);
or UO_836 (O_836,N_24646,N_24091);
or UO_837 (O_837,N_24491,N_24804);
nor UO_838 (O_838,N_24048,N_24462);
nand UO_839 (O_839,N_24755,N_24905);
xnor UO_840 (O_840,N_24774,N_24881);
and UO_841 (O_841,N_24111,N_24236);
xnor UO_842 (O_842,N_24926,N_24459);
nor UO_843 (O_843,N_24573,N_24716);
nor UO_844 (O_844,N_24106,N_24731);
xor UO_845 (O_845,N_24660,N_24084);
or UO_846 (O_846,N_24539,N_24545);
and UO_847 (O_847,N_24844,N_24476);
and UO_848 (O_848,N_24746,N_24938);
xnor UO_849 (O_849,N_24509,N_24821);
nor UO_850 (O_850,N_24504,N_24847);
xnor UO_851 (O_851,N_24475,N_24403);
and UO_852 (O_852,N_24419,N_24516);
nor UO_853 (O_853,N_24057,N_24156);
xor UO_854 (O_854,N_24762,N_24085);
and UO_855 (O_855,N_24055,N_24455);
and UO_856 (O_856,N_24892,N_24273);
xnor UO_857 (O_857,N_24026,N_24683);
nand UO_858 (O_858,N_24992,N_24090);
nor UO_859 (O_859,N_24358,N_24269);
and UO_860 (O_860,N_24958,N_24336);
or UO_861 (O_861,N_24474,N_24599);
and UO_862 (O_862,N_24903,N_24303);
or UO_863 (O_863,N_24910,N_24486);
xnor UO_864 (O_864,N_24761,N_24924);
and UO_865 (O_865,N_24005,N_24304);
nand UO_866 (O_866,N_24568,N_24487);
nor UO_867 (O_867,N_24191,N_24007);
xnor UO_868 (O_868,N_24561,N_24784);
nor UO_869 (O_869,N_24288,N_24471);
or UO_870 (O_870,N_24314,N_24800);
and UO_871 (O_871,N_24676,N_24264);
nor UO_872 (O_872,N_24796,N_24337);
nor UO_873 (O_873,N_24203,N_24127);
and UO_874 (O_874,N_24896,N_24972);
and UO_875 (O_875,N_24222,N_24069);
nor UO_876 (O_876,N_24191,N_24974);
nand UO_877 (O_877,N_24530,N_24323);
nand UO_878 (O_878,N_24186,N_24236);
and UO_879 (O_879,N_24389,N_24229);
nand UO_880 (O_880,N_24514,N_24677);
nor UO_881 (O_881,N_24216,N_24828);
nor UO_882 (O_882,N_24548,N_24416);
nor UO_883 (O_883,N_24421,N_24911);
nand UO_884 (O_884,N_24375,N_24579);
nor UO_885 (O_885,N_24052,N_24819);
or UO_886 (O_886,N_24028,N_24232);
or UO_887 (O_887,N_24356,N_24789);
and UO_888 (O_888,N_24667,N_24211);
nand UO_889 (O_889,N_24739,N_24166);
nor UO_890 (O_890,N_24850,N_24813);
nor UO_891 (O_891,N_24748,N_24453);
or UO_892 (O_892,N_24224,N_24541);
nor UO_893 (O_893,N_24720,N_24345);
and UO_894 (O_894,N_24165,N_24724);
and UO_895 (O_895,N_24566,N_24985);
nor UO_896 (O_896,N_24228,N_24863);
xnor UO_897 (O_897,N_24059,N_24098);
nand UO_898 (O_898,N_24708,N_24678);
and UO_899 (O_899,N_24365,N_24126);
and UO_900 (O_900,N_24142,N_24256);
and UO_901 (O_901,N_24153,N_24971);
and UO_902 (O_902,N_24264,N_24535);
nor UO_903 (O_903,N_24111,N_24482);
or UO_904 (O_904,N_24415,N_24298);
or UO_905 (O_905,N_24522,N_24777);
or UO_906 (O_906,N_24903,N_24760);
or UO_907 (O_907,N_24074,N_24919);
and UO_908 (O_908,N_24572,N_24817);
nor UO_909 (O_909,N_24993,N_24705);
or UO_910 (O_910,N_24125,N_24062);
or UO_911 (O_911,N_24927,N_24224);
xnor UO_912 (O_912,N_24883,N_24136);
nor UO_913 (O_913,N_24021,N_24683);
and UO_914 (O_914,N_24237,N_24655);
xor UO_915 (O_915,N_24687,N_24733);
or UO_916 (O_916,N_24282,N_24907);
and UO_917 (O_917,N_24409,N_24848);
nor UO_918 (O_918,N_24869,N_24204);
and UO_919 (O_919,N_24380,N_24157);
and UO_920 (O_920,N_24463,N_24378);
nor UO_921 (O_921,N_24906,N_24405);
and UO_922 (O_922,N_24675,N_24991);
and UO_923 (O_923,N_24702,N_24894);
and UO_924 (O_924,N_24477,N_24482);
xnor UO_925 (O_925,N_24688,N_24941);
xor UO_926 (O_926,N_24409,N_24389);
nand UO_927 (O_927,N_24309,N_24276);
nand UO_928 (O_928,N_24159,N_24847);
xor UO_929 (O_929,N_24575,N_24009);
nor UO_930 (O_930,N_24932,N_24731);
or UO_931 (O_931,N_24032,N_24736);
or UO_932 (O_932,N_24967,N_24724);
or UO_933 (O_933,N_24232,N_24283);
or UO_934 (O_934,N_24230,N_24911);
xnor UO_935 (O_935,N_24147,N_24750);
or UO_936 (O_936,N_24363,N_24680);
nor UO_937 (O_937,N_24331,N_24008);
or UO_938 (O_938,N_24577,N_24897);
and UO_939 (O_939,N_24290,N_24342);
nand UO_940 (O_940,N_24027,N_24207);
and UO_941 (O_941,N_24583,N_24850);
xor UO_942 (O_942,N_24455,N_24222);
and UO_943 (O_943,N_24780,N_24814);
xor UO_944 (O_944,N_24676,N_24261);
or UO_945 (O_945,N_24774,N_24372);
xnor UO_946 (O_946,N_24415,N_24271);
nor UO_947 (O_947,N_24128,N_24775);
and UO_948 (O_948,N_24515,N_24719);
xor UO_949 (O_949,N_24737,N_24395);
and UO_950 (O_950,N_24530,N_24843);
and UO_951 (O_951,N_24971,N_24574);
nor UO_952 (O_952,N_24740,N_24881);
or UO_953 (O_953,N_24481,N_24745);
and UO_954 (O_954,N_24506,N_24577);
nor UO_955 (O_955,N_24641,N_24581);
nand UO_956 (O_956,N_24150,N_24797);
xnor UO_957 (O_957,N_24071,N_24898);
and UO_958 (O_958,N_24561,N_24530);
nor UO_959 (O_959,N_24363,N_24709);
nor UO_960 (O_960,N_24036,N_24171);
nor UO_961 (O_961,N_24618,N_24449);
nor UO_962 (O_962,N_24307,N_24456);
or UO_963 (O_963,N_24979,N_24784);
or UO_964 (O_964,N_24477,N_24051);
or UO_965 (O_965,N_24300,N_24091);
and UO_966 (O_966,N_24908,N_24142);
or UO_967 (O_967,N_24850,N_24799);
nand UO_968 (O_968,N_24376,N_24304);
xnor UO_969 (O_969,N_24813,N_24651);
and UO_970 (O_970,N_24665,N_24921);
nor UO_971 (O_971,N_24379,N_24940);
and UO_972 (O_972,N_24225,N_24882);
xnor UO_973 (O_973,N_24388,N_24653);
and UO_974 (O_974,N_24234,N_24364);
or UO_975 (O_975,N_24070,N_24435);
or UO_976 (O_976,N_24685,N_24189);
nor UO_977 (O_977,N_24575,N_24759);
and UO_978 (O_978,N_24632,N_24147);
and UO_979 (O_979,N_24438,N_24377);
nor UO_980 (O_980,N_24461,N_24495);
and UO_981 (O_981,N_24379,N_24825);
or UO_982 (O_982,N_24882,N_24425);
or UO_983 (O_983,N_24510,N_24537);
and UO_984 (O_984,N_24610,N_24270);
xnor UO_985 (O_985,N_24369,N_24849);
nor UO_986 (O_986,N_24180,N_24488);
nor UO_987 (O_987,N_24554,N_24472);
nor UO_988 (O_988,N_24612,N_24129);
nand UO_989 (O_989,N_24281,N_24801);
nand UO_990 (O_990,N_24553,N_24639);
or UO_991 (O_991,N_24983,N_24647);
nor UO_992 (O_992,N_24601,N_24753);
and UO_993 (O_993,N_24304,N_24979);
and UO_994 (O_994,N_24052,N_24572);
or UO_995 (O_995,N_24228,N_24358);
or UO_996 (O_996,N_24280,N_24579);
xor UO_997 (O_997,N_24950,N_24095);
and UO_998 (O_998,N_24156,N_24369);
and UO_999 (O_999,N_24990,N_24944);
or UO_1000 (O_1000,N_24983,N_24215);
nand UO_1001 (O_1001,N_24624,N_24051);
or UO_1002 (O_1002,N_24104,N_24281);
nand UO_1003 (O_1003,N_24650,N_24443);
nor UO_1004 (O_1004,N_24253,N_24458);
and UO_1005 (O_1005,N_24161,N_24342);
and UO_1006 (O_1006,N_24461,N_24360);
xnor UO_1007 (O_1007,N_24777,N_24786);
and UO_1008 (O_1008,N_24180,N_24726);
or UO_1009 (O_1009,N_24069,N_24716);
or UO_1010 (O_1010,N_24754,N_24727);
xnor UO_1011 (O_1011,N_24304,N_24271);
nand UO_1012 (O_1012,N_24939,N_24393);
nand UO_1013 (O_1013,N_24694,N_24610);
or UO_1014 (O_1014,N_24162,N_24932);
nor UO_1015 (O_1015,N_24187,N_24396);
or UO_1016 (O_1016,N_24327,N_24385);
xor UO_1017 (O_1017,N_24421,N_24668);
and UO_1018 (O_1018,N_24669,N_24352);
nor UO_1019 (O_1019,N_24520,N_24665);
or UO_1020 (O_1020,N_24503,N_24735);
or UO_1021 (O_1021,N_24555,N_24560);
and UO_1022 (O_1022,N_24785,N_24027);
and UO_1023 (O_1023,N_24865,N_24182);
and UO_1024 (O_1024,N_24918,N_24920);
and UO_1025 (O_1025,N_24460,N_24553);
xnor UO_1026 (O_1026,N_24309,N_24541);
nand UO_1027 (O_1027,N_24437,N_24845);
xnor UO_1028 (O_1028,N_24053,N_24153);
or UO_1029 (O_1029,N_24133,N_24791);
or UO_1030 (O_1030,N_24237,N_24635);
and UO_1031 (O_1031,N_24316,N_24188);
and UO_1032 (O_1032,N_24446,N_24605);
nand UO_1033 (O_1033,N_24292,N_24690);
nor UO_1034 (O_1034,N_24134,N_24995);
xnor UO_1035 (O_1035,N_24302,N_24698);
xnor UO_1036 (O_1036,N_24104,N_24017);
nor UO_1037 (O_1037,N_24156,N_24566);
nand UO_1038 (O_1038,N_24128,N_24057);
nor UO_1039 (O_1039,N_24986,N_24761);
nand UO_1040 (O_1040,N_24282,N_24048);
nand UO_1041 (O_1041,N_24733,N_24780);
nor UO_1042 (O_1042,N_24189,N_24002);
nor UO_1043 (O_1043,N_24388,N_24568);
nand UO_1044 (O_1044,N_24945,N_24688);
xor UO_1045 (O_1045,N_24567,N_24811);
xnor UO_1046 (O_1046,N_24893,N_24494);
xnor UO_1047 (O_1047,N_24733,N_24537);
xnor UO_1048 (O_1048,N_24408,N_24543);
xor UO_1049 (O_1049,N_24855,N_24956);
xnor UO_1050 (O_1050,N_24226,N_24758);
nor UO_1051 (O_1051,N_24299,N_24568);
xnor UO_1052 (O_1052,N_24140,N_24536);
xor UO_1053 (O_1053,N_24598,N_24030);
nor UO_1054 (O_1054,N_24844,N_24893);
and UO_1055 (O_1055,N_24506,N_24650);
nand UO_1056 (O_1056,N_24791,N_24532);
and UO_1057 (O_1057,N_24750,N_24082);
xor UO_1058 (O_1058,N_24461,N_24386);
and UO_1059 (O_1059,N_24940,N_24226);
and UO_1060 (O_1060,N_24953,N_24262);
xor UO_1061 (O_1061,N_24688,N_24056);
nand UO_1062 (O_1062,N_24217,N_24913);
xor UO_1063 (O_1063,N_24068,N_24300);
nand UO_1064 (O_1064,N_24420,N_24859);
nand UO_1065 (O_1065,N_24277,N_24115);
xnor UO_1066 (O_1066,N_24592,N_24839);
nor UO_1067 (O_1067,N_24552,N_24397);
nand UO_1068 (O_1068,N_24442,N_24045);
xnor UO_1069 (O_1069,N_24300,N_24174);
nor UO_1070 (O_1070,N_24052,N_24755);
xor UO_1071 (O_1071,N_24859,N_24062);
or UO_1072 (O_1072,N_24182,N_24605);
xnor UO_1073 (O_1073,N_24941,N_24024);
nand UO_1074 (O_1074,N_24683,N_24979);
xnor UO_1075 (O_1075,N_24528,N_24194);
xnor UO_1076 (O_1076,N_24832,N_24849);
and UO_1077 (O_1077,N_24218,N_24478);
or UO_1078 (O_1078,N_24609,N_24601);
nand UO_1079 (O_1079,N_24344,N_24608);
or UO_1080 (O_1080,N_24454,N_24393);
xnor UO_1081 (O_1081,N_24710,N_24511);
nor UO_1082 (O_1082,N_24591,N_24249);
and UO_1083 (O_1083,N_24985,N_24650);
nor UO_1084 (O_1084,N_24194,N_24474);
nand UO_1085 (O_1085,N_24357,N_24870);
nand UO_1086 (O_1086,N_24873,N_24964);
and UO_1087 (O_1087,N_24989,N_24843);
or UO_1088 (O_1088,N_24516,N_24858);
and UO_1089 (O_1089,N_24985,N_24407);
xnor UO_1090 (O_1090,N_24108,N_24167);
nand UO_1091 (O_1091,N_24052,N_24126);
and UO_1092 (O_1092,N_24774,N_24412);
or UO_1093 (O_1093,N_24784,N_24169);
nand UO_1094 (O_1094,N_24516,N_24079);
or UO_1095 (O_1095,N_24559,N_24729);
xnor UO_1096 (O_1096,N_24348,N_24401);
and UO_1097 (O_1097,N_24294,N_24211);
xnor UO_1098 (O_1098,N_24130,N_24343);
nand UO_1099 (O_1099,N_24827,N_24322);
nand UO_1100 (O_1100,N_24880,N_24650);
and UO_1101 (O_1101,N_24895,N_24684);
and UO_1102 (O_1102,N_24612,N_24618);
nand UO_1103 (O_1103,N_24978,N_24733);
xnor UO_1104 (O_1104,N_24286,N_24153);
and UO_1105 (O_1105,N_24390,N_24739);
xnor UO_1106 (O_1106,N_24970,N_24056);
nand UO_1107 (O_1107,N_24420,N_24943);
nand UO_1108 (O_1108,N_24543,N_24446);
xnor UO_1109 (O_1109,N_24613,N_24939);
and UO_1110 (O_1110,N_24059,N_24698);
xor UO_1111 (O_1111,N_24991,N_24447);
nand UO_1112 (O_1112,N_24807,N_24096);
or UO_1113 (O_1113,N_24457,N_24256);
nor UO_1114 (O_1114,N_24793,N_24250);
and UO_1115 (O_1115,N_24559,N_24826);
and UO_1116 (O_1116,N_24278,N_24497);
and UO_1117 (O_1117,N_24776,N_24978);
xor UO_1118 (O_1118,N_24773,N_24279);
nor UO_1119 (O_1119,N_24363,N_24940);
nand UO_1120 (O_1120,N_24498,N_24713);
nand UO_1121 (O_1121,N_24655,N_24300);
and UO_1122 (O_1122,N_24679,N_24191);
and UO_1123 (O_1123,N_24370,N_24124);
or UO_1124 (O_1124,N_24496,N_24152);
and UO_1125 (O_1125,N_24600,N_24575);
nand UO_1126 (O_1126,N_24377,N_24810);
or UO_1127 (O_1127,N_24915,N_24619);
nand UO_1128 (O_1128,N_24276,N_24025);
nand UO_1129 (O_1129,N_24847,N_24799);
nor UO_1130 (O_1130,N_24461,N_24637);
or UO_1131 (O_1131,N_24466,N_24106);
nand UO_1132 (O_1132,N_24779,N_24332);
nand UO_1133 (O_1133,N_24793,N_24200);
or UO_1134 (O_1134,N_24686,N_24889);
nor UO_1135 (O_1135,N_24099,N_24914);
xnor UO_1136 (O_1136,N_24092,N_24897);
xnor UO_1137 (O_1137,N_24294,N_24365);
and UO_1138 (O_1138,N_24043,N_24186);
nand UO_1139 (O_1139,N_24297,N_24108);
nor UO_1140 (O_1140,N_24658,N_24394);
and UO_1141 (O_1141,N_24677,N_24374);
xnor UO_1142 (O_1142,N_24387,N_24193);
or UO_1143 (O_1143,N_24269,N_24488);
or UO_1144 (O_1144,N_24192,N_24960);
nor UO_1145 (O_1145,N_24206,N_24216);
nor UO_1146 (O_1146,N_24939,N_24900);
nor UO_1147 (O_1147,N_24224,N_24493);
and UO_1148 (O_1148,N_24780,N_24386);
or UO_1149 (O_1149,N_24528,N_24931);
and UO_1150 (O_1150,N_24305,N_24596);
nand UO_1151 (O_1151,N_24428,N_24890);
and UO_1152 (O_1152,N_24846,N_24416);
xnor UO_1153 (O_1153,N_24234,N_24989);
xor UO_1154 (O_1154,N_24337,N_24740);
nand UO_1155 (O_1155,N_24036,N_24363);
nor UO_1156 (O_1156,N_24349,N_24761);
nor UO_1157 (O_1157,N_24902,N_24607);
nor UO_1158 (O_1158,N_24595,N_24582);
nand UO_1159 (O_1159,N_24382,N_24522);
or UO_1160 (O_1160,N_24213,N_24393);
nor UO_1161 (O_1161,N_24519,N_24511);
or UO_1162 (O_1162,N_24611,N_24501);
or UO_1163 (O_1163,N_24047,N_24692);
nand UO_1164 (O_1164,N_24519,N_24014);
nor UO_1165 (O_1165,N_24425,N_24839);
xor UO_1166 (O_1166,N_24290,N_24569);
and UO_1167 (O_1167,N_24717,N_24162);
or UO_1168 (O_1168,N_24811,N_24027);
nor UO_1169 (O_1169,N_24933,N_24093);
or UO_1170 (O_1170,N_24044,N_24587);
and UO_1171 (O_1171,N_24782,N_24515);
nand UO_1172 (O_1172,N_24999,N_24606);
nand UO_1173 (O_1173,N_24173,N_24315);
nand UO_1174 (O_1174,N_24359,N_24062);
nand UO_1175 (O_1175,N_24398,N_24705);
xnor UO_1176 (O_1176,N_24018,N_24637);
nor UO_1177 (O_1177,N_24649,N_24371);
nor UO_1178 (O_1178,N_24861,N_24469);
or UO_1179 (O_1179,N_24394,N_24075);
or UO_1180 (O_1180,N_24375,N_24856);
and UO_1181 (O_1181,N_24338,N_24077);
and UO_1182 (O_1182,N_24280,N_24216);
nand UO_1183 (O_1183,N_24405,N_24710);
and UO_1184 (O_1184,N_24240,N_24008);
nor UO_1185 (O_1185,N_24647,N_24785);
nand UO_1186 (O_1186,N_24258,N_24537);
nor UO_1187 (O_1187,N_24739,N_24695);
xor UO_1188 (O_1188,N_24652,N_24318);
or UO_1189 (O_1189,N_24536,N_24301);
or UO_1190 (O_1190,N_24542,N_24439);
nor UO_1191 (O_1191,N_24797,N_24428);
or UO_1192 (O_1192,N_24966,N_24068);
or UO_1193 (O_1193,N_24473,N_24963);
xnor UO_1194 (O_1194,N_24532,N_24833);
nor UO_1195 (O_1195,N_24351,N_24129);
nand UO_1196 (O_1196,N_24110,N_24260);
nand UO_1197 (O_1197,N_24446,N_24137);
or UO_1198 (O_1198,N_24247,N_24575);
and UO_1199 (O_1199,N_24069,N_24715);
and UO_1200 (O_1200,N_24501,N_24978);
xnor UO_1201 (O_1201,N_24987,N_24752);
and UO_1202 (O_1202,N_24231,N_24837);
or UO_1203 (O_1203,N_24789,N_24835);
and UO_1204 (O_1204,N_24890,N_24256);
nand UO_1205 (O_1205,N_24825,N_24218);
xnor UO_1206 (O_1206,N_24778,N_24273);
xor UO_1207 (O_1207,N_24840,N_24071);
and UO_1208 (O_1208,N_24211,N_24913);
nor UO_1209 (O_1209,N_24207,N_24014);
and UO_1210 (O_1210,N_24559,N_24366);
nor UO_1211 (O_1211,N_24642,N_24127);
and UO_1212 (O_1212,N_24304,N_24174);
xor UO_1213 (O_1213,N_24108,N_24242);
or UO_1214 (O_1214,N_24904,N_24878);
nand UO_1215 (O_1215,N_24135,N_24342);
xor UO_1216 (O_1216,N_24559,N_24289);
xnor UO_1217 (O_1217,N_24411,N_24734);
xor UO_1218 (O_1218,N_24362,N_24541);
xnor UO_1219 (O_1219,N_24771,N_24593);
and UO_1220 (O_1220,N_24563,N_24771);
nor UO_1221 (O_1221,N_24792,N_24111);
or UO_1222 (O_1222,N_24998,N_24764);
or UO_1223 (O_1223,N_24338,N_24632);
or UO_1224 (O_1224,N_24927,N_24467);
xor UO_1225 (O_1225,N_24717,N_24464);
or UO_1226 (O_1226,N_24155,N_24689);
xnor UO_1227 (O_1227,N_24752,N_24377);
and UO_1228 (O_1228,N_24302,N_24914);
or UO_1229 (O_1229,N_24838,N_24320);
xnor UO_1230 (O_1230,N_24006,N_24830);
nor UO_1231 (O_1231,N_24449,N_24258);
nor UO_1232 (O_1232,N_24136,N_24970);
or UO_1233 (O_1233,N_24470,N_24965);
nand UO_1234 (O_1234,N_24549,N_24313);
nand UO_1235 (O_1235,N_24859,N_24535);
nor UO_1236 (O_1236,N_24671,N_24625);
nand UO_1237 (O_1237,N_24878,N_24427);
xor UO_1238 (O_1238,N_24402,N_24575);
or UO_1239 (O_1239,N_24722,N_24457);
nand UO_1240 (O_1240,N_24137,N_24048);
and UO_1241 (O_1241,N_24343,N_24346);
xnor UO_1242 (O_1242,N_24076,N_24336);
nand UO_1243 (O_1243,N_24793,N_24013);
xnor UO_1244 (O_1244,N_24723,N_24875);
and UO_1245 (O_1245,N_24066,N_24891);
xnor UO_1246 (O_1246,N_24491,N_24266);
and UO_1247 (O_1247,N_24891,N_24909);
and UO_1248 (O_1248,N_24790,N_24872);
and UO_1249 (O_1249,N_24496,N_24124);
xor UO_1250 (O_1250,N_24851,N_24493);
nand UO_1251 (O_1251,N_24461,N_24889);
xor UO_1252 (O_1252,N_24884,N_24493);
and UO_1253 (O_1253,N_24573,N_24519);
or UO_1254 (O_1254,N_24828,N_24063);
or UO_1255 (O_1255,N_24955,N_24070);
xor UO_1256 (O_1256,N_24649,N_24625);
or UO_1257 (O_1257,N_24231,N_24527);
nor UO_1258 (O_1258,N_24411,N_24024);
or UO_1259 (O_1259,N_24099,N_24482);
nand UO_1260 (O_1260,N_24047,N_24396);
and UO_1261 (O_1261,N_24115,N_24308);
nor UO_1262 (O_1262,N_24199,N_24957);
nor UO_1263 (O_1263,N_24109,N_24851);
nand UO_1264 (O_1264,N_24348,N_24213);
or UO_1265 (O_1265,N_24004,N_24258);
nand UO_1266 (O_1266,N_24294,N_24861);
and UO_1267 (O_1267,N_24179,N_24101);
nand UO_1268 (O_1268,N_24131,N_24911);
xor UO_1269 (O_1269,N_24086,N_24792);
or UO_1270 (O_1270,N_24655,N_24752);
or UO_1271 (O_1271,N_24318,N_24912);
and UO_1272 (O_1272,N_24880,N_24948);
and UO_1273 (O_1273,N_24534,N_24450);
and UO_1274 (O_1274,N_24530,N_24023);
and UO_1275 (O_1275,N_24765,N_24629);
xnor UO_1276 (O_1276,N_24573,N_24999);
or UO_1277 (O_1277,N_24873,N_24475);
nor UO_1278 (O_1278,N_24214,N_24773);
nor UO_1279 (O_1279,N_24933,N_24331);
nor UO_1280 (O_1280,N_24059,N_24271);
and UO_1281 (O_1281,N_24895,N_24251);
or UO_1282 (O_1282,N_24156,N_24554);
nand UO_1283 (O_1283,N_24464,N_24465);
or UO_1284 (O_1284,N_24975,N_24765);
nor UO_1285 (O_1285,N_24510,N_24151);
nand UO_1286 (O_1286,N_24452,N_24973);
nor UO_1287 (O_1287,N_24648,N_24852);
nand UO_1288 (O_1288,N_24591,N_24212);
nor UO_1289 (O_1289,N_24672,N_24996);
or UO_1290 (O_1290,N_24074,N_24025);
xor UO_1291 (O_1291,N_24178,N_24808);
xor UO_1292 (O_1292,N_24908,N_24368);
and UO_1293 (O_1293,N_24401,N_24639);
nand UO_1294 (O_1294,N_24348,N_24404);
xnor UO_1295 (O_1295,N_24405,N_24697);
and UO_1296 (O_1296,N_24142,N_24928);
nor UO_1297 (O_1297,N_24603,N_24797);
and UO_1298 (O_1298,N_24206,N_24410);
xnor UO_1299 (O_1299,N_24236,N_24395);
xnor UO_1300 (O_1300,N_24854,N_24982);
nor UO_1301 (O_1301,N_24156,N_24495);
and UO_1302 (O_1302,N_24565,N_24560);
nor UO_1303 (O_1303,N_24852,N_24485);
or UO_1304 (O_1304,N_24442,N_24999);
xor UO_1305 (O_1305,N_24017,N_24576);
nor UO_1306 (O_1306,N_24833,N_24414);
and UO_1307 (O_1307,N_24814,N_24829);
or UO_1308 (O_1308,N_24785,N_24835);
or UO_1309 (O_1309,N_24372,N_24033);
xor UO_1310 (O_1310,N_24807,N_24932);
or UO_1311 (O_1311,N_24615,N_24342);
and UO_1312 (O_1312,N_24372,N_24132);
xor UO_1313 (O_1313,N_24217,N_24807);
nand UO_1314 (O_1314,N_24818,N_24810);
nor UO_1315 (O_1315,N_24530,N_24691);
xnor UO_1316 (O_1316,N_24490,N_24803);
and UO_1317 (O_1317,N_24713,N_24081);
or UO_1318 (O_1318,N_24267,N_24260);
nand UO_1319 (O_1319,N_24140,N_24937);
or UO_1320 (O_1320,N_24263,N_24615);
xnor UO_1321 (O_1321,N_24360,N_24482);
nand UO_1322 (O_1322,N_24814,N_24403);
nor UO_1323 (O_1323,N_24673,N_24470);
or UO_1324 (O_1324,N_24858,N_24324);
nand UO_1325 (O_1325,N_24973,N_24750);
xor UO_1326 (O_1326,N_24994,N_24684);
and UO_1327 (O_1327,N_24720,N_24667);
nor UO_1328 (O_1328,N_24223,N_24961);
xnor UO_1329 (O_1329,N_24538,N_24561);
and UO_1330 (O_1330,N_24960,N_24293);
xnor UO_1331 (O_1331,N_24046,N_24277);
xnor UO_1332 (O_1332,N_24887,N_24234);
or UO_1333 (O_1333,N_24790,N_24596);
xor UO_1334 (O_1334,N_24683,N_24524);
and UO_1335 (O_1335,N_24891,N_24566);
nand UO_1336 (O_1336,N_24027,N_24294);
and UO_1337 (O_1337,N_24684,N_24495);
xor UO_1338 (O_1338,N_24880,N_24233);
or UO_1339 (O_1339,N_24020,N_24873);
xnor UO_1340 (O_1340,N_24360,N_24203);
and UO_1341 (O_1341,N_24892,N_24332);
xnor UO_1342 (O_1342,N_24742,N_24386);
nor UO_1343 (O_1343,N_24881,N_24382);
nor UO_1344 (O_1344,N_24790,N_24945);
nand UO_1345 (O_1345,N_24634,N_24650);
nor UO_1346 (O_1346,N_24432,N_24558);
xor UO_1347 (O_1347,N_24342,N_24702);
nor UO_1348 (O_1348,N_24202,N_24756);
and UO_1349 (O_1349,N_24721,N_24404);
and UO_1350 (O_1350,N_24969,N_24383);
xor UO_1351 (O_1351,N_24925,N_24882);
nand UO_1352 (O_1352,N_24616,N_24418);
xnor UO_1353 (O_1353,N_24917,N_24231);
xor UO_1354 (O_1354,N_24770,N_24685);
xor UO_1355 (O_1355,N_24618,N_24759);
xor UO_1356 (O_1356,N_24719,N_24605);
nor UO_1357 (O_1357,N_24536,N_24585);
nor UO_1358 (O_1358,N_24668,N_24390);
nor UO_1359 (O_1359,N_24733,N_24388);
xnor UO_1360 (O_1360,N_24093,N_24555);
xnor UO_1361 (O_1361,N_24777,N_24366);
and UO_1362 (O_1362,N_24444,N_24601);
xor UO_1363 (O_1363,N_24865,N_24370);
or UO_1364 (O_1364,N_24956,N_24473);
and UO_1365 (O_1365,N_24467,N_24509);
and UO_1366 (O_1366,N_24170,N_24470);
nand UO_1367 (O_1367,N_24978,N_24251);
and UO_1368 (O_1368,N_24685,N_24398);
and UO_1369 (O_1369,N_24584,N_24746);
or UO_1370 (O_1370,N_24960,N_24265);
nor UO_1371 (O_1371,N_24496,N_24957);
and UO_1372 (O_1372,N_24770,N_24730);
nor UO_1373 (O_1373,N_24053,N_24210);
nor UO_1374 (O_1374,N_24124,N_24952);
or UO_1375 (O_1375,N_24758,N_24189);
nand UO_1376 (O_1376,N_24811,N_24343);
nor UO_1377 (O_1377,N_24258,N_24329);
nand UO_1378 (O_1378,N_24590,N_24441);
and UO_1379 (O_1379,N_24878,N_24539);
nor UO_1380 (O_1380,N_24780,N_24083);
or UO_1381 (O_1381,N_24750,N_24770);
nor UO_1382 (O_1382,N_24427,N_24681);
xor UO_1383 (O_1383,N_24806,N_24312);
nor UO_1384 (O_1384,N_24871,N_24851);
nor UO_1385 (O_1385,N_24723,N_24294);
or UO_1386 (O_1386,N_24433,N_24842);
nor UO_1387 (O_1387,N_24799,N_24459);
and UO_1388 (O_1388,N_24990,N_24537);
and UO_1389 (O_1389,N_24517,N_24349);
nand UO_1390 (O_1390,N_24103,N_24725);
and UO_1391 (O_1391,N_24935,N_24018);
or UO_1392 (O_1392,N_24321,N_24841);
and UO_1393 (O_1393,N_24767,N_24405);
or UO_1394 (O_1394,N_24317,N_24363);
xor UO_1395 (O_1395,N_24358,N_24512);
xor UO_1396 (O_1396,N_24475,N_24363);
nor UO_1397 (O_1397,N_24296,N_24334);
xor UO_1398 (O_1398,N_24383,N_24055);
nor UO_1399 (O_1399,N_24298,N_24126);
or UO_1400 (O_1400,N_24725,N_24732);
nand UO_1401 (O_1401,N_24658,N_24375);
and UO_1402 (O_1402,N_24767,N_24741);
nor UO_1403 (O_1403,N_24144,N_24309);
nor UO_1404 (O_1404,N_24121,N_24878);
xor UO_1405 (O_1405,N_24851,N_24870);
and UO_1406 (O_1406,N_24634,N_24852);
nand UO_1407 (O_1407,N_24909,N_24415);
nand UO_1408 (O_1408,N_24287,N_24715);
nand UO_1409 (O_1409,N_24097,N_24777);
and UO_1410 (O_1410,N_24481,N_24268);
nor UO_1411 (O_1411,N_24228,N_24295);
nor UO_1412 (O_1412,N_24727,N_24189);
nand UO_1413 (O_1413,N_24404,N_24909);
nor UO_1414 (O_1414,N_24476,N_24932);
and UO_1415 (O_1415,N_24762,N_24235);
nor UO_1416 (O_1416,N_24933,N_24358);
nand UO_1417 (O_1417,N_24478,N_24513);
xnor UO_1418 (O_1418,N_24973,N_24712);
xnor UO_1419 (O_1419,N_24356,N_24824);
and UO_1420 (O_1420,N_24817,N_24443);
or UO_1421 (O_1421,N_24168,N_24298);
xnor UO_1422 (O_1422,N_24691,N_24548);
or UO_1423 (O_1423,N_24436,N_24594);
xnor UO_1424 (O_1424,N_24202,N_24721);
or UO_1425 (O_1425,N_24340,N_24075);
or UO_1426 (O_1426,N_24297,N_24267);
xor UO_1427 (O_1427,N_24627,N_24158);
nor UO_1428 (O_1428,N_24485,N_24283);
nand UO_1429 (O_1429,N_24601,N_24141);
nand UO_1430 (O_1430,N_24126,N_24137);
nand UO_1431 (O_1431,N_24344,N_24311);
and UO_1432 (O_1432,N_24632,N_24656);
nand UO_1433 (O_1433,N_24629,N_24300);
xor UO_1434 (O_1434,N_24722,N_24493);
nor UO_1435 (O_1435,N_24419,N_24128);
xnor UO_1436 (O_1436,N_24129,N_24223);
or UO_1437 (O_1437,N_24036,N_24577);
nor UO_1438 (O_1438,N_24170,N_24967);
nand UO_1439 (O_1439,N_24466,N_24974);
or UO_1440 (O_1440,N_24739,N_24598);
or UO_1441 (O_1441,N_24178,N_24105);
xnor UO_1442 (O_1442,N_24792,N_24347);
or UO_1443 (O_1443,N_24947,N_24759);
xnor UO_1444 (O_1444,N_24431,N_24559);
nor UO_1445 (O_1445,N_24138,N_24612);
nor UO_1446 (O_1446,N_24562,N_24695);
nor UO_1447 (O_1447,N_24326,N_24104);
xnor UO_1448 (O_1448,N_24059,N_24269);
nor UO_1449 (O_1449,N_24795,N_24763);
nand UO_1450 (O_1450,N_24830,N_24364);
nand UO_1451 (O_1451,N_24161,N_24406);
and UO_1452 (O_1452,N_24398,N_24521);
nor UO_1453 (O_1453,N_24748,N_24072);
xnor UO_1454 (O_1454,N_24730,N_24184);
and UO_1455 (O_1455,N_24359,N_24690);
xor UO_1456 (O_1456,N_24462,N_24472);
or UO_1457 (O_1457,N_24316,N_24373);
and UO_1458 (O_1458,N_24873,N_24444);
xor UO_1459 (O_1459,N_24058,N_24772);
nand UO_1460 (O_1460,N_24243,N_24817);
nand UO_1461 (O_1461,N_24134,N_24677);
and UO_1462 (O_1462,N_24172,N_24772);
and UO_1463 (O_1463,N_24887,N_24997);
xor UO_1464 (O_1464,N_24356,N_24448);
nand UO_1465 (O_1465,N_24273,N_24953);
nor UO_1466 (O_1466,N_24362,N_24754);
nand UO_1467 (O_1467,N_24458,N_24501);
nand UO_1468 (O_1468,N_24760,N_24973);
and UO_1469 (O_1469,N_24296,N_24778);
and UO_1470 (O_1470,N_24721,N_24582);
or UO_1471 (O_1471,N_24361,N_24199);
xor UO_1472 (O_1472,N_24944,N_24830);
nand UO_1473 (O_1473,N_24251,N_24160);
xor UO_1474 (O_1474,N_24809,N_24515);
xnor UO_1475 (O_1475,N_24808,N_24376);
xnor UO_1476 (O_1476,N_24957,N_24232);
and UO_1477 (O_1477,N_24784,N_24393);
nor UO_1478 (O_1478,N_24982,N_24445);
nor UO_1479 (O_1479,N_24643,N_24838);
xnor UO_1480 (O_1480,N_24748,N_24942);
nor UO_1481 (O_1481,N_24437,N_24579);
and UO_1482 (O_1482,N_24261,N_24084);
or UO_1483 (O_1483,N_24592,N_24910);
xnor UO_1484 (O_1484,N_24794,N_24497);
and UO_1485 (O_1485,N_24556,N_24894);
or UO_1486 (O_1486,N_24752,N_24081);
xnor UO_1487 (O_1487,N_24923,N_24527);
xor UO_1488 (O_1488,N_24416,N_24483);
or UO_1489 (O_1489,N_24069,N_24327);
nand UO_1490 (O_1490,N_24183,N_24400);
xor UO_1491 (O_1491,N_24421,N_24284);
or UO_1492 (O_1492,N_24352,N_24017);
xor UO_1493 (O_1493,N_24793,N_24565);
nand UO_1494 (O_1494,N_24532,N_24445);
or UO_1495 (O_1495,N_24357,N_24094);
nand UO_1496 (O_1496,N_24939,N_24596);
xnor UO_1497 (O_1497,N_24507,N_24222);
xor UO_1498 (O_1498,N_24742,N_24716);
and UO_1499 (O_1499,N_24302,N_24894);
xor UO_1500 (O_1500,N_24066,N_24556);
xor UO_1501 (O_1501,N_24719,N_24813);
nor UO_1502 (O_1502,N_24630,N_24126);
xor UO_1503 (O_1503,N_24154,N_24877);
and UO_1504 (O_1504,N_24086,N_24216);
nand UO_1505 (O_1505,N_24682,N_24919);
nand UO_1506 (O_1506,N_24977,N_24805);
nand UO_1507 (O_1507,N_24491,N_24236);
or UO_1508 (O_1508,N_24490,N_24265);
and UO_1509 (O_1509,N_24155,N_24350);
or UO_1510 (O_1510,N_24708,N_24168);
xnor UO_1511 (O_1511,N_24925,N_24908);
and UO_1512 (O_1512,N_24838,N_24654);
and UO_1513 (O_1513,N_24518,N_24207);
nor UO_1514 (O_1514,N_24082,N_24574);
xor UO_1515 (O_1515,N_24864,N_24878);
nor UO_1516 (O_1516,N_24241,N_24824);
or UO_1517 (O_1517,N_24754,N_24181);
or UO_1518 (O_1518,N_24405,N_24063);
nor UO_1519 (O_1519,N_24862,N_24035);
nand UO_1520 (O_1520,N_24025,N_24591);
and UO_1521 (O_1521,N_24222,N_24798);
nor UO_1522 (O_1522,N_24044,N_24225);
nand UO_1523 (O_1523,N_24796,N_24817);
or UO_1524 (O_1524,N_24336,N_24086);
or UO_1525 (O_1525,N_24524,N_24811);
or UO_1526 (O_1526,N_24790,N_24913);
nor UO_1527 (O_1527,N_24639,N_24340);
nand UO_1528 (O_1528,N_24489,N_24353);
or UO_1529 (O_1529,N_24710,N_24107);
and UO_1530 (O_1530,N_24108,N_24442);
nor UO_1531 (O_1531,N_24754,N_24349);
or UO_1532 (O_1532,N_24880,N_24304);
and UO_1533 (O_1533,N_24108,N_24922);
or UO_1534 (O_1534,N_24074,N_24911);
nand UO_1535 (O_1535,N_24257,N_24642);
and UO_1536 (O_1536,N_24573,N_24096);
xnor UO_1537 (O_1537,N_24361,N_24115);
or UO_1538 (O_1538,N_24209,N_24067);
xor UO_1539 (O_1539,N_24940,N_24182);
xnor UO_1540 (O_1540,N_24139,N_24572);
xor UO_1541 (O_1541,N_24247,N_24760);
and UO_1542 (O_1542,N_24606,N_24100);
or UO_1543 (O_1543,N_24608,N_24610);
nor UO_1544 (O_1544,N_24326,N_24952);
nor UO_1545 (O_1545,N_24509,N_24525);
xor UO_1546 (O_1546,N_24521,N_24423);
nand UO_1547 (O_1547,N_24288,N_24858);
nand UO_1548 (O_1548,N_24004,N_24494);
or UO_1549 (O_1549,N_24990,N_24380);
and UO_1550 (O_1550,N_24163,N_24627);
or UO_1551 (O_1551,N_24927,N_24569);
xnor UO_1552 (O_1552,N_24321,N_24473);
or UO_1553 (O_1553,N_24792,N_24198);
xor UO_1554 (O_1554,N_24153,N_24984);
or UO_1555 (O_1555,N_24522,N_24441);
or UO_1556 (O_1556,N_24924,N_24753);
or UO_1557 (O_1557,N_24457,N_24228);
and UO_1558 (O_1558,N_24642,N_24586);
or UO_1559 (O_1559,N_24951,N_24264);
or UO_1560 (O_1560,N_24732,N_24059);
nand UO_1561 (O_1561,N_24937,N_24698);
xor UO_1562 (O_1562,N_24216,N_24373);
nand UO_1563 (O_1563,N_24832,N_24996);
nor UO_1564 (O_1564,N_24416,N_24736);
nand UO_1565 (O_1565,N_24740,N_24186);
nand UO_1566 (O_1566,N_24315,N_24532);
and UO_1567 (O_1567,N_24013,N_24373);
and UO_1568 (O_1568,N_24383,N_24590);
nand UO_1569 (O_1569,N_24466,N_24057);
nor UO_1570 (O_1570,N_24678,N_24627);
nand UO_1571 (O_1571,N_24412,N_24060);
or UO_1572 (O_1572,N_24939,N_24369);
nand UO_1573 (O_1573,N_24466,N_24989);
nor UO_1574 (O_1574,N_24117,N_24199);
nand UO_1575 (O_1575,N_24665,N_24470);
nor UO_1576 (O_1576,N_24590,N_24328);
nand UO_1577 (O_1577,N_24891,N_24097);
nand UO_1578 (O_1578,N_24258,N_24103);
xor UO_1579 (O_1579,N_24930,N_24271);
xor UO_1580 (O_1580,N_24567,N_24718);
nor UO_1581 (O_1581,N_24956,N_24234);
and UO_1582 (O_1582,N_24886,N_24887);
nor UO_1583 (O_1583,N_24005,N_24793);
or UO_1584 (O_1584,N_24283,N_24291);
nor UO_1585 (O_1585,N_24390,N_24136);
nor UO_1586 (O_1586,N_24728,N_24661);
and UO_1587 (O_1587,N_24339,N_24072);
and UO_1588 (O_1588,N_24902,N_24891);
xor UO_1589 (O_1589,N_24414,N_24417);
and UO_1590 (O_1590,N_24322,N_24926);
xor UO_1591 (O_1591,N_24465,N_24495);
nand UO_1592 (O_1592,N_24223,N_24768);
and UO_1593 (O_1593,N_24909,N_24899);
nand UO_1594 (O_1594,N_24047,N_24483);
xnor UO_1595 (O_1595,N_24440,N_24466);
nor UO_1596 (O_1596,N_24648,N_24416);
or UO_1597 (O_1597,N_24344,N_24546);
xnor UO_1598 (O_1598,N_24668,N_24245);
nor UO_1599 (O_1599,N_24805,N_24698);
or UO_1600 (O_1600,N_24790,N_24590);
xor UO_1601 (O_1601,N_24147,N_24530);
nand UO_1602 (O_1602,N_24270,N_24441);
nand UO_1603 (O_1603,N_24612,N_24769);
or UO_1604 (O_1604,N_24022,N_24622);
xor UO_1605 (O_1605,N_24071,N_24543);
nor UO_1606 (O_1606,N_24451,N_24281);
and UO_1607 (O_1607,N_24291,N_24357);
and UO_1608 (O_1608,N_24949,N_24760);
and UO_1609 (O_1609,N_24779,N_24794);
or UO_1610 (O_1610,N_24600,N_24499);
nor UO_1611 (O_1611,N_24826,N_24528);
or UO_1612 (O_1612,N_24545,N_24437);
xnor UO_1613 (O_1613,N_24696,N_24331);
or UO_1614 (O_1614,N_24322,N_24250);
or UO_1615 (O_1615,N_24902,N_24665);
nor UO_1616 (O_1616,N_24996,N_24539);
and UO_1617 (O_1617,N_24860,N_24003);
and UO_1618 (O_1618,N_24700,N_24343);
nand UO_1619 (O_1619,N_24658,N_24484);
and UO_1620 (O_1620,N_24477,N_24008);
or UO_1621 (O_1621,N_24680,N_24272);
or UO_1622 (O_1622,N_24135,N_24907);
and UO_1623 (O_1623,N_24140,N_24156);
and UO_1624 (O_1624,N_24976,N_24503);
nor UO_1625 (O_1625,N_24046,N_24821);
xor UO_1626 (O_1626,N_24504,N_24313);
xor UO_1627 (O_1627,N_24377,N_24056);
xor UO_1628 (O_1628,N_24499,N_24061);
nand UO_1629 (O_1629,N_24451,N_24146);
xor UO_1630 (O_1630,N_24950,N_24088);
nand UO_1631 (O_1631,N_24247,N_24009);
or UO_1632 (O_1632,N_24076,N_24978);
or UO_1633 (O_1633,N_24926,N_24794);
and UO_1634 (O_1634,N_24757,N_24304);
nand UO_1635 (O_1635,N_24435,N_24159);
and UO_1636 (O_1636,N_24322,N_24075);
or UO_1637 (O_1637,N_24969,N_24167);
nor UO_1638 (O_1638,N_24053,N_24909);
nor UO_1639 (O_1639,N_24151,N_24047);
nand UO_1640 (O_1640,N_24555,N_24106);
or UO_1641 (O_1641,N_24433,N_24723);
or UO_1642 (O_1642,N_24521,N_24211);
xor UO_1643 (O_1643,N_24471,N_24594);
and UO_1644 (O_1644,N_24651,N_24379);
and UO_1645 (O_1645,N_24823,N_24358);
and UO_1646 (O_1646,N_24765,N_24287);
xor UO_1647 (O_1647,N_24920,N_24149);
nand UO_1648 (O_1648,N_24467,N_24176);
nor UO_1649 (O_1649,N_24595,N_24593);
nor UO_1650 (O_1650,N_24077,N_24580);
or UO_1651 (O_1651,N_24461,N_24436);
xor UO_1652 (O_1652,N_24269,N_24430);
xor UO_1653 (O_1653,N_24842,N_24895);
or UO_1654 (O_1654,N_24655,N_24279);
nor UO_1655 (O_1655,N_24477,N_24473);
xnor UO_1656 (O_1656,N_24804,N_24246);
and UO_1657 (O_1657,N_24155,N_24078);
or UO_1658 (O_1658,N_24587,N_24590);
and UO_1659 (O_1659,N_24594,N_24824);
xnor UO_1660 (O_1660,N_24293,N_24612);
xnor UO_1661 (O_1661,N_24055,N_24407);
xor UO_1662 (O_1662,N_24950,N_24161);
nor UO_1663 (O_1663,N_24769,N_24023);
xnor UO_1664 (O_1664,N_24905,N_24819);
or UO_1665 (O_1665,N_24912,N_24911);
nor UO_1666 (O_1666,N_24040,N_24680);
xor UO_1667 (O_1667,N_24574,N_24912);
nor UO_1668 (O_1668,N_24707,N_24358);
and UO_1669 (O_1669,N_24538,N_24834);
xnor UO_1670 (O_1670,N_24297,N_24083);
or UO_1671 (O_1671,N_24521,N_24685);
xnor UO_1672 (O_1672,N_24995,N_24274);
xnor UO_1673 (O_1673,N_24987,N_24747);
nor UO_1674 (O_1674,N_24080,N_24178);
nand UO_1675 (O_1675,N_24242,N_24931);
nand UO_1676 (O_1676,N_24351,N_24583);
or UO_1677 (O_1677,N_24298,N_24520);
or UO_1678 (O_1678,N_24636,N_24092);
or UO_1679 (O_1679,N_24995,N_24032);
and UO_1680 (O_1680,N_24577,N_24099);
nand UO_1681 (O_1681,N_24050,N_24152);
nand UO_1682 (O_1682,N_24242,N_24319);
or UO_1683 (O_1683,N_24095,N_24509);
nor UO_1684 (O_1684,N_24546,N_24451);
nand UO_1685 (O_1685,N_24935,N_24555);
xor UO_1686 (O_1686,N_24869,N_24456);
or UO_1687 (O_1687,N_24205,N_24392);
xnor UO_1688 (O_1688,N_24670,N_24039);
nor UO_1689 (O_1689,N_24669,N_24834);
and UO_1690 (O_1690,N_24823,N_24211);
nor UO_1691 (O_1691,N_24935,N_24317);
xnor UO_1692 (O_1692,N_24916,N_24051);
nand UO_1693 (O_1693,N_24811,N_24423);
xor UO_1694 (O_1694,N_24128,N_24481);
and UO_1695 (O_1695,N_24957,N_24356);
xnor UO_1696 (O_1696,N_24873,N_24451);
or UO_1697 (O_1697,N_24714,N_24722);
and UO_1698 (O_1698,N_24992,N_24795);
nand UO_1699 (O_1699,N_24752,N_24660);
nor UO_1700 (O_1700,N_24700,N_24882);
xor UO_1701 (O_1701,N_24584,N_24919);
or UO_1702 (O_1702,N_24486,N_24968);
or UO_1703 (O_1703,N_24850,N_24081);
nor UO_1704 (O_1704,N_24548,N_24296);
and UO_1705 (O_1705,N_24700,N_24130);
nor UO_1706 (O_1706,N_24154,N_24999);
nand UO_1707 (O_1707,N_24779,N_24224);
nand UO_1708 (O_1708,N_24380,N_24907);
nor UO_1709 (O_1709,N_24075,N_24762);
or UO_1710 (O_1710,N_24640,N_24216);
nand UO_1711 (O_1711,N_24568,N_24862);
nor UO_1712 (O_1712,N_24504,N_24169);
and UO_1713 (O_1713,N_24573,N_24811);
and UO_1714 (O_1714,N_24696,N_24863);
nor UO_1715 (O_1715,N_24849,N_24243);
xnor UO_1716 (O_1716,N_24622,N_24377);
nor UO_1717 (O_1717,N_24880,N_24902);
xnor UO_1718 (O_1718,N_24521,N_24383);
xor UO_1719 (O_1719,N_24274,N_24549);
and UO_1720 (O_1720,N_24163,N_24114);
xor UO_1721 (O_1721,N_24008,N_24517);
nor UO_1722 (O_1722,N_24819,N_24146);
xnor UO_1723 (O_1723,N_24581,N_24277);
nor UO_1724 (O_1724,N_24376,N_24674);
nand UO_1725 (O_1725,N_24145,N_24013);
or UO_1726 (O_1726,N_24474,N_24795);
nor UO_1727 (O_1727,N_24833,N_24270);
xnor UO_1728 (O_1728,N_24588,N_24719);
nand UO_1729 (O_1729,N_24047,N_24015);
and UO_1730 (O_1730,N_24480,N_24754);
and UO_1731 (O_1731,N_24511,N_24727);
and UO_1732 (O_1732,N_24678,N_24682);
and UO_1733 (O_1733,N_24133,N_24529);
xnor UO_1734 (O_1734,N_24746,N_24497);
and UO_1735 (O_1735,N_24590,N_24637);
and UO_1736 (O_1736,N_24017,N_24753);
or UO_1737 (O_1737,N_24783,N_24365);
or UO_1738 (O_1738,N_24539,N_24291);
xnor UO_1739 (O_1739,N_24924,N_24157);
xor UO_1740 (O_1740,N_24081,N_24873);
or UO_1741 (O_1741,N_24920,N_24775);
and UO_1742 (O_1742,N_24752,N_24952);
xor UO_1743 (O_1743,N_24388,N_24140);
nor UO_1744 (O_1744,N_24192,N_24214);
xnor UO_1745 (O_1745,N_24690,N_24142);
and UO_1746 (O_1746,N_24399,N_24078);
nor UO_1747 (O_1747,N_24944,N_24389);
or UO_1748 (O_1748,N_24909,N_24279);
or UO_1749 (O_1749,N_24155,N_24386);
nor UO_1750 (O_1750,N_24313,N_24690);
and UO_1751 (O_1751,N_24953,N_24172);
or UO_1752 (O_1752,N_24127,N_24982);
xnor UO_1753 (O_1753,N_24698,N_24224);
xor UO_1754 (O_1754,N_24252,N_24023);
and UO_1755 (O_1755,N_24574,N_24638);
nor UO_1756 (O_1756,N_24462,N_24165);
nand UO_1757 (O_1757,N_24286,N_24049);
nand UO_1758 (O_1758,N_24402,N_24781);
nor UO_1759 (O_1759,N_24895,N_24174);
nand UO_1760 (O_1760,N_24556,N_24788);
xnor UO_1761 (O_1761,N_24360,N_24067);
xor UO_1762 (O_1762,N_24582,N_24062);
and UO_1763 (O_1763,N_24083,N_24480);
nor UO_1764 (O_1764,N_24064,N_24710);
and UO_1765 (O_1765,N_24328,N_24525);
nor UO_1766 (O_1766,N_24653,N_24348);
or UO_1767 (O_1767,N_24825,N_24170);
nor UO_1768 (O_1768,N_24985,N_24857);
and UO_1769 (O_1769,N_24659,N_24132);
and UO_1770 (O_1770,N_24680,N_24511);
or UO_1771 (O_1771,N_24429,N_24562);
and UO_1772 (O_1772,N_24689,N_24635);
nand UO_1773 (O_1773,N_24915,N_24214);
or UO_1774 (O_1774,N_24069,N_24340);
nor UO_1775 (O_1775,N_24405,N_24813);
nor UO_1776 (O_1776,N_24706,N_24769);
and UO_1777 (O_1777,N_24670,N_24151);
nand UO_1778 (O_1778,N_24176,N_24835);
and UO_1779 (O_1779,N_24211,N_24178);
xor UO_1780 (O_1780,N_24033,N_24783);
nand UO_1781 (O_1781,N_24517,N_24800);
xnor UO_1782 (O_1782,N_24639,N_24347);
and UO_1783 (O_1783,N_24698,N_24950);
or UO_1784 (O_1784,N_24630,N_24327);
nor UO_1785 (O_1785,N_24185,N_24658);
and UO_1786 (O_1786,N_24264,N_24928);
and UO_1787 (O_1787,N_24282,N_24715);
or UO_1788 (O_1788,N_24937,N_24602);
xnor UO_1789 (O_1789,N_24677,N_24845);
nor UO_1790 (O_1790,N_24546,N_24101);
xor UO_1791 (O_1791,N_24938,N_24778);
or UO_1792 (O_1792,N_24844,N_24635);
and UO_1793 (O_1793,N_24092,N_24976);
or UO_1794 (O_1794,N_24516,N_24429);
nor UO_1795 (O_1795,N_24295,N_24456);
nor UO_1796 (O_1796,N_24354,N_24642);
or UO_1797 (O_1797,N_24218,N_24677);
or UO_1798 (O_1798,N_24871,N_24170);
nand UO_1799 (O_1799,N_24123,N_24040);
xnor UO_1800 (O_1800,N_24644,N_24921);
xnor UO_1801 (O_1801,N_24370,N_24083);
xor UO_1802 (O_1802,N_24819,N_24851);
nor UO_1803 (O_1803,N_24935,N_24835);
xnor UO_1804 (O_1804,N_24568,N_24798);
nand UO_1805 (O_1805,N_24848,N_24754);
nand UO_1806 (O_1806,N_24478,N_24723);
or UO_1807 (O_1807,N_24322,N_24384);
or UO_1808 (O_1808,N_24889,N_24439);
and UO_1809 (O_1809,N_24170,N_24517);
nand UO_1810 (O_1810,N_24080,N_24051);
xor UO_1811 (O_1811,N_24281,N_24131);
xnor UO_1812 (O_1812,N_24167,N_24316);
nor UO_1813 (O_1813,N_24354,N_24388);
and UO_1814 (O_1814,N_24169,N_24447);
nand UO_1815 (O_1815,N_24696,N_24234);
and UO_1816 (O_1816,N_24793,N_24732);
nand UO_1817 (O_1817,N_24541,N_24012);
and UO_1818 (O_1818,N_24651,N_24842);
and UO_1819 (O_1819,N_24106,N_24975);
or UO_1820 (O_1820,N_24102,N_24010);
xnor UO_1821 (O_1821,N_24192,N_24851);
nand UO_1822 (O_1822,N_24680,N_24644);
or UO_1823 (O_1823,N_24942,N_24762);
xnor UO_1824 (O_1824,N_24995,N_24103);
nor UO_1825 (O_1825,N_24240,N_24469);
nor UO_1826 (O_1826,N_24337,N_24868);
and UO_1827 (O_1827,N_24060,N_24256);
xor UO_1828 (O_1828,N_24168,N_24955);
xor UO_1829 (O_1829,N_24927,N_24528);
and UO_1830 (O_1830,N_24966,N_24625);
xnor UO_1831 (O_1831,N_24498,N_24304);
and UO_1832 (O_1832,N_24631,N_24238);
or UO_1833 (O_1833,N_24844,N_24287);
nand UO_1834 (O_1834,N_24472,N_24381);
nor UO_1835 (O_1835,N_24027,N_24631);
nor UO_1836 (O_1836,N_24327,N_24813);
nor UO_1837 (O_1837,N_24880,N_24690);
and UO_1838 (O_1838,N_24452,N_24051);
or UO_1839 (O_1839,N_24498,N_24336);
xnor UO_1840 (O_1840,N_24058,N_24996);
and UO_1841 (O_1841,N_24102,N_24512);
xnor UO_1842 (O_1842,N_24824,N_24443);
or UO_1843 (O_1843,N_24617,N_24687);
xnor UO_1844 (O_1844,N_24270,N_24447);
or UO_1845 (O_1845,N_24681,N_24468);
and UO_1846 (O_1846,N_24400,N_24276);
and UO_1847 (O_1847,N_24614,N_24995);
or UO_1848 (O_1848,N_24478,N_24710);
xnor UO_1849 (O_1849,N_24655,N_24664);
xor UO_1850 (O_1850,N_24907,N_24730);
or UO_1851 (O_1851,N_24950,N_24683);
or UO_1852 (O_1852,N_24814,N_24922);
and UO_1853 (O_1853,N_24705,N_24925);
xnor UO_1854 (O_1854,N_24893,N_24650);
and UO_1855 (O_1855,N_24605,N_24548);
nor UO_1856 (O_1856,N_24753,N_24696);
or UO_1857 (O_1857,N_24433,N_24438);
and UO_1858 (O_1858,N_24133,N_24022);
nand UO_1859 (O_1859,N_24160,N_24710);
nand UO_1860 (O_1860,N_24743,N_24508);
xor UO_1861 (O_1861,N_24021,N_24663);
nor UO_1862 (O_1862,N_24563,N_24597);
xnor UO_1863 (O_1863,N_24955,N_24872);
nand UO_1864 (O_1864,N_24727,N_24634);
and UO_1865 (O_1865,N_24461,N_24324);
or UO_1866 (O_1866,N_24244,N_24089);
nor UO_1867 (O_1867,N_24327,N_24890);
nor UO_1868 (O_1868,N_24406,N_24228);
or UO_1869 (O_1869,N_24340,N_24380);
or UO_1870 (O_1870,N_24981,N_24107);
or UO_1871 (O_1871,N_24622,N_24214);
and UO_1872 (O_1872,N_24346,N_24659);
xnor UO_1873 (O_1873,N_24771,N_24224);
nand UO_1874 (O_1874,N_24434,N_24581);
and UO_1875 (O_1875,N_24388,N_24422);
or UO_1876 (O_1876,N_24135,N_24419);
nand UO_1877 (O_1877,N_24257,N_24670);
nand UO_1878 (O_1878,N_24248,N_24743);
nor UO_1879 (O_1879,N_24017,N_24496);
or UO_1880 (O_1880,N_24188,N_24149);
xnor UO_1881 (O_1881,N_24409,N_24317);
nor UO_1882 (O_1882,N_24658,N_24224);
or UO_1883 (O_1883,N_24743,N_24607);
xor UO_1884 (O_1884,N_24276,N_24600);
nand UO_1885 (O_1885,N_24498,N_24631);
or UO_1886 (O_1886,N_24654,N_24335);
and UO_1887 (O_1887,N_24407,N_24530);
or UO_1888 (O_1888,N_24742,N_24462);
nand UO_1889 (O_1889,N_24940,N_24944);
or UO_1890 (O_1890,N_24057,N_24485);
xnor UO_1891 (O_1891,N_24065,N_24139);
or UO_1892 (O_1892,N_24948,N_24093);
nor UO_1893 (O_1893,N_24516,N_24177);
and UO_1894 (O_1894,N_24940,N_24792);
or UO_1895 (O_1895,N_24215,N_24837);
nor UO_1896 (O_1896,N_24362,N_24565);
and UO_1897 (O_1897,N_24972,N_24969);
nor UO_1898 (O_1898,N_24708,N_24860);
and UO_1899 (O_1899,N_24907,N_24965);
nor UO_1900 (O_1900,N_24620,N_24507);
or UO_1901 (O_1901,N_24221,N_24541);
xor UO_1902 (O_1902,N_24518,N_24991);
and UO_1903 (O_1903,N_24230,N_24343);
or UO_1904 (O_1904,N_24247,N_24145);
xor UO_1905 (O_1905,N_24778,N_24591);
nor UO_1906 (O_1906,N_24175,N_24515);
xor UO_1907 (O_1907,N_24040,N_24063);
xor UO_1908 (O_1908,N_24505,N_24762);
and UO_1909 (O_1909,N_24831,N_24765);
or UO_1910 (O_1910,N_24098,N_24635);
nand UO_1911 (O_1911,N_24215,N_24886);
xor UO_1912 (O_1912,N_24645,N_24145);
and UO_1913 (O_1913,N_24443,N_24359);
nor UO_1914 (O_1914,N_24349,N_24855);
nor UO_1915 (O_1915,N_24523,N_24050);
or UO_1916 (O_1916,N_24910,N_24360);
nand UO_1917 (O_1917,N_24457,N_24461);
or UO_1918 (O_1918,N_24663,N_24291);
and UO_1919 (O_1919,N_24010,N_24998);
and UO_1920 (O_1920,N_24194,N_24581);
nand UO_1921 (O_1921,N_24334,N_24107);
and UO_1922 (O_1922,N_24173,N_24923);
or UO_1923 (O_1923,N_24457,N_24624);
and UO_1924 (O_1924,N_24127,N_24917);
and UO_1925 (O_1925,N_24296,N_24402);
nor UO_1926 (O_1926,N_24392,N_24787);
or UO_1927 (O_1927,N_24011,N_24466);
nand UO_1928 (O_1928,N_24635,N_24374);
or UO_1929 (O_1929,N_24164,N_24233);
nor UO_1930 (O_1930,N_24897,N_24472);
xnor UO_1931 (O_1931,N_24246,N_24094);
and UO_1932 (O_1932,N_24775,N_24549);
nand UO_1933 (O_1933,N_24284,N_24856);
or UO_1934 (O_1934,N_24319,N_24156);
or UO_1935 (O_1935,N_24850,N_24044);
xnor UO_1936 (O_1936,N_24788,N_24197);
and UO_1937 (O_1937,N_24718,N_24781);
nor UO_1938 (O_1938,N_24762,N_24099);
or UO_1939 (O_1939,N_24847,N_24003);
xor UO_1940 (O_1940,N_24495,N_24568);
xor UO_1941 (O_1941,N_24412,N_24351);
and UO_1942 (O_1942,N_24327,N_24569);
and UO_1943 (O_1943,N_24862,N_24863);
nand UO_1944 (O_1944,N_24914,N_24917);
nor UO_1945 (O_1945,N_24509,N_24705);
nor UO_1946 (O_1946,N_24927,N_24865);
nor UO_1947 (O_1947,N_24278,N_24563);
nand UO_1948 (O_1948,N_24612,N_24680);
nand UO_1949 (O_1949,N_24703,N_24625);
and UO_1950 (O_1950,N_24284,N_24437);
or UO_1951 (O_1951,N_24235,N_24823);
or UO_1952 (O_1952,N_24587,N_24311);
nand UO_1953 (O_1953,N_24960,N_24819);
or UO_1954 (O_1954,N_24853,N_24829);
xnor UO_1955 (O_1955,N_24516,N_24022);
nor UO_1956 (O_1956,N_24092,N_24926);
xnor UO_1957 (O_1957,N_24561,N_24495);
xor UO_1958 (O_1958,N_24570,N_24105);
nand UO_1959 (O_1959,N_24608,N_24601);
nor UO_1960 (O_1960,N_24922,N_24725);
nor UO_1961 (O_1961,N_24525,N_24879);
nor UO_1962 (O_1962,N_24608,N_24983);
xnor UO_1963 (O_1963,N_24338,N_24846);
and UO_1964 (O_1964,N_24471,N_24703);
nand UO_1965 (O_1965,N_24695,N_24814);
nor UO_1966 (O_1966,N_24441,N_24899);
nand UO_1967 (O_1967,N_24983,N_24812);
or UO_1968 (O_1968,N_24242,N_24733);
and UO_1969 (O_1969,N_24247,N_24531);
and UO_1970 (O_1970,N_24580,N_24374);
and UO_1971 (O_1971,N_24173,N_24988);
xnor UO_1972 (O_1972,N_24011,N_24599);
xor UO_1973 (O_1973,N_24913,N_24595);
nand UO_1974 (O_1974,N_24438,N_24253);
nor UO_1975 (O_1975,N_24295,N_24666);
or UO_1976 (O_1976,N_24771,N_24322);
xnor UO_1977 (O_1977,N_24634,N_24601);
and UO_1978 (O_1978,N_24833,N_24509);
nand UO_1979 (O_1979,N_24335,N_24709);
and UO_1980 (O_1980,N_24199,N_24453);
xor UO_1981 (O_1981,N_24697,N_24440);
nor UO_1982 (O_1982,N_24152,N_24941);
xor UO_1983 (O_1983,N_24528,N_24398);
nand UO_1984 (O_1984,N_24015,N_24196);
and UO_1985 (O_1985,N_24427,N_24122);
xnor UO_1986 (O_1986,N_24846,N_24930);
nor UO_1987 (O_1987,N_24623,N_24055);
and UO_1988 (O_1988,N_24837,N_24323);
nand UO_1989 (O_1989,N_24537,N_24991);
or UO_1990 (O_1990,N_24863,N_24734);
or UO_1991 (O_1991,N_24104,N_24053);
and UO_1992 (O_1992,N_24884,N_24176);
nand UO_1993 (O_1993,N_24958,N_24260);
nor UO_1994 (O_1994,N_24819,N_24475);
nor UO_1995 (O_1995,N_24484,N_24276);
or UO_1996 (O_1996,N_24417,N_24639);
or UO_1997 (O_1997,N_24355,N_24230);
nand UO_1998 (O_1998,N_24948,N_24857);
nand UO_1999 (O_1999,N_24790,N_24779);
nand UO_2000 (O_2000,N_24208,N_24591);
nand UO_2001 (O_2001,N_24897,N_24274);
xnor UO_2002 (O_2002,N_24531,N_24898);
xor UO_2003 (O_2003,N_24032,N_24898);
nand UO_2004 (O_2004,N_24104,N_24517);
or UO_2005 (O_2005,N_24427,N_24139);
nand UO_2006 (O_2006,N_24680,N_24455);
xnor UO_2007 (O_2007,N_24811,N_24342);
and UO_2008 (O_2008,N_24948,N_24217);
nand UO_2009 (O_2009,N_24893,N_24390);
nand UO_2010 (O_2010,N_24621,N_24453);
and UO_2011 (O_2011,N_24023,N_24560);
nor UO_2012 (O_2012,N_24079,N_24529);
or UO_2013 (O_2013,N_24115,N_24339);
nor UO_2014 (O_2014,N_24980,N_24665);
nor UO_2015 (O_2015,N_24097,N_24784);
nand UO_2016 (O_2016,N_24257,N_24519);
or UO_2017 (O_2017,N_24073,N_24975);
xor UO_2018 (O_2018,N_24153,N_24842);
nand UO_2019 (O_2019,N_24470,N_24838);
and UO_2020 (O_2020,N_24559,N_24967);
nand UO_2021 (O_2021,N_24292,N_24473);
or UO_2022 (O_2022,N_24742,N_24717);
or UO_2023 (O_2023,N_24658,N_24320);
and UO_2024 (O_2024,N_24751,N_24081);
nand UO_2025 (O_2025,N_24085,N_24385);
or UO_2026 (O_2026,N_24603,N_24627);
nand UO_2027 (O_2027,N_24489,N_24785);
xnor UO_2028 (O_2028,N_24862,N_24479);
nor UO_2029 (O_2029,N_24073,N_24439);
and UO_2030 (O_2030,N_24689,N_24020);
nand UO_2031 (O_2031,N_24662,N_24263);
and UO_2032 (O_2032,N_24452,N_24181);
nor UO_2033 (O_2033,N_24458,N_24797);
and UO_2034 (O_2034,N_24834,N_24232);
xor UO_2035 (O_2035,N_24890,N_24170);
xnor UO_2036 (O_2036,N_24789,N_24477);
or UO_2037 (O_2037,N_24178,N_24359);
nand UO_2038 (O_2038,N_24360,N_24692);
nor UO_2039 (O_2039,N_24356,N_24712);
or UO_2040 (O_2040,N_24942,N_24429);
xnor UO_2041 (O_2041,N_24068,N_24647);
nand UO_2042 (O_2042,N_24983,N_24895);
nor UO_2043 (O_2043,N_24999,N_24223);
nand UO_2044 (O_2044,N_24333,N_24596);
nand UO_2045 (O_2045,N_24905,N_24437);
or UO_2046 (O_2046,N_24424,N_24414);
xnor UO_2047 (O_2047,N_24026,N_24396);
and UO_2048 (O_2048,N_24071,N_24932);
xor UO_2049 (O_2049,N_24014,N_24151);
nand UO_2050 (O_2050,N_24912,N_24727);
xor UO_2051 (O_2051,N_24961,N_24488);
nor UO_2052 (O_2052,N_24785,N_24852);
or UO_2053 (O_2053,N_24098,N_24032);
xor UO_2054 (O_2054,N_24049,N_24270);
nand UO_2055 (O_2055,N_24447,N_24922);
nand UO_2056 (O_2056,N_24578,N_24853);
or UO_2057 (O_2057,N_24168,N_24184);
or UO_2058 (O_2058,N_24891,N_24815);
nor UO_2059 (O_2059,N_24843,N_24808);
and UO_2060 (O_2060,N_24133,N_24303);
xor UO_2061 (O_2061,N_24163,N_24596);
or UO_2062 (O_2062,N_24475,N_24860);
or UO_2063 (O_2063,N_24434,N_24145);
nand UO_2064 (O_2064,N_24249,N_24050);
nand UO_2065 (O_2065,N_24195,N_24646);
and UO_2066 (O_2066,N_24203,N_24915);
nor UO_2067 (O_2067,N_24748,N_24133);
nand UO_2068 (O_2068,N_24400,N_24815);
nand UO_2069 (O_2069,N_24686,N_24897);
nand UO_2070 (O_2070,N_24309,N_24890);
xnor UO_2071 (O_2071,N_24327,N_24817);
nor UO_2072 (O_2072,N_24526,N_24942);
xnor UO_2073 (O_2073,N_24336,N_24935);
nor UO_2074 (O_2074,N_24346,N_24122);
or UO_2075 (O_2075,N_24614,N_24115);
nor UO_2076 (O_2076,N_24668,N_24439);
or UO_2077 (O_2077,N_24754,N_24725);
xor UO_2078 (O_2078,N_24381,N_24279);
or UO_2079 (O_2079,N_24253,N_24701);
xnor UO_2080 (O_2080,N_24621,N_24068);
nor UO_2081 (O_2081,N_24643,N_24225);
nor UO_2082 (O_2082,N_24218,N_24053);
nor UO_2083 (O_2083,N_24537,N_24975);
xnor UO_2084 (O_2084,N_24483,N_24693);
or UO_2085 (O_2085,N_24046,N_24183);
and UO_2086 (O_2086,N_24608,N_24557);
nand UO_2087 (O_2087,N_24380,N_24941);
nand UO_2088 (O_2088,N_24031,N_24731);
or UO_2089 (O_2089,N_24348,N_24439);
or UO_2090 (O_2090,N_24776,N_24782);
and UO_2091 (O_2091,N_24867,N_24748);
nor UO_2092 (O_2092,N_24606,N_24495);
and UO_2093 (O_2093,N_24928,N_24356);
and UO_2094 (O_2094,N_24785,N_24059);
and UO_2095 (O_2095,N_24498,N_24425);
or UO_2096 (O_2096,N_24341,N_24452);
nand UO_2097 (O_2097,N_24368,N_24405);
nand UO_2098 (O_2098,N_24046,N_24288);
nor UO_2099 (O_2099,N_24976,N_24595);
xor UO_2100 (O_2100,N_24031,N_24880);
nand UO_2101 (O_2101,N_24408,N_24944);
and UO_2102 (O_2102,N_24307,N_24585);
nor UO_2103 (O_2103,N_24892,N_24584);
xnor UO_2104 (O_2104,N_24199,N_24551);
and UO_2105 (O_2105,N_24101,N_24497);
nand UO_2106 (O_2106,N_24846,N_24309);
nand UO_2107 (O_2107,N_24714,N_24833);
xnor UO_2108 (O_2108,N_24594,N_24677);
xor UO_2109 (O_2109,N_24874,N_24357);
and UO_2110 (O_2110,N_24718,N_24577);
xor UO_2111 (O_2111,N_24380,N_24149);
or UO_2112 (O_2112,N_24878,N_24752);
nand UO_2113 (O_2113,N_24776,N_24248);
xor UO_2114 (O_2114,N_24117,N_24894);
nor UO_2115 (O_2115,N_24910,N_24389);
or UO_2116 (O_2116,N_24552,N_24314);
and UO_2117 (O_2117,N_24304,N_24189);
or UO_2118 (O_2118,N_24073,N_24641);
nand UO_2119 (O_2119,N_24857,N_24349);
nand UO_2120 (O_2120,N_24714,N_24997);
nand UO_2121 (O_2121,N_24685,N_24836);
xor UO_2122 (O_2122,N_24008,N_24137);
nor UO_2123 (O_2123,N_24817,N_24649);
nor UO_2124 (O_2124,N_24606,N_24879);
and UO_2125 (O_2125,N_24284,N_24525);
nor UO_2126 (O_2126,N_24378,N_24842);
nor UO_2127 (O_2127,N_24038,N_24234);
and UO_2128 (O_2128,N_24916,N_24711);
nor UO_2129 (O_2129,N_24836,N_24313);
xor UO_2130 (O_2130,N_24263,N_24077);
nor UO_2131 (O_2131,N_24939,N_24913);
nand UO_2132 (O_2132,N_24454,N_24506);
and UO_2133 (O_2133,N_24571,N_24897);
nand UO_2134 (O_2134,N_24654,N_24738);
nor UO_2135 (O_2135,N_24104,N_24496);
xnor UO_2136 (O_2136,N_24547,N_24891);
xor UO_2137 (O_2137,N_24827,N_24775);
xor UO_2138 (O_2138,N_24966,N_24938);
nor UO_2139 (O_2139,N_24458,N_24477);
or UO_2140 (O_2140,N_24781,N_24516);
nor UO_2141 (O_2141,N_24741,N_24460);
xnor UO_2142 (O_2142,N_24080,N_24995);
nor UO_2143 (O_2143,N_24523,N_24407);
nor UO_2144 (O_2144,N_24448,N_24760);
xnor UO_2145 (O_2145,N_24678,N_24710);
nand UO_2146 (O_2146,N_24858,N_24773);
nand UO_2147 (O_2147,N_24329,N_24004);
or UO_2148 (O_2148,N_24962,N_24521);
or UO_2149 (O_2149,N_24261,N_24106);
nor UO_2150 (O_2150,N_24537,N_24365);
xnor UO_2151 (O_2151,N_24957,N_24845);
and UO_2152 (O_2152,N_24844,N_24768);
xnor UO_2153 (O_2153,N_24312,N_24301);
xor UO_2154 (O_2154,N_24499,N_24090);
nand UO_2155 (O_2155,N_24626,N_24269);
nor UO_2156 (O_2156,N_24799,N_24332);
nand UO_2157 (O_2157,N_24123,N_24535);
xnor UO_2158 (O_2158,N_24625,N_24476);
xnor UO_2159 (O_2159,N_24513,N_24052);
xnor UO_2160 (O_2160,N_24344,N_24175);
nor UO_2161 (O_2161,N_24241,N_24268);
or UO_2162 (O_2162,N_24465,N_24214);
and UO_2163 (O_2163,N_24170,N_24099);
xnor UO_2164 (O_2164,N_24484,N_24452);
or UO_2165 (O_2165,N_24924,N_24655);
nor UO_2166 (O_2166,N_24608,N_24090);
nand UO_2167 (O_2167,N_24681,N_24590);
or UO_2168 (O_2168,N_24425,N_24141);
or UO_2169 (O_2169,N_24426,N_24774);
or UO_2170 (O_2170,N_24557,N_24142);
xnor UO_2171 (O_2171,N_24556,N_24073);
xnor UO_2172 (O_2172,N_24275,N_24164);
nand UO_2173 (O_2173,N_24971,N_24805);
nand UO_2174 (O_2174,N_24273,N_24957);
and UO_2175 (O_2175,N_24191,N_24448);
or UO_2176 (O_2176,N_24931,N_24825);
and UO_2177 (O_2177,N_24158,N_24167);
or UO_2178 (O_2178,N_24162,N_24425);
nand UO_2179 (O_2179,N_24782,N_24639);
nand UO_2180 (O_2180,N_24466,N_24467);
nand UO_2181 (O_2181,N_24162,N_24389);
nand UO_2182 (O_2182,N_24831,N_24418);
nand UO_2183 (O_2183,N_24359,N_24708);
nand UO_2184 (O_2184,N_24199,N_24386);
nand UO_2185 (O_2185,N_24420,N_24915);
xnor UO_2186 (O_2186,N_24840,N_24671);
nand UO_2187 (O_2187,N_24065,N_24602);
xnor UO_2188 (O_2188,N_24303,N_24774);
and UO_2189 (O_2189,N_24546,N_24218);
nor UO_2190 (O_2190,N_24522,N_24306);
and UO_2191 (O_2191,N_24092,N_24842);
or UO_2192 (O_2192,N_24406,N_24893);
and UO_2193 (O_2193,N_24564,N_24731);
nor UO_2194 (O_2194,N_24902,N_24270);
nand UO_2195 (O_2195,N_24707,N_24806);
and UO_2196 (O_2196,N_24780,N_24712);
or UO_2197 (O_2197,N_24594,N_24689);
nand UO_2198 (O_2198,N_24744,N_24479);
and UO_2199 (O_2199,N_24850,N_24319);
or UO_2200 (O_2200,N_24903,N_24542);
and UO_2201 (O_2201,N_24931,N_24235);
nand UO_2202 (O_2202,N_24998,N_24840);
or UO_2203 (O_2203,N_24815,N_24590);
nand UO_2204 (O_2204,N_24317,N_24037);
nand UO_2205 (O_2205,N_24078,N_24896);
and UO_2206 (O_2206,N_24250,N_24731);
nor UO_2207 (O_2207,N_24939,N_24410);
and UO_2208 (O_2208,N_24745,N_24774);
nor UO_2209 (O_2209,N_24238,N_24103);
nand UO_2210 (O_2210,N_24970,N_24519);
and UO_2211 (O_2211,N_24712,N_24537);
and UO_2212 (O_2212,N_24768,N_24105);
and UO_2213 (O_2213,N_24556,N_24865);
or UO_2214 (O_2214,N_24702,N_24531);
and UO_2215 (O_2215,N_24342,N_24030);
nor UO_2216 (O_2216,N_24434,N_24641);
xnor UO_2217 (O_2217,N_24400,N_24423);
nor UO_2218 (O_2218,N_24559,N_24179);
and UO_2219 (O_2219,N_24482,N_24551);
or UO_2220 (O_2220,N_24895,N_24004);
or UO_2221 (O_2221,N_24330,N_24377);
and UO_2222 (O_2222,N_24765,N_24624);
nand UO_2223 (O_2223,N_24614,N_24471);
or UO_2224 (O_2224,N_24136,N_24349);
xor UO_2225 (O_2225,N_24039,N_24858);
xnor UO_2226 (O_2226,N_24023,N_24567);
xor UO_2227 (O_2227,N_24399,N_24071);
xnor UO_2228 (O_2228,N_24044,N_24595);
nand UO_2229 (O_2229,N_24496,N_24555);
xor UO_2230 (O_2230,N_24084,N_24546);
and UO_2231 (O_2231,N_24766,N_24282);
and UO_2232 (O_2232,N_24720,N_24625);
or UO_2233 (O_2233,N_24083,N_24270);
nor UO_2234 (O_2234,N_24651,N_24704);
xnor UO_2235 (O_2235,N_24295,N_24719);
and UO_2236 (O_2236,N_24433,N_24208);
nand UO_2237 (O_2237,N_24697,N_24448);
xnor UO_2238 (O_2238,N_24861,N_24939);
and UO_2239 (O_2239,N_24260,N_24370);
and UO_2240 (O_2240,N_24684,N_24502);
xor UO_2241 (O_2241,N_24501,N_24537);
and UO_2242 (O_2242,N_24817,N_24131);
xor UO_2243 (O_2243,N_24733,N_24468);
nor UO_2244 (O_2244,N_24356,N_24081);
xnor UO_2245 (O_2245,N_24589,N_24775);
and UO_2246 (O_2246,N_24785,N_24313);
nor UO_2247 (O_2247,N_24080,N_24150);
or UO_2248 (O_2248,N_24662,N_24949);
and UO_2249 (O_2249,N_24400,N_24835);
nand UO_2250 (O_2250,N_24834,N_24126);
xor UO_2251 (O_2251,N_24998,N_24187);
nand UO_2252 (O_2252,N_24021,N_24612);
nor UO_2253 (O_2253,N_24563,N_24708);
or UO_2254 (O_2254,N_24839,N_24678);
or UO_2255 (O_2255,N_24586,N_24976);
nand UO_2256 (O_2256,N_24855,N_24462);
or UO_2257 (O_2257,N_24204,N_24202);
nand UO_2258 (O_2258,N_24471,N_24304);
and UO_2259 (O_2259,N_24384,N_24730);
or UO_2260 (O_2260,N_24171,N_24905);
nand UO_2261 (O_2261,N_24828,N_24075);
or UO_2262 (O_2262,N_24989,N_24058);
and UO_2263 (O_2263,N_24960,N_24706);
nand UO_2264 (O_2264,N_24799,N_24526);
xor UO_2265 (O_2265,N_24308,N_24058);
xnor UO_2266 (O_2266,N_24474,N_24370);
nand UO_2267 (O_2267,N_24618,N_24072);
xor UO_2268 (O_2268,N_24574,N_24860);
or UO_2269 (O_2269,N_24640,N_24929);
nand UO_2270 (O_2270,N_24465,N_24792);
or UO_2271 (O_2271,N_24989,N_24065);
xor UO_2272 (O_2272,N_24176,N_24058);
nand UO_2273 (O_2273,N_24392,N_24099);
xnor UO_2274 (O_2274,N_24878,N_24135);
nor UO_2275 (O_2275,N_24747,N_24371);
nand UO_2276 (O_2276,N_24610,N_24753);
nand UO_2277 (O_2277,N_24311,N_24406);
or UO_2278 (O_2278,N_24095,N_24499);
nand UO_2279 (O_2279,N_24591,N_24553);
nand UO_2280 (O_2280,N_24870,N_24774);
or UO_2281 (O_2281,N_24735,N_24052);
or UO_2282 (O_2282,N_24385,N_24769);
nor UO_2283 (O_2283,N_24217,N_24002);
nor UO_2284 (O_2284,N_24257,N_24928);
xor UO_2285 (O_2285,N_24640,N_24977);
xnor UO_2286 (O_2286,N_24583,N_24675);
nand UO_2287 (O_2287,N_24392,N_24182);
nand UO_2288 (O_2288,N_24591,N_24722);
nand UO_2289 (O_2289,N_24141,N_24000);
or UO_2290 (O_2290,N_24444,N_24361);
and UO_2291 (O_2291,N_24426,N_24888);
nand UO_2292 (O_2292,N_24463,N_24524);
nand UO_2293 (O_2293,N_24948,N_24932);
nor UO_2294 (O_2294,N_24259,N_24178);
or UO_2295 (O_2295,N_24308,N_24617);
or UO_2296 (O_2296,N_24996,N_24158);
xor UO_2297 (O_2297,N_24579,N_24407);
nor UO_2298 (O_2298,N_24712,N_24329);
xnor UO_2299 (O_2299,N_24398,N_24402);
xnor UO_2300 (O_2300,N_24001,N_24432);
xor UO_2301 (O_2301,N_24511,N_24173);
nor UO_2302 (O_2302,N_24290,N_24194);
xnor UO_2303 (O_2303,N_24957,N_24518);
or UO_2304 (O_2304,N_24044,N_24638);
nand UO_2305 (O_2305,N_24327,N_24536);
or UO_2306 (O_2306,N_24243,N_24377);
and UO_2307 (O_2307,N_24087,N_24106);
or UO_2308 (O_2308,N_24231,N_24853);
xnor UO_2309 (O_2309,N_24854,N_24676);
nand UO_2310 (O_2310,N_24554,N_24823);
xor UO_2311 (O_2311,N_24107,N_24097);
or UO_2312 (O_2312,N_24806,N_24230);
and UO_2313 (O_2313,N_24667,N_24834);
or UO_2314 (O_2314,N_24379,N_24315);
or UO_2315 (O_2315,N_24650,N_24060);
and UO_2316 (O_2316,N_24235,N_24233);
or UO_2317 (O_2317,N_24089,N_24919);
and UO_2318 (O_2318,N_24207,N_24031);
nor UO_2319 (O_2319,N_24815,N_24648);
nand UO_2320 (O_2320,N_24799,N_24650);
and UO_2321 (O_2321,N_24965,N_24499);
nor UO_2322 (O_2322,N_24799,N_24959);
nand UO_2323 (O_2323,N_24052,N_24569);
xnor UO_2324 (O_2324,N_24950,N_24134);
and UO_2325 (O_2325,N_24532,N_24967);
nand UO_2326 (O_2326,N_24583,N_24886);
xor UO_2327 (O_2327,N_24303,N_24750);
or UO_2328 (O_2328,N_24008,N_24234);
xnor UO_2329 (O_2329,N_24569,N_24132);
nor UO_2330 (O_2330,N_24712,N_24699);
nand UO_2331 (O_2331,N_24068,N_24284);
xor UO_2332 (O_2332,N_24592,N_24032);
xor UO_2333 (O_2333,N_24852,N_24700);
xnor UO_2334 (O_2334,N_24038,N_24278);
nand UO_2335 (O_2335,N_24325,N_24142);
or UO_2336 (O_2336,N_24083,N_24840);
xor UO_2337 (O_2337,N_24478,N_24437);
and UO_2338 (O_2338,N_24212,N_24571);
or UO_2339 (O_2339,N_24992,N_24791);
or UO_2340 (O_2340,N_24265,N_24133);
or UO_2341 (O_2341,N_24325,N_24989);
and UO_2342 (O_2342,N_24983,N_24472);
or UO_2343 (O_2343,N_24628,N_24127);
or UO_2344 (O_2344,N_24659,N_24502);
and UO_2345 (O_2345,N_24610,N_24758);
nand UO_2346 (O_2346,N_24852,N_24943);
or UO_2347 (O_2347,N_24332,N_24318);
or UO_2348 (O_2348,N_24869,N_24445);
nor UO_2349 (O_2349,N_24168,N_24960);
nor UO_2350 (O_2350,N_24314,N_24143);
nand UO_2351 (O_2351,N_24707,N_24438);
nor UO_2352 (O_2352,N_24346,N_24304);
and UO_2353 (O_2353,N_24974,N_24715);
and UO_2354 (O_2354,N_24304,N_24827);
nand UO_2355 (O_2355,N_24806,N_24884);
and UO_2356 (O_2356,N_24886,N_24119);
or UO_2357 (O_2357,N_24336,N_24090);
or UO_2358 (O_2358,N_24659,N_24296);
xnor UO_2359 (O_2359,N_24087,N_24917);
nor UO_2360 (O_2360,N_24222,N_24141);
xor UO_2361 (O_2361,N_24245,N_24917);
xor UO_2362 (O_2362,N_24943,N_24710);
xnor UO_2363 (O_2363,N_24005,N_24871);
and UO_2364 (O_2364,N_24799,N_24745);
nand UO_2365 (O_2365,N_24164,N_24200);
nand UO_2366 (O_2366,N_24973,N_24190);
nand UO_2367 (O_2367,N_24801,N_24566);
nor UO_2368 (O_2368,N_24552,N_24477);
and UO_2369 (O_2369,N_24122,N_24054);
xnor UO_2370 (O_2370,N_24515,N_24093);
or UO_2371 (O_2371,N_24042,N_24497);
xnor UO_2372 (O_2372,N_24880,N_24939);
nand UO_2373 (O_2373,N_24453,N_24393);
or UO_2374 (O_2374,N_24275,N_24079);
xor UO_2375 (O_2375,N_24689,N_24063);
nor UO_2376 (O_2376,N_24143,N_24698);
nand UO_2377 (O_2377,N_24741,N_24939);
or UO_2378 (O_2378,N_24052,N_24486);
or UO_2379 (O_2379,N_24586,N_24524);
or UO_2380 (O_2380,N_24821,N_24792);
and UO_2381 (O_2381,N_24994,N_24254);
nand UO_2382 (O_2382,N_24450,N_24922);
or UO_2383 (O_2383,N_24999,N_24690);
and UO_2384 (O_2384,N_24343,N_24966);
xnor UO_2385 (O_2385,N_24599,N_24556);
nand UO_2386 (O_2386,N_24822,N_24988);
nor UO_2387 (O_2387,N_24060,N_24125);
xor UO_2388 (O_2388,N_24109,N_24267);
and UO_2389 (O_2389,N_24212,N_24638);
nand UO_2390 (O_2390,N_24000,N_24344);
or UO_2391 (O_2391,N_24524,N_24206);
nor UO_2392 (O_2392,N_24885,N_24456);
and UO_2393 (O_2393,N_24144,N_24538);
nand UO_2394 (O_2394,N_24651,N_24988);
and UO_2395 (O_2395,N_24632,N_24347);
xor UO_2396 (O_2396,N_24517,N_24609);
and UO_2397 (O_2397,N_24260,N_24065);
and UO_2398 (O_2398,N_24403,N_24096);
nor UO_2399 (O_2399,N_24035,N_24068);
xnor UO_2400 (O_2400,N_24988,N_24993);
xor UO_2401 (O_2401,N_24996,N_24408);
and UO_2402 (O_2402,N_24074,N_24758);
or UO_2403 (O_2403,N_24742,N_24697);
or UO_2404 (O_2404,N_24045,N_24227);
xnor UO_2405 (O_2405,N_24541,N_24262);
or UO_2406 (O_2406,N_24504,N_24840);
nor UO_2407 (O_2407,N_24626,N_24684);
nor UO_2408 (O_2408,N_24372,N_24370);
xor UO_2409 (O_2409,N_24897,N_24404);
nand UO_2410 (O_2410,N_24961,N_24131);
or UO_2411 (O_2411,N_24994,N_24143);
nor UO_2412 (O_2412,N_24042,N_24255);
and UO_2413 (O_2413,N_24452,N_24793);
nand UO_2414 (O_2414,N_24943,N_24595);
and UO_2415 (O_2415,N_24717,N_24562);
or UO_2416 (O_2416,N_24210,N_24807);
nand UO_2417 (O_2417,N_24301,N_24872);
nor UO_2418 (O_2418,N_24560,N_24006);
or UO_2419 (O_2419,N_24609,N_24718);
or UO_2420 (O_2420,N_24857,N_24130);
nor UO_2421 (O_2421,N_24055,N_24961);
xnor UO_2422 (O_2422,N_24953,N_24348);
and UO_2423 (O_2423,N_24444,N_24296);
nand UO_2424 (O_2424,N_24759,N_24036);
nand UO_2425 (O_2425,N_24538,N_24099);
nand UO_2426 (O_2426,N_24388,N_24261);
nor UO_2427 (O_2427,N_24876,N_24031);
or UO_2428 (O_2428,N_24047,N_24042);
nand UO_2429 (O_2429,N_24606,N_24136);
nand UO_2430 (O_2430,N_24099,N_24345);
and UO_2431 (O_2431,N_24030,N_24703);
nand UO_2432 (O_2432,N_24548,N_24383);
or UO_2433 (O_2433,N_24327,N_24908);
and UO_2434 (O_2434,N_24932,N_24586);
nand UO_2435 (O_2435,N_24488,N_24509);
xor UO_2436 (O_2436,N_24997,N_24662);
nand UO_2437 (O_2437,N_24291,N_24610);
or UO_2438 (O_2438,N_24009,N_24382);
xnor UO_2439 (O_2439,N_24854,N_24558);
nor UO_2440 (O_2440,N_24816,N_24860);
or UO_2441 (O_2441,N_24119,N_24559);
and UO_2442 (O_2442,N_24239,N_24121);
and UO_2443 (O_2443,N_24417,N_24065);
nand UO_2444 (O_2444,N_24485,N_24205);
nand UO_2445 (O_2445,N_24665,N_24523);
nand UO_2446 (O_2446,N_24929,N_24342);
nor UO_2447 (O_2447,N_24816,N_24005);
nand UO_2448 (O_2448,N_24320,N_24359);
nand UO_2449 (O_2449,N_24039,N_24208);
and UO_2450 (O_2450,N_24681,N_24878);
or UO_2451 (O_2451,N_24291,N_24588);
or UO_2452 (O_2452,N_24227,N_24571);
xnor UO_2453 (O_2453,N_24541,N_24363);
and UO_2454 (O_2454,N_24765,N_24444);
xor UO_2455 (O_2455,N_24298,N_24880);
nor UO_2456 (O_2456,N_24088,N_24607);
xnor UO_2457 (O_2457,N_24887,N_24282);
nand UO_2458 (O_2458,N_24978,N_24351);
nor UO_2459 (O_2459,N_24788,N_24297);
or UO_2460 (O_2460,N_24281,N_24788);
nand UO_2461 (O_2461,N_24576,N_24834);
and UO_2462 (O_2462,N_24561,N_24588);
nand UO_2463 (O_2463,N_24786,N_24788);
nor UO_2464 (O_2464,N_24596,N_24668);
or UO_2465 (O_2465,N_24338,N_24971);
nor UO_2466 (O_2466,N_24088,N_24618);
nor UO_2467 (O_2467,N_24058,N_24680);
nand UO_2468 (O_2468,N_24972,N_24044);
and UO_2469 (O_2469,N_24150,N_24130);
nand UO_2470 (O_2470,N_24651,N_24428);
xnor UO_2471 (O_2471,N_24931,N_24773);
xor UO_2472 (O_2472,N_24016,N_24058);
nand UO_2473 (O_2473,N_24911,N_24112);
xor UO_2474 (O_2474,N_24233,N_24197);
xnor UO_2475 (O_2475,N_24498,N_24753);
and UO_2476 (O_2476,N_24477,N_24715);
nand UO_2477 (O_2477,N_24091,N_24414);
xnor UO_2478 (O_2478,N_24795,N_24500);
xor UO_2479 (O_2479,N_24104,N_24361);
nand UO_2480 (O_2480,N_24232,N_24677);
and UO_2481 (O_2481,N_24817,N_24779);
or UO_2482 (O_2482,N_24160,N_24757);
or UO_2483 (O_2483,N_24035,N_24386);
xnor UO_2484 (O_2484,N_24331,N_24537);
xor UO_2485 (O_2485,N_24903,N_24905);
nor UO_2486 (O_2486,N_24950,N_24750);
xor UO_2487 (O_2487,N_24951,N_24850);
xnor UO_2488 (O_2488,N_24005,N_24168);
or UO_2489 (O_2489,N_24650,N_24123);
or UO_2490 (O_2490,N_24093,N_24144);
xnor UO_2491 (O_2491,N_24581,N_24021);
and UO_2492 (O_2492,N_24970,N_24228);
nand UO_2493 (O_2493,N_24645,N_24668);
and UO_2494 (O_2494,N_24708,N_24019);
nor UO_2495 (O_2495,N_24785,N_24483);
and UO_2496 (O_2496,N_24972,N_24336);
nand UO_2497 (O_2497,N_24340,N_24605);
nor UO_2498 (O_2498,N_24874,N_24802);
nand UO_2499 (O_2499,N_24905,N_24271);
and UO_2500 (O_2500,N_24457,N_24602);
nand UO_2501 (O_2501,N_24722,N_24678);
or UO_2502 (O_2502,N_24120,N_24877);
xnor UO_2503 (O_2503,N_24545,N_24715);
and UO_2504 (O_2504,N_24511,N_24955);
or UO_2505 (O_2505,N_24284,N_24313);
nor UO_2506 (O_2506,N_24816,N_24081);
nor UO_2507 (O_2507,N_24034,N_24206);
nor UO_2508 (O_2508,N_24631,N_24890);
xnor UO_2509 (O_2509,N_24202,N_24484);
xor UO_2510 (O_2510,N_24756,N_24658);
nor UO_2511 (O_2511,N_24024,N_24600);
xor UO_2512 (O_2512,N_24250,N_24997);
xor UO_2513 (O_2513,N_24391,N_24556);
or UO_2514 (O_2514,N_24880,N_24459);
nor UO_2515 (O_2515,N_24402,N_24544);
or UO_2516 (O_2516,N_24024,N_24367);
and UO_2517 (O_2517,N_24707,N_24429);
or UO_2518 (O_2518,N_24568,N_24068);
nor UO_2519 (O_2519,N_24257,N_24826);
xnor UO_2520 (O_2520,N_24560,N_24420);
nor UO_2521 (O_2521,N_24966,N_24783);
and UO_2522 (O_2522,N_24872,N_24896);
or UO_2523 (O_2523,N_24360,N_24922);
nor UO_2524 (O_2524,N_24616,N_24095);
nand UO_2525 (O_2525,N_24872,N_24804);
nand UO_2526 (O_2526,N_24693,N_24866);
xor UO_2527 (O_2527,N_24926,N_24594);
xor UO_2528 (O_2528,N_24874,N_24235);
nand UO_2529 (O_2529,N_24505,N_24919);
nand UO_2530 (O_2530,N_24537,N_24237);
and UO_2531 (O_2531,N_24972,N_24030);
and UO_2532 (O_2532,N_24817,N_24406);
nor UO_2533 (O_2533,N_24582,N_24294);
nor UO_2534 (O_2534,N_24459,N_24072);
and UO_2535 (O_2535,N_24982,N_24172);
and UO_2536 (O_2536,N_24945,N_24836);
nor UO_2537 (O_2537,N_24275,N_24545);
nand UO_2538 (O_2538,N_24273,N_24755);
nand UO_2539 (O_2539,N_24412,N_24190);
and UO_2540 (O_2540,N_24840,N_24709);
and UO_2541 (O_2541,N_24821,N_24764);
xor UO_2542 (O_2542,N_24590,N_24748);
xor UO_2543 (O_2543,N_24246,N_24123);
and UO_2544 (O_2544,N_24614,N_24228);
xnor UO_2545 (O_2545,N_24007,N_24701);
nand UO_2546 (O_2546,N_24132,N_24937);
nand UO_2547 (O_2547,N_24227,N_24269);
nand UO_2548 (O_2548,N_24907,N_24633);
and UO_2549 (O_2549,N_24664,N_24457);
nor UO_2550 (O_2550,N_24257,N_24087);
and UO_2551 (O_2551,N_24881,N_24957);
nand UO_2552 (O_2552,N_24368,N_24189);
nand UO_2553 (O_2553,N_24436,N_24490);
or UO_2554 (O_2554,N_24467,N_24656);
or UO_2555 (O_2555,N_24754,N_24940);
or UO_2556 (O_2556,N_24313,N_24198);
nand UO_2557 (O_2557,N_24645,N_24308);
xor UO_2558 (O_2558,N_24574,N_24512);
or UO_2559 (O_2559,N_24251,N_24805);
or UO_2560 (O_2560,N_24974,N_24237);
nand UO_2561 (O_2561,N_24696,N_24031);
nand UO_2562 (O_2562,N_24521,N_24833);
nor UO_2563 (O_2563,N_24259,N_24098);
nand UO_2564 (O_2564,N_24894,N_24790);
nand UO_2565 (O_2565,N_24122,N_24539);
or UO_2566 (O_2566,N_24705,N_24888);
nor UO_2567 (O_2567,N_24009,N_24353);
and UO_2568 (O_2568,N_24619,N_24245);
nand UO_2569 (O_2569,N_24079,N_24850);
and UO_2570 (O_2570,N_24230,N_24485);
xnor UO_2571 (O_2571,N_24388,N_24010);
xor UO_2572 (O_2572,N_24939,N_24032);
xor UO_2573 (O_2573,N_24979,N_24602);
and UO_2574 (O_2574,N_24238,N_24672);
nor UO_2575 (O_2575,N_24935,N_24536);
nor UO_2576 (O_2576,N_24680,N_24656);
nand UO_2577 (O_2577,N_24642,N_24982);
nor UO_2578 (O_2578,N_24178,N_24818);
xnor UO_2579 (O_2579,N_24079,N_24570);
or UO_2580 (O_2580,N_24587,N_24828);
nor UO_2581 (O_2581,N_24211,N_24009);
xor UO_2582 (O_2582,N_24011,N_24269);
nand UO_2583 (O_2583,N_24773,N_24489);
nand UO_2584 (O_2584,N_24703,N_24877);
nor UO_2585 (O_2585,N_24703,N_24602);
xnor UO_2586 (O_2586,N_24972,N_24681);
or UO_2587 (O_2587,N_24632,N_24321);
xor UO_2588 (O_2588,N_24216,N_24379);
xnor UO_2589 (O_2589,N_24401,N_24591);
nor UO_2590 (O_2590,N_24413,N_24016);
nand UO_2591 (O_2591,N_24370,N_24019);
nor UO_2592 (O_2592,N_24721,N_24162);
nor UO_2593 (O_2593,N_24060,N_24823);
xnor UO_2594 (O_2594,N_24671,N_24270);
nor UO_2595 (O_2595,N_24322,N_24183);
and UO_2596 (O_2596,N_24396,N_24717);
nand UO_2597 (O_2597,N_24554,N_24256);
or UO_2598 (O_2598,N_24925,N_24791);
or UO_2599 (O_2599,N_24606,N_24093);
and UO_2600 (O_2600,N_24748,N_24216);
nor UO_2601 (O_2601,N_24048,N_24369);
and UO_2602 (O_2602,N_24603,N_24375);
or UO_2603 (O_2603,N_24607,N_24156);
nor UO_2604 (O_2604,N_24267,N_24299);
nand UO_2605 (O_2605,N_24105,N_24396);
or UO_2606 (O_2606,N_24708,N_24312);
nand UO_2607 (O_2607,N_24883,N_24338);
nor UO_2608 (O_2608,N_24936,N_24300);
xnor UO_2609 (O_2609,N_24140,N_24108);
or UO_2610 (O_2610,N_24004,N_24911);
or UO_2611 (O_2611,N_24671,N_24759);
nand UO_2612 (O_2612,N_24592,N_24402);
nand UO_2613 (O_2613,N_24636,N_24417);
xnor UO_2614 (O_2614,N_24660,N_24208);
or UO_2615 (O_2615,N_24446,N_24685);
nand UO_2616 (O_2616,N_24152,N_24970);
and UO_2617 (O_2617,N_24403,N_24632);
nor UO_2618 (O_2618,N_24815,N_24518);
nor UO_2619 (O_2619,N_24775,N_24734);
nor UO_2620 (O_2620,N_24752,N_24932);
or UO_2621 (O_2621,N_24639,N_24105);
or UO_2622 (O_2622,N_24819,N_24404);
nor UO_2623 (O_2623,N_24698,N_24529);
nand UO_2624 (O_2624,N_24547,N_24675);
xnor UO_2625 (O_2625,N_24789,N_24753);
nand UO_2626 (O_2626,N_24292,N_24031);
and UO_2627 (O_2627,N_24179,N_24825);
or UO_2628 (O_2628,N_24725,N_24933);
or UO_2629 (O_2629,N_24064,N_24949);
nand UO_2630 (O_2630,N_24743,N_24531);
nand UO_2631 (O_2631,N_24805,N_24596);
or UO_2632 (O_2632,N_24640,N_24755);
xor UO_2633 (O_2633,N_24064,N_24432);
and UO_2634 (O_2634,N_24265,N_24155);
xnor UO_2635 (O_2635,N_24423,N_24328);
and UO_2636 (O_2636,N_24632,N_24262);
or UO_2637 (O_2637,N_24628,N_24798);
xnor UO_2638 (O_2638,N_24868,N_24734);
nand UO_2639 (O_2639,N_24245,N_24716);
xor UO_2640 (O_2640,N_24793,N_24049);
or UO_2641 (O_2641,N_24766,N_24324);
xnor UO_2642 (O_2642,N_24521,N_24920);
nand UO_2643 (O_2643,N_24987,N_24406);
or UO_2644 (O_2644,N_24329,N_24350);
or UO_2645 (O_2645,N_24034,N_24083);
and UO_2646 (O_2646,N_24034,N_24625);
nand UO_2647 (O_2647,N_24065,N_24215);
nor UO_2648 (O_2648,N_24373,N_24972);
xor UO_2649 (O_2649,N_24985,N_24490);
nor UO_2650 (O_2650,N_24237,N_24516);
and UO_2651 (O_2651,N_24702,N_24433);
nor UO_2652 (O_2652,N_24595,N_24544);
xor UO_2653 (O_2653,N_24510,N_24844);
and UO_2654 (O_2654,N_24445,N_24950);
nor UO_2655 (O_2655,N_24229,N_24976);
and UO_2656 (O_2656,N_24386,N_24204);
xnor UO_2657 (O_2657,N_24993,N_24182);
and UO_2658 (O_2658,N_24860,N_24081);
nor UO_2659 (O_2659,N_24761,N_24489);
nand UO_2660 (O_2660,N_24486,N_24939);
nand UO_2661 (O_2661,N_24106,N_24517);
nor UO_2662 (O_2662,N_24897,N_24525);
xnor UO_2663 (O_2663,N_24274,N_24687);
or UO_2664 (O_2664,N_24466,N_24126);
nand UO_2665 (O_2665,N_24835,N_24214);
or UO_2666 (O_2666,N_24193,N_24229);
xor UO_2667 (O_2667,N_24918,N_24376);
or UO_2668 (O_2668,N_24768,N_24599);
nor UO_2669 (O_2669,N_24625,N_24147);
or UO_2670 (O_2670,N_24767,N_24461);
and UO_2671 (O_2671,N_24279,N_24350);
nor UO_2672 (O_2672,N_24677,N_24168);
nor UO_2673 (O_2673,N_24964,N_24532);
nor UO_2674 (O_2674,N_24193,N_24838);
xnor UO_2675 (O_2675,N_24133,N_24174);
nor UO_2676 (O_2676,N_24183,N_24338);
nor UO_2677 (O_2677,N_24675,N_24460);
nor UO_2678 (O_2678,N_24949,N_24701);
nand UO_2679 (O_2679,N_24748,N_24120);
nand UO_2680 (O_2680,N_24038,N_24518);
or UO_2681 (O_2681,N_24403,N_24136);
or UO_2682 (O_2682,N_24113,N_24141);
nor UO_2683 (O_2683,N_24690,N_24212);
xnor UO_2684 (O_2684,N_24991,N_24102);
and UO_2685 (O_2685,N_24628,N_24235);
nor UO_2686 (O_2686,N_24154,N_24984);
nand UO_2687 (O_2687,N_24556,N_24776);
and UO_2688 (O_2688,N_24901,N_24035);
nor UO_2689 (O_2689,N_24767,N_24119);
nand UO_2690 (O_2690,N_24816,N_24503);
and UO_2691 (O_2691,N_24485,N_24752);
nor UO_2692 (O_2692,N_24443,N_24345);
or UO_2693 (O_2693,N_24829,N_24609);
or UO_2694 (O_2694,N_24207,N_24069);
and UO_2695 (O_2695,N_24046,N_24287);
or UO_2696 (O_2696,N_24386,N_24561);
and UO_2697 (O_2697,N_24179,N_24977);
xnor UO_2698 (O_2698,N_24754,N_24152);
nor UO_2699 (O_2699,N_24215,N_24495);
xnor UO_2700 (O_2700,N_24403,N_24495);
or UO_2701 (O_2701,N_24314,N_24548);
nor UO_2702 (O_2702,N_24949,N_24448);
nand UO_2703 (O_2703,N_24779,N_24394);
and UO_2704 (O_2704,N_24586,N_24605);
and UO_2705 (O_2705,N_24333,N_24108);
nand UO_2706 (O_2706,N_24749,N_24371);
and UO_2707 (O_2707,N_24918,N_24670);
or UO_2708 (O_2708,N_24387,N_24383);
nand UO_2709 (O_2709,N_24259,N_24999);
nor UO_2710 (O_2710,N_24375,N_24244);
nor UO_2711 (O_2711,N_24258,N_24216);
and UO_2712 (O_2712,N_24798,N_24646);
nor UO_2713 (O_2713,N_24757,N_24303);
nand UO_2714 (O_2714,N_24792,N_24585);
xnor UO_2715 (O_2715,N_24293,N_24850);
nor UO_2716 (O_2716,N_24186,N_24711);
and UO_2717 (O_2717,N_24693,N_24549);
or UO_2718 (O_2718,N_24253,N_24755);
xnor UO_2719 (O_2719,N_24404,N_24347);
xnor UO_2720 (O_2720,N_24311,N_24380);
and UO_2721 (O_2721,N_24725,N_24779);
xnor UO_2722 (O_2722,N_24690,N_24927);
or UO_2723 (O_2723,N_24723,N_24859);
and UO_2724 (O_2724,N_24539,N_24209);
or UO_2725 (O_2725,N_24235,N_24067);
xor UO_2726 (O_2726,N_24267,N_24305);
or UO_2727 (O_2727,N_24823,N_24818);
and UO_2728 (O_2728,N_24307,N_24426);
and UO_2729 (O_2729,N_24434,N_24431);
or UO_2730 (O_2730,N_24171,N_24189);
xor UO_2731 (O_2731,N_24730,N_24842);
or UO_2732 (O_2732,N_24739,N_24040);
nor UO_2733 (O_2733,N_24814,N_24112);
and UO_2734 (O_2734,N_24776,N_24924);
or UO_2735 (O_2735,N_24167,N_24413);
xnor UO_2736 (O_2736,N_24432,N_24473);
xnor UO_2737 (O_2737,N_24227,N_24266);
and UO_2738 (O_2738,N_24921,N_24525);
and UO_2739 (O_2739,N_24135,N_24290);
nand UO_2740 (O_2740,N_24121,N_24194);
xor UO_2741 (O_2741,N_24164,N_24238);
nand UO_2742 (O_2742,N_24606,N_24549);
nand UO_2743 (O_2743,N_24571,N_24396);
and UO_2744 (O_2744,N_24763,N_24302);
or UO_2745 (O_2745,N_24659,N_24986);
and UO_2746 (O_2746,N_24432,N_24654);
xnor UO_2747 (O_2747,N_24130,N_24469);
or UO_2748 (O_2748,N_24158,N_24758);
and UO_2749 (O_2749,N_24009,N_24723);
nor UO_2750 (O_2750,N_24052,N_24990);
nor UO_2751 (O_2751,N_24371,N_24316);
nor UO_2752 (O_2752,N_24274,N_24735);
nand UO_2753 (O_2753,N_24466,N_24023);
and UO_2754 (O_2754,N_24700,N_24458);
nor UO_2755 (O_2755,N_24945,N_24369);
nand UO_2756 (O_2756,N_24808,N_24242);
nor UO_2757 (O_2757,N_24238,N_24023);
nand UO_2758 (O_2758,N_24463,N_24301);
xnor UO_2759 (O_2759,N_24549,N_24618);
xnor UO_2760 (O_2760,N_24736,N_24260);
nand UO_2761 (O_2761,N_24057,N_24548);
xor UO_2762 (O_2762,N_24378,N_24065);
xnor UO_2763 (O_2763,N_24853,N_24467);
nand UO_2764 (O_2764,N_24963,N_24607);
nand UO_2765 (O_2765,N_24405,N_24703);
xor UO_2766 (O_2766,N_24677,N_24306);
xor UO_2767 (O_2767,N_24560,N_24504);
nand UO_2768 (O_2768,N_24852,N_24601);
and UO_2769 (O_2769,N_24373,N_24274);
nand UO_2770 (O_2770,N_24699,N_24291);
or UO_2771 (O_2771,N_24290,N_24579);
and UO_2772 (O_2772,N_24549,N_24887);
and UO_2773 (O_2773,N_24261,N_24814);
xor UO_2774 (O_2774,N_24773,N_24074);
nand UO_2775 (O_2775,N_24801,N_24141);
xnor UO_2776 (O_2776,N_24488,N_24785);
xor UO_2777 (O_2777,N_24514,N_24696);
and UO_2778 (O_2778,N_24131,N_24261);
or UO_2779 (O_2779,N_24844,N_24689);
nand UO_2780 (O_2780,N_24346,N_24858);
or UO_2781 (O_2781,N_24814,N_24860);
xnor UO_2782 (O_2782,N_24096,N_24882);
nand UO_2783 (O_2783,N_24546,N_24777);
nand UO_2784 (O_2784,N_24962,N_24129);
or UO_2785 (O_2785,N_24480,N_24298);
and UO_2786 (O_2786,N_24380,N_24982);
nor UO_2787 (O_2787,N_24112,N_24862);
xor UO_2788 (O_2788,N_24898,N_24649);
or UO_2789 (O_2789,N_24432,N_24204);
nor UO_2790 (O_2790,N_24523,N_24677);
and UO_2791 (O_2791,N_24334,N_24100);
nor UO_2792 (O_2792,N_24188,N_24686);
or UO_2793 (O_2793,N_24832,N_24630);
xnor UO_2794 (O_2794,N_24156,N_24505);
and UO_2795 (O_2795,N_24817,N_24453);
and UO_2796 (O_2796,N_24681,N_24346);
xor UO_2797 (O_2797,N_24894,N_24997);
nand UO_2798 (O_2798,N_24337,N_24516);
or UO_2799 (O_2799,N_24396,N_24478);
and UO_2800 (O_2800,N_24039,N_24106);
or UO_2801 (O_2801,N_24603,N_24619);
and UO_2802 (O_2802,N_24519,N_24863);
nand UO_2803 (O_2803,N_24029,N_24524);
nor UO_2804 (O_2804,N_24063,N_24589);
xor UO_2805 (O_2805,N_24214,N_24144);
nor UO_2806 (O_2806,N_24303,N_24128);
or UO_2807 (O_2807,N_24744,N_24047);
xnor UO_2808 (O_2808,N_24854,N_24840);
xnor UO_2809 (O_2809,N_24457,N_24989);
and UO_2810 (O_2810,N_24262,N_24145);
nor UO_2811 (O_2811,N_24194,N_24467);
or UO_2812 (O_2812,N_24743,N_24213);
and UO_2813 (O_2813,N_24827,N_24987);
or UO_2814 (O_2814,N_24170,N_24866);
and UO_2815 (O_2815,N_24001,N_24167);
nor UO_2816 (O_2816,N_24401,N_24758);
xor UO_2817 (O_2817,N_24723,N_24068);
and UO_2818 (O_2818,N_24814,N_24317);
nand UO_2819 (O_2819,N_24593,N_24692);
xnor UO_2820 (O_2820,N_24268,N_24167);
and UO_2821 (O_2821,N_24805,N_24103);
nor UO_2822 (O_2822,N_24259,N_24229);
nor UO_2823 (O_2823,N_24061,N_24238);
and UO_2824 (O_2824,N_24667,N_24147);
xnor UO_2825 (O_2825,N_24649,N_24091);
or UO_2826 (O_2826,N_24233,N_24687);
nand UO_2827 (O_2827,N_24090,N_24396);
xor UO_2828 (O_2828,N_24976,N_24975);
nor UO_2829 (O_2829,N_24610,N_24993);
or UO_2830 (O_2830,N_24737,N_24306);
nor UO_2831 (O_2831,N_24069,N_24004);
nand UO_2832 (O_2832,N_24642,N_24461);
nor UO_2833 (O_2833,N_24228,N_24102);
xor UO_2834 (O_2834,N_24637,N_24671);
nor UO_2835 (O_2835,N_24694,N_24018);
xor UO_2836 (O_2836,N_24470,N_24008);
nand UO_2837 (O_2837,N_24512,N_24741);
or UO_2838 (O_2838,N_24155,N_24063);
or UO_2839 (O_2839,N_24978,N_24806);
nor UO_2840 (O_2840,N_24032,N_24284);
xnor UO_2841 (O_2841,N_24315,N_24328);
nor UO_2842 (O_2842,N_24628,N_24616);
nor UO_2843 (O_2843,N_24833,N_24117);
or UO_2844 (O_2844,N_24040,N_24938);
or UO_2845 (O_2845,N_24032,N_24260);
or UO_2846 (O_2846,N_24212,N_24602);
nor UO_2847 (O_2847,N_24952,N_24045);
or UO_2848 (O_2848,N_24991,N_24364);
or UO_2849 (O_2849,N_24439,N_24197);
xor UO_2850 (O_2850,N_24732,N_24811);
or UO_2851 (O_2851,N_24390,N_24874);
and UO_2852 (O_2852,N_24147,N_24516);
and UO_2853 (O_2853,N_24081,N_24962);
xnor UO_2854 (O_2854,N_24029,N_24198);
nor UO_2855 (O_2855,N_24531,N_24151);
nor UO_2856 (O_2856,N_24428,N_24108);
nor UO_2857 (O_2857,N_24217,N_24442);
or UO_2858 (O_2858,N_24831,N_24725);
or UO_2859 (O_2859,N_24126,N_24202);
or UO_2860 (O_2860,N_24719,N_24891);
or UO_2861 (O_2861,N_24570,N_24101);
or UO_2862 (O_2862,N_24997,N_24070);
nand UO_2863 (O_2863,N_24457,N_24935);
and UO_2864 (O_2864,N_24800,N_24739);
nor UO_2865 (O_2865,N_24845,N_24653);
xnor UO_2866 (O_2866,N_24562,N_24661);
nand UO_2867 (O_2867,N_24116,N_24402);
nand UO_2868 (O_2868,N_24317,N_24669);
nor UO_2869 (O_2869,N_24403,N_24293);
nor UO_2870 (O_2870,N_24182,N_24413);
nand UO_2871 (O_2871,N_24833,N_24221);
or UO_2872 (O_2872,N_24185,N_24056);
and UO_2873 (O_2873,N_24231,N_24126);
and UO_2874 (O_2874,N_24664,N_24614);
or UO_2875 (O_2875,N_24956,N_24688);
xor UO_2876 (O_2876,N_24269,N_24046);
nor UO_2877 (O_2877,N_24881,N_24938);
or UO_2878 (O_2878,N_24084,N_24266);
xor UO_2879 (O_2879,N_24446,N_24634);
nor UO_2880 (O_2880,N_24231,N_24339);
or UO_2881 (O_2881,N_24576,N_24331);
xor UO_2882 (O_2882,N_24291,N_24638);
or UO_2883 (O_2883,N_24132,N_24568);
nor UO_2884 (O_2884,N_24183,N_24225);
nand UO_2885 (O_2885,N_24865,N_24884);
nor UO_2886 (O_2886,N_24151,N_24269);
and UO_2887 (O_2887,N_24018,N_24704);
nor UO_2888 (O_2888,N_24511,N_24888);
and UO_2889 (O_2889,N_24539,N_24344);
nand UO_2890 (O_2890,N_24925,N_24894);
nor UO_2891 (O_2891,N_24468,N_24645);
nor UO_2892 (O_2892,N_24581,N_24569);
and UO_2893 (O_2893,N_24056,N_24913);
xnor UO_2894 (O_2894,N_24161,N_24498);
nor UO_2895 (O_2895,N_24191,N_24420);
nand UO_2896 (O_2896,N_24270,N_24706);
nor UO_2897 (O_2897,N_24431,N_24634);
nor UO_2898 (O_2898,N_24224,N_24236);
nand UO_2899 (O_2899,N_24431,N_24909);
nand UO_2900 (O_2900,N_24086,N_24126);
and UO_2901 (O_2901,N_24929,N_24980);
xnor UO_2902 (O_2902,N_24255,N_24450);
or UO_2903 (O_2903,N_24796,N_24321);
nand UO_2904 (O_2904,N_24723,N_24681);
or UO_2905 (O_2905,N_24962,N_24747);
nand UO_2906 (O_2906,N_24591,N_24530);
xnor UO_2907 (O_2907,N_24428,N_24977);
or UO_2908 (O_2908,N_24068,N_24768);
and UO_2909 (O_2909,N_24421,N_24279);
xnor UO_2910 (O_2910,N_24507,N_24543);
and UO_2911 (O_2911,N_24584,N_24879);
nand UO_2912 (O_2912,N_24067,N_24742);
nand UO_2913 (O_2913,N_24742,N_24746);
and UO_2914 (O_2914,N_24371,N_24222);
and UO_2915 (O_2915,N_24395,N_24005);
nand UO_2916 (O_2916,N_24990,N_24801);
nor UO_2917 (O_2917,N_24324,N_24838);
and UO_2918 (O_2918,N_24076,N_24885);
or UO_2919 (O_2919,N_24167,N_24165);
and UO_2920 (O_2920,N_24999,N_24070);
nor UO_2921 (O_2921,N_24294,N_24814);
nor UO_2922 (O_2922,N_24391,N_24406);
and UO_2923 (O_2923,N_24117,N_24475);
and UO_2924 (O_2924,N_24087,N_24248);
xor UO_2925 (O_2925,N_24678,N_24137);
or UO_2926 (O_2926,N_24530,N_24668);
xnor UO_2927 (O_2927,N_24989,N_24312);
xnor UO_2928 (O_2928,N_24823,N_24359);
nand UO_2929 (O_2929,N_24440,N_24675);
xnor UO_2930 (O_2930,N_24925,N_24040);
nand UO_2931 (O_2931,N_24490,N_24359);
nor UO_2932 (O_2932,N_24195,N_24030);
nor UO_2933 (O_2933,N_24043,N_24729);
or UO_2934 (O_2934,N_24870,N_24638);
nor UO_2935 (O_2935,N_24077,N_24924);
nor UO_2936 (O_2936,N_24214,N_24913);
nand UO_2937 (O_2937,N_24042,N_24839);
or UO_2938 (O_2938,N_24194,N_24127);
nor UO_2939 (O_2939,N_24200,N_24221);
nand UO_2940 (O_2940,N_24510,N_24232);
and UO_2941 (O_2941,N_24374,N_24187);
nor UO_2942 (O_2942,N_24743,N_24086);
nor UO_2943 (O_2943,N_24650,N_24144);
xnor UO_2944 (O_2944,N_24476,N_24007);
nor UO_2945 (O_2945,N_24335,N_24683);
nor UO_2946 (O_2946,N_24353,N_24995);
nor UO_2947 (O_2947,N_24912,N_24443);
xor UO_2948 (O_2948,N_24590,N_24365);
or UO_2949 (O_2949,N_24615,N_24112);
nand UO_2950 (O_2950,N_24706,N_24772);
nand UO_2951 (O_2951,N_24770,N_24673);
or UO_2952 (O_2952,N_24790,N_24914);
nor UO_2953 (O_2953,N_24647,N_24141);
or UO_2954 (O_2954,N_24052,N_24761);
nand UO_2955 (O_2955,N_24692,N_24745);
xor UO_2956 (O_2956,N_24012,N_24784);
nor UO_2957 (O_2957,N_24173,N_24208);
nand UO_2958 (O_2958,N_24777,N_24309);
nand UO_2959 (O_2959,N_24165,N_24155);
and UO_2960 (O_2960,N_24096,N_24281);
nand UO_2961 (O_2961,N_24792,N_24446);
or UO_2962 (O_2962,N_24367,N_24259);
nand UO_2963 (O_2963,N_24470,N_24895);
nand UO_2964 (O_2964,N_24178,N_24737);
and UO_2965 (O_2965,N_24169,N_24548);
nor UO_2966 (O_2966,N_24706,N_24152);
or UO_2967 (O_2967,N_24432,N_24066);
or UO_2968 (O_2968,N_24265,N_24930);
nor UO_2969 (O_2969,N_24898,N_24641);
and UO_2970 (O_2970,N_24509,N_24431);
nand UO_2971 (O_2971,N_24651,N_24401);
nand UO_2972 (O_2972,N_24374,N_24311);
nor UO_2973 (O_2973,N_24658,N_24990);
and UO_2974 (O_2974,N_24454,N_24935);
nand UO_2975 (O_2975,N_24357,N_24080);
xnor UO_2976 (O_2976,N_24924,N_24608);
nor UO_2977 (O_2977,N_24948,N_24707);
nor UO_2978 (O_2978,N_24734,N_24605);
and UO_2979 (O_2979,N_24712,N_24630);
or UO_2980 (O_2980,N_24230,N_24031);
or UO_2981 (O_2981,N_24611,N_24196);
nand UO_2982 (O_2982,N_24377,N_24326);
and UO_2983 (O_2983,N_24250,N_24736);
nand UO_2984 (O_2984,N_24758,N_24667);
nor UO_2985 (O_2985,N_24194,N_24768);
nand UO_2986 (O_2986,N_24714,N_24576);
nand UO_2987 (O_2987,N_24147,N_24849);
nand UO_2988 (O_2988,N_24374,N_24995);
nor UO_2989 (O_2989,N_24688,N_24762);
nand UO_2990 (O_2990,N_24905,N_24071);
or UO_2991 (O_2991,N_24164,N_24810);
nor UO_2992 (O_2992,N_24451,N_24787);
and UO_2993 (O_2993,N_24980,N_24337);
nand UO_2994 (O_2994,N_24246,N_24064);
nand UO_2995 (O_2995,N_24483,N_24623);
xor UO_2996 (O_2996,N_24396,N_24185);
or UO_2997 (O_2997,N_24816,N_24777);
xor UO_2998 (O_2998,N_24450,N_24759);
xor UO_2999 (O_2999,N_24789,N_24402);
endmodule