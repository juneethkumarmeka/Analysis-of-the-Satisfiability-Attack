module basic_1000_10000_1500_50_levels_5xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
nor U0 (N_0,In_629,In_66);
nand U1 (N_1,In_210,In_87);
nor U2 (N_2,In_774,In_498);
xor U3 (N_3,In_638,In_471);
nor U4 (N_4,In_712,In_955);
nand U5 (N_5,In_903,In_331);
nand U6 (N_6,In_50,In_879);
or U7 (N_7,In_573,In_404);
nor U8 (N_8,In_613,In_634);
xnor U9 (N_9,In_457,In_109);
and U10 (N_10,In_939,In_162);
or U11 (N_11,In_298,In_342);
and U12 (N_12,In_691,In_98);
and U13 (N_13,In_891,In_385);
nor U14 (N_14,In_606,In_697);
nand U15 (N_15,In_520,In_172);
nor U16 (N_16,In_2,In_578);
or U17 (N_17,In_330,In_124);
nor U18 (N_18,In_390,In_149);
and U19 (N_19,In_301,In_846);
nand U20 (N_20,In_374,In_899);
and U21 (N_21,In_365,In_394);
or U22 (N_22,In_243,In_73);
xor U23 (N_23,In_798,In_770);
and U24 (N_24,In_459,In_384);
or U25 (N_25,In_536,In_541);
and U26 (N_26,In_917,In_57);
nor U27 (N_27,In_26,In_554);
nand U28 (N_28,In_853,In_991);
nand U29 (N_29,In_995,In_277);
nor U30 (N_30,In_362,In_960);
nor U31 (N_31,In_183,In_242);
nand U32 (N_32,In_503,In_418);
nor U33 (N_33,In_725,In_4);
nand U34 (N_34,In_300,In_969);
and U35 (N_35,In_211,In_169);
xor U36 (N_36,In_440,In_618);
nor U37 (N_37,In_364,In_681);
nor U38 (N_38,In_347,In_926);
xnor U39 (N_39,In_888,In_781);
or U40 (N_40,In_88,In_212);
xnor U41 (N_41,In_664,In_84);
nor U42 (N_42,In_21,In_892);
nor U43 (N_43,In_225,In_624);
or U44 (N_44,In_647,In_469);
nand U45 (N_45,In_906,In_462);
nand U46 (N_46,In_890,In_561);
nand U47 (N_47,In_549,In_114);
or U48 (N_48,In_942,In_830);
and U49 (N_49,In_274,In_768);
nor U50 (N_50,In_645,In_265);
nor U51 (N_51,In_376,In_810);
and U52 (N_52,In_333,In_945);
xnor U53 (N_53,In_420,In_68);
nor U54 (N_54,In_31,In_751);
and U55 (N_55,In_978,In_924);
xor U56 (N_56,In_154,In_22);
and U57 (N_57,In_95,In_894);
nor U58 (N_58,In_56,In_354);
or U59 (N_59,In_828,In_389);
xnor U60 (N_60,In_730,In_53);
nor U61 (N_61,In_249,In_270);
nand U62 (N_62,In_295,In_623);
or U63 (N_63,In_264,In_927);
xor U64 (N_64,In_334,In_657);
nand U65 (N_65,In_91,In_148);
and U66 (N_66,In_108,In_864);
or U67 (N_67,In_959,In_728);
or U68 (N_68,In_644,In_359);
or U69 (N_69,In_706,In_870);
nor U70 (N_70,In_332,In_209);
nor U71 (N_71,In_0,In_858);
nor U72 (N_72,In_948,In_757);
and U73 (N_73,In_405,In_314);
xnor U74 (N_74,In_788,In_262);
xnor U75 (N_75,In_219,In_399);
nor U76 (N_76,In_860,In_696);
nand U77 (N_77,In_723,In_878);
or U78 (N_78,In_106,In_610);
or U79 (N_79,In_248,In_366);
nor U80 (N_80,In_463,In_152);
xor U81 (N_81,In_233,In_736);
and U82 (N_82,In_373,In_519);
nand U83 (N_83,In_121,In_715);
or U84 (N_84,In_603,In_543);
or U85 (N_85,In_952,In_783);
nor U86 (N_86,In_827,In_448);
and U87 (N_87,In_61,In_216);
nand U88 (N_88,In_717,In_253);
or U89 (N_89,In_302,In_893);
or U90 (N_90,In_85,In_428);
xor U91 (N_91,In_682,In_532);
nand U92 (N_92,In_59,In_29);
nand U93 (N_93,In_458,In_982);
and U94 (N_94,In_28,In_693);
nor U95 (N_95,In_648,In_522);
and U96 (N_96,In_72,In_276);
nand U97 (N_97,In_658,In_542);
nor U98 (N_98,In_83,In_383);
or U99 (N_99,In_69,In_983);
or U100 (N_100,In_583,In_854);
nor U101 (N_101,In_821,In_55);
or U102 (N_102,In_151,In_466);
or U103 (N_103,In_642,In_628);
nand U104 (N_104,In_962,In_586);
or U105 (N_105,In_178,In_556);
or U106 (N_106,In_320,In_229);
or U107 (N_107,In_475,In_547);
nand U108 (N_108,In_305,In_646);
nor U109 (N_109,In_263,In_911);
nand U110 (N_110,In_143,In_241);
nor U111 (N_111,In_445,In_741);
or U112 (N_112,In_131,In_395);
xnor U113 (N_113,In_386,In_292);
nor U114 (N_114,In_614,In_407);
nand U115 (N_115,In_677,In_382);
nor U116 (N_116,In_269,In_857);
nor U117 (N_117,In_485,In_401);
nand U118 (N_118,In_461,In_165);
or U119 (N_119,In_280,In_156);
or U120 (N_120,In_739,In_758);
or U121 (N_121,In_823,In_815);
nor U122 (N_122,In_589,In_661);
nor U123 (N_123,In_166,In_848);
or U124 (N_124,In_254,In_453);
xnor U125 (N_125,In_370,In_60);
or U126 (N_126,In_703,In_987);
nand U127 (N_127,In_527,In_968);
nand U128 (N_128,In_800,In_246);
nand U129 (N_129,In_790,In_297);
or U130 (N_130,In_958,In_585);
and U131 (N_131,In_594,In_468);
nand U132 (N_132,In_616,In_431);
nor U133 (N_133,In_692,In_766);
xor U134 (N_134,In_579,In_643);
nor U135 (N_135,In_444,In_832);
and U136 (N_136,In_311,In_78);
xnor U137 (N_137,In_487,In_46);
or U138 (N_138,In_372,In_325);
nor U139 (N_139,In_255,In_943);
nand U140 (N_140,In_19,In_173);
nor U141 (N_141,In_632,In_432);
nor U142 (N_142,In_339,In_763);
nor U143 (N_143,In_222,In_437);
xnor U144 (N_144,In_799,In_361);
or U145 (N_145,In_318,In_592);
xor U146 (N_146,In_136,In_455);
or U147 (N_147,In_48,In_611);
nor U148 (N_148,In_306,In_438);
nand U149 (N_149,In_819,In_540);
nor U150 (N_150,In_601,In_922);
nand U151 (N_151,In_479,In_1);
nor U152 (N_152,In_737,In_36);
and U153 (N_153,In_450,In_198);
or U154 (N_154,In_49,In_34);
and U155 (N_155,In_378,In_12);
or U156 (N_156,In_313,In_67);
nor U157 (N_157,In_371,In_869);
or U158 (N_158,In_294,In_811);
and U159 (N_159,In_240,In_282);
nand U160 (N_160,In_587,In_283);
and U161 (N_161,In_925,In_550);
nand U162 (N_162,In_187,In_804);
nor U163 (N_163,In_731,In_593);
or U164 (N_164,In_836,In_335);
nand U165 (N_165,In_633,In_257);
nand U166 (N_166,In_729,In_627);
or U167 (N_167,In_630,In_825);
nor U168 (N_168,In_886,In_621);
nand U169 (N_169,In_826,In_147);
nor U170 (N_170,In_898,In_882);
and U171 (N_171,In_533,In_876);
nor U172 (N_172,In_493,In_805);
or U173 (N_173,In_489,In_705);
or U174 (N_174,In_904,In_289);
xor U175 (N_175,In_414,In_186);
and U176 (N_176,In_180,In_285);
and U177 (N_177,In_488,In_913);
nor U178 (N_178,In_700,In_901);
nor U179 (N_179,In_308,In_234);
or U180 (N_180,In_363,In_337);
and U181 (N_181,In_317,In_416);
and U182 (N_182,In_607,In_900);
nor U183 (N_183,In_244,In_524);
and U184 (N_184,In_517,In_473);
and U185 (N_185,In_284,In_350);
nand U186 (N_186,In_921,In_761);
or U187 (N_187,In_954,In_743);
nor U188 (N_188,In_410,In_964);
nand U189 (N_189,In_107,In_797);
or U190 (N_190,In_135,In_668);
or U191 (N_191,In_970,In_423);
or U192 (N_192,In_531,In_406);
nand U193 (N_193,In_785,In_51);
and U194 (N_194,In_612,In_912);
xor U195 (N_195,In_230,In_833);
nand U196 (N_196,In_841,In_82);
nor U197 (N_197,In_567,In_529);
nor U198 (N_198,In_734,In_44);
or U199 (N_199,In_231,In_396);
nand U200 (N_200,In_118,N_7);
and U201 (N_201,In_196,In_427);
nand U202 (N_202,In_167,In_224);
nand U203 (N_203,N_31,N_22);
or U204 (N_204,N_43,N_185);
and U205 (N_205,N_4,In_974);
and U206 (N_206,In_574,In_936);
nor U207 (N_207,In_769,In_851);
xor U208 (N_208,In_345,In_287);
xor U209 (N_209,In_516,In_765);
and U210 (N_210,N_118,In_54);
nand U211 (N_211,In_940,In_581);
and U212 (N_212,In_58,In_683);
and U213 (N_213,In_80,In_546);
nor U214 (N_214,N_18,In_738);
nand U215 (N_215,In_862,In_637);
nor U216 (N_216,In_140,In_120);
nand U217 (N_217,In_62,In_42);
nand U218 (N_218,N_75,In_938);
or U219 (N_219,In_708,In_659);
xor U220 (N_220,In_247,N_35);
or U221 (N_221,N_70,In_368);
nand U222 (N_222,In_865,In_640);
and U223 (N_223,In_780,N_105);
xnor U224 (N_224,N_110,In_33);
nand U225 (N_225,N_71,In_965);
nor U226 (N_226,In_946,In_75);
nand U227 (N_227,In_133,In_673);
nor U228 (N_228,In_852,In_30);
nand U229 (N_229,In_429,In_873);
and U230 (N_230,N_25,In_102);
nand U231 (N_231,In_137,In_992);
and U232 (N_232,In_934,In_500);
or U233 (N_233,N_50,N_122);
nor U234 (N_234,N_95,N_147);
or U235 (N_235,In_171,N_30);
or U236 (N_236,In_275,In_90);
or U237 (N_237,In_393,N_170);
nand U238 (N_238,N_26,In_273);
or U239 (N_239,In_338,In_669);
or U240 (N_240,In_433,In_93);
xnor U241 (N_241,N_183,In_772);
or U242 (N_242,In_570,In_460);
or U243 (N_243,In_63,In_387);
xor U244 (N_244,In_663,In_784);
nand U245 (N_245,In_636,In_181);
or U246 (N_246,N_103,In_651);
or U247 (N_247,In_575,In_483);
xor U248 (N_248,N_161,In_41);
and U249 (N_249,In_111,In_980);
nand U250 (N_250,In_713,N_186);
or U251 (N_251,In_122,In_565);
nand U252 (N_252,In_202,In_679);
and U253 (N_253,In_312,In_474);
nand U254 (N_254,In_989,In_144);
or U255 (N_255,In_675,In_351);
and U256 (N_256,In_464,In_115);
nor U257 (N_257,N_16,In_245);
and U258 (N_258,In_125,In_191);
xor U259 (N_259,In_123,In_443);
and U260 (N_260,In_796,In_674);
or U261 (N_261,N_188,In_14);
or U262 (N_262,In_792,In_650);
nand U263 (N_263,In_718,In_591);
nand U264 (N_264,In_732,N_44);
nor U265 (N_265,N_139,In_928);
nor U266 (N_266,N_117,In_18);
or U267 (N_267,N_116,In_250);
or U268 (N_268,N_97,In_771);
nand U269 (N_269,In_839,In_695);
or U270 (N_270,In_348,N_175);
and U271 (N_271,In_595,In_710);
xor U272 (N_272,In_625,In_808);
or U273 (N_273,N_143,In_874);
xor U274 (N_274,N_135,In_963);
nor U275 (N_275,In_490,N_58);
xnor U276 (N_276,In_844,In_923);
and U277 (N_277,In_355,N_166);
nor U278 (N_278,In_988,In_128);
and U279 (N_279,In_973,In_272);
xnor U280 (N_280,In_930,N_160);
nand U281 (N_281,N_190,In_507);
nand U282 (N_282,In_199,In_367);
nand U283 (N_283,In_6,In_8);
or U284 (N_284,In_195,N_77);
nand U285 (N_285,In_146,In_806);
nand U286 (N_286,In_711,N_67);
xor U287 (N_287,In_74,In_545);
nand U288 (N_288,In_426,In_716);
nand U289 (N_289,In_641,In_92);
or U290 (N_290,In_486,N_114);
and U291 (N_291,In_81,In_15);
or U292 (N_292,N_61,In_20);
or U293 (N_293,In_304,In_494);
and U294 (N_294,In_190,In_829);
and U295 (N_295,In_793,N_191);
and U296 (N_296,In_446,In_484);
and U297 (N_297,In_235,In_662);
and U298 (N_298,In_492,N_72);
and U299 (N_299,In_391,In_976);
or U300 (N_300,In_476,In_113);
nor U301 (N_301,In_508,In_727);
xor U302 (N_302,N_151,N_112);
nand U303 (N_303,N_146,In_495);
or U304 (N_304,N_179,N_163);
nor U305 (N_305,In_604,In_867);
and U306 (N_306,In_497,In_528);
nor U307 (N_307,In_185,In_377);
nor U308 (N_308,In_316,In_947);
nor U309 (N_309,N_76,In_357);
nor U310 (N_310,In_961,In_950);
nand U311 (N_311,In_905,In_45);
xnor U312 (N_312,In_597,N_49);
nand U313 (N_313,In_271,In_268);
nand U314 (N_314,In_984,In_812);
or U315 (N_315,In_380,In_237);
and U316 (N_316,In_478,In_261);
nand U317 (N_317,N_40,N_140);
nand U318 (N_318,In_303,In_649);
or U319 (N_319,In_177,N_193);
nand U320 (N_320,In_801,In_467);
and U321 (N_321,In_129,In_949);
and U322 (N_322,In_290,In_724);
or U323 (N_323,N_159,In_560);
nand U324 (N_324,In_481,N_167);
nand U325 (N_325,In_755,In_782);
or U326 (N_326,In_760,In_232);
and U327 (N_327,In_667,In_795);
nand U328 (N_328,In_599,In_105);
nand U329 (N_329,In_813,N_59);
and U330 (N_330,N_73,In_721);
and U331 (N_331,N_198,N_158);
or U332 (N_332,In_207,In_820);
and U333 (N_333,N_144,In_236);
and U334 (N_334,In_293,In_789);
nand U335 (N_335,In_910,In_704);
nand U336 (N_336,In_941,In_439);
nor U337 (N_337,In_510,In_134);
nor U338 (N_338,In_116,In_847);
nand U339 (N_339,In_566,N_56);
xnor U340 (N_340,In_220,N_38);
or U341 (N_341,In_145,N_150);
and U342 (N_342,In_65,In_990);
or U343 (N_343,In_807,In_559);
nor U344 (N_344,In_435,In_759);
nand U345 (N_345,N_94,In_605);
xor U346 (N_346,In_518,In_319);
or U347 (N_347,In_885,In_620);
nand U348 (N_348,In_477,In_326);
and U349 (N_349,In_887,N_194);
and U350 (N_350,In_600,In_824);
nor U351 (N_351,In_850,In_877);
or U352 (N_352,In_786,In_746);
and U353 (N_353,In_141,In_267);
xor U354 (N_354,N_173,In_96);
nand U355 (N_355,In_748,In_975);
or U356 (N_356,N_102,N_87);
and U357 (N_357,In_505,In_9);
and U358 (N_358,In_513,In_182);
or U359 (N_359,In_548,In_323);
or U360 (N_360,In_684,N_145);
nand U361 (N_361,In_24,In_834);
and U362 (N_362,N_45,In_309);
or U363 (N_363,N_109,In_534);
nand U364 (N_364,In_310,In_944);
or U365 (N_365,In_328,N_187);
or U366 (N_366,In_170,In_972);
xor U367 (N_367,In_747,N_164);
and U368 (N_368,In_442,In_472);
nand U369 (N_369,In_501,In_764);
or U370 (N_370,In_206,In_881);
nand U371 (N_371,In_159,N_184);
nor U372 (N_372,In_698,In_164);
nor U373 (N_373,In_756,N_171);
nor U374 (N_374,In_117,In_266);
and U375 (N_375,N_99,In_470);
and U376 (N_376,In_535,N_123);
nand U377 (N_377,In_94,N_182);
or U378 (N_378,N_64,In_112);
or U379 (N_379,In_184,In_809);
nand U380 (N_380,N_168,In_110);
or U381 (N_381,In_449,N_17);
nand U382 (N_382,N_127,In_340);
and U383 (N_383,N_42,N_81);
xor U384 (N_384,In_25,N_93);
nand U385 (N_385,In_324,In_336);
or U386 (N_386,In_5,In_142);
nor U387 (N_387,In_203,In_157);
and U388 (N_388,N_189,In_441);
xnor U389 (N_389,In_557,In_97);
xnor U390 (N_390,In_767,In_840);
and U391 (N_391,In_179,In_103);
and U392 (N_392,N_142,In_932);
xor U393 (N_393,In_896,In_670);
nor U394 (N_394,In_176,In_189);
and U395 (N_395,In_863,In_126);
nor U396 (N_396,In_699,N_12);
nand U397 (N_397,In_153,In_831);
and U398 (N_398,In_421,In_552);
and U399 (N_399,In_571,In_39);
and U400 (N_400,N_275,N_126);
nand U401 (N_401,In_37,In_880);
or U402 (N_402,N_19,N_259);
and U403 (N_403,In_197,N_291);
and U404 (N_404,N_201,In_719);
nor U405 (N_405,N_236,In_895);
and U406 (N_406,In_866,N_215);
and U407 (N_407,In_787,N_232);
nand U408 (N_408,In_523,In_915);
nand U409 (N_409,N_258,In_776);
and U410 (N_410,N_233,N_227);
and U411 (N_411,N_218,N_51);
or U412 (N_412,In_871,N_383);
and U413 (N_413,N_263,N_338);
nor U414 (N_414,N_245,N_148);
and U415 (N_415,N_226,In_506);
and U416 (N_416,In_929,In_872);
nor U417 (N_417,In_299,In_617);
nor U418 (N_418,N_69,In_935);
or U419 (N_419,N_389,In_859);
or U420 (N_420,N_14,N_52);
nor U421 (N_421,N_195,In_909);
nand U422 (N_422,N_362,In_100);
or U423 (N_423,N_261,In_544);
nor U424 (N_424,In_86,In_259);
and U425 (N_425,In_931,N_352);
or U426 (N_426,N_129,N_131);
or U427 (N_427,N_107,N_152);
xnor U428 (N_428,N_269,N_172);
nand U429 (N_429,N_321,In_584);
or U430 (N_430,In_193,N_176);
or U431 (N_431,N_20,N_279);
or U432 (N_432,In_977,N_228);
or U433 (N_433,In_346,In_419);
or U434 (N_434,N_369,N_339);
nand U435 (N_435,N_244,N_331);
xor U436 (N_436,In_889,In_349);
nand U437 (N_437,In_201,In_861);
nor U438 (N_438,N_390,N_346);
and U439 (N_439,N_222,N_386);
nand U440 (N_440,N_378,In_150);
or U441 (N_441,N_395,In_775);
xor U442 (N_442,N_124,In_260);
nor U443 (N_443,N_260,N_305);
xnor U444 (N_444,In_482,N_157);
or U445 (N_445,N_192,N_250);
nand U446 (N_446,N_1,N_231);
and U447 (N_447,N_276,In_307);
nand U448 (N_448,In_686,N_327);
nor U449 (N_449,In_496,N_128);
nand U450 (N_450,N_375,N_83);
nand U451 (N_451,In_555,In_215);
or U452 (N_452,In_322,In_953);
and U453 (N_453,N_13,In_754);
nand U454 (N_454,In_933,N_221);
and U455 (N_455,N_224,N_11);
xor U456 (N_456,N_80,In_530);
nand U457 (N_457,N_48,In_596);
nor U458 (N_458,N_397,In_842);
nand U459 (N_459,In_409,N_210);
or U460 (N_460,In_71,N_8);
or U461 (N_461,N_57,N_169);
nand U462 (N_462,In_653,In_563);
nand U463 (N_463,N_46,In_572);
nor U464 (N_464,In_551,In_127);
nand U465 (N_465,In_569,N_391);
and U466 (N_466,In_375,N_205);
nand U467 (N_467,N_308,N_377);
or U468 (N_468,In_919,In_465);
nand U469 (N_469,In_239,N_86);
and U470 (N_470,N_138,N_319);
nand U471 (N_471,In_689,N_197);
nand U472 (N_472,N_24,In_329);
or U473 (N_473,N_262,In_957);
nand U474 (N_474,In_411,N_65);
or U475 (N_475,In_38,N_312);
and U476 (N_476,N_396,In_856);
or U477 (N_477,N_322,In_908);
or U478 (N_478,N_3,In_981);
nor U479 (N_479,N_91,N_254);
xor U480 (N_480,N_208,In_762);
xnor U481 (N_481,In_907,N_399);
or U482 (N_482,N_180,In_27);
or U483 (N_483,In_161,N_302);
nand U484 (N_484,N_363,In_436);
nand U485 (N_485,N_253,N_341);
xnor U486 (N_486,N_287,In_752);
or U487 (N_487,In_937,In_403);
nand U488 (N_488,N_177,N_199);
xor U489 (N_489,In_902,N_246);
and U490 (N_490,N_303,In_791);
nor U491 (N_491,N_353,In_422);
and U492 (N_492,In_678,N_130);
and U493 (N_493,In_918,In_822);
or U494 (N_494,N_304,N_241);
or U495 (N_495,N_153,In_291);
nand U496 (N_496,N_256,In_194);
nand U497 (N_497,N_394,N_360);
or U498 (N_498,N_273,N_267);
xor U499 (N_499,In_979,N_92);
nand U500 (N_500,In_694,In_163);
or U501 (N_501,N_337,In_258);
nand U502 (N_502,In_511,N_90);
xor U503 (N_503,In_369,In_343);
nand U504 (N_504,In_32,In_360);
and U505 (N_505,In_688,In_217);
xor U506 (N_506,N_379,In_687);
and U507 (N_507,In_916,In_454);
nor U508 (N_508,In_735,In_740);
and U509 (N_509,In_256,In_226);
and U510 (N_510,In_883,In_296);
xor U511 (N_511,In_452,In_327);
xnor U512 (N_512,In_251,In_994);
nor U513 (N_513,In_400,In_175);
xor U514 (N_514,In_227,In_562);
and U515 (N_515,N_320,N_243);
and U516 (N_516,N_342,N_108);
nor U517 (N_517,In_588,In_660);
or U518 (N_518,N_156,N_230);
nor U519 (N_519,N_100,N_47);
or U520 (N_520,In_480,N_217);
xnor U521 (N_521,N_340,In_381);
or U522 (N_522,N_272,N_332);
nand U523 (N_523,N_211,In_208);
nor U524 (N_524,In_456,N_311);
nand U525 (N_525,N_121,N_149);
or U526 (N_526,N_125,N_137);
or U527 (N_527,N_364,N_10);
or U528 (N_528,In_971,In_998);
or U529 (N_529,In_779,N_21);
and U530 (N_530,N_181,In_286);
or U531 (N_531,N_355,In_701);
xnor U532 (N_532,In_749,N_292);
xnor U533 (N_533,In_252,In_130);
or U534 (N_534,N_301,N_132);
xor U535 (N_535,N_225,In_602);
or U536 (N_536,N_219,N_203);
and U537 (N_537,In_119,In_64);
nor U538 (N_538,N_5,N_27);
nor U539 (N_539,In_835,In_818);
or U540 (N_540,In_773,In_794);
nand U541 (N_541,N_0,In_413);
nor U542 (N_542,N_174,In_192);
or U543 (N_543,In_726,N_101);
and U544 (N_544,In_77,N_111);
nand U545 (N_545,In_76,In_635);
xnor U546 (N_546,In_666,In_714);
nor U547 (N_547,In_392,In_228);
or U548 (N_548,N_285,N_133);
and U549 (N_549,N_372,In_447);
nor U550 (N_550,N_325,N_336);
xor U551 (N_551,N_238,In_408);
or U552 (N_552,N_380,N_104);
and U553 (N_553,N_89,N_209);
nand U554 (N_554,In_843,In_993);
xnor U555 (N_555,N_206,In_514);
or U556 (N_556,N_293,N_74);
or U557 (N_557,N_78,In_35);
xor U558 (N_558,N_264,In_680);
nand U559 (N_559,N_34,N_376);
or U560 (N_560,In_16,In_356);
or U561 (N_561,In_3,N_289);
nor U562 (N_562,N_357,In_434);
nand U563 (N_563,N_366,N_265);
xor U564 (N_564,In_47,In_685);
and U565 (N_565,In_914,N_365);
nand U566 (N_566,N_317,N_315);
nand U567 (N_567,In_837,N_286);
xor U568 (N_568,N_358,N_324);
and U569 (N_569,N_370,In_690);
nand U570 (N_570,N_15,N_96);
and U571 (N_571,N_310,In_985);
or U572 (N_572,In_996,In_101);
nor U573 (N_573,N_334,In_174);
and U574 (N_574,In_553,In_951);
nor U575 (N_575,N_297,In_967);
nand U576 (N_576,N_384,In_200);
nand U577 (N_577,In_564,N_344);
nand U578 (N_578,In_816,N_278);
nor U579 (N_579,In_722,N_242);
or U580 (N_580,In_504,In_515);
nor U581 (N_581,N_2,N_326);
nor U582 (N_582,N_234,In_344);
nor U583 (N_583,N_354,In_745);
xor U584 (N_584,In_491,In_639);
nor U585 (N_585,N_212,In_849);
nor U586 (N_586,N_202,In_160);
nor U587 (N_587,N_252,In_353);
and U588 (N_588,N_361,In_278);
nand U589 (N_589,In_654,N_141);
or U590 (N_590,In_526,In_676);
or U591 (N_591,N_300,N_313);
nor U592 (N_592,In_238,N_39);
nand U593 (N_593,N_120,N_359);
xnor U594 (N_594,In_626,In_652);
and U595 (N_595,N_374,N_204);
nand U596 (N_596,In_288,In_997);
nand U597 (N_597,N_398,N_290);
nand U598 (N_598,N_79,In_750);
xnor U599 (N_599,N_367,In_709);
nand U600 (N_600,In_188,N_460);
xor U601 (N_601,N_248,N_486);
nor U602 (N_602,N_569,N_540);
and U603 (N_603,N_330,In_590);
nand U604 (N_604,In_204,In_609);
and U605 (N_605,N_510,N_54);
xnor U606 (N_606,N_583,N_554);
nor U607 (N_607,N_6,N_519);
or U608 (N_608,N_373,N_425);
nand U609 (N_609,N_527,In_138);
nand U610 (N_610,In_213,In_656);
or U611 (N_611,N_520,N_501);
and U612 (N_612,N_472,N_473);
or U613 (N_613,N_277,N_490);
or U614 (N_614,N_282,N_483);
xnor U615 (N_615,N_284,N_409);
nor U616 (N_616,N_596,N_451);
nand U617 (N_617,N_539,In_598);
nor U618 (N_618,N_270,N_573);
nor U619 (N_619,N_523,N_434);
xnor U620 (N_620,In_168,N_500);
nand U621 (N_621,N_442,N_387);
nand U622 (N_622,N_200,N_400);
nor U623 (N_623,N_240,N_590);
or U624 (N_624,N_466,N_33);
or U625 (N_625,N_478,N_298);
and U626 (N_626,N_538,N_588);
nand U627 (N_627,N_423,N_555);
nand U628 (N_628,N_251,N_410);
and U629 (N_629,N_463,In_802);
and U630 (N_630,N_512,N_504);
or U631 (N_631,N_599,In_956);
nand U632 (N_632,N_445,N_446);
nor U633 (N_633,N_29,N_552);
or U634 (N_634,N_511,N_561);
xor U635 (N_635,N_577,N_514);
xor U636 (N_636,N_481,In_777);
xnor U637 (N_637,In_884,N_494);
nand U638 (N_638,In_11,N_407);
or U639 (N_639,N_579,In_582);
and U640 (N_640,N_348,N_581);
nand U641 (N_641,N_522,N_411);
and U642 (N_642,N_487,In_608);
nand U643 (N_643,N_543,In_868);
and U644 (N_644,N_274,N_480);
or U645 (N_645,N_485,N_491);
nor U646 (N_646,In_702,N_586);
or U647 (N_647,N_424,N_382);
and U648 (N_648,In_845,N_84);
nor U649 (N_649,N_207,In_424);
nor U650 (N_650,N_271,N_448);
and U651 (N_651,N_414,In_742);
nand U652 (N_652,In_10,N_592);
nor U653 (N_653,In_720,N_517);
xor U654 (N_654,N_558,N_568);
or U655 (N_655,N_461,N_484);
or U656 (N_656,In_521,N_385);
or U657 (N_657,In_512,N_439);
and U658 (N_658,N_492,In_315);
and U659 (N_659,N_443,N_235);
nor U660 (N_660,N_318,N_476);
nor U661 (N_661,N_593,N_280);
and U662 (N_662,N_532,N_597);
or U663 (N_663,N_531,In_52);
nand U664 (N_664,In_744,N_63);
or U665 (N_665,In_398,In_388);
or U666 (N_666,In_321,In_875);
and U667 (N_667,N_408,N_493);
or U668 (N_668,N_462,N_413);
and U669 (N_669,In_538,N_415);
or U670 (N_670,In_753,N_82);
nand U671 (N_671,N_429,In_79);
or U672 (N_672,N_541,N_66);
nor U673 (N_673,N_165,N_60);
xnor U674 (N_674,In_104,N_388);
nor U675 (N_675,N_328,N_41);
or U676 (N_676,N_450,N_566);
nor U677 (N_677,N_247,N_371);
nand U678 (N_678,In_379,N_314);
or U679 (N_679,In_430,N_316);
or U680 (N_680,N_406,In_281);
and U681 (N_681,N_55,N_495);
nand U682 (N_682,In_412,In_838);
nor U683 (N_683,N_594,N_582);
nor U684 (N_684,N_136,In_397);
nor U685 (N_685,N_106,In_580);
nor U686 (N_686,In_814,N_268);
and U687 (N_687,N_421,In_214);
and U688 (N_688,N_435,N_575);
and U689 (N_689,N_530,N_468);
or U690 (N_690,In_279,N_437);
nor U691 (N_691,N_323,N_513);
and U692 (N_692,N_589,N_598);
nand U693 (N_693,In_223,N_266);
and U694 (N_694,N_556,N_550);
xor U695 (N_695,N_562,N_62);
nor U696 (N_696,In_655,In_622);
nand U697 (N_697,N_440,In_451);
nor U698 (N_698,N_405,In_920);
or U699 (N_699,N_349,N_426);
nor U700 (N_700,N_452,N_119);
or U701 (N_701,N_419,N_470);
nand U702 (N_702,In_502,In_966);
nand U703 (N_703,N_237,In_417);
and U704 (N_704,N_155,In_817);
nor U705 (N_705,In_40,N_574);
nand U706 (N_706,N_294,N_546);
and U707 (N_707,In_576,In_221);
nor U708 (N_708,In_43,In_672);
and U709 (N_709,N_518,N_23);
nand U710 (N_710,In_733,N_553);
nand U711 (N_711,N_489,N_515);
xor U712 (N_712,N_503,N_335);
or U713 (N_713,In_537,N_565);
nor U714 (N_714,N_548,N_420);
and U715 (N_715,N_496,In_615);
or U716 (N_716,N_459,In_425);
nor U717 (N_717,N_239,N_393);
xnor U718 (N_718,In_155,N_528);
nand U719 (N_719,N_392,N_416);
xnor U720 (N_720,In_986,N_436);
or U721 (N_721,N_433,N_549);
nand U722 (N_722,N_438,N_220);
nor U723 (N_723,N_526,N_457);
nor U724 (N_724,N_368,N_585);
nand U725 (N_725,N_505,N_113);
nand U726 (N_726,N_535,N_295);
and U727 (N_727,N_281,In_70);
or U728 (N_728,N_557,N_32);
or U729 (N_729,In_205,In_539);
or U730 (N_730,N_288,N_509);
xor U731 (N_731,N_402,N_524);
xnor U732 (N_732,N_255,N_283);
or U733 (N_733,N_453,In_631);
and U734 (N_734,In_577,N_544);
nor U735 (N_735,N_196,N_533);
nand U736 (N_736,N_403,N_563);
nor U737 (N_737,N_595,N_422);
nand U738 (N_738,In_23,In_803);
nor U739 (N_739,N_477,N_551);
nor U740 (N_740,N_497,N_455);
and U741 (N_741,N_85,N_257);
or U742 (N_742,N_28,N_449);
nand U743 (N_743,N_537,N_345);
or U744 (N_744,N_329,In_897);
and U745 (N_745,N_68,N_229);
or U746 (N_746,N_506,N_430);
nand U747 (N_747,N_428,N_115);
nand U748 (N_748,N_564,N_567);
nor U749 (N_749,N_214,In_139);
nand U750 (N_750,In_17,N_525);
nor U751 (N_751,N_508,N_499);
nor U752 (N_752,N_333,N_482);
or U753 (N_753,N_444,In_558);
and U754 (N_754,In_415,In_99);
xor U755 (N_755,N_521,In_13);
nor U756 (N_756,N_572,N_474);
nor U757 (N_757,N_296,N_507);
and U758 (N_758,In_999,In_855);
or U759 (N_759,In_158,N_576);
nor U760 (N_760,N_465,N_178);
nor U761 (N_761,N_9,N_134);
nand U762 (N_762,N_587,In_358);
or U763 (N_763,N_223,N_356);
nand U764 (N_764,N_427,N_580);
nor U765 (N_765,N_307,N_417);
xor U766 (N_766,In_218,N_570);
nand U767 (N_767,N_454,In_568);
and U768 (N_768,N_542,In_352);
and U769 (N_769,N_404,N_547);
nand U770 (N_770,N_464,N_432);
and U771 (N_771,N_216,N_498);
or U772 (N_772,N_98,N_213);
nand U773 (N_773,In_778,N_591);
nand U774 (N_774,N_502,N_571);
or U775 (N_775,N_381,In_402);
nor U776 (N_776,N_343,N_469);
nand U777 (N_777,N_559,N_441);
or U778 (N_778,N_471,In_341);
nand U779 (N_779,N_309,N_401);
xnor U780 (N_780,In_619,N_351);
nor U781 (N_781,N_529,N_475);
nand U782 (N_782,N_306,N_456);
nand U783 (N_783,N_578,In_509);
or U784 (N_784,In_525,In_665);
or U785 (N_785,N_431,In_132);
or U786 (N_786,N_53,N_447);
or U787 (N_787,N_347,N_479);
nand U788 (N_788,In_7,N_458);
nand U789 (N_789,N_488,N_249);
nand U790 (N_790,N_299,N_536);
xor U791 (N_791,N_560,N_37);
nor U792 (N_792,In_707,N_467);
or U793 (N_793,N_162,N_584);
nand U794 (N_794,N_418,In_671);
and U795 (N_795,N_534,N_154);
nor U796 (N_796,N_36,N_350);
and U797 (N_797,In_499,N_88);
or U798 (N_798,In_89,N_412);
and U799 (N_799,N_545,N_516);
xnor U800 (N_800,N_713,N_608);
or U801 (N_801,N_790,N_648);
and U802 (N_802,N_634,N_653);
and U803 (N_803,N_787,N_646);
nand U804 (N_804,N_728,N_707);
xnor U805 (N_805,N_665,N_690);
nand U806 (N_806,N_610,N_701);
or U807 (N_807,N_737,N_699);
or U808 (N_808,N_775,N_606);
and U809 (N_809,N_745,N_674);
nor U810 (N_810,N_658,N_789);
and U811 (N_811,N_672,N_709);
or U812 (N_812,N_733,N_666);
or U813 (N_813,N_786,N_760);
nor U814 (N_814,N_623,N_627);
nor U815 (N_815,N_630,N_724);
or U816 (N_816,N_652,N_732);
or U817 (N_817,N_711,N_720);
and U818 (N_818,N_761,N_619);
and U819 (N_819,N_793,N_773);
and U820 (N_820,N_697,N_643);
xnor U821 (N_821,N_651,N_694);
nor U822 (N_822,N_647,N_783);
nor U823 (N_823,N_788,N_785);
nor U824 (N_824,N_691,N_603);
or U825 (N_825,N_784,N_675);
nand U826 (N_826,N_611,N_725);
or U827 (N_827,N_659,N_722);
xnor U828 (N_828,N_750,N_680);
xor U829 (N_829,N_792,N_695);
and U830 (N_830,N_799,N_747);
or U831 (N_831,N_729,N_777);
nor U832 (N_832,N_757,N_769);
nor U833 (N_833,N_657,N_686);
xnor U834 (N_834,N_614,N_743);
nand U835 (N_835,N_748,N_764);
and U836 (N_836,N_628,N_708);
or U837 (N_837,N_780,N_735);
nor U838 (N_838,N_626,N_719);
or U839 (N_839,N_604,N_684);
or U840 (N_840,N_796,N_736);
or U841 (N_841,N_681,N_758);
nor U842 (N_842,N_734,N_704);
and U843 (N_843,N_678,N_727);
and U844 (N_844,N_640,N_632);
nor U845 (N_845,N_746,N_631);
nand U846 (N_846,N_609,N_739);
nor U847 (N_847,N_616,N_767);
or U848 (N_848,N_602,N_676);
or U849 (N_849,N_685,N_752);
nor U850 (N_850,N_638,N_782);
xor U851 (N_851,N_794,N_762);
or U852 (N_852,N_759,N_618);
or U853 (N_853,N_622,N_650);
or U854 (N_854,N_601,N_664);
nor U855 (N_855,N_677,N_741);
nand U856 (N_856,N_629,N_798);
nand U857 (N_857,N_714,N_781);
and U858 (N_858,N_765,N_740);
xnor U859 (N_859,N_772,N_776);
and U860 (N_860,N_703,N_742);
and U861 (N_861,N_755,N_668);
and U862 (N_862,N_661,N_687);
or U863 (N_863,N_669,N_730);
nand U864 (N_864,N_621,N_778);
and U865 (N_865,N_663,N_731);
or U866 (N_866,N_692,N_667);
nand U867 (N_867,N_607,N_637);
or U868 (N_868,N_797,N_771);
nor U869 (N_869,N_779,N_670);
and U870 (N_870,N_768,N_710);
nor U871 (N_871,N_744,N_749);
nand U872 (N_872,N_656,N_645);
or U873 (N_873,N_766,N_688);
nand U874 (N_874,N_624,N_620);
nand U875 (N_875,N_756,N_726);
or U876 (N_876,N_754,N_639);
nor U877 (N_877,N_721,N_615);
or U878 (N_878,N_612,N_649);
and U879 (N_879,N_683,N_642);
nor U880 (N_880,N_605,N_716);
or U881 (N_881,N_763,N_662);
or U882 (N_882,N_706,N_641);
and U883 (N_883,N_671,N_660);
or U884 (N_884,N_673,N_738);
nand U885 (N_885,N_700,N_774);
nor U886 (N_886,N_654,N_613);
nor U887 (N_887,N_717,N_753);
and U888 (N_888,N_617,N_689);
nand U889 (N_889,N_644,N_635);
xnor U890 (N_890,N_791,N_636);
nor U891 (N_891,N_693,N_705);
and U892 (N_892,N_718,N_600);
or U893 (N_893,N_751,N_712);
or U894 (N_894,N_698,N_679);
and U895 (N_895,N_770,N_625);
and U896 (N_896,N_795,N_715);
and U897 (N_897,N_696,N_723);
nand U898 (N_898,N_655,N_682);
nand U899 (N_899,N_702,N_633);
or U900 (N_900,N_785,N_673);
and U901 (N_901,N_791,N_752);
xor U902 (N_902,N_726,N_682);
nor U903 (N_903,N_753,N_794);
nand U904 (N_904,N_743,N_682);
and U905 (N_905,N_690,N_626);
xnor U906 (N_906,N_609,N_799);
or U907 (N_907,N_704,N_612);
nand U908 (N_908,N_786,N_652);
and U909 (N_909,N_765,N_705);
and U910 (N_910,N_637,N_729);
and U911 (N_911,N_602,N_610);
or U912 (N_912,N_629,N_792);
and U913 (N_913,N_652,N_708);
or U914 (N_914,N_786,N_635);
nor U915 (N_915,N_602,N_603);
and U916 (N_916,N_740,N_600);
nand U917 (N_917,N_657,N_795);
nor U918 (N_918,N_797,N_639);
nand U919 (N_919,N_772,N_662);
nand U920 (N_920,N_753,N_788);
and U921 (N_921,N_713,N_755);
nor U922 (N_922,N_608,N_670);
or U923 (N_923,N_702,N_767);
nand U924 (N_924,N_674,N_619);
nand U925 (N_925,N_751,N_704);
nand U926 (N_926,N_677,N_783);
and U927 (N_927,N_718,N_770);
or U928 (N_928,N_633,N_635);
xnor U929 (N_929,N_711,N_773);
and U930 (N_930,N_731,N_675);
or U931 (N_931,N_710,N_629);
nor U932 (N_932,N_794,N_667);
or U933 (N_933,N_626,N_752);
nor U934 (N_934,N_699,N_690);
or U935 (N_935,N_654,N_678);
nand U936 (N_936,N_762,N_747);
and U937 (N_937,N_759,N_754);
nand U938 (N_938,N_766,N_730);
nand U939 (N_939,N_688,N_793);
xnor U940 (N_940,N_647,N_643);
or U941 (N_941,N_738,N_600);
nor U942 (N_942,N_792,N_666);
and U943 (N_943,N_794,N_602);
or U944 (N_944,N_684,N_719);
and U945 (N_945,N_703,N_667);
nor U946 (N_946,N_681,N_789);
nand U947 (N_947,N_600,N_673);
xnor U948 (N_948,N_601,N_672);
and U949 (N_949,N_649,N_629);
and U950 (N_950,N_691,N_703);
nand U951 (N_951,N_726,N_685);
nand U952 (N_952,N_701,N_707);
nor U953 (N_953,N_696,N_778);
or U954 (N_954,N_703,N_639);
or U955 (N_955,N_669,N_701);
nor U956 (N_956,N_709,N_669);
xnor U957 (N_957,N_771,N_709);
xnor U958 (N_958,N_779,N_648);
or U959 (N_959,N_656,N_753);
nor U960 (N_960,N_675,N_795);
or U961 (N_961,N_725,N_742);
nand U962 (N_962,N_649,N_687);
nand U963 (N_963,N_661,N_664);
or U964 (N_964,N_752,N_686);
or U965 (N_965,N_786,N_736);
nand U966 (N_966,N_669,N_613);
xor U967 (N_967,N_728,N_651);
or U968 (N_968,N_714,N_616);
or U969 (N_969,N_710,N_644);
or U970 (N_970,N_749,N_772);
nor U971 (N_971,N_782,N_680);
nor U972 (N_972,N_721,N_646);
nor U973 (N_973,N_718,N_737);
nand U974 (N_974,N_741,N_748);
or U975 (N_975,N_606,N_612);
nor U976 (N_976,N_609,N_719);
and U977 (N_977,N_700,N_765);
nand U978 (N_978,N_735,N_710);
or U979 (N_979,N_697,N_797);
nor U980 (N_980,N_727,N_751);
nor U981 (N_981,N_719,N_694);
and U982 (N_982,N_774,N_685);
nor U983 (N_983,N_738,N_724);
nor U984 (N_984,N_773,N_742);
nor U985 (N_985,N_621,N_646);
nand U986 (N_986,N_613,N_614);
or U987 (N_987,N_707,N_770);
nand U988 (N_988,N_632,N_624);
xnor U989 (N_989,N_710,N_663);
and U990 (N_990,N_715,N_769);
and U991 (N_991,N_788,N_692);
and U992 (N_992,N_734,N_611);
nand U993 (N_993,N_713,N_658);
or U994 (N_994,N_697,N_722);
or U995 (N_995,N_787,N_666);
nor U996 (N_996,N_722,N_711);
nand U997 (N_997,N_754,N_773);
nor U998 (N_998,N_610,N_638);
nor U999 (N_999,N_606,N_721);
or U1000 (N_1000,N_822,N_988);
and U1001 (N_1001,N_889,N_957);
or U1002 (N_1002,N_844,N_964);
xnor U1003 (N_1003,N_953,N_963);
nand U1004 (N_1004,N_854,N_909);
nand U1005 (N_1005,N_917,N_955);
nor U1006 (N_1006,N_873,N_939);
nor U1007 (N_1007,N_856,N_995);
or U1008 (N_1008,N_803,N_813);
and U1009 (N_1009,N_884,N_934);
and U1010 (N_1010,N_930,N_949);
or U1011 (N_1011,N_859,N_851);
or U1012 (N_1012,N_872,N_912);
nor U1013 (N_1013,N_970,N_935);
and U1014 (N_1014,N_863,N_877);
nor U1015 (N_1015,N_978,N_868);
and U1016 (N_1016,N_981,N_924);
or U1017 (N_1017,N_907,N_829);
or U1018 (N_1018,N_800,N_881);
and U1019 (N_1019,N_804,N_850);
nor U1020 (N_1020,N_918,N_911);
or U1021 (N_1021,N_897,N_853);
or U1022 (N_1022,N_842,N_906);
xor U1023 (N_1023,N_910,N_815);
and U1024 (N_1024,N_967,N_836);
nand U1025 (N_1025,N_893,N_885);
and U1026 (N_1026,N_802,N_807);
nand U1027 (N_1027,N_811,N_938);
or U1028 (N_1028,N_913,N_952);
nor U1029 (N_1029,N_847,N_867);
nor U1030 (N_1030,N_905,N_892);
and U1031 (N_1031,N_895,N_979);
xor U1032 (N_1032,N_834,N_846);
nand U1033 (N_1033,N_996,N_965);
or U1034 (N_1034,N_878,N_990);
or U1035 (N_1035,N_820,N_936);
or U1036 (N_1036,N_933,N_870);
xnor U1037 (N_1037,N_971,N_941);
nor U1038 (N_1038,N_968,N_886);
nand U1039 (N_1039,N_828,N_824);
or U1040 (N_1040,N_984,N_942);
and U1041 (N_1041,N_969,N_814);
or U1042 (N_1042,N_843,N_810);
and U1043 (N_1043,N_945,N_864);
nand U1044 (N_1044,N_901,N_931);
and U1045 (N_1045,N_992,N_899);
nand U1046 (N_1046,N_927,N_920);
or U1047 (N_1047,N_922,N_840);
nor U1048 (N_1048,N_919,N_801);
nand U1049 (N_1049,N_972,N_821);
or U1050 (N_1050,N_929,N_940);
nand U1051 (N_1051,N_923,N_977);
nor U1052 (N_1052,N_894,N_999);
xor U1053 (N_1053,N_947,N_986);
nor U1054 (N_1054,N_966,N_879);
nor U1055 (N_1055,N_830,N_944);
xnor U1056 (N_1056,N_812,N_914);
and U1057 (N_1057,N_874,N_982);
nor U1058 (N_1058,N_985,N_831);
nor U1059 (N_1059,N_862,N_825);
or U1060 (N_1060,N_816,N_852);
nor U1061 (N_1061,N_943,N_841);
xnor U1062 (N_1062,N_823,N_980);
nand U1063 (N_1063,N_950,N_860);
and U1064 (N_1064,N_805,N_908);
and U1065 (N_1065,N_926,N_875);
nand U1066 (N_1066,N_838,N_855);
nand U1067 (N_1067,N_991,N_809);
and U1068 (N_1068,N_898,N_975);
and U1069 (N_1069,N_989,N_900);
or U1070 (N_1070,N_951,N_865);
and U1071 (N_1071,N_983,N_976);
or U1072 (N_1072,N_904,N_994);
nor U1073 (N_1073,N_937,N_849);
and U1074 (N_1074,N_987,N_956);
xor U1075 (N_1075,N_880,N_890);
and U1076 (N_1076,N_959,N_876);
or U1077 (N_1077,N_848,N_818);
nor U1078 (N_1078,N_857,N_932);
nand U1079 (N_1079,N_946,N_998);
nor U1080 (N_1080,N_888,N_866);
nor U1081 (N_1081,N_961,N_835);
and U1082 (N_1082,N_858,N_887);
nand U1083 (N_1083,N_993,N_826);
or U1084 (N_1084,N_921,N_832);
and U1085 (N_1085,N_839,N_962);
xor U1086 (N_1086,N_861,N_837);
nand U1087 (N_1087,N_954,N_974);
or U1088 (N_1088,N_960,N_916);
or U1089 (N_1089,N_845,N_833);
and U1090 (N_1090,N_808,N_973);
nor U1091 (N_1091,N_903,N_928);
and U1092 (N_1092,N_869,N_997);
xor U1093 (N_1093,N_948,N_871);
nor U1094 (N_1094,N_882,N_958);
and U1095 (N_1095,N_817,N_925);
and U1096 (N_1096,N_891,N_827);
and U1097 (N_1097,N_819,N_902);
nor U1098 (N_1098,N_806,N_883);
xnor U1099 (N_1099,N_915,N_896);
xnor U1100 (N_1100,N_906,N_968);
nand U1101 (N_1101,N_817,N_864);
or U1102 (N_1102,N_848,N_878);
or U1103 (N_1103,N_922,N_890);
or U1104 (N_1104,N_895,N_994);
nand U1105 (N_1105,N_938,N_996);
nor U1106 (N_1106,N_803,N_808);
nor U1107 (N_1107,N_804,N_830);
nand U1108 (N_1108,N_914,N_827);
nor U1109 (N_1109,N_937,N_886);
nor U1110 (N_1110,N_938,N_857);
and U1111 (N_1111,N_809,N_995);
nand U1112 (N_1112,N_916,N_926);
xor U1113 (N_1113,N_945,N_950);
or U1114 (N_1114,N_937,N_823);
nor U1115 (N_1115,N_992,N_998);
nor U1116 (N_1116,N_995,N_816);
xnor U1117 (N_1117,N_873,N_945);
nand U1118 (N_1118,N_825,N_885);
nand U1119 (N_1119,N_835,N_980);
or U1120 (N_1120,N_894,N_992);
or U1121 (N_1121,N_876,N_974);
nor U1122 (N_1122,N_899,N_964);
nor U1123 (N_1123,N_980,N_902);
nand U1124 (N_1124,N_997,N_973);
nand U1125 (N_1125,N_914,N_883);
nor U1126 (N_1126,N_848,N_815);
and U1127 (N_1127,N_938,N_997);
nor U1128 (N_1128,N_910,N_801);
nor U1129 (N_1129,N_812,N_946);
and U1130 (N_1130,N_940,N_813);
nor U1131 (N_1131,N_814,N_914);
nor U1132 (N_1132,N_887,N_816);
nor U1133 (N_1133,N_825,N_849);
nor U1134 (N_1134,N_830,N_875);
and U1135 (N_1135,N_995,N_843);
or U1136 (N_1136,N_947,N_970);
nand U1137 (N_1137,N_981,N_849);
and U1138 (N_1138,N_808,N_993);
xor U1139 (N_1139,N_820,N_918);
nand U1140 (N_1140,N_925,N_932);
or U1141 (N_1141,N_816,N_891);
and U1142 (N_1142,N_857,N_870);
and U1143 (N_1143,N_888,N_971);
nor U1144 (N_1144,N_818,N_923);
or U1145 (N_1145,N_812,N_803);
nand U1146 (N_1146,N_872,N_891);
or U1147 (N_1147,N_965,N_820);
xnor U1148 (N_1148,N_858,N_840);
and U1149 (N_1149,N_956,N_884);
nor U1150 (N_1150,N_885,N_923);
and U1151 (N_1151,N_997,N_834);
or U1152 (N_1152,N_970,N_823);
nor U1153 (N_1153,N_924,N_867);
nand U1154 (N_1154,N_842,N_877);
or U1155 (N_1155,N_929,N_800);
or U1156 (N_1156,N_807,N_908);
xor U1157 (N_1157,N_881,N_882);
nor U1158 (N_1158,N_831,N_901);
xor U1159 (N_1159,N_923,N_893);
or U1160 (N_1160,N_984,N_979);
nor U1161 (N_1161,N_812,N_945);
nor U1162 (N_1162,N_863,N_996);
nand U1163 (N_1163,N_860,N_879);
nor U1164 (N_1164,N_829,N_821);
xnor U1165 (N_1165,N_876,N_948);
nor U1166 (N_1166,N_817,N_877);
or U1167 (N_1167,N_967,N_899);
nand U1168 (N_1168,N_864,N_998);
and U1169 (N_1169,N_828,N_948);
or U1170 (N_1170,N_970,N_882);
nand U1171 (N_1171,N_838,N_871);
nand U1172 (N_1172,N_840,N_998);
and U1173 (N_1173,N_802,N_867);
nand U1174 (N_1174,N_949,N_896);
nor U1175 (N_1175,N_810,N_978);
nor U1176 (N_1176,N_928,N_904);
or U1177 (N_1177,N_871,N_961);
or U1178 (N_1178,N_898,N_951);
or U1179 (N_1179,N_819,N_985);
or U1180 (N_1180,N_926,N_811);
nor U1181 (N_1181,N_870,N_830);
or U1182 (N_1182,N_918,N_881);
and U1183 (N_1183,N_862,N_997);
and U1184 (N_1184,N_934,N_966);
xor U1185 (N_1185,N_804,N_809);
and U1186 (N_1186,N_954,N_934);
nor U1187 (N_1187,N_881,N_887);
and U1188 (N_1188,N_921,N_893);
xor U1189 (N_1189,N_964,N_890);
nor U1190 (N_1190,N_888,N_944);
or U1191 (N_1191,N_931,N_993);
and U1192 (N_1192,N_944,N_850);
or U1193 (N_1193,N_953,N_834);
nand U1194 (N_1194,N_969,N_862);
nand U1195 (N_1195,N_888,N_917);
or U1196 (N_1196,N_839,N_904);
or U1197 (N_1197,N_999,N_961);
nand U1198 (N_1198,N_854,N_917);
nor U1199 (N_1199,N_828,N_991);
nor U1200 (N_1200,N_1159,N_1088);
nand U1201 (N_1201,N_1005,N_1051);
nand U1202 (N_1202,N_1151,N_1139);
nor U1203 (N_1203,N_1161,N_1099);
xnor U1204 (N_1204,N_1008,N_1022);
nand U1205 (N_1205,N_1020,N_1191);
xnor U1206 (N_1206,N_1030,N_1172);
or U1207 (N_1207,N_1169,N_1019);
and U1208 (N_1208,N_1187,N_1110);
nand U1209 (N_1209,N_1112,N_1186);
and U1210 (N_1210,N_1098,N_1055);
nor U1211 (N_1211,N_1084,N_1001);
nor U1212 (N_1212,N_1121,N_1115);
nand U1213 (N_1213,N_1081,N_1085);
and U1214 (N_1214,N_1128,N_1093);
and U1215 (N_1215,N_1165,N_1127);
nor U1216 (N_1216,N_1185,N_1190);
xnor U1217 (N_1217,N_1177,N_1188);
xor U1218 (N_1218,N_1181,N_1077);
nand U1219 (N_1219,N_1122,N_1074);
nand U1220 (N_1220,N_1152,N_1029);
or U1221 (N_1221,N_1164,N_1064);
nor U1222 (N_1222,N_1025,N_1068);
and U1223 (N_1223,N_1036,N_1111);
and U1224 (N_1224,N_1134,N_1009);
and U1225 (N_1225,N_1150,N_1070);
and U1226 (N_1226,N_1061,N_1082);
and U1227 (N_1227,N_1028,N_1129);
or U1228 (N_1228,N_1196,N_1079);
and U1229 (N_1229,N_1044,N_1045);
or U1230 (N_1230,N_1075,N_1078);
or U1231 (N_1231,N_1083,N_1021);
or U1232 (N_1232,N_1080,N_1087);
xor U1233 (N_1233,N_1014,N_1076);
nor U1234 (N_1234,N_1089,N_1059);
nor U1235 (N_1235,N_1194,N_1090);
and U1236 (N_1236,N_1086,N_1016);
or U1237 (N_1237,N_1138,N_1026);
or U1238 (N_1238,N_1038,N_1032);
nor U1239 (N_1239,N_1096,N_1040);
nand U1240 (N_1240,N_1178,N_1092);
and U1241 (N_1241,N_1120,N_1058);
nor U1242 (N_1242,N_1097,N_1133);
nor U1243 (N_1243,N_1149,N_1141);
nor U1244 (N_1244,N_1153,N_1124);
and U1245 (N_1245,N_1163,N_1066);
or U1246 (N_1246,N_1140,N_1174);
nor U1247 (N_1247,N_1173,N_1195);
nand U1248 (N_1248,N_1100,N_1067);
and U1249 (N_1249,N_1002,N_1039);
nor U1250 (N_1250,N_1105,N_1130);
nor U1251 (N_1251,N_1156,N_1154);
and U1252 (N_1252,N_1011,N_1006);
nor U1253 (N_1253,N_1109,N_1046);
nand U1254 (N_1254,N_1146,N_1160);
or U1255 (N_1255,N_1091,N_1108);
or U1256 (N_1256,N_1147,N_1062);
and U1257 (N_1257,N_1031,N_1175);
nand U1258 (N_1258,N_1012,N_1157);
or U1259 (N_1259,N_1117,N_1037);
nand U1260 (N_1260,N_1007,N_1048);
nand U1261 (N_1261,N_1198,N_1000);
and U1262 (N_1262,N_1018,N_1072);
and U1263 (N_1263,N_1167,N_1142);
and U1264 (N_1264,N_1182,N_1170);
or U1265 (N_1265,N_1095,N_1073);
nor U1266 (N_1266,N_1176,N_1015);
nor U1267 (N_1267,N_1053,N_1107);
and U1268 (N_1268,N_1023,N_1057);
and U1269 (N_1269,N_1101,N_1123);
xor U1270 (N_1270,N_1171,N_1199);
or U1271 (N_1271,N_1183,N_1158);
nor U1272 (N_1272,N_1118,N_1113);
or U1273 (N_1273,N_1010,N_1114);
and U1274 (N_1274,N_1003,N_1179);
and U1275 (N_1275,N_1047,N_1056);
or U1276 (N_1276,N_1197,N_1126);
nand U1277 (N_1277,N_1033,N_1049);
nor U1278 (N_1278,N_1004,N_1162);
nand U1279 (N_1279,N_1024,N_1103);
nand U1280 (N_1280,N_1054,N_1052);
and U1281 (N_1281,N_1168,N_1119);
nor U1282 (N_1282,N_1148,N_1069);
and U1283 (N_1283,N_1184,N_1144);
and U1284 (N_1284,N_1094,N_1017);
nand U1285 (N_1285,N_1180,N_1131);
or U1286 (N_1286,N_1145,N_1132);
nand U1287 (N_1287,N_1166,N_1034);
nand U1288 (N_1288,N_1104,N_1135);
and U1289 (N_1289,N_1035,N_1155);
or U1290 (N_1290,N_1137,N_1136);
or U1291 (N_1291,N_1106,N_1041);
nor U1292 (N_1292,N_1065,N_1189);
and U1293 (N_1293,N_1042,N_1192);
nor U1294 (N_1294,N_1043,N_1013);
or U1295 (N_1295,N_1143,N_1050);
nand U1296 (N_1296,N_1063,N_1071);
nand U1297 (N_1297,N_1125,N_1116);
nand U1298 (N_1298,N_1027,N_1102);
or U1299 (N_1299,N_1060,N_1193);
and U1300 (N_1300,N_1038,N_1035);
or U1301 (N_1301,N_1172,N_1057);
nand U1302 (N_1302,N_1148,N_1111);
and U1303 (N_1303,N_1151,N_1086);
xor U1304 (N_1304,N_1099,N_1011);
or U1305 (N_1305,N_1063,N_1037);
and U1306 (N_1306,N_1179,N_1086);
xor U1307 (N_1307,N_1125,N_1096);
nand U1308 (N_1308,N_1140,N_1032);
nand U1309 (N_1309,N_1157,N_1196);
nand U1310 (N_1310,N_1090,N_1131);
nand U1311 (N_1311,N_1029,N_1112);
or U1312 (N_1312,N_1108,N_1069);
xor U1313 (N_1313,N_1074,N_1010);
or U1314 (N_1314,N_1057,N_1080);
and U1315 (N_1315,N_1141,N_1196);
and U1316 (N_1316,N_1116,N_1108);
and U1317 (N_1317,N_1001,N_1015);
nand U1318 (N_1318,N_1008,N_1087);
or U1319 (N_1319,N_1089,N_1006);
or U1320 (N_1320,N_1087,N_1199);
nor U1321 (N_1321,N_1078,N_1021);
nor U1322 (N_1322,N_1090,N_1177);
or U1323 (N_1323,N_1105,N_1033);
and U1324 (N_1324,N_1129,N_1094);
nor U1325 (N_1325,N_1100,N_1182);
nand U1326 (N_1326,N_1068,N_1106);
or U1327 (N_1327,N_1149,N_1000);
or U1328 (N_1328,N_1082,N_1192);
or U1329 (N_1329,N_1057,N_1025);
nor U1330 (N_1330,N_1053,N_1157);
or U1331 (N_1331,N_1171,N_1053);
and U1332 (N_1332,N_1041,N_1043);
xnor U1333 (N_1333,N_1141,N_1107);
or U1334 (N_1334,N_1183,N_1008);
xnor U1335 (N_1335,N_1111,N_1009);
or U1336 (N_1336,N_1041,N_1120);
and U1337 (N_1337,N_1055,N_1019);
or U1338 (N_1338,N_1073,N_1074);
nor U1339 (N_1339,N_1093,N_1024);
xor U1340 (N_1340,N_1126,N_1027);
and U1341 (N_1341,N_1018,N_1189);
or U1342 (N_1342,N_1067,N_1132);
or U1343 (N_1343,N_1102,N_1021);
or U1344 (N_1344,N_1158,N_1124);
nand U1345 (N_1345,N_1081,N_1170);
nand U1346 (N_1346,N_1064,N_1028);
nand U1347 (N_1347,N_1158,N_1071);
nor U1348 (N_1348,N_1193,N_1061);
nand U1349 (N_1349,N_1151,N_1190);
and U1350 (N_1350,N_1139,N_1089);
nor U1351 (N_1351,N_1087,N_1108);
or U1352 (N_1352,N_1180,N_1076);
or U1353 (N_1353,N_1092,N_1124);
nor U1354 (N_1354,N_1182,N_1033);
nor U1355 (N_1355,N_1130,N_1152);
nor U1356 (N_1356,N_1078,N_1127);
or U1357 (N_1357,N_1025,N_1036);
nor U1358 (N_1358,N_1090,N_1082);
nor U1359 (N_1359,N_1132,N_1035);
or U1360 (N_1360,N_1167,N_1058);
or U1361 (N_1361,N_1015,N_1112);
or U1362 (N_1362,N_1158,N_1060);
nand U1363 (N_1363,N_1078,N_1146);
nand U1364 (N_1364,N_1156,N_1149);
and U1365 (N_1365,N_1173,N_1092);
xnor U1366 (N_1366,N_1173,N_1005);
nor U1367 (N_1367,N_1123,N_1007);
nor U1368 (N_1368,N_1189,N_1011);
and U1369 (N_1369,N_1169,N_1173);
or U1370 (N_1370,N_1031,N_1024);
nand U1371 (N_1371,N_1104,N_1194);
or U1372 (N_1372,N_1157,N_1006);
nor U1373 (N_1373,N_1012,N_1148);
nand U1374 (N_1374,N_1055,N_1199);
nand U1375 (N_1375,N_1195,N_1107);
nand U1376 (N_1376,N_1068,N_1031);
nor U1377 (N_1377,N_1093,N_1179);
xor U1378 (N_1378,N_1044,N_1122);
and U1379 (N_1379,N_1062,N_1042);
or U1380 (N_1380,N_1018,N_1009);
nor U1381 (N_1381,N_1139,N_1036);
xnor U1382 (N_1382,N_1058,N_1098);
nand U1383 (N_1383,N_1188,N_1158);
and U1384 (N_1384,N_1194,N_1057);
nor U1385 (N_1385,N_1063,N_1082);
and U1386 (N_1386,N_1142,N_1189);
nand U1387 (N_1387,N_1020,N_1014);
or U1388 (N_1388,N_1036,N_1028);
and U1389 (N_1389,N_1015,N_1100);
or U1390 (N_1390,N_1187,N_1194);
and U1391 (N_1391,N_1078,N_1080);
or U1392 (N_1392,N_1168,N_1192);
nor U1393 (N_1393,N_1199,N_1142);
nor U1394 (N_1394,N_1141,N_1033);
nor U1395 (N_1395,N_1187,N_1096);
and U1396 (N_1396,N_1016,N_1109);
nor U1397 (N_1397,N_1117,N_1040);
nand U1398 (N_1398,N_1119,N_1190);
nor U1399 (N_1399,N_1034,N_1014);
and U1400 (N_1400,N_1234,N_1318);
nand U1401 (N_1401,N_1364,N_1214);
nor U1402 (N_1402,N_1356,N_1309);
nor U1403 (N_1403,N_1218,N_1388);
and U1404 (N_1404,N_1263,N_1334);
nand U1405 (N_1405,N_1368,N_1355);
or U1406 (N_1406,N_1217,N_1300);
or U1407 (N_1407,N_1286,N_1369);
xnor U1408 (N_1408,N_1324,N_1264);
nand U1409 (N_1409,N_1289,N_1261);
nand U1410 (N_1410,N_1345,N_1235);
xor U1411 (N_1411,N_1223,N_1222);
xor U1412 (N_1412,N_1249,N_1239);
or U1413 (N_1413,N_1238,N_1276);
xnor U1414 (N_1414,N_1308,N_1287);
or U1415 (N_1415,N_1332,N_1314);
nand U1416 (N_1416,N_1266,N_1328);
nor U1417 (N_1417,N_1383,N_1321);
nand U1418 (N_1418,N_1273,N_1386);
and U1419 (N_1419,N_1357,N_1336);
nand U1420 (N_1420,N_1269,N_1335);
or U1421 (N_1421,N_1379,N_1394);
nor U1422 (N_1422,N_1327,N_1359);
nand U1423 (N_1423,N_1397,N_1208);
and U1424 (N_1424,N_1225,N_1325);
or U1425 (N_1425,N_1272,N_1320);
or U1426 (N_1426,N_1277,N_1306);
nor U1427 (N_1427,N_1201,N_1285);
nand U1428 (N_1428,N_1230,N_1343);
nand U1429 (N_1429,N_1274,N_1329);
nor U1430 (N_1430,N_1268,N_1212);
nor U1431 (N_1431,N_1293,N_1341);
xor U1432 (N_1432,N_1295,N_1310);
nor U1433 (N_1433,N_1250,N_1221);
nor U1434 (N_1434,N_1372,N_1279);
nor U1435 (N_1435,N_1311,N_1202);
and U1436 (N_1436,N_1305,N_1354);
or U1437 (N_1437,N_1302,N_1389);
xor U1438 (N_1438,N_1290,N_1387);
nand U1439 (N_1439,N_1256,N_1232);
nand U1440 (N_1440,N_1315,N_1304);
xnor U1441 (N_1441,N_1252,N_1203);
and U1442 (N_1442,N_1366,N_1330);
and U1443 (N_1443,N_1262,N_1317);
xor U1444 (N_1444,N_1391,N_1224);
nand U1445 (N_1445,N_1378,N_1226);
nor U1446 (N_1446,N_1245,N_1283);
and U1447 (N_1447,N_1278,N_1381);
nand U1448 (N_1448,N_1301,N_1384);
or U1449 (N_1449,N_1361,N_1339);
nand U1450 (N_1450,N_1367,N_1253);
nand U1451 (N_1451,N_1288,N_1242);
nor U1452 (N_1452,N_1303,N_1382);
and U1453 (N_1453,N_1292,N_1231);
nor U1454 (N_1454,N_1370,N_1284);
nand U1455 (N_1455,N_1348,N_1377);
and U1456 (N_1456,N_1349,N_1312);
or U1457 (N_1457,N_1322,N_1319);
nand U1458 (N_1458,N_1346,N_1390);
and U1459 (N_1459,N_1326,N_1342);
and U1460 (N_1460,N_1257,N_1371);
and U1461 (N_1461,N_1229,N_1265);
nor U1462 (N_1462,N_1271,N_1204);
nand U1463 (N_1463,N_1243,N_1258);
nor U1464 (N_1464,N_1236,N_1375);
or U1465 (N_1465,N_1362,N_1240);
xor U1466 (N_1466,N_1393,N_1313);
nand U1467 (N_1467,N_1244,N_1352);
xnor U1468 (N_1468,N_1281,N_1259);
or U1469 (N_1469,N_1206,N_1316);
xor U1470 (N_1470,N_1219,N_1215);
nor U1471 (N_1471,N_1351,N_1228);
nand U1472 (N_1472,N_1248,N_1254);
and U1473 (N_1473,N_1251,N_1376);
nor U1474 (N_1474,N_1363,N_1331);
nand U1475 (N_1475,N_1385,N_1233);
nand U1476 (N_1476,N_1396,N_1373);
and U1477 (N_1477,N_1358,N_1275);
nand U1478 (N_1478,N_1220,N_1260);
or U1479 (N_1479,N_1237,N_1307);
nor U1480 (N_1480,N_1323,N_1347);
xor U1481 (N_1481,N_1210,N_1211);
nor U1482 (N_1482,N_1360,N_1380);
nor U1483 (N_1483,N_1216,N_1207);
and U1484 (N_1484,N_1344,N_1298);
and U1485 (N_1485,N_1209,N_1255);
or U1486 (N_1486,N_1267,N_1392);
nand U1487 (N_1487,N_1399,N_1294);
nor U1488 (N_1488,N_1333,N_1270);
or U1489 (N_1489,N_1213,N_1340);
and U1490 (N_1490,N_1365,N_1291);
and U1491 (N_1491,N_1282,N_1205);
and U1492 (N_1492,N_1200,N_1227);
nand U1493 (N_1493,N_1350,N_1280);
nor U1494 (N_1494,N_1241,N_1338);
and U1495 (N_1495,N_1247,N_1374);
xnor U1496 (N_1496,N_1296,N_1337);
nor U1497 (N_1497,N_1297,N_1395);
and U1498 (N_1498,N_1353,N_1398);
and U1499 (N_1499,N_1246,N_1299);
nand U1500 (N_1500,N_1394,N_1332);
nor U1501 (N_1501,N_1250,N_1331);
nand U1502 (N_1502,N_1264,N_1249);
nor U1503 (N_1503,N_1335,N_1278);
nand U1504 (N_1504,N_1337,N_1292);
nand U1505 (N_1505,N_1308,N_1280);
and U1506 (N_1506,N_1311,N_1249);
and U1507 (N_1507,N_1369,N_1365);
nor U1508 (N_1508,N_1365,N_1383);
nor U1509 (N_1509,N_1249,N_1363);
and U1510 (N_1510,N_1229,N_1302);
or U1511 (N_1511,N_1399,N_1329);
or U1512 (N_1512,N_1224,N_1357);
nand U1513 (N_1513,N_1255,N_1216);
or U1514 (N_1514,N_1303,N_1397);
or U1515 (N_1515,N_1353,N_1347);
and U1516 (N_1516,N_1304,N_1373);
nand U1517 (N_1517,N_1205,N_1386);
and U1518 (N_1518,N_1264,N_1273);
nor U1519 (N_1519,N_1337,N_1210);
and U1520 (N_1520,N_1331,N_1371);
nor U1521 (N_1521,N_1254,N_1391);
nand U1522 (N_1522,N_1352,N_1234);
or U1523 (N_1523,N_1309,N_1313);
or U1524 (N_1524,N_1290,N_1281);
and U1525 (N_1525,N_1373,N_1279);
or U1526 (N_1526,N_1258,N_1314);
nand U1527 (N_1527,N_1398,N_1239);
nor U1528 (N_1528,N_1260,N_1363);
and U1529 (N_1529,N_1301,N_1356);
and U1530 (N_1530,N_1265,N_1268);
xor U1531 (N_1531,N_1322,N_1379);
nand U1532 (N_1532,N_1386,N_1240);
or U1533 (N_1533,N_1293,N_1383);
or U1534 (N_1534,N_1277,N_1320);
and U1535 (N_1535,N_1283,N_1352);
or U1536 (N_1536,N_1377,N_1303);
or U1537 (N_1537,N_1241,N_1367);
nor U1538 (N_1538,N_1360,N_1252);
nor U1539 (N_1539,N_1238,N_1323);
or U1540 (N_1540,N_1369,N_1268);
nand U1541 (N_1541,N_1380,N_1323);
nor U1542 (N_1542,N_1250,N_1206);
and U1543 (N_1543,N_1398,N_1375);
nor U1544 (N_1544,N_1208,N_1219);
nand U1545 (N_1545,N_1247,N_1237);
xnor U1546 (N_1546,N_1348,N_1313);
nand U1547 (N_1547,N_1376,N_1246);
xor U1548 (N_1548,N_1387,N_1360);
nor U1549 (N_1549,N_1299,N_1217);
and U1550 (N_1550,N_1361,N_1352);
and U1551 (N_1551,N_1275,N_1259);
nor U1552 (N_1552,N_1203,N_1310);
or U1553 (N_1553,N_1385,N_1278);
or U1554 (N_1554,N_1295,N_1309);
xnor U1555 (N_1555,N_1227,N_1267);
and U1556 (N_1556,N_1321,N_1297);
nand U1557 (N_1557,N_1208,N_1237);
nand U1558 (N_1558,N_1379,N_1296);
xor U1559 (N_1559,N_1306,N_1336);
nor U1560 (N_1560,N_1386,N_1375);
nand U1561 (N_1561,N_1323,N_1217);
nand U1562 (N_1562,N_1364,N_1341);
or U1563 (N_1563,N_1368,N_1223);
nand U1564 (N_1564,N_1211,N_1203);
and U1565 (N_1565,N_1316,N_1293);
nor U1566 (N_1566,N_1300,N_1381);
nand U1567 (N_1567,N_1394,N_1229);
and U1568 (N_1568,N_1327,N_1262);
and U1569 (N_1569,N_1308,N_1298);
nand U1570 (N_1570,N_1399,N_1308);
or U1571 (N_1571,N_1271,N_1364);
xor U1572 (N_1572,N_1370,N_1237);
nand U1573 (N_1573,N_1250,N_1308);
or U1574 (N_1574,N_1248,N_1341);
nand U1575 (N_1575,N_1316,N_1241);
and U1576 (N_1576,N_1365,N_1212);
nor U1577 (N_1577,N_1283,N_1370);
nor U1578 (N_1578,N_1374,N_1264);
and U1579 (N_1579,N_1295,N_1329);
xnor U1580 (N_1580,N_1330,N_1351);
nand U1581 (N_1581,N_1379,N_1335);
nand U1582 (N_1582,N_1355,N_1333);
or U1583 (N_1583,N_1217,N_1342);
nand U1584 (N_1584,N_1203,N_1279);
and U1585 (N_1585,N_1278,N_1344);
or U1586 (N_1586,N_1238,N_1298);
or U1587 (N_1587,N_1269,N_1361);
and U1588 (N_1588,N_1363,N_1351);
xnor U1589 (N_1589,N_1306,N_1221);
nand U1590 (N_1590,N_1235,N_1211);
or U1591 (N_1591,N_1376,N_1357);
xor U1592 (N_1592,N_1311,N_1316);
or U1593 (N_1593,N_1205,N_1293);
and U1594 (N_1594,N_1354,N_1348);
or U1595 (N_1595,N_1389,N_1364);
or U1596 (N_1596,N_1276,N_1392);
xor U1597 (N_1597,N_1367,N_1360);
nor U1598 (N_1598,N_1391,N_1220);
nand U1599 (N_1599,N_1254,N_1269);
nor U1600 (N_1600,N_1428,N_1500);
or U1601 (N_1601,N_1462,N_1510);
nand U1602 (N_1602,N_1528,N_1536);
or U1603 (N_1603,N_1522,N_1457);
nand U1604 (N_1604,N_1424,N_1423);
nand U1605 (N_1605,N_1456,N_1474);
or U1606 (N_1606,N_1592,N_1453);
or U1607 (N_1607,N_1465,N_1575);
nor U1608 (N_1608,N_1443,N_1440);
or U1609 (N_1609,N_1559,N_1485);
or U1610 (N_1610,N_1526,N_1556);
or U1611 (N_1611,N_1468,N_1501);
and U1612 (N_1612,N_1405,N_1496);
nor U1613 (N_1613,N_1553,N_1422);
nor U1614 (N_1614,N_1434,N_1557);
or U1615 (N_1615,N_1596,N_1475);
or U1616 (N_1616,N_1432,N_1525);
nand U1617 (N_1617,N_1472,N_1545);
nor U1618 (N_1618,N_1551,N_1566);
or U1619 (N_1619,N_1498,N_1558);
nand U1620 (N_1620,N_1590,N_1438);
and U1621 (N_1621,N_1582,N_1463);
and U1622 (N_1622,N_1452,N_1574);
nand U1623 (N_1623,N_1448,N_1524);
or U1624 (N_1624,N_1563,N_1447);
and U1625 (N_1625,N_1597,N_1517);
and U1626 (N_1626,N_1598,N_1503);
and U1627 (N_1627,N_1469,N_1460);
or U1628 (N_1628,N_1504,N_1535);
and U1629 (N_1629,N_1408,N_1539);
and U1630 (N_1630,N_1415,N_1430);
and U1631 (N_1631,N_1568,N_1550);
or U1632 (N_1632,N_1519,N_1418);
and U1633 (N_1633,N_1426,N_1402);
nor U1634 (N_1634,N_1527,N_1455);
nor U1635 (N_1635,N_1555,N_1546);
or U1636 (N_1636,N_1491,N_1466);
nor U1637 (N_1637,N_1492,N_1571);
nor U1638 (N_1638,N_1565,N_1483);
nand U1639 (N_1639,N_1581,N_1441);
and U1640 (N_1640,N_1508,N_1533);
nor U1641 (N_1641,N_1547,N_1413);
xor U1642 (N_1642,N_1437,N_1406);
nand U1643 (N_1643,N_1529,N_1537);
and U1644 (N_1644,N_1593,N_1461);
and U1645 (N_1645,N_1407,N_1587);
nor U1646 (N_1646,N_1481,N_1477);
nand U1647 (N_1647,N_1464,N_1499);
or U1648 (N_1648,N_1420,N_1490);
and U1649 (N_1649,N_1467,N_1417);
and U1650 (N_1650,N_1512,N_1534);
nand U1651 (N_1651,N_1564,N_1591);
or U1652 (N_1652,N_1589,N_1482);
nor U1653 (N_1653,N_1538,N_1531);
and U1654 (N_1654,N_1506,N_1540);
nand U1655 (N_1655,N_1480,N_1541);
or U1656 (N_1656,N_1567,N_1409);
nor U1657 (N_1657,N_1521,N_1403);
or U1658 (N_1658,N_1542,N_1509);
and U1659 (N_1659,N_1523,N_1450);
nor U1660 (N_1660,N_1442,N_1552);
or U1661 (N_1661,N_1431,N_1594);
and U1662 (N_1662,N_1404,N_1549);
or U1663 (N_1663,N_1507,N_1572);
xor U1664 (N_1664,N_1458,N_1532);
nand U1665 (N_1665,N_1562,N_1488);
nor U1666 (N_1666,N_1494,N_1416);
or U1667 (N_1667,N_1561,N_1451);
or U1668 (N_1668,N_1580,N_1454);
or U1669 (N_1669,N_1576,N_1502);
or U1670 (N_1670,N_1459,N_1435);
and U1671 (N_1671,N_1530,N_1414);
nor U1672 (N_1672,N_1439,N_1436);
nand U1673 (N_1673,N_1470,N_1515);
and U1674 (N_1674,N_1513,N_1419);
and U1675 (N_1675,N_1511,N_1505);
or U1676 (N_1676,N_1595,N_1493);
nor U1677 (N_1677,N_1544,N_1577);
and U1678 (N_1678,N_1449,N_1444);
or U1679 (N_1679,N_1445,N_1518);
nand U1680 (N_1680,N_1586,N_1497);
nand U1681 (N_1681,N_1573,N_1429);
nand U1682 (N_1682,N_1516,N_1548);
xor U1683 (N_1683,N_1484,N_1478);
xor U1684 (N_1684,N_1412,N_1411);
nand U1685 (N_1685,N_1476,N_1570);
or U1686 (N_1686,N_1520,N_1579);
nor U1687 (N_1687,N_1421,N_1479);
or U1688 (N_1688,N_1446,N_1486);
and U1689 (N_1689,N_1471,N_1588);
nor U1690 (N_1690,N_1514,N_1569);
or U1691 (N_1691,N_1400,N_1584);
or U1692 (N_1692,N_1487,N_1427);
nor U1693 (N_1693,N_1578,N_1560);
nand U1694 (N_1694,N_1473,N_1401);
and U1695 (N_1695,N_1585,N_1495);
nor U1696 (N_1696,N_1489,N_1425);
or U1697 (N_1697,N_1433,N_1554);
nand U1698 (N_1698,N_1599,N_1583);
nor U1699 (N_1699,N_1410,N_1543);
nor U1700 (N_1700,N_1470,N_1412);
and U1701 (N_1701,N_1532,N_1583);
and U1702 (N_1702,N_1462,N_1488);
or U1703 (N_1703,N_1558,N_1536);
nand U1704 (N_1704,N_1577,N_1507);
and U1705 (N_1705,N_1587,N_1418);
nand U1706 (N_1706,N_1429,N_1478);
and U1707 (N_1707,N_1478,N_1475);
nor U1708 (N_1708,N_1413,N_1488);
or U1709 (N_1709,N_1521,N_1407);
and U1710 (N_1710,N_1493,N_1471);
or U1711 (N_1711,N_1410,N_1532);
and U1712 (N_1712,N_1545,N_1499);
nor U1713 (N_1713,N_1429,N_1462);
nor U1714 (N_1714,N_1442,N_1532);
xnor U1715 (N_1715,N_1572,N_1462);
or U1716 (N_1716,N_1485,N_1404);
nor U1717 (N_1717,N_1469,N_1596);
nand U1718 (N_1718,N_1481,N_1474);
nor U1719 (N_1719,N_1452,N_1587);
and U1720 (N_1720,N_1531,N_1447);
nor U1721 (N_1721,N_1476,N_1538);
and U1722 (N_1722,N_1470,N_1463);
or U1723 (N_1723,N_1533,N_1400);
nor U1724 (N_1724,N_1431,N_1500);
or U1725 (N_1725,N_1531,N_1440);
nor U1726 (N_1726,N_1508,N_1541);
and U1727 (N_1727,N_1519,N_1469);
or U1728 (N_1728,N_1433,N_1463);
and U1729 (N_1729,N_1584,N_1542);
or U1730 (N_1730,N_1573,N_1402);
xor U1731 (N_1731,N_1585,N_1466);
xnor U1732 (N_1732,N_1506,N_1580);
and U1733 (N_1733,N_1480,N_1419);
nor U1734 (N_1734,N_1504,N_1430);
and U1735 (N_1735,N_1482,N_1445);
and U1736 (N_1736,N_1442,N_1468);
nor U1737 (N_1737,N_1479,N_1584);
nand U1738 (N_1738,N_1584,N_1453);
nor U1739 (N_1739,N_1545,N_1430);
nor U1740 (N_1740,N_1596,N_1420);
nor U1741 (N_1741,N_1595,N_1406);
nor U1742 (N_1742,N_1494,N_1444);
nand U1743 (N_1743,N_1492,N_1543);
and U1744 (N_1744,N_1489,N_1517);
nor U1745 (N_1745,N_1538,N_1521);
or U1746 (N_1746,N_1558,N_1507);
or U1747 (N_1747,N_1472,N_1492);
or U1748 (N_1748,N_1417,N_1469);
or U1749 (N_1749,N_1450,N_1499);
and U1750 (N_1750,N_1531,N_1410);
nor U1751 (N_1751,N_1417,N_1439);
or U1752 (N_1752,N_1484,N_1548);
nor U1753 (N_1753,N_1557,N_1595);
and U1754 (N_1754,N_1570,N_1463);
nor U1755 (N_1755,N_1408,N_1440);
and U1756 (N_1756,N_1459,N_1584);
nor U1757 (N_1757,N_1529,N_1560);
nand U1758 (N_1758,N_1597,N_1532);
nand U1759 (N_1759,N_1413,N_1556);
and U1760 (N_1760,N_1518,N_1585);
nand U1761 (N_1761,N_1436,N_1494);
nor U1762 (N_1762,N_1499,N_1521);
nor U1763 (N_1763,N_1492,N_1446);
nand U1764 (N_1764,N_1504,N_1402);
nand U1765 (N_1765,N_1562,N_1426);
xor U1766 (N_1766,N_1561,N_1433);
or U1767 (N_1767,N_1595,N_1413);
or U1768 (N_1768,N_1502,N_1425);
or U1769 (N_1769,N_1582,N_1581);
and U1770 (N_1770,N_1471,N_1426);
xor U1771 (N_1771,N_1513,N_1532);
and U1772 (N_1772,N_1527,N_1541);
nand U1773 (N_1773,N_1425,N_1524);
xnor U1774 (N_1774,N_1496,N_1559);
or U1775 (N_1775,N_1437,N_1524);
and U1776 (N_1776,N_1548,N_1545);
nand U1777 (N_1777,N_1566,N_1453);
or U1778 (N_1778,N_1424,N_1594);
and U1779 (N_1779,N_1445,N_1426);
nor U1780 (N_1780,N_1585,N_1514);
or U1781 (N_1781,N_1533,N_1503);
nand U1782 (N_1782,N_1427,N_1594);
and U1783 (N_1783,N_1550,N_1408);
nand U1784 (N_1784,N_1548,N_1568);
and U1785 (N_1785,N_1599,N_1419);
xnor U1786 (N_1786,N_1453,N_1527);
xnor U1787 (N_1787,N_1475,N_1484);
or U1788 (N_1788,N_1541,N_1427);
nor U1789 (N_1789,N_1413,N_1572);
nor U1790 (N_1790,N_1596,N_1539);
nor U1791 (N_1791,N_1459,N_1449);
nand U1792 (N_1792,N_1557,N_1535);
xnor U1793 (N_1793,N_1585,N_1435);
nor U1794 (N_1794,N_1515,N_1519);
and U1795 (N_1795,N_1439,N_1558);
xnor U1796 (N_1796,N_1457,N_1506);
and U1797 (N_1797,N_1527,N_1469);
xor U1798 (N_1798,N_1448,N_1468);
nand U1799 (N_1799,N_1509,N_1413);
or U1800 (N_1800,N_1708,N_1742);
xnor U1801 (N_1801,N_1770,N_1658);
or U1802 (N_1802,N_1747,N_1710);
nor U1803 (N_1803,N_1703,N_1721);
nor U1804 (N_1804,N_1741,N_1711);
and U1805 (N_1805,N_1751,N_1725);
or U1806 (N_1806,N_1672,N_1784);
nand U1807 (N_1807,N_1772,N_1613);
and U1808 (N_1808,N_1763,N_1686);
or U1809 (N_1809,N_1637,N_1798);
nand U1810 (N_1810,N_1673,N_1759);
or U1811 (N_1811,N_1638,N_1702);
or U1812 (N_1812,N_1715,N_1746);
nand U1813 (N_1813,N_1714,N_1642);
nand U1814 (N_1814,N_1651,N_1609);
or U1815 (N_1815,N_1768,N_1753);
nor U1816 (N_1816,N_1756,N_1779);
or U1817 (N_1817,N_1719,N_1707);
xor U1818 (N_1818,N_1773,N_1631);
and U1819 (N_1819,N_1762,N_1688);
or U1820 (N_1820,N_1643,N_1644);
or U1821 (N_1821,N_1740,N_1749);
nand U1822 (N_1822,N_1668,N_1620);
or U1823 (N_1823,N_1696,N_1692);
nand U1824 (N_1824,N_1752,N_1743);
nand U1825 (N_1825,N_1664,N_1694);
nand U1826 (N_1826,N_1775,N_1611);
nand U1827 (N_1827,N_1723,N_1698);
or U1828 (N_1828,N_1717,N_1640);
xnor U1829 (N_1829,N_1755,N_1706);
nand U1830 (N_1830,N_1704,N_1757);
or U1831 (N_1831,N_1774,N_1685);
and U1832 (N_1832,N_1782,N_1799);
xor U1833 (N_1833,N_1649,N_1602);
nor U1834 (N_1834,N_1610,N_1671);
or U1835 (N_1835,N_1623,N_1736);
nand U1836 (N_1836,N_1699,N_1728);
and U1837 (N_1837,N_1712,N_1661);
nand U1838 (N_1838,N_1683,N_1679);
nand U1839 (N_1839,N_1786,N_1669);
nor U1840 (N_1840,N_1787,N_1633);
and U1841 (N_1841,N_1795,N_1760);
or U1842 (N_1842,N_1769,N_1713);
and U1843 (N_1843,N_1793,N_1629);
or U1844 (N_1844,N_1734,N_1607);
nand U1845 (N_1845,N_1767,N_1652);
xnor U1846 (N_1846,N_1785,N_1670);
nor U1847 (N_1847,N_1635,N_1701);
nor U1848 (N_1848,N_1691,N_1745);
nor U1849 (N_1849,N_1656,N_1733);
nand U1850 (N_1850,N_1695,N_1781);
or U1851 (N_1851,N_1606,N_1627);
or U1852 (N_1852,N_1617,N_1632);
or U1853 (N_1853,N_1709,N_1700);
nor U1854 (N_1854,N_1771,N_1738);
and U1855 (N_1855,N_1729,N_1615);
nor U1856 (N_1856,N_1720,N_1639);
and U1857 (N_1857,N_1618,N_1648);
nand U1858 (N_1858,N_1687,N_1744);
or U1859 (N_1859,N_1605,N_1797);
nor U1860 (N_1860,N_1657,N_1777);
xor U1861 (N_1861,N_1748,N_1612);
nand U1862 (N_1862,N_1601,N_1682);
nand U1863 (N_1863,N_1677,N_1645);
xnor U1864 (N_1864,N_1783,N_1614);
nand U1865 (N_1865,N_1680,N_1667);
nor U1866 (N_1866,N_1666,N_1655);
nand U1867 (N_1867,N_1675,N_1663);
or U1868 (N_1868,N_1624,N_1761);
nor U1869 (N_1869,N_1735,N_1754);
and U1870 (N_1870,N_1684,N_1791);
nand U1871 (N_1871,N_1674,N_1764);
or U1872 (N_1872,N_1660,N_1716);
or U1873 (N_1873,N_1780,N_1727);
and U1874 (N_1874,N_1730,N_1665);
xnor U1875 (N_1875,N_1788,N_1776);
nor U1876 (N_1876,N_1689,N_1619);
xnor U1877 (N_1877,N_1636,N_1603);
nand U1878 (N_1878,N_1600,N_1678);
and U1879 (N_1879,N_1778,N_1718);
or U1880 (N_1880,N_1739,N_1724);
or U1881 (N_1881,N_1737,N_1681);
nor U1882 (N_1882,N_1622,N_1621);
and U1883 (N_1883,N_1731,N_1650);
nor U1884 (N_1884,N_1790,N_1676);
nand U1885 (N_1885,N_1690,N_1626);
xor U1886 (N_1886,N_1634,N_1604);
and U1887 (N_1887,N_1726,N_1766);
nor U1888 (N_1888,N_1796,N_1765);
nand U1889 (N_1889,N_1625,N_1616);
xnor U1890 (N_1890,N_1722,N_1641);
or U1891 (N_1891,N_1693,N_1705);
and U1892 (N_1892,N_1662,N_1750);
or U1893 (N_1893,N_1654,N_1732);
and U1894 (N_1894,N_1653,N_1792);
nor U1895 (N_1895,N_1628,N_1630);
xor U1896 (N_1896,N_1646,N_1659);
and U1897 (N_1897,N_1789,N_1697);
nand U1898 (N_1898,N_1758,N_1608);
xnor U1899 (N_1899,N_1794,N_1647);
and U1900 (N_1900,N_1717,N_1646);
nand U1901 (N_1901,N_1660,N_1729);
or U1902 (N_1902,N_1615,N_1767);
or U1903 (N_1903,N_1644,N_1691);
or U1904 (N_1904,N_1764,N_1680);
nor U1905 (N_1905,N_1735,N_1648);
nand U1906 (N_1906,N_1789,N_1713);
or U1907 (N_1907,N_1758,N_1689);
nor U1908 (N_1908,N_1725,N_1642);
and U1909 (N_1909,N_1624,N_1724);
nand U1910 (N_1910,N_1790,N_1620);
xor U1911 (N_1911,N_1624,N_1614);
nand U1912 (N_1912,N_1707,N_1795);
xnor U1913 (N_1913,N_1714,N_1611);
and U1914 (N_1914,N_1632,N_1756);
or U1915 (N_1915,N_1769,N_1680);
or U1916 (N_1916,N_1752,N_1662);
and U1917 (N_1917,N_1703,N_1669);
nand U1918 (N_1918,N_1722,N_1625);
or U1919 (N_1919,N_1630,N_1688);
and U1920 (N_1920,N_1666,N_1771);
or U1921 (N_1921,N_1725,N_1789);
or U1922 (N_1922,N_1793,N_1687);
nor U1923 (N_1923,N_1730,N_1710);
xor U1924 (N_1924,N_1714,N_1790);
and U1925 (N_1925,N_1618,N_1719);
nor U1926 (N_1926,N_1639,N_1605);
or U1927 (N_1927,N_1645,N_1753);
and U1928 (N_1928,N_1776,N_1619);
nor U1929 (N_1929,N_1646,N_1705);
nor U1930 (N_1930,N_1738,N_1640);
and U1931 (N_1931,N_1745,N_1782);
or U1932 (N_1932,N_1746,N_1731);
nor U1933 (N_1933,N_1719,N_1772);
nand U1934 (N_1934,N_1601,N_1795);
nor U1935 (N_1935,N_1764,N_1622);
and U1936 (N_1936,N_1755,N_1698);
or U1937 (N_1937,N_1733,N_1675);
and U1938 (N_1938,N_1694,N_1783);
nand U1939 (N_1939,N_1720,N_1715);
nor U1940 (N_1940,N_1790,N_1602);
nor U1941 (N_1941,N_1612,N_1778);
or U1942 (N_1942,N_1627,N_1799);
and U1943 (N_1943,N_1709,N_1607);
and U1944 (N_1944,N_1755,N_1759);
nand U1945 (N_1945,N_1649,N_1657);
nor U1946 (N_1946,N_1740,N_1739);
xnor U1947 (N_1947,N_1683,N_1636);
nand U1948 (N_1948,N_1682,N_1691);
or U1949 (N_1949,N_1791,N_1751);
nor U1950 (N_1950,N_1728,N_1683);
or U1951 (N_1951,N_1654,N_1697);
nand U1952 (N_1952,N_1755,N_1617);
and U1953 (N_1953,N_1797,N_1667);
nand U1954 (N_1954,N_1675,N_1637);
and U1955 (N_1955,N_1742,N_1790);
and U1956 (N_1956,N_1668,N_1728);
nor U1957 (N_1957,N_1792,N_1729);
nor U1958 (N_1958,N_1605,N_1779);
and U1959 (N_1959,N_1649,N_1655);
nand U1960 (N_1960,N_1711,N_1681);
nand U1961 (N_1961,N_1709,N_1600);
xnor U1962 (N_1962,N_1775,N_1733);
nor U1963 (N_1963,N_1738,N_1767);
xnor U1964 (N_1964,N_1787,N_1685);
nor U1965 (N_1965,N_1615,N_1738);
nor U1966 (N_1966,N_1611,N_1788);
xor U1967 (N_1967,N_1780,N_1666);
or U1968 (N_1968,N_1706,N_1764);
xnor U1969 (N_1969,N_1680,N_1722);
or U1970 (N_1970,N_1655,N_1674);
nand U1971 (N_1971,N_1792,N_1716);
and U1972 (N_1972,N_1673,N_1642);
or U1973 (N_1973,N_1790,N_1651);
and U1974 (N_1974,N_1640,N_1698);
nor U1975 (N_1975,N_1610,N_1766);
xnor U1976 (N_1976,N_1733,N_1799);
and U1977 (N_1977,N_1696,N_1665);
or U1978 (N_1978,N_1780,N_1622);
and U1979 (N_1979,N_1652,N_1655);
or U1980 (N_1980,N_1700,N_1725);
nor U1981 (N_1981,N_1745,N_1642);
nor U1982 (N_1982,N_1651,N_1689);
and U1983 (N_1983,N_1660,N_1768);
or U1984 (N_1984,N_1714,N_1720);
and U1985 (N_1985,N_1672,N_1660);
or U1986 (N_1986,N_1739,N_1737);
or U1987 (N_1987,N_1638,N_1684);
nand U1988 (N_1988,N_1630,N_1758);
or U1989 (N_1989,N_1766,N_1723);
nor U1990 (N_1990,N_1797,N_1729);
nand U1991 (N_1991,N_1779,N_1659);
xnor U1992 (N_1992,N_1601,N_1778);
nor U1993 (N_1993,N_1796,N_1759);
nor U1994 (N_1994,N_1773,N_1678);
nand U1995 (N_1995,N_1790,N_1746);
and U1996 (N_1996,N_1758,N_1767);
or U1997 (N_1997,N_1618,N_1621);
nand U1998 (N_1998,N_1679,N_1609);
nor U1999 (N_1999,N_1734,N_1627);
or U2000 (N_2000,N_1903,N_1940);
xnor U2001 (N_2001,N_1906,N_1883);
nand U2002 (N_2002,N_1913,N_1810);
nor U2003 (N_2003,N_1801,N_1980);
and U2004 (N_2004,N_1986,N_1994);
nor U2005 (N_2005,N_1944,N_1802);
xnor U2006 (N_2006,N_1925,N_1975);
and U2007 (N_2007,N_1952,N_1857);
nor U2008 (N_2008,N_1886,N_1837);
nor U2009 (N_2009,N_1951,N_1965);
nand U2010 (N_2010,N_1891,N_1998);
nand U2011 (N_2011,N_1938,N_1909);
nand U2012 (N_2012,N_1989,N_1895);
nand U2013 (N_2013,N_1863,N_1880);
nand U2014 (N_2014,N_1996,N_1820);
or U2015 (N_2015,N_1889,N_1967);
and U2016 (N_2016,N_1814,N_1833);
nand U2017 (N_2017,N_1867,N_1845);
nor U2018 (N_2018,N_1842,N_1958);
nand U2019 (N_2019,N_1907,N_1868);
nand U2020 (N_2020,N_1969,N_1804);
nor U2021 (N_2021,N_1920,N_1834);
nand U2022 (N_2022,N_1847,N_1990);
nand U2023 (N_2023,N_1873,N_1841);
nor U2024 (N_2024,N_1946,N_1878);
nor U2025 (N_2025,N_1840,N_1849);
and U2026 (N_2026,N_1932,N_1968);
nor U2027 (N_2027,N_1861,N_1928);
nor U2028 (N_2028,N_1827,N_1914);
nand U2029 (N_2029,N_1901,N_1872);
or U2030 (N_2030,N_1978,N_1874);
and U2031 (N_2031,N_1950,N_1904);
or U2032 (N_2032,N_1830,N_1890);
and U2033 (N_2033,N_1809,N_1995);
nor U2034 (N_2034,N_1806,N_1936);
nor U2035 (N_2035,N_1821,N_1915);
or U2036 (N_2036,N_1937,N_1910);
nand U2037 (N_2037,N_1985,N_1858);
nor U2038 (N_2038,N_1959,N_1977);
nand U2039 (N_2039,N_1853,N_1972);
nand U2040 (N_2040,N_1999,N_1973);
or U2041 (N_2041,N_1875,N_1905);
and U2042 (N_2042,N_1939,N_1817);
xor U2043 (N_2043,N_1988,N_1921);
nand U2044 (N_2044,N_1930,N_1976);
or U2045 (N_2045,N_1902,N_1927);
and U2046 (N_2046,N_1819,N_1803);
nor U2047 (N_2047,N_1933,N_1960);
nor U2048 (N_2048,N_1865,N_1974);
or U2049 (N_2049,N_1851,N_1822);
or U2050 (N_2050,N_1979,N_1839);
and U2051 (N_2051,N_1924,N_1815);
or U2052 (N_2052,N_1898,N_1825);
xnor U2053 (N_2053,N_1911,N_1919);
and U2054 (N_2054,N_1981,N_1860);
nand U2055 (N_2055,N_1983,N_1900);
xor U2056 (N_2056,N_1897,N_1934);
nor U2057 (N_2057,N_1871,N_1956);
nor U2058 (N_2058,N_1943,N_1881);
nor U2059 (N_2059,N_1870,N_1843);
and U2060 (N_2060,N_1823,N_1836);
nor U2061 (N_2061,N_1953,N_1963);
nand U2062 (N_2062,N_1882,N_1917);
and U2063 (N_2063,N_1838,N_1879);
or U2064 (N_2064,N_1829,N_1844);
nor U2065 (N_2065,N_1805,N_1899);
nand U2066 (N_2066,N_1987,N_1923);
xnor U2067 (N_2067,N_1855,N_1947);
and U2068 (N_2068,N_1856,N_1888);
xnor U2069 (N_2069,N_1876,N_1929);
nand U2070 (N_2070,N_1997,N_1945);
or U2071 (N_2071,N_1970,N_1892);
xnor U2072 (N_2072,N_1811,N_1852);
or U2073 (N_2073,N_1912,N_1826);
nor U2074 (N_2074,N_1846,N_1926);
or U2075 (N_2075,N_1908,N_1931);
nor U2076 (N_2076,N_1885,N_1954);
or U2077 (N_2077,N_1866,N_1854);
and U2078 (N_2078,N_1877,N_1948);
or U2079 (N_2079,N_1800,N_1984);
and U2080 (N_2080,N_1894,N_1828);
and U2081 (N_2081,N_1961,N_1962);
and U2082 (N_2082,N_1832,N_1916);
nand U2083 (N_2083,N_1884,N_1992);
nor U2084 (N_2084,N_1864,N_1808);
and U2085 (N_2085,N_1941,N_1942);
nor U2086 (N_2086,N_1991,N_1955);
nand U2087 (N_2087,N_1824,N_1982);
or U2088 (N_2088,N_1848,N_1964);
nand U2089 (N_2089,N_1813,N_1831);
nor U2090 (N_2090,N_1993,N_1807);
nand U2091 (N_2091,N_1918,N_1816);
nand U2092 (N_2092,N_1893,N_1966);
nand U2093 (N_2093,N_1887,N_1922);
or U2094 (N_2094,N_1949,N_1835);
or U2095 (N_2095,N_1818,N_1862);
nand U2096 (N_2096,N_1896,N_1971);
nor U2097 (N_2097,N_1859,N_1869);
or U2098 (N_2098,N_1957,N_1812);
nor U2099 (N_2099,N_1935,N_1850);
nand U2100 (N_2100,N_1836,N_1807);
or U2101 (N_2101,N_1924,N_1994);
nand U2102 (N_2102,N_1852,N_1862);
nor U2103 (N_2103,N_1809,N_1847);
and U2104 (N_2104,N_1990,N_1899);
or U2105 (N_2105,N_1969,N_1847);
xnor U2106 (N_2106,N_1862,N_1957);
xnor U2107 (N_2107,N_1849,N_1932);
nor U2108 (N_2108,N_1806,N_1818);
nand U2109 (N_2109,N_1839,N_1892);
and U2110 (N_2110,N_1974,N_1904);
and U2111 (N_2111,N_1886,N_1820);
nor U2112 (N_2112,N_1944,N_1950);
and U2113 (N_2113,N_1990,N_1957);
nand U2114 (N_2114,N_1805,N_1940);
nand U2115 (N_2115,N_1967,N_1912);
or U2116 (N_2116,N_1815,N_1974);
nor U2117 (N_2117,N_1876,N_1948);
nand U2118 (N_2118,N_1908,N_1903);
or U2119 (N_2119,N_1847,N_1926);
xnor U2120 (N_2120,N_1901,N_1937);
nor U2121 (N_2121,N_1877,N_1965);
nand U2122 (N_2122,N_1829,N_1860);
nand U2123 (N_2123,N_1907,N_1944);
or U2124 (N_2124,N_1836,N_1834);
nor U2125 (N_2125,N_1903,N_1841);
and U2126 (N_2126,N_1875,N_1965);
and U2127 (N_2127,N_1877,N_1972);
and U2128 (N_2128,N_1962,N_1832);
and U2129 (N_2129,N_1967,N_1890);
xnor U2130 (N_2130,N_1822,N_1886);
or U2131 (N_2131,N_1910,N_1825);
and U2132 (N_2132,N_1806,N_1980);
and U2133 (N_2133,N_1881,N_1805);
nand U2134 (N_2134,N_1958,N_1900);
nand U2135 (N_2135,N_1825,N_1882);
xor U2136 (N_2136,N_1889,N_1860);
xnor U2137 (N_2137,N_1882,N_1900);
or U2138 (N_2138,N_1997,N_1803);
nand U2139 (N_2139,N_1988,N_1994);
nor U2140 (N_2140,N_1830,N_1876);
nand U2141 (N_2141,N_1912,N_1875);
xnor U2142 (N_2142,N_1937,N_1822);
or U2143 (N_2143,N_1909,N_1882);
or U2144 (N_2144,N_1830,N_1862);
nand U2145 (N_2145,N_1983,N_1935);
nor U2146 (N_2146,N_1823,N_1928);
nor U2147 (N_2147,N_1962,N_1822);
nor U2148 (N_2148,N_1919,N_1807);
nand U2149 (N_2149,N_1800,N_1822);
nand U2150 (N_2150,N_1917,N_1974);
or U2151 (N_2151,N_1886,N_1887);
or U2152 (N_2152,N_1829,N_1938);
or U2153 (N_2153,N_1817,N_1905);
and U2154 (N_2154,N_1977,N_1881);
xor U2155 (N_2155,N_1814,N_1988);
nor U2156 (N_2156,N_1884,N_1989);
and U2157 (N_2157,N_1984,N_1838);
and U2158 (N_2158,N_1906,N_1840);
nand U2159 (N_2159,N_1806,N_1834);
nor U2160 (N_2160,N_1998,N_1890);
and U2161 (N_2161,N_1819,N_1924);
nand U2162 (N_2162,N_1945,N_1831);
xnor U2163 (N_2163,N_1824,N_1898);
or U2164 (N_2164,N_1958,N_1820);
nor U2165 (N_2165,N_1971,N_1982);
nor U2166 (N_2166,N_1894,N_1903);
xnor U2167 (N_2167,N_1915,N_1854);
or U2168 (N_2168,N_1976,N_1937);
nor U2169 (N_2169,N_1945,N_1902);
and U2170 (N_2170,N_1875,N_1864);
or U2171 (N_2171,N_1842,N_1949);
nand U2172 (N_2172,N_1831,N_1904);
nand U2173 (N_2173,N_1843,N_1875);
nand U2174 (N_2174,N_1874,N_1816);
and U2175 (N_2175,N_1998,N_1985);
nand U2176 (N_2176,N_1911,N_1873);
and U2177 (N_2177,N_1844,N_1910);
or U2178 (N_2178,N_1938,N_1896);
and U2179 (N_2179,N_1899,N_1818);
nand U2180 (N_2180,N_1874,N_1940);
or U2181 (N_2181,N_1947,N_1995);
or U2182 (N_2182,N_1958,N_1830);
nor U2183 (N_2183,N_1933,N_1999);
and U2184 (N_2184,N_1930,N_1862);
nand U2185 (N_2185,N_1893,N_1849);
xnor U2186 (N_2186,N_1915,N_1976);
or U2187 (N_2187,N_1963,N_1973);
nand U2188 (N_2188,N_1840,N_1819);
and U2189 (N_2189,N_1810,N_1886);
or U2190 (N_2190,N_1943,N_1829);
nor U2191 (N_2191,N_1951,N_1876);
nand U2192 (N_2192,N_1971,N_1809);
nand U2193 (N_2193,N_1894,N_1898);
and U2194 (N_2194,N_1865,N_1858);
or U2195 (N_2195,N_1974,N_1960);
or U2196 (N_2196,N_1822,N_1895);
nor U2197 (N_2197,N_1860,N_1903);
or U2198 (N_2198,N_1948,N_1907);
nand U2199 (N_2199,N_1879,N_1867);
nor U2200 (N_2200,N_2104,N_2008);
and U2201 (N_2201,N_2080,N_2061);
nand U2202 (N_2202,N_2180,N_2033);
nor U2203 (N_2203,N_2006,N_2060);
or U2204 (N_2204,N_2148,N_2076);
or U2205 (N_2205,N_2025,N_2197);
nand U2206 (N_2206,N_2102,N_2103);
or U2207 (N_2207,N_2055,N_2020);
xnor U2208 (N_2208,N_2154,N_2046);
xor U2209 (N_2209,N_2163,N_2040);
nor U2210 (N_2210,N_2065,N_2053);
nand U2211 (N_2211,N_2098,N_2023);
nor U2212 (N_2212,N_2035,N_2017);
nand U2213 (N_2213,N_2031,N_2089);
nor U2214 (N_2214,N_2131,N_2042);
nor U2215 (N_2215,N_2097,N_2018);
or U2216 (N_2216,N_2110,N_2185);
nand U2217 (N_2217,N_2192,N_2118);
nand U2218 (N_2218,N_2028,N_2013);
nor U2219 (N_2219,N_2059,N_2187);
nand U2220 (N_2220,N_2157,N_2128);
and U2221 (N_2221,N_2156,N_2134);
or U2222 (N_2222,N_2123,N_2054);
nor U2223 (N_2223,N_2041,N_2147);
and U2224 (N_2224,N_2144,N_2078);
nand U2225 (N_2225,N_2198,N_2005);
and U2226 (N_2226,N_2051,N_2047);
and U2227 (N_2227,N_2093,N_2058);
xor U2228 (N_2228,N_2133,N_2090);
nor U2229 (N_2229,N_2159,N_2056);
nand U2230 (N_2230,N_2083,N_2009);
or U2231 (N_2231,N_2146,N_2100);
nor U2232 (N_2232,N_2038,N_2048);
and U2233 (N_2233,N_2044,N_2193);
and U2234 (N_2234,N_2138,N_2043);
or U2235 (N_2235,N_2030,N_2137);
and U2236 (N_2236,N_2049,N_2099);
nor U2237 (N_2237,N_2139,N_2149);
and U2238 (N_2238,N_2062,N_2127);
and U2239 (N_2239,N_2140,N_2145);
or U2240 (N_2240,N_2000,N_2153);
and U2241 (N_2241,N_2165,N_2002);
nand U2242 (N_2242,N_2113,N_2088);
nor U2243 (N_2243,N_2195,N_2050);
xor U2244 (N_2244,N_2072,N_2112);
nor U2245 (N_2245,N_2122,N_2191);
nor U2246 (N_2246,N_2116,N_2177);
and U2247 (N_2247,N_2001,N_2096);
nand U2248 (N_2248,N_2019,N_2079);
and U2249 (N_2249,N_2036,N_2007);
and U2250 (N_2250,N_2160,N_2011);
nor U2251 (N_2251,N_2179,N_2012);
nand U2252 (N_2252,N_2039,N_2081);
nand U2253 (N_2253,N_2064,N_2027);
nor U2254 (N_2254,N_2164,N_2057);
nand U2255 (N_2255,N_2052,N_2092);
nor U2256 (N_2256,N_2120,N_2190);
nor U2257 (N_2257,N_2015,N_2106);
and U2258 (N_2258,N_2114,N_2168);
and U2259 (N_2259,N_2129,N_2150);
nor U2260 (N_2260,N_2094,N_2143);
or U2261 (N_2261,N_2085,N_2166);
nor U2262 (N_2262,N_2124,N_2178);
nor U2263 (N_2263,N_2024,N_2175);
nor U2264 (N_2264,N_2125,N_2158);
and U2265 (N_2265,N_2174,N_2010);
nor U2266 (N_2266,N_2152,N_2022);
nand U2267 (N_2267,N_2181,N_2091);
nand U2268 (N_2268,N_2109,N_2014);
xor U2269 (N_2269,N_2073,N_2173);
nor U2270 (N_2270,N_2066,N_2029);
or U2271 (N_2271,N_2171,N_2069);
and U2272 (N_2272,N_2142,N_2075);
nor U2273 (N_2273,N_2037,N_2135);
nand U2274 (N_2274,N_2087,N_2107);
or U2275 (N_2275,N_2034,N_2183);
nand U2276 (N_2276,N_2108,N_2045);
nand U2277 (N_2277,N_2184,N_2132);
and U2278 (N_2278,N_2199,N_2136);
or U2279 (N_2279,N_2141,N_2082);
and U2280 (N_2280,N_2115,N_2117);
nor U2281 (N_2281,N_2074,N_2155);
nor U2282 (N_2282,N_2084,N_2182);
or U2283 (N_2283,N_2021,N_2194);
nand U2284 (N_2284,N_2176,N_2095);
xnor U2285 (N_2285,N_2077,N_2101);
nand U2286 (N_2286,N_2063,N_2188);
nor U2287 (N_2287,N_2121,N_2170);
or U2288 (N_2288,N_2070,N_2126);
or U2289 (N_2289,N_2086,N_2026);
or U2290 (N_2290,N_2105,N_2151);
nand U2291 (N_2291,N_2196,N_2167);
and U2292 (N_2292,N_2172,N_2111);
or U2293 (N_2293,N_2186,N_2119);
and U2294 (N_2294,N_2169,N_2004);
nand U2295 (N_2295,N_2161,N_2068);
nor U2296 (N_2296,N_2162,N_2016);
nand U2297 (N_2297,N_2003,N_2189);
nor U2298 (N_2298,N_2032,N_2067);
nand U2299 (N_2299,N_2130,N_2071);
or U2300 (N_2300,N_2173,N_2016);
xor U2301 (N_2301,N_2141,N_2013);
nand U2302 (N_2302,N_2094,N_2069);
nor U2303 (N_2303,N_2068,N_2104);
nand U2304 (N_2304,N_2156,N_2066);
or U2305 (N_2305,N_2091,N_2082);
and U2306 (N_2306,N_2002,N_2150);
or U2307 (N_2307,N_2002,N_2135);
and U2308 (N_2308,N_2032,N_2114);
or U2309 (N_2309,N_2016,N_2138);
nor U2310 (N_2310,N_2125,N_2179);
xnor U2311 (N_2311,N_2135,N_2051);
nand U2312 (N_2312,N_2059,N_2141);
nand U2313 (N_2313,N_2198,N_2090);
and U2314 (N_2314,N_2044,N_2008);
nor U2315 (N_2315,N_2103,N_2038);
xor U2316 (N_2316,N_2074,N_2183);
and U2317 (N_2317,N_2152,N_2168);
nand U2318 (N_2318,N_2049,N_2118);
nand U2319 (N_2319,N_2007,N_2088);
nand U2320 (N_2320,N_2026,N_2184);
or U2321 (N_2321,N_2154,N_2013);
xor U2322 (N_2322,N_2077,N_2062);
nand U2323 (N_2323,N_2046,N_2162);
and U2324 (N_2324,N_2122,N_2177);
nand U2325 (N_2325,N_2134,N_2030);
nor U2326 (N_2326,N_2120,N_2040);
nand U2327 (N_2327,N_2126,N_2035);
nand U2328 (N_2328,N_2024,N_2169);
or U2329 (N_2329,N_2103,N_2143);
xnor U2330 (N_2330,N_2042,N_2043);
or U2331 (N_2331,N_2091,N_2137);
and U2332 (N_2332,N_2187,N_2054);
or U2333 (N_2333,N_2073,N_2049);
and U2334 (N_2334,N_2142,N_2081);
and U2335 (N_2335,N_2035,N_2144);
and U2336 (N_2336,N_2182,N_2016);
or U2337 (N_2337,N_2007,N_2112);
and U2338 (N_2338,N_2021,N_2049);
nor U2339 (N_2339,N_2044,N_2052);
nor U2340 (N_2340,N_2025,N_2174);
xnor U2341 (N_2341,N_2080,N_2164);
nor U2342 (N_2342,N_2088,N_2065);
nand U2343 (N_2343,N_2030,N_2096);
and U2344 (N_2344,N_2032,N_2145);
nand U2345 (N_2345,N_2104,N_2053);
xnor U2346 (N_2346,N_2013,N_2155);
and U2347 (N_2347,N_2148,N_2124);
and U2348 (N_2348,N_2017,N_2113);
nand U2349 (N_2349,N_2025,N_2010);
or U2350 (N_2350,N_2043,N_2139);
nand U2351 (N_2351,N_2142,N_2045);
nor U2352 (N_2352,N_2190,N_2199);
nand U2353 (N_2353,N_2192,N_2163);
nor U2354 (N_2354,N_2143,N_2181);
nor U2355 (N_2355,N_2169,N_2047);
or U2356 (N_2356,N_2155,N_2048);
or U2357 (N_2357,N_2169,N_2150);
or U2358 (N_2358,N_2198,N_2140);
and U2359 (N_2359,N_2057,N_2149);
xor U2360 (N_2360,N_2186,N_2020);
and U2361 (N_2361,N_2050,N_2116);
nor U2362 (N_2362,N_2193,N_2084);
nand U2363 (N_2363,N_2051,N_2148);
and U2364 (N_2364,N_2084,N_2176);
nand U2365 (N_2365,N_2102,N_2022);
and U2366 (N_2366,N_2037,N_2170);
nor U2367 (N_2367,N_2088,N_2125);
xnor U2368 (N_2368,N_2094,N_2085);
nor U2369 (N_2369,N_2079,N_2031);
nor U2370 (N_2370,N_2183,N_2085);
nand U2371 (N_2371,N_2049,N_2038);
nand U2372 (N_2372,N_2160,N_2069);
nand U2373 (N_2373,N_2071,N_2008);
or U2374 (N_2374,N_2068,N_2029);
or U2375 (N_2375,N_2040,N_2131);
nand U2376 (N_2376,N_2092,N_2141);
and U2377 (N_2377,N_2138,N_2110);
and U2378 (N_2378,N_2120,N_2185);
nand U2379 (N_2379,N_2189,N_2179);
or U2380 (N_2380,N_2139,N_2046);
xnor U2381 (N_2381,N_2000,N_2119);
nor U2382 (N_2382,N_2105,N_2022);
nor U2383 (N_2383,N_2164,N_2129);
and U2384 (N_2384,N_2155,N_2041);
xnor U2385 (N_2385,N_2198,N_2102);
and U2386 (N_2386,N_2128,N_2107);
and U2387 (N_2387,N_2011,N_2134);
or U2388 (N_2388,N_2153,N_2195);
nand U2389 (N_2389,N_2175,N_2058);
nand U2390 (N_2390,N_2180,N_2045);
xnor U2391 (N_2391,N_2191,N_2065);
nor U2392 (N_2392,N_2119,N_2125);
nand U2393 (N_2393,N_2154,N_2171);
nor U2394 (N_2394,N_2187,N_2008);
or U2395 (N_2395,N_2093,N_2188);
nor U2396 (N_2396,N_2026,N_2009);
or U2397 (N_2397,N_2197,N_2078);
and U2398 (N_2398,N_2195,N_2181);
and U2399 (N_2399,N_2195,N_2101);
or U2400 (N_2400,N_2339,N_2269);
or U2401 (N_2401,N_2349,N_2201);
or U2402 (N_2402,N_2312,N_2305);
xnor U2403 (N_2403,N_2272,N_2381);
or U2404 (N_2404,N_2294,N_2225);
nand U2405 (N_2405,N_2355,N_2326);
nor U2406 (N_2406,N_2376,N_2316);
or U2407 (N_2407,N_2341,N_2394);
nand U2408 (N_2408,N_2315,N_2310);
and U2409 (N_2409,N_2287,N_2254);
nor U2410 (N_2410,N_2226,N_2369);
and U2411 (N_2411,N_2260,N_2237);
or U2412 (N_2412,N_2211,N_2290);
and U2413 (N_2413,N_2398,N_2219);
nor U2414 (N_2414,N_2368,N_2214);
or U2415 (N_2415,N_2324,N_2243);
or U2416 (N_2416,N_2302,N_2277);
and U2417 (N_2417,N_2357,N_2221);
nor U2418 (N_2418,N_2207,N_2220);
xor U2419 (N_2419,N_2328,N_2213);
nor U2420 (N_2420,N_2300,N_2329);
nor U2421 (N_2421,N_2227,N_2340);
and U2422 (N_2422,N_2318,N_2370);
and U2423 (N_2423,N_2388,N_2297);
nand U2424 (N_2424,N_2250,N_2224);
nand U2425 (N_2425,N_2395,N_2331);
nand U2426 (N_2426,N_2251,N_2330);
nand U2427 (N_2427,N_2333,N_2258);
and U2428 (N_2428,N_2230,N_2314);
nor U2429 (N_2429,N_2342,N_2375);
nand U2430 (N_2430,N_2255,N_2206);
nor U2431 (N_2431,N_2261,N_2262);
or U2432 (N_2432,N_2390,N_2229);
nor U2433 (N_2433,N_2292,N_2244);
nand U2434 (N_2434,N_2309,N_2374);
and U2435 (N_2435,N_2284,N_2320);
and U2436 (N_2436,N_2371,N_2285);
nand U2437 (N_2437,N_2233,N_2271);
and U2438 (N_2438,N_2210,N_2345);
nand U2439 (N_2439,N_2307,N_2313);
nand U2440 (N_2440,N_2325,N_2346);
and U2441 (N_2441,N_2264,N_2337);
nor U2442 (N_2442,N_2317,N_2336);
and U2443 (N_2443,N_2274,N_2391);
or U2444 (N_2444,N_2343,N_2378);
and U2445 (N_2445,N_2335,N_2279);
nand U2446 (N_2446,N_2200,N_2218);
or U2447 (N_2447,N_2319,N_2372);
nand U2448 (N_2448,N_2334,N_2383);
and U2449 (N_2449,N_2373,N_2273);
or U2450 (N_2450,N_2234,N_2270);
nand U2451 (N_2451,N_2281,N_2363);
nand U2452 (N_2452,N_2379,N_2240);
and U2453 (N_2453,N_2367,N_2321);
nor U2454 (N_2454,N_2205,N_2382);
nor U2455 (N_2455,N_2257,N_2298);
and U2456 (N_2456,N_2362,N_2323);
nand U2457 (N_2457,N_2286,N_2364);
and U2458 (N_2458,N_2223,N_2295);
nor U2459 (N_2459,N_2311,N_2392);
nor U2460 (N_2460,N_2386,N_2282);
nor U2461 (N_2461,N_2380,N_2275);
nor U2462 (N_2462,N_2288,N_2253);
nor U2463 (N_2463,N_2265,N_2266);
and U2464 (N_2464,N_2247,N_2338);
and U2465 (N_2465,N_2202,N_2289);
or U2466 (N_2466,N_2389,N_2301);
or U2467 (N_2467,N_2203,N_2353);
or U2468 (N_2468,N_2327,N_2365);
nand U2469 (N_2469,N_2216,N_2228);
nand U2470 (N_2470,N_2252,N_2209);
nand U2471 (N_2471,N_2354,N_2397);
or U2472 (N_2472,N_2242,N_2387);
nor U2473 (N_2473,N_2236,N_2280);
or U2474 (N_2474,N_2344,N_2238);
or U2475 (N_2475,N_2322,N_2351);
or U2476 (N_2476,N_2222,N_2246);
or U2477 (N_2477,N_2256,N_2268);
nand U2478 (N_2478,N_2249,N_2204);
nand U2479 (N_2479,N_2208,N_2293);
and U2480 (N_2480,N_2267,N_2215);
nand U2481 (N_2481,N_2259,N_2359);
or U2482 (N_2482,N_2347,N_2361);
or U2483 (N_2483,N_2348,N_2217);
and U2484 (N_2484,N_2291,N_2384);
or U2485 (N_2485,N_2360,N_2352);
and U2486 (N_2486,N_2396,N_2278);
xnor U2487 (N_2487,N_2304,N_2232);
and U2488 (N_2488,N_2385,N_2332);
nor U2489 (N_2489,N_2356,N_2299);
nand U2490 (N_2490,N_2283,N_2231);
or U2491 (N_2491,N_2358,N_2235);
or U2492 (N_2492,N_2366,N_2248);
nor U2493 (N_2493,N_2212,N_2241);
nor U2494 (N_2494,N_2239,N_2276);
nor U2495 (N_2495,N_2308,N_2350);
nor U2496 (N_2496,N_2263,N_2377);
nand U2497 (N_2497,N_2245,N_2393);
and U2498 (N_2498,N_2306,N_2296);
or U2499 (N_2499,N_2399,N_2303);
nand U2500 (N_2500,N_2348,N_2295);
and U2501 (N_2501,N_2299,N_2292);
and U2502 (N_2502,N_2320,N_2286);
and U2503 (N_2503,N_2308,N_2277);
nand U2504 (N_2504,N_2274,N_2320);
nor U2505 (N_2505,N_2312,N_2398);
nand U2506 (N_2506,N_2330,N_2391);
nand U2507 (N_2507,N_2206,N_2260);
and U2508 (N_2508,N_2242,N_2273);
or U2509 (N_2509,N_2304,N_2369);
or U2510 (N_2510,N_2384,N_2395);
nand U2511 (N_2511,N_2337,N_2349);
or U2512 (N_2512,N_2285,N_2229);
or U2513 (N_2513,N_2203,N_2336);
nand U2514 (N_2514,N_2356,N_2385);
nand U2515 (N_2515,N_2358,N_2279);
xor U2516 (N_2516,N_2255,N_2310);
nand U2517 (N_2517,N_2306,N_2348);
or U2518 (N_2518,N_2396,N_2348);
nand U2519 (N_2519,N_2248,N_2331);
nand U2520 (N_2520,N_2235,N_2350);
nand U2521 (N_2521,N_2264,N_2207);
and U2522 (N_2522,N_2390,N_2240);
and U2523 (N_2523,N_2316,N_2347);
and U2524 (N_2524,N_2203,N_2310);
nor U2525 (N_2525,N_2274,N_2330);
nor U2526 (N_2526,N_2320,N_2238);
nor U2527 (N_2527,N_2356,N_2275);
nor U2528 (N_2528,N_2383,N_2222);
nand U2529 (N_2529,N_2353,N_2322);
or U2530 (N_2530,N_2239,N_2283);
and U2531 (N_2531,N_2293,N_2385);
and U2532 (N_2532,N_2230,N_2355);
nor U2533 (N_2533,N_2330,N_2203);
nand U2534 (N_2534,N_2237,N_2231);
nand U2535 (N_2535,N_2284,N_2254);
or U2536 (N_2536,N_2219,N_2254);
nand U2537 (N_2537,N_2394,N_2245);
nor U2538 (N_2538,N_2307,N_2221);
or U2539 (N_2539,N_2317,N_2221);
xnor U2540 (N_2540,N_2331,N_2315);
or U2541 (N_2541,N_2306,N_2352);
and U2542 (N_2542,N_2233,N_2322);
nor U2543 (N_2543,N_2382,N_2310);
and U2544 (N_2544,N_2361,N_2371);
and U2545 (N_2545,N_2203,N_2321);
nand U2546 (N_2546,N_2290,N_2384);
nand U2547 (N_2547,N_2293,N_2383);
or U2548 (N_2548,N_2201,N_2234);
nor U2549 (N_2549,N_2375,N_2383);
nor U2550 (N_2550,N_2379,N_2204);
and U2551 (N_2551,N_2341,N_2380);
or U2552 (N_2552,N_2353,N_2282);
nor U2553 (N_2553,N_2353,N_2393);
or U2554 (N_2554,N_2280,N_2363);
nor U2555 (N_2555,N_2322,N_2212);
nor U2556 (N_2556,N_2392,N_2286);
and U2557 (N_2557,N_2292,N_2341);
nand U2558 (N_2558,N_2369,N_2292);
and U2559 (N_2559,N_2264,N_2229);
nand U2560 (N_2560,N_2379,N_2273);
and U2561 (N_2561,N_2238,N_2307);
nand U2562 (N_2562,N_2209,N_2255);
nand U2563 (N_2563,N_2264,N_2272);
and U2564 (N_2564,N_2369,N_2373);
nand U2565 (N_2565,N_2249,N_2247);
or U2566 (N_2566,N_2302,N_2333);
or U2567 (N_2567,N_2249,N_2210);
nor U2568 (N_2568,N_2367,N_2339);
or U2569 (N_2569,N_2386,N_2260);
xor U2570 (N_2570,N_2221,N_2283);
or U2571 (N_2571,N_2305,N_2349);
nand U2572 (N_2572,N_2271,N_2258);
xnor U2573 (N_2573,N_2335,N_2390);
and U2574 (N_2574,N_2279,N_2231);
nor U2575 (N_2575,N_2206,N_2247);
nand U2576 (N_2576,N_2266,N_2248);
nor U2577 (N_2577,N_2273,N_2339);
or U2578 (N_2578,N_2325,N_2394);
nor U2579 (N_2579,N_2346,N_2254);
nand U2580 (N_2580,N_2256,N_2284);
nor U2581 (N_2581,N_2228,N_2273);
nand U2582 (N_2582,N_2388,N_2331);
nand U2583 (N_2583,N_2292,N_2231);
or U2584 (N_2584,N_2302,N_2332);
and U2585 (N_2585,N_2261,N_2219);
nor U2586 (N_2586,N_2383,N_2373);
xnor U2587 (N_2587,N_2281,N_2276);
nand U2588 (N_2588,N_2361,N_2234);
or U2589 (N_2589,N_2385,N_2281);
or U2590 (N_2590,N_2275,N_2308);
nor U2591 (N_2591,N_2236,N_2365);
or U2592 (N_2592,N_2288,N_2330);
or U2593 (N_2593,N_2313,N_2378);
or U2594 (N_2594,N_2273,N_2322);
and U2595 (N_2595,N_2279,N_2384);
nor U2596 (N_2596,N_2269,N_2392);
or U2597 (N_2597,N_2302,N_2271);
nand U2598 (N_2598,N_2286,N_2273);
nor U2599 (N_2599,N_2314,N_2213);
nand U2600 (N_2600,N_2468,N_2532);
or U2601 (N_2601,N_2444,N_2569);
and U2602 (N_2602,N_2463,N_2575);
and U2603 (N_2603,N_2441,N_2531);
nand U2604 (N_2604,N_2427,N_2501);
or U2605 (N_2605,N_2402,N_2409);
nor U2606 (N_2606,N_2503,N_2457);
nand U2607 (N_2607,N_2488,N_2432);
nand U2608 (N_2608,N_2527,N_2418);
nor U2609 (N_2609,N_2589,N_2474);
nor U2610 (N_2610,N_2491,N_2573);
and U2611 (N_2611,N_2563,N_2526);
xor U2612 (N_2612,N_2570,N_2593);
or U2613 (N_2613,N_2449,N_2597);
nand U2614 (N_2614,N_2485,N_2492);
nand U2615 (N_2615,N_2464,N_2562);
or U2616 (N_2616,N_2410,N_2486);
or U2617 (N_2617,N_2401,N_2433);
and U2618 (N_2618,N_2590,N_2546);
nand U2619 (N_2619,N_2514,N_2524);
nor U2620 (N_2620,N_2484,N_2435);
nand U2621 (N_2621,N_2460,N_2549);
or U2622 (N_2622,N_2594,N_2477);
and U2623 (N_2623,N_2446,N_2447);
xor U2624 (N_2624,N_2541,N_2442);
nand U2625 (N_2625,N_2583,N_2480);
or U2626 (N_2626,N_2494,N_2574);
and U2627 (N_2627,N_2408,N_2415);
nand U2628 (N_2628,N_2538,N_2424);
nor U2629 (N_2629,N_2515,N_2499);
and U2630 (N_2630,N_2506,N_2553);
nand U2631 (N_2631,N_2542,N_2584);
nor U2632 (N_2632,N_2568,N_2596);
nand U2633 (N_2633,N_2496,N_2555);
nor U2634 (N_2634,N_2577,N_2564);
and U2635 (N_2635,N_2565,N_2417);
and U2636 (N_2636,N_2430,N_2426);
or U2637 (N_2637,N_2445,N_2411);
nand U2638 (N_2638,N_2523,N_2414);
and U2639 (N_2639,N_2529,N_2407);
nand U2640 (N_2640,N_2448,N_2483);
nand U2641 (N_2641,N_2475,N_2454);
nor U2642 (N_2642,N_2592,N_2455);
and U2643 (N_2643,N_2498,N_2516);
or U2644 (N_2644,N_2462,N_2412);
or U2645 (N_2645,N_2453,N_2511);
or U2646 (N_2646,N_2581,N_2481);
nand U2647 (N_2647,N_2478,N_2451);
and U2648 (N_2648,N_2466,N_2440);
nand U2649 (N_2649,N_2517,N_2434);
and U2650 (N_2650,N_2576,N_2487);
or U2651 (N_2651,N_2428,N_2582);
xnor U2652 (N_2652,N_2425,N_2560);
nor U2653 (N_2653,N_2545,N_2509);
and U2654 (N_2654,N_2572,N_2493);
nand U2655 (N_2655,N_2465,N_2458);
nor U2656 (N_2656,N_2482,N_2554);
nand U2657 (N_2657,N_2406,N_2547);
nand U2658 (N_2658,N_2537,N_2591);
nor U2659 (N_2659,N_2507,N_2467);
nor U2660 (N_2660,N_2400,N_2405);
and U2661 (N_2661,N_2530,N_2520);
or U2662 (N_2662,N_2479,N_2586);
nand U2663 (N_2663,N_2513,N_2490);
or U2664 (N_2664,N_2436,N_2571);
nand U2665 (N_2665,N_2557,N_2443);
nor U2666 (N_2666,N_2518,N_2512);
or U2667 (N_2667,N_2595,N_2534);
nand U2668 (N_2668,N_2450,N_2550);
or U2669 (N_2669,N_2533,N_2598);
xnor U2670 (N_2670,N_2566,N_2437);
nor U2671 (N_2671,N_2508,N_2422);
nor U2672 (N_2672,N_2495,N_2497);
and U2673 (N_2673,N_2471,N_2543);
nor U2674 (N_2674,N_2510,N_2588);
nand U2675 (N_2675,N_2579,N_2535);
nand U2676 (N_2676,N_2504,N_2431);
xor U2677 (N_2677,N_2540,N_2404);
nand U2678 (N_2678,N_2519,N_2423);
or U2679 (N_2679,N_2521,N_2544);
nand U2680 (N_2680,N_2552,N_2528);
and U2681 (N_2681,N_2419,N_2472);
or U2682 (N_2682,N_2551,N_2585);
nor U2683 (N_2683,N_2578,N_2429);
nor U2684 (N_2684,N_2438,N_2500);
nand U2685 (N_2685,N_2439,N_2473);
nand U2686 (N_2686,N_2522,N_2452);
nand U2687 (N_2687,N_2548,N_2416);
and U2688 (N_2688,N_2461,N_2525);
xnor U2689 (N_2689,N_2413,N_2502);
nand U2690 (N_2690,N_2599,N_2470);
xnor U2691 (N_2691,N_2505,N_2456);
nand U2692 (N_2692,N_2558,N_2489);
and U2693 (N_2693,N_2403,N_2459);
xnor U2694 (N_2694,N_2536,N_2421);
nor U2695 (N_2695,N_2539,N_2556);
or U2696 (N_2696,N_2567,N_2580);
or U2697 (N_2697,N_2476,N_2420);
nand U2698 (N_2698,N_2559,N_2469);
nor U2699 (N_2699,N_2587,N_2561);
nor U2700 (N_2700,N_2529,N_2547);
nand U2701 (N_2701,N_2570,N_2584);
nor U2702 (N_2702,N_2458,N_2456);
nor U2703 (N_2703,N_2472,N_2484);
nand U2704 (N_2704,N_2405,N_2446);
and U2705 (N_2705,N_2523,N_2469);
and U2706 (N_2706,N_2412,N_2591);
or U2707 (N_2707,N_2576,N_2442);
or U2708 (N_2708,N_2500,N_2538);
and U2709 (N_2709,N_2447,N_2547);
nor U2710 (N_2710,N_2522,N_2413);
or U2711 (N_2711,N_2562,N_2411);
and U2712 (N_2712,N_2434,N_2483);
nor U2713 (N_2713,N_2411,N_2465);
xor U2714 (N_2714,N_2517,N_2538);
or U2715 (N_2715,N_2599,N_2585);
and U2716 (N_2716,N_2422,N_2432);
and U2717 (N_2717,N_2567,N_2589);
nand U2718 (N_2718,N_2514,N_2534);
nand U2719 (N_2719,N_2455,N_2548);
nand U2720 (N_2720,N_2523,N_2470);
or U2721 (N_2721,N_2574,N_2565);
or U2722 (N_2722,N_2556,N_2468);
or U2723 (N_2723,N_2529,N_2421);
or U2724 (N_2724,N_2503,N_2597);
and U2725 (N_2725,N_2477,N_2550);
nand U2726 (N_2726,N_2520,N_2565);
and U2727 (N_2727,N_2579,N_2571);
nor U2728 (N_2728,N_2477,N_2426);
or U2729 (N_2729,N_2448,N_2420);
nand U2730 (N_2730,N_2511,N_2541);
nand U2731 (N_2731,N_2485,N_2465);
and U2732 (N_2732,N_2517,N_2591);
nand U2733 (N_2733,N_2571,N_2417);
or U2734 (N_2734,N_2452,N_2458);
or U2735 (N_2735,N_2543,N_2576);
or U2736 (N_2736,N_2417,N_2476);
nor U2737 (N_2737,N_2500,N_2528);
xor U2738 (N_2738,N_2578,N_2555);
nand U2739 (N_2739,N_2435,N_2442);
nor U2740 (N_2740,N_2454,N_2594);
nor U2741 (N_2741,N_2547,N_2577);
nand U2742 (N_2742,N_2404,N_2548);
xnor U2743 (N_2743,N_2582,N_2555);
or U2744 (N_2744,N_2407,N_2566);
nand U2745 (N_2745,N_2471,N_2556);
and U2746 (N_2746,N_2509,N_2595);
nor U2747 (N_2747,N_2599,N_2487);
nand U2748 (N_2748,N_2528,N_2490);
nor U2749 (N_2749,N_2530,N_2489);
or U2750 (N_2750,N_2472,N_2537);
nor U2751 (N_2751,N_2539,N_2555);
nor U2752 (N_2752,N_2498,N_2477);
nor U2753 (N_2753,N_2458,N_2472);
and U2754 (N_2754,N_2504,N_2452);
and U2755 (N_2755,N_2529,N_2578);
or U2756 (N_2756,N_2419,N_2465);
nor U2757 (N_2757,N_2523,N_2495);
or U2758 (N_2758,N_2507,N_2551);
and U2759 (N_2759,N_2484,N_2526);
and U2760 (N_2760,N_2521,N_2595);
nor U2761 (N_2761,N_2474,N_2433);
xor U2762 (N_2762,N_2530,N_2498);
or U2763 (N_2763,N_2494,N_2469);
and U2764 (N_2764,N_2530,N_2416);
or U2765 (N_2765,N_2430,N_2583);
nand U2766 (N_2766,N_2589,N_2408);
and U2767 (N_2767,N_2521,N_2432);
or U2768 (N_2768,N_2562,N_2475);
or U2769 (N_2769,N_2458,N_2568);
nand U2770 (N_2770,N_2570,N_2532);
or U2771 (N_2771,N_2430,N_2401);
nor U2772 (N_2772,N_2546,N_2481);
and U2773 (N_2773,N_2442,N_2463);
or U2774 (N_2774,N_2464,N_2520);
nor U2775 (N_2775,N_2463,N_2512);
and U2776 (N_2776,N_2511,N_2543);
xnor U2777 (N_2777,N_2438,N_2461);
and U2778 (N_2778,N_2571,N_2547);
nor U2779 (N_2779,N_2537,N_2511);
nor U2780 (N_2780,N_2501,N_2412);
and U2781 (N_2781,N_2433,N_2535);
or U2782 (N_2782,N_2496,N_2423);
and U2783 (N_2783,N_2564,N_2532);
nor U2784 (N_2784,N_2465,N_2537);
and U2785 (N_2785,N_2561,N_2552);
and U2786 (N_2786,N_2521,N_2400);
or U2787 (N_2787,N_2415,N_2403);
nor U2788 (N_2788,N_2479,N_2562);
or U2789 (N_2789,N_2408,N_2525);
or U2790 (N_2790,N_2541,N_2538);
nand U2791 (N_2791,N_2470,N_2493);
xor U2792 (N_2792,N_2521,N_2541);
nor U2793 (N_2793,N_2569,N_2449);
nand U2794 (N_2794,N_2591,N_2489);
and U2795 (N_2795,N_2409,N_2565);
nand U2796 (N_2796,N_2455,N_2507);
nor U2797 (N_2797,N_2531,N_2558);
or U2798 (N_2798,N_2472,N_2454);
or U2799 (N_2799,N_2503,N_2406);
nand U2800 (N_2800,N_2689,N_2785);
xor U2801 (N_2801,N_2677,N_2736);
nand U2802 (N_2802,N_2648,N_2760);
nor U2803 (N_2803,N_2656,N_2657);
and U2804 (N_2804,N_2733,N_2678);
nand U2805 (N_2805,N_2682,N_2680);
nand U2806 (N_2806,N_2691,N_2703);
nand U2807 (N_2807,N_2706,N_2730);
or U2808 (N_2808,N_2796,N_2718);
and U2809 (N_2809,N_2734,N_2647);
or U2810 (N_2810,N_2675,N_2600);
nor U2811 (N_2811,N_2726,N_2779);
or U2812 (N_2812,N_2731,N_2757);
xnor U2813 (N_2813,N_2741,N_2776);
and U2814 (N_2814,N_2719,N_2729);
xnor U2815 (N_2815,N_2694,N_2725);
and U2816 (N_2816,N_2684,N_2655);
and U2817 (N_2817,N_2609,N_2645);
or U2818 (N_2818,N_2636,N_2697);
or U2819 (N_2819,N_2753,N_2659);
nand U2820 (N_2820,N_2640,N_2637);
and U2821 (N_2821,N_2782,N_2607);
and U2822 (N_2822,N_2673,N_2763);
and U2823 (N_2823,N_2794,N_2781);
and U2824 (N_2824,N_2611,N_2769);
nor U2825 (N_2825,N_2668,N_2700);
or U2826 (N_2826,N_2759,N_2728);
nand U2827 (N_2827,N_2739,N_2625);
and U2828 (N_2828,N_2654,N_2617);
or U2829 (N_2829,N_2652,N_2798);
nand U2830 (N_2830,N_2662,N_2799);
and U2831 (N_2831,N_2755,N_2681);
nor U2832 (N_2832,N_2644,N_2727);
or U2833 (N_2833,N_2787,N_2724);
xor U2834 (N_2834,N_2768,N_2783);
and U2835 (N_2835,N_2714,N_2784);
nor U2836 (N_2836,N_2777,N_2751);
and U2837 (N_2837,N_2710,N_2674);
nor U2838 (N_2838,N_2616,N_2721);
nand U2839 (N_2839,N_2643,N_2650);
or U2840 (N_2840,N_2692,N_2702);
or U2841 (N_2841,N_2601,N_2651);
and U2842 (N_2842,N_2638,N_2797);
xor U2843 (N_2843,N_2778,N_2676);
xnor U2844 (N_2844,N_2606,N_2693);
and U2845 (N_2845,N_2790,N_2632);
and U2846 (N_2846,N_2610,N_2613);
nand U2847 (N_2847,N_2707,N_2788);
or U2848 (N_2848,N_2765,N_2618);
nor U2849 (N_2849,N_2716,N_2631);
and U2850 (N_2850,N_2634,N_2775);
or U2851 (N_2851,N_2671,N_2756);
nand U2852 (N_2852,N_2683,N_2602);
nand U2853 (N_2853,N_2738,N_2771);
nor U2854 (N_2854,N_2770,N_2639);
and U2855 (N_2855,N_2661,N_2764);
nand U2856 (N_2856,N_2791,N_2722);
and U2857 (N_2857,N_2774,N_2605);
or U2858 (N_2858,N_2704,N_2633);
xnor U2859 (N_2859,N_2687,N_2740);
nor U2860 (N_2860,N_2603,N_2629);
and U2861 (N_2861,N_2732,N_2641);
and U2862 (N_2862,N_2747,N_2630);
nor U2863 (N_2863,N_2743,N_2735);
nor U2864 (N_2864,N_2766,N_2686);
nand U2865 (N_2865,N_2646,N_2758);
or U2866 (N_2866,N_2663,N_2748);
nand U2867 (N_2867,N_2717,N_2695);
and U2868 (N_2868,N_2698,N_2628);
xor U2869 (N_2869,N_2786,N_2701);
and U2870 (N_2870,N_2793,N_2619);
and U2871 (N_2871,N_2622,N_2615);
or U2872 (N_2872,N_2709,N_2665);
nand U2873 (N_2873,N_2612,N_2664);
nor U2874 (N_2874,N_2754,N_2623);
and U2875 (N_2875,N_2749,N_2742);
and U2876 (N_2876,N_2627,N_2653);
or U2877 (N_2877,N_2620,N_2696);
nand U2878 (N_2878,N_2614,N_2708);
nor U2879 (N_2879,N_2745,N_2649);
nor U2880 (N_2880,N_2780,N_2737);
and U2881 (N_2881,N_2604,N_2772);
and U2882 (N_2882,N_2705,N_2688);
nand U2883 (N_2883,N_2746,N_2712);
nand U2884 (N_2884,N_2795,N_2744);
or U2885 (N_2885,N_2669,N_2711);
and U2886 (N_2886,N_2666,N_2690);
nor U2887 (N_2887,N_2608,N_2792);
xor U2888 (N_2888,N_2789,N_2762);
nand U2889 (N_2889,N_2667,N_2752);
or U2890 (N_2890,N_2761,N_2624);
nand U2891 (N_2891,N_2699,N_2670);
and U2892 (N_2892,N_2658,N_2642);
or U2893 (N_2893,N_2715,N_2621);
nor U2894 (N_2894,N_2679,N_2767);
nor U2895 (N_2895,N_2773,N_2723);
nand U2896 (N_2896,N_2626,N_2672);
and U2897 (N_2897,N_2685,N_2713);
nand U2898 (N_2898,N_2720,N_2750);
nor U2899 (N_2899,N_2660,N_2635);
and U2900 (N_2900,N_2658,N_2703);
nor U2901 (N_2901,N_2694,N_2776);
or U2902 (N_2902,N_2669,N_2667);
nor U2903 (N_2903,N_2617,N_2713);
or U2904 (N_2904,N_2685,N_2692);
and U2905 (N_2905,N_2691,N_2733);
or U2906 (N_2906,N_2621,N_2651);
nor U2907 (N_2907,N_2798,N_2678);
or U2908 (N_2908,N_2644,N_2702);
and U2909 (N_2909,N_2709,N_2754);
or U2910 (N_2910,N_2796,N_2664);
or U2911 (N_2911,N_2709,N_2619);
or U2912 (N_2912,N_2697,N_2712);
nand U2913 (N_2913,N_2726,N_2782);
or U2914 (N_2914,N_2646,N_2694);
nand U2915 (N_2915,N_2775,N_2696);
nand U2916 (N_2916,N_2689,N_2748);
or U2917 (N_2917,N_2764,N_2641);
nor U2918 (N_2918,N_2785,N_2767);
or U2919 (N_2919,N_2677,N_2669);
nand U2920 (N_2920,N_2630,N_2706);
nor U2921 (N_2921,N_2683,N_2675);
nand U2922 (N_2922,N_2644,N_2604);
and U2923 (N_2923,N_2765,N_2652);
nor U2924 (N_2924,N_2701,N_2705);
or U2925 (N_2925,N_2711,N_2778);
nand U2926 (N_2926,N_2645,N_2611);
and U2927 (N_2927,N_2718,N_2738);
or U2928 (N_2928,N_2615,N_2618);
nand U2929 (N_2929,N_2607,N_2765);
nand U2930 (N_2930,N_2645,N_2638);
nand U2931 (N_2931,N_2607,N_2769);
and U2932 (N_2932,N_2683,N_2785);
or U2933 (N_2933,N_2796,N_2673);
nor U2934 (N_2934,N_2697,N_2606);
nor U2935 (N_2935,N_2670,N_2671);
nand U2936 (N_2936,N_2738,N_2685);
nor U2937 (N_2937,N_2648,N_2766);
and U2938 (N_2938,N_2644,N_2690);
nor U2939 (N_2939,N_2759,N_2716);
nand U2940 (N_2940,N_2666,N_2729);
nor U2941 (N_2941,N_2782,N_2611);
nand U2942 (N_2942,N_2734,N_2707);
and U2943 (N_2943,N_2644,N_2739);
and U2944 (N_2944,N_2757,N_2666);
and U2945 (N_2945,N_2708,N_2642);
nor U2946 (N_2946,N_2758,N_2676);
nor U2947 (N_2947,N_2718,N_2628);
nand U2948 (N_2948,N_2683,N_2615);
or U2949 (N_2949,N_2798,N_2656);
nor U2950 (N_2950,N_2751,N_2647);
or U2951 (N_2951,N_2775,N_2631);
and U2952 (N_2952,N_2776,N_2748);
nor U2953 (N_2953,N_2798,N_2758);
and U2954 (N_2954,N_2767,N_2752);
xnor U2955 (N_2955,N_2792,N_2747);
or U2956 (N_2956,N_2655,N_2622);
nor U2957 (N_2957,N_2692,N_2701);
nor U2958 (N_2958,N_2799,N_2732);
nand U2959 (N_2959,N_2735,N_2616);
and U2960 (N_2960,N_2608,N_2758);
nand U2961 (N_2961,N_2632,N_2652);
nor U2962 (N_2962,N_2711,N_2772);
nor U2963 (N_2963,N_2779,N_2660);
and U2964 (N_2964,N_2747,N_2741);
or U2965 (N_2965,N_2770,N_2756);
nand U2966 (N_2966,N_2674,N_2705);
xnor U2967 (N_2967,N_2692,N_2636);
or U2968 (N_2968,N_2636,N_2624);
nand U2969 (N_2969,N_2739,N_2603);
or U2970 (N_2970,N_2689,N_2791);
nor U2971 (N_2971,N_2713,N_2739);
nand U2972 (N_2972,N_2749,N_2796);
nand U2973 (N_2973,N_2655,N_2751);
and U2974 (N_2974,N_2679,N_2659);
and U2975 (N_2975,N_2735,N_2732);
or U2976 (N_2976,N_2788,N_2669);
or U2977 (N_2977,N_2773,N_2677);
and U2978 (N_2978,N_2730,N_2692);
xnor U2979 (N_2979,N_2726,N_2729);
nor U2980 (N_2980,N_2601,N_2783);
xnor U2981 (N_2981,N_2609,N_2766);
nand U2982 (N_2982,N_2773,N_2760);
and U2983 (N_2983,N_2608,N_2719);
nand U2984 (N_2984,N_2682,N_2775);
and U2985 (N_2985,N_2793,N_2622);
and U2986 (N_2986,N_2759,N_2610);
and U2987 (N_2987,N_2710,N_2771);
or U2988 (N_2988,N_2639,N_2662);
or U2989 (N_2989,N_2715,N_2703);
or U2990 (N_2990,N_2791,N_2691);
or U2991 (N_2991,N_2728,N_2797);
nor U2992 (N_2992,N_2790,N_2782);
nand U2993 (N_2993,N_2710,N_2648);
and U2994 (N_2994,N_2787,N_2696);
or U2995 (N_2995,N_2706,N_2715);
nor U2996 (N_2996,N_2702,N_2788);
nor U2997 (N_2997,N_2776,N_2649);
and U2998 (N_2998,N_2752,N_2694);
nor U2999 (N_2999,N_2797,N_2686);
and U3000 (N_3000,N_2958,N_2898);
nand U3001 (N_3001,N_2830,N_2906);
nand U3002 (N_3002,N_2977,N_2846);
nand U3003 (N_3003,N_2952,N_2911);
and U3004 (N_3004,N_2812,N_2818);
and U3005 (N_3005,N_2996,N_2983);
and U3006 (N_3006,N_2974,N_2847);
nor U3007 (N_3007,N_2832,N_2934);
and U3008 (N_3008,N_2853,N_2935);
and U3009 (N_3009,N_2834,N_2875);
nor U3010 (N_3010,N_2872,N_2884);
xnor U3011 (N_3011,N_2950,N_2960);
nor U3012 (N_3012,N_2809,N_2863);
nand U3013 (N_3013,N_2838,N_2989);
nor U3014 (N_3014,N_2870,N_2929);
and U3015 (N_3015,N_2959,N_2821);
nand U3016 (N_3016,N_2808,N_2909);
nand U3017 (N_3017,N_2997,N_2990);
xor U3018 (N_3018,N_2845,N_2860);
or U3019 (N_3019,N_2877,N_2856);
xor U3020 (N_3020,N_2948,N_2970);
nand U3021 (N_3021,N_2849,N_2878);
nand U3022 (N_3022,N_2865,N_2936);
nand U3023 (N_3023,N_2814,N_2888);
or U3024 (N_3024,N_2973,N_2918);
xnor U3025 (N_3025,N_2994,N_2859);
or U3026 (N_3026,N_2943,N_2927);
and U3027 (N_3027,N_2882,N_2879);
nor U3028 (N_3028,N_2967,N_2984);
nor U3029 (N_3029,N_2925,N_2941);
nand U3030 (N_3030,N_2914,N_2858);
nand U3031 (N_3031,N_2968,N_2889);
nand U3032 (N_3032,N_2833,N_2905);
nand U3033 (N_3033,N_2811,N_2823);
and U3034 (N_3034,N_2864,N_2907);
xnor U3035 (N_3035,N_2890,N_2944);
and U3036 (N_3036,N_2981,N_2947);
nor U3037 (N_3037,N_2966,N_2957);
and U3038 (N_3038,N_2988,N_2810);
or U3039 (N_3039,N_2901,N_2922);
nor U3040 (N_3040,N_2937,N_2949);
nor U3041 (N_3041,N_2807,N_2965);
and U3042 (N_3042,N_2822,N_2825);
and U3043 (N_3043,N_2908,N_2826);
nand U3044 (N_3044,N_2978,N_2939);
nor U3045 (N_3045,N_2940,N_2931);
and U3046 (N_3046,N_2992,N_2816);
or U3047 (N_3047,N_2850,N_2902);
nor U3048 (N_3048,N_2956,N_2962);
and U3049 (N_3049,N_2913,N_2801);
and U3050 (N_3050,N_2857,N_2837);
and U3051 (N_3051,N_2932,N_2971);
nor U3052 (N_3052,N_2806,N_2903);
or U3053 (N_3053,N_2881,N_2964);
nor U3054 (N_3054,N_2919,N_2891);
or U3055 (N_3055,N_2924,N_2910);
and U3056 (N_3056,N_2900,N_2915);
and U3057 (N_3057,N_2861,N_2986);
and U3058 (N_3058,N_2840,N_2897);
nor U3059 (N_3059,N_2800,N_2923);
nor U3060 (N_3060,N_2876,N_2895);
nand U3061 (N_3061,N_2855,N_2928);
and U3062 (N_3062,N_2843,N_2862);
xor U3063 (N_3063,N_2987,N_2802);
nand U3064 (N_3064,N_2969,N_2815);
nor U3065 (N_3065,N_2893,N_2824);
nor U3066 (N_3066,N_2839,N_2813);
or U3067 (N_3067,N_2921,N_2883);
or U3068 (N_3068,N_2955,N_2896);
and U3069 (N_3069,N_2887,N_2842);
and U3070 (N_3070,N_2972,N_2844);
nor U3071 (N_3071,N_2993,N_2835);
and U3072 (N_3072,N_2999,N_2828);
nor U3073 (N_3073,N_2942,N_2836);
nor U3074 (N_3074,N_2885,N_2980);
nand U3075 (N_3075,N_2874,N_2873);
and U3076 (N_3076,N_2912,N_2841);
and U3077 (N_3077,N_2926,N_2854);
xor U3078 (N_3078,N_2886,N_2829);
or U3079 (N_3079,N_2985,N_2945);
nand U3080 (N_3080,N_2946,N_2904);
nor U3081 (N_3081,N_2961,N_2998);
nand U3082 (N_3082,N_2976,N_2963);
and U3083 (N_3083,N_2916,N_2868);
xnor U3084 (N_3084,N_2871,N_2979);
nor U3085 (N_3085,N_2938,N_2852);
or U3086 (N_3086,N_2869,N_2995);
nand U3087 (N_3087,N_2848,N_2803);
xor U3088 (N_3088,N_2917,N_2899);
and U3089 (N_3089,N_2867,N_2819);
nor U3090 (N_3090,N_2805,N_2827);
nor U3091 (N_3091,N_2866,N_2951);
and U3092 (N_3092,N_2930,N_2820);
or U3093 (N_3093,N_2991,N_2851);
or U3094 (N_3094,N_2831,N_2892);
and U3095 (N_3095,N_2982,N_2954);
nand U3096 (N_3096,N_2894,N_2975);
and U3097 (N_3097,N_2804,N_2953);
and U3098 (N_3098,N_2880,N_2933);
nor U3099 (N_3099,N_2920,N_2817);
nor U3100 (N_3100,N_2960,N_2892);
nand U3101 (N_3101,N_2818,N_2911);
nand U3102 (N_3102,N_2989,N_2917);
nand U3103 (N_3103,N_2956,N_2929);
or U3104 (N_3104,N_2994,N_2988);
nand U3105 (N_3105,N_2857,N_2976);
and U3106 (N_3106,N_2981,N_2984);
nor U3107 (N_3107,N_2947,N_2848);
nand U3108 (N_3108,N_2971,N_2876);
nand U3109 (N_3109,N_2844,N_2971);
nand U3110 (N_3110,N_2944,N_2803);
or U3111 (N_3111,N_2800,N_2998);
xor U3112 (N_3112,N_2987,N_2925);
and U3113 (N_3113,N_2916,N_2832);
and U3114 (N_3114,N_2963,N_2917);
or U3115 (N_3115,N_2807,N_2941);
and U3116 (N_3116,N_2979,N_2997);
and U3117 (N_3117,N_2892,N_2828);
nand U3118 (N_3118,N_2840,N_2913);
nand U3119 (N_3119,N_2835,N_2827);
and U3120 (N_3120,N_2835,N_2919);
xor U3121 (N_3121,N_2895,N_2841);
and U3122 (N_3122,N_2881,N_2882);
nor U3123 (N_3123,N_2838,N_2801);
nand U3124 (N_3124,N_2991,N_2830);
or U3125 (N_3125,N_2804,N_2930);
and U3126 (N_3126,N_2848,N_2847);
or U3127 (N_3127,N_2897,N_2916);
nand U3128 (N_3128,N_2947,N_2860);
nor U3129 (N_3129,N_2878,N_2911);
nor U3130 (N_3130,N_2825,N_2902);
nand U3131 (N_3131,N_2881,N_2896);
and U3132 (N_3132,N_2802,N_2889);
and U3133 (N_3133,N_2917,N_2935);
and U3134 (N_3134,N_2883,N_2926);
nand U3135 (N_3135,N_2878,N_2833);
nand U3136 (N_3136,N_2872,N_2953);
or U3137 (N_3137,N_2810,N_2841);
or U3138 (N_3138,N_2822,N_2820);
nand U3139 (N_3139,N_2967,N_2827);
nand U3140 (N_3140,N_2838,N_2984);
and U3141 (N_3141,N_2871,N_2976);
xor U3142 (N_3142,N_2997,N_2819);
nor U3143 (N_3143,N_2841,N_2921);
xnor U3144 (N_3144,N_2937,N_2896);
xnor U3145 (N_3145,N_2902,N_2905);
or U3146 (N_3146,N_2897,N_2898);
or U3147 (N_3147,N_2849,N_2848);
xor U3148 (N_3148,N_2881,N_2968);
or U3149 (N_3149,N_2974,N_2975);
or U3150 (N_3150,N_2976,N_2822);
nor U3151 (N_3151,N_2944,N_2992);
or U3152 (N_3152,N_2968,N_2802);
nor U3153 (N_3153,N_2817,N_2901);
nor U3154 (N_3154,N_2945,N_2814);
or U3155 (N_3155,N_2982,N_2983);
and U3156 (N_3156,N_2981,N_2930);
nand U3157 (N_3157,N_2813,N_2853);
nor U3158 (N_3158,N_2967,N_2896);
nor U3159 (N_3159,N_2992,N_2990);
nand U3160 (N_3160,N_2977,N_2978);
and U3161 (N_3161,N_2846,N_2911);
xor U3162 (N_3162,N_2845,N_2893);
xor U3163 (N_3163,N_2971,N_2828);
nor U3164 (N_3164,N_2897,N_2948);
or U3165 (N_3165,N_2961,N_2806);
nor U3166 (N_3166,N_2872,N_2979);
or U3167 (N_3167,N_2945,N_2976);
and U3168 (N_3168,N_2953,N_2962);
nand U3169 (N_3169,N_2922,N_2845);
nand U3170 (N_3170,N_2804,N_2954);
xor U3171 (N_3171,N_2846,N_2865);
nor U3172 (N_3172,N_2822,N_2906);
or U3173 (N_3173,N_2895,N_2972);
xor U3174 (N_3174,N_2888,N_2913);
or U3175 (N_3175,N_2804,N_2872);
or U3176 (N_3176,N_2910,N_2888);
nor U3177 (N_3177,N_2868,N_2939);
xor U3178 (N_3178,N_2965,N_2985);
or U3179 (N_3179,N_2852,N_2877);
nand U3180 (N_3180,N_2807,N_2961);
and U3181 (N_3181,N_2950,N_2985);
nor U3182 (N_3182,N_2867,N_2829);
nand U3183 (N_3183,N_2960,N_2906);
nor U3184 (N_3184,N_2952,N_2995);
nor U3185 (N_3185,N_2899,N_2808);
nor U3186 (N_3186,N_2986,N_2857);
and U3187 (N_3187,N_2883,N_2808);
and U3188 (N_3188,N_2854,N_2829);
and U3189 (N_3189,N_2943,N_2870);
nand U3190 (N_3190,N_2820,N_2805);
or U3191 (N_3191,N_2872,N_2824);
and U3192 (N_3192,N_2852,N_2835);
nand U3193 (N_3193,N_2930,N_2862);
and U3194 (N_3194,N_2937,N_2883);
xor U3195 (N_3195,N_2805,N_2962);
nand U3196 (N_3196,N_2949,N_2884);
or U3197 (N_3197,N_2963,N_2897);
or U3198 (N_3198,N_2936,N_2990);
or U3199 (N_3199,N_2976,N_2952);
nor U3200 (N_3200,N_3096,N_3046);
nand U3201 (N_3201,N_3159,N_3006);
or U3202 (N_3202,N_3131,N_3011);
nor U3203 (N_3203,N_3118,N_3008);
and U3204 (N_3204,N_3107,N_3061);
and U3205 (N_3205,N_3149,N_3026);
nand U3206 (N_3206,N_3122,N_3100);
and U3207 (N_3207,N_3174,N_3013);
nor U3208 (N_3208,N_3058,N_3111);
nand U3209 (N_3209,N_3037,N_3195);
or U3210 (N_3210,N_3151,N_3005);
nand U3211 (N_3211,N_3190,N_3176);
nor U3212 (N_3212,N_3080,N_3041);
or U3213 (N_3213,N_3101,N_3106);
nor U3214 (N_3214,N_3139,N_3145);
nand U3215 (N_3215,N_3133,N_3084);
or U3216 (N_3216,N_3188,N_3171);
and U3217 (N_3217,N_3091,N_3082);
and U3218 (N_3218,N_3124,N_3199);
or U3219 (N_3219,N_3040,N_3023);
and U3220 (N_3220,N_3088,N_3090);
or U3221 (N_3221,N_3198,N_3194);
or U3222 (N_3222,N_3057,N_3170);
and U3223 (N_3223,N_3132,N_3183);
or U3224 (N_3224,N_3113,N_3087);
or U3225 (N_3225,N_3186,N_3126);
nor U3226 (N_3226,N_3014,N_3157);
nand U3227 (N_3227,N_3116,N_3038);
or U3228 (N_3228,N_3044,N_3189);
nor U3229 (N_3229,N_3004,N_3079);
nor U3230 (N_3230,N_3155,N_3108);
nand U3231 (N_3231,N_3102,N_3127);
xnor U3232 (N_3232,N_3056,N_3003);
nor U3233 (N_3233,N_3172,N_3016);
xnor U3234 (N_3234,N_3134,N_3192);
or U3235 (N_3235,N_3156,N_3060);
or U3236 (N_3236,N_3062,N_3121);
nor U3237 (N_3237,N_3064,N_3020);
and U3238 (N_3238,N_3077,N_3076);
nor U3239 (N_3239,N_3138,N_3068);
xnor U3240 (N_3240,N_3150,N_3117);
nor U3241 (N_3241,N_3146,N_3018);
xnor U3242 (N_3242,N_3162,N_3153);
nor U3243 (N_3243,N_3009,N_3180);
or U3244 (N_3244,N_3182,N_3109);
nor U3245 (N_3245,N_3161,N_3184);
nand U3246 (N_3246,N_3065,N_3066);
nand U3247 (N_3247,N_3166,N_3035);
and U3248 (N_3248,N_3104,N_3051);
nand U3249 (N_3249,N_3179,N_3167);
or U3250 (N_3250,N_3094,N_3019);
and U3251 (N_3251,N_3073,N_3081);
and U3252 (N_3252,N_3070,N_3095);
nand U3253 (N_3253,N_3173,N_3142);
and U3254 (N_3254,N_3007,N_3158);
and U3255 (N_3255,N_3093,N_3032);
nor U3256 (N_3256,N_3181,N_3053);
nand U3257 (N_3257,N_3017,N_3169);
or U3258 (N_3258,N_3141,N_3120);
or U3259 (N_3259,N_3074,N_3078);
nor U3260 (N_3260,N_3030,N_3130);
and U3261 (N_3261,N_3175,N_3148);
nor U3262 (N_3262,N_3123,N_3164);
nand U3263 (N_3263,N_3027,N_3128);
or U3264 (N_3264,N_3152,N_3031);
or U3265 (N_3265,N_3002,N_3000);
and U3266 (N_3266,N_3129,N_3136);
and U3267 (N_3267,N_3097,N_3045);
and U3268 (N_3268,N_3054,N_3177);
and U3269 (N_3269,N_3024,N_3034);
and U3270 (N_3270,N_3025,N_3193);
or U3271 (N_3271,N_3039,N_3168);
nand U3272 (N_3272,N_3110,N_3028);
and U3273 (N_3273,N_3050,N_3021);
or U3274 (N_3274,N_3143,N_3144);
xor U3275 (N_3275,N_3185,N_3059);
nor U3276 (N_3276,N_3047,N_3135);
nand U3277 (N_3277,N_3071,N_3187);
nor U3278 (N_3278,N_3114,N_3015);
nor U3279 (N_3279,N_3012,N_3165);
nand U3280 (N_3280,N_3160,N_3036);
nor U3281 (N_3281,N_3063,N_3085);
and U3282 (N_3282,N_3052,N_3049);
nor U3283 (N_3283,N_3163,N_3103);
or U3284 (N_3284,N_3098,N_3010);
and U3285 (N_3285,N_3029,N_3055);
nor U3286 (N_3286,N_3042,N_3086);
nor U3287 (N_3287,N_3022,N_3119);
xor U3288 (N_3288,N_3112,N_3001);
and U3289 (N_3289,N_3043,N_3197);
nor U3290 (N_3290,N_3105,N_3196);
nor U3291 (N_3291,N_3137,N_3140);
nor U3292 (N_3292,N_3178,N_3125);
or U3293 (N_3293,N_3115,N_3154);
xor U3294 (N_3294,N_3083,N_3147);
nor U3295 (N_3295,N_3048,N_3033);
nor U3296 (N_3296,N_3089,N_3075);
nor U3297 (N_3297,N_3067,N_3191);
nand U3298 (N_3298,N_3072,N_3069);
nor U3299 (N_3299,N_3099,N_3092);
nor U3300 (N_3300,N_3191,N_3114);
or U3301 (N_3301,N_3072,N_3160);
nor U3302 (N_3302,N_3064,N_3157);
nor U3303 (N_3303,N_3101,N_3086);
nor U3304 (N_3304,N_3127,N_3105);
and U3305 (N_3305,N_3012,N_3018);
nor U3306 (N_3306,N_3061,N_3098);
nand U3307 (N_3307,N_3052,N_3085);
nand U3308 (N_3308,N_3059,N_3094);
or U3309 (N_3309,N_3064,N_3189);
xnor U3310 (N_3310,N_3047,N_3067);
nand U3311 (N_3311,N_3104,N_3137);
nand U3312 (N_3312,N_3041,N_3025);
nand U3313 (N_3313,N_3028,N_3040);
xor U3314 (N_3314,N_3120,N_3078);
or U3315 (N_3315,N_3192,N_3011);
or U3316 (N_3316,N_3026,N_3059);
and U3317 (N_3317,N_3141,N_3008);
nand U3318 (N_3318,N_3120,N_3087);
or U3319 (N_3319,N_3117,N_3039);
nor U3320 (N_3320,N_3062,N_3035);
or U3321 (N_3321,N_3152,N_3046);
or U3322 (N_3322,N_3088,N_3066);
nor U3323 (N_3323,N_3004,N_3105);
nand U3324 (N_3324,N_3008,N_3191);
nor U3325 (N_3325,N_3157,N_3100);
nor U3326 (N_3326,N_3059,N_3071);
nand U3327 (N_3327,N_3081,N_3079);
or U3328 (N_3328,N_3188,N_3118);
nand U3329 (N_3329,N_3180,N_3112);
and U3330 (N_3330,N_3159,N_3090);
and U3331 (N_3331,N_3043,N_3012);
and U3332 (N_3332,N_3019,N_3084);
or U3333 (N_3333,N_3029,N_3151);
xnor U3334 (N_3334,N_3182,N_3151);
or U3335 (N_3335,N_3143,N_3102);
and U3336 (N_3336,N_3107,N_3038);
or U3337 (N_3337,N_3056,N_3135);
xor U3338 (N_3338,N_3078,N_3119);
nand U3339 (N_3339,N_3066,N_3074);
nand U3340 (N_3340,N_3005,N_3117);
or U3341 (N_3341,N_3093,N_3152);
or U3342 (N_3342,N_3051,N_3070);
and U3343 (N_3343,N_3072,N_3019);
or U3344 (N_3344,N_3145,N_3117);
or U3345 (N_3345,N_3031,N_3090);
and U3346 (N_3346,N_3031,N_3198);
xnor U3347 (N_3347,N_3186,N_3055);
and U3348 (N_3348,N_3111,N_3154);
xor U3349 (N_3349,N_3074,N_3052);
nor U3350 (N_3350,N_3158,N_3124);
and U3351 (N_3351,N_3144,N_3105);
and U3352 (N_3352,N_3013,N_3195);
and U3353 (N_3353,N_3119,N_3069);
or U3354 (N_3354,N_3048,N_3183);
nand U3355 (N_3355,N_3138,N_3133);
nor U3356 (N_3356,N_3129,N_3147);
xnor U3357 (N_3357,N_3089,N_3193);
nand U3358 (N_3358,N_3076,N_3196);
or U3359 (N_3359,N_3136,N_3032);
or U3360 (N_3360,N_3184,N_3179);
xor U3361 (N_3361,N_3080,N_3118);
nor U3362 (N_3362,N_3101,N_3156);
xnor U3363 (N_3363,N_3103,N_3156);
or U3364 (N_3364,N_3124,N_3052);
xor U3365 (N_3365,N_3162,N_3012);
nor U3366 (N_3366,N_3063,N_3021);
nor U3367 (N_3367,N_3006,N_3109);
or U3368 (N_3368,N_3005,N_3015);
or U3369 (N_3369,N_3048,N_3036);
nand U3370 (N_3370,N_3168,N_3146);
or U3371 (N_3371,N_3081,N_3020);
nor U3372 (N_3372,N_3090,N_3177);
nand U3373 (N_3373,N_3070,N_3012);
nand U3374 (N_3374,N_3127,N_3038);
nor U3375 (N_3375,N_3155,N_3103);
or U3376 (N_3376,N_3060,N_3135);
nand U3377 (N_3377,N_3187,N_3122);
and U3378 (N_3378,N_3096,N_3036);
and U3379 (N_3379,N_3153,N_3053);
nor U3380 (N_3380,N_3069,N_3135);
nor U3381 (N_3381,N_3007,N_3148);
and U3382 (N_3382,N_3026,N_3065);
or U3383 (N_3383,N_3098,N_3181);
nand U3384 (N_3384,N_3071,N_3146);
or U3385 (N_3385,N_3179,N_3122);
nand U3386 (N_3386,N_3116,N_3114);
nor U3387 (N_3387,N_3173,N_3051);
nand U3388 (N_3388,N_3171,N_3098);
nor U3389 (N_3389,N_3008,N_3108);
or U3390 (N_3390,N_3106,N_3130);
or U3391 (N_3391,N_3151,N_3138);
and U3392 (N_3392,N_3179,N_3020);
or U3393 (N_3393,N_3038,N_3180);
and U3394 (N_3394,N_3054,N_3068);
nand U3395 (N_3395,N_3144,N_3006);
or U3396 (N_3396,N_3138,N_3196);
and U3397 (N_3397,N_3105,N_3176);
xor U3398 (N_3398,N_3030,N_3118);
nor U3399 (N_3399,N_3130,N_3109);
nand U3400 (N_3400,N_3234,N_3213);
nand U3401 (N_3401,N_3245,N_3385);
xnor U3402 (N_3402,N_3229,N_3310);
nand U3403 (N_3403,N_3386,N_3216);
and U3404 (N_3404,N_3241,N_3200);
nand U3405 (N_3405,N_3206,N_3299);
or U3406 (N_3406,N_3355,N_3357);
nor U3407 (N_3407,N_3228,N_3373);
nor U3408 (N_3408,N_3350,N_3238);
nor U3409 (N_3409,N_3290,N_3361);
or U3410 (N_3410,N_3230,N_3237);
and U3411 (N_3411,N_3278,N_3204);
nor U3412 (N_3412,N_3332,N_3240);
nor U3413 (N_3413,N_3390,N_3320);
xnor U3414 (N_3414,N_3341,N_3340);
nand U3415 (N_3415,N_3377,N_3263);
nand U3416 (N_3416,N_3287,N_3369);
and U3417 (N_3417,N_3217,N_3335);
or U3418 (N_3418,N_3328,N_3397);
or U3419 (N_3419,N_3313,N_3382);
nor U3420 (N_3420,N_3211,N_3391);
or U3421 (N_3421,N_3317,N_3265);
or U3422 (N_3422,N_3381,N_3285);
or U3423 (N_3423,N_3318,N_3380);
xor U3424 (N_3424,N_3275,N_3280);
nor U3425 (N_3425,N_3333,N_3337);
xnor U3426 (N_3426,N_3349,N_3288);
and U3427 (N_3427,N_3364,N_3254);
or U3428 (N_3428,N_3376,N_3273);
and U3429 (N_3429,N_3319,N_3259);
or U3430 (N_3430,N_3272,N_3243);
nor U3431 (N_3431,N_3306,N_3329);
or U3432 (N_3432,N_3345,N_3283);
nor U3433 (N_3433,N_3388,N_3284);
or U3434 (N_3434,N_3304,N_3221);
or U3435 (N_3435,N_3220,N_3356);
xnor U3436 (N_3436,N_3399,N_3247);
xnor U3437 (N_3437,N_3365,N_3351);
or U3438 (N_3438,N_3311,N_3224);
and U3439 (N_3439,N_3251,N_3294);
nor U3440 (N_3440,N_3363,N_3322);
or U3441 (N_3441,N_3253,N_3286);
nor U3442 (N_3442,N_3352,N_3316);
xnor U3443 (N_3443,N_3256,N_3279);
or U3444 (N_3444,N_3342,N_3331);
and U3445 (N_3445,N_3362,N_3210);
nand U3446 (N_3446,N_3274,N_3346);
or U3447 (N_3447,N_3338,N_3249);
nor U3448 (N_3448,N_3270,N_3225);
nor U3449 (N_3449,N_3354,N_3242);
and U3450 (N_3450,N_3326,N_3314);
nor U3451 (N_3451,N_3336,N_3323);
and U3452 (N_3452,N_3269,N_3293);
and U3453 (N_3453,N_3375,N_3261);
or U3454 (N_3454,N_3348,N_3396);
and U3455 (N_3455,N_3343,N_3393);
nand U3456 (N_3456,N_3218,N_3360);
or U3457 (N_3457,N_3372,N_3392);
and U3458 (N_3458,N_3233,N_3308);
nor U3459 (N_3459,N_3394,N_3267);
xor U3460 (N_3460,N_3383,N_3389);
nand U3461 (N_3461,N_3276,N_3260);
or U3462 (N_3462,N_3207,N_3324);
and U3463 (N_3463,N_3203,N_3258);
nand U3464 (N_3464,N_3277,N_3297);
and U3465 (N_3465,N_3370,N_3300);
or U3466 (N_3466,N_3339,N_3327);
nand U3467 (N_3467,N_3374,N_3371);
nor U3468 (N_3468,N_3387,N_3295);
nand U3469 (N_3469,N_3222,N_3264);
and U3470 (N_3470,N_3305,N_3321);
xnor U3471 (N_3471,N_3208,N_3303);
or U3472 (N_3472,N_3271,N_3291);
and U3473 (N_3473,N_3367,N_3359);
and U3474 (N_3474,N_3257,N_3255);
nand U3475 (N_3475,N_3301,N_3366);
or U3476 (N_3476,N_3282,N_3289);
and U3477 (N_3477,N_3398,N_3268);
nor U3478 (N_3478,N_3201,N_3231);
nand U3479 (N_3479,N_3292,N_3325);
nor U3480 (N_3480,N_3239,N_3296);
xor U3481 (N_3481,N_3212,N_3209);
xnor U3482 (N_3482,N_3202,N_3236);
nand U3483 (N_3483,N_3315,N_3309);
or U3484 (N_3484,N_3232,N_3298);
and U3485 (N_3485,N_3378,N_3246);
xnor U3486 (N_3486,N_3227,N_3353);
nor U3487 (N_3487,N_3266,N_3252);
or U3488 (N_3488,N_3244,N_3223);
nand U3489 (N_3489,N_3205,N_3235);
or U3490 (N_3490,N_3226,N_3307);
xnor U3491 (N_3491,N_3302,N_3214);
or U3492 (N_3492,N_3250,N_3262);
nand U3493 (N_3493,N_3344,N_3219);
or U3494 (N_3494,N_3347,N_3358);
nand U3495 (N_3495,N_3384,N_3215);
nor U3496 (N_3496,N_3330,N_3368);
and U3497 (N_3497,N_3395,N_3379);
or U3498 (N_3498,N_3248,N_3281);
nor U3499 (N_3499,N_3312,N_3334);
and U3500 (N_3500,N_3349,N_3292);
nand U3501 (N_3501,N_3325,N_3216);
nand U3502 (N_3502,N_3251,N_3224);
or U3503 (N_3503,N_3362,N_3374);
and U3504 (N_3504,N_3350,N_3308);
nand U3505 (N_3505,N_3371,N_3373);
nand U3506 (N_3506,N_3300,N_3289);
or U3507 (N_3507,N_3325,N_3352);
or U3508 (N_3508,N_3354,N_3376);
nor U3509 (N_3509,N_3292,N_3254);
nor U3510 (N_3510,N_3315,N_3352);
and U3511 (N_3511,N_3215,N_3290);
nand U3512 (N_3512,N_3352,N_3278);
nor U3513 (N_3513,N_3277,N_3317);
and U3514 (N_3514,N_3331,N_3333);
or U3515 (N_3515,N_3301,N_3296);
or U3516 (N_3516,N_3319,N_3284);
nor U3517 (N_3517,N_3347,N_3330);
or U3518 (N_3518,N_3279,N_3331);
or U3519 (N_3519,N_3297,N_3359);
xor U3520 (N_3520,N_3398,N_3376);
or U3521 (N_3521,N_3222,N_3312);
and U3522 (N_3522,N_3285,N_3249);
or U3523 (N_3523,N_3370,N_3219);
and U3524 (N_3524,N_3230,N_3250);
or U3525 (N_3525,N_3386,N_3262);
nor U3526 (N_3526,N_3347,N_3288);
nand U3527 (N_3527,N_3394,N_3289);
or U3528 (N_3528,N_3328,N_3210);
and U3529 (N_3529,N_3284,N_3234);
nand U3530 (N_3530,N_3377,N_3212);
or U3531 (N_3531,N_3218,N_3385);
or U3532 (N_3532,N_3344,N_3284);
and U3533 (N_3533,N_3290,N_3263);
and U3534 (N_3534,N_3328,N_3204);
and U3535 (N_3535,N_3355,N_3218);
and U3536 (N_3536,N_3340,N_3280);
or U3537 (N_3537,N_3241,N_3282);
and U3538 (N_3538,N_3262,N_3215);
xor U3539 (N_3539,N_3393,N_3222);
and U3540 (N_3540,N_3393,N_3212);
and U3541 (N_3541,N_3399,N_3372);
or U3542 (N_3542,N_3235,N_3232);
and U3543 (N_3543,N_3369,N_3311);
nand U3544 (N_3544,N_3375,N_3336);
or U3545 (N_3545,N_3215,N_3355);
nand U3546 (N_3546,N_3395,N_3295);
or U3547 (N_3547,N_3260,N_3286);
and U3548 (N_3548,N_3257,N_3200);
or U3549 (N_3549,N_3327,N_3376);
xor U3550 (N_3550,N_3312,N_3348);
nor U3551 (N_3551,N_3220,N_3238);
or U3552 (N_3552,N_3347,N_3244);
or U3553 (N_3553,N_3384,N_3232);
or U3554 (N_3554,N_3308,N_3234);
nor U3555 (N_3555,N_3307,N_3203);
or U3556 (N_3556,N_3253,N_3340);
or U3557 (N_3557,N_3301,N_3266);
nand U3558 (N_3558,N_3234,N_3348);
nand U3559 (N_3559,N_3385,N_3237);
nor U3560 (N_3560,N_3231,N_3304);
nand U3561 (N_3561,N_3331,N_3251);
or U3562 (N_3562,N_3210,N_3214);
nor U3563 (N_3563,N_3260,N_3298);
nor U3564 (N_3564,N_3337,N_3290);
or U3565 (N_3565,N_3203,N_3265);
nand U3566 (N_3566,N_3271,N_3388);
xnor U3567 (N_3567,N_3235,N_3213);
nor U3568 (N_3568,N_3294,N_3297);
and U3569 (N_3569,N_3276,N_3296);
nor U3570 (N_3570,N_3256,N_3339);
nand U3571 (N_3571,N_3214,N_3296);
and U3572 (N_3572,N_3393,N_3256);
xor U3573 (N_3573,N_3260,N_3398);
nor U3574 (N_3574,N_3266,N_3399);
and U3575 (N_3575,N_3214,N_3258);
nor U3576 (N_3576,N_3319,N_3356);
or U3577 (N_3577,N_3382,N_3200);
or U3578 (N_3578,N_3256,N_3262);
and U3579 (N_3579,N_3221,N_3369);
and U3580 (N_3580,N_3226,N_3298);
nor U3581 (N_3581,N_3311,N_3266);
nand U3582 (N_3582,N_3372,N_3394);
nand U3583 (N_3583,N_3384,N_3262);
nand U3584 (N_3584,N_3220,N_3228);
xor U3585 (N_3585,N_3389,N_3296);
xnor U3586 (N_3586,N_3262,N_3246);
nor U3587 (N_3587,N_3367,N_3330);
xor U3588 (N_3588,N_3260,N_3346);
and U3589 (N_3589,N_3234,N_3298);
nand U3590 (N_3590,N_3312,N_3292);
and U3591 (N_3591,N_3394,N_3253);
and U3592 (N_3592,N_3347,N_3379);
and U3593 (N_3593,N_3298,N_3209);
nand U3594 (N_3594,N_3299,N_3285);
and U3595 (N_3595,N_3243,N_3386);
or U3596 (N_3596,N_3200,N_3227);
or U3597 (N_3597,N_3298,N_3348);
nand U3598 (N_3598,N_3299,N_3292);
and U3599 (N_3599,N_3396,N_3310);
nand U3600 (N_3600,N_3547,N_3450);
and U3601 (N_3601,N_3409,N_3591);
or U3602 (N_3602,N_3536,N_3468);
or U3603 (N_3603,N_3554,N_3436);
nor U3604 (N_3604,N_3434,N_3574);
or U3605 (N_3605,N_3576,N_3597);
nand U3606 (N_3606,N_3529,N_3505);
nor U3607 (N_3607,N_3420,N_3590);
nor U3608 (N_3608,N_3526,N_3470);
nor U3609 (N_3609,N_3485,N_3501);
and U3610 (N_3610,N_3568,N_3534);
nand U3611 (N_3611,N_3564,N_3511);
xor U3612 (N_3612,N_3431,N_3588);
nor U3613 (N_3613,N_3415,N_3522);
and U3614 (N_3614,N_3419,N_3479);
nand U3615 (N_3615,N_3455,N_3477);
or U3616 (N_3616,N_3571,N_3425);
nor U3617 (N_3617,N_3586,N_3592);
xor U3618 (N_3618,N_3475,N_3558);
nand U3619 (N_3619,N_3553,N_3555);
and U3620 (N_3620,N_3512,N_3570);
nor U3621 (N_3621,N_3427,N_3565);
nand U3622 (N_3622,N_3444,N_3423);
nor U3623 (N_3623,N_3500,N_3561);
xor U3624 (N_3624,N_3451,N_3441);
nand U3625 (N_3625,N_3412,N_3486);
or U3626 (N_3626,N_3416,N_3566);
nand U3627 (N_3627,N_3429,N_3438);
nand U3628 (N_3628,N_3514,N_3482);
and U3629 (N_3629,N_3594,N_3580);
nand U3630 (N_3630,N_3499,N_3532);
and U3631 (N_3631,N_3466,N_3593);
and U3632 (N_3632,N_3445,N_3569);
nor U3633 (N_3633,N_3460,N_3575);
and U3634 (N_3634,N_3405,N_3469);
or U3635 (N_3635,N_3464,N_3497);
or U3636 (N_3636,N_3521,N_3516);
or U3637 (N_3637,N_3454,N_3480);
or U3638 (N_3638,N_3559,N_3573);
or U3639 (N_3639,N_3404,N_3546);
or U3640 (N_3640,N_3463,N_3458);
xor U3641 (N_3641,N_3528,N_3540);
nor U3642 (N_3642,N_3489,N_3513);
xor U3643 (N_3643,N_3467,N_3471);
and U3644 (N_3644,N_3448,N_3401);
nand U3645 (N_3645,N_3520,N_3579);
and U3646 (N_3646,N_3457,N_3437);
and U3647 (N_3647,N_3421,N_3541);
nand U3648 (N_3648,N_3407,N_3446);
nand U3649 (N_3649,N_3556,N_3449);
and U3650 (N_3650,N_3430,N_3495);
nand U3651 (N_3651,N_3508,N_3461);
nand U3652 (N_3652,N_3402,N_3465);
nor U3653 (N_3653,N_3518,N_3414);
xor U3654 (N_3654,N_3583,N_3542);
and U3655 (N_3655,N_3453,N_3435);
and U3656 (N_3656,N_3572,N_3488);
nand U3657 (N_3657,N_3426,N_3549);
or U3658 (N_3658,N_3452,N_3599);
nor U3659 (N_3659,N_3494,N_3524);
and U3660 (N_3660,N_3490,N_3525);
nor U3661 (N_3661,N_3424,N_3584);
nand U3662 (N_3662,N_3413,N_3531);
xnor U3663 (N_3663,N_3504,N_3492);
nor U3664 (N_3664,N_3535,N_3509);
xor U3665 (N_3665,N_3496,N_3507);
and U3666 (N_3666,N_3483,N_3519);
nor U3667 (N_3667,N_3474,N_3523);
and U3668 (N_3668,N_3582,N_3447);
or U3669 (N_3669,N_3567,N_3563);
nand U3670 (N_3670,N_3598,N_3442);
nor U3671 (N_3671,N_3577,N_3510);
or U3672 (N_3672,N_3403,N_3585);
or U3673 (N_3673,N_3506,N_3550);
nor U3674 (N_3674,N_3543,N_3472);
or U3675 (N_3675,N_3443,N_3493);
nand U3676 (N_3676,N_3551,N_3481);
or U3677 (N_3677,N_3462,N_3400);
or U3678 (N_3678,N_3596,N_3406);
nor U3679 (N_3679,N_3498,N_3491);
xor U3680 (N_3680,N_3478,N_3545);
or U3681 (N_3681,N_3581,N_3539);
or U3682 (N_3682,N_3502,N_3537);
or U3683 (N_3683,N_3418,N_3432);
and U3684 (N_3684,N_3517,N_3503);
and U3685 (N_3685,N_3440,N_3557);
nor U3686 (N_3686,N_3562,N_3589);
nor U3687 (N_3687,N_3422,N_3408);
and U3688 (N_3688,N_3433,N_3439);
nand U3689 (N_3689,N_3533,N_3484);
xor U3690 (N_3690,N_3487,N_3459);
nand U3691 (N_3691,N_3456,N_3411);
nor U3692 (N_3692,N_3530,N_3548);
or U3693 (N_3693,N_3515,N_3544);
and U3694 (N_3694,N_3428,N_3552);
nand U3695 (N_3695,N_3476,N_3417);
and U3696 (N_3696,N_3560,N_3538);
or U3697 (N_3697,N_3595,N_3587);
and U3698 (N_3698,N_3578,N_3473);
and U3699 (N_3699,N_3410,N_3527);
and U3700 (N_3700,N_3527,N_3540);
nand U3701 (N_3701,N_3566,N_3595);
nor U3702 (N_3702,N_3531,N_3434);
and U3703 (N_3703,N_3531,N_3573);
xnor U3704 (N_3704,N_3456,N_3407);
and U3705 (N_3705,N_3571,N_3567);
nor U3706 (N_3706,N_3457,N_3431);
and U3707 (N_3707,N_3504,N_3584);
xnor U3708 (N_3708,N_3443,N_3594);
nor U3709 (N_3709,N_3491,N_3511);
nand U3710 (N_3710,N_3581,N_3559);
nor U3711 (N_3711,N_3582,N_3504);
and U3712 (N_3712,N_3410,N_3544);
and U3713 (N_3713,N_3568,N_3439);
nand U3714 (N_3714,N_3458,N_3405);
nand U3715 (N_3715,N_3499,N_3486);
nor U3716 (N_3716,N_3494,N_3527);
nor U3717 (N_3717,N_3557,N_3598);
nand U3718 (N_3718,N_3501,N_3537);
xor U3719 (N_3719,N_3503,N_3479);
and U3720 (N_3720,N_3476,N_3594);
or U3721 (N_3721,N_3470,N_3412);
xnor U3722 (N_3722,N_3570,N_3579);
nand U3723 (N_3723,N_3585,N_3474);
nor U3724 (N_3724,N_3459,N_3494);
nor U3725 (N_3725,N_3586,N_3596);
nand U3726 (N_3726,N_3546,N_3459);
nor U3727 (N_3727,N_3581,N_3547);
and U3728 (N_3728,N_3488,N_3537);
nand U3729 (N_3729,N_3482,N_3577);
and U3730 (N_3730,N_3520,N_3463);
and U3731 (N_3731,N_3530,N_3460);
nand U3732 (N_3732,N_3559,N_3411);
and U3733 (N_3733,N_3431,N_3427);
xor U3734 (N_3734,N_3568,N_3458);
or U3735 (N_3735,N_3429,N_3557);
nor U3736 (N_3736,N_3571,N_3599);
nand U3737 (N_3737,N_3495,N_3591);
or U3738 (N_3738,N_3534,N_3560);
nand U3739 (N_3739,N_3430,N_3579);
nor U3740 (N_3740,N_3484,N_3464);
and U3741 (N_3741,N_3500,N_3598);
nand U3742 (N_3742,N_3470,N_3414);
nor U3743 (N_3743,N_3517,N_3541);
nor U3744 (N_3744,N_3597,N_3589);
nand U3745 (N_3745,N_3514,N_3502);
nor U3746 (N_3746,N_3550,N_3493);
nor U3747 (N_3747,N_3532,N_3405);
or U3748 (N_3748,N_3542,N_3520);
and U3749 (N_3749,N_3566,N_3518);
nand U3750 (N_3750,N_3441,N_3458);
or U3751 (N_3751,N_3477,N_3559);
and U3752 (N_3752,N_3417,N_3495);
nor U3753 (N_3753,N_3453,N_3470);
xnor U3754 (N_3754,N_3533,N_3437);
nand U3755 (N_3755,N_3536,N_3451);
and U3756 (N_3756,N_3446,N_3469);
or U3757 (N_3757,N_3465,N_3460);
and U3758 (N_3758,N_3598,N_3514);
nand U3759 (N_3759,N_3589,N_3507);
xnor U3760 (N_3760,N_3550,N_3401);
xnor U3761 (N_3761,N_3441,N_3523);
and U3762 (N_3762,N_3588,N_3558);
and U3763 (N_3763,N_3401,N_3506);
and U3764 (N_3764,N_3529,N_3487);
or U3765 (N_3765,N_3553,N_3490);
nand U3766 (N_3766,N_3404,N_3518);
nand U3767 (N_3767,N_3564,N_3501);
nand U3768 (N_3768,N_3415,N_3549);
and U3769 (N_3769,N_3570,N_3456);
nand U3770 (N_3770,N_3486,N_3514);
and U3771 (N_3771,N_3433,N_3518);
and U3772 (N_3772,N_3597,N_3418);
nand U3773 (N_3773,N_3456,N_3553);
nand U3774 (N_3774,N_3530,N_3537);
xor U3775 (N_3775,N_3465,N_3483);
or U3776 (N_3776,N_3568,N_3517);
nor U3777 (N_3777,N_3571,N_3538);
nand U3778 (N_3778,N_3404,N_3461);
and U3779 (N_3779,N_3572,N_3460);
nor U3780 (N_3780,N_3437,N_3534);
and U3781 (N_3781,N_3566,N_3471);
nand U3782 (N_3782,N_3570,N_3481);
xnor U3783 (N_3783,N_3584,N_3528);
or U3784 (N_3784,N_3582,N_3567);
or U3785 (N_3785,N_3489,N_3480);
or U3786 (N_3786,N_3536,N_3467);
or U3787 (N_3787,N_3413,N_3465);
xor U3788 (N_3788,N_3437,N_3585);
and U3789 (N_3789,N_3592,N_3580);
and U3790 (N_3790,N_3486,N_3495);
and U3791 (N_3791,N_3538,N_3594);
or U3792 (N_3792,N_3502,N_3584);
nand U3793 (N_3793,N_3417,N_3431);
and U3794 (N_3794,N_3589,N_3538);
nor U3795 (N_3795,N_3570,N_3404);
or U3796 (N_3796,N_3473,N_3482);
and U3797 (N_3797,N_3427,N_3493);
nor U3798 (N_3798,N_3431,N_3470);
nand U3799 (N_3799,N_3508,N_3468);
and U3800 (N_3800,N_3773,N_3713);
and U3801 (N_3801,N_3780,N_3601);
nand U3802 (N_3802,N_3705,N_3633);
nor U3803 (N_3803,N_3638,N_3767);
nand U3804 (N_3804,N_3600,N_3646);
nor U3805 (N_3805,N_3726,N_3753);
nand U3806 (N_3806,N_3655,N_3623);
nand U3807 (N_3807,N_3759,N_3724);
or U3808 (N_3808,N_3630,N_3793);
nand U3809 (N_3809,N_3653,N_3708);
nand U3810 (N_3810,N_3668,N_3722);
nand U3811 (N_3811,N_3607,N_3747);
or U3812 (N_3812,N_3671,N_3789);
or U3813 (N_3813,N_3661,N_3717);
nand U3814 (N_3814,N_3704,N_3718);
xor U3815 (N_3815,N_3613,N_3691);
nor U3816 (N_3816,N_3687,N_3775);
nor U3817 (N_3817,N_3751,N_3795);
nor U3818 (N_3818,N_3690,N_3725);
or U3819 (N_3819,N_3602,N_3647);
or U3820 (N_3820,N_3664,N_3683);
xor U3821 (N_3821,N_3714,N_3673);
or U3822 (N_3822,N_3741,N_3783);
and U3823 (N_3823,N_3766,N_3701);
nor U3824 (N_3824,N_3744,N_3743);
or U3825 (N_3825,N_3626,N_3731);
nor U3826 (N_3826,N_3720,N_3635);
nor U3827 (N_3827,N_3659,N_3707);
nand U3828 (N_3828,N_3643,N_3697);
xnor U3829 (N_3829,N_3644,N_3778);
or U3830 (N_3830,N_3700,N_3636);
and U3831 (N_3831,N_3648,N_3791);
or U3832 (N_3832,N_3693,N_3641);
xor U3833 (N_3833,N_3663,N_3674);
nand U3834 (N_3834,N_3675,N_3618);
or U3835 (N_3835,N_3728,N_3712);
nand U3836 (N_3836,N_3672,N_3763);
or U3837 (N_3837,N_3740,N_3651);
xor U3838 (N_3838,N_3606,N_3739);
nand U3839 (N_3839,N_3614,N_3629);
or U3840 (N_3840,N_3696,N_3684);
nor U3841 (N_3841,N_3620,N_3616);
nor U3842 (N_3842,N_3694,N_3709);
nor U3843 (N_3843,N_3757,N_3615);
nand U3844 (N_3844,N_3733,N_3730);
or U3845 (N_3845,N_3667,N_3645);
and U3846 (N_3846,N_3605,N_3665);
xnor U3847 (N_3847,N_3760,N_3721);
or U3848 (N_3848,N_3699,N_3686);
and U3849 (N_3849,N_3662,N_3734);
and U3850 (N_3850,N_3627,N_3609);
or U3851 (N_3851,N_3611,N_3772);
nor U3852 (N_3852,N_3634,N_3603);
or U3853 (N_3853,N_3732,N_3770);
nor U3854 (N_3854,N_3755,N_3764);
nor U3855 (N_3855,N_3631,N_3790);
and U3856 (N_3856,N_3695,N_3677);
nand U3857 (N_3857,N_3797,N_3666);
or U3858 (N_3858,N_3688,N_3769);
nand U3859 (N_3859,N_3658,N_3782);
and U3860 (N_3860,N_3679,N_3754);
nor U3861 (N_3861,N_3727,N_3737);
nor U3862 (N_3862,N_3762,N_3774);
and U3863 (N_3863,N_3779,N_3756);
or U3864 (N_3864,N_3637,N_3738);
nor U3865 (N_3865,N_3608,N_3624);
nor U3866 (N_3866,N_3736,N_3792);
nand U3867 (N_3867,N_3715,N_3660);
nor U3868 (N_3868,N_3702,N_3621);
and U3869 (N_3869,N_3716,N_3656);
and U3870 (N_3870,N_3610,N_3604);
nand U3871 (N_3871,N_3681,N_3682);
and U3872 (N_3872,N_3676,N_3796);
and U3873 (N_3873,N_3669,N_3640);
and U3874 (N_3874,N_3776,N_3703);
or U3875 (N_3875,N_3617,N_3649);
nor U3876 (N_3876,N_3729,N_3784);
nor U3877 (N_3877,N_3632,N_3750);
xor U3878 (N_3878,N_3788,N_3761);
and U3879 (N_3879,N_3711,N_3685);
nand U3880 (N_3880,N_3748,N_3698);
or U3881 (N_3881,N_3678,N_3628);
nand U3882 (N_3882,N_3771,N_3619);
and U3883 (N_3883,N_3787,N_3799);
nand U3884 (N_3884,N_3652,N_3777);
and U3885 (N_3885,N_3719,N_3785);
nand U3886 (N_3886,N_3752,N_3765);
and U3887 (N_3887,N_3735,N_3706);
nand U3888 (N_3888,N_3798,N_3746);
nor U3889 (N_3889,N_3749,N_3723);
nand U3890 (N_3890,N_3742,N_3639);
or U3891 (N_3891,N_3670,N_3622);
nand U3892 (N_3892,N_3680,N_3786);
nor U3893 (N_3893,N_3625,N_3781);
or U3894 (N_3894,N_3758,N_3657);
nor U3895 (N_3895,N_3710,N_3642);
or U3896 (N_3896,N_3650,N_3612);
or U3897 (N_3897,N_3794,N_3692);
nand U3898 (N_3898,N_3768,N_3654);
nor U3899 (N_3899,N_3745,N_3689);
nand U3900 (N_3900,N_3611,N_3683);
nor U3901 (N_3901,N_3711,N_3744);
or U3902 (N_3902,N_3752,N_3619);
and U3903 (N_3903,N_3779,N_3614);
xnor U3904 (N_3904,N_3738,N_3665);
or U3905 (N_3905,N_3636,N_3618);
nand U3906 (N_3906,N_3600,N_3711);
or U3907 (N_3907,N_3669,N_3762);
or U3908 (N_3908,N_3620,N_3724);
nor U3909 (N_3909,N_3738,N_3640);
nand U3910 (N_3910,N_3730,N_3783);
and U3911 (N_3911,N_3606,N_3782);
nor U3912 (N_3912,N_3739,N_3744);
nand U3913 (N_3913,N_3672,N_3610);
and U3914 (N_3914,N_3602,N_3777);
nand U3915 (N_3915,N_3678,N_3640);
and U3916 (N_3916,N_3747,N_3743);
and U3917 (N_3917,N_3645,N_3604);
and U3918 (N_3918,N_3721,N_3692);
nor U3919 (N_3919,N_3747,N_3706);
or U3920 (N_3920,N_3748,N_3710);
nor U3921 (N_3921,N_3685,N_3663);
or U3922 (N_3922,N_3601,N_3656);
and U3923 (N_3923,N_3672,N_3773);
or U3924 (N_3924,N_3660,N_3652);
or U3925 (N_3925,N_3654,N_3739);
and U3926 (N_3926,N_3646,N_3643);
or U3927 (N_3927,N_3673,N_3795);
and U3928 (N_3928,N_3647,N_3694);
nand U3929 (N_3929,N_3658,N_3704);
and U3930 (N_3930,N_3697,N_3683);
and U3931 (N_3931,N_3781,N_3747);
and U3932 (N_3932,N_3727,N_3665);
xor U3933 (N_3933,N_3709,N_3730);
nor U3934 (N_3934,N_3692,N_3704);
nor U3935 (N_3935,N_3727,N_3641);
nor U3936 (N_3936,N_3780,N_3774);
nand U3937 (N_3937,N_3671,N_3759);
or U3938 (N_3938,N_3609,N_3653);
nand U3939 (N_3939,N_3619,N_3721);
nor U3940 (N_3940,N_3674,N_3741);
xnor U3941 (N_3941,N_3671,N_3765);
and U3942 (N_3942,N_3716,N_3765);
or U3943 (N_3943,N_3723,N_3744);
and U3944 (N_3944,N_3748,N_3785);
or U3945 (N_3945,N_3773,N_3768);
or U3946 (N_3946,N_3648,N_3675);
and U3947 (N_3947,N_3636,N_3721);
xor U3948 (N_3948,N_3703,N_3634);
nor U3949 (N_3949,N_3621,N_3602);
and U3950 (N_3950,N_3776,N_3799);
and U3951 (N_3951,N_3698,N_3771);
nand U3952 (N_3952,N_3664,N_3611);
or U3953 (N_3953,N_3798,N_3731);
or U3954 (N_3954,N_3662,N_3616);
nor U3955 (N_3955,N_3786,N_3678);
and U3956 (N_3956,N_3676,N_3782);
and U3957 (N_3957,N_3624,N_3770);
nand U3958 (N_3958,N_3604,N_3629);
nand U3959 (N_3959,N_3652,N_3731);
and U3960 (N_3960,N_3796,N_3702);
or U3961 (N_3961,N_3777,N_3747);
or U3962 (N_3962,N_3761,N_3755);
and U3963 (N_3963,N_3730,N_3779);
nor U3964 (N_3964,N_3750,N_3652);
xnor U3965 (N_3965,N_3787,N_3762);
and U3966 (N_3966,N_3699,N_3659);
or U3967 (N_3967,N_3731,N_3673);
or U3968 (N_3968,N_3763,N_3621);
or U3969 (N_3969,N_3621,N_3752);
and U3970 (N_3970,N_3600,N_3747);
xnor U3971 (N_3971,N_3770,N_3695);
nor U3972 (N_3972,N_3786,N_3739);
nand U3973 (N_3973,N_3601,N_3614);
and U3974 (N_3974,N_3671,N_3626);
nor U3975 (N_3975,N_3729,N_3624);
xor U3976 (N_3976,N_3652,N_3656);
or U3977 (N_3977,N_3626,N_3793);
and U3978 (N_3978,N_3668,N_3720);
nor U3979 (N_3979,N_3646,N_3798);
nand U3980 (N_3980,N_3690,N_3669);
xor U3981 (N_3981,N_3741,N_3790);
or U3982 (N_3982,N_3680,N_3698);
xor U3983 (N_3983,N_3743,N_3726);
or U3984 (N_3984,N_3702,N_3635);
and U3985 (N_3985,N_3789,N_3621);
xor U3986 (N_3986,N_3687,N_3737);
and U3987 (N_3987,N_3642,N_3711);
or U3988 (N_3988,N_3713,N_3731);
or U3989 (N_3989,N_3785,N_3794);
and U3990 (N_3990,N_3638,N_3664);
nor U3991 (N_3991,N_3703,N_3700);
xor U3992 (N_3992,N_3718,N_3683);
nor U3993 (N_3993,N_3793,N_3687);
and U3994 (N_3994,N_3676,N_3754);
or U3995 (N_3995,N_3623,N_3753);
nor U3996 (N_3996,N_3703,N_3677);
and U3997 (N_3997,N_3767,N_3646);
nand U3998 (N_3998,N_3601,N_3615);
nor U3999 (N_3999,N_3669,N_3786);
and U4000 (N_4000,N_3812,N_3912);
nand U4001 (N_4001,N_3897,N_3985);
or U4002 (N_4002,N_3884,N_3929);
nor U4003 (N_4003,N_3847,N_3854);
nand U4004 (N_4004,N_3963,N_3954);
xor U4005 (N_4005,N_3953,N_3896);
nor U4006 (N_4006,N_3969,N_3907);
xnor U4007 (N_4007,N_3801,N_3885);
and U4008 (N_4008,N_3879,N_3876);
nor U4009 (N_4009,N_3807,N_3823);
or U4010 (N_4010,N_3966,N_3889);
nand U4011 (N_4011,N_3899,N_3970);
nor U4012 (N_4012,N_3974,N_3883);
and U4013 (N_4013,N_3851,N_3874);
and U4014 (N_4014,N_3856,N_3916);
nand U4015 (N_4015,N_3837,N_3928);
and U4016 (N_4016,N_3943,N_3880);
nor U4017 (N_4017,N_3902,N_3861);
nor U4018 (N_4018,N_3841,N_3961);
or U4019 (N_4019,N_3891,N_3852);
xor U4020 (N_4020,N_3833,N_3934);
or U4021 (N_4021,N_3829,N_3815);
or U4022 (N_4022,N_3831,N_3982);
nor U4023 (N_4023,N_3992,N_3957);
or U4024 (N_4024,N_3976,N_3855);
nand U4025 (N_4025,N_3864,N_3910);
nor U4026 (N_4026,N_3956,N_3993);
nor U4027 (N_4027,N_3981,N_3830);
or U4028 (N_4028,N_3933,N_3828);
nor U4029 (N_4029,N_3816,N_3932);
or U4030 (N_4030,N_3806,N_3835);
and U4031 (N_4031,N_3834,N_3922);
xnor U4032 (N_4032,N_3820,N_3848);
nor U4033 (N_4033,N_3809,N_3908);
and U4034 (N_4034,N_3893,N_3983);
and U4035 (N_4035,N_3898,N_3877);
nor U4036 (N_4036,N_3827,N_3814);
nor U4037 (N_4037,N_3886,N_3904);
and U4038 (N_4038,N_3824,N_3973);
nor U4039 (N_4039,N_3931,N_3914);
and U4040 (N_4040,N_3839,N_3958);
or U4041 (N_4041,N_3924,N_3865);
nand U4042 (N_4042,N_3842,N_3903);
or U4043 (N_4043,N_3918,N_3972);
or U4044 (N_4044,N_3964,N_3800);
and U4045 (N_4045,N_3936,N_3959);
nand U4046 (N_4046,N_3890,N_3810);
or U4047 (N_4047,N_3948,N_3952);
nand U4048 (N_4048,N_3975,N_3962);
or U4049 (N_4049,N_3906,N_3887);
nor U4050 (N_4050,N_3968,N_3860);
nor U4051 (N_4051,N_3870,N_3926);
xnor U4052 (N_4052,N_3875,N_3939);
or U4053 (N_4053,N_3868,N_3905);
xor U4054 (N_4054,N_3979,N_3871);
nand U4055 (N_4055,N_3917,N_3878);
or U4056 (N_4056,N_3930,N_3987);
and U4057 (N_4057,N_3978,N_3941);
nand U4058 (N_4058,N_3997,N_3832);
or U4059 (N_4059,N_3846,N_3980);
xor U4060 (N_4060,N_3927,N_3988);
nand U4061 (N_4061,N_3911,N_3951);
xnor U4062 (N_4062,N_3935,N_3817);
nand U4063 (N_4063,N_3950,N_3862);
or U4064 (N_4064,N_3999,N_3892);
nand U4065 (N_4065,N_3849,N_3996);
nand U4066 (N_4066,N_3894,N_3913);
nor U4067 (N_4067,N_3803,N_3822);
or U4068 (N_4068,N_3804,N_3945);
nor U4069 (N_4069,N_3826,N_3863);
nor U4070 (N_4070,N_3802,N_3881);
xor U4071 (N_4071,N_3949,N_3967);
and U4072 (N_4072,N_3990,N_3836);
nand U4073 (N_4073,N_3811,N_3971);
and U4074 (N_4074,N_3938,N_3984);
and U4075 (N_4075,N_3920,N_3844);
xnor U4076 (N_4076,N_3901,N_3843);
nor U4077 (N_4077,N_3977,N_3859);
nand U4078 (N_4078,N_3915,N_3940);
nor U4079 (N_4079,N_3947,N_3838);
nor U4080 (N_4080,N_3946,N_3873);
nor U4081 (N_4081,N_3869,N_3995);
xnor U4082 (N_4082,N_3986,N_3989);
and U4083 (N_4083,N_3867,N_3937);
or U4084 (N_4084,N_3813,N_3925);
xnor U4085 (N_4085,N_3872,N_3994);
nor U4086 (N_4086,N_3942,N_3923);
nand U4087 (N_4087,N_3955,N_3882);
and U4088 (N_4088,N_3909,N_3866);
xor U4089 (N_4089,N_3991,N_3805);
nand U4090 (N_4090,N_3819,N_3850);
nand U4091 (N_4091,N_3944,N_3960);
nand U4092 (N_4092,N_3895,N_3821);
nor U4093 (N_4093,N_3921,N_3857);
xnor U4094 (N_4094,N_3900,N_3858);
nand U4095 (N_4095,N_3825,N_3919);
nand U4096 (N_4096,N_3965,N_3853);
nor U4097 (N_4097,N_3998,N_3845);
nor U4098 (N_4098,N_3818,N_3808);
or U4099 (N_4099,N_3888,N_3840);
nand U4100 (N_4100,N_3877,N_3968);
nor U4101 (N_4101,N_3956,N_3981);
and U4102 (N_4102,N_3822,N_3924);
and U4103 (N_4103,N_3835,N_3952);
nand U4104 (N_4104,N_3996,N_3885);
and U4105 (N_4105,N_3992,N_3970);
nor U4106 (N_4106,N_3954,N_3858);
nand U4107 (N_4107,N_3917,N_3890);
nor U4108 (N_4108,N_3837,N_3817);
nand U4109 (N_4109,N_3845,N_3887);
nand U4110 (N_4110,N_3807,N_3969);
or U4111 (N_4111,N_3989,N_3853);
and U4112 (N_4112,N_3916,N_3901);
nand U4113 (N_4113,N_3869,N_3899);
and U4114 (N_4114,N_3903,N_3889);
nor U4115 (N_4115,N_3993,N_3922);
nand U4116 (N_4116,N_3825,N_3856);
xor U4117 (N_4117,N_3897,N_3836);
and U4118 (N_4118,N_3991,N_3998);
or U4119 (N_4119,N_3919,N_3876);
nor U4120 (N_4120,N_3872,N_3823);
nand U4121 (N_4121,N_3996,N_3993);
nor U4122 (N_4122,N_3935,N_3829);
nor U4123 (N_4123,N_3894,N_3855);
or U4124 (N_4124,N_3921,N_3802);
and U4125 (N_4125,N_3932,N_3897);
and U4126 (N_4126,N_3978,N_3859);
nor U4127 (N_4127,N_3846,N_3933);
or U4128 (N_4128,N_3879,N_3828);
nor U4129 (N_4129,N_3921,N_3828);
and U4130 (N_4130,N_3987,N_3982);
and U4131 (N_4131,N_3926,N_3822);
nand U4132 (N_4132,N_3997,N_3906);
xnor U4133 (N_4133,N_3835,N_3931);
xor U4134 (N_4134,N_3933,N_3927);
xnor U4135 (N_4135,N_3809,N_3838);
nor U4136 (N_4136,N_3868,N_3912);
or U4137 (N_4137,N_3946,N_3947);
or U4138 (N_4138,N_3867,N_3915);
and U4139 (N_4139,N_3833,N_3815);
and U4140 (N_4140,N_3845,N_3830);
or U4141 (N_4141,N_3921,N_3948);
or U4142 (N_4142,N_3948,N_3859);
and U4143 (N_4143,N_3886,N_3965);
nor U4144 (N_4144,N_3887,N_3969);
or U4145 (N_4145,N_3947,N_3989);
and U4146 (N_4146,N_3980,N_3871);
nor U4147 (N_4147,N_3936,N_3878);
nand U4148 (N_4148,N_3853,N_3970);
and U4149 (N_4149,N_3896,N_3911);
and U4150 (N_4150,N_3850,N_3858);
and U4151 (N_4151,N_3871,N_3848);
or U4152 (N_4152,N_3882,N_3959);
and U4153 (N_4153,N_3942,N_3986);
nor U4154 (N_4154,N_3917,N_3992);
and U4155 (N_4155,N_3985,N_3853);
or U4156 (N_4156,N_3922,N_3830);
and U4157 (N_4157,N_3942,N_3909);
nor U4158 (N_4158,N_3958,N_3806);
or U4159 (N_4159,N_3849,N_3882);
or U4160 (N_4160,N_3983,N_3956);
or U4161 (N_4161,N_3835,N_3991);
and U4162 (N_4162,N_3851,N_3991);
and U4163 (N_4163,N_3946,N_3842);
or U4164 (N_4164,N_3809,N_3892);
nor U4165 (N_4165,N_3945,N_3801);
nor U4166 (N_4166,N_3850,N_3966);
nand U4167 (N_4167,N_3960,N_3986);
nand U4168 (N_4168,N_3836,N_3874);
or U4169 (N_4169,N_3908,N_3962);
nand U4170 (N_4170,N_3992,N_3800);
nor U4171 (N_4171,N_3941,N_3897);
or U4172 (N_4172,N_3958,N_3902);
nand U4173 (N_4173,N_3971,N_3859);
or U4174 (N_4174,N_3881,N_3968);
nand U4175 (N_4175,N_3950,N_3885);
xnor U4176 (N_4176,N_3803,N_3961);
nor U4177 (N_4177,N_3965,N_3988);
nand U4178 (N_4178,N_3932,N_3869);
and U4179 (N_4179,N_3892,N_3915);
xnor U4180 (N_4180,N_3975,N_3997);
or U4181 (N_4181,N_3823,N_3802);
or U4182 (N_4182,N_3920,N_3864);
and U4183 (N_4183,N_3941,N_3985);
xor U4184 (N_4184,N_3907,N_3852);
or U4185 (N_4185,N_3981,N_3942);
nor U4186 (N_4186,N_3901,N_3847);
nand U4187 (N_4187,N_3814,N_3802);
nand U4188 (N_4188,N_3949,N_3925);
or U4189 (N_4189,N_3946,N_3859);
and U4190 (N_4190,N_3843,N_3885);
or U4191 (N_4191,N_3868,N_3858);
and U4192 (N_4192,N_3871,N_3978);
nand U4193 (N_4193,N_3817,N_3979);
and U4194 (N_4194,N_3872,N_3827);
nor U4195 (N_4195,N_3895,N_3912);
nor U4196 (N_4196,N_3876,N_3970);
nor U4197 (N_4197,N_3884,N_3895);
nand U4198 (N_4198,N_3913,N_3926);
nor U4199 (N_4199,N_3875,N_3897);
and U4200 (N_4200,N_4172,N_4132);
or U4201 (N_4201,N_4013,N_4144);
nand U4202 (N_4202,N_4021,N_4161);
or U4203 (N_4203,N_4163,N_4155);
nand U4204 (N_4204,N_4184,N_4199);
or U4205 (N_4205,N_4188,N_4056);
nand U4206 (N_4206,N_4140,N_4129);
and U4207 (N_4207,N_4041,N_4150);
or U4208 (N_4208,N_4093,N_4146);
and U4209 (N_4209,N_4009,N_4044);
nor U4210 (N_4210,N_4076,N_4198);
nand U4211 (N_4211,N_4101,N_4166);
nand U4212 (N_4212,N_4114,N_4112);
xor U4213 (N_4213,N_4080,N_4136);
or U4214 (N_4214,N_4089,N_4177);
or U4215 (N_4215,N_4157,N_4168);
nor U4216 (N_4216,N_4178,N_4067);
nor U4217 (N_4217,N_4014,N_4045);
nand U4218 (N_4218,N_4191,N_4180);
nor U4219 (N_4219,N_4171,N_4143);
or U4220 (N_4220,N_4027,N_4109);
nand U4221 (N_4221,N_4190,N_4043);
or U4222 (N_4222,N_4128,N_4094);
or U4223 (N_4223,N_4092,N_4105);
nor U4224 (N_4224,N_4147,N_4182);
and U4225 (N_4225,N_4079,N_4074);
nand U4226 (N_4226,N_4110,N_4126);
and U4227 (N_4227,N_4040,N_4106);
nor U4228 (N_4228,N_4058,N_4137);
and U4229 (N_4229,N_4010,N_4141);
or U4230 (N_4230,N_4158,N_4059);
nor U4231 (N_4231,N_4169,N_4176);
nor U4232 (N_4232,N_4090,N_4037);
nor U4233 (N_4233,N_4064,N_4164);
and U4234 (N_4234,N_4052,N_4096);
xnor U4235 (N_4235,N_4099,N_4173);
nand U4236 (N_4236,N_4115,N_4193);
nand U4237 (N_4237,N_4032,N_4004);
and U4238 (N_4238,N_4015,N_4098);
and U4239 (N_4239,N_4035,N_4102);
or U4240 (N_4240,N_4117,N_4125);
nand U4241 (N_4241,N_4165,N_4138);
and U4242 (N_4242,N_4148,N_4159);
nand U4243 (N_4243,N_4030,N_4025);
nand U4244 (N_4244,N_4063,N_4108);
or U4245 (N_4245,N_4123,N_4072);
nor U4246 (N_4246,N_4154,N_4012);
or U4247 (N_4247,N_4195,N_4156);
or U4248 (N_4248,N_4005,N_4042);
nand U4249 (N_4249,N_4057,N_4175);
or U4250 (N_4250,N_4019,N_4055);
nor U4251 (N_4251,N_4062,N_4091);
nor U4252 (N_4252,N_4026,N_4111);
or U4253 (N_4253,N_4085,N_4075);
and U4254 (N_4254,N_4185,N_4061);
xnor U4255 (N_4255,N_4120,N_4088);
nor U4256 (N_4256,N_4008,N_4001);
nand U4257 (N_4257,N_4007,N_4186);
and U4258 (N_4258,N_4139,N_4086);
or U4259 (N_4259,N_4068,N_4082);
nand U4260 (N_4260,N_4153,N_4135);
or U4261 (N_4261,N_4073,N_4145);
nor U4262 (N_4262,N_4018,N_4000);
and U4263 (N_4263,N_4071,N_4187);
and U4264 (N_4264,N_4060,N_4031);
nor U4265 (N_4265,N_4049,N_4036);
and U4266 (N_4266,N_4124,N_4084);
and U4267 (N_4267,N_4130,N_4107);
nand U4268 (N_4268,N_4103,N_4083);
nor U4269 (N_4269,N_4160,N_4039);
nand U4270 (N_4270,N_4053,N_4116);
or U4271 (N_4271,N_4192,N_4174);
or U4272 (N_4272,N_4016,N_4077);
or U4273 (N_4273,N_4152,N_4038);
or U4274 (N_4274,N_4194,N_4149);
and U4275 (N_4275,N_4065,N_4162);
or U4276 (N_4276,N_4196,N_4029);
nand U4277 (N_4277,N_4087,N_4011);
and U4278 (N_4278,N_4070,N_4142);
or U4279 (N_4279,N_4151,N_4003);
xnor U4280 (N_4280,N_4017,N_4133);
nand U4281 (N_4281,N_4050,N_4183);
xor U4282 (N_4282,N_4119,N_4069);
and U4283 (N_4283,N_4034,N_4167);
nand U4284 (N_4284,N_4048,N_4113);
nor U4285 (N_4285,N_4118,N_4179);
and U4286 (N_4286,N_4054,N_4020);
and U4287 (N_4287,N_4127,N_4046);
or U4288 (N_4288,N_4066,N_4181);
or U4289 (N_4289,N_4100,N_4097);
nor U4290 (N_4290,N_4047,N_4022);
or U4291 (N_4291,N_4170,N_4197);
nor U4292 (N_4292,N_4095,N_4024);
and U4293 (N_4293,N_4131,N_4104);
xor U4294 (N_4294,N_4121,N_4122);
nand U4295 (N_4295,N_4002,N_4033);
and U4296 (N_4296,N_4078,N_4189);
nand U4297 (N_4297,N_4081,N_4028);
and U4298 (N_4298,N_4023,N_4006);
and U4299 (N_4299,N_4051,N_4134);
nor U4300 (N_4300,N_4167,N_4115);
and U4301 (N_4301,N_4137,N_4099);
or U4302 (N_4302,N_4051,N_4020);
nand U4303 (N_4303,N_4190,N_4104);
nand U4304 (N_4304,N_4198,N_4110);
nor U4305 (N_4305,N_4103,N_4178);
nor U4306 (N_4306,N_4056,N_4052);
nor U4307 (N_4307,N_4029,N_4191);
nand U4308 (N_4308,N_4073,N_4112);
or U4309 (N_4309,N_4023,N_4126);
and U4310 (N_4310,N_4102,N_4045);
or U4311 (N_4311,N_4079,N_4103);
xor U4312 (N_4312,N_4146,N_4152);
and U4313 (N_4313,N_4165,N_4174);
nand U4314 (N_4314,N_4141,N_4113);
and U4315 (N_4315,N_4043,N_4132);
or U4316 (N_4316,N_4013,N_4056);
or U4317 (N_4317,N_4093,N_4057);
nand U4318 (N_4318,N_4038,N_4030);
nand U4319 (N_4319,N_4028,N_4147);
xnor U4320 (N_4320,N_4102,N_4193);
and U4321 (N_4321,N_4095,N_4114);
and U4322 (N_4322,N_4064,N_4066);
and U4323 (N_4323,N_4156,N_4017);
and U4324 (N_4324,N_4165,N_4105);
nand U4325 (N_4325,N_4031,N_4086);
and U4326 (N_4326,N_4042,N_4095);
nand U4327 (N_4327,N_4137,N_4095);
nor U4328 (N_4328,N_4017,N_4114);
or U4329 (N_4329,N_4168,N_4110);
or U4330 (N_4330,N_4145,N_4090);
nor U4331 (N_4331,N_4096,N_4083);
nor U4332 (N_4332,N_4099,N_4022);
nand U4333 (N_4333,N_4179,N_4036);
or U4334 (N_4334,N_4165,N_4163);
nand U4335 (N_4335,N_4012,N_4171);
xnor U4336 (N_4336,N_4097,N_4045);
nor U4337 (N_4337,N_4018,N_4148);
nor U4338 (N_4338,N_4108,N_4127);
or U4339 (N_4339,N_4014,N_4148);
and U4340 (N_4340,N_4197,N_4069);
xnor U4341 (N_4341,N_4138,N_4176);
nor U4342 (N_4342,N_4080,N_4198);
and U4343 (N_4343,N_4039,N_4121);
or U4344 (N_4344,N_4114,N_4158);
nand U4345 (N_4345,N_4126,N_4042);
nor U4346 (N_4346,N_4111,N_4016);
and U4347 (N_4347,N_4151,N_4002);
and U4348 (N_4348,N_4113,N_4063);
nand U4349 (N_4349,N_4020,N_4079);
or U4350 (N_4350,N_4064,N_4073);
and U4351 (N_4351,N_4065,N_4168);
nand U4352 (N_4352,N_4048,N_4085);
xor U4353 (N_4353,N_4165,N_4087);
nand U4354 (N_4354,N_4078,N_4092);
nand U4355 (N_4355,N_4112,N_4138);
and U4356 (N_4356,N_4197,N_4081);
xnor U4357 (N_4357,N_4055,N_4108);
and U4358 (N_4358,N_4110,N_4018);
and U4359 (N_4359,N_4180,N_4181);
xor U4360 (N_4360,N_4147,N_4058);
xnor U4361 (N_4361,N_4154,N_4133);
nor U4362 (N_4362,N_4148,N_4096);
or U4363 (N_4363,N_4113,N_4139);
nand U4364 (N_4364,N_4001,N_4051);
nor U4365 (N_4365,N_4178,N_4044);
and U4366 (N_4366,N_4108,N_4085);
nand U4367 (N_4367,N_4040,N_4091);
nor U4368 (N_4368,N_4043,N_4140);
or U4369 (N_4369,N_4078,N_4193);
nand U4370 (N_4370,N_4021,N_4002);
or U4371 (N_4371,N_4105,N_4160);
or U4372 (N_4372,N_4041,N_4174);
nor U4373 (N_4373,N_4095,N_4183);
or U4374 (N_4374,N_4053,N_4124);
or U4375 (N_4375,N_4157,N_4063);
nor U4376 (N_4376,N_4083,N_4143);
and U4377 (N_4377,N_4090,N_4164);
nand U4378 (N_4378,N_4013,N_4182);
nand U4379 (N_4379,N_4024,N_4142);
nor U4380 (N_4380,N_4189,N_4172);
nand U4381 (N_4381,N_4037,N_4197);
nand U4382 (N_4382,N_4173,N_4152);
nor U4383 (N_4383,N_4185,N_4034);
and U4384 (N_4384,N_4034,N_4088);
and U4385 (N_4385,N_4114,N_4108);
nor U4386 (N_4386,N_4152,N_4001);
nand U4387 (N_4387,N_4180,N_4160);
and U4388 (N_4388,N_4011,N_4100);
and U4389 (N_4389,N_4029,N_4144);
nor U4390 (N_4390,N_4030,N_4026);
or U4391 (N_4391,N_4030,N_4144);
or U4392 (N_4392,N_4126,N_4097);
and U4393 (N_4393,N_4080,N_4121);
nand U4394 (N_4394,N_4066,N_4140);
and U4395 (N_4395,N_4185,N_4030);
nor U4396 (N_4396,N_4184,N_4019);
and U4397 (N_4397,N_4021,N_4194);
and U4398 (N_4398,N_4094,N_4145);
and U4399 (N_4399,N_4041,N_4126);
and U4400 (N_4400,N_4224,N_4273);
and U4401 (N_4401,N_4350,N_4364);
or U4402 (N_4402,N_4369,N_4231);
and U4403 (N_4403,N_4377,N_4287);
or U4404 (N_4404,N_4356,N_4264);
or U4405 (N_4405,N_4204,N_4380);
xnor U4406 (N_4406,N_4324,N_4368);
or U4407 (N_4407,N_4329,N_4366);
and U4408 (N_4408,N_4278,N_4254);
and U4409 (N_4409,N_4298,N_4221);
nand U4410 (N_4410,N_4385,N_4372);
or U4411 (N_4411,N_4265,N_4210);
and U4412 (N_4412,N_4227,N_4341);
nand U4413 (N_4413,N_4344,N_4219);
and U4414 (N_4414,N_4330,N_4226);
and U4415 (N_4415,N_4381,N_4216);
and U4416 (N_4416,N_4253,N_4268);
nand U4417 (N_4417,N_4388,N_4367);
or U4418 (N_4418,N_4242,N_4211);
xnor U4419 (N_4419,N_4349,N_4267);
nor U4420 (N_4420,N_4257,N_4359);
or U4421 (N_4421,N_4371,N_4235);
xnor U4422 (N_4422,N_4256,N_4378);
and U4423 (N_4423,N_4345,N_4310);
or U4424 (N_4424,N_4335,N_4201);
or U4425 (N_4425,N_4374,N_4326);
or U4426 (N_4426,N_4357,N_4382);
nor U4427 (N_4427,N_4203,N_4259);
or U4428 (N_4428,N_4260,N_4280);
or U4429 (N_4429,N_4343,N_4331);
and U4430 (N_4430,N_4296,N_4395);
nand U4431 (N_4431,N_4248,N_4337);
and U4432 (N_4432,N_4397,N_4236);
nand U4433 (N_4433,N_4272,N_4288);
nand U4434 (N_4434,N_4354,N_4342);
and U4435 (N_4435,N_4399,N_4347);
or U4436 (N_4436,N_4328,N_4286);
nand U4437 (N_4437,N_4233,N_4293);
and U4438 (N_4438,N_4361,N_4214);
and U4439 (N_4439,N_4322,N_4396);
or U4440 (N_4440,N_4338,N_4234);
nand U4441 (N_4441,N_4391,N_4303);
nor U4442 (N_4442,N_4353,N_4222);
and U4443 (N_4443,N_4244,N_4229);
nand U4444 (N_4444,N_4301,N_4237);
or U4445 (N_4445,N_4336,N_4276);
nand U4446 (N_4446,N_4289,N_4284);
nor U4447 (N_4447,N_4375,N_4304);
nand U4448 (N_4448,N_4376,N_4258);
and U4449 (N_4449,N_4320,N_4394);
nand U4450 (N_4450,N_4299,N_4306);
or U4451 (N_4451,N_4393,N_4277);
xor U4452 (N_4452,N_4362,N_4250);
nor U4453 (N_4453,N_4285,N_4302);
nand U4454 (N_4454,N_4240,N_4212);
or U4455 (N_4455,N_4358,N_4238);
nand U4456 (N_4456,N_4398,N_4307);
or U4457 (N_4457,N_4274,N_4266);
xnor U4458 (N_4458,N_4239,N_4271);
or U4459 (N_4459,N_4213,N_4282);
and U4460 (N_4460,N_4355,N_4262);
and U4461 (N_4461,N_4220,N_4389);
and U4462 (N_4462,N_4241,N_4319);
nor U4463 (N_4463,N_4215,N_4251);
and U4464 (N_4464,N_4261,N_4346);
and U4465 (N_4465,N_4255,N_4205);
xnor U4466 (N_4466,N_4247,N_4313);
nand U4467 (N_4467,N_4243,N_4325);
xor U4468 (N_4468,N_4283,N_4316);
xnor U4469 (N_4469,N_4352,N_4202);
and U4470 (N_4470,N_4246,N_4245);
nand U4471 (N_4471,N_4269,N_4200);
xnor U4472 (N_4472,N_4392,N_4332);
and U4473 (N_4473,N_4311,N_4312);
nand U4474 (N_4474,N_4275,N_4340);
and U4475 (N_4475,N_4360,N_4290);
and U4476 (N_4476,N_4223,N_4305);
nand U4477 (N_4477,N_4339,N_4217);
xor U4478 (N_4478,N_4323,N_4387);
nand U4479 (N_4479,N_4383,N_4384);
or U4480 (N_4480,N_4252,N_4309);
nand U4481 (N_4481,N_4270,N_4225);
or U4482 (N_4482,N_4300,N_4390);
nand U4483 (N_4483,N_4263,N_4365);
and U4484 (N_4484,N_4249,N_4206);
nand U4485 (N_4485,N_4348,N_4297);
nand U4486 (N_4486,N_4315,N_4317);
or U4487 (N_4487,N_4207,N_4209);
and U4488 (N_4488,N_4363,N_4318);
or U4489 (N_4489,N_4370,N_4228);
and U4490 (N_4490,N_4292,N_4308);
nand U4491 (N_4491,N_4281,N_4386);
and U4492 (N_4492,N_4295,N_4218);
nand U4493 (N_4493,N_4327,N_4314);
nand U4494 (N_4494,N_4321,N_4232);
nand U4495 (N_4495,N_4291,N_4208);
nand U4496 (N_4496,N_4279,N_4294);
and U4497 (N_4497,N_4351,N_4373);
and U4498 (N_4498,N_4379,N_4334);
or U4499 (N_4499,N_4230,N_4333);
and U4500 (N_4500,N_4291,N_4202);
and U4501 (N_4501,N_4237,N_4296);
and U4502 (N_4502,N_4352,N_4338);
nand U4503 (N_4503,N_4202,N_4246);
or U4504 (N_4504,N_4320,N_4248);
and U4505 (N_4505,N_4285,N_4353);
or U4506 (N_4506,N_4293,N_4333);
nor U4507 (N_4507,N_4223,N_4362);
or U4508 (N_4508,N_4264,N_4255);
or U4509 (N_4509,N_4279,N_4270);
or U4510 (N_4510,N_4269,N_4320);
or U4511 (N_4511,N_4341,N_4312);
or U4512 (N_4512,N_4311,N_4292);
or U4513 (N_4513,N_4352,N_4284);
xnor U4514 (N_4514,N_4224,N_4258);
nor U4515 (N_4515,N_4311,N_4261);
nand U4516 (N_4516,N_4349,N_4257);
and U4517 (N_4517,N_4201,N_4283);
nor U4518 (N_4518,N_4297,N_4311);
nor U4519 (N_4519,N_4331,N_4312);
nor U4520 (N_4520,N_4390,N_4240);
nor U4521 (N_4521,N_4322,N_4318);
xor U4522 (N_4522,N_4299,N_4281);
nor U4523 (N_4523,N_4365,N_4270);
nor U4524 (N_4524,N_4228,N_4305);
and U4525 (N_4525,N_4322,N_4319);
or U4526 (N_4526,N_4235,N_4336);
and U4527 (N_4527,N_4394,N_4377);
and U4528 (N_4528,N_4232,N_4330);
and U4529 (N_4529,N_4398,N_4375);
nor U4530 (N_4530,N_4333,N_4376);
nand U4531 (N_4531,N_4379,N_4307);
and U4532 (N_4532,N_4256,N_4309);
nor U4533 (N_4533,N_4296,N_4202);
nand U4534 (N_4534,N_4348,N_4357);
nor U4535 (N_4535,N_4279,N_4316);
nor U4536 (N_4536,N_4295,N_4294);
nand U4537 (N_4537,N_4209,N_4389);
xor U4538 (N_4538,N_4302,N_4239);
nor U4539 (N_4539,N_4245,N_4232);
and U4540 (N_4540,N_4266,N_4221);
or U4541 (N_4541,N_4317,N_4286);
and U4542 (N_4542,N_4227,N_4270);
nor U4543 (N_4543,N_4221,N_4218);
or U4544 (N_4544,N_4365,N_4238);
xor U4545 (N_4545,N_4291,N_4362);
nor U4546 (N_4546,N_4320,N_4365);
xor U4547 (N_4547,N_4315,N_4300);
nand U4548 (N_4548,N_4356,N_4230);
or U4549 (N_4549,N_4369,N_4366);
nor U4550 (N_4550,N_4343,N_4356);
or U4551 (N_4551,N_4245,N_4356);
nor U4552 (N_4552,N_4346,N_4258);
nor U4553 (N_4553,N_4215,N_4384);
nor U4554 (N_4554,N_4209,N_4324);
nor U4555 (N_4555,N_4392,N_4257);
xor U4556 (N_4556,N_4237,N_4295);
and U4557 (N_4557,N_4297,N_4212);
nand U4558 (N_4558,N_4330,N_4325);
nand U4559 (N_4559,N_4247,N_4389);
nand U4560 (N_4560,N_4202,N_4383);
or U4561 (N_4561,N_4265,N_4264);
or U4562 (N_4562,N_4352,N_4331);
nand U4563 (N_4563,N_4381,N_4218);
or U4564 (N_4564,N_4254,N_4343);
nor U4565 (N_4565,N_4396,N_4212);
nand U4566 (N_4566,N_4385,N_4391);
and U4567 (N_4567,N_4334,N_4225);
and U4568 (N_4568,N_4210,N_4342);
or U4569 (N_4569,N_4396,N_4226);
and U4570 (N_4570,N_4328,N_4273);
or U4571 (N_4571,N_4232,N_4383);
or U4572 (N_4572,N_4384,N_4283);
or U4573 (N_4573,N_4392,N_4210);
nand U4574 (N_4574,N_4211,N_4245);
nand U4575 (N_4575,N_4343,N_4316);
or U4576 (N_4576,N_4306,N_4368);
nor U4577 (N_4577,N_4320,N_4363);
nor U4578 (N_4578,N_4200,N_4222);
or U4579 (N_4579,N_4243,N_4264);
nand U4580 (N_4580,N_4358,N_4221);
nand U4581 (N_4581,N_4310,N_4340);
or U4582 (N_4582,N_4248,N_4355);
and U4583 (N_4583,N_4259,N_4285);
or U4584 (N_4584,N_4220,N_4342);
xor U4585 (N_4585,N_4212,N_4202);
nand U4586 (N_4586,N_4296,N_4267);
or U4587 (N_4587,N_4277,N_4337);
and U4588 (N_4588,N_4342,N_4274);
and U4589 (N_4589,N_4373,N_4200);
nand U4590 (N_4590,N_4338,N_4365);
or U4591 (N_4591,N_4333,N_4295);
and U4592 (N_4592,N_4351,N_4278);
or U4593 (N_4593,N_4240,N_4340);
nand U4594 (N_4594,N_4222,N_4334);
or U4595 (N_4595,N_4249,N_4269);
or U4596 (N_4596,N_4389,N_4372);
nor U4597 (N_4597,N_4336,N_4290);
or U4598 (N_4598,N_4383,N_4221);
xnor U4599 (N_4599,N_4376,N_4355);
and U4600 (N_4600,N_4453,N_4419);
nand U4601 (N_4601,N_4538,N_4413);
or U4602 (N_4602,N_4442,N_4591);
nor U4603 (N_4603,N_4564,N_4422);
or U4604 (N_4604,N_4416,N_4411);
or U4605 (N_4605,N_4496,N_4487);
or U4606 (N_4606,N_4575,N_4465);
and U4607 (N_4607,N_4503,N_4596);
and U4608 (N_4608,N_4435,N_4414);
nand U4609 (N_4609,N_4433,N_4463);
nand U4610 (N_4610,N_4527,N_4502);
or U4611 (N_4611,N_4511,N_4499);
nor U4612 (N_4612,N_4535,N_4532);
or U4613 (N_4613,N_4461,N_4512);
nand U4614 (N_4614,N_4425,N_4500);
nand U4615 (N_4615,N_4428,N_4405);
and U4616 (N_4616,N_4450,N_4521);
nand U4617 (N_4617,N_4448,N_4455);
or U4618 (N_4618,N_4477,N_4597);
nand U4619 (N_4619,N_4529,N_4451);
nor U4620 (N_4620,N_4443,N_4436);
or U4621 (N_4621,N_4548,N_4545);
nor U4622 (N_4622,N_4452,N_4472);
nor U4623 (N_4623,N_4546,N_4558);
or U4624 (N_4624,N_4404,N_4526);
or U4625 (N_4625,N_4515,N_4439);
and U4626 (N_4626,N_4480,N_4508);
nand U4627 (N_4627,N_4454,N_4509);
nor U4628 (N_4628,N_4506,N_4458);
or U4629 (N_4629,N_4534,N_4491);
nand U4630 (N_4630,N_4549,N_4479);
and U4631 (N_4631,N_4577,N_4468);
nand U4632 (N_4632,N_4493,N_4434);
or U4633 (N_4633,N_4584,N_4449);
and U4634 (N_4634,N_4483,N_4554);
or U4635 (N_4635,N_4482,N_4424);
or U4636 (N_4636,N_4557,N_4423);
or U4637 (N_4637,N_4542,N_4516);
and U4638 (N_4638,N_4490,N_4498);
nor U4639 (N_4639,N_4444,N_4523);
xor U4640 (N_4640,N_4410,N_4488);
and U4641 (N_4641,N_4562,N_4589);
xnor U4642 (N_4642,N_4580,N_4570);
nor U4643 (N_4643,N_4486,N_4525);
nand U4644 (N_4644,N_4456,N_4569);
xnor U4645 (N_4645,N_4406,N_4581);
nand U4646 (N_4646,N_4524,N_4447);
nor U4647 (N_4647,N_4478,N_4530);
or U4648 (N_4648,N_4507,N_4550);
nor U4649 (N_4649,N_4494,N_4475);
xor U4650 (N_4650,N_4553,N_4528);
and U4651 (N_4651,N_4418,N_4537);
and U4652 (N_4652,N_4421,N_4407);
or U4653 (N_4653,N_4539,N_4441);
xnor U4654 (N_4654,N_4544,N_4573);
and U4655 (N_4655,N_4565,N_4552);
or U4656 (N_4656,N_4420,N_4590);
or U4657 (N_4657,N_4531,N_4547);
nand U4658 (N_4658,N_4430,N_4586);
or U4659 (N_4659,N_4576,N_4473);
nor U4660 (N_4660,N_4559,N_4466);
xor U4661 (N_4661,N_4476,N_4540);
nand U4662 (N_4662,N_4460,N_4459);
nand U4663 (N_4663,N_4464,N_4440);
or U4664 (N_4664,N_4401,N_4536);
or U4665 (N_4665,N_4415,N_4403);
or U4666 (N_4666,N_4594,N_4560);
nor U4667 (N_4667,N_4431,N_4595);
and U4668 (N_4668,N_4568,N_4574);
xnor U4669 (N_4669,N_4518,N_4501);
nand U4670 (N_4670,N_4481,N_4582);
and U4671 (N_4671,N_4438,N_4513);
nor U4672 (N_4672,N_4572,N_4563);
or U4673 (N_4673,N_4543,N_4571);
and U4674 (N_4674,N_4587,N_4519);
nand U4675 (N_4675,N_4445,N_4588);
nor U4676 (N_4676,N_4599,N_4583);
xor U4677 (N_4677,N_4432,N_4426);
and U4678 (N_4678,N_4514,N_4485);
and U4679 (N_4679,N_4578,N_4400);
or U4680 (N_4680,N_4593,N_4489);
or U4681 (N_4681,N_4427,N_4592);
and U4682 (N_4682,N_4522,N_4495);
and U4683 (N_4683,N_4505,N_4470);
and U4684 (N_4684,N_4541,N_4492);
nor U4685 (N_4685,N_4484,N_4408);
and U4686 (N_4686,N_4497,N_4504);
nand U4687 (N_4687,N_4412,N_4417);
and U4688 (N_4688,N_4520,N_4471);
and U4689 (N_4689,N_4533,N_4579);
or U4690 (N_4690,N_4561,N_4517);
and U4691 (N_4691,N_4556,N_4467);
xor U4692 (N_4692,N_4566,N_4437);
and U4693 (N_4693,N_4598,N_4402);
nand U4694 (N_4694,N_4409,N_4585);
or U4695 (N_4695,N_4474,N_4555);
and U4696 (N_4696,N_4429,N_4551);
nor U4697 (N_4697,N_4446,N_4510);
or U4698 (N_4698,N_4462,N_4469);
or U4699 (N_4699,N_4567,N_4457);
nand U4700 (N_4700,N_4519,N_4422);
or U4701 (N_4701,N_4403,N_4534);
or U4702 (N_4702,N_4416,N_4413);
xor U4703 (N_4703,N_4543,N_4558);
and U4704 (N_4704,N_4549,N_4469);
nand U4705 (N_4705,N_4539,N_4578);
xor U4706 (N_4706,N_4462,N_4465);
xor U4707 (N_4707,N_4572,N_4496);
or U4708 (N_4708,N_4423,N_4519);
and U4709 (N_4709,N_4453,N_4416);
nor U4710 (N_4710,N_4508,N_4488);
nor U4711 (N_4711,N_4500,N_4419);
and U4712 (N_4712,N_4558,N_4429);
xnor U4713 (N_4713,N_4492,N_4573);
nor U4714 (N_4714,N_4424,N_4471);
and U4715 (N_4715,N_4588,N_4491);
nor U4716 (N_4716,N_4472,N_4590);
nand U4717 (N_4717,N_4571,N_4501);
and U4718 (N_4718,N_4490,N_4520);
or U4719 (N_4719,N_4590,N_4520);
and U4720 (N_4720,N_4472,N_4489);
and U4721 (N_4721,N_4410,N_4526);
nand U4722 (N_4722,N_4584,N_4516);
nor U4723 (N_4723,N_4542,N_4409);
nand U4724 (N_4724,N_4486,N_4595);
nand U4725 (N_4725,N_4553,N_4441);
nand U4726 (N_4726,N_4454,N_4516);
or U4727 (N_4727,N_4495,N_4413);
or U4728 (N_4728,N_4456,N_4453);
and U4729 (N_4729,N_4415,N_4422);
nor U4730 (N_4730,N_4458,N_4500);
xor U4731 (N_4731,N_4436,N_4575);
xor U4732 (N_4732,N_4535,N_4439);
or U4733 (N_4733,N_4530,N_4552);
and U4734 (N_4734,N_4590,N_4497);
and U4735 (N_4735,N_4470,N_4556);
xnor U4736 (N_4736,N_4580,N_4445);
or U4737 (N_4737,N_4518,N_4410);
and U4738 (N_4738,N_4448,N_4559);
nand U4739 (N_4739,N_4529,N_4560);
nor U4740 (N_4740,N_4509,N_4561);
nand U4741 (N_4741,N_4421,N_4584);
nor U4742 (N_4742,N_4587,N_4555);
xnor U4743 (N_4743,N_4419,N_4546);
or U4744 (N_4744,N_4518,N_4546);
xnor U4745 (N_4745,N_4565,N_4424);
nand U4746 (N_4746,N_4460,N_4413);
and U4747 (N_4747,N_4554,N_4503);
nor U4748 (N_4748,N_4456,N_4441);
nand U4749 (N_4749,N_4575,N_4596);
xnor U4750 (N_4750,N_4452,N_4536);
xnor U4751 (N_4751,N_4422,N_4456);
or U4752 (N_4752,N_4484,N_4556);
nand U4753 (N_4753,N_4541,N_4510);
or U4754 (N_4754,N_4528,N_4590);
xnor U4755 (N_4755,N_4480,N_4494);
and U4756 (N_4756,N_4442,N_4456);
and U4757 (N_4757,N_4451,N_4417);
xor U4758 (N_4758,N_4525,N_4574);
or U4759 (N_4759,N_4466,N_4409);
nor U4760 (N_4760,N_4430,N_4587);
nand U4761 (N_4761,N_4568,N_4466);
and U4762 (N_4762,N_4523,N_4405);
xnor U4763 (N_4763,N_4556,N_4580);
and U4764 (N_4764,N_4466,N_4480);
nor U4765 (N_4765,N_4423,N_4469);
xor U4766 (N_4766,N_4407,N_4513);
or U4767 (N_4767,N_4481,N_4432);
nand U4768 (N_4768,N_4539,N_4533);
nor U4769 (N_4769,N_4502,N_4591);
nor U4770 (N_4770,N_4404,N_4462);
nand U4771 (N_4771,N_4414,N_4517);
nand U4772 (N_4772,N_4482,N_4531);
xnor U4773 (N_4773,N_4445,N_4581);
nand U4774 (N_4774,N_4475,N_4491);
and U4775 (N_4775,N_4410,N_4470);
nand U4776 (N_4776,N_4539,N_4553);
nor U4777 (N_4777,N_4547,N_4500);
nand U4778 (N_4778,N_4586,N_4434);
xor U4779 (N_4779,N_4416,N_4531);
nand U4780 (N_4780,N_4451,N_4516);
or U4781 (N_4781,N_4516,N_4559);
and U4782 (N_4782,N_4569,N_4424);
and U4783 (N_4783,N_4541,N_4444);
or U4784 (N_4784,N_4589,N_4487);
nor U4785 (N_4785,N_4514,N_4403);
nor U4786 (N_4786,N_4415,N_4458);
nor U4787 (N_4787,N_4422,N_4527);
xnor U4788 (N_4788,N_4403,N_4417);
nor U4789 (N_4789,N_4518,N_4539);
and U4790 (N_4790,N_4477,N_4542);
nor U4791 (N_4791,N_4429,N_4421);
nand U4792 (N_4792,N_4482,N_4581);
or U4793 (N_4793,N_4447,N_4592);
and U4794 (N_4794,N_4569,N_4564);
nand U4795 (N_4795,N_4554,N_4446);
or U4796 (N_4796,N_4549,N_4448);
or U4797 (N_4797,N_4507,N_4466);
nand U4798 (N_4798,N_4538,N_4427);
nand U4799 (N_4799,N_4554,N_4478);
or U4800 (N_4800,N_4761,N_4782);
nand U4801 (N_4801,N_4726,N_4693);
and U4802 (N_4802,N_4680,N_4634);
nor U4803 (N_4803,N_4718,N_4626);
nor U4804 (N_4804,N_4749,N_4662);
or U4805 (N_4805,N_4724,N_4796);
and U4806 (N_4806,N_4739,N_4745);
or U4807 (N_4807,N_4741,N_4672);
nor U4808 (N_4808,N_4678,N_4635);
nand U4809 (N_4809,N_4661,N_4648);
nor U4810 (N_4810,N_4689,N_4729);
or U4811 (N_4811,N_4752,N_4730);
or U4812 (N_4812,N_4631,N_4719);
nor U4813 (N_4813,N_4751,N_4688);
nand U4814 (N_4814,N_4600,N_4740);
xnor U4815 (N_4815,N_4673,N_4628);
nand U4816 (N_4816,N_4615,N_4613);
and U4817 (N_4817,N_4647,N_4696);
and U4818 (N_4818,N_4799,N_4694);
nand U4819 (N_4819,N_4715,N_4797);
nor U4820 (N_4820,N_4731,N_4670);
nand U4821 (N_4821,N_4620,N_4775);
nor U4822 (N_4822,N_4649,N_4706);
and U4823 (N_4823,N_4603,N_4608);
nand U4824 (N_4824,N_4792,N_4607);
and U4825 (N_4825,N_4742,N_4777);
and U4826 (N_4826,N_4760,N_4612);
nand U4827 (N_4827,N_4755,N_4747);
nand U4828 (N_4828,N_4733,N_4703);
and U4829 (N_4829,N_4734,N_4683);
nand U4830 (N_4830,N_4714,N_4707);
and U4831 (N_4831,N_4687,N_4666);
nor U4832 (N_4832,N_4682,N_4723);
and U4833 (N_4833,N_4676,N_4643);
or U4834 (N_4834,N_4681,N_4767);
nand U4835 (N_4835,N_4717,N_4786);
or U4836 (N_4836,N_4732,N_4757);
nand U4837 (N_4837,N_4765,N_4646);
or U4838 (N_4838,N_4675,N_4667);
and U4839 (N_4839,N_4785,N_4686);
xor U4840 (N_4840,N_4651,N_4737);
and U4841 (N_4841,N_4617,N_4788);
or U4842 (N_4842,N_4669,N_4611);
and U4843 (N_4843,N_4602,N_4684);
and U4844 (N_4844,N_4779,N_4754);
nand U4845 (N_4845,N_4787,N_4633);
or U4846 (N_4846,N_4618,N_4708);
nor U4847 (N_4847,N_4798,N_4795);
and U4848 (N_4848,N_4790,N_4710);
nand U4849 (N_4849,N_4699,N_4709);
and U4850 (N_4850,N_4697,N_4623);
nor U4851 (N_4851,N_4606,N_4664);
xnor U4852 (N_4852,N_4776,N_4770);
and U4853 (N_4853,N_4654,N_4627);
nor U4854 (N_4854,N_4698,N_4748);
nand U4855 (N_4855,N_4789,N_4690);
nor U4856 (N_4856,N_4668,N_4711);
nor U4857 (N_4857,N_4639,N_4636);
xnor U4858 (N_4858,N_4658,N_4625);
nand U4859 (N_4859,N_4736,N_4728);
nand U4860 (N_4860,N_4665,N_4783);
nor U4861 (N_4861,N_4605,N_4604);
nand U4862 (N_4862,N_4660,N_4705);
nand U4863 (N_4863,N_4624,N_4771);
nand U4864 (N_4864,N_4677,N_4663);
or U4865 (N_4865,N_4614,N_4784);
and U4866 (N_4866,N_4691,N_4721);
and U4867 (N_4867,N_4794,N_4743);
and U4868 (N_4868,N_4645,N_4629);
nor U4869 (N_4869,N_4657,N_4764);
nand U4870 (N_4870,N_4685,N_4762);
and U4871 (N_4871,N_4632,N_4656);
or U4872 (N_4872,N_4744,N_4753);
and U4873 (N_4873,N_4641,N_4701);
or U4874 (N_4874,N_4778,N_4791);
nand U4875 (N_4875,N_4758,N_4713);
xor U4876 (N_4876,N_4781,N_4652);
and U4877 (N_4877,N_4712,N_4769);
nor U4878 (N_4878,N_4746,N_4735);
nand U4879 (N_4879,N_4638,N_4637);
and U4880 (N_4880,N_4716,N_4601);
nand U4881 (N_4881,N_4619,N_4610);
or U4882 (N_4882,N_4702,N_4609);
and U4883 (N_4883,N_4679,N_4642);
xnor U4884 (N_4884,N_4750,N_4738);
nand U4885 (N_4885,N_4630,N_4756);
and U4886 (N_4886,N_4704,N_4759);
nor U4887 (N_4887,N_4720,N_4700);
nand U4888 (N_4888,N_4722,N_4793);
xnor U4889 (N_4889,N_4616,N_4780);
or U4890 (N_4890,N_4659,N_4766);
and U4891 (N_4891,N_4727,N_4621);
nor U4892 (N_4892,N_4692,N_4653);
nand U4893 (N_4893,N_4725,N_4644);
nor U4894 (N_4894,N_4772,N_4674);
nor U4895 (N_4895,N_4695,N_4768);
nor U4896 (N_4896,N_4671,N_4640);
nor U4897 (N_4897,N_4763,N_4655);
xnor U4898 (N_4898,N_4622,N_4773);
nor U4899 (N_4899,N_4774,N_4650);
nand U4900 (N_4900,N_4662,N_4774);
xor U4901 (N_4901,N_4688,N_4651);
xnor U4902 (N_4902,N_4757,N_4746);
xor U4903 (N_4903,N_4769,N_4612);
nor U4904 (N_4904,N_4674,N_4715);
and U4905 (N_4905,N_4766,N_4783);
or U4906 (N_4906,N_4632,N_4792);
or U4907 (N_4907,N_4681,N_4755);
and U4908 (N_4908,N_4709,N_4778);
nor U4909 (N_4909,N_4712,N_4632);
nand U4910 (N_4910,N_4626,N_4794);
nor U4911 (N_4911,N_4720,N_4704);
nor U4912 (N_4912,N_4655,N_4600);
xnor U4913 (N_4913,N_4685,N_4642);
or U4914 (N_4914,N_4641,N_4700);
nor U4915 (N_4915,N_4663,N_4669);
nor U4916 (N_4916,N_4630,N_4746);
nor U4917 (N_4917,N_4699,N_4668);
and U4918 (N_4918,N_4769,N_4747);
xnor U4919 (N_4919,N_4647,N_4633);
or U4920 (N_4920,N_4797,N_4649);
or U4921 (N_4921,N_4667,N_4700);
nor U4922 (N_4922,N_4609,N_4666);
and U4923 (N_4923,N_4773,N_4629);
or U4924 (N_4924,N_4734,N_4702);
or U4925 (N_4925,N_4657,N_4627);
nand U4926 (N_4926,N_4770,N_4797);
or U4927 (N_4927,N_4725,N_4733);
or U4928 (N_4928,N_4727,N_4729);
and U4929 (N_4929,N_4639,N_4764);
or U4930 (N_4930,N_4623,N_4720);
nand U4931 (N_4931,N_4702,N_4790);
and U4932 (N_4932,N_4740,N_4790);
or U4933 (N_4933,N_4662,N_4778);
or U4934 (N_4934,N_4757,N_4794);
nor U4935 (N_4935,N_4694,N_4731);
nand U4936 (N_4936,N_4629,N_4664);
and U4937 (N_4937,N_4752,N_4635);
nor U4938 (N_4938,N_4775,N_4788);
nand U4939 (N_4939,N_4610,N_4713);
nand U4940 (N_4940,N_4613,N_4702);
nor U4941 (N_4941,N_4762,N_4733);
or U4942 (N_4942,N_4711,N_4783);
or U4943 (N_4943,N_4645,N_4678);
nand U4944 (N_4944,N_4610,N_4699);
xor U4945 (N_4945,N_4636,N_4733);
nand U4946 (N_4946,N_4732,N_4799);
nand U4947 (N_4947,N_4794,N_4701);
nor U4948 (N_4948,N_4692,N_4694);
nor U4949 (N_4949,N_4701,N_4681);
or U4950 (N_4950,N_4754,N_4756);
nand U4951 (N_4951,N_4666,N_4665);
nand U4952 (N_4952,N_4774,N_4784);
xor U4953 (N_4953,N_4637,N_4757);
or U4954 (N_4954,N_4653,N_4668);
nor U4955 (N_4955,N_4771,N_4789);
nand U4956 (N_4956,N_4657,N_4646);
or U4957 (N_4957,N_4780,N_4625);
nor U4958 (N_4958,N_4703,N_4766);
and U4959 (N_4959,N_4772,N_4773);
and U4960 (N_4960,N_4775,N_4659);
and U4961 (N_4961,N_4607,N_4681);
nor U4962 (N_4962,N_4681,N_4673);
nor U4963 (N_4963,N_4672,N_4601);
nand U4964 (N_4964,N_4616,N_4715);
nand U4965 (N_4965,N_4694,N_4729);
nand U4966 (N_4966,N_4706,N_4743);
and U4967 (N_4967,N_4693,N_4706);
nand U4968 (N_4968,N_4711,N_4754);
nor U4969 (N_4969,N_4786,N_4619);
nand U4970 (N_4970,N_4687,N_4639);
nor U4971 (N_4971,N_4765,N_4652);
xnor U4972 (N_4972,N_4673,N_4760);
or U4973 (N_4973,N_4626,N_4665);
xor U4974 (N_4974,N_4786,N_4711);
xor U4975 (N_4975,N_4775,N_4785);
and U4976 (N_4976,N_4722,N_4682);
nor U4977 (N_4977,N_4703,N_4634);
and U4978 (N_4978,N_4688,N_4659);
nand U4979 (N_4979,N_4667,N_4737);
and U4980 (N_4980,N_4687,N_4637);
xor U4981 (N_4981,N_4714,N_4679);
nand U4982 (N_4982,N_4626,N_4732);
nand U4983 (N_4983,N_4636,N_4611);
xnor U4984 (N_4984,N_4643,N_4686);
xnor U4985 (N_4985,N_4733,N_4635);
or U4986 (N_4986,N_4679,N_4767);
nand U4987 (N_4987,N_4744,N_4738);
nor U4988 (N_4988,N_4637,N_4773);
and U4989 (N_4989,N_4739,N_4666);
and U4990 (N_4990,N_4646,N_4618);
or U4991 (N_4991,N_4683,N_4639);
or U4992 (N_4992,N_4741,N_4770);
nor U4993 (N_4993,N_4613,N_4771);
and U4994 (N_4994,N_4718,N_4708);
xor U4995 (N_4995,N_4698,N_4625);
nor U4996 (N_4996,N_4662,N_4739);
nand U4997 (N_4997,N_4733,N_4795);
xnor U4998 (N_4998,N_4725,N_4711);
or U4999 (N_4999,N_4702,N_4616);
or U5000 (N_5000,N_4880,N_4941);
and U5001 (N_5001,N_4949,N_4802);
and U5002 (N_5002,N_4887,N_4938);
nor U5003 (N_5003,N_4857,N_4839);
or U5004 (N_5004,N_4813,N_4803);
and U5005 (N_5005,N_4851,N_4969);
nor U5006 (N_5006,N_4807,N_4928);
nor U5007 (N_5007,N_4906,N_4821);
nor U5008 (N_5008,N_4934,N_4800);
and U5009 (N_5009,N_4873,N_4988);
and U5010 (N_5010,N_4832,N_4844);
nand U5011 (N_5011,N_4859,N_4817);
nand U5012 (N_5012,N_4852,N_4916);
or U5013 (N_5013,N_4840,N_4862);
nand U5014 (N_5014,N_4885,N_4995);
nor U5015 (N_5015,N_4897,N_4868);
and U5016 (N_5016,N_4922,N_4948);
nor U5017 (N_5017,N_4875,N_4984);
and U5018 (N_5018,N_4828,N_4831);
or U5019 (N_5019,N_4804,N_4894);
nor U5020 (N_5020,N_4900,N_4842);
nor U5021 (N_5021,N_4892,N_4838);
nand U5022 (N_5022,N_4856,N_4958);
and U5023 (N_5023,N_4972,N_4964);
nor U5024 (N_5024,N_4991,N_4836);
or U5025 (N_5025,N_4891,N_4915);
xor U5026 (N_5026,N_4952,N_4884);
xnor U5027 (N_5027,N_4912,N_4823);
nand U5028 (N_5028,N_4886,N_4858);
and U5029 (N_5029,N_4945,N_4806);
or U5030 (N_5030,N_4975,N_4933);
and U5031 (N_5031,N_4968,N_4983);
nor U5032 (N_5032,N_4872,N_4827);
xor U5033 (N_5033,N_4919,N_4937);
nor U5034 (N_5034,N_4911,N_4973);
nor U5035 (N_5035,N_4965,N_4888);
nor U5036 (N_5036,N_4801,N_4951);
or U5037 (N_5037,N_4986,N_4850);
nor U5038 (N_5038,N_4895,N_4942);
nand U5039 (N_5039,N_4847,N_4816);
or U5040 (N_5040,N_4960,N_4898);
nand U5041 (N_5041,N_4905,N_4819);
and U5042 (N_5042,N_4917,N_4955);
and U5043 (N_5043,N_4853,N_4864);
and U5044 (N_5044,N_4870,N_4910);
nor U5045 (N_5045,N_4902,N_4878);
nand U5046 (N_5046,N_4861,N_4904);
nand U5047 (N_5047,N_4876,N_4914);
and U5048 (N_5048,N_4987,N_4849);
or U5049 (N_5049,N_4907,N_4953);
nor U5050 (N_5050,N_4971,N_4903);
nor U5051 (N_5051,N_4855,N_4996);
and U5052 (N_5052,N_4967,N_4976);
xor U5053 (N_5053,N_4963,N_4959);
nand U5054 (N_5054,N_4982,N_4820);
nor U5055 (N_5055,N_4863,N_4989);
nor U5056 (N_5056,N_4814,N_4909);
or U5057 (N_5057,N_4981,N_4860);
nand U5058 (N_5058,N_4822,N_4883);
or U5059 (N_5059,N_4843,N_4815);
nand U5060 (N_5060,N_4936,N_4829);
nor U5061 (N_5061,N_4825,N_4923);
nor U5062 (N_5062,N_4935,N_4845);
xor U5063 (N_5063,N_4824,N_4833);
and U5064 (N_5064,N_4961,N_4956);
and U5065 (N_5065,N_4834,N_4871);
nor U5066 (N_5066,N_4882,N_4990);
xor U5067 (N_5067,N_4893,N_4865);
xnor U5068 (N_5068,N_4966,N_4946);
or U5069 (N_5069,N_4826,N_4947);
nor U5070 (N_5070,N_4877,N_4970);
or U5071 (N_5071,N_4921,N_4978);
or U5072 (N_5072,N_4944,N_4908);
nor U5073 (N_5073,N_4889,N_4927);
and U5074 (N_5074,N_4818,N_4931);
xnor U5075 (N_5075,N_4929,N_4930);
and U5076 (N_5076,N_4866,N_4925);
and U5077 (N_5077,N_4962,N_4950);
and U5078 (N_5078,N_4854,N_4993);
or U5079 (N_5079,N_4837,N_4998);
nor U5080 (N_5080,N_4899,N_4901);
xnor U5081 (N_5081,N_4999,N_4874);
nor U5082 (N_5082,N_4943,N_4805);
and U5083 (N_5083,N_4939,N_4997);
nand U5084 (N_5084,N_4810,N_4812);
and U5085 (N_5085,N_4830,N_4926);
nor U5086 (N_5086,N_4835,N_4924);
nand U5087 (N_5087,N_4977,N_4867);
xor U5088 (N_5088,N_4980,N_4974);
and U5089 (N_5089,N_4881,N_4811);
and U5090 (N_5090,N_4841,N_4954);
nand U5091 (N_5091,N_4869,N_4879);
nor U5092 (N_5092,N_4932,N_4846);
nor U5093 (N_5093,N_4809,N_4985);
or U5094 (N_5094,N_4913,N_4992);
nand U5095 (N_5095,N_4896,N_4808);
xor U5096 (N_5096,N_4848,N_4890);
nor U5097 (N_5097,N_4994,N_4979);
nor U5098 (N_5098,N_4957,N_4918);
and U5099 (N_5099,N_4940,N_4920);
nand U5100 (N_5100,N_4968,N_4887);
nand U5101 (N_5101,N_4847,N_4899);
nor U5102 (N_5102,N_4952,N_4843);
and U5103 (N_5103,N_4829,N_4831);
nor U5104 (N_5104,N_4992,N_4889);
or U5105 (N_5105,N_4841,N_4990);
xor U5106 (N_5106,N_4988,N_4944);
nand U5107 (N_5107,N_4911,N_4838);
nand U5108 (N_5108,N_4857,N_4897);
nor U5109 (N_5109,N_4803,N_4901);
and U5110 (N_5110,N_4976,N_4895);
nand U5111 (N_5111,N_4975,N_4962);
and U5112 (N_5112,N_4826,N_4813);
and U5113 (N_5113,N_4890,N_4873);
or U5114 (N_5114,N_4953,N_4938);
xnor U5115 (N_5115,N_4895,N_4947);
and U5116 (N_5116,N_4818,N_4988);
or U5117 (N_5117,N_4955,N_4910);
xor U5118 (N_5118,N_4806,N_4876);
nand U5119 (N_5119,N_4946,N_4836);
or U5120 (N_5120,N_4991,N_4980);
nand U5121 (N_5121,N_4955,N_4957);
nand U5122 (N_5122,N_4976,N_4857);
xor U5123 (N_5123,N_4810,N_4802);
and U5124 (N_5124,N_4971,N_4872);
and U5125 (N_5125,N_4843,N_4908);
or U5126 (N_5126,N_4872,N_4940);
nand U5127 (N_5127,N_4898,N_4837);
and U5128 (N_5128,N_4854,N_4930);
nand U5129 (N_5129,N_4914,N_4815);
xor U5130 (N_5130,N_4884,N_4988);
nand U5131 (N_5131,N_4807,N_4980);
or U5132 (N_5132,N_4912,N_4887);
xor U5133 (N_5133,N_4804,N_4810);
and U5134 (N_5134,N_4868,N_4960);
nand U5135 (N_5135,N_4845,N_4996);
xnor U5136 (N_5136,N_4893,N_4873);
nor U5137 (N_5137,N_4915,N_4800);
xor U5138 (N_5138,N_4954,N_4884);
and U5139 (N_5139,N_4810,N_4821);
or U5140 (N_5140,N_4875,N_4828);
and U5141 (N_5141,N_4993,N_4841);
xor U5142 (N_5142,N_4852,N_4859);
nand U5143 (N_5143,N_4959,N_4972);
xor U5144 (N_5144,N_4849,N_4914);
or U5145 (N_5145,N_4892,N_4992);
xor U5146 (N_5146,N_4907,N_4854);
nor U5147 (N_5147,N_4802,N_4820);
nand U5148 (N_5148,N_4980,N_4978);
and U5149 (N_5149,N_4853,N_4841);
nor U5150 (N_5150,N_4998,N_4846);
or U5151 (N_5151,N_4948,N_4845);
or U5152 (N_5152,N_4991,N_4822);
xor U5153 (N_5153,N_4962,N_4969);
or U5154 (N_5154,N_4882,N_4843);
nor U5155 (N_5155,N_4808,N_4871);
xnor U5156 (N_5156,N_4882,N_4809);
and U5157 (N_5157,N_4815,N_4885);
nand U5158 (N_5158,N_4814,N_4873);
and U5159 (N_5159,N_4971,N_4926);
and U5160 (N_5160,N_4918,N_4844);
nand U5161 (N_5161,N_4988,N_4859);
xnor U5162 (N_5162,N_4912,N_4892);
and U5163 (N_5163,N_4804,N_4952);
and U5164 (N_5164,N_4995,N_4841);
or U5165 (N_5165,N_4870,N_4980);
xor U5166 (N_5166,N_4927,N_4899);
or U5167 (N_5167,N_4942,N_4823);
nor U5168 (N_5168,N_4812,N_4963);
nor U5169 (N_5169,N_4879,N_4948);
xor U5170 (N_5170,N_4921,N_4992);
and U5171 (N_5171,N_4999,N_4905);
nand U5172 (N_5172,N_4922,N_4923);
nand U5173 (N_5173,N_4866,N_4845);
nand U5174 (N_5174,N_4992,N_4950);
nand U5175 (N_5175,N_4807,N_4931);
nor U5176 (N_5176,N_4842,N_4963);
nor U5177 (N_5177,N_4965,N_4926);
nor U5178 (N_5178,N_4988,N_4906);
or U5179 (N_5179,N_4903,N_4949);
or U5180 (N_5180,N_4891,N_4971);
nand U5181 (N_5181,N_4929,N_4822);
or U5182 (N_5182,N_4928,N_4861);
xnor U5183 (N_5183,N_4990,N_4970);
or U5184 (N_5184,N_4946,N_4835);
and U5185 (N_5185,N_4802,N_4849);
or U5186 (N_5186,N_4902,N_4837);
and U5187 (N_5187,N_4929,N_4990);
and U5188 (N_5188,N_4945,N_4801);
nand U5189 (N_5189,N_4825,N_4872);
and U5190 (N_5190,N_4866,N_4917);
nor U5191 (N_5191,N_4821,N_4948);
nand U5192 (N_5192,N_4964,N_4896);
and U5193 (N_5193,N_4912,N_4895);
nor U5194 (N_5194,N_4922,N_4975);
or U5195 (N_5195,N_4931,N_4922);
and U5196 (N_5196,N_4870,N_4873);
and U5197 (N_5197,N_4879,N_4935);
nor U5198 (N_5198,N_4948,N_4907);
nand U5199 (N_5199,N_4981,N_4922);
and U5200 (N_5200,N_5004,N_5139);
nor U5201 (N_5201,N_5006,N_5007);
or U5202 (N_5202,N_5110,N_5131);
or U5203 (N_5203,N_5099,N_5072);
nor U5204 (N_5204,N_5050,N_5146);
nand U5205 (N_5205,N_5136,N_5065);
or U5206 (N_5206,N_5103,N_5085);
nor U5207 (N_5207,N_5002,N_5119);
or U5208 (N_5208,N_5156,N_5032);
or U5209 (N_5209,N_5198,N_5039);
nand U5210 (N_5210,N_5121,N_5056);
and U5211 (N_5211,N_5143,N_5134);
or U5212 (N_5212,N_5080,N_5083);
and U5213 (N_5213,N_5074,N_5003);
nand U5214 (N_5214,N_5116,N_5027);
xor U5215 (N_5215,N_5190,N_5167);
nand U5216 (N_5216,N_5114,N_5186);
or U5217 (N_5217,N_5015,N_5047);
xor U5218 (N_5218,N_5055,N_5071);
and U5219 (N_5219,N_5158,N_5035);
or U5220 (N_5220,N_5140,N_5057);
xor U5221 (N_5221,N_5070,N_5175);
xor U5222 (N_5222,N_5177,N_5097);
nor U5223 (N_5223,N_5094,N_5008);
or U5224 (N_5224,N_5126,N_5076);
nand U5225 (N_5225,N_5092,N_5081);
and U5226 (N_5226,N_5033,N_5005);
xor U5227 (N_5227,N_5090,N_5195);
or U5228 (N_5228,N_5107,N_5012);
nor U5229 (N_5229,N_5061,N_5191);
nand U5230 (N_5230,N_5066,N_5113);
and U5231 (N_5231,N_5171,N_5182);
and U5232 (N_5232,N_5095,N_5051);
nor U5233 (N_5233,N_5170,N_5180);
and U5234 (N_5234,N_5105,N_5043);
nand U5235 (N_5235,N_5154,N_5155);
nand U5236 (N_5236,N_5045,N_5001);
nor U5237 (N_5237,N_5168,N_5135);
nor U5238 (N_5238,N_5075,N_5166);
and U5239 (N_5239,N_5049,N_5188);
or U5240 (N_5240,N_5069,N_5160);
nand U5241 (N_5241,N_5023,N_5029);
xnor U5242 (N_5242,N_5184,N_5125);
nand U5243 (N_5243,N_5054,N_5174);
nand U5244 (N_5244,N_5151,N_5025);
nor U5245 (N_5245,N_5009,N_5152);
and U5246 (N_5246,N_5123,N_5102);
and U5247 (N_5247,N_5179,N_5141);
or U5248 (N_5248,N_5082,N_5109);
nand U5249 (N_5249,N_5117,N_5089);
nand U5250 (N_5250,N_5017,N_5138);
nand U5251 (N_5251,N_5041,N_5178);
nor U5252 (N_5252,N_5010,N_5192);
nor U5253 (N_5253,N_5064,N_5145);
or U5254 (N_5254,N_5062,N_5127);
xnor U5255 (N_5255,N_5079,N_5000);
nor U5256 (N_5256,N_5181,N_5014);
nand U5257 (N_5257,N_5060,N_5196);
or U5258 (N_5258,N_5164,N_5162);
nor U5259 (N_5259,N_5077,N_5144);
and U5260 (N_5260,N_5183,N_5129);
nor U5261 (N_5261,N_5120,N_5030);
nor U5262 (N_5262,N_5028,N_5172);
nor U5263 (N_5263,N_5068,N_5058);
nand U5264 (N_5264,N_5034,N_5037);
and U5265 (N_5265,N_5091,N_5124);
nand U5266 (N_5266,N_5086,N_5148);
and U5267 (N_5267,N_5026,N_5096);
and U5268 (N_5268,N_5053,N_5147);
or U5269 (N_5269,N_5165,N_5020);
nor U5270 (N_5270,N_5104,N_5031);
or U5271 (N_5271,N_5189,N_5087);
nand U5272 (N_5272,N_5016,N_5197);
nand U5273 (N_5273,N_5022,N_5133);
and U5274 (N_5274,N_5036,N_5169);
nand U5275 (N_5275,N_5024,N_5046);
nor U5276 (N_5276,N_5048,N_5193);
nor U5277 (N_5277,N_5163,N_5059);
or U5278 (N_5278,N_5137,N_5132);
or U5279 (N_5279,N_5159,N_5149);
or U5280 (N_5280,N_5093,N_5044);
and U5281 (N_5281,N_5112,N_5106);
and U5282 (N_5282,N_5173,N_5122);
nand U5283 (N_5283,N_5161,N_5078);
nand U5284 (N_5284,N_5118,N_5052);
or U5285 (N_5285,N_5021,N_5130);
nor U5286 (N_5286,N_5019,N_5115);
and U5287 (N_5287,N_5011,N_5063);
or U5288 (N_5288,N_5018,N_5150);
or U5289 (N_5289,N_5176,N_5042);
or U5290 (N_5290,N_5088,N_5194);
nand U5291 (N_5291,N_5101,N_5108);
or U5292 (N_5292,N_5098,N_5157);
or U5293 (N_5293,N_5067,N_5013);
and U5294 (N_5294,N_5142,N_5187);
nand U5295 (N_5295,N_5084,N_5111);
nand U5296 (N_5296,N_5100,N_5153);
nand U5297 (N_5297,N_5038,N_5073);
or U5298 (N_5298,N_5185,N_5128);
nand U5299 (N_5299,N_5040,N_5199);
nor U5300 (N_5300,N_5101,N_5130);
xnor U5301 (N_5301,N_5002,N_5000);
or U5302 (N_5302,N_5151,N_5125);
xor U5303 (N_5303,N_5064,N_5197);
and U5304 (N_5304,N_5087,N_5123);
nand U5305 (N_5305,N_5106,N_5186);
or U5306 (N_5306,N_5050,N_5168);
nor U5307 (N_5307,N_5164,N_5054);
and U5308 (N_5308,N_5151,N_5044);
nand U5309 (N_5309,N_5089,N_5186);
and U5310 (N_5310,N_5107,N_5102);
and U5311 (N_5311,N_5116,N_5063);
nor U5312 (N_5312,N_5027,N_5098);
nor U5313 (N_5313,N_5086,N_5033);
nand U5314 (N_5314,N_5104,N_5108);
or U5315 (N_5315,N_5085,N_5118);
or U5316 (N_5316,N_5133,N_5026);
and U5317 (N_5317,N_5119,N_5183);
nor U5318 (N_5318,N_5072,N_5151);
nand U5319 (N_5319,N_5147,N_5041);
and U5320 (N_5320,N_5186,N_5079);
nor U5321 (N_5321,N_5065,N_5183);
nor U5322 (N_5322,N_5171,N_5057);
nand U5323 (N_5323,N_5104,N_5128);
and U5324 (N_5324,N_5128,N_5043);
nor U5325 (N_5325,N_5098,N_5022);
xnor U5326 (N_5326,N_5180,N_5159);
nor U5327 (N_5327,N_5134,N_5067);
or U5328 (N_5328,N_5033,N_5012);
xnor U5329 (N_5329,N_5139,N_5195);
nor U5330 (N_5330,N_5183,N_5144);
xnor U5331 (N_5331,N_5008,N_5130);
and U5332 (N_5332,N_5084,N_5072);
nand U5333 (N_5333,N_5072,N_5148);
and U5334 (N_5334,N_5028,N_5070);
nand U5335 (N_5335,N_5052,N_5191);
or U5336 (N_5336,N_5004,N_5044);
and U5337 (N_5337,N_5186,N_5067);
nand U5338 (N_5338,N_5133,N_5163);
or U5339 (N_5339,N_5118,N_5016);
xor U5340 (N_5340,N_5062,N_5031);
or U5341 (N_5341,N_5175,N_5010);
or U5342 (N_5342,N_5131,N_5178);
nor U5343 (N_5343,N_5097,N_5125);
or U5344 (N_5344,N_5155,N_5059);
or U5345 (N_5345,N_5199,N_5042);
nand U5346 (N_5346,N_5056,N_5131);
or U5347 (N_5347,N_5142,N_5092);
or U5348 (N_5348,N_5177,N_5157);
or U5349 (N_5349,N_5134,N_5177);
or U5350 (N_5350,N_5185,N_5142);
and U5351 (N_5351,N_5149,N_5133);
or U5352 (N_5352,N_5035,N_5054);
nor U5353 (N_5353,N_5082,N_5161);
nor U5354 (N_5354,N_5124,N_5148);
nor U5355 (N_5355,N_5071,N_5113);
or U5356 (N_5356,N_5134,N_5062);
and U5357 (N_5357,N_5047,N_5084);
nand U5358 (N_5358,N_5016,N_5196);
or U5359 (N_5359,N_5124,N_5008);
nand U5360 (N_5360,N_5157,N_5156);
and U5361 (N_5361,N_5134,N_5074);
xor U5362 (N_5362,N_5141,N_5148);
nor U5363 (N_5363,N_5106,N_5175);
nand U5364 (N_5364,N_5107,N_5145);
xor U5365 (N_5365,N_5111,N_5016);
nor U5366 (N_5366,N_5073,N_5008);
nor U5367 (N_5367,N_5026,N_5185);
nand U5368 (N_5368,N_5038,N_5095);
and U5369 (N_5369,N_5190,N_5031);
and U5370 (N_5370,N_5184,N_5163);
and U5371 (N_5371,N_5088,N_5016);
nand U5372 (N_5372,N_5192,N_5026);
nand U5373 (N_5373,N_5011,N_5072);
nand U5374 (N_5374,N_5105,N_5025);
nor U5375 (N_5375,N_5079,N_5081);
and U5376 (N_5376,N_5012,N_5034);
nand U5377 (N_5377,N_5117,N_5061);
nor U5378 (N_5378,N_5003,N_5097);
or U5379 (N_5379,N_5072,N_5106);
nor U5380 (N_5380,N_5119,N_5071);
nor U5381 (N_5381,N_5090,N_5057);
or U5382 (N_5382,N_5046,N_5109);
nand U5383 (N_5383,N_5038,N_5108);
xor U5384 (N_5384,N_5184,N_5086);
nand U5385 (N_5385,N_5082,N_5081);
and U5386 (N_5386,N_5184,N_5166);
or U5387 (N_5387,N_5047,N_5043);
or U5388 (N_5388,N_5034,N_5133);
and U5389 (N_5389,N_5172,N_5125);
nand U5390 (N_5390,N_5138,N_5021);
nor U5391 (N_5391,N_5115,N_5174);
nand U5392 (N_5392,N_5076,N_5137);
xnor U5393 (N_5393,N_5069,N_5122);
nor U5394 (N_5394,N_5030,N_5091);
and U5395 (N_5395,N_5127,N_5123);
or U5396 (N_5396,N_5108,N_5006);
and U5397 (N_5397,N_5054,N_5091);
nor U5398 (N_5398,N_5066,N_5185);
nor U5399 (N_5399,N_5163,N_5085);
nor U5400 (N_5400,N_5395,N_5236);
nand U5401 (N_5401,N_5372,N_5388);
and U5402 (N_5402,N_5349,N_5359);
nor U5403 (N_5403,N_5323,N_5383);
and U5404 (N_5404,N_5282,N_5275);
and U5405 (N_5405,N_5342,N_5231);
and U5406 (N_5406,N_5272,N_5271);
nor U5407 (N_5407,N_5295,N_5308);
nor U5408 (N_5408,N_5370,N_5256);
xor U5409 (N_5409,N_5255,N_5226);
or U5410 (N_5410,N_5373,N_5316);
and U5411 (N_5411,N_5322,N_5362);
nor U5412 (N_5412,N_5235,N_5312);
or U5413 (N_5413,N_5343,N_5205);
nand U5414 (N_5414,N_5259,N_5267);
xor U5415 (N_5415,N_5212,N_5348);
xor U5416 (N_5416,N_5218,N_5330);
nand U5417 (N_5417,N_5345,N_5305);
and U5418 (N_5418,N_5274,N_5356);
or U5419 (N_5419,N_5380,N_5306);
and U5420 (N_5420,N_5392,N_5302);
nand U5421 (N_5421,N_5357,N_5368);
nand U5422 (N_5422,N_5332,N_5320);
and U5423 (N_5423,N_5374,N_5394);
nor U5424 (N_5424,N_5281,N_5230);
or U5425 (N_5425,N_5331,N_5228);
and U5426 (N_5426,N_5232,N_5303);
nand U5427 (N_5427,N_5387,N_5384);
and U5428 (N_5428,N_5214,N_5352);
and U5429 (N_5429,N_5240,N_5341);
and U5430 (N_5430,N_5311,N_5333);
nor U5431 (N_5431,N_5225,N_5381);
and U5432 (N_5432,N_5365,N_5293);
or U5433 (N_5433,N_5200,N_5344);
nor U5434 (N_5434,N_5298,N_5215);
and U5435 (N_5435,N_5346,N_5210);
nor U5436 (N_5436,N_5393,N_5340);
nor U5437 (N_5437,N_5337,N_5287);
xnor U5438 (N_5438,N_5277,N_5389);
or U5439 (N_5439,N_5304,N_5278);
and U5440 (N_5440,N_5246,N_5292);
or U5441 (N_5441,N_5309,N_5244);
nor U5442 (N_5442,N_5276,N_5290);
and U5443 (N_5443,N_5334,N_5223);
or U5444 (N_5444,N_5284,N_5329);
nor U5445 (N_5445,N_5375,N_5268);
nor U5446 (N_5446,N_5241,N_5326);
nand U5447 (N_5447,N_5360,N_5251);
nor U5448 (N_5448,N_5361,N_5324);
or U5449 (N_5449,N_5325,N_5297);
nor U5450 (N_5450,N_5310,N_5209);
and U5451 (N_5451,N_5234,N_5318);
or U5452 (N_5452,N_5358,N_5307);
xor U5453 (N_5453,N_5213,N_5364);
or U5454 (N_5454,N_5279,N_5224);
xnor U5455 (N_5455,N_5396,N_5353);
and U5456 (N_5456,N_5204,N_5371);
nand U5457 (N_5457,N_5258,N_5386);
xnor U5458 (N_5458,N_5347,N_5263);
nor U5459 (N_5459,N_5238,N_5203);
and U5460 (N_5460,N_5379,N_5288);
and U5461 (N_5461,N_5296,N_5327);
or U5462 (N_5462,N_5239,N_5222);
nor U5463 (N_5463,N_5350,N_5319);
or U5464 (N_5464,N_5338,N_5206);
nand U5465 (N_5465,N_5243,N_5221);
or U5466 (N_5466,N_5315,N_5351);
or U5467 (N_5467,N_5249,N_5254);
nor U5468 (N_5468,N_5248,N_5207);
nand U5469 (N_5469,N_5314,N_5264);
nand U5470 (N_5470,N_5291,N_5369);
or U5471 (N_5471,N_5220,N_5237);
nand U5472 (N_5472,N_5216,N_5233);
nand U5473 (N_5473,N_5299,N_5300);
nand U5474 (N_5474,N_5313,N_5283);
or U5475 (N_5475,N_5229,N_5363);
xnor U5476 (N_5476,N_5219,N_5266);
nor U5477 (N_5477,N_5398,N_5253);
xnor U5478 (N_5478,N_5382,N_5294);
or U5479 (N_5479,N_5376,N_5366);
nand U5480 (N_5480,N_5257,N_5399);
nor U5481 (N_5481,N_5317,N_5211);
and U5482 (N_5482,N_5367,N_5269);
and U5483 (N_5483,N_5378,N_5335);
and U5484 (N_5484,N_5261,N_5270);
nor U5485 (N_5485,N_5355,N_5289);
nor U5486 (N_5486,N_5201,N_5260);
nor U5487 (N_5487,N_5265,N_5377);
nor U5488 (N_5488,N_5242,N_5202);
nor U5489 (N_5489,N_5247,N_5286);
or U5490 (N_5490,N_5301,N_5250);
and U5491 (N_5491,N_5390,N_5262);
nor U5492 (N_5492,N_5321,N_5285);
and U5493 (N_5493,N_5354,N_5339);
xor U5494 (N_5494,N_5280,N_5245);
xnor U5495 (N_5495,N_5217,N_5397);
and U5496 (N_5496,N_5385,N_5336);
nand U5497 (N_5497,N_5227,N_5252);
or U5498 (N_5498,N_5273,N_5391);
nand U5499 (N_5499,N_5328,N_5208);
nand U5500 (N_5500,N_5377,N_5384);
nor U5501 (N_5501,N_5247,N_5217);
nor U5502 (N_5502,N_5250,N_5314);
nor U5503 (N_5503,N_5252,N_5250);
or U5504 (N_5504,N_5230,N_5381);
or U5505 (N_5505,N_5327,N_5215);
nand U5506 (N_5506,N_5228,N_5374);
and U5507 (N_5507,N_5246,N_5247);
and U5508 (N_5508,N_5319,N_5308);
or U5509 (N_5509,N_5264,N_5277);
nand U5510 (N_5510,N_5280,N_5249);
and U5511 (N_5511,N_5330,N_5333);
or U5512 (N_5512,N_5344,N_5334);
and U5513 (N_5513,N_5365,N_5294);
nand U5514 (N_5514,N_5255,N_5384);
nor U5515 (N_5515,N_5378,N_5345);
or U5516 (N_5516,N_5292,N_5201);
nand U5517 (N_5517,N_5311,N_5349);
and U5518 (N_5518,N_5300,N_5398);
nor U5519 (N_5519,N_5382,N_5231);
or U5520 (N_5520,N_5281,N_5398);
and U5521 (N_5521,N_5261,N_5332);
nor U5522 (N_5522,N_5354,N_5256);
xor U5523 (N_5523,N_5213,N_5246);
or U5524 (N_5524,N_5251,N_5336);
or U5525 (N_5525,N_5200,N_5272);
and U5526 (N_5526,N_5350,N_5216);
nor U5527 (N_5527,N_5338,N_5356);
nand U5528 (N_5528,N_5302,N_5293);
nor U5529 (N_5529,N_5383,N_5385);
and U5530 (N_5530,N_5319,N_5237);
and U5531 (N_5531,N_5267,N_5366);
and U5532 (N_5532,N_5207,N_5381);
nand U5533 (N_5533,N_5394,N_5373);
nand U5534 (N_5534,N_5398,N_5342);
or U5535 (N_5535,N_5355,N_5299);
nand U5536 (N_5536,N_5236,N_5228);
xnor U5537 (N_5537,N_5224,N_5380);
or U5538 (N_5538,N_5261,N_5387);
and U5539 (N_5539,N_5287,N_5362);
nand U5540 (N_5540,N_5365,N_5351);
and U5541 (N_5541,N_5268,N_5250);
nor U5542 (N_5542,N_5209,N_5395);
and U5543 (N_5543,N_5218,N_5372);
nor U5544 (N_5544,N_5326,N_5386);
and U5545 (N_5545,N_5358,N_5382);
nor U5546 (N_5546,N_5374,N_5287);
xor U5547 (N_5547,N_5270,N_5236);
or U5548 (N_5548,N_5332,N_5280);
nor U5549 (N_5549,N_5291,N_5390);
nor U5550 (N_5550,N_5293,N_5321);
nor U5551 (N_5551,N_5266,N_5366);
nor U5552 (N_5552,N_5300,N_5236);
nor U5553 (N_5553,N_5398,N_5202);
xor U5554 (N_5554,N_5211,N_5338);
or U5555 (N_5555,N_5236,N_5282);
nor U5556 (N_5556,N_5387,N_5209);
nor U5557 (N_5557,N_5347,N_5209);
nand U5558 (N_5558,N_5227,N_5258);
nand U5559 (N_5559,N_5216,N_5239);
nor U5560 (N_5560,N_5318,N_5265);
nand U5561 (N_5561,N_5240,N_5229);
nand U5562 (N_5562,N_5283,N_5261);
nor U5563 (N_5563,N_5272,N_5263);
and U5564 (N_5564,N_5203,N_5207);
and U5565 (N_5565,N_5239,N_5284);
nor U5566 (N_5566,N_5373,N_5266);
nand U5567 (N_5567,N_5372,N_5303);
nand U5568 (N_5568,N_5378,N_5237);
and U5569 (N_5569,N_5288,N_5265);
or U5570 (N_5570,N_5384,N_5346);
and U5571 (N_5571,N_5381,N_5274);
nor U5572 (N_5572,N_5380,N_5240);
and U5573 (N_5573,N_5211,N_5264);
and U5574 (N_5574,N_5304,N_5224);
and U5575 (N_5575,N_5343,N_5326);
or U5576 (N_5576,N_5326,N_5324);
xnor U5577 (N_5577,N_5309,N_5276);
nand U5578 (N_5578,N_5271,N_5295);
xnor U5579 (N_5579,N_5263,N_5229);
or U5580 (N_5580,N_5367,N_5285);
nand U5581 (N_5581,N_5258,N_5292);
or U5582 (N_5582,N_5258,N_5389);
nor U5583 (N_5583,N_5251,N_5388);
or U5584 (N_5584,N_5383,N_5285);
and U5585 (N_5585,N_5347,N_5317);
and U5586 (N_5586,N_5375,N_5334);
nand U5587 (N_5587,N_5356,N_5364);
xor U5588 (N_5588,N_5334,N_5237);
nand U5589 (N_5589,N_5366,N_5293);
nand U5590 (N_5590,N_5395,N_5377);
or U5591 (N_5591,N_5388,N_5364);
or U5592 (N_5592,N_5256,N_5316);
and U5593 (N_5593,N_5336,N_5249);
and U5594 (N_5594,N_5205,N_5341);
nor U5595 (N_5595,N_5307,N_5315);
xnor U5596 (N_5596,N_5310,N_5396);
or U5597 (N_5597,N_5298,N_5274);
nand U5598 (N_5598,N_5335,N_5270);
nor U5599 (N_5599,N_5350,N_5364);
nand U5600 (N_5600,N_5581,N_5531);
xor U5601 (N_5601,N_5482,N_5539);
xnor U5602 (N_5602,N_5576,N_5597);
or U5603 (N_5603,N_5588,N_5402);
or U5604 (N_5604,N_5459,N_5544);
and U5605 (N_5605,N_5553,N_5518);
nor U5606 (N_5606,N_5509,N_5444);
and U5607 (N_5607,N_5571,N_5551);
nand U5608 (N_5608,N_5525,N_5593);
nand U5609 (N_5609,N_5421,N_5467);
or U5610 (N_5610,N_5453,N_5503);
or U5611 (N_5611,N_5542,N_5433);
nor U5612 (N_5612,N_5471,N_5489);
xnor U5613 (N_5613,N_5594,N_5549);
and U5614 (N_5614,N_5428,N_5498);
xor U5615 (N_5615,N_5423,N_5454);
or U5616 (N_5616,N_5511,N_5506);
or U5617 (N_5617,N_5592,N_5409);
or U5618 (N_5618,N_5406,N_5480);
xnor U5619 (N_5619,N_5478,N_5439);
nor U5620 (N_5620,N_5432,N_5537);
or U5621 (N_5621,N_5580,N_5475);
or U5622 (N_5622,N_5437,N_5515);
nand U5623 (N_5623,N_5464,N_5570);
and U5624 (N_5624,N_5586,N_5486);
nor U5625 (N_5625,N_5420,N_5513);
or U5626 (N_5626,N_5585,N_5440);
and U5627 (N_5627,N_5441,N_5485);
nand U5628 (N_5628,N_5436,N_5565);
nand U5629 (N_5629,N_5493,N_5410);
and U5630 (N_5630,N_5430,N_5598);
xor U5631 (N_5631,N_5595,N_5448);
nand U5632 (N_5632,N_5522,N_5569);
nand U5633 (N_5633,N_5495,N_5599);
or U5634 (N_5634,N_5589,N_5562);
nand U5635 (N_5635,N_5474,N_5535);
nor U5636 (N_5636,N_5523,N_5465);
xor U5637 (N_5637,N_5443,N_5434);
and U5638 (N_5638,N_5422,N_5456);
and U5639 (N_5639,N_5487,N_5528);
nand U5640 (N_5640,N_5460,N_5527);
nor U5641 (N_5641,N_5572,N_5446);
or U5642 (N_5642,N_5500,N_5488);
and U5643 (N_5643,N_5405,N_5591);
nor U5644 (N_5644,N_5520,N_5529);
or U5645 (N_5645,N_5435,N_5530);
and U5646 (N_5646,N_5419,N_5490);
or U5647 (N_5647,N_5574,N_5557);
or U5648 (N_5648,N_5502,N_5508);
nor U5649 (N_5649,N_5548,N_5533);
and U5650 (N_5650,N_5470,N_5563);
or U5651 (N_5651,N_5554,N_5416);
nand U5652 (N_5652,N_5550,N_5426);
xnor U5653 (N_5653,N_5573,N_5587);
or U5654 (N_5654,N_5457,N_5466);
or U5655 (N_5655,N_5575,N_5479);
and U5656 (N_5656,N_5472,N_5546);
or U5657 (N_5657,N_5558,N_5566);
nor U5658 (N_5658,N_5473,N_5596);
nand U5659 (N_5659,N_5469,N_5510);
xnor U5660 (N_5660,N_5452,N_5438);
or U5661 (N_5661,N_5519,N_5524);
and U5662 (N_5662,N_5484,N_5552);
or U5663 (N_5663,N_5413,N_5564);
nor U5664 (N_5664,N_5577,N_5578);
nor U5665 (N_5665,N_5540,N_5407);
or U5666 (N_5666,N_5494,N_5491);
nor U5667 (N_5667,N_5504,N_5516);
or U5668 (N_5668,N_5497,N_5455);
and U5669 (N_5669,N_5425,N_5538);
nand U5670 (N_5670,N_5481,N_5404);
or U5671 (N_5671,N_5517,N_5555);
nand U5672 (N_5672,N_5417,N_5543);
xor U5673 (N_5673,N_5547,N_5411);
or U5674 (N_5674,N_5477,N_5476);
and U5675 (N_5675,N_5584,N_5521);
nand U5676 (N_5676,N_5496,N_5499);
nand U5677 (N_5677,N_5561,N_5536);
and U5678 (N_5678,N_5445,N_5568);
nor U5679 (N_5679,N_5463,N_5505);
nor U5680 (N_5680,N_5579,N_5458);
and U5681 (N_5681,N_5450,N_5424);
nor U5682 (N_5682,N_5556,N_5451);
nand U5683 (N_5683,N_5461,N_5418);
nor U5684 (N_5684,N_5514,N_5431);
and U5685 (N_5685,N_5449,N_5429);
nor U5686 (N_5686,N_5534,N_5492);
and U5687 (N_5687,N_5501,N_5442);
nand U5688 (N_5688,N_5590,N_5583);
and U5689 (N_5689,N_5415,N_5541);
and U5690 (N_5690,N_5468,N_5427);
nor U5691 (N_5691,N_5462,N_5567);
nor U5692 (N_5692,N_5532,N_5447);
and U5693 (N_5693,N_5400,N_5545);
xnor U5694 (N_5694,N_5403,N_5408);
and U5695 (N_5695,N_5582,N_5526);
nand U5696 (N_5696,N_5512,N_5412);
and U5697 (N_5697,N_5401,N_5559);
or U5698 (N_5698,N_5414,N_5483);
or U5699 (N_5699,N_5560,N_5507);
or U5700 (N_5700,N_5569,N_5515);
nor U5701 (N_5701,N_5464,N_5565);
xnor U5702 (N_5702,N_5400,N_5574);
xnor U5703 (N_5703,N_5435,N_5509);
or U5704 (N_5704,N_5596,N_5531);
and U5705 (N_5705,N_5492,N_5471);
nor U5706 (N_5706,N_5532,N_5482);
or U5707 (N_5707,N_5422,N_5575);
nand U5708 (N_5708,N_5438,N_5434);
nor U5709 (N_5709,N_5526,N_5544);
or U5710 (N_5710,N_5566,N_5501);
or U5711 (N_5711,N_5439,N_5422);
nand U5712 (N_5712,N_5420,N_5593);
nor U5713 (N_5713,N_5428,N_5403);
or U5714 (N_5714,N_5489,N_5453);
nor U5715 (N_5715,N_5507,N_5403);
nand U5716 (N_5716,N_5592,N_5403);
nand U5717 (N_5717,N_5454,N_5583);
or U5718 (N_5718,N_5431,N_5487);
nand U5719 (N_5719,N_5457,N_5558);
xnor U5720 (N_5720,N_5442,N_5467);
or U5721 (N_5721,N_5479,N_5404);
nor U5722 (N_5722,N_5417,N_5435);
or U5723 (N_5723,N_5576,N_5487);
or U5724 (N_5724,N_5504,N_5576);
and U5725 (N_5725,N_5532,N_5491);
and U5726 (N_5726,N_5476,N_5594);
nand U5727 (N_5727,N_5515,N_5480);
and U5728 (N_5728,N_5539,N_5485);
and U5729 (N_5729,N_5585,N_5491);
or U5730 (N_5730,N_5593,N_5572);
nor U5731 (N_5731,N_5516,N_5561);
and U5732 (N_5732,N_5590,N_5440);
or U5733 (N_5733,N_5457,N_5447);
or U5734 (N_5734,N_5460,N_5506);
nor U5735 (N_5735,N_5483,N_5417);
or U5736 (N_5736,N_5548,N_5485);
xnor U5737 (N_5737,N_5457,N_5430);
and U5738 (N_5738,N_5460,N_5491);
or U5739 (N_5739,N_5408,N_5597);
xnor U5740 (N_5740,N_5535,N_5460);
nor U5741 (N_5741,N_5578,N_5583);
nand U5742 (N_5742,N_5522,N_5526);
nand U5743 (N_5743,N_5517,N_5456);
and U5744 (N_5744,N_5585,N_5470);
nand U5745 (N_5745,N_5495,N_5468);
nor U5746 (N_5746,N_5447,N_5445);
and U5747 (N_5747,N_5468,N_5428);
nand U5748 (N_5748,N_5412,N_5453);
nand U5749 (N_5749,N_5554,N_5506);
and U5750 (N_5750,N_5524,N_5561);
nand U5751 (N_5751,N_5448,N_5582);
nor U5752 (N_5752,N_5427,N_5483);
or U5753 (N_5753,N_5428,N_5515);
nor U5754 (N_5754,N_5526,N_5529);
nor U5755 (N_5755,N_5533,N_5411);
or U5756 (N_5756,N_5534,N_5547);
nand U5757 (N_5757,N_5502,N_5593);
and U5758 (N_5758,N_5539,N_5519);
nor U5759 (N_5759,N_5536,N_5502);
xnor U5760 (N_5760,N_5407,N_5430);
nor U5761 (N_5761,N_5486,N_5410);
or U5762 (N_5762,N_5583,N_5421);
nor U5763 (N_5763,N_5481,N_5453);
nor U5764 (N_5764,N_5550,N_5572);
and U5765 (N_5765,N_5403,N_5436);
or U5766 (N_5766,N_5510,N_5417);
nand U5767 (N_5767,N_5455,N_5510);
and U5768 (N_5768,N_5520,N_5464);
xnor U5769 (N_5769,N_5556,N_5421);
and U5770 (N_5770,N_5521,N_5524);
or U5771 (N_5771,N_5541,N_5449);
nand U5772 (N_5772,N_5514,N_5475);
xor U5773 (N_5773,N_5409,N_5560);
and U5774 (N_5774,N_5509,N_5505);
and U5775 (N_5775,N_5529,N_5518);
and U5776 (N_5776,N_5589,N_5466);
and U5777 (N_5777,N_5417,N_5463);
or U5778 (N_5778,N_5482,N_5590);
and U5779 (N_5779,N_5557,N_5595);
nand U5780 (N_5780,N_5576,N_5476);
or U5781 (N_5781,N_5516,N_5434);
nand U5782 (N_5782,N_5524,N_5467);
nor U5783 (N_5783,N_5416,N_5522);
or U5784 (N_5784,N_5580,N_5402);
xnor U5785 (N_5785,N_5511,N_5482);
nand U5786 (N_5786,N_5551,N_5569);
nor U5787 (N_5787,N_5544,N_5470);
nor U5788 (N_5788,N_5461,N_5512);
nor U5789 (N_5789,N_5542,N_5550);
nor U5790 (N_5790,N_5535,N_5523);
nand U5791 (N_5791,N_5588,N_5549);
and U5792 (N_5792,N_5402,N_5533);
or U5793 (N_5793,N_5461,N_5444);
and U5794 (N_5794,N_5412,N_5592);
nand U5795 (N_5795,N_5533,N_5476);
or U5796 (N_5796,N_5555,N_5471);
or U5797 (N_5797,N_5416,N_5583);
or U5798 (N_5798,N_5586,N_5402);
or U5799 (N_5799,N_5574,N_5516);
nor U5800 (N_5800,N_5649,N_5674);
and U5801 (N_5801,N_5710,N_5608);
xor U5802 (N_5802,N_5745,N_5668);
or U5803 (N_5803,N_5645,N_5754);
and U5804 (N_5804,N_5666,N_5619);
xor U5805 (N_5805,N_5627,N_5766);
nand U5806 (N_5806,N_5779,N_5671);
nor U5807 (N_5807,N_5631,N_5798);
nand U5808 (N_5808,N_5615,N_5607);
and U5809 (N_5809,N_5698,N_5688);
nand U5810 (N_5810,N_5634,N_5741);
nand U5811 (N_5811,N_5697,N_5767);
xor U5812 (N_5812,N_5792,N_5647);
nor U5813 (N_5813,N_5667,N_5703);
xnor U5814 (N_5814,N_5772,N_5791);
and U5815 (N_5815,N_5689,N_5675);
xor U5816 (N_5816,N_5795,N_5714);
or U5817 (N_5817,N_5636,N_5611);
and U5818 (N_5818,N_5707,N_5763);
or U5819 (N_5819,N_5764,N_5702);
or U5820 (N_5820,N_5724,N_5782);
xor U5821 (N_5821,N_5635,N_5793);
or U5822 (N_5822,N_5721,N_5693);
or U5823 (N_5823,N_5628,N_5717);
and U5824 (N_5824,N_5663,N_5759);
xnor U5825 (N_5825,N_5643,N_5722);
xnor U5826 (N_5826,N_5650,N_5797);
nand U5827 (N_5827,N_5727,N_5657);
nand U5828 (N_5828,N_5747,N_5659);
nand U5829 (N_5829,N_5736,N_5673);
and U5830 (N_5830,N_5730,N_5774);
or U5831 (N_5831,N_5733,N_5796);
or U5832 (N_5832,N_5648,N_5709);
nor U5833 (N_5833,N_5604,N_5756);
and U5834 (N_5834,N_5755,N_5771);
nand U5835 (N_5835,N_5706,N_5769);
and U5836 (N_5836,N_5713,N_5672);
nor U5837 (N_5837,N_5744,N_5656);
or U5838 (N_5838,N_5732,N_5639);
nor U5839 (N_5839,N_5711,N_5652);
nand U5840 (N_5840,N_5699,N_5638);
xnor U5841 (N_5841,N_5655,N_5644);
nor U5842 (N_5842,N_5662,N_5758);
or U5843 (N_5843,N_5752,N_5790);
or U5844 (N_5844,N_5781,N_5725);
nand U5845 (N_5845,N_5624,N_5614);
and U5846 (N_5846,N_5609,N_5728);
nor U5847 (N_5847,N_5761,N_5603);
nor U5848 (N_5848,N_5762,N_5778);
nor U5849 (N_5849,N_5642,N_5665);
nand U5850 (N_5850,N_5661,N_5632);
xnor U5851 (N_5851,N_5613,N_5677);
nor U5852 (N_5852,N_5687,N_5726);
or U5853 (N_5853,N_5743,N_5640);
and U5854 (N_5854,N_5749,N_5660);
or U5855 (N_5855,N_5770,N_5760);
xnor U5856 (N_5856,N_5601,N_5775);
or U5857 (N_5857,N_5765,N_5701);
or U5858 (N_5858,N_5664,N_5700);
or U5859 (N_5859,N_5641,N_5704);
or U5860 (N_5860,N_5685,N_5718);
nand U5861 (N_5861,N_5794,N_5787);
or U5862 (N_5862,N_5676,N_5788);
and U5863 (N_5863,N_5653,N_5716);
and U5864 (N_5864,N_5626,N_5623);
and U5865 (N_5865,N_5750,N_5696);
nor U5866 (N_5866,N_5786,N_5731);
and U5867 (N_5867,N_5625,N_5637);
nand U5868 (N_5868,N_5669,N_5629);
or U5869 (N_5869,N_5753,N_5684);
nand U5870 (N_5870,N_5633,N_5600);
and U5871 (N_5871,N_5739,N_5683);
nand U5872 (N_5872,N_5617,N_5720);
nor U5873 (N_5873,N_5610,N_5691);
nor U5874 (N_5874,N_5777,N_5602);
or U5875 (N_5875,N_5715,N_5719);
and U5876 (N_5876,N_5692,N_5735);
or U5877 (N_5877,N_5799,N_5751);
nor U5878 (N_5878,N_5646,N_5680);
nand U5879 (N_5879,N_5658,N_5768);
nand U5880 (N_5880,N_5737,N_5682);
nor U5881 (N_5881,N_5738,N_5606);
nand U5882 (N_5882,N_5686,N_5734);
and U5883 (N_5883,N_5748,N_5742);
and U5884 (N_5884,N_5746,N_5776);
and U5885 (N_5885,N_5679,N_5757);
and U5886 (N_5886,N_5740,N_5612);
xnor U5887 (N_5887,N_5705,N_5784);
or U5888 (N_5888,N_5651,N_5780);
nand U5889 (N_5889,N_5681,N_5708);
nor U5890 (N_5890,N_5605,N_5789);
nand U5891 (N_5891,N_5773,N_5618);
nand U5892 (N_5892,N_5622,N_5630);
and U5893 (N_5893,N_5620,N_5723);
or U5894 (N_5894,N_5694,N_5712);
and U5895 (N_5895,N_5654,N_5670);
and U5896 (N_5896,N_5695,N_5783);
or U5897 (N_5897,N_5785,N_5729);
nor U5898 (N_5898,N_5678,N_5690);
nor U5899 (N_5899,N_5616,N_5621);
nand U5900 (N_5900,N_5759,N_5708);
xnor U5901 (N_5901,N_5657,N_5777);
or U5902 (N_5902,N_5723,N_5739);
or U5903 (N_5903,N_5749,N_5738);
and U5904 (N_5904,N_5761,N_5790);
and U5905 (N_5905,N_5722,N_5747);
and U5906 (N_5906,N_5789,N_5780);
and U5907 (N_5907,N_5649,N_5642);
or U5908 (N_5908,N_5741,N_5602);
nand U5909 (N_5909,N_5782,N_5671);
xor U5910 (N_5910,N_5670,N_5655);
nor U5911 (N_5911,N_5663,N_5646);
nor U5912 (N_5912,N_5635,N_5770);
nor U5913 (N_5913,N_5677,N_5744);
or U5914 (N_5914,N_5623,N_5699);
nor U5915 (N_5915,N_5634,N_5734);
nor U5916 (N_5916,N_5705,N_5632);
and U5917 (N_5917,N_5712,N_5732);
and U5918 (N_5918,N_5658,N_5680);
and U5919 (N_5919,N_5728,N_5661);
and U5920 (N_5920,N_5640,N_5656);
and U5921 (N_5921,N_5673,N_5681);
nor U5922 (N_5922,N_5773,N_5783);
nand U5923 (N_5923,N_5608,N_5763);
nand U5924 (N_5924,N_5700,N_5713);
or U5925 (N_5925,N_5772,N_5658);
or U5926 (N_5926,N_5683,N_5790);
nand U5927 (N_5927,N_5698,N_5755);
and U5928 (N_5928,N_5664,N_5654);
nor U5929 (N_5929,N_5747,N_5642);
nor U5930 (N_5930,N_5731,N_5710);
or U5931 (N_5931,N_5742,N_5611);
xor U5932 (N_5932,N_5636,N_5605);
or U5933 (N_5933,N_5696,N_5798);
nor U5934 (N_5934,N_5773,N_5611);
or U5935 (N_5935,N_5678,N_5738);
and U5936 (N_5936,N_5746,N_5605);
nor U5937 (N_5937,N_5726,N_5611);
nor U5938 (N_5938,N_5636,N_5604);
nand U5939 (N_5939,N_5639,N_5711);
nand U5940 (N_5940,N_5706,N_5668);
nand U5941 (N_5941,N_5716,N_5707);
nand U5942 (N_5942,N_5696,N_5714);
or U5943 (N_5943,N_5656,N_5769);
nor U5944 (N_5944,N_5724,N_5720);
and U5945 (N_5945,N_5747,N_5775);
xnor U5946 (N_5946,N_5603,N_5608);
nor U5947 (N_5947,N_5737,N_5733);
or U5948 (N_5948,N_5704,N_5736);
or U5949 (N_5949,N_5647,N_5643);
and U5950 (N_5950,N_5606,N_5720);
nand U5951 (N_5951,N_5631,N_5799);
nor U5952 (N_5952,N_5749,N_5624);
or U5953 (N_5953,N_5737,N_5683);
nor U5954 (N_5954,N_5606,N_5648);
and U5955 (N_5955,N_5638,N_5793);
nor U5956 (N_5956,N_5673,N_5640);
nand U5957 (N_5957,N_5612,N_5689);
nor U5958 (N_5958,N_5689,N_5772);
or U5959 (N_5959,N_5738,N_5788);
and U5960 (N_5960,N_5635,N_5613);
or U5961 (N_5961,N_5621,N_5600);
xor U5962 (N_5962,N_5610,N_5735);
nor U5963 (N_5963,N_5737,N_5639);
and U5964 (N_5964,N_5673,N_5675);
or U5965 (N_5965,N_5668,N_5755);
nor U5966 (N_5966,N_5690,N_5620);
nor U5967 (N_5967,N_5604,N_5798);
nand U5968 (N_5968,N_5602,N_5719);
nand U5969 (N_5969,N_5754,N_5746);
or U5970 (N_5970,N_5686,N_5749);
or U5971 (N_5971,N_5768,N_5665);
nor U5972 (N_5972,N_5701,N_5780);
nor U5973 (N_5973,N_5744,N_5680);
nand U5974 (N_5974,N_5638,N_5652);
nand U5975 (N_5975,N_5702,N_5659);
or U5976 (N_5976,N_5693,N_5731);
nand U5977 (N_5977,N_5775,N_5672);
or U5978 (N_5978,N_5674,N_5774);
and U5979 (N_5979,N_5642,N_5777);
nand U5980 (N_5980,N_5760,N_5757);
and U5981 (N_5981,N_5742,N_5634);
or U5982 (N_5982,N_5798,N_5612);
and U5983 (N_5983,N_5680,N_5677);
or U5984 (N_5984,N_5776,N_5683);
and U5985 (N_5985,N_5699,N_5788);
nor U5986 (N_5986,N_5682,N_5613);
or U5987 (N_5987,N_5612,N_5746);
nor U5988 (N_5988,N_5625,N_5687);
nand U5989 (N_5989,N_5666,N_5716);
nor U5990 (N_5990,N_5713,N_5665);
nor U5991 (N_5991,N_5723,N_5610);
and U5992 (N_5992,N_5772,N_5715);
and U5993 (N_5993,N_5794,N_5620);
nand U5994 (N_5994,N_5626,N_5763);
or U5995 (N_5995,N_5738,N_5780);
nor U5996 (N_5996,N_5611,N_5609);
or U5997 (N_5997,N_5772,N_5759);
nor U5998 (N_5998,N_5730,N_5760);
nand U5999 (N_5999,N_5696,N_5659);
xor U6000 (N_6000,N_5943,N_5908);
xnor U6001 (N_6001,N_5934,N_5832);
or U6002 (N_6002,N_5800,N_5978);
nor U6003 (N_6003,N_5966,N_5801);
nor U6004 (N_6004,N_5836,N_5947);
and U6005 (N_6005,N_5992,N_5925);
nand U6006 (N_6006,N_5887,N_5989);
and U6007 (N_6007,N_5892,N_5927);
and U6008 (N_6008,N_5864,N_5909);
and U6009 (N_6009,N_5866,N_5830);
or U6010 (N_6010,N_5855,N_5842);
and U6011 (N_6011,N_5826,N_5962);
xnor U6012 (N_6012,N_5902,N_5815);
nand U6013 (N_6013,N_5827,N_5813);
and U6014 (N_6014,N_5935,N_5967);
or U6015 (N_6015,N_5999,N_5841);
xnor U6016 (N_6016,N_5984,N_5923);
and U6017 (N_6017,N_5814,N_5876);
or U6018 (N_6018,N_5920,N_5973);
nor U6019 (N_6019,N_5833,N_5901);
nor U6020 (N_6020,N_5911,N_5968);
or U6021 (N_6021,N_5821,N_5904);
and U6022 (N_6022,N_5917,N_5946);
nand U6023 (N_6023,N_5898,N_5955);
nor U6024 (N_6024,N_5959,N_5916);
or U6025 (N_6025,N_5818,N_5961);
nand U6026 (N_6026,N_5964,N_5886);
and U6027 (N_6027,N_5903,N_5996);
nand U6028 (N_6028,N_5882,N_5981);
and U6029 (N_6029,N_5954,N_5912);
xnor U6030 (N_6030,N_5858,N_5806);
nor U6031 (N_6031,N_5867,N_5808);
or U6032 (N_6032,N_5985,N_5889);
nor U6033 (N_6033,N_5939,N_5931);
nor U6034 (N_6034,N_5944,N_5834);
nand U6035 (N_6035,N_5972,N_5899);
nor U6036 (N_6036,N_5915,N_5997);
xor U6037 (N_6037,N_5945,N_5926);
nor U6038 (N_6038,N_5913,N_5872);
nor U6039 (N_6039,N_5822,N_5900);
nor U6040 (N_6040,N_5951,N_5819);
or U6041 (N_6041,N_5845,N_5874);
and U6042 (N_6042,N_5849,N_5844);
or U6043 (N_6043,N_5910,N_5885);
and U6044 (N_6044,N_5896,N_5988);
or U6045 (N_6045,N_5958,N_5879);
nand U6046 (N_6046,N_5969,N_5880);
nand U6047 (N_6047,N_5924,N_5843);
nand U6048 (N_6048,N_5873,N_5853);
nand U6049 (N_6049,N_5930,N_5937);
nand U6050 (N_6050,N_5861,N_5811);
nor U6051 (N_6051,N_5828,N_5809);
nor U6052 (N_6052,N_5979,N_5986);
and U6053 (N_6053,N_5847,N_5825);
and U6054 (N_6054,N_5928,N_5839);
and U6055 (N_6055,N_5810,N_5802);
nand U6056 (N_6056,N_5890,N_5963);
nand U6057 (N_6057,N_5829,N_5871);
nand U6058 (N_6058,N_5993,N_5870);
and U6059 (N_6059,N_5919,N_5998);
or U6060 (N_6060,N_5994,N_5805);
nand U6061 (N_6061,N_5863,N_5938);
and U6062 (N_6062,N_5846,N_5854);
nand U6063 (N_6063,N_5991,N_5862);
nor U6064 (N_6064,N_5893,N_5850);
nor U6065 (N_6065,N_5816,N_5932);
nor U6066 (N_6066,N_5869,N_5953);
nand U6067 (N_6067,N_5990,N_5980);
and U6068 (N_6068,N_5941,N_5949);
nand U6069 (N_6069,N_5987,N_5914);
and U6070 (N_6070,N_5940,N_5965);
nor U6071 (N_6071,N_5976,N_5952);
or U6072 (N_6072,N_5950,N_5868);
nor U6073 (N_6073,N_5957,N_5852);
nand U6074 (N_6074,N_5983,N_5888);
nor U6075 (N_6075,N_5948,N_5936);
or U6076 (N_6076,N_5856,N_5883);
xnor U6077 (N_6077,N_5960,N_5982);
and U6078 (N_6078,N_5831,N_5933);
and U6079 (N_6079,N_5956,N_5977);
nor U6080 (N_6080,N_5812,N_5817);
nor U6081 (N_6081,N_5820,N_5906);
or U6082 (N_6082,N_5881,N_5891);
and U6083 (N_6083,N_5995,N_5974);
xnor U6084 (N_6084,N_5905,N_5851);
and U6085 (N_6085,N_5971,N_5877);
nor U6086 (N_6086,N_5875,N_5895);
or U6087 (N_6087,N_5942,N_5857);
or U6088 (N_6088,N_5838,N_5918);
xnor U6089 (N_6089,N_5929,N_5970);
nand U6090 (N_6090,N_5807,N_5897);
and U6091 (N_6091,N_5884,N_5975);
and U6092 (N_6092,N_5837,N_5894);
or U6093 (N_6093,N_5922,N_5865);
nand U6094 (N_6094,N_5835,N_5859);
and U6095 (N_6095,N_5848,N_5804);
nand U6096 (N_6096,N_5840,N_5823);
nand U6097 (N_6097,N_5803,N_5921);
nand U6098 (N_6098,N_5907,N_5860);
nand U6099 (N_6099,N_5824,N_5878);
or U6100 (N_6100,N_5987,N_5824);
or U6101 (N_6101,N_5886,N_5973);
and U6102 (N_6102,N_5941,N_5861);
or U6103 (N_6103,N_5931,N_5957);
or U6104 (N_6104,N_5903,N_5853);
nand U6105 (N_6105,N_5860,N_5948);
nor U6106 (N_6106,N_5926,N_5993);
or U6107 (N_6107,N_5901,N_5831);
nor U6108 (N_6108,N_5940,N_5869);
or U6109 (N_6109,N_5881,N_5875);
or U6110 (N_6110,N_5848,N_5876);
or U6111 (N_6111,N_5931,N_5947);
or U6112 (N_6112,N_5933,N_5962);
and U6113 (N_6113,N_5906,N_5988);
or U6114 (N_6114,N_5853,N_5886);
and U6115 (N_6115,N_5879,N_5924);
or U6116 (N_6116,N_5809,N_5899);
and U6117 (N_6117,N_5991,N_5841);
or U6118 (N_6118,N_5817,N_5823);
nand U6119 (N_6119,N_5887,N_5964);
xnor U6120 (N_6120,N_5864,N_5980);
or U6121 (N_6121,N_5806,N_5987);
nor U6122 (N_6122,N_5865,N_5990);
or U6123 (N_6123,N_5900,N_5805);
nor U6124 (N_6124,N_5985,N_5965);
nor U6125 (N_6125,N_5953,N_5982);
nor U6126 (N_6126,N_5924,N_5892);
and U6127 (N_6127,N_5964,N_5907);
nand U6128 (N_6128,N_5883,N_5853);
or U6129 (N_6129,N_5816,N_5887);
nand U6130 (N_6130,N_5860,N_5822);
and U6131 (N_6131,N_5840,N_5880);
nor U6132 (N_6132,N_5896,N_5862);
nand U6133 (N_6133,N_5906,N_5807);
nand U6134 (N_6134,N_5944,N_5843);
nand U6135 (N_6135,N_5882,N_5922);
and U6136 (N_6136,N_5878,N_5966);
and U6137 (N_6137,N_5857,N_5807);
nor U6138 (N_6138,N_5915,N_5967);
xnor U6139 (N_6139,N_5934,N_5928);
and U6140 (N_6140,N_5867,N_5963);
nand U6141 (N_6141,N_5952,N_5843);
nand U6142 (N_6142,N_5964,N_5893);
or U6143 (N_6143,N_5835,N_5830);
xor U6144 (N_6144,N_5978,N_5905);
and U6145 (N_6145,N_5805,N_5892);
or U6146 (N_6146,N_5813,N_5976);
or U6147 (N_6147,N_5866,N_5974);
nor U6148 (N_6148,N_5984,N_5840);
or U6149 (N_6149,N_5873,N_5988);
and U6150 (N_6150,N_5821,N_5973);
nand U6151 (N_6151,N_5967,N_5985);
or U6152 (N_6152,N_5899,N_5939);
or U6153 (N_6153,N_5946,N_5891);
and U6154 (N_6154,N_5910,N_5842);
nand U6155 (N_6155,N_5990,N_5910);
or U6156 (N_6156,N_5933,N_5835);
and U6157 (N_6157,N_5865,N_5980);
nand U6158 (N_6158,N_5875,N_5810);
nand U6159 (N_6159,N_5898,N_5897);
xnor U6160 (N_6160,N_5867,N_5930);
nand U6161 (N_6161,N_5880,N_5860);
xnor U6162 (N_6162,N_5940,N_5882);
nor U6163 (N_6163,N_5910,N_5807);
or U6164 (N_6164,N_5817,N_5981);
and U6165 (N_6165,N_5824,N_5932);
or U6166 (N_6166,N_5804,N_5844);
nor U6167 (N_6167,N_5922,N_5927);
or U6168 (N_6168,N_5912,N_5922);
or U6169 (N_6169,N_5924,N_5917);
and U6170 (N_6170,N_5879,N_5830);
and U6171 (N_6171,N_5833,N_5801);
nand U6172 (N_6172,N_5937,N_5886);
nor U6173 (N_6173,N_5945,N_5901);
nor U6174 (N_6174,N_5976,N_5938);
nor U6175 (N_6175,N_5829,N_5873);
nand U6176 (N_6176,N_5897,N_5837);
or U6177 (N_6177,N_5840,N_5992);
nand U6178 (N_6178,N_5922,N_5854);
nor U6179 (N_6179,N_5990,N_5876);
xor U6180 (N_6180,N_5803,N_5814);
or U6181 (N_6181,N_5939,N_5833);
or U6182 (N_6182,N_5820,N_5818);
nor U6183 (N_6183,N_5864,N_5969);
nand U6184 (N_6184,N_5806,N_5995);
and U6185 (N_6185,N_5972,N_5810);
nand U6186 (N_6186,N_5896,N_5949);
or U6187 (N_6187,N_5979,N_5893);
nor U6188 (N_6188,N_5896,N_5893);
or U6189 (N_6189,N_5856,N_5925);
and U6190 (N_6190,N_5921,N_5941);
and U6191 (N_6191,N_5939,N_5821);
nor U6192 (N_6192,N_5913,N_5925);
or U6193 (N_6193,N_5807,N_5934);
or U6194 (N_6194,N_5884,N_5928);
and U6195 (N_6195,N_5886,N_5884);
and U6196 (N_6196,N_5836,N_5869);
xor U6197 (N_6197,N_5943,N_5995);
nand U6198 (N_6198,N_5937,N_5811);
nor U6199 (N_6199,N_5919,N_5894);
and U6200 (N_6200,N_6083,N_6025);
or U6201 (N_6201,N_6153,N_6197);
xor U6202 (N_6202,N_6099,N_6168);
and U6203 (N_6203,N_6034,N_6125);
and U6204 (N_6204,N_6106,N_6118);
nor U6205 (N_6205,N_6045,N_6170);
and U6206 (N_6206,N_6126,N_6088);
xnor U6207 (N_6207,N_6111,N_6130);
nand U6208 (N_6208,N_6049,N_6159);
or U6209 (N_6209,N_6132,N_6003);
nand U6210 (N_6210,N_6007,N_6072);
nor U6211 (N_6211,N_6199,N_6057);
nor U6212 (N_6212,N_6185,N_6009);
nand U6213 (N_6213,N_6037,N_6019);
and U6214 (N_6214,N_6195,N_6128);
or U6215 (N_6215,N_6137,N_6142);
nor U6216 (N_6216,N_6151,N_6114);
nor U6217 (N_6217,N_6056,N_6051);
or U6218 (N_6218,N_6038,N_6116);
nand U6219 (N_6219,N_6115,N_6157);
nor U6220 (N_6220,N_6066,N_6127);
xor U6221 (N_6221,N_6027,N_6053);
nand U6222 (N_6222,N_6140,N_6054);
or U6223 (N_6223,N_6131,N_6065);
nor U6224 (N_6224,N_6187,N_6188);
nor U6225 (N_6225,N_6107,N_6067);
nand U6226 (N_6226,N_6117,N_6184);
nor U6227 (N_6227,N_6143,N_6041);
or U6228 (N_6228,N_6108,N_6110);
xnor U6229 (N_6229,N_6050,N_6180);
or U6230 (N_6230,N_6136,N_6160);
and U6231 (N_6231,N_6103,N_6036);
or U6232 (N_6232,N_6102,N_6091);
and U6233 (N_6233,N_6084,N_6055);
or U6234 (N_6234,N_6120,N_6040);
and U6235 (N_6235,N_6169,N_6109);
nor U6236 (N_6236,N_6030,N_6146);
xnor U6237 (N_6237,N_6161,N_6058);
xor U6238 (N_6238,N_6135,N_6152);
or U6239 (N_6239,N_6074,N_6171);
nand U6240 (N_6240,N_6035,N_6062);
nor U6241 (N_6241,N_6133,N_6178);
xnor U6242 (N_6242,N_6089,N_6069);
and U6243 (N_6243,N_6121,N_6022);
and U6244 (N_6244,N_6061,N_6181);
nor U6245 (N_6245,N_6060,N_6174);
or U6246 (N_6246,N_6176,N_6182);
and U6247 (N_6247,N_6085,N_6064);
xnor U6248 (N_6248,N_6154,N_6194);
nor U6249 (N_6249,N_6001,N_6098);
and U6250 (N_6250,N_6101,N_6073);
and U6251 (N_6251,N_6097,N_6015);
and U6252 (N_6252,N_6092,N_6164);
and U6253 (N_6253,N_6129,N_6096);
or U6254 (N_6254,N_6113,N_6082);
nor U6255 (N_6255,N_6059,N_6005);
or U6256 (N_6256,N_6013,N_6147);
nor U6257 (N_6257,N_6112,N_6002);
nor U6258 (N_6258,N_6145,N_6190);
or U6259 (N_6259,N_6177,N_6076);
xor U6260 (N_6260,N_6141,N_6094);
nor U6261 (N_6261,N_6018,N_6078);
nand U6262 (N_6262,N_6077,N_6032);
nor U6263 (N_6263,N_6004,N_6079);
nor U6264 (N_6264,N_6029,N_6048);
and U6265 (N_6265,N_6063,N_6198);
or U6266 (N_6266,N_6031,N_6104);
and U6267 (N_6267,N_6021,N_6052);
nor U6268 (N_6268,N_6014,N_6043);
xnor U6269 (N_6269,N_6155,N_6046);
nor U6270 (N_6270,N_6012,N_6179);
nor U6271 (N_6271,N_6173,N_6162);
and U6272 (N_6272,N_6191,N_6039);
nand U6273 (N_6273,N_6163,N_6068);
nor U6274 (N_6274,N_6186,N_6086);
nand U6275 (N_6275,N_6175,N_6149);
and U6276 (N_6276,N_6010,N_6172);
nand U6277 (N_6277,N_6167,N_6070);
and U6278 (N_6278,N_6044,N_6134);
or U6279 (N_6279,N_6196,N_6148);
nor U6280 (N_6280,N_6008,N_6192);
or U6281 (N_6281,N_6122,N_6006);
nand U6282 (N_6282,N_6080,N_6087);
nand U6283 (N_6283,N_6033,N_6139);
nand U6284 (N_6284,N_6123,N_6189);
xor U6285 (N_6285,N_6119,N_6158);
and U6286 (N_6286,N_6028,N_6093);
or U6287 (N_6287,N_6144,N_6105);
nor U6288 (N_6288,N_6095,N_6017);
nand U6289 (N_6289,N_6024,N_6193);
nand U6290 (N_6290,N_6150,N_6075);
nor U6291 (N_6291,N_6081,N_6020);
nor U6292 (N_6292,N_6000,N_6026);
and U6293 (N_6293,N_6023,N_6071);
and U6294 (N_6294,N_6042,N_6183);
and U6295 (N_6295,N_6166,N_6156);
nor U6296 (N_6296,N_6100,N_6138);
xnor U6297 (N_6297,N_6016,N_6047);
and U6298 (N_6298,N_6090,N_6165);
nor U6299 (N_6299,N_6011,N_6124);
xnor U6300 (N_6300,N_6058,N_6108);
nor U6301 (N_6301,N_6101,N_6022);
nand U6302 (N_6302,N_6041,N_6020);
and U6303 (N_6303,N_6140,N_6130);
xnor U6304 (N_6304,N_6173,N_6023);
nand U6305 (N_6305,N_6126,N_6130);
or U6306 (N_6306,N_6108,N_6100);
or U6307 (N_6307,N_6040,N_6038);
and U6308 (N_6308,N_6180,N_6086);
and U6309 (N_6309,N_6105,N_6177);
and U6310 (N_6310,N_6008,N_6197);
xnor U6311 (N_6311,N_6076,N_6027);
and U6312 (N_6312,N_6107,N_6019);
nand U6313 (N_6313,N_6042,N_6150);
nor U6314 (N_6314,N_6061,N_6162);
and U6315 (N_6315,N_6032,N_6080);
or U6316 (N_6316,N_6173,N_6155);
nand U6317 (N_6317,N_6102,N_6142);
or U6318 (N_6318,N_6050,N_6195);
nor U6319 (N_6319,N_6183,N_6055);
nor U6320 (N_6320,N_6019,N_6002);
and U6321 (N_6321,N_6093,N_6097);
xor U6322 (N_6322,N_6153,N_6184);
and U6323 (N_6323,N_6015,N_6031);
nand U6324 (N_6324,N_6005,N_6117);
and U6325 (N_6325,N_6093,N_6155);
xor U6326 (N_6326,N_6034,N_6055);
nor U6327 (N_6327,N_6026,N_6169);
nor U6328 (N_6328,N_6199,N_6164);
nand U6329 (N_6329,N_6048,N_6109);
nor U6330 (N_6330,N_6105,N_6159);
nor U6331 (N_6331,N_6101,N_6091);
nor U6332 (N_6332,N_6198,N_6192);
and U6333 (N_6333,N_6170,N_6017);
or U6334 (N_6334,N_6157,N_6141);
and U6335 (N_6335,N_6057,N_6082);
nand U6336 (N_6336,N_6111,N_6141);
nor U6337 (N_6337,N_6024,N_6109);
nand U6338 (N_6338,N_6097,N_6199);
nor U6339 (N_6339,N_6058,N_6182);
nor U6340 (N_6340,N_6175,N_6152);
xnor U6341 (N_6341,N_6028,N_6082);
nand U6342 (N_6342,N_6072,N_6117);
xnor U6343 (N_6343,N_6188,N_6102);
nand U6344 (N_6344,N_6142,N_6074);
nor U6345 (N_6345,N_6022,N_6125);
or U6346 (N_6346,N_6117,N_6063);
nor U6347 (N_6347,N_6005,N_6112);
nand U6348 (N_6348,N_6111,N_6144);
nor U6349 (N_6349,N_6163,N_6102);
xnor U6350 (N_6350,N_6197,N_6012);
nor U6351 (N_6351,N_6145,N_6131);
and U6352 (N_6352,N_6057,N_6103);
xnor U6353 (N_6353,N_6196,N_6142);
or U6354 (N_6354,N_6079,N_6063);
nand U6355 (N_6355,N_6125,N_6156);
nand U6356 (N_6356,N_6049,N_6135);
nand U6357 (N_6357,N_6150,N_6082);
or U6358 (N_6358,N_6089,N_6019);
nand U6359 (N_6359,N_6021,N_6151);
and U6360 (N_6360,N_6194,N_6053);
and U6361 (N_6361,N_6188,N_6100);
nor U6362 (N_6362,N_6054,N_6064);
or U6363 (N_6363,N_6188,N_6148);
or U6364 (N_6364,N_6124,N_6067);
or U6365 (N_6365,N_6177,N_6154);
nor U6366 (N_6366,N_6069,N_6168);
or U6367 (N_6367,N_6006,N_6011);
nand U6368 (N_6368,N_6005,N_6167);
nor U6369 (N_6369,N_6090,N_6198);
and U6370 (N_6370,N_6135,N_6156);
nand U6371 (N_6371,N_6041,N_6169);
and U6372 (N_6372,N_6025,N_6081);
or U6373 (N_6373,N_6167,N_6145);
and U6374 (N_6374,N_6157,N_6147);
nor U6375 (N_6375,N_6171,N_6114);
nand U6376 (N_6376,N_6121,N_6062);
and U6377 (N_6377,N_6056,N_6064);
xor U6378 (N_6378,N_6008,N_6044);
and U6379 (N_6379,N_6173,N_6026);
and U6380 (N_6380,N_6144,N_6097);
and U6381 (N_6381,N_6175,N_6167);
nand U6382 (N_6382,N_6045,N_6080);
and U6383 (N_6383,N_6166,N_6062);
nand U6384 (N_6384,N_6115,N_6159);
and U6385 (N_6385,N_6012,N_6022);
or U6386 (N_6386,N_6089,N_6171);
xor U6387 (N_6387,N_6015,N_6108);
nand U6388 (N_6388,N_6192,N_6040);
or U6389 (N_6389,N_6161,N_6137);
nand U6390 (N_6390,N_6109,N_6063);
nor U6391 (N_6391,N_6181,N_6158);
or U6392 (N_6392,N_6175,N_6172);
xnor U6393 (N_6393,N_6193,N_6167);
nand U6394 (N_6394,N_6158,N_6195);
nand U6395 (N_6395,N_6157,N_6154);
xor U6396 (N_6396,N_6020,N_6065);
or U6397 (N_6397,N_6087,N_6058);
nand U6398 (N_6398,N_6105,N_6034);
nand U6399 (N_6399,N_6038,N_6146);
nand U6400 (N_6400,N_6256,N_6212);
or U6401 (N_6401,N_6340,N_6398);
nand U6402 (N_6402,N_6375,N_6261);
nand U6403 (N_6403,N_6293,N_6255);
or U6404 (N_6404,N_6393,N_6231);
nand U6405 (N_6405,N_6392,N_6358);
nor U6406 (N_6406,N_6205,N_6384);
and U6407 (N_6407,N_6371,N_6221);
or U6408 (N_6408,N_6292,N_6272);
nor U6409 (N_6409,N_6352,N_6342);
nor U6410 (N_6410,N_6209,N_6222);
or U6411 (N_6411,N_6319,N_6217);
and U6412 (N_6412,N_6381,N_6287);
or U6413 (N_6413,N_6328,N_6326);
or U6414 (N_6414,N_6244,N_6320);
xnor U6415 (N_6415,N_6330,N_6344);
or U6416 (N_6416,N_6203,N_6397);
nor U6417 (N_6417,N_6373,N_6368);
or U6418 (N_6418,N_6376,N_6369);
nand U6419 (N_6419,N_6236,N_6241);
nand U6420 (N_6420,N_6388,N_6289);
nor U6421 (N_6421,N_6211,N_6247);
xnor U6422 (N_6422,N_6239,N_6338);
and U6423 (N_6423,N_6207,N_6286);
nor U6424 (N_6424,N_6279,N_6232);
and U6425 (N_6425,N_6240,N_6225);
nand U6426 (N_6426,N_6308,N_6366);
and U6427 (N_6427,N_6389,N_6312);
or U6428 (N_6428,N_6306,N_6331);
xor U6429 (N_6429,N_6324,N_6285);
or U6430 (N_6430,N_6396,N_6283);
or U6431 (N_6431,N_6210,N_6313);
nor U6432 (N_6432,N_6380,N_6233);
and U6433 (N_6433,N_6359,N_6281);
and U6434 (N_6434,N_6206,N_6355);
nor U6435 (N_6435,N_6323,N_6335);
or U6436 (N_6436,N_6214,N_6298);
nor U6437 (N_6437,N_6327,N_6242);
nor U6438 (N_6438,N_6277,N_6235);
and U6439 (N_6439,N_6391,N_6341);
xnor U6440 (N_6440,N_6300,N_6284);
or U6441 (N_6441,N_6374,N_6248);
nor U6442 (N_6442,N_6337,N_6317);
nor U6443 (N_6443,N_6297,N_6224);
and U6444 (N_6444,N_6386,N_6260);
and U6445 (N_6445,N_6234,N_6223);
nor U6446 (N_6446,N_6316,N_6302);
or U6447 (N_6447,N_6215,N_6348);
or U6448 (N_6448,N_6349,N_6267);
and U6449 (N_6449,N_6385,N_6201);
nor U6450 (N_6450,N_6322,N_6254);
and U6451 (N_6451,N_6325,N_6332);
and U6452 (N_6452,N_6357,N_6294);
nor U6453 (N_6453,N_6238,N_6315);
nor U6454 (N_6454,N_6343,N_6258);
or U6455 (N_6455,N_6301,N_6365);
or U6456 (N_6456,N_6257,N_6246);
nor U6457 (N_6457,N_6216,N_6367);
nor U6458 (N_6458,N_6290,N_6226);
nor U6459 (N_6459,N_6351,N_6307);
and U6460 (N_6460,N_6364,N_6311);
nand U6461 (N_6461,N_6299,N_6346);
nor U6462 (N_6462,N_6399,N_6360);
and U6463 (N_6463,N_6345,N_6382);
nand U6464 (N_6464,N_6268,N_6252);
and U6465 (N_6465,N_6249,N_6394);
xnor U6466 (N_6466,N_6270,N_6304);
nor U6467 (N_6467,N_6303,N_6329);
and U6468 (N_6468,N_6245,N_6347);
or U6469 (N_6469,N_6339,N_6377);
nor U6470 (N_6470,N_6280,N_6295);
or U6471 (N_6471,N_6305,N_6219);
or U6472 (N_6472,N_6229,N_6333);
or U6473 (N_6473,N_6314,N_6291);
and U6474 (N_6474,N_6200,N_6353);
and U6475 (N_6475,N_6288,N_6309);
nand U6476 (N_6476,N_6227,N_6218);
and U6477 (N_6477,N_6237,N_6263);
nand U6478 (N_6478,N_6276,N_6273);
nor U6479 (N_6479,N_6269,N_6213);
nor U6480 (N_6480,N_6265,N_6379);
and U6481 (N_6481,N_6253,N_6310);
and U6482 (N_6482,N_6208,N_6250);
nor U6483 (N_6483,N_6204,N_6266);
nor U6484 (N_6484,N_6336,N_6356);
and U6485 (N_6485,N_6243,N_6259);
and U6486 (N_6486,N_6282,N_6395);
nand U6487 (N_6487,N_6251,N_6354);
or U6488 (N_6488,N_6321,N_6296);
nor U6489 (N_6489,N_6275,N_6278);
and U6490 (N_6490,N_6378,N_6318);
and U6491 (N_6491,N_6264,N_6271);
xor U6492 (N_6492,N_6383,N_6362);
and U6493 (N_6493,N_6372,N_6361);
nand U6494 (N_6494,N_6350,N_6334);
and U6495 (N_6495,N_6363,N_6370);
xnor U6496 (N_6496,N_6387,N_6220);
or U6497 (N_6497,N_6262,N_6202);
nor U6498 (N_6498,N_6228,N_6230);
nor U6499 (N_6499,N_6274,N_6390);
xnor U6500 (N_6500,N_6228,N_6333);
xor U6501 (N_6501,N_6229,N_6319);
nand U6502 (N_6502,N_6266,N_6378);
nor U6503 (N_6503,N_6255,N_6397);
and U6504 (N_6504,N_6206,N_6216);
nand U6505 (N_6505,N_6273,N_6383);
nand U6506 (N_6506,N_6258,N_6296);
nand U6507 (N_6507,N_6210,N_6318);
xor U6508 (N_6508,N_6206,N_6373);
xor U6509 (N_6509,N_6324,N_6286);
nand U6510 (N_6510,N_6307,N_6201);
nand U6511 (N_6511,N_6202,N_6337);
nand U6512 (N_6512,N_6257,N_6363);
nor U6513 (N_6513,N_6380,N_6214);
nor U6514 (N_6514,N_6237,N_6213);
and U6515 (N_6515,N_6202,N_6275);
nor U6516 (N_6516,N_6357,N_6232);
nand U6517 (N_6517,N_6241,N_6262);
nand U6518 (N_6518,N_6234,N_6378);
and U6519 (N_6519,N_6318,N_6367);
or U6520 (N_6520,N_6299,N_6336);
or U6521 (N_6521,N_6238,N_6205);
and U6522 (N_6522,N_6291,N_6210);
and U6523 (N_6523,N_6260,N_6324);
nor U6524 (N_6524,N_6275,N_6341);
nor U6525 (N_6525,N_6230,N_6368);
nor U6526 (N_6526,N_6217,N_6345);
or U6527 (N_6527,N_6364,N_6323);
and U6528 (N_6528,N_6298,N_6348);
nor U6529 (N_6529,N_6212,N_6213);
or U6530 (N_6530,N_6276,N_6235);
and U6531 (N_6531,N_6257,N_6347);
or U6532 (N_6532,N_6222,N_6389);
nor U6533 (N_6533,N_6346,N_6394);
nand U6534 (N_6534,N_6342,N_6319);
or U6535 (N_6535,N_6239,N_6233);
and U6536 (N_6536,N_6355,N_6280);
nor U6537 (N_6537,N_6223,N_6200);
or U6538 (N_6538,N_6281,N_6202);
nor U6539 (N_6539,N_6359,N_6224);
or U6540 (N_6540,N_6226,N_6221);
and U6541 (N_6541,N_6305,N_6215);
nor U6542 (N_6542,N_6386,N_6299);
or U6543 (N_6543,N_6288,N_6395);
nand U6544 (N_6544,N_6347,N_6365);
nand U6545 (N_6545,N_6289,N_6359);
nor U6546 (N_6546,N_6382,N_6210);
and U6547 (N_6547,N_6263,N_6323);
nand U6548 (N_6548,N_6361,N_6305);
nor U6549 (N_6549,N_6297,N_6258);
and U6550 (N_6550,N_6245,N_6391);
nor U6551 (N_6551,N_6311,N_6238);
nand U6552 (N_6552,N_6381,N_6356);
nand U6553 (N_6553,N_6321,N_6225);
nor U6554 (N_6554,N_6305,N_6292);
nor U6555 (N_6555,N_6248,N_6345);
and U6556 (N_6556,N_6364,N_6211);
nand U6557 (N_6557,N_6223,N_6267);
or U6558 (N_6558,N_6333,N_6219);
or U6559 (N_6559,N_6360,N_6259);
nor U6560 (N_6560,N_6313,N_6255);
and U6561 (N_6561,N_6207,N_6387);
nor U6562 (N_6562,N_6325,N_6357);
and U6563 (N_6563,N_6203,N_6214);
and U6564 (N_6564,N_6375,N_6354);
and U6565 (N_6565,N_6363,N_6344);
and U6566 (N_6566,N_6351,N_6263);
or U6567 (N_6567,N_6232,N_6272);
nor U6568 (N_6568,N_6386,N_6245);
nor U6569 (N_6569,N_6242,N_6285);
xor U6570 (N_6570,N_6249,N_6354);
xnor U6571 (N_6571,N_6301,N_6298);
and U6572 (N_6572,N_6214,N_6307);
or U6573 (N_6573,N_6371,N_6260);
nand U6574 (N_6574,N_6306,N_6271);
nand U6575 (N_6575,N_6291,N_6268);
and U6576 (N_6576,N_6321,N_6342);
nand U6577 (N_6577,N_6223,N_6247);
nand U6578 (N_6578,N_6368,N_6393);
xor U6579 (N_6579,N_6332,N_6340);
nand U6580 (N_6580,N_6306,N_6384);
and U6581 (N_6581,N_6386,N_6365);
nand U6582 (N_6582,N_6351,N_6244);
nand U6583 (N_6583,N_6327,N_6348);
nand U6584 (N_6584,N_6264,N_6218);
nor U6585 (N_6585,N_6396,N_6373);
and U6586 (N_6586,N_6223,N_6208);
nor U6587 (N_6587,N_6340,N_6371);
nor U6588 (N_6588,N_6316,N_6276);
nand U6589 (N_6589,N_6208,N_6292);
xnor U6590 (N_6590,N_6324,N_6222);
and U6591 (N_6591,N_6314,N_6251);
nand U6592 (N_6592,N_6377,N_6396);
nand U6593 (N_6593,N_6215,N_6293);
or U6594 (N_6594,N_6295,N_6230);
and U6595 (N_6595,N_6319,N_6324);
xor U6596 (N_6596,N_6281,N_6249);
or U6597 (N_6597,N_6399,N_6208);
or U6598 (N_6598,N_6357,N_6344);
nand U6599 (N_6599,N_6204,N_6290);
and U6600 (N_6600,N_6528,N_6547);
nand U6601 (N_6601,N_6478,N_6503);
nor U6602 (N_6602,N_6562,N_6495);
nor U6603 (N_6603,N_6443,N_6542);
and U6604 (N_6604,N_6446,N_6577);
nor U6605 (N_6605,N_6551,N_6406);
nand U6606 (N_6606,N_6440,N_6566);
and U6607 (N_6607,N_6438,N_6582);
nor U6608 (N_6608,N_6593,N_6554);
and U6609 (N_6609,N_6448,N_6525);
and U6610 (N_6610,N_6511,N_6591);
and U6611 (N_6611,N_6480,N_6460);
nand U6612 (N_6612,N_6471,N_6423);
or U6613 (N_6613,N_6453,N_6450);
xnor U6614 (N_6614,N_6517,N_6524);
nand U6615 (N_6615,N_6575,N_6428);
nor U6616 (N_6616,N_6421,N_6437);
nor U6617 (N_6617,N_6579,N_6498);
nand U6618 (N_6618,N_6584,N_6518);
or U6619 (N_6619,N_6516,N_6484);
or U6620 (N_6620,N_6519,N_6409);
nor U6621 (N_6621,N_6514,N_6489);
or U6622 (N_6622,N_6549,N_6580);
nor U6623 (N_6623,N_6539,N_6544);
xor U6624 (N_6624,N_6465,N_6429);
nand U6625 (N_6625,N_6550,N_6581);
or U6626 (N_6626,N_6463,N_6491);
nand U6627 (N_6627,N_6537,N_6400);
nand U6628 (N_6628,N_6492,N_6538);
nand U6629 (N_6629,N_6472,N_6499);
or U6630 (N_6630,N_6559,N_6595);
and U6631 (N_6631,N_6455,N_6546);
and U6632 (N_6632,N_6413,N_6599);
and U6633 (N_6633,N_6500,N_6456);
xor U6634 (N_6634,N_6597,N_6494);
or U6635 (N_6635,N_6441,N_6535);
nand U6636 (N_6636,N_6442,N_6435);
and U6637 (N_6637,N_6447,N_6572);
or U6638 (N_6638,N_6475,N_6523);
and U6639 (N_6639,N_6416,N_6504);
nand U6640 (N_6640,N_6461,N_6462);
xnor U6641 (N_6641,N_6508,N_6563);
nor U6642 (N_6642,N_6553,N_6405);
or U6643 (N_6643,N_6587,N_6401);
nand U6644 (N_6644,N_6417,N_6481);
nand U6645 (N_6645,N_6585,N_6430);
or U6646 (N_6646,N_6479,N_6596);
nand U6647 (N_6647,N_6513,N_6592);
and U6648 (N_6648,N_6526,N_6564);
nor U6649 (N_6649,N_6439,N_6473);
nand U6650 (N_6650,N_6436,N_6434);
nor U6651 (N_6651,N_6502,N_6474);
or U6652 (N_6652,N_6578,N_6427);
nor U6653 (N_6653,N_6541,N_6402);
and U6654 (N_6654,N_6557,N_6509);
nand U6655 (N_6655,N_6565,N_6458);
nor U6656 (N_6656,N_6555,N_6433);
nand U6657 (N_6657,N_6467,N_6505);
and U6658 (N_6658,N_6573,N_6588);
or U6659 (N_6659,N_6403,N_6420);
and U6660 (N_6660,N_6527,N_6533);
and U6661 (N_6661,N_6510,N_6457);
nor U6662 (N_6662,N_6431,N_6497);
or U6663 (N_6663,N_6530,N_6444);
nand U6664 (N_6664,N_6422,N_6536);
nand U6665 (N_6665,N_6445,N_6469);
xnor U6666 (N_6666,N_6449,N_6486);
or U6667 (N_6667,N_6468,N_6419);
or U6668 (N_6668,N_6432,N_6490);
nand U6669 (N_6669,N_6410,N_6548);
nand U6670 (N_6670,N_6561,N_6568);
nand U6671 (N_6671,N_6560,N_6496);
or U6672 (N_6672,N_6594,N_6451);
nor U6673 (N_6673,N_6532,N_6545);
and U6674 (N_6674,N_6506,N_6408);
or U6675 (N_6675,N_6493,N_6586);
and U6676 (N_6676,N_6570,N_6464);
or U6677 (N_6677,N_6576,N_6520);
nor U6678 (N_6678,N_6534,N_6482);
and U6679 (N_6679,N_6543,N_6529);
and U6680 (N_6680,N_6507,N_6558);
nand U6681 (N_6681,N_6590,N_6501);
and U6682 (N_6682,N_6552,N_6598);
and U6683 (N_6683,N_6407,N_6412);
and U6684 (N_6684,N_6415,N_6418);
nor U6685 (N_6685,N_6531,N_6404);
nor U6686 (N_6686,N_6512,N_6574);
or U6687 (N_6687,N_6425,N_6426);
or U6688 (N_6688,N_6454,N_6411);
and U6689 (N_6689,N_6567,N_6569);
and U6690 (N_6690,N_6414,N_6556);
and U6691 (N_6691,N_6522,N_6540);
nor U6692 (N_6692,N_6476,N_6424);
or U6693 (N_6693,N_6515,N_6452);
or U6694 (N_6694,N_6487,N_6589);
nor U6695 (N_6695,N_6521,N_6466);
or U6696 (N_6696,N_6583,N_6470);
nand U6697 (N_6697,N_6483,N_6477);
xor U6698 (N_6698,N_6571,N_6488);
xor U6699 (N_6699,N_6459,N_6485);
xnor U6700 (N_6700,N_6550,N_6506);
xnor U6701 (N_6701,N_6557,N_6598);
or U6702 (N_6702,N_6595,N_6510);
or U6703 (N_6703,N_6545,N_6582);
nand U6704 (N_6704,N_6542,N_6441);
xor U6705 (N_6705,N_6485,N_6533);
or U6706 (N_6706,N_6412,N_6414);
nand U6707 (N_6707,N_6430,N_6501);
or U6708 (N_6708,N_6400,N_6492);
nor U6709 (N_6709,N_6513,N_6435);
or U6710 (N_6710,N_6404,N_6570);
and U6711 (N_6711,N_6433,N_6584);
nand U6712 (N_6712,N_6589,N_6505);
and U6713 (N_6713,N_6502,N_6522);
nand U6714 (N_6714,N_6597,N_6563);
and U6715 (N_6715,N_6459,N_6405);
nor U6716 (N_6716,N_6581,N_6504);
and U6717 (N_6717,N_6574,N_6455);
or U6718 (N_6718,N_6431,N_6571);
nand U6719 (N_6719,N_6429,N_6552);
or U6720 (N_6720,N_6450,N_6413);
nand U6721 (N_6721,N_6596,N_6476);
and U6722 (N_6722,N_6402,N_6594);
or U6723 (N_6723,N_6506,N_6569);
nor U6724 (N_6724,N_6474,N_6436);
nand U6725 (N_6725,N_6513,N_6400);
or U6726 (N_6726,N_6536,N_6449);
or U6727 (N_6727,N_6496,N_6579);
or U6728 (N_6728,N_6400,N_6427);
nand U6729 (N_6729,N_6428,N_6557);
xnor U6730 (N_6730,N_6583,N_6473);
nand U6731 (N_6731,N_6513,N_6468);
and U6732 (N_6732,N_6594,N_6523);
and U6733 (N_6733,N_6597,N_6408);
nor U6734 (N_6734,N_6499,N_6502);
or U6735 (N_6735,N_6509,N_6524);
and U6736 (N_6736,N_6484,N_6528);
and U6737 (N_6737,N_6488,N_6570);
nor U6738 (N_6738,N_6401,N_6468);
xor U6739 (N_6739,N_6447,N_6471);
or U6740 (N_6740,N_6432,N_6503);
or U6741 (N_6741,N_6419,N_6444);
nand U6742 (N_6742,N_6482,N_6462);
and U6743 (N_6743,N_6532,N_6430);
nand U6744 (N_6744,N_6474,N_6452);
xnor U6745 (N_6745,N_6400,N_6466);
or U6746 (N_6746,N_6493,N_6551);
and U6747 (N_6747,N_6458,N_6411);
or U6748 (N_6748,N_6581,N_6450);
nand U6749 (N_6749,N_6448,N_6526);
nand U6750 (N_6750,N_6478,N_6593);
and U6751 (N_6751,N_6548,N_6553);
nor U6752 (N_6752,N_6486,N_6529);
or U6753 (N_6753,N_6529,N_6464);
and U6754 (N_6754,N_6419,N_6520);
or U6755 (N_6755,N_6518,N_6488);
nand U6756 (N_6756,N_6582,N_6479);
nand U6757 (N_6757,N_6424,N_6436);
or U6758 (N_6758,N_6518,N_6495);
or U6759 (N_6759,N_6469,N_6558);
nor U6760 (N_6760,N_6426,N_6421);
nand U6761 (N_6761,N_6458,N_6477);
xor U6762 (N_6762,N_6586,N_6558);
nor U6763 (N_6763,N_6444,N_6429);
nand U6764 (N_6764,N_6529,N_6560);
or U6765 (N_6765,N_6489,N_6423);
and U6766 (N_6766,N_6570,N_6427);
xor U6767 (N_6767,N_6411,N_6433);
xor U6768 (N_6768,N_6491,N_6560);
and U6769 (N_6769,N_6478,N_6434);
nand U6770 (N_6770,N_6493,N_6429);
nor U6771 (N_6771,N_6508,N_6443);
nand U6772 (N_6772,N_6444,N_6541);
and U6773 (N_6773,N_6497,N_6452);
and U6774 (N_6774,N_6467,N_6559);
or U6775 (N_6775,N_6574,N_6416);
xor U6776 (N_6776,N_6410,N_6494);
xor U6777 (N_6777,N_6424,N_6572);
and U6778 (N_6778,N_6537,N_6477);
xnor U6779 (N_6779,N_6449,N_6413);
nand U6780 (N_6780,N_6515,N_6402);
and U6781 (N_6781,N_6597,N_6546);
xor U6782 (N_6782,N_6565,N_6483);
nor U6783 (N_6783,N_6574,N_6499);
nor U6784 (N_6784,N_6411,N_6529);
nor U6785 (N_6785,N_6536,N_6595);
nand U6786 (N_6786,N_6433,N_6456);
xnor U6787 (N_6787,N_6497,N_6460);
and U6788 (N_6788,N_6585,N_6567);
nand U6789 (N_6789,N_6505,N_6424);
or U6790 (N_6790,N_6517,N_6557);
nor U6791 (N_6791,N_6500,N_6535);
or U6792 (N_6792,N_6580,N_6515);
nor U6793 (N_6793,N_6455,N_6498);
nand U6794 (N_6794,N_6512,N_6515);
nor U6795 (N_6795,N_6488,N_6526);
and U6796 (N_6796,N_6487,N_6465);
nand U6797 (N_6797,N_6531,N_6468);
nor U6798 (N_6798,N_6495,N_6416);
nand U6799 (N_6799,N_6500,N_6568);
nand U6800 (N_6800,N_6781,N_6728);
nand U6801 (N_6801,N_6632,N_6670);
and U6802 (N_6802,N_6611,N_6714);
nand U6803 (N_6803,N_6796,N_6673);
nor U6804 (N_6804,N_6751,N_6686);
or U6805 (N_6805,N_6715,N_6706);
xnor U6806 (N_6806,N_6660,N_6766);
or U6807 (N_6807,N_6687,N_6691);
nor U6808 (N_6808,N_6666,N_6791);
nor U6809 (N_6809,N_6759,N_6635);
xor U6810 (N_6810,N_6616,N_6733);
and U6811 (N_6811,N_6737,N_6639);
nor U6812 (N_6812,N_6647,N_6762);
nand U6813 (N_6813,N_6790,N_6665);
nor U6814 (N_6814,N_6780,N_6768);
or U6815 (N_6815,N_6757,N_6717);
nor U6816 (N_6816,N_6705,N_6797);
nor U6817 (N_6817,N_6702,N_6697);
or U6818 (N_6818,N_6692,N_6655);
and U6819 (N_6819,N_6723,N_6689);
nor U6820 (N_6820,N_6718,N_6710);
and U6821 (N_6821,N_6649,N_6618);
xnor U6822 (N_6822,N_6645,N_6664);
and U6823 (N_6823,N_6708,N_6600);
xnor U6824 (N_6824,N_6617,N_6661);
and U6825 (N_6825,N_6669,N_6631);
or U6826 (N_6826,N_6739,N_6799);
nand U6827 (N_6827,N_6761,N_6668);
or U6828 (N_6828,N_6711,N_6651);
or U6829 (N_6829,N_6758,N_6746);
nor U6830 (N_6830,N_6760,N_6671);
nor U6831 (N_6831,N_6638,N_6778);
or U6832 (N_6832,N_6676,N_6755);
and U6833 (N_6833,N_6628,N_6732);
and U6834 (N_6834,N_6633,N_6750);
or U6835 (N_6835,N_6725,N_6741);
and U6836 (N_6836,N_6744,N_6672);
and U6837 (N_6837,N_6641,N_6623);
and U6838 (N_6838,N_6730,N_6696);
nor U6839 (N_6839,N_6636,N_6688);
nor U6840 (N_6840,N_6629,N_6716);
nand U6841 (N_6841,N_6704,N_6784);
nand U6842 (N_6842,N_6776,N_6612);
or U6843 (N_6843,N_6677,N_6650);
nor U6844 (N_6844,N_6674,N_6783);
nand U6845 (N_6845,N_6752,N_6622);
or U6846 (N_6846,N_6720,N_6734);
xor U6847 (N_6847,N_6662,N_6606);
or U6848 (N_6848,N_6727,N_6603);
nand U6849 (N_6849,N_6625,N_6738);
xor U6850 (N_6850,N_6608,N_6743);
nand U6851 (N_6851,N_6794,N_6788);
and U6852 (N_6852,N_6634,N_6642);
nand U6853 (N_6853,N_6694,N_6724);
xor U6854 (N_6854,N_6756,N_6602);
and U6855 (N_6855,N_6747,N_6729);
or U6856 (N_6856,N_6604,N_6767);
nand U6857 (N_6857,N_6626,N_6749);
nand U6858 (N_6858,N_6701,N_6624);
nand U6859 (N_6859,N_6695,N_6745);
and U6860 (N_6860,N_6748,N_6798);
nor U6861 (N_6861,N_6630,N_6698);
or U6862 (N_6862,N_6786,N_6787);
nor U6863 (N_6863,N_6709,N_6726);
and U6864 (N_6864,N_6653,N_6680);
nand U6865 (N_6865,N_6646,N_6699);
nor U6866 (N_6866,N_6773,N_6679);
nand U6867 (N_6867,N_6782,N_6619);
nand U6868 (N_6868,N_6735,N_6621);
xor U6869 (N_6869,N_6667,N_6722);
or U6870 (N_6870,N_6644,N_6678);
nand U6871 (N_6871,N_6610,N_6683);
nand U6872 (N_6872,N_6792,N_6620);
nor U6873 (N_6873,N_6763,N_6659);
or U6874 (N_6874,N_6615,N_6656);
nor U6875 (N_6875,N_6795,N_6765);
nand U6876 (N_6876,N_6736,N_6627);
nor U6877 (N_6877,N_6713,N_6789);
nor U6878 (N_6878,N_6605,N_6640);
or U6879 (N_6879,N_6643,N_6770);
and U6880 (N_6880,N_6607,N_6682);
nand U6881 (N_6881,N_6775,N_6779);
nand U6882 (N_6882,N_6764,N_6652);
and U6883 (N_6883,N_6654,N_6707);
nand U6884 (N_6884,N_6681,N_6648);
or U6885 (N_6885,N_6769,N_6793);
nand U6886 (N_6886,N_6675,N_6740);
nor U6887 (N_6887,N_6693,N_6684);
nand U6888 (N_6888,N_6614,N_6772);
and U6889 (N_6889,N_6742,N_6685);
xnor U6890 (N_6890,N_6658,N_6721);
xor U6891 (N_6891,N_6771,N_6712);
nand U6892 (N_6892,N_6609,N_6785);
nor U6893 (N_6893,N_6663,N_6601);
nand U6894 (N_6894,N_6731,N_6719);
nor U6895 (N_6895,N_6754,N_6690);
nand U6896 (N_6896,N_6777,N_6753);
and U6897 (N_6897,N_6613,N_6774);
or U6898 (N_6898,N_6700,N_6657);
xor U6899 (N_6899,N_6637,N_6703);
or U6900 (N_6900,N_6712,N_6724);
nor U6901 (N_6901,N_6747,N_6625);
or U6902 (N_6902,N_6771,N_6747);
nand U6903 (N_6903,N_6673,N_6604);
or U6904 (N_6904,N_6722,N_6666);
nor U6905 (N_6905,N_6741,N_6654);
or U6906 (N_6906,N_6637,N_6789);
nand U6907 (N_6907,N_6695,N_6779);
and U6908 (N_6908,N_6740,N_6695);
xor U6909 (N_6909,N_6758,N_6744);
and U6910 (N_6910,N_6686,N_6620);
nor U6911 (N_6911,N_6626,N_6615);
nand U6912 (N_6912,N_6766,N_6602);
and U6913 (N_6913,N_6651,N_6799);
nor U6914 (N_6914,N_6644,N_6763);
nor U6915 (N_6915,N_6619,N_6738);
or U6916 (N_6916,N_6781,N_6685);
and U6917 (N_6917,N_6680,N_6700);
or U6918 (N_6918,N_6611,N_6743);
or U6919 (N_6919,N_6630,N_6703);
and U6920 (N_6920,N_6754,N_6607);
xnor U6921 (N_6921,N_6716,N_6646);
nand U6922 (N_6922,N_6719,N_6686);
or U6923 (N_6923,N_6691,N_6669);
and U6924 (N_6924,N_6692,N_6758);
nand U6925 (N_6925,N_6696,N_6727);
or U6926 (N_6926,N_6681,N_6630);
xor U6927 (N_6927,N_6610,N_6764);
or U6928 (N_6928,N_6774,N_6695);
nor U6929 (N_6929,N_6785,N_6758);
and U6930 (N_6930,N_6746,N_6668);
and U6931 (N_6931,N_6764,N_6725);
nand U6932 (N_6932,N_6750,N_6614);
nor U6933 (N_6933,N_6631,N_6620);
nand U6934 (N_6934,N_6677,N_6672);
or U6935 (N_6935,N_6689,N_6791);
or U6936 (N_6936,N_6781,N_6751);
nor U6937 (N_6937,N_6685,N_6704);
and U6938 (N_6938,N_6697,N_6653);
xnor U6939 (N_6939,N_6785,N_6678);
nor U6940 (N_6940,N_6668,N_6661);
or U6941 (N_6941,N_6606,N_6799);
and U6942 (N_6942,N_6668,N_6606);
nor U6943 (N_6943,N_6624,N_6759);
and U6944 (N_6944,N_6796,N_6710);
and U6945 (N_6945,N_6643,N_6628);
nor U6946 (N_6946,N_6655,N_6772);
nor U6947 (N_6947,N_6771,N_6627);
and U6948 (N_6948,N_6678,N_6649);
xor U6949 (N_6949,N_6616,N_6694);
nand U6950 (N_6950,N_6608,N_6689);
nand U6951 (N_6951,N_6790,N_6723);
nand U6952 (N_6952,N_6664,N_6610);
or U6953 (N_6953,N_6780,N_6613);
nand U6954 (N_6954,N_6680,N_6635);
nand U6955 (N_6955,N_6718,N_6631);
nand U6956 (N_6956,N_6784,N_6759);
or U6957 (N_6957,N_6725,N_6679);
or U6958 (N_6958,N_6765,N_6732);
nor U6959 (N_6959,N_6613,N_6756);
and U6960 (N_6960,N_6726,N_6782);
nand U6961 (N_6961,N_6695,N_6768);
nor U6962 (N_6962,N_6789,N_6656);
nor U6963 (N_6963,N_6738,N_6764);
and U6964 (N_6964,N_6705,N_6716);
xnor U6965 (N_6965,N_6612,N_6728);
nand U6966 (N_6966,N_6642,N_6697);
nor U6967 (N_6967,N_6635,N_6689);
nand U6968 (N_6968,N_6744,N_6718);
nor U6969 (N_6969,N_6680,N_6641);
or U6970 (N_6970,N_6777,N_6645);
and U6971 (N_6971,N_6682,N_6783);
nor U6972 (N_6972,N_6708,N_6707);
or U6973 (N_6973,N_6735,N_6723);
nand U6974 (N_6974,N_6660,N_6645);
nor U6975 (N_6975,N_6798,N_6778);
or U6976 (N_6976,N_6769,N_6729);
or U6977 (N_6977,N_6666,N_6751);
or U6978 (N_6978,N_6664,N_6642);
and U6979 (N_6979,N_6689,N_6749);
xor U6980 (N_6980,N_6703,N_6737);
nand U6981 (N_6981,N_6650,N_6787);
nand U6982 (N_6982,N_6693,N_6644);
and U6983 (N_6983,N_6735,N_6685);
nor U6984 (N_6984,N_6630,N_6676);
nor U6985 (N_6985,N_6684,N_6774);
or U6986 (N_6986,N_6628,N_6695);
or U6987 (N_6987,N_6742,N_6735);
nand U6988 (N_6988,N_6637,N_6790);
nand U6989 (N_6989,N_6649,N_6635);
nor U6990 (N_6990,N_6758,N_6691);
nor U6991 (N_6991,N_6720,N_6719);
or U6992 (N_6992,N_6738,N_6792);
xor U6993 (N_6993,N_6669,N_6677);
and U6994 (N_6994,N_6795,N_6603);
and U6995 (N_6995,N_6715,N_6680);
and U6996 (N_6996,N_6672,N_6662);
or U6997 (N_6997,N_6696,N_6685);
nand U6998 (N_6998,N_6708,N_6793);
or U6999 (N_6999,N_6748,N_6653);
or U7000 (N_7000,N_6801,N_6991);
nor U7001 (N_7001,N_6805,N_6917);
and U7002 (N_7002,N_6838,N_6987);
nor U7003 (N_7003,N_6944,N_6909);
and U7004 (N_7004,N_6979,N_6880);
nor U7005 (N_7005,N_6901,N_6952);
nor U7006 (N_7006,N_6886,N_6922);
nand U7007 (N_7007,N_6861,N_6937);
xnor U7008 (N_7008,N_6932,N_6845);
nand U7009 (N_7009,N_6832,N_6808);
or U7010 (N_7010,N_6940,N_6936);
and U7011 (N_7011,N_6891,N_6853);
nand U7012 (N_7012,N_6864,N_6883);
nand U7013 (N_7013,N_6918,N_6995);
nor U7014 (N_7014,N_6807,N_6975);
or U7015 (N_7015,N_6976,N_6914);
nor U7016 (N_7016,N_6986,N_6850);
nor U7017 (N_7017,N_6800,N_6950);
xnor U7018 (N_7018,N_6802,N_6817);
and U7019 (N_7019,N_6806,N_6980);
and U7020 (N_7020,N_6865,N_6847);
nor U7021 (N_7021,N_6958,N_6997);
or U7022 (N_7022,N_6825,N_6947);
or U7023 (N_7023,N_6935,N_6905);
xor U7024 (N_7024,N_6870,N_6829);
or U7025 (N_7025,N_6814,N_6874);
or U7026 (N_7026,N_6894,N_6959);
and U7027 (N_7027,N_6966,N_6961);
or U7028 (N_7028,N_6854,N_6994);
nor U7029 (N_7029,N_6823,N_6942);
or U7030 (N_7030,N_6971,N_6873);
xnor U7031 (N_7031,N_6820,N_6809);
and U7032 (N_7032,N_6871,N_6907);
and U7033 (N_7033,N_6928,N_6960);
nor U7034 (N_7034,N_6813,N_6811);
and U7035 (N_7035,N_6903,N_6925);
nor U7036 (N_7036,N_6924,N_6858);
nor U7037 (N_7037,N_6892,N_6983);
or U7038 (N_7038,N_6985,N_6893);
or U7039 (N_7039,N_6876,N_6819);
nor U7040 (N_7040,N_6996,N_6881);
or U7041 (N_7041,N_6890,N_6951);
nand U7042 (N_7042,N_6954,N_6906);
or U7043 (N_7043,N_6849,N_6842);
xnor U7044 (N_7044,N_6869,N_6929);
or U7045 (N_7045,N_6988,N_6839);
xor U7046 (N_7046,N_6884,N_6982);
nand U7047 (N_7047,N_6939,N_6934);
nand U7048 (N_7048,N_6834,N_6859);
nor U7049 (N_7049,N_6810,N_6855);
xnor U7050 (N_7050,N_6913,N_6945);
nor U7051 (N_7051,N_6836,N_6999);
or U7052 (N_7052,N_6815,N_6931);
nand U7053 (N_7053,N_6846,N_6878);
nand U7054 (N_7054,N_6993,N_6948);
xor U7055 (N_7055,N_6956,N_6866);
nand U7056 (N_7056,N_6827,N_6927);
and U7057 (N_7057,N_6989,N_6848);
nand U7058 (N_7058,N_6926,N_6856);
and U7059 (N_7059,N_6998,N_6803);
or U7060 (N_7060,N_6885,N_6888);
and U7061 (N_7061,N_6974,N_6860);
nand U7062 (N_7062,N_6930,N_6938);
or U7063 (N_7063,N_6816,N_6818);
nor U7064 (N_7064,N_6933,N_6946);
nor U7065 (N_7065,N_6835,N_6920);
nor U7066 (N_7066,N_6978,N_6923);
nor U7067 (N_7067,N_6899,N_6862);
nor U7068 (N_7068,N_6882,N_6900);
and U7069 (N_7069,N_6868,N_6972);
nor U7070 (N_7070,N_6898,N_6812);
or U7071 (N_7071,N_6904,N_6828);
xor U7072 (N_7072,N_6841,N_6826);
or U7073 (N_7073,N_6895,N_6837);
and U7074 (N_7074,N_6857,N_6912);
nor U7075 (N_7075,N_6964,N_6970);
or U7076 (N_7076,N_6897,N_6887);
or U7077 (N_7077,N_6910,N_6969);
nor U7078 (N_7078,N_6822,N_6915);
or U7079 (N_7079,N_6973,N_6968);
and U7080 (N_7080,N_6911,N_6977);
xor U7081 (N_7081,N_6875,N_6902);
or U7082 (N_7082,N_6962,N_6941);
nor U7083 (N_7083,N_6908,N_6821);
nor U7084 (N_7084,N_6844,N_6967);
nor U7085 (N_7085,N_6830,N_6863);
nand U7086 (N_7086,N_6889,N_6824);
nand U7087 (N_7087,N_6992,N_6981);
and U7088 (N_7088,N_6896,N_6955);
nor U7089 (N_7089,N_6843,N_6921);
nor U7090 (N_7090,N_6916,N_6851);
or U7091 (N_7091,N_6831,N_6949);
nor U7092 (N_7092,N_6990,N_6957);
nor U7093 (N_7093,N_6877,N_6965);
nor U7094 (N_7094,N_6984,N_6852);
nor U7095 (N_7095,N_6919,N_6804);
or U7096 (N_7096,N_6867,N_6872);
and U7097 (N_7097,N_6953,N_6879);
and U7098 (N_7098,N_6943,N_6833);
and U7099 (N_7099,N_6840,N_6963);
and U7100 (N_7100,N_6929,N_6915);
or U7101 (N_7101,N_6852,N_6802);
xnor U7102 (N_7102,N_6822,N_6922);
nand U7103 (N_7103,N_6847,N_6963);
nand U7104 (N_7104,N_6942,N_6948);
xor U7105 (N_7105,N_6985,N_6810);
or U7106 (N_7106,N_6876,N_6829);
nand U7107 (N_7107,N_6842,N_6872);
nor U7108 (N_7108,N_6817,N_6890);
and U7109 (N_7109,N_6920,N_6810);
and U7110 (N_7110,N_6945,N_6858);
xor U7111 (N_7111,N_6943,N_6992);
xor U7112 (N_7112,N_6942,N_6986);
and U7113 (N_7113,N_6878,N_6990);
nand U7114 (N_7114,N_6989,N_6945);
and U7115 (N_7115,N_6951,N_6901);
and U7116 (N_7116,N_6883,N_6935);
and U7117 (N_7117,N_6943,N_6832);
nand U7118 (N_7118,N_6935,N_6890);
or U7119 (N_7119,N_6868,N_6982);
and U7120 (N_7120,N_6889,N_6877);
nor U7121 (N_7121,N_6843,N_6844);
or U7122 (N_7122,N_6870,N_6862);
or U7123 (N_7123,N_6804,N_6853);
or U7124 (N_7124,N_6874,N_6820);
and U7125 (N_7125,N_6802,N_6988);
or U7126 (N_7126,N_6971,N_6819);
and U7127 (N_7127,N_6963,N_6857);
xnor U7128 (N_7128,N_6948,N_6997);
nor U7129 (N_7129,N_6885,N_6843);
nand U7130 (N_7130,N_6806,N_6851);
nor U7131 (N_7131,N_6918,N_6986);
and U7132 (N_7132,N_6935,N_6838);
or U7133 (N_7133,N_6944,N_6927);
or U7134 (N_7134,N_6809,N_6877);
nor U7135 (N_7135,N_6858,N_6970);
or U7136 (N_7136,N_6905,N_6954);
and U7137 (N_7137,N_6991,N_6934);
and U7138 (N_7138,N_6956,N_6800);
nor U7139 (N_7139,N_6934,N_6984);
nand U7140 (N_7140,N_6875,N_6865);
or U7141 (N_7141,N_6867,N_6885);
nor U7142 (N_7142,N_6905,N_6805);
nand U7143 (N_7143,N_6991,N_6883);
nor U7144 (N_7144,N_6806,N_6826);
nand U7145 (N_7145,N_6877,N_6903);
nor U7146 (N_7146,N_6906,N_6870);
or U7147 (N_7147,N_6993,N_6971);
and U7148 (N_7148,N_6840,N_6918);
or U7149 (N_7149,N_6992,N_6909);
and U7150 (N_7150,N_6952,N_6882);
nor U7151 (N_7151,N_6885,N_6914);
and U7152 (N_7152,N_6927,N_6925);
or U7153 (N_7153,N_6899,N_6859);
nand U7154 (N_7154,N_6843,N_6966);
nand U7155 (N_7155,N_6940,N_6916);
or U7156 (N_7156,N_6890,N_6986);
or U7157 (N_7157,N_6913,N_6905);
or U7158 (N_7158,N_6826,N_6922);
and U7159 (N_7159,N_6871,N_6819);
and U7160 (N_7160,N_6878,N_6958);
nor U7161 (N_7161,N_6846,N_6853);
or U7162 (N_7162,N_6992,N_6802);
nor U7163 (N_7163,N_6800,N_6868);
and U7164 (N_7164,N_6976,N_6869);
nor U7165 (N_7165,N_6806,N_6968);
nor U7166 (N_7166,N_6834,N_6974);
and U7167 (N_7167,N_6868,N_6941);
nor U7168 (N_7168,N_6977,N_6807);
nor U7169 (N_7169,N_6868,N_6954);
nand U7170 (N_7170,N_6847,N_6884);
nand U7171 (N_7171,N_6854,N_6876);
nor U7172 (N_7172,N_6808,N_6910);
or U7173 (N_7173,N_6884,N_6929);
nor U7174 (N_7174,N_6984,N_6905);
and U7175 (N_7175,N_6853,N_6979);
and U7176 (N_7176,N_6970,N_6952);
and U7177 (N_7177,N_6933,N_6866);
or U7178 (N_7178,N_6843,N_6802);
and U7179 (N_7179,N_6804,N_6815);
and U7180 (N_7180,N_6891,N_6899);
or U7181 (N_7181,N_6867,N_6836);
and U7182 (N_7182,N_6869,N_6883);
xnor U7183 (N_7183,N_6881,N_6872);
nand U7184 (N_7184,N_6848,N_6822);
xor U7185 (N_7185,N_6971,N_6973);
or U7186 (N_7186,N_6995,N_6960);
nand U7187 (N_7187,N_6947,N_6896);
or U7188 (N_7188,N_6872,N_6857);
and U7189 (N_7189,N_6942,N_6931);
nor U7190 (N_7190,N_6862,N_6806);
nor U7191 (N_7191,N_6919,N_6876);
xnor U7192 (N_7192,N_6883,N_6829);
and U7193 (N_7193,N_6949,N_6810);
nand U7194 (N_7194,N_6803,N_6870);
and U7195 (N_7195,N_6917,N_6923);
nand U7196 (N_7196,N_6917,N_6921);
xnor U7197 (N_7197,N_6948,N_6928);
nand U7198 (N_7198,N_6834,N_6821);
nand U7199 (N_7199,N_6917,N_6848);
nor U7200 (N_7200,N_7002,N_7027);
or U7201 (N_7201,N_7028,N_7171);
nor U7202 (N_7202,N_7158,N_7029);
or U7203 (N_7203,N_7089,N_7142);
nor U7204 (N_7204,N_7129,N_7099);
nor U7205 (N_7205,N_7172,N_7088);
nand U7206 (N_7206,N_7052,N_7065);
and U7207 (N_7207,N_7127,N_7067);
and U7208 (N_7208,N_7097,N_7141);
nor U7209 (N_7209,N_7133,N_7020);
nand U7210 (N_7210,N_7149,N_7177);
xor U7211 (N_7211,N_7125,N_7160);
or U7212 (N_7212,N_7163,N_7139);
nand U7213 (N_7213,N_7024,N_7076);
nand U7214 (N_7214,N_7032,N_7012);
and U7215 (N_7215,N_7086,N_7015);
and U7216 (N_7216,N_7140,N_7055);
and U7217 (N_7217,N_7187,N_7084);
or U7218 (N_7218,N_7073,N_7131);
or U7219 (N_7219,N_7041,N_7103);
xor U7220 (N_7220,N_7046,N_7036);
and U7221 (N_7221,N_7011,N_7197);
nor U7222 (N_7222,N_7175,N_7098);
nand U7223 (N_7223,N_7121,N_7116);
and U7224 (N_7224,N_7143,N_7115);
nand U7225 (N_7225,N_7092,N_7010);
nand U7226 (N_7226,N_7075,N_7014);
and U7227 (N_7227,N_7007,N_7189);
xnor U7228 (N_7228,N_7164,N_7157);
xor U7229 (N_7229,N_7077,N_7080);
nand U7230 (N_7230,N_7119,N_7057);
nor U7231 (N_7231,N_7153,N_7144);
nor U7232 (N_7232,N_7025,N_7062);
nor U7233 (N_7233,N_7083,N_7078);
or U7234 (N_7234,N_7043,N_7009);
or U7235 (N_7235,N_7174,N_7165);
or U7236 (N_7236,N_7019,N_7048);
or U7237 (N_7237,N_7114,N_7108);
xnor U7238 (N_7238,N_7136,N_7182);
nor U7239 (N_7239,N_7094,N_7045);
nand U7240 (N_7240,N_7072,N_7156);
xor U7241 (N_7241,N_7060,N_7179);
or U7242 (N_7242,N_7022,N_7113);
nor U7243 (N_7243,N_7054,N_7190);
or U7244 (N_7244,N_7017,N_7066);
or U7245 (N_7245,N_7069,N_7071);
nand U7246 (N_7246,N_7008,N_7162);
nor U7247 (N_7247,N_7124,N_7035);
nand U7248 (N_7248,N_7150,N_7167);
nor U7249 (N_7249,N_7111,N_7159);
or U7250 (N_7250,N_7166,N_7102);
nand U7251 (N_7251,N_7181,N_7056);
or U7252 (N_7252,N_7090,N_7037);
xnor U7253 (N_7253,N_7064,N_7161);
nor U7254 (N_7254,N_7132,N_7180);
and U7255 (N_7255,N_7001,N_7130);
or U7256 (N_7256,N_7034,N_7155);
nand U7257 (N_7257,N_7018,N_7151);
and U7258 (N_7258,N_7061,N_7118);
nand U7259 (N_7259,N_7152,N_7199);
xnor U7260 (N_7260,N_7100,N_7039);
or U7261 (N_7261,N_7185,N_7138);
xor U7262 (N_7262,N_7194,N_7112);
nor U7263 (N_7263,N_7068,N_7148);
and U7264 (N_7264,N_7146,N_7154);
and U7265 (N_7265,N_7091,N_7195);
or U7266 (N_7266,N_7169,N_7042);
xor U7267 (N_7267,N_7135,N_7079);
nand U7268 (N_7268,N_7176,N_7003);
nor U7269 (N_7269,N_7059,N_7074);
and U7270 (N_7270,N_7147,N_7110);
and U7271 (N_7271,N_7081,N_7040);
or U7272 (N_7272,N_7053,N_7168);
nor U7273 (N_7273,N_7109,N_7122);
and U7274 (N_7274,N_7106,N_7023);
and U7275 (N_7275,N_7026,N_7050);
or U7276 (N_7276,N_7093,N_7101);
and U7277 (N_7277,N_7193,N_7047);
nor U7278 (N_7278,N_7192,N_7123);
nor U7279 (N_7279,N_7038,N_7087);
and U7280 (N_7280,N_7004,N_7196);
and U7281 (N_7281,N_7082,N_7191);
or U7282 (N_7282,N_7031,N_7096);
xnor U7283 (N_7283,N_7051,N_7005);
and U7284 (N_7284,N_7044,N_7006);
or U7285 (N_7285,N_7120,N_7016);
or U7286 (N_7286,N_7145,N_7178);
or U7287 (N_7287,N_7198,N_7188);
nand U7288 (N_7288,N_7128,N_7049);
and U7289 (N_7289,N_7170,N_7104);
and U7290 (N_7290,N_7013,N_7021);
nor U7291 (N_7291,N_7184,N_7058);
nor U7292 (N_7292,N_7030,N_7063);
and U7293 (N_7293,N_7137,N_7126);
nand U7294 (N_7294,N_7095,N_7033);
nor U7295 (N_7295,N_7107,N_7117);
nand U7296 (N_7296,N_7000,N_7173);
nor U7297 (N_7297,N_7183,N_7134);
and U7298 (N_7298,N_7085,N_7105);
nor U7299 (N_7299,N_7186,N_7070);
xnor U7300 (N_7300,N_7064,N_7075);
and U7301 (N_7301,N_7112,N_7123);
nand U7302 (N_7302,N_7001,N_7005);
or U7303 (N_7303,N_7022,N_7019);
xnor U7304 (N_7304,N_7017,N_7008);
nor U7305 (N_7305,N_7003,N_7173);
and U7306 (N_7306,N_7148,N_7096);
and U7307 (N_7307,N_7052,N_7081);
or U7308 (N_7308,N_7141,N_7167);
nand U7309 (N_7309,N_7106,N_7010);
nor U7310 (N_7310,N_7044,N_7154);
or U7311 (N_7311,N_7018,N_7060);
xnor U7312 (N_7312,N_7108,N_7191);
or U7313 (N_7313,N_7153,N_7141);
nor U7314 (N_7314,N_7057,N_7006);
xnor U7315 (N_7315,N_7077,N_7020);
xor U7316 (N_7316,N_7084,N_7040);
nand U7317 (N_7317,N_7081,N_7086);
and U7318 (N_7318,N_7147,N_7015);
nand U7319 (N_7319,N_7109,N_7057);
and U7320 (N_7320,N_7198,N_7032);
or U7321 (N_7321,N_7004,N_7068);
and U7322 (N_7322,N_7176,N_7159);
nand U7323 (N_7323,N_7177,N_7195);
and U7324 (N_7324,N_7037,N_7045);
nor U7325 (N_7325,N_7142,N_7155);
nand U7326 (N_7326,N_7131,N_7048);
xor U7327 (N_7327,N_7040,N_7048);
nand U7328 (N_7328,N_7135,N_7004);
nand U7329 (N_7329,N_7131,N_7199);
and U7330 (N_7330,N_7177,N_7168);
nand U7331 (N_7331,N_7164,N_7174);
or U7332 (N_7332,N_7029,N_7047);
nand U7333 (N_7333,N_7197,N_7054);
nand U7334 (N_7334,N_7113,N_7083);
nand U7335 (N_7335,N_7185,N_7057);
nand U7336 (N_7336,N_7106,N_7070);
nor U7337 (N_7337,N_7055,N_7071);
or U7338 (N_7338,N_7098,N_7178);
nand U7339 (N_7339,N_7107,N_7140);
nor U7340 (N_7340,N_7154,N_7040);
or U7341 (N_7341,N_7181,N_7044);
and U7342 (N_7342,N_7044,N_7182);
nor U7343 (N_7343,N_7163,N_7090);
xor U7344 (N_7344,N_7006,N_7039);
nand U7345 (N_7345,N_7033,N_7082);
nand U7346 (N_7346,N_7172,N_7197);
nand U7347 (N_7347,N_7147,N_7166);
and U7348 (N_7348,N_7165,N_7077);
nand U7349 (N_7349,N_7078,N_7000);
or U7350 (N_7350,N_7100,N_7001);
xnor U7351 (N_7351,N_7185,N_7014);
or U7352 (N_7352,N_7184,N_7198);
xnor U7353 (N_7353,N_7017,N_7098);
and U7354 (N_7354,N_7159,N_7098);
nand U7355 (N_7355,N_7068,N_7009);
and U7356 (N_7356,N_7101,N_7153);
or U7357 (N_7357,N_7034,N_7045);
nand U7358 (N_7358,N_7037,N_7043);
nor U7359 (N_7359,N_7116,N_7103);
nor U7360 (N_7360,N_7172,N_7017);
nand U7361 (N_7361,N_7007,N_7084);
or U7362 (N_7362,N_7001,N_7056);
xor U7363 (N_7363,N_7001,N_7031);
nand U7364 (N_7364,N_7002,N_7190);
and U7365 (N_7365,N_7091,N_7175);
or U7366 (N_7366,N_7145,N_7057);
and U7367 (N_7367,N_7121,N_7190);
nand U7368 (N_7368,N_7062,N_7108);
nor U7369 (N_7369,N_7011,N_7176);
and U7370 (N_7370,N_7012,N_7080);
or U7371 (N_7371,N_7059,N_7134);
xor U7372 (N_7372,N_7108,N_7077);
nand U7373 (N_7373,N_7011,N_7136);
nor U7374 (N_7374,N_7141,N_7195);
or U7375 (N_7375,N_7196,N_7084);
and U7376 (N_7376,N_7158,N_7197);
nor U7377 (N_7377,N_7101,N_7107);
and U7378 (N_7378,N_7058,N_7016);
nand U7379 (N_7379,N_7129,N_7053);
or U7380 (N_7380,N_7012,N_7120);
and U7381 (N_7381,N_7141,N_7046);
or U7382 (N_7382,N_7129,N_7112);
or U7383 (N_7383,N_7122,N_7198);
or U7384 (N_7384,N_7128,N_7160);
xnor U7385 (N_7385,N_7199,N_7195);
nor U7386 (N_7386,N_7066,N_7169);
xnor U7387 (N_7387,N_7153,N_7158);
nor U7388 (N_7388,N_7144,N_7139);
nor U7389 (N_7389,N_7196,N_7074);
or U7390 (N_7390,N_7070,N_7147);
or U7391 (N_7391,N_7186,N_7045);
and U7392 (N_7392,N_7097,N_7011);
and U7393 (N_7393,N_7023,N_7112);
and U7394 (N_7394,N_7079,N_7016);
nand U7395 (N_7395,N_7003,N_7140);
nand U7396 (N_7396,N_7097,N_7134);
and U7397 (N_7397,N_7128,N_7070);
or U7398 (N_7398,N_7054,N_7053);
and U7399 (N_7399,N_7120,N_7172);
and U7400 (N_7400,N_7361,N_7215);
or U7401 (N_7401,N_7203,N_7341);
nor U7402 (N_7402,N_7373,N_7248);
nand U7403 (N_7403,N_7290,N_7340);
and U7404 (N_7404,N_7278,N_7320);
nand U7405 (N_7405,N_7225,N_7224);
nor U7406 (N_7406,N_7277,N_7398);
or U7407 (N_7407,N_7218,N_7210);
nor U7408 (N_7408,N_7307,N_7217);
nand U7409 (N_7409,N_7253,N_7230);
or U7410 (N_7410,N_7383,N_7310);
and U7411 (N_7411,N_7243,N_7232);
or U7412 (N_7412,N_7319,N_7212);
nand U7413 (N_7413,N_7365,N_7234);
nand U7414 (N_7414,N_7297,N_7386);
xor U7415 (N_7415,N_7244,N_7282);
nand U7416 (N_7416,N_7357,N_7255);
and U7417 (N_7417,N_7382,N_7350);
and U7418 (N_7418,N_7270,N_7273);
or U7419 (N_7419,N_7304,N_7385);
and U7420 (N_7420,N_7211,N_7393);
or U7421 (N_7421,N_7342,N_7262);
and U7422 (N_7422,N_7374,N_7266);
nand U7423 (N_7423,N_7205,N_7301);
nor U7424 (N_7424,N_7242,N_7275);
nand U7425 (N_7425,N_7269,N_7387);
and U7426 (N_7426,N_7256,N_7376);
or U7427 (N_7427,N_7254,N_7207);
or U7428 (N_7428,N_7231,N_7292);
nor U7429 (N_7429,N_7209,N_7330);
or U7430 (N_7430,N_7293,N_7276);
and U7431 (N_7431,N_7285,N_7399);
or U7432 (N_7432,N_7344,N_7337);
xor U7433 (N_7433,N_7368,N_7331);
nor U7434 (N_7434,N_7363,N_7332);
and U7435 (N_7435,N_7206,N_7287);
xor U7436 (N_7436,N_7325,N_7298);
nor U7437 (N_7437,N_7247,N_7346);
nand U7438 (N_7438,N_7226,N_7371);
nor U7439 (N_7439,N_7334,N_7321);
and U7440 (N_7440,N_7313,N_7216);
or U7441 (N_7441,N_7221,N_7267);
or U7442 (N_7442,N_7351,N_7388);
nor U7443 (N_7443,N_7263,N_7309);
xnor U7444 (N_7444,N_7349,N_7366);
nor U7445 (N_7445,N_7359,N_7397);
or U7446 (N_7446,N_7348,N_7236);
nand U7447 (N_7447,N_7245,N_7239);
nand U7448 (N_7448,N_7360,N_7324);
nand U7449 (N_7449,N_7315,N_7312);
nand U7450 (N_7450,N_7335,N_7364);
nor U7451 (N_7451,N_7272,N_7302);
or U7452 (N_7452,N_7378,N_7289);
xnor U7453 (N_7453,N_7392,N_7294);
nand U7454 (N_7454,N_7229,N_7260);
and U7455 (N_7455,N_7258,N_7201);
and U7456 (N_7456,N_7317,N_7326);
xnor U7457 (N_7457,N_7252,N_7384);
or U7458 (N_7458,N_7303,N_7327);
nand U7459 (N_7459,N_7264,N_7235);
or U7460 (N_7460,N_7299,N_7339);
xnor U7461 (N_7461,N_7358,N_7316);
nand U7462 (N_7462,N_7271,N_7246);
nor U7463 (N_7463,N_7333,N_7250);
nand U7464 (N_7464,N_7311,N_7370);
nand U7465 (N_7465,N_7259,N_7338);
or U7466 (N_7466,N_7240,N_7222);
nor U7467 (N_7467,N_7377,N_7306);
nand U7468 (N_7468,N_7261,N_7295);
nor U7469 (N_7469,N_7268,N_7214);
and U7470 (N_7470,N_7355,N_7237);
nand U7471 (N_7471,N_7228,N_7202);
nor U7472 (N_7472,N_7362,N_7322);
nor U7473 (N_7473,N_7395,N_7227);
or U7474 (N_7474,N_7219,N_7329);
nand U7475 (N_7475,N_7233,N_7208);
nand U7476 (N_7476,N_7291,N_7220);
nand U7477 (N_7477,N_7249,N_7394);
nand U7478 (N_7478,N_7318,N_7354);
or U7479 (N_7479,N_7390,N_7391);
or U7480 (N_7480,N_7381,N_7204);
or U7481 (N_7481,N_7300,N_7389);
or U7482 (N_7482,N_7367,N_7265);
and U7483 (N_7483,N_7336,N_7352);
or U7484 (N_7484,N_7279,N_7251);
or U7485 (N_7485,N_7288,N_7328);
nor U7486 (N_7486,N_7286,N_7241);
nand U7487 (N_7487,N_7296,N_7345);
nor U7488 (N_7488,N_7200,N_7396);
nor U7489 (N_7489,N_7343,N_7283);
and U7490 (N_7490,N_7284,N_7356);
or U7491 (N_7491,N_7281,N_7379);
nor U7492 (N_7492,N_7274,N_7314);
and U7493 (N_7493,N_7380,N_7308);
nand U7494 (N_7494,N_7353,N_7257);
nor U7495 (N_7495,N_7238,N_7369);
nor U7496 (N_7496,N_7305,N_7223);
or U7497 (N_7497,N_7280,N_7347);
nor U7498 (N_7498,N_7213,N_7375);
and U7499 (N_7499,N_7372,N_7323);
nor U7500 (N_7500,N_7285,N_7204);
nor U7501 (N_7501,N_7228,N_7367);
nor U7502 (N_7502,N_7324,N_7215);
or U7503 (N_7503,N_7217,N_7319);
and U7504 (N_7504,N_7281,N_7372);
or U7505 (N_7505,N_7325,N_7282);
and U7506 (N_7506,N_7356,N_7366);
or U7507 (N_7507,N_7310,N_7238);
nor U7508 (N_7508,N_7350,N_7222);
and U7509 (N_7509,N_7207,N_7244);
nor U7510 (N_7510,N_7270,N_7250);
nand U7511 (N_7511,N_7242,N_7204);
nand U7512 (N_7512,N_7319,N_7317);
nor U7513 (N_7513,N_7221,N_7329);
and U7514 (N_7514,N_7344,N_7235);
and U7515 (N_7515,N_7245,N_7398);
or U7516 (N_7516,N_7306,N_7244);
or U7517 (N_7517,N_7208,N_7252);
nand U7518 (N_7518,N_7277,N_7286);
nand U7519 (N_7519,N_7254,N_7230);
or U7520 (N_7520,N_7393,N_7336);
and U7521 (N_7521,N_7354,N_7323);
or U7522 (N_7522,N_7237,N_7343);
nand U7523 (N_7523,N_7263,N_7217);
nand U7524 (N_7524,N_7319,N_7293);
nand U7525 (N_7525,N_7298,N_7280);
nor U7526 (N_7526,N_7363,N_7276);
nor U7527 (N_7527,N_7388,N_7390);
and U7528 (N_7528,N_7393,N_7338);
or U7529 (N_7529,N_7313,N_7309);
nand U7530 (N_7530,N_7325,N_7365);
nor U7531 (N_7531,N_7202,N_7264);
or U7532 (N_7532,N_7328,N_7210);
or U7533 (N_7533,N_7250,N_7393);
xor U7534 (N_7534,N_7311,N_7230);
nor U7535 (N_7535,N_7327,N_7202);
nor U7536 (N_7536,N_7216,N_7353);
nand U7537 (N_7537,N_7391,N_7396);
nor U7538 (N_7538,N_7282,N_7338);
nor U7539 (N_7539,N_7239,N_7295);
nand U7540 (N_7540,N_7283,N_7339);
nor U7541 (N_7541,N_7309,N_7259);
nor U7542 (N_7542,N_7259,N_7213);
or U7543 (N_7543,N_7362,N_7235);
nand U7544 (N_7544,N_7398,N_7268);
nand U7545 (N_7545,N_7320,N_7398);
nand U7546 (N_7546,N_7346,N_7249);
xnor U7547 (N_7547,N_7215,N_7344);
and U7548 (N_7548,N_7274,N_7300);
nand U7549 (N_7549,N_7302,N_7200);
nor U7550 (N_7550,N_7381,N_7242);
or U7551 (N_7551,N_7227,N_7239);
nor U7552 (N_7552,N_7202,N_7225);
or U7553 (N_7553,N_7383,N_7277);
nor U7554 (N_7554,N_7211,N_7205);
or U7555 (N_7555,N_7216,N_7295);
nand U7556 (N_7556,N_7389,N_7269);
or U7557 (N_7557,N_7229,N_7366);
nor U7558 (N_7558,N_7371,N_7379);
nor U7559 (N_7559,N_7323,N_7394);
and U7560 (N_7560,N_7298,N_7305);
nand U7561 (N_7561,N_7275,N_7254);
nor U7562 (N_7562,N_7269,N_7203);
nand U7563 (N_7563,N_7211,N_7369);
and U7564 (N_7564,N_7351,N_7315);
nor U7565 (N_7565,N_7372,N_7321);
or U7566 (N_7566,N_7371,N_7307);
xor U7567 (N_7567,N_7390,N_7220);
xor U7568 (N_7568,N_7346,N_7318);
xnor U7569 (N_7569,N_7312,N_7268);
nand U7570 (N_7570,N_7355,N_7333);
and U7571 (N_7571,N_7293,N_7214);
and U7572 (N_7572,N_7275,N_7371);
and U7573 (N_7573,N_7263,N_7291);
or U7574 (N_7574,N_7390,N_7291);
xnor U7575 (N_7575,N_7337,N_7270);
and U7576 (N_7576,N_7398,N_7330);
xnor U7577 (N_7577,N_7251,N_7392);
xnor U7578 (N_7578,N_7303,N_7309);
xor U7579 (N_7579,N_7244,N_7317);
nand U7580 (N_7580,N_7293,N_7344);
or U7581 (N_7581,N_7326,N_7348);
nand U7582 (N_7582,N_7385,N_7332);
nand U7583 (N_7583,N_7314,N_7397);
nor U7584 (N_7584,N_7368,N_7353);
or U7585 (N_7585,N_7223,N_7369);
nor U7586 (N_7586,N_7282,N_7395);
xnor U7587 (N_7587,N_7335,N_7274);
nand U7588 (N_7588,N_7226,N_7297);
nor U7589 (N_7589,N_7211,N_7228);
and U7590 (N_7590,N_7306,N_7379);
or U7591 (N_7591,N_7295,N_7343);
or U7592 (N_7592,N_7374,N_7371);
nor U7593 (N_7593,N_7242,N_7370);
and U7594 (N_7594,N_7300,N_7204);
and U7595 (N_7595,N_7242,N_7327);
or U7596 (N_7596,N_7284,N_7303);
and U7597 (N_7597,N_7309,N_7256);
nor U7598 (N_7598,N_7389,N_7351);
nand U7599 (N_7599,N_7359,N_7299);
nor U7600 (N_7600,N_7559,N_7427);
xnor U7601 (N_7601,N_7403,N_7520);
and U7602 (N_7602,N_7540,N_7517);
and U7603 (N_7603,N_7407,N_7417);
or U7604 (N_7604,N_7422,N_7414);
or U7605 (N_7605,N_7584,N_7457);
and U7606 (N_7606,N_7502,N_7596);
nand U7607 (N_7607,N_7454,N_7558);
nand U7608 (N_7608,N_7587,N_7419);
nor U7609 (N_7609,N_7543,N_7553);
nor U7610 (N_7610,N_7595,N_7577);
or U7611 (N_7611,N_7442,N_7489);
or U7612 (N_7612,N_7556,N_7477);
and U7613 (N_7613,N_7592,N_7416);
xnor U7614 (N_7614,N_7463,N_7492);
xor U7615 (N_7615,N_7515,N_7598);
and U7616 (N_7616,N_7519,N_7464);
nand U7617 (N_7617,N_7410,N_7538);
and U7618 (N_7618,N_7514,N_7567);
nor U7619 (N_7619,N_7491,N_7572);
and U7620 (N_7620,N_7579,N_7445);
nand U7621 (N_7621,N_7505,N_7420);
nor U7622 (N_7622,N_7508,N_7503);
xor U7623 (N_7623,N_7441,N_7495);
and U7624 (N_7624,N_7458,N_7487);
nand U7625 (N_7625,N_7561,N_7466);
and U7626 (N_7626,N_7449,N_7448);
xor U7627 (N_7627,N_7560,N_7440);
or U7628 (N_7628,N_7435,N_7564);
nor U7629 (N_7629,N_7479,N_7493);
nor U7630 (N_7630,N_7524,N_7428);
or U7631 (N_7631,N_7462,N_7548);
and U7632 (N_7632,N_7451,N_7532);
nor U7633 (N_7633,N_7480,N_7537);
and U7634 (N_7634,N_7574,N_7573);
nand U7635 (N_7635,N_7534,N_7585);
xnor U7636 (N_7636,N_7578,N_7599);
nand U7637 (N_7637,N_7405,N_7406);
and U7638 (N_7638,N_7516,N_7562);
xor U7639 (N_7639,N_7402,N_7588);
nand U7640 (N_7640,N_7507,N_7437);
or U7641 (N_7641,N_7409,N_7460);
nor U7642 (N_7642,N_7575,N_7509);
nor U7643 (N_7643,N_7597,N_7455);
or U7644 (N_7644,N_7552,N_7412);
xor U7645 (N_7645,N_7468,N_7506);
nor U7646 (N_7646,N_7533,N_7484);
or U7647 (N_7647,N_7496,N_7467);
nand U7648 (N_7648,N_7539,N_7518);
nor U7649 (N_7649,N_7404,N_7485);
and U7650 (N_7650,N_7513,N_7408);
xor U7651 (N_7651,N_7446,N_7433);
nor U7652 (N_7652,N_7547,N_7541);
or U7653 (N_7653,N_7554,N_7447);
nor U7654 (N_7654,N_7499,N_7498);
nand U7655 (N_7655,N_7456,N_7418);
nor U7656 (N_7656,N_7424,N_7400);
and U7657 (N_7657,N_7443,N_7583);
or U7658 (N_7658,N_7415,N_7571);
nor U7659 (N_7659,N_7581,N_7545);
or U7660 (N_7660,N_7555,N_7565);
or U7661 (N_7661,N_7531,N_7476);
and U7662 (N_7662,N_7439,N_7459);
xnor U7663 (N_7663,N_7486,N_7526);
nor U7664 (N_7664,N_7472,N_7490);
nor U7665 (N_7665,N_7401,N_7474);
nor U7666 (N_7666,N_7557,N_7542);
or U7667 (N_7667,N_7551,N_7528);
and U7668 (N_7668,N_7434,N_7501);
nor U7669 (N_7669,N_7510,N_7421);
nand U7670 (N_7670,N_7453,N_7594);
and U7671 (N_7671,N_7494,N_7527);
nand U7672 (N_7672,N_7444,N_7580);
nand U7673 (N_7673,N_7576,N_7593);
nor U7674 (N_7674,N_7563,N_7500);
nor U7675 (N_7675,N_7429,N_7469);
and U7676 (N_7676,N_7525,N_7550);
or U7677 (N_7677,N_7530,N_7478);
or U7678 (N_7678,N_7461,N_7436);
nor U7679 (N_7679,N_7452,N_7522);
or U7680 (N_7680,N_7566,N_7582);
or U7681 (N_7681,N_7423,N_7497);
nor U7682 (N_7682,N_7512,N_7529);
and U7683 (N_7683,N_7483,N_7504);
or U7684 (N_7684,N_7569,N_7590);
xor U7685 (N_7685,N_7535,N_7426);
or U7686 (N_7686,N_7411,N_7536);
or U7687 (N_7687,N_7438,N_7430);
or U7688 (N_7688,N_7568,N_7570);
or U7689 (N_7689,N_7471,N_7549);
nor U7690 (N_7690,N_7511,N_7470);
or U7691 (N_7691,N_7586,N_7432);
nand U7692 (N_7692,N_7482,N_7521);
or U7693 (N_7693,N_7589,N_7431);
nor U7694 (N_7694,N_7488,N_7523);
nor U7695 (N_7695,N_7544,N_7546);
nand U7696 (N_7696,N_7425,N_7591);
and U7697 (N_7697,N_7481,N_7475);
and U7698 (N_7698,N_7450,N_7413);
nand U7699 (N_7699,N_7473,N_7465);
and U7700 (N_7700,N_7511,N_7552);
and U7701 (N_7701,N_7578,N_7421);
nor U7702 (N_7702,N_7555,N_7536);
nor U7703 (N_7703,N_7404,N_7542);
and U7704 (N_7704,N_7524,N_7514);
and U7705 (N_7705,N_7478,N_7519);
or U7706 (N_7706,N_7407,N_7475);
nand U7707 (N_7707,N_7480,N_7498);
nand U7708 (N_7708,N_7453,N_7460);
nor U7709 (N_7709,N_7597,N_7400);
nor U7710 (N_7710,N_7538,N_7404);
xnor U7711 (N_7711,N_7449,N_7531);
xnor U7712 (N_7712,N_7413,N_7578);
xor U7713 (N_7713,N_7542,N_7550);
and U7714 (N_7714,N_7409,N_7468);
or U7715 (N_7715,N_7520,N_7531);
or U7716 (N_7716,N_7494,N_7525);
nor U7717 (N_7717,N_7539,N_7417);
or U7718 (N_7718,N_7476,N_7551);
nor U7719 (N_7719,N_7568,N_7452);
or U7720 (N_7720,N_7556,N_7501);
and U7721 (N_7721,N_7476,N_7546);
nor U7722 (N_7722,N_7498,N_7421);
nor U7723 (N_7723,N_7511,N_7503);
xnor U7724 (N_7724,N_7589,N_7424);
or U7725 (N_7725,N_7436,N_7574);
nor U7726 (N_7726,N_7515,N_7505);
or U7727 (N_7727,N_7446,N_7532);
nor U7728 (N_7728,N_7565,N_7473);
xor U7729 (N_7729,N_7493,N_7454);
and U7730 (N_7730,N_7529,N_7508);
or U7731 (N_7731,N_7550,N_7452);
nand U7732 (N_7732,N_7545,N_7582);
or U7733 (N_7733,N_7568,N_7544);
nor U7734 (N_7734,N_7441,N_7498);
nand U7735 (N_7735,N_7550,N_7497);
nand U7736 (N_7736,N_7528,N_7501);
nand U7737 (N_7737,N_7523,N_7532);
xor U7738 (N_7738,N_7512,N_7517);
xor U7739 (N_7739,N_7455,N_7432);
or U7740 (N_7740,N_7579,N_7454);
nand U7741 (N_7741,N_7414,N_7568);
and U7742 (N_7742,N_7406,N_7545);
and U7743 (N_7743,N_7513,N_7511);
or U7744 (N_7744,N_7586,N_7427);
nand U7745 (N_7745,N_7487,N_7420);
nand U7746 (N_7746,N_7446,N_7459);
nor U7747 (N_7747,N_7449,N_7480);
xor U7748 (N_7748,N_7480,N_7543);
nor U7749 (N_7749,N_7407,N_7504);
nor U7750 (N_7750,N_7550,N_7444);
nor U7751 (N_7751,N_7498,N_7431);
xor U7752 (N_7752,N_7547,N_7577);
nand U7753 (N_7753,N_7487,N_7412);
xor U7754 (N_7754,N_7469,N_7512);
nand U7755 (N_7755,N_7496,N_7460);
and U7756 (N_7756,N_7485,N_7417);
and U7757 (N_7757,N_7468,N_7436);
and U7758 (N_7758,N_7507,N_7596);
nand U7759 (N_7759,N_7460,N_7438);
nand U7760 (N_7760,N_7582,N_7515);
nor U7761 (N_7761,N_7413,N_7576);
and U7762 (N_7762,N_7590,N_7492);
xor U7763 (N_7763,N_7508,N_7534);
nor U7764 (N_7764,N_7451,N_7538);
xnor U7765 (N_7765,N_7429,N_7502);
or U7766 (N_7766,N_7468,N_7559);
and U7767 (N_7767,N_7570,N_7438);
xnor U7768 (N_7768,N_7584,N_7505);
or U7769 (N_7769,N_7400,N_7402);
nor U7770 (N_7770,N_7596,N_7524);
and U7771 (N_7771,N_7525,N_7539);
xor U7772 (N_7772,N_7486,N_7417);
and U7773 (N_7773,N_7592,N_7472);
nor U7774 (N_7774,N_7595,N_7427);
nand U7775 (N_7775,N_7529,N_7546);
nor U7776 (N_7776,N_7521,N_7492);
nor U7777 (N_7777,N_7502,N_7571);
nand U7778 (N_7778,N_7544,N_7487);
or U7779 (N_7779,N_7491,N_7521);
nor U7780 (N_7780,N_7509,N_7411);
and U7781 (N_7781,N_7424,N_7587);
nand U7782 (N_7782,N_7410,N_7455);
xor U7783 (N_7783,N_7416,N_7443);
and U7784 (N_7784,N_7445,N_7556);
and U7785 (N_7785,N_7563,N_7440);
nand U7786 (N_7786,N_7554,N_7559);
nand U7787 (N_7787,N_7472,N_7433);
nor U7788 (N_7788,N_7400,N_7408);
nand U7789 (N_7789,N_7511,N_7455);
xnor U7790 (N_7790,N_7497,N_7475);
or U7791 (N_7791,N_7463,N_7490);
xnor U7792 (N_7792,N_7439,N_7410);
nor U7793 (N_7793,N_7474,N_7590);
and U7794 (N_7794,N_7483,N_7555);
nand U7795 (N_7795,N_7494,N_7587);
nor U7796 (N_7796,N_7585,N_7439);
nand U7797 (N_7797,N_7424,N_7481);
nor U7798 (N_7798,N_7575,N_7475);
or U7799 (N_7799,N_7418,N_7521);
and U7800 (N_7800,N_7767,N_7774);
nor U7801 (N_7801,N_7699,N_7729);
nand U7802 (N_7802,N_7702,N_7704);
and U7803 (N_7803,N_7621,N_7694);
nand U7804 (N_7804,N_7790,N_7656);
nand U7805 (N_7805,N_7770,N_7691);
and U7806 (N_7806,N_7666,N_7635);
nand U7807 (N_7807,N_7605,N_7636);
or U7808 (N_7808,N_7752,N_7646);
and U7809 (N_7809,N_7747,N_7756);
nand U7810 (N_7810,N_7692,N_7670);
xor U7811 (N_7811,N_7630,N_7719);
or U7812 (N_7812,N_7687,N_7640);
and U7813 (N_7813,N_7654,N_7686);
xor U7814 (N_7814,N_7758,N_7781);
nand U7815 (N_7815,N_7768,N_7753);
or U7816 (N_7816,N_7754,N_7784);
nor U7817 (N_7817,N_7705,N_7649);
xor U7818 (N_7818,N_7678,N_7736);
nand U7819 (N_7819,N_7602,N_7671);
nand U7820 (N_7820,N_7600,N_7771);
and U7821 (N_7821,N_7603,N_7657);
and U7822 (N_7822,N_7759,N_7718);
or U7823 (N_7823,N_7628,N_7651);
or U7824 (N_7824,N_7742,N_7608);
xor U7825 (N_7825,N_7609,N_7750);
nand U7826 (N_7826,N_7757,N_7737);
and U7827 (N_7827,N_7785,N_7783);
and U7828 (N_7828,N_7761,N_7683);
and U7829 (N_7829,N_7776,N_7786);
nor U7830 (N_7830,N_7763,N_7659);
nand U7831 (N_7831,N_7732,N_7633);
or U7832 (N_7832,N_7798,N_7795);
nand U7833 (N_7833,N_7637,N_7679);
nor U7834 (N_7834,N_7658,N_7741);
nand U7835 (N_7835,N_7780,N_7764);
nand U7836 (N_7836,N_7645,N_7601);
or U7837 (N_7837,N_7669,N_7690);
and U7838 (N_7838,N_7662,N_7748);
nor U7839 (N_7839,N_7665,N_7627);
and U7840 (N_7840,N_7625,N_7725);
nor U7841 (N_7841,N_7643,N_7778);
and U7842 (N_7842,N_7751,N_7641);
nor U7843 (N_7843,N_7755,N_7744);
nor U7844 (N_7844,N_7782,N_7639);
and U7845 (N_7845,N_7762,N_7723);
and U7846 (N_7846,N_7619,N_7675);
xnor U7847 (N_7847,N_7617,N_7726);
nor U7848 (N_7848,N_7700,N_7722);
nor U7849 (N_7849,N_7735,N_7655);
and U7850 (N_7850,N_7697,N_7799);
nand U7851 (N_7851,N_7611,N_7624);
and U7852 (N_7852,N_7733,N_7703);
or U7853 (N_7853,N_7727,N_7728);
xor U7854 (N_7854,N_7673,N_7779);
or U7855 (N_7855,N_7710,N_7769);
nand U7856 (N_7856,N_7707,N_7745);
nand U7857 (N_7857,N_7661,N_7650);
nand U7858 (N_7858,N_7731,N_7613);
or U7859 (N_7859,N_7631,N_7775);
xnor U7860 (N_7860,N_7652,N_7711);
nor U7861 (N_7861,N_7701,N_7629);
or U7862 (N_7862,N_7712,N_7743);
nand U7863 (N_7863,N_7715,N_7680);
nor U7864 (N_7864,N_7668,N_7787);
or U7865 (N_7865,N_7653,N_7738);
nor U7866 (N_7866,N_7794,N_7713);
nand U7867 (N_7867,N_7615,N_7777);
nand U7868 (N_7868,N_7667,N_7664);
or U7869 (N_7869,N_7695,N_7724);
nor U7870 (N_7870,N_7638,N_7610);
xor U7871 (N_7871,N_7663,N_7720);
and U7872 (N_7872,N_7788,N_7672);
or U7873 (N_7873,N_7616,N_7730);
nor U7874 (N_7874,N_7689,N_7717);
or U7875 (N_7875,N_7674,N_7676);
and U7876 (N_7876,N_7688,N_7708);
xnor U7877 (N_7877,N_7706,N_7772);
and U7878 (N_7878,N_7791,N_7620);
nor U7879 (N_7879,N_7714,N_7740);
nand U7880 (N_7880,N_7749,N_7622);
and U7881 (N_7881,N_7793,N_7696);
and U7882 (N_7882,N_7614,N_7623);
or U7883 (N_7883,N_7648,N_7739);
nand U7884 (N_7884,N_7765,N_7685);
xor U7885 (N_7885,N_7681,N_7660);
or U7886 (N_7886,N_7607,N_7682);
nand U7887 (N_7887,N_7766,N_7684);
nor U7888 (N_7888,N_7721,N_7632);
or U7889 (N_7889,N_7644,N_7693);
nand U7890 (N_7890,N_7773,N_7606);
nand U7891 (N_7891,N_7698,N_7677);
nor U7892 (N_7892,N_7716,N_7789);
and U7893 (N_7893,N_7647,N_7797);
nor U7894 (N_7894,N_7760,N_7618);
or U7895 (N_7895,N_7612,N_7734);
nor U7896 (N_7896,N_7746,N_7626);
nor U7897 (N_7897,N_7796,N_7634);
nor U7898 (N_7898,N_7642,N_7792);
or U7899 (N_7899,N_7604,N_7709);
and U7900 (N_7900,N_7600,N_7726);
nand U7901 (N_7901,N_7664,N_7762);
nand U7902 (N_7902,N_7735,N_7798);
nand U7903 (N_7903,N_7617,N_7745);
nor U7904 (N_7904,N_7783,N_7698);
and U7905 (N_7905,N_7667,N_7710);
and U7906 (N_7906,N_7753,N_7640);
or U7907 (N_7907,N_7669,N_7634);
xnor U7908 (N_7908,N_7739,N_7742);
or U7909 (N_7909,N_7655,N_7629);
xnor U7910 (N_7910,N_7645,N_7618);
and U7911 (N_7911,N_7795,N_7742);
or U7912 (N_7912,N_7770,N_7678);
and U7913 (N_7913,N_7644,N_7672);
or U7914 (N_7914,N_7716,N_7680);
and U7915 (N_7915,N_7757,N_7655);
nor U7916 (N_7916,N_7736,N_7751);
and U7917 (N_7917,N_7648,N_7760);
nor U7918 (N_7918,N_7726,N_7671);
xnor U7919 (N_7919,N_7767,N_7654);
or U7920 (N_7920,N_7715,N_7666);
nor U7921 (N_7921,N_7750,N_7739);
xnor U7922 (N_7922,N_7754,N_7686);
or U7923 (N_7923,N_7691,N_7736);
and U7924 (N_7924,N_7729,N_7669);
and U7925 (N_7925,N_7629,N_7625);
nand U7926 (N_7926,N_7709,N_7608);
nand U7927 (N_7927,N_7662,N_7718);
nor U7928 (N_7928,N_7614,N_7625);
and U7929 (N_7929,N_7790,N_7792);
xnor U7930 (N_7930,N_7724,N_7775);
xnor U7931 (N_7931,N_7657,N_7609);
nor U7932 (N_7932,N_7696,N_7792);
and U7933 (N_7933,N_7763,N_7781);
nand U7934 (N_7934,N_7711,N_7681);
and U7935 (N_7935,N_7717,N_7715);
or U7936 (N_7936,N_7637,N_7728);
and U7937 (N_7937,N_7706,N_7674);
nand U7938 (N_7938,N_7666,N_7604);
or U7939 (N_7939,N_7796,N_7639);
and U7940 (N_7940,N_7793,N_7645);
and U7941 (N_7941,N_7710,N_7670);
and U7942 (N_7942,N_7626,N_7685);
and U7943 (N_7943,N_7628,N_7721);
or U7944 (N_7944,N_7697,N_7666);
or U7945 (N_7945,N_7622,N_7637);
and U7946 (N_7946,N_7667,N_7758);
nand U7947 (N_7947,N_7683,N_7622);
nor U7948 (N_7948,N_7769,N_7670);
nor U7949 (N_7949,N_7749,N_7620);
and U7950 (N_7950,N_7695,N_7665);
nor U7951 (N_7951,N_7682,N_7659);
nand U7952 (N_7952,N_7654,N_7603);
or U7953 (N_7953,N_7767,N_7629);
and U7954 (N_7954,N_7716,N_7732);
and U7955 (N_7955,N_7643,N_7733);
nand U7956 (N_7956,N_7622,N_7746);
and U7957 (N_7957,N_7760,N_7748);
nor U7958 (N_7958,N_7731,N_7745);
and U7959 (N_7959,N_7663,N_7761);
or U7960 (N_7960,N_7649,N_7636);
nand U7961 (N_7961,N_7741,N_7614);
and U7962 (N_7962,N_7779,N_7798);
or U7963 (N_7963,N_7617,N_7681);
xnor U7964 (N_7964,N_7679,N_7786);
and U7965 (N_7965,N_7696,N_7649);
xor U7966 (N_7966,N_7735,N_7729);
nand U7967 (N_7967,N_7611,N_7767);
and U7968 (N_7968,N_7720,N_7625);
nand U7969 (N_7969,N_7762,N_7674);
and U7970 (N_7970,N_7670,N_7790);
nand U7971 (N_7971,N_7741,N_7674);
xor U7972 (N_7972,N_7717,N_7670);
nor U7973 (N_7973,N_7604,N_7605);
and U7974 (N_7974,N_7771,N_7674);
nor U7975 (N_7975,N_7752,N_7715);
or U7976 (N_7976,N_7662,N_7702);
nor U7977 (N_7977,N_7680,N_7781);
and U7978 (N_7978,N_7632,N_7761);
nand U7979 (N_7979,N_7770,N_7695);
or U7980 (N_7980,N_7726,N_7618);
xor U7981 (N_7981,N_7681,N_7637);
and U7982 (N_7982,N_7667,N_7766);
nor U7983 (N_7983,N_7718,N_7712);
or U7984 (N_7984,N_7778,N_7792);
nor U7985 (N_7985,N_7688,N_7682);
or U7986 (N_7986,N_7606,N_7729);
and U7987 (N_7987,N_7605,N_7755);
nor U7988 (N_7988,N_7784,N_7748);
nand U7989 (N_7989,N_7676,N_7606);
and U7990 (N_7990,N_7757,N_7797);
or U7991 (N_7991,N_7673,N_7781);
nand U7992 (N_7992,N_7796,N_7717);
nor U7993 (N_7993,N_7784,N_7739);
or U7994 (N_7994,N_7749,N_7606);
and U7995 (N_7995,N_7615,N_7700);
nor U7996 (N_7996,N_7689,N_7612);
nand U7997 (N_7997,N_7781,N_7618);
nor U7998 (N_7998,N_7615,N_7742);
nand U7999 (N_7999,N_7625,N_7645);
nand U8000 (N_8000,N_7955,N_7843);
and U8001 (N_8001,N_7855,N_7967);
nand U8002 (N_8002,N_7889,N_7859);
nor U8003 (N_8003,N_7875,N_7869);
nand U8004 (N_8004,N_7901,N_7835);
or U8005 (N_8005,N_7982,N_7958);
or U8006 (N_8006,N_7913,N_7962);
and U8007 (N_8007,N_7810,N_7910);
or U8008 (N_8008,N_7840,N_7842);
or U8009 (N_8009,N_7872,N_7856);
xnor U8010 (N_8010,N_7919,N_7989);
nor U8011 (N_8011,N_7960,N_7884);
nor U8012 (N_8012,N_7828,N_7905);
nand U8013 (N_8013,N_7801,N_7921);
and U8014 (N_8014,N_7870,N_7871);
or U8015 (N_8015,N_7980,N_7922);
and U8016 (N_8016,N_7914,N_7864);
nor U8017 (N_8017,N_7857,N_7945);
xnor U8018 (N_8018,N_7890,N_7811);
or U8019 (N_8019,N_7839,N_7924);
and U8020 (N_8020,N_7994,N_7819);
or U8021 (N_8021,N_7820,N_7821);
and U8022 (N_8022,N_7966,N_7954);
and U8023 (N_8023,N_7943,N_7888);
or U8024 (N_8024,N_7808,N_7834);
nor U8025 (N_8025,N_7934,N_7918);
and U8026 (N_8026,N_7882,N_7876);
nor U8027 (N_8027,N_7847,N_7813);
or U8028 (N_8028,N_7867,N_7946);
nand U8029 (N_8029,N_7981,N_7825);
and U8030 (N_8030,N_7963,N_7949);
nor U8031 (N_8031,N_7827,N_7833);
nor U8032 (N_8032,N_7902,N_7858);
xor U8033 (N_8033,N_7978,N_7997);
xor U8034 (N_8034,N_7920,N_7831);
nand U8035 (N_8035,N_7817,N_7935);
nand U8036 (N_8036,N_7909,N_7942);
and U8037 (N_8037,N_7937,N_7806);
and U8038 (N_8038,N_7950,N_7933);
or U8039 (N_8039,N_7930,N_7927);
nand U8040 (N_8040,N_7973,N_7939);
nand U8041 (N_8041,N_7908,N_7892);
or U8042 (N_8042,N_7815,N_7826);
and U8043 (N_8043,N_7907,N_7837);
nor U8044 (N_8044,N_7818,N_7932);
nand U8045 (N_8045,N_7986,N_7968);
or U8046 (N_8046,N_7929,N_7800);
and U8047 (N_8047,N_7860,N_7906);
nor U8048 (N_8048,N_7883,N_7990);
nand U8049 (N_8049,N_7915,N_7999);
and U8050 (N_8050,N_7976,N_7879);
nor U8051 (N_8051,N_7987,N_7926);
or U8052 (N_8052,N_7899,N_7970);
and U8053 (N_8053,N_7886,N_7802);
xnor U8054 (N_8054,N_7832,N_7900);
or U8055 (N_8055,N_7851,N_7969);
nand U8056 (N_8056,N_7938,N_7972);
nor U8057 (N_8057,N_7977,N_7911);
or U8058 (N_8058,N_7863,N_7814);
or U8059 (N_8059,N_7894,N_7993);
or U8060 (N_8060,N_7995,N_7885);
nand U8061 (N_8061,N_7931,N_7804);
xor U8062 (N_8062,N_7844,N_7957);
nand U8063 (N_8063,N_7928,N_7865);
nor U8064 (N_8064,N_7936,N_7961);
and U8065 (N_8065,N_7904,N_7984);
and U8066 (N_8066,N_7878,N_7971);
or U8067 (N_8067,N_7898,N_7992);
xor U8068 (N_8068,N_7874,N_7891);
nand U8069 (N_8069,N_7824,N_7956);
nand U8070 (N_8070,N_7948,N_7985);
xnor U8071 (N_8071,N_7893,N_7923);
and U8072 (N_8072,N_7895,N_7916);
nor U8073 (N_8073,N_7809,N_7941);
or U8074 (N_8074,N_7964,N_7841);
nor U8075 (N_8075,N_7836,N_7848);
and U8076 (N_8076,N_7998,N_7880);
nand U8077 (N_8077,N_7965,N_7873);
nor U8078 (N_8078,N_7959,N_7996);
nand U8079 (N_8079,N_7974,N_7897);
nor U8080 (N_8080,N_7979,N_7917);
and U8081 (N_8081,N_7868,N_7854);
nand U8082 (N_8082,N_7877,N_7953);
nand U8083 (N_8083,N_7862,N_7887);
or U8084 (N_8084,N_7991,N_7983);
and U8085 (N_8085,N_7951,N_7925);
xnor U8086 (N_8086,N_7853,N_7896);
or U8087 (N_8087,N_7944,N_7845);
nor U8088 (N_8088,N_7852,N_7988);
nor U8089 (N_8089,N_7807,N_7952);
or U8090 (N_8090,N_7829,N_7903);
xor U8091 (N_8091,N_7838,N_7830);
xnor U8092 (N_8092,N_7805,N_7861);
or U8093 (N_8093,N_7975,N_7822);
and U8094 (N_8094,N_7947,N_7849);
or U8095 (N_8095,N_7912,N_7823);
nand U8096 (N_8096,N_7881,N_7850);
and U8097 (N_8097,N_7803,N_7816);
xnor U8098 (N_8098,N_7866,N_7846);
and U8099 (N_8099,N_7812,N_7940);
nand U8100 (N_8100,N_7952,N_7962);
and U8101 (N_8101,N_7900,N_7861);
or U8102 (N_8102,N_7929,N_7943);
nor U8103 (N_8103,N_7917,N_7853);
nor U8104 (N_8104,N_7801,N_7994);
nor U8105 (N_8105,N_7929,N_7913);
nand U8106 (N_8106,N_7809,N_7913);
or U8107 (N_8107,N_7868,N_7841);
nand U8108 (N_8108,N_7965,N_7800);
and U8109 (N_8109,N_7961,N_7800);
or U8110 (N_8110,N_7956,N_7869);
nand U8111 (N_8111,N_7942,N_7978);
or U8112 (N_8112,N_7860,N_7966);
and U8113 (N_8113,N_7839,N_7889);
or U8114 (N_8114,N_7935,N_7866);
xnor U8115 (N_8115,N_7933,N_7809);
nand U8116 (N_8116,N_7904,N_7913);
and U8117 (N_8117,N_7955,N_7823);
nor U8118 (N_8118,N_7825,N_7916);
nand U8119 (N_8119,N_7837,N_7949);
and U8120 (N_8120,N_7984,N_7840);
xor U8121 (N_8121,N_7975,N_7903);
nor U8122 (N_8122,N_7980,N_7872);
nand U8123 (N_8123,N_7812,N_7855);
xnor U8124 (N_8124,N_7886,N_7881);
nor U8125 (N_8125,N_7854,N_7836);
nand U8126 (N_8126,N_7891,N_7824);
nand U8127 (N_8127,N_7935,N_7912);
nand U8128 (N_8128,N_7944,N_7809);
and U8129 (N_8129,N_7894,N_7826);
and U8130 (N_8130,N_7989,N_7885);
and U8131 (N_8131,N_7963,N_7896);
and U8132 (N_8132,N_7897,N_7968);
and U8133 (N_8133,N_7965,N_7980);
nand U8134 (N_8134,N_7845,N_7812);
nor U8135 (N_8135,N_7956,N_7811);
nor U8136 (N_8136,N_7819,N_7990);
and U8137 (N_8137,N_7883,N_7959);
or U8138 (N_8138,N_7883,N_7885);
nor U8139 (N_8139,N_7958,N_7970);
or U8140 (N_8140,N_7855,N_7971);
or U8141 (N_8141,N_7996,N_7938);
nor U8142 (N_8142,N_7970,N_7947);
nor U8143 (N_8143,N_7882,N_7804);
nor U8144 (N_8144,N_7848,N_7814);
nor U8145 (N_8145,N_7884,N_7870);
and U8146 (N_8146,N_7921,N_7901);
xor U8147 (N_8147,N_7854,N_7990);
and U8148 (N_8148,N_7952,N_7827);
nand U8149 (N_8149,N_7979,N_7941);
nand U8150 (N_8150,N_7899,N_7967);
or U8151 (N_8151,N_7831,N_7855);
xnor U8152 (N_8152,N_7805,N_7858);
nand U8153 (N_8153,N_7818,N_7940);
or U8154 (N_8154,N_7964,N_7838);
and U8155 (N_8155,N_7869,N_7824);
and U8156 (N_8156,N_7821,N_7877);
and U8157 (N_8157,N_7880,N_7994);
or U8158 (N_8158,N_7874,N_7837);
nand U8159 (N_8159,N_7945,N_7950);
nand U8160 (N_8160,N_7921,N_7858);
xnor U8161 (N_8161,N_7907,N_7923);
or U8162 (N_8162,N_7972,N_7828);
nand U8163 (N_8163,N_7832,N_7918);
nor U8164 (N_8164,N_7817,N_7949);
or U8165 (N_8165,N_7852,N_7879);
xor U8166 (N_8166,N_7835,N_7874);
nand U8167 (N_8167,N_7888,N_7866);
or U8168 (N_8168,N_7805,N_7863);
nand U8169 (N_8169,N_7906,N_7827);
nor U8170 (N_8170,N_7945,N_7830);
or U8171 (N_8171,N_7825,N_7996);
nand U8172 (N_8172,N_7853,N_7860);
nand U8173 (N_8173,N_7804,N_7989);
nor U8174 (N_8174,N_7836,N_7905);
or U8175 (N_8175,N_7890,N_7969);
or U8176 (N_8176,N_7834,N_7858);
and U8177 (N_8177,N_7967,N_7947);
nand U8178 (N_8178,N_7841,N_7826);
and U8179 (N_8179,N_7933,N_7826);
nand U8180 (N_8180,N_7913,N_7902);
nor U8181 (N_8181,N_7997,N_7926);
xor U8182 (N_8182,N_7985,N_7951);
xor U8183 (N_8183,N_7801,N_7813);
nand U8184 (N_8184,N_7956,N_7862);
and U8185 (N_8185,N_7998,N_7984);
nor U8186 (N_8186,N_7843,N_7815);
or U8187 (N_8187,N_7813,N_7902);
and U8188 (N_8188,N_7855,N_7981);
and U8189 (N_8189,N_7936,N_7827);
and U8190 (N_8190,N_7896,N_7805);
nand U8191 (N_8191,N_7851,N_7965);
nor U8192 (N_8192,N_7916,N_7802);
nor U8193 (N_8193,N_7882,N_7917);
nor U8194 (N_8194,N_7938,N_7819);
and U8195 (N_8195,N_7841,N_7894);
nor U8196 (N_8196,N_7960,N_7867);
and U8197 (N_8197,N_7982,N_7983);
or U8198 (N_8198,N_7880,N_7850);
nor U8199 (N_8199,N_7984,N_7886);
nand U8200 (N_8200,N_8071,N_8117);
nor U8201 (N_8201,N_8018,N_8128);
nor U8202 (N_8202,N_8145,N_8051);
and U8203 (N_8203,N_8195,N_8199);
and U8204 (N_8204,N_8036,N_8008);
xnor U8205 (N_8205,N_8026,N_8092);
nand U8206 (N_8206,N_8037,N_8108);
or U8207 (N_8207,N_8140,N_8028);
nand U8208 (N_8208,N_8144,N_8047);
nand U8209 (N_8209,N_8127,N_8001);
and U8210 (N_8210,N_8107,N_8084);
nand U8211 (N_8211,N_8073,N_8049);
or U8212 (N_8212,N_8087,N_8134);
nor U8213 (N_8213,N_8136,N_8115);
nor U8214 (N_8214,N_8017,N_8033);
or U8215 (N_8215,N_8014,N_8074);
or U8216 (N_8216,N_8160,N_8039);
and U8217 (N_8217,N_8067,N_8152);
and U8218 (N_8218,N_8198,N_8006);
nand U8219 (N_8219,N_8041,N_8110);
nor U8220 (N_8220,N_8129,N_8002);
nor U8221 (N_8221,N_8019,N_8054);
xnor U8222 (N_8222,N_8161,N_8013);
and U8223 (N_8223,N_8099,N_8125);
or U8224 (N_8224,N_8076,N_8095);
nor U8225 (N_8225,N_8097,N_8162);
nor U8226 (N_8226,N_8090,N_8101);
and U8227 (N_8227,N_8089,N_8122);
or U8228 (N_8228,N_8082,N_8086);
and U8229 (N_8229,N_8011,N_8070);
or U8230 (N_8230,N_8126,N_8069);
and U8231 (N_8231,N_8009,N_8171);
nor U8232 (N_8232,N_8148,N_8046);
and U8233 (N_8233,N_8159,N_8100);
or U8234 (N_8234,N_8029,N_8179);
or U8235 (N_8235,N_8055,N_8177);
or U8236 (N_8236,N_8163,N_8170);
and U8237 (N_8237,N_8143,N_8147);
and U8238 (N_8238,N_8175,N_8061);
and U8239 (N_8239,N_8053,N_8156);
or U8240 (N_8240,N_8158,N_8135);
and U8241 (N_8241,N_8112,N_8155);
and U8242 (N_8242,N_8080,N_8141);
nor U8243 (N_8243,N_8012,N_8000);
and U8244 (N_8244,N_8058,N_8088);
or U8245 (N_8245,N_8094,N_8178);
nand U8246 (N_8246,N_8114,N_8131);
nand U8247 (N_8247,N_8188,N_8075);
nor U8248 (N_8248,N_8166,N_8121);
nand U8249 (N_8249,N_8120,N_8103);
or U8250 (N_8250,N_8169,N_8035);
nor U8251 (N_8251,N_8190,N_8016);
and U8252 (N_8252,N_8007,N_8176);
nor U8253 (N_8253,N_8106,N_8072);
nand U8254 (N_8254,N_8068,N_8015);
or U8255 (N_8255,N_8124,N_8042);
or U8256 (N_8256,N_8123,N_8185);
and U8257 (N_8257,N_8081,N_8174);
or U8258 (N_8258,N_8146,N_8192);
nand U8259 (N_8259,N_8193,N_8184);
or U8260 (N_8260,N_8023,N_8142);
xnor U8261 (N_8261,N_8077,N_8083);
or U8262 (N_8262,N_8091,N_8196);
or U8263 (N_8263,N_8064,N_8109);
nor U8264 (N_8264,N_8181,N_8021);
or U8265 (N_8265,N_8048,N_8062);
nand U8266 (N_8266,N_8032,N_8025);
xnor U8267 (N_8267,N_8183,N_8005);
xnor U8268 (N_8268,N_8057,N_8104);
nand U8269 (N_8269,N_8186,N_8003);
and U8270 (N_8270,N_8105,N_8022);
and U8271 (N_8271,N_8085,N_8189);
nand U8272 (N_8272,N_8132,N_8024);
and U8273 (N_8273,N_8004,N_8167);
xnor U8274 (N_8274,N_8034,N_8187);
and U8275 (N_8275,N_8157,N_8096);
xnor U8276 (N_8276,N_8038,N_8044);
and U8277 (N_8277,N_8079,N_8027);
and U8278 (N_8278,N_8040,N_8113);
nand U8279 (N_8279,N_8045,N_8139);
nor U8280 (N_8280,N_8031,N_8150);
or U8281 (N_8281,N_8066,N_8116);
and U8282 (N_8282,N_8111,N_8133);
and U8283 (N_8283,N_8102,N_8020);
xnor U8284 (N_8284,N_8165,N_8078);
nand U8285 (N_8285,N_8098,N_8153);
nand U8286 (N_8286,N_8093,N_8149);
and U8287 (N_8287,N_8197,N_8060);
nand U8288 (N_8288,N_8043,N_8063);
nand U8289 (N_8289,N_8137,N_8056);
nand U8290 (N_8290,N_8173,N_8194);
or U8291 (N_8291,N_8154,N_8050);
nor U8292 (N_8292,N_8130,N_8052);
nor U8293 (N_8293,N_8118,N_8182);
nor U8294 (N_8294,N_8059,N_8138);
nand U8295 (N_8295,N_8151,N_8010);
nor U8296 (N_8296,N_8191,N_8168);
nand U8297 (N_8297,N_8172,N_8065);
nand U8298 (N_8298,N_8119,N_8164);
and U8299 (N_8299,N_8180,N_8030);
and U8300 (N_8300,N_8134,N_8197);
and U8301 (N_8301,N_8021,N_8157);
nor U8302 (N_8302,N_8030,N_8074);
or U8303 (N_8303,N_8079,N_8092);
and U8304 (N_8304,N_8166,N_8052);
or U8305 (N_8305,N_8195,N_8099);
xnor U8306 (N_8306,N_8169,N_8193);
nor U8307 (N_8307,N_8084,N_8056);
and U8308 (N_8308,N_8023,N_8127);
and U8309 (N_8309,N_8076,N_8130);
nand U8310 (N_8310,N_8016,N_8008);
nand U8311 (N_8311,N_8124,N_8056);
nand U8312 (N_8312,N_8013,N_8146);
nor U8313 (N_8313,N_8161,N_8023);
or U8314 (N_8314,N_8089,N_8187);
nand U8315 (N_8315,N_8184,N_8024);
or U8316 (N_8316,N_8104,N_8194);
nand U8317 (N_8317,N_8089,N_8177);
and U8318 (N_8318,N_8130,N_8142);
or U8319 (N_8319,N_8147,N_8087);
and U8320 (N_8320,N_8018,N_8010);
nor U8321 (N_8321,N_8022,N_8083);
and U8322 (N_8322,N_8171,N_8092);
nor U8323 (N_8323,N_8000,N_8112);
xor U8324 (N_8324,N_8057,N_8016);
nand U8325 (N_8325,N_8017,N_8073);
or U8326 (N_8326,N_8154,N_8111);
nand U8327 (N_8327,N_8093,N_8087);
nand U8328 (N_8328,N_8046,N_8047);
nor U8329 (N_8329,N_8055,N_8114);
and U8330 (N_8330,N_8077,N_8026);
nor U8331 (N_8331,N_8008,N_8050);
xor U8332 (N_8332,N_8101,N_8102);
nand U8333 (N_8333,N_8008,N_8068);
nor U8334 (N_8334,N_8041,N_8073);
nor U8335 (N_8335,N_8114,N_8062);
and U8336 (N_8336,N_8103,N_8038);
xnor U8337 (N_8337,N_8066,N_8082);
xor U8338 (N_8338,N_8104,N_8183);
and U8339 (N_8339,N_8099,N_8171);
or U8340 (N_8340,N_8034,N_8076);
nand U8341 (N_8341,N_8039,N_8058);
nor U8342 (N_8342,N_8143,N_8096);
nand U8343 (N_8343,N_8081,N_8180);
and U8344 (N_8344,N_8064,N_8145);
and U8345 (N_8345,N_8102,N_8012);
nor U8346 (N_8346,N_8050,N_8029);
nand U8347 (N_8347,N_8147,N_8145);
and U8348 (N_8348,N_8050,N_8026);
and U8349 (N_8349,N_8069,N_8096);
nor U8350 (N_8350,N_8057,N_8190);
nand U8351 (N_8351,N_8185,N_8044);
nand U8352 (N_8352,N_8071,N_8143);
or U8353 (N_8353,N_8132,N_8141);
xor U8354 (N_8354,N_8173,N_8145);
nor U8355 (N_8355,N_8190,N_8086);
or U8356 (N_8356,N_8109,N_8166);
nor U8357 (N_8357,N_8075,N_8149);
or U8358 (N_8358,N_8191,N_8120);
and U8359 (N_8359,N_8155,N_8165);
or U8360 (N_8360,N_8153,N_8083);
nand U8361 (N_8361,N_8023,N_8095);
and U8362 (N_8362,N_8038,N_8050);
or U8363 (N_8363,N_8031,N_8070);
or U8364 (N_8364,N_8057,N_8108);
nor U8365 (N_8365,N_8047,N_8043);
or U8366 (N_8366,N_8042,N_8012);
nor U8367 (N_8367,N_8069,N_8002);
nor U8368 (N_8368,N_8121,N_8097);
nor U8369 (N_8369,N_8039,N_8183);
nor U8370 (N_8370,N_8013,N_8188);
xor U8371 (N_8371,N_8093,N_8173);
nand U8372 (N_8372,N_8015,N_8091);
and U8373 (N_8373,N_8192,N_8013);
or U8374 (N_8374,N_8038,N_8068);
or U8375 (N_8375,N_8047,N_8053);
and U8376 (N_8376,N_8026,N_8083);
xnor U8377 (N_8377,N_8025,N_8002);
or U8378 (N_8378,N_8173,N_8142);
nand U8379 (N_8379,N_8098,N_8038);
xnor U8380 (N_8380,N_8101,N_8153);
or U8381 (N_8381,N_8057,N_8153);
and U8382 (N_8382,N_8194,N_8031);
and U8383 (N_8383,N_8106,N_8039);
nand U8384 (N_8384,N_8168,N_8011);
and U8385 (N_8385,N_8170,N_8181);
and U8386 (N_8386,N_8140,N_8155);
or U8387 (N_8387,N_8041,N_8109);
or U8388 (N_8388,N_8051,N_8072);
nor U8389 (N_8389,N_8130,N_8116);
nand U8390 (N_8390,N_8181,N_8135);
nor U8391 (N_8391,N_8069,N_8016);
nor U8392 (N_8392,N_8138,N_8127);
nor U8393 (N_8393,N_8072,N_8055);
nand U8394 (N_8394,N_8134,N_8055);
and U8395 (N_8395,N_8017,N_8099);
nand U8396 (N_8396,N_8030,N_8122);
xnor U8397 (N_8397,N_8073,N_8053);
nor U8398 (N_8398,N_8189,N_8065);
and U8399 (N_8399,N_8197,N_8029);
nand U8400 (N_8400,N_8221,N_8269);
and U8401 (N_8401,N_8380,N_8251);
nor U8402 (N_8402,N_8260,N_8206);
nor U8403 (N_8403,N_8285,N_8200);
and U8404 (N_8404,N_8369,N_8204);
nor U8405 (N_8405,N_8334,N_8265);
or U8406 (N_8406,N_8388,N_8348);
nor U8407 (N_8407,N_8313,N_8398);
nor U8408 (N_8408,N_8223,N_8248);
nand U8409 (N_8409,N_8328,N_8362);
or U8410 (N_8410,N_8232,N_8335);
and U8411 (N_8411,N_8214,N_8235);
and U8412 (N_8412,N_8297,N_8366);
or U8413 (N_8413,N_8257,N_8290);
nand U8414 (N_8414,N_8360,N_8311);
or U8415 (N_8415,N_8300,N_8296);
and U8416 (N_8416,N_8222,N_8233);
nand U8417 (N_8417,N_8294,N_8263);
nor U8418 (N_8418,N_8386,N_8322);
nor U8419 (N_8419,N_8371,N_8215);
nor U8420 (N_8420,N_8308,N_8341);
or U8421 (N_8421,N_8319,N_8318);
xor U8422 (N_8422,N_8320,N_8342);
nor U8423 (N_8423,N_8270,N_8337);
or U8424 (N_8424,N_8391,N_8310);
and U8425 (N_8425,N_8306,N_8346);
nand U8426 (N_8426,N_8280,N_8385);
nand U8427 (N_8427,N_8379,N_8262);
xnor U8428 (N_8428,N_8228,N_8317);
and U8429 (N_8429,N_8253,N_8392);
and U8430 (N_8430,N_8340,N_8329);
and U8431 (N_8431,N_8275,N_8227);
nor U8432 (N_8432,N_8396,N_8286);
or U8433 (N_8433,N_8243,N_8315);
xnor U8434 (N_8434,N_8343,N_8301);
nand U8435 (N_8435,N_8210,N_8247);
nor U8436 (N_8436,N_8212,N_8330);
or U8437 (N_8437,N_8220,N_8283);
or U8438 (N_8438,N_8273,N_8378);
or U8439 (N_8439,N_8332,N_8229);
nand U8440 (N_8440,N_8254,N_8207);
and U8441 (N_8441,N_8325,N_8327);
and U8442 (N_8442,N_8305,N_8359);
nor U8443 (N_8443,N_8356,N_8357);
and U8444 (N_8444,N_8338,N_8287);
and U8445 (N_8445,N_8234,N_8373);
nor U8446 (N_8446,N_8365,N_8244);
nor U8447 (N_8447,N_8231,N_8339);
nor U8448 (N_8448,N_8397,N_8226);
nand U8449 (N_8449,N_8303,N_8237);
and U8450 (N_8450,N_8390,N_8271);
nor U8451 (N_8451,N_8213,N_8321);
nand U8452 (N_8452,N_8208,N_8238);
xor U8453 (N_8453,N_8304,N_8282);
nor U8454 (N_8454,N_8268,N_8389);
nand U8455 (N_8455,N_8384,N_8224);
nand U8456 (N_8456,N_8250,N_8395);
or U8457 (N_8457,N_8381,N_8347);
nand U8458 (N_8458,N_8218,N_8387);
nand U8459 (N_8459,N_8267,N_8350);
nand U8460 (N_8460,N_8364,N_8225);
and U8461 (N_8461,N_8331,N_8324);
and U8462 (N_8462,N_8230,N_8323);
nand U8463 (N_8463,N_8284,N_8393);
or U8464 (N_8464,N_8370,N_8363);
or U8465 (N_8465,N_8399,N_8292);
nand U8466 (N_8466,N_8372,N_8349);
or U8467 (N_8467,N_8358,N_8314);
and U8468 (N_8468,N_8295,N_8246);
or U8469 (N_8469,N_8368,N_8376);
or U8470 (N_8470,N_8236,N_8291);
or U8471 (N_8471,N_8316,N_8361);
nor U8472 (N_8472,N_8377,N_8255);
nand U8473 (N_8473,N_8383,N_8279);
nand U8474 (N_8474,N_8276,N_8245);
or U8475 (N_8475,N_8205,N_8307);
or U8476 (N_8476,N_8293,N_8374);
nor U8477 (N_8477,N_8394,N_8256);
nor U8478 (N_8478,N_8239,N_8266);
nand U8479 (N_8479,N_8289,N_8258);
or U8480 (N_8480,N_8259,N_8203);
nand U8481 (N_8481,N_8274,N_8252);
nand U8482 (N_8482,N_8375,N_8355);
or U8483 (N_8483,N_8367,N_8272);
nand U8484 (N_8484,N_8298,N_8242);
nand U8485 (N_8485,N_8240,N_8299);
nor U8486 (N_8486,N_8261,N_8344);
xnor U8487 (N_8487,N_8241,N_8249);
or U8488 (N_8488,N_8216,N_8302);
or U8489 (N_8489,N_8211,N_8353);
or U8490 (N_8490,N_8209,N_8333);
or U8491 (N_8491,N_8352,N_8219);
nand U8492 (N_8492,N_8345,N_8277);
nor U8493 (N_8493,N_8202,N_8354);
or U8494 (N_8494,N_8312,N_8288);
nand U8495 (N_8495,N_8336,N_8281);
nand U8496 (N_8496,N_8201,N_8278);
or U8497 (N_8497,N_8351,N_8309);
nand U8498 (N_8498,N_8382,N_8326);
and U8499 (N_8499,N_8264,N_8217);
or U8500 (N_8500,N_8370,N_8206);
nand U8501 (N_8501,N_8360,N_8215);
nor U8502 (N_8502,N_8322,N_8302);
or U8503 (N_8503,N_8347,N_8262);
nand U8504 (N_8504,N_8234,N_8389);
or U8505 (N_8505,N_8262,N_8392);
xnor U8506 (N_8506,N_8364,N_8367);
and U8507 (N_8507,N_8253,N_8284);
nand U8508 (N_8508,N_8207,N_8375);
nand U8509 (N_8509,N_8243,N_8277);
or U8510 (N_8510,N_8380,N_8258);
nor U8511 (N_8511,N_8221,N_8371);
nor U8512 (N_8512,N_8300,N_8323);
nand U8513 (N_8513,N_8229,N_8330);
nor U8514 (N_8514,N_8200,N_8289);
and U8515 (N_8515,N_8282,N_8318);
nand U8516 (N_8516,N_8297,N_8290);
or U8517 (N_8517,N_8316,N_8303);
and U8518 (N_8518,N_8264,N_8368);
and U8519 (N_8519,N_8275,N_8252);
and U8520 (N_8520,N_8206,N_8286);
nand U8521 (N_8521,N_8344,N_8207);
or U8522 (N_8522,N_8272,N_8386);
and U8523 (N_8523,N_8303,N_8366);
nor U8524 (N_8524,N_8326,N_8315);
nor U8525 (N_8525,N_8321,N_8222);
and U8526 (N_8526,N_8214,N_8360);
and U8527 (N_8527,N_8271,N_8306);
or U8528 (N_8528,N_8243,N_8213);
and U8529 (N_8529,N_8394,N_8230);
nor U8530 (N_8530,N_8391,N_8335);
or U8531 (N_8531,N_8388,N_8394);
and U8532 (N_8532,N_8275,N_8338);
nand U8533 (N_8533,N_8383,N_8264);
or U8534 (N_8534,N_8366,N_8374);
or U8535 (N_8535,N_8244,N_8277);
nor U8536 (N_8536,N_8298,N_8232);
xnor U8537 (N_8537,N_8213,N_8365);
or U8538 (N_8538,N_8231,N_8212);
nand U8539 (N_8539,N_8225,N_8359);
nand U8540 (N_8540,N_8236,N_8257);
nor U8541 (N_8541,N_8330,N_8312);
nand U8542 (N_8542,N_8355,N_8395);
or U8543 (N_8543,N_8270,N_8382);
and U8544 (N_8544,N_8349,N_8352);
nand U8545 (N_8545,N_8372,N_8334);
or U8546 (N_8546,N_8271,N_8304);
or U8547 (N_8547,N_8363,N_8336);
or U8548 (N_8548,N_8304,N_8207);
nand U8549 (N_8549,N_8363,N_8302);
or U8550 (N_8550,N_8221,N_8218);
nand U8551 (N_8551,N_8367,N_8334);
nor U8552 (N_8552,N_8284,N_8392);
nor U8553 (N_8553,N_8237,N_8375);
or U8554 (N_8554,N_8352,N_8369);
nor U8555 (N_8555,N_8210,N_8319);
nand U8556 (N_8556,N_8261,N_8340);
or U8557 (N_8557,N_8257,N_8390);
and U8558 (N_8558,N_8264,N_8258);
or U8559 (N_8559,N_8223,N_8353);
nor U8560 (N_8560,N_8279,N_8309);
or U8561 (N_8561,N_8237,N_8225);
xor U8562 (N_8562,N_8322,N_8332);
and U8563 (N_8563,N_8354,N_8301);
nand U8564 (N_8564,N_8229,N_8239);
nor U8565 (N_8565,N_8387,N_8326);
nor U8566 (N_8566,N_8237,N_8227);
or U8567 (N_8567,N_8380,N_8373);
or U8568 (N_8568,N_8340,N_8278);
nor U8569 (N_8569,N_8355,N_8275);
or U8570 (N_8570,N_8278,N_8205);
and U8571 (N_8571,N_8232,N_8268);
or U8572 (N_8572,N_8362,N_8348);
and U8573 (N_8573,N_8226,N_8257);
or U8574 (N_8574,N_8261,N_8294);
nand U8575 (N_8575,N_8333,N_8326);
nand U8576 (N_8576,N_8316,N_8334);
and U8577 (N_8577,N_8283,N_8377);
or U8578 (N_8578,N_8217,N_8293);
xor U8579 (N_8579,N_8315,N_8383);
or U8580 (N_8580,N_8257,N_8302);
nor U8581 (N_8581,N_8377,N_8304);
and U8582 (N_8582,N_8316,N_8258);
and U8583 (N_8583,N_8209,N_8352);
or U8584 (N_8584,N_8305,N_8207);
and U8585 (N_8585,N_8331,N_8307);
xor U8586 (N_8586,N_8397,N_8220);
or U8587 (N_8587,N_8255,N_8231);
nand U8588 (N_8588,N_8366,N_8272);
or U8589 (N_8589,N_8383,N_8378);
nand U8590 (N_8590,N_8299,N_8224);
or U8591 (N_8591,N_8306,N_8246);
and U8592 (N_8592,N_8310,N_8280);
nand U8593 (N_8593,N_8320,N_8226);
nor U8594 (N_8594,N_8369,N_8264);
and U8595 (N_8595,N_8269,N_8279);
or U8596 (N_8596,N_8388,N_8362);
or U8597 (N_8597,N_8301,N_8242);
and U8598 (N_8598,N_8380,N_8330);
and U8599 (N_8599,N_8394,N_8298);
nand U8600 (N_8600,N_8469,N_8432);
nand U8601 (N_8601,N_8477,N_8445);
nand U8602 (N_8602,N_8576,N_8535);
xor U8603 (N_8603,N_8541,N_8454);
nor U8604 (N_8604,N_8404,N_8507);
and U8605 (N_8605,N_8510,N_8441);
nor U8606 (N_8606,N_8482,N_8470);
nand U8607 (N_8607,N_8557,N_8409);
or U8608 (N_8608,N_8542,N_8419);
and U8609 (N_8609,N_8460,N_8439);
nor U8610 (N_8610,N_8586,N_8570);
nand U8611 (N_8611,N_8580,N_8564);
nand U8612 (N_8612,N_8483,N_8485);
nand U8613 (N_8613,N_8559,N_8591);
nor U8614 (N_8614,N_8436,N_8598);
nor U8615 (N_8615,N_8501,N_8506);
or U8616 (N_8616,N_8571,N_8514);
and U8617 (N_8617,N_8426,N_8400);
nand U8618 (N_8618,N_8408,N_8446);
nor U8619 (N_8619,N_8547,N_8498);
nand U8620 (N_8620,N_8462,N_8548);
xor U8621 (N_8621,N_8471,N_8539);
and U8622 (N_8622,N_8573,N_8488);
xor U8623 (N_8623,N_8447,N_8588);
or U8624 (N_8624,N_8517,N_8556);
xnor U8625 (N_8625,N_8518,N_8582);
nand U8626 (N_8626,N_8533,N_8508);
nor U8627 (N_8627,N_8414,N_8532);
or U8628 (N_8628,N_8560,N_8512);
and U8629 (N_8629,N_8401,N_8458);
and U8630 (N_8630,N_8567,N_8599);
nand U8631 (N_8631,N_8420,N_8523);
nand U8632 (N_8632,N_8428,N_8467);
nor U8633 (N_8633,N_8421,N_8534);
and U8634 (N_8634,N_8527,N_8417);
xor U8635 (N_8635,N_8451,N_8522);
xnor U8636 (N_8636,N_8424,N_8457);
or U8637 (N_8637,N_8497,N_8434);
nand U8638 (N_8638,N_8475,N_8511);
nor U8639 (N_8639,N_8415,N_8438);
nor U8640 (N_8640,N_8416,N_8587);
and U8641 (N_8641,N_8526,N_8450);
nand U8642 (N_8642,N_8545,N_8544);
nand U8643 (N_8643,N_8551,N_8558);
xnor U8644 (N_8644,N_8524,N_8521);
nor U8645 (N_8645,N_8405,N_8466);
nand U8646 (N_8646,N_8442,N_8538);
or U8647 (N_8647,N_8464,N_8569);
and U8648 (N_8648,N_8499,N_8520);
nor U8649 (N_8649,N_8537,N_8515);
xor U8650 (N_8650,N_8490,N_8500);
and U8651 (N_8651,N_8423,N_8562);
or U8652 (N_8652,N_8584,N_8430);
nand U8653 (N_8653,N_8554,N_8592);
nor U8654 (N_8654,N_8536,N_8516);
and U8655 (N_8655,N_8581,N_8585);
nor U8656 (N_8656,N_8481,N_8449);
and U8657 (N_8657,N_8444,N_8473);
or U8658 (N_8658,N_8410,N_8504);
or U8659 (N_8659,N_8465,N_8577);
nor U8660 (N_8660,N_8566,N_8412);
and U8661 (N_8661,N_8595,N_8452);
nand U8662 (N_8662,N_8578,N_8509);
or U8663 (N_8663,N_8583,N_8574);
nand U8664 (N_8664,N_8406,N_8572);
xor U8665 (N_8665,N_8596,N_8494);
or U8666 (N_8666,N_8448,N_8463);
nor U8667 (N_8667,N_8443,N_8429);
or U8668 (N_8668,N_8502,N_8403);
and U8669 (N_8669,N_8435,N_8505);
nor U8670 (N_8670,N_8402,N_8540);
and U8671 (N_8671,N_8422,N_8552);
nand U8672 (N_8672,N_8553,N_8597);
nand U8673 (N_8673,N_8525,N_8487);
or U8674 (N_8674,N_8461,N_8486);
nand U8675 (N_8675,N_8484,N_8550);
or U8676 (N_8676,N_8549,N_8593);
or U8677 (N_8677,N_8433,N_8575);
nand U8678 (N_8678,N_8489,N_8479);
and U8679 (N_8679,N_8480,N_8529);
and U8680 (N_8680,N_8468,N_8427);
or U8681 (N_8681,N_8546,N_8418);
nor U8682 (N_8682,N_8495,N_8568);
nor U8683 (N_8683,N_8472,N_8425);
xnor U8684 (N_8684,N_8456,N_8503);
xor U8685 (N_8685,N_8459,N_8543);
nor U8686 (N_8686,N_8513,N_8519);
or U8687 (N_8687,N_8493,N_8437);
nand U8688 (N_8688,N_8589,N_8440);
and U8689 (N_8689,N_8431,N_8579);
xnor U8690 (N_8690,N_8530,N_8478);
nand U8691 (N_8691,N_8455,N_8413);
or U8692 (N_8692,N_8565,N_8411);
nand U8693 (N_8693,N_8492,N_8496);
nand U8694 (N_8694,N_8476,N_8474);
xor U8695 (N_8695,N_8528,N_8594);
and U8696 (N_8696,N_8407,N_8531);
or U8697 (N_8697,N_8563,N_8453);
and U8698 (N_8698,N_8491,N_8555);
and U8699 (N_8699,N_8561,N_8590);
nor U8700 (N_8700,N_8585,N_8461);
nor U8701 (N_8701,N_8493,N_8453);
nand U8702 (N_8702,N_8524,N_8559);
nand U8703 (N_8703,N_8443,N_8536);
and U8704 (N_8704,N_8416,N_8442);
xor U8705 (N_8705,N_8429,N_8423);
nand U8706 (N_8706,N_8572,N_8446);
nand U8707 (N_8707,N_8543,N_8405);
or U8708 (N_8708,N_8514,N_8565);
nand U8709 (N_8709,N_8444,N_8515);
nand U8710 (N_8710,N_8507,N_8426);
nor U8711 (N_8711,N_8531,N_8447);
nor U8712 (N_8712,N_8503,N_8488);
nand U8713 (N_8713,N_8511,N_8592);
or U8714 (N_8714,N_8597,N_8479);
and U8715 (N_8715,N_8415,N_8505);
xnor U8716 (N_8716,N_8416,N_8412);
and U8717 (N_8717,N_8514,N_8467);
nor U8718 (N_8718,N_8449,N_8494);
and U8719 (N_8719,N_8490,N_8433);
or U8720 (N_8720,N_8405,N_8419);
or U8721 (N_8721,N_8445,N_8594);
or U8722 (N_8722,N_8522,N_8474);
nand U8723 (N_8723,N_8531,N_8448);
or U8724 (N_8724,N_8426,N_8479);
nand U8725 (N_8725,N_8493,N_8465);
and U8726 (N_8726,N_8580,N_8431);
and U8727 (N_8727,N_8442,N_8524);
or U8728 (N_8728,N_8571,N_8445);
and U8729 (N_8729,N_8420,N_8492);
xnor U8730 (N_8730,N_8416,N_8491);
nand U8731 (N_8731,N_8475,N_8501);
and U8732 (N_8732,N_8585,N_8529);
nand U8733 (N_8733,N_8463,N_8430);
and U8734 (N_8734,N_8480,N_8463);
or U8735 (N_8735,N_8582,N_8505);
or U8736 (N_8736,N_8403,N_8551);
or U8737 (N_8737,N_8456,N_8532);
xor U8738 (N_8738,N_8477,N_8536);
or U8739 (N_8739,N_8478,N_8580);
nor U8740 (N_8740,N_8462,N_8584);
nand U8741 (N_8741,N_8552,N_8441);
nand U8742 (N_8742,N_8543,N_8458);
or U8743 (N_8743,N_8416,N_8488);
and U8744 (N_8744,N_8463,N_8522);
or U8745 (N_8745,N_8582,N_8586);
or U8746 (N_8746,N_8511,N_8588);
nand U8747 (N_8747,N_8425,N_8413);
nor U8748 (N_8748,N_8464,N_8577);
nand U8749 (N_8749,N_8499,N_8488);
and U8750 (N_8750,N_8436,N_8470);
nand U8751 (N_8751,N_8404,N_8523);
and U8752 (N_8752,N_8411,N_8452);
nor U8753 (N_8753,N_8429,N_8523);
nor U8754 (N_8754,N_8525,N_8473);
or U8755 (N_8755,N_8559,N_8534);
and U8756 (N_8756,N_8463,N_8589);
nor U8757 (N_8757,N_8414,N_8582);
xor U8758 (N_8758,N_8571,N_8498);
nor U8759 (N_8759,N_8598,N_8418);
or U8760 (N_8760,N_8437,N_8480);
nor U8761 (N_8761,N_8472,N_8439);
and U8762 (N_8762,N_8581,N_8440);
nor U8763 (N_8763,N_8505,N_8593);
and U8764 (N_8764,N_8412,N_8557);
nor U8765 (N_8765,N_8542,N_8428);
nand U8766 (N_8766,N_8559,N_8595);
or U8767 (N_8767,N_8566,N_8502);
nor U8768 (N_8768,N_8518,N_8461);
or U8769 (N_8769,N_8400,N_8554);
and U8770 (N_8770,N_8486,N_8533);
nor U8771 (N_8771,N_8581,N_8527);
and U8772 (N_8772,N_8476,N_8417);
nor U8773 (N_8773,N_8591,N_8401);
nand U8774 (N_8774,N_8594,N_8486);
and U8775 (N_8775,N_8414,N_8444);
and U8776 (N_8776,N_8421,N_8404);
nor U8777 (N_8777,N_8581,N_8587);
or U8778 (N_8778,N_8532,N_8440);
nand U8779 (N_8779,N_8451,N_8488);
nand U8780 (N_8780,N_8486,N_8503);
nor U8781 (N_8781,N_8454,N_8406);
nor U8782 (N_8782,N_8465,N_8536);
nand U8783 (N_8783,N_8557,N_8581);
nand U8784 (N_8784,N_8586,N_8537);
nor U8785 (N_8785,N_8565,N_8450);
and U8786 (N_8786,N_8480,N_8499);
and U8787 (N_8787,N_8548,N_8450);
or U8788 (N_8788,N_8450,N_8409);
nor U8789 (N_8789,N_8415,N_8531);
and U8790 (N_8790,N_8563,N_8597);
or U8791 (N_8791,N_8550,N_8516);
and U8792 (N_8792,N_8489,N_8525);
and U8793 (N_8793,N_8439,N_8486);
nor U8794 (N_8794,N_8406,N_8539);
nor U8795 (N_8795,N_8473,N_8466);
nor U8796 (N_8796,N_8453,N_8424);
xor U8797 (N_8797,N_8449,N_8513);
or U8798 (N_8798,N_8522,N_8490);
nand U8799 (N_8799,N_8552,N_8541);
and U8800 (N_8800,N_8713,N_8659);
nor U8801 (N_8801,N_8791,N_8660);
or U8802 (N_8802,N_8663,N_8619);
xnor U8803 (N_8803,N_8750,N_8722);
nand U8804 (N_8804,N_8754,N_8741);
xor U8805 (N_8805,N_8773,N_8796);
and U8806 (N_8806,N_8744,N_8789);
and U8807 (N_8807,N_8687,N_8633);
nor U8808 (N_8808,N_8678,N_8606);
or U8809 (N_8809,N_8757,N_8664);
or U8810 (N_8810,N_8748,N_8753);
and U8811 (N_8811,N_8710,N_8622);
and U8812 (N_8812,N_8761,N_8695);
or U8813 (N_8813,N_8679,N_8641);
xnor U8814 (N_8814,N_8698,N_8772);
nor U8815 (N_8815,N_8740,N_8600);
or U8816 (N_8816,N_8603,N_8661);
nand U8817 (N_8817,N_8666,N_8645);
and U8818 (N_8818,N_8605,N_8670);
or U8819 (N_8819,N_8604,N_8732);
and U8820 (N_8820,N_8702,N_8655);
nor U8821 (N_8821,N_8712,N_8683);
and U8822 (N_8822,N_8762,N_8721);
or U8823 (N_8823,N_8718,N_8682);
or U8824 (N_8824,N_8684,N_8730);
and U8825 (N_8825,N_8787,N_8743);
or U8826 (N_8826,N_8639,N_8771);
xnor U8827 (N_8827,N_8715,N_8674);
nor U8828 (N_8828,N_8671,N_8775);
nor U8829 (N_8829,N_8711,N_8745);
xnor U8830 (N_8830,N_8708,N_8630);
nor U8831 (N_8831,N_8786,N_8613);
nor U8832 (N_8832,N_8681,N_8785);
or U8833 (N_8833,N_8617,N_8676);
xnor U8834 (N_8834,N_8643,N_8662);
or U8835 (N_8835,N_8781,N_8727);
or U8836 (N_8836,N_8640,N_8624);
and U8837 (N_8837,N_8729,N_8707);
xnor U8838 (N_8838,N_8642,N_8657);
nand U8839 (N_8839,N_8653,N_8742);
nand U8840 (N_8840,N_8788,N_8767);
or U8841 (N_8841,N_8689,N_8615);
nand U8842 (N_8842,N_8709,N_8669);
xnor U8843 (N_8843,N_8714,N_8675);
and U8844 (N_8844,N_8607,N_8609);
and U8845 (N_8845,N_8716,N_8618);
or U8846 (N_8846,N_8765,N_8783);
nor U8847 (N_8847,N_8779,N_8636);
or U8848 (N_8848,N_8752,N_8638);
and U8849 (N_8849,N_8737,N_8621);
xnor U8850 (N_8850,N_8686,N_8747);
and U8851 (N_8851,N_8749,N_8790);
or U8852 (N_8852,N_8733,N_8672);
nor U8853 (N_8853,N_8667,N_8608);
or U8854 (N_8854,N_8736,N_8625);
nand U8855 (N_8855,N_8764,N_8652);
nand U8856 (N_8856,N_8632,N_8628);
and U8857 (N_8857,N_8739,N_8784);
nor U8858 (N_8858,N_8646,N_8797);
nor U8859 (N_8859,N_8717,N_8650);
nand U8860 (N_8860,N_8692,N_8769);
or U8861 (N_8861,N_8726,N_8658);
nand U8862 (N_8862,N_8760,N_8616);
nand U8863 (N_8863,N_8756,N_8777);
or U8864 (N_8864,N_8697,N_8701);
nor U8865 (N_8865,N_8629,N_8793);
nor U8866 (N_8866,N_8623,N_8734);
and U8867 (N_8867,N_8759,N_8723);
nor U8868 (N_8868,N_8651,N_8795);
or U8869 (N_8869,N_8656,N_8706);
nor U8870 (N_8870,N_8626,N_8610);
xor U8871 (N_8871,N_8799,N_8794);
and U8872 (N_8872,N_8768,N_8738);
nand U8873 (N_8873,N_8798,N_8735);
nor U8874 (N_8874,N_8755,N_8668);
nor U8875 (N_8875,N_8685,N_8700);
and U8876 (N_8876,N_8719,N_8637);
nor U8877 (N_8877,N_8688,N_8654);
or U8878 (N_8878,N_8694,N_8770);
nor U8879 (N_8879,N_8792,N_8634);
nor U8880 (N_8880,N_8780,N_8703);
and U8881 (N_8881,N_8631,N_8649);
or U8882 (N_8882,N_8763,N_8782);
or U8883 (N_8883,N_8680,N_8647);
nand U8884 (N_8884,N_8705,N_8746);
or U8885 (N_8885,N_8620,N_8673);
or U8886 (N_8886,N_8728,N_8731);
xnor U8887 (N_8887,N_8766,N_8612);
nand U8888 (N_8888,N_8758,N_8635);
and U8889 (N_8889,N_8648,N_8776);
and U8890 (N_8890,N_8725,N_8720);
nand U8891 (N_8891,N_8691,N_8774);
xnor U8892 (N_8892,N_8611,N_8665);
nor U8893 (N_8893,N_8627,N_8696);
or U8894 (N_8894,N_8602,N_8677);
nor U8895 (N_8895,N_8704,N_8644);
nor U8896 (N_8896,N_8614,N_8601);
or U8897 (N_8897,N_8751,N_8724);
xor U8898 (N_8898,N_8699,N_8778);
or U8899 (N_8899,N_8693,N_8690);
nand U8900 (N_8900,N_8705,N_8656);
or U8901 (N_8901,N_8772,N_8789);
and U8902 (N_8902,N_8679,N_8710);
and U8903 (N_8903,N_8735,N_8703);
xnor U8904 (N_8904,N_8675,N_8643);
or U8905 (N_8905,N_8778,N_8681);
and U8906 (N_8906,N_8771,N_8736);
or U8907 (N_8907,N_8700,N_8659);
and U8908 (N_8908,N_8686,N_8623);
nor U8909 (N_8909,N_8645,N_8784);
nand U8910 (N_8910,N_8767,N_8684);
nor U8911 (N_8911,N_8684,N_8631);
nand U8912 (N_8912,N_8707,N_8640);
or U8913 (N_8913,N_8719,N_8704);
and U8914 (N_8914,N_8748,N_8764);
xnor U8915 (N_8915,N_8642,N_8765);
nor U8916 (N_8916,N_8679,N_8621);
nand U8917 (N_8917,N_8629,N_8686);
or U8918 (N_8918,N_8635,N_8735);
and U8919 (N_8919,N_8720,N_8705);
or U8920 (N_8920,N_8637,N_8609);
nand U8921 (N_8921,N_8727,N_8780);
nand U8922 (N_8922,N_8699,N_8640);
and U8923 (N_8923,N_8644,N_8695);
and U8924 (N_8924,N_8673,N_8744);
and U8925 (N_8925,N_8647,N_8630);
nor U8926 (N_8926,N_8616,N_8729);
nor U8927 (N_8927,N_8780,N_8711);
nor U8928 (N_8928,N_8611,N_8720);
and U8929 (N_8929,N_8705,N_8671);
nor U8930 (N_8930,N_8681,N_8783);
or U8931 (N_8931,N_8783,N_8671);
nor U8932 (N_8932,N_8763,N_8613);
xor U8933 (N_8933,N_8704,N_8757);
nor U8934 (N_8934,N_8794,N_8728);
xnor U8935 (N_8935,N_8676,N_8658);
nor U8936 (N_8936,N_8740,N_8643);
nor U8937 (N_8937,N_8761,N_8628);
and U8938 (N_8938,N_8614,N_8687);
nor U8939 (N_8939,N_8648,N_8643);
xor U8940 (N_8940,N_8600,N_8724);
or U8941 (N_8941,N_8689,N_8700);
nor U8942 (N_8942,N_8631,N_8738);
and U8943 (N_8943,N_8655,N_8740);
or U8944 (N_8944,N_8750,N_8730);
nor U8945 (N_8945,N_8665,N_8692);
and U8946 (N_8946,N_8620,N_8765);
or U8947 (N_8947,N_8736,N_8660);
xnor U8948 (N_8948,N_8742,N_8674);
and U8949 (N_8949,N_8789,N_8661);
nand U8950 (N_8950,N_8741,N_8710);
nor U8951 (N_8951,N_8737,N_8670);
xnor U8952 (N_8952,N_8674,N_8795);
or U8953 (N_8953,N_8774,N_8769);
and U8954 (N_8954,N_8732,N_8631);
nand U8955 (N_8955,N_8643,N_8697);
nor U8956 (N_8956,N_8667,N_8751);
and U8957 (N_8957,N_8754,N_8625);
nor U8958 (N_8958,N_8771,N_8756);
nand U8959 (N_8959,N_8737,N_8606);
xor U8960 (N_8960,N_8754,N_8776);
nand U8961 (N_8961,N_8665,N_8733);
nand U8962 (N_8962,N_8711,N_8795);
and U8963 (N_8963,N_8736,N_8694);
nand U8964 (N_8964,N_8646,N_8661);
or U8965 (N_8965,N_8705,N_8719);
nor U8966 (N_8966,N_8635,N_8600);
nor U8967 (N_8967,N_8631,N_8644);
or U8968 (N_8968,N_8625,N_8722);
or U8969 (N_8969,N_8683,N_8797);
nand U8970 (N_8970,N_8775,N_8660);
and U8971 (N_8971,N_8645,N_8610);
or U8972 (N_8972,N_8608,N_8619);
or U8973 (N_8973,N_8651,N_8670);
and U8974 (N_8974,N_8784,N_8756);
or U8975 (N_8975,N_8677,N_8625);
and U8976 (N_8976,N_8720,N_8686);
xnor U8977 (N_8977,N_8622,N_8731);
nor U8978 (N_8978,N_8623,N_8799);
or U8979 (N_8979,N_8645,N_8786);
nand U8980 (N_8980,N_8780,N_8647);
or U8981 (N_8981,N_8653,N_8791);
and U8982 (N_8982,N_8737,N_8658);
nand U8983 (N_8983,N_8758,N_8677);
xor U8984 (N_8984,N_8793,N_8691);
nand U8985 (N_8985,N_8706,N_8643);
nor U8986 (N_8986,N_8748,N_8660);
nor U8987 (N_8987,N_8734,N_8606);
nand U8988 (N_8988,N_8694,N_8713);
nand U8989 (N_8989,N_8756,N_8626);
nand U8990 (N_8990,N_8766,N_8757);
nand U8991 (N_8991,N_8668,N_8724);
or U8992 (N_8992,N_8611,N_8612);
or U8993 (N_8993,N_8783,N_8609);
nand U8994 (N_8994,N_8751,N_8712);
nor U8995 (N_8995,N_8691,N_8663);
nor U8996 (N_8996,N_8741,N_8607);
or U8997 (N_8997,N_8715,N_8600);
and U8998 (N_8998,N_8600,N_8752);
nor U8999 (N_8999,N_8610,N_8685);
or U9000 (N_9000,N_8984,N_8833);
or U9001 (N_9001,N_8853,N_8926);
nor U9002 (N_9002,N_8965,N_8937);
nand U9003 (N_9003,N_8959,N_8826);
or U9004 (N_9004,N_8838,N_8943);
and U9005 (N_9005,N_8946,N_8989);
nor U9006 (N_9006,N_8875,N_8818);
nor U9007 (N_9007,N_8848,N_8842);
or U9008 (N_9008,N_8877,N_8806);
nor U9009 (N_9009,N_8867,N_8814);
nand U9010 (N_9010,N_8961,N_8908);
xor U9011 (N_9011,N_8973,N_8841);
and U9012 (N_9012,N_8930,N_8804);
and U9013 (N_9013,N_8944,N_8888);
or U9014 (N_9014,N_8822,N_8932);
nor U9015 (N_9015,N_8820,N_8846);
nor U9016 (N_9016,N_8917,N_8947);
nor U9017 (N_9017,N_8900,N_8898);
nor U9018 (N_9018,N_8985,N_8992);
nor U9019 (N_9019,N_8987,N_8873);
nor U9020 (N_9020,N_8843,N_8956);
nor U9021 (N_9021,N_8828,N_8864);
nor U9022 (N_9022,N_8810,N_8816);
nand U9023 (N_9023,N_8954,N_8881);
xnor U9024 (N_9024,N_8983,N_8845);
and U9025 (N_9025,N_8868,N_8981);
and U9026 (N_9026,N_8861,N_8976);
or U9027 (N_9027,N_8974,N_8837);
nor U9028 (N_9028,N_8817,N_8883);
or U9029 (N_9029,N_8966,N_8830);
nand U9030 (N_9030,N_8894,N_8948);
or U9031 (N_9031,N_8825,N_8986);
and U9032 (N_9032,N_8933,N_8805);
nor U9033 (N_9033,N_8887,N_8803);
nand U9034 (N_9034,N_8823,N_8870);
nand U9035 (N_9035,N_8844,N_8935);
or U9036 (N_9036,N_8949,N_8879);
xor U9037 (N_9037,N_8978,N_8811);
nand U9038 (N_9038,N_8960,N_8902);
nor U9039 (N_9039,N_8847,N_8945);
or U9040 (N_9040,N_8899,N_8855);
and U9041 (N_9041,N_8871,N_8852);
nand U9042 (N_9042,N_8982,N_8851);
nand U9043 (N_9043,N_8931,N_8800);
and U9044 (N_9044,N_8904,N_8880);
nand U9045 (N_9045,N_8807,N_8963);
nand U9046 (N_9046,N_8969,N_8874);
nand U9047 (N_9047,N_8957,N_8882);
nand U9048 (N_9048,N_8849,N_8907);
xnor U9049 (N_9049,N_8928,N_8850);
and U9050 (N_9050,N_8919,N_8953);
nor U9051 (N_9051,N_8920,N_8921);
nor U9052 (N_9052,N_8934,N_8952);
xor U9053 (N_9053,N_8942,N_8940);
or U9054 (N_9054,N_8834,N_8922);
and U9055 (N_9055,N_8859,N_8962);
or U9056 (N_9056,N_8821,N_8909);
nor U9057 (N_9057,N_8812,N_8975);
xnor U9058 (N_9058,N_8980,N_8813);
or U9059 (N_9059,N_8801,N_8808);
and U9060 (N_9060,N_8964,N_8896);
nor U9061 (N_9061,N_8872,N_8906);
nor U9062 (N_9062,N_8839,N_8835);
nor U9063 (N_9063,N_8829,N_8912);
or U9064 (N_9064,N_8990,N_8876);
xnor U9065 (N_9065,N_8911,N_8967);
or U9066 (N_9066,N_8941,N_8938);
nand U9067 (N_9067,N_8998,N_8955);
nor U9068 (N_9068,N_8802,N_8939);
nand U9069 (N_9069,N_8892,N_8815);
or U9070 (N_9070,N_8903,N_8905);
nand U9071 (N_9071,N_8856,N_8809);
xnor U9072 (N_9072,N_8950,N_8854);
or U9073 (N_9073,N_8878,N_8893);
nand U9074 (N_9074,N_8866,N_8977);
nor U9075 (N_9075,N_8840,N_8889);
and U9076 (N_9076,N_8913,N_8890);
nand U9077 (N_9077,N_8991,N_8885);
nor U9078 (N_9078,N_8999,N_8824);
and U9079 (N_9079,N_8884,N_8897);
and U9080 (N_9080,N_8972,N_8971);
and U9081 (N_9081,N_8958,N_8869);
nand U9082 (N_9082,N_8979,N_8832);
xnor U9083 (N_9083,N_8988,N_8923);
nor U9084 (N_9084,N_8994,N_8927);
nor U9085 (N_9085,N_8970,N_8997);
nand U9086 (N_9086,N_8993,N_8916);
nand U9087 (N_9087,N_8929,N_8901);
nor U9088 (N_9088,N_8936,N_8910);
nand U9089 (N_9089,N_8995,N_8925);
and U9090 (N_9090,N_8915,N_8860);
and U9091 (N_9091,N_8858,N_8996);
nand U9092 (N_9092,N_8863,N_8831);
nor U9093 (N_9093,N_8865,N_8914);
nor U9094 (N_9094,N_8836,N_8827);
xnor U9095 (N_9095,N_8968,N_8951);
nand U9096 (N_9096,N_8862,N_8918);
or U9097 (N_9097,N_8891,N_8857);
nand U9098 (N_9098,N_8895,N_8924);
and U9099 (N_9099,N_8819,N_8886);
nor U9100 (N_9100,N_8837,N_8828);
or U9101 (N_9101,N_8865,N_8839);
xor U9102 (N_9102,N_8854,N_8869);
xnor U9103 (N_9103,N_8814,N_8998);
or U9104 (N_9104,N_8992,N_8990);
and U9105 (N_9105,N_8914,N_8896);
and U9106 (N_9106,N_8912,N_8874);
or U9107 (N_9107,N_8993,N_8955);
nor U9108 (N_9108,N_8951,N_8894);
nor U9109 (N_9109,N_8924,N_8893);
xor U9110 (N_9110,N_8957,N_8997);
nor U9111 (N_9111,N_8809,N_8992);
or U9112 (N_9112,N_8978,N_8873);
and U9113 (N_9113,N_8931,N_8882);
and U9114 (N_9114,N_8845,N_8895);
and U9115 (N_9115,N_8826,N_8883);
or U9116 (N_9116,N_8941,N_8911);
or U9117 (N_9117,N_8943,N_8898);
and U9118 (N_9118,N_8824,N_8811);
and U9119 (N_9119,N_8845,N_8847);
or U9120 (N_9120,N_8895,N_8888);
xor U9121 (N_9121,N_8920,N_8891);
nand U9122 (N_9122,N_8827,N_8898);
xor U9123 (N_9123,N_8907,N_8864);
or U9124 (N_9124,N_8941,N_8983);
nor U9125 (N_9125,N_8932,N_8859);
nor U9126 (N_9126,N_8879,N_8980);
or U9127 (N_9127,N_8911,N_8814);
nor U9128 (N_9128,N_8991,N_8926);
nand U9129 (N_9129,N_8982,N_8899);
and U9130 (N_9130,N_8919,N_8940);
xnor U9131 (N_9131,N_8889,N_8991);
and U9132 (N_9132,N_8870,N_8827);
nand U9133 (N_9133,N_8958,N_8984);
or U9134 (N_9134,N_8976,N_8855);
nor U9135 (N_9135,N_8817,N_8995);
nor U9136 (N_9136,N_8894,N_8879);
nand U9137 (N_9137,N_8812,N_8919);
nor U9138 (N_9138,N_8901,N_8969);
nand U9139 (N_9139,N_8823,N_8990);
xnor U9140 (N_9140,N_8974,N_8911);
and U9141 (N_9141,N_8911,N_8896);
and U9142 (N_9142,N_8977,N_8999);
or U9143 (N_9143,N_8873,N_8953);
and U9144 (N_9144,N_8972,N_8970);
and U9145 (N_9145,N_8949,N_8876);
and U9146 (N_9146,N_8939,N_8910);
nor U9147 (N_9147,N_8850,N_8836);
and U9148 (N_9148,N_8984,N_8955);
nor U9149 (N_9149,N_8994,N_8905);
nor U9150 (N_9150,N_8991,N_8951);
nand U9151 (N_9151,N_8978,N_8960);
nand U9152 (N_9152,N_8998,N_8951);
and U9153 (N_9153,N_8958,N_8886);
and U9154 (N_9154,N_8953,N_8858);
and U9155 (N_9155,N_8848,N_8975);
and U9156 (N_9156,N_8832,N_8905);
nand U9157 (N_9157,N_8950,N_8866);
nand U9158 (N_9158,N_8904,N_8997);
and U9159 (N_9159,N_8953,N_8962);
and U9160 (N_9160,N_8949,N_8859);
or U9161 (N_9161,N_8855,N_8809);
and U9162 (N_9162,N_8993,N_8961);
nor U9163 (N_9163,N_8935,N_8883);
and U9164 (N_9164,N_8906,N_8905);
nor U9165 (N_9165,N_8979,N_8969);
nor U9166 (N_9166,N_8845,N_8987);
or U9167 (N_9167,N_8881,N_8862);
nor U9168 (N_9168,N_8942,N_8907);
or U9169 (N_9169,N_8975,N_8911);
and U9170 (N_9170,N_8862,N_8831);
and U9171 (N_9171,N_8882,N_8951);
nand U9172 (N_9172,N_8813,N_8811);
and U9173 (N_9173,N_8867,N_8853);
and U9174 (N_9174,N_8925,N_8994);
nor U9175 (N_9175,N_8939,N_8800);
or U9176 (N_9176,N_8852,N_8861);
xnor U9177 (N_9177,N_8834,N_8831);
nand U9178 (N_9178,N_8801,N_8928);
and U9179 (N_9179,N_8967,N_8943);
and U9180 (N_9180,N_8876,N_8852);
and U9181 (N_9181,N_8891,N_8801);
nor U9182 (N_9182,N_8874,N_8980);
nor U9183 (N_9183,N_8866,N_8914);
and U9184 (N_9184,N_8873,N_8989);
and U9185 (N_9185,N_8870,N_8808);
or U9186 (N_9186,N_8896,N_8856);
nor U9187 (N_9187,N_8860,N_8938);
nor U9188 (N_9188,N_8960,N_8923);
or U9189 (N_9189,N_8949,N_8816);
xnor U9190 (N_9190,N_8829,N_8889);
or U9191 (N_9191,N_8879,N_8830);
or U9192 (N_9192,N_8956,N_8891);
and U9193 (N_9193,N_8845,N_8804);
nor U9194 (N_9194,N_8924,N_8813);
and U9195 (N_9195,N_8989,N_8841);
and U9196 (N_9196,N_8813,N_8905);
nor U9197 (N_9197,N_8960,N_8979);
nand U9198 (N_9198,N_8883,N_8981);
xnor U9199 (N_9199,N_8987,N_8911);
nor U9200 (N_9200,N_9087,N_9167);
nand U9201 (N_9201,N_9063,N_9059);
xnor U9202 (N_9202,N_9173,N_9036);
or U9203 (N_9203,N_9004,N_9190);
or U9204 (N_9204,N_9155,N_9006);
and U9205 (N_9205,N_9189,N_9079);
nand U9206 (N_9206,N_9081,N_9102);
or U9207 (N_9207,N_9181,N_9027);
nor U9208 (N_9208,N_9135,N_9095);
nor U9209 (N_9209,N_9172,N_9051);
or U9210 (N_9210,N_9157,N_9021);
nor U9211 (N_9211,N_9066,N_9024);
nand U9212 (N_9212,N_9074,N_9048);
nor U9213 (N_9213,N_9179,N_9086);
xnor U9214 (N_9214,N_9065,N_9057);
or U9215 (N_9215,N_9075,N_9182);
nor U9216 (N_9216,N_9114,N_9023);
nand U9217 (N_9217,N_9145,N_9105);
or U9218 (N_9218,N_9144,N_9185);
or U9219 (N_9219,N_9191,N_9045);
or U9220 (N_9220,N_9106,N_9003);
nand U9221 (N_9221,N_9025,N_9168);
or U9222 (N_9222,N_9198,N_9110);
nand U9223 (N_9223,N_9089,N_9118);
nand U9224 (N_9224,N_9115,N_9124);
xnor U9225 (N_9225,N_9097,N_9064);
nor U9226 (N_9226,N_9177,N_9180);
nand U9227 (N_9227,N_9176,N_9119);
xor U9228 (N_9228,N_9037,N_9033);
and U9229 (N_9229,N_9088,N_9002);
nor U9230 (N_9230,N_9160,N_9090);
nand U9231 (N_9231,N_9158,N_9055);
nor U9232 (N_9232,N_9132,N_9111);
nor U9233 (N_9233,N_9101,N_9053);
and U9234 (N_9234,N_9136,N_9121);
xor U9235 (N_9235,N_9142,N_9193);
nand U9236 (N_9236,N_9017,N_9125);
nand U9237 (N_9237,N_9060,N_9197);
nand U9238 (N_9238,N_9152,N_9164);
and U9239 (N_9239,N_9034,N_9195);
xnor U9240 (N_9240,N_9031,N_9032);
nand U9241 (N_9241,N_9013,N_9153);
nand U9242 (N_9242,N_9183,N_9016);
and U9243 (N_9243,N_9163,N_9073);
nand U9244 (N_9244,N_9096,N_9161);
xnor U9245 (N_9245,N_9169,N_9188);
nand U9246 (N_9246,N_9151,N_9147);
nand U9247 (N_9247,N_9078,N_9137);
nand U9248 (N_9248,N_9149,N_9071);
nor U9249 (N_9249,N_9170,N_9103);
xnor U9250 (N_9250,N_9082,N_9046);
and U9251 (N_9251,N_9120,N_9056);
and U9252 (N_9252,N_9099,N_9122);
and U9253 (N_9253,N_9113,N_9070);
and U9254 (N_9254,N_9194,N_9139);
and U9255 (N_9255,N_9062,N_9148);
nor U9256 (N_9256,N_9008,N_9196);
nand U9257 (N_9257,N_9159,N_9133);
or U9258 (N_9258,N_9035,N_9117);
and U9259 (N_9259,N_9038,N_9007);
or U9260 (N_9260,N_9192,N_9041);
nand U9261 (N_9261,N_9058,N_9043);
nor U9262 (N_9262,N_9026,N_9108);
nor U9263 (N_9263,N_9014,N_9022);
or U9264 (N_9264,N_9029,N_9116);
or U9265 (N_9265,N_9085,N_9175);
nand U9266 (N_9266,N_9165,N_9112);
nand U9267 (N_9267,N_9156,N_9083);
xnor U9268 (N_9268,N_9011,N_9130);
and U9269 (N_9269,N_9077,N_9084);
nand U9270 (N_9270,N_9104,N_9109);
xnor U9271 (N_9271,N_9049,N_9123);
nand U9272 (N_9272,N_9098,N_9171);
or U9273 (N_9273,N_9072,N_9001);
nand U9274 (N_9274,N_9092,N_9107);
nand U9275 (N_9275,N_9000,N_9044);
or U9276 (N_9276,N_9174,N_9186);
nand U9277 (N_9277,N_9067,N_9146);
or U9278 (N_9278,N_9020,N_9100);
nor U9279 (N_9279,N_9128,N_9050);
or U9280 (N_9280,N_9134,N_9140);
nor U9281 (N_9281,N_9030,N_9080);
or U9282 (N_9282,N_9061,N_9131);
nand U9283 (N_9283,N_9047,N_9039);
and U9284 (N_9284,N_9094,N_9005);
nand U9285 (N_9285,N_9091,N_9150);
nand U9286 (N_9286,N_9138,N_9199);
or U9287 (N_9287,N_9069,N_9178);
xnor U9288 (N_9288,N_9154,N_9010);
and U9289 (N_9289,N_9052,N_9068);
nand U9290 (N_9290,N_9019,N_9042);
nand U9291 (N_9291,N_9184,N_9166);
nand U9292 (N_9292,N_9012,N_9076);
or U9293 (N_9293,N_9015,N_9028);
nand U9294 (N_9294,N_9018,N_9040);
nor U9295 (N_9295,N_9162,N_9187);
xnor U9296 (N_9296,N_9143,N_9009);
or U9297 (N_9297,N_9093,N_9141);
xor U9298 (N_9298,N_9127,N_9126);
nand U9299 (N_9299,N_9129,N_9054);
or U9300 (N_9300,N_9169,N_9084);
nor U9301 (N_9301,N_9191,N_9027);
nand U9302 (N_9302,N_9034,N_9166);
nand U9303 (N_9303,N_9099,N_9027);
nor U9304 (N_9304,N_9074,N_9092);
and U9305 (N_9305,N_9063,N_9175);
or U9306 (N_9306,N_9175,N_9144);
nand U9307 (N_9307,N_9040,N_9073);
or U9308 (N_9308,N_9019,N_9016);
nand U9309 (N_9309,N_9045,N_9048);
or U9310 (N_9310,N_9120,N_9021);
nor U9311 (N_9311,N_9173,N_9155);
xnor U9312 (N_9312,N_9049,N_9009);
and U9313 (N_9313,N_9142,N_9035);
and U9314 (N_9314,N_9031,N_9009);
or U9315 (N_9315,N_9010,N_9067);
nand U9316 (N_9316,N_9128,N_9015);
and U9317 (N_9317,N_9117,N_9154);
xnor U9318 (N_9318,N_9081,N_9073);
and U9319 (N_9319,N_9068,N_9099);
and U9320 (N_9320,N_9131,N_9102);
nand U9321 (N_9321,N_9038,N_9009);
xor U9322 (N_9322,N_9103,N_9130);
and U9323 (N_9323,N_9134,N_9120);
and U9324 (N_9324,N_9079,N_9159);
and U9325 (N_9325,N_9150,N_9083);
and U9326 (N_9326,N_9072,N_9192);
or U9327 (N_9327,N_9151,N_9177);
or U9328 (N_9328,N_9192,N_9163);
nand U9329 (N_9329,N_9016,N_9077);
or U9330 (N_9330,N_9061,N_9115);
nor U9331 (N_9331,N_9060,N_9028);
nand U9332 (N_9332,N_9066,N_9145);
nor U9333 (N_9333,N_9050,N_9148);
and U9334 (N_9334,N_9041,N_9154);
nor U9335 (N_9335,N_9095,N_9077);
or U9336 (N_9336,N_9169,N_9026);
nand U9337 (N_9337,N_9082,N_9149);
nand U9338 (N_9338,N_9048,N_9193);
and U9339 (N_9339,N_9088,N_9114);
and U9340 (N_9340,N_9089,N_9122);
nor U9341 (N_9341,N_9055,N_9000);
and U9342 (N_9342,N_9177,N_9083);
nand U9343 (N_9343,N_9155,N_9109);
nand U9344 (N_9344,N_9021,N_9108);
xor U9345 (N_9345,N_9032,N_9132);
nand U9346 (N_9346,N_9053,N_9183);
nor U9347 (N_9347,N_9148,N_9198);
nand U9348 (N_9348,N_9000,N_9164);
xnor U9349 (N_9349,N_9113,N_9066);
and U9350 (N_9350,N_9131,N_9029);
or U9351 (N_9351,N_9047,N_9023);
nand U9352 (N_9352,N_9111,N_9043);
nand U9353 (N_9353,N_9089,N_9019);
nor U9354 (N_9354,N_9031,N_9125);
nor U9355 (N_9355,N_9077,N_9151);
nand U9356 (N_9356,N_9085,N_9118);
and U9357 (N_9357,N_9131,N_9088);
and U9358 (N_9358,N_9114,N_9150);
nor U9359 (N_9359,N_9018,N_9082);
nand U9360 (N_9360,N_9187,N_9025);
or U9361 (N_9361,N_9117,N_9181);
xor U9362 (N_9362,N_9197,N_9187);
and U9363 (N_9363,N_9178,N_9131);
and U9364 (N_9364,N_9157,N_9184);
nand U9365 (N_9365,N_9073,N_9052);
or U9366 (N_9366,N_9081,N_9046);
nor U9367 (N_9367,N_9036,N_9199);
xor U9368 (N_9368,N_9181,N_9047);
nor U9369 (N_9369,N_9015,N_9036);
xnor U9370 (N_9370,N_9008,N_9168);
and U9371 (N_9371,N_9113,N_9182);
or U9372 (N_9372,N_9139,N_9009);
nand U9373 (N_9373,N_9181,N_9053);
nor U9374 (N_9374,N_9049,N_9164);
nand U9375 (N_9375,N_9027,N_9124);
and U9376 (N_9376,N_9052,N_9140);
and U9377 (N_9377,N_9096,N_9076);
or U9378 (N_9378,N_9034,N_9040);
or U9379 (N_9379,N_9112,N_9000);
nand U9380 (N_9380,N_9088,N_9124);
nand U9381 (N_9381,N_9059,N_9147);
nor U9382 (N_9382,N_9163,N_9058);
and U9383 (N_9383,N_9122,N_9108);
nor U9384 (N_9384,N_9078,N_9047);
and U9385 (N_9385,N_9172,N_9043);
nor U9386 (N_9386,N_9005,N_9105);
nor U9387 (N_9387,N_9191,N_9183);
and U9388 (N_9388,N_9047,N_9028);
nor U9389 (N_9389,N_9008,N_9050);
or U9390 (N_9390,N_9049,N_9158);
xnor U9391 (N_9391,N_9175,N_9139);
xnor U9392 (N_9392,N_9094,N_9191);
or U9393 (N_9393,N_9082,N_9052);
or U9394 (N_9394,N_9144,N_9081);
or U9395 (N_9395,N_9084,N_9008);
and U9396 (N_9396,N_9070,N_9087);
nand U9397 (N_9397,N_9049,N_9139);
nor U9398 (N_9398,N_9012,N_9087);
nor U9399 (N_9399,N_9047,N_9184);
nand U9400 (N_9400,N_9213,N_9387);
nand U9401 (N_9401,N_9251,N_9377);
xor U9402 (N_9402,N_9384,N_9262);
xor U9403 (N_9403,N_9295,N_9289);
and U9404 (N_9404,N_9224,N_9381);
nor U9405 (N_9405,N_9243,N_9278);
and U9406 (N_9406,N_9332,N_9327);
nor U9407 (N_9407,N_9385,N_9312);
nand U9408 (N_9408,N_9306,N_9275);
or U9409 (N_9409,N_9282,N_9394);
nor U9410 (N_9410,N_9247,N_9216);
or U9411 (N_9411,N_9211,N_9283);
or U9412 (N_9412,N_9374,N_9218);
nor U9413 (N_9413,N_9348,N_9212);
and U9414 (N_9414,N_9205,N_9279);
nor U9415 (N_9415,N_9305,N_9241);
nor U9416 (N_9416,N_9227,N_9366);
nand U9417 (N_9417,N_9353,N_9274);
and U9418 (N_9418,N_9233,N_9370);
nand U9419 (N_9419,N_9378,N_9259);
nand U9420 (N_9420,N_9389,N_9393);
nor U9421 (N_9421,N_9362,N_9313);
and U9422 (N_9422,N_9386,N_9284);
xor U9423 (N_9423,N_9256,N_9300);
nor U9424 (N_9424,N_9225,N_9215);
nor U9425 (N_9425,N_9323,N_9331);
nand U9426 (N_9426,N_9214,N_9268);
or U9427 (N_9427,N_9201,N_9238);
nand U9428 (N_9428,N_9302,N_9292);
or U9429 (N_9429,N_9263,N_9254);
nand U9430 (N_9430,N_9342,N_9363);
or U9431 (N_9431,N_9367,N_9203);
or U9432 (N_9432,N_9288,N_9336);
and U9433 (N_9433,N_9217,N_9337);
nand U9434 (N_9434,N_9317,N_9258);
nor U9435 (N_9435,N_9286,N_9221);
nor U9436 (N_9436,N_9349,N_9294);
or U9437 (N_9437,N_9299,N_9209);
nor U9438 (N_9438,N_9310,N_9273);
nand U9439 (N_9439,N_9388,N_9356);
and U9440 (N_9440,N_9340,N_9333);
nor U9441 (N_9441,N_9298,N_9272);
nand U9442 (N_9442,N_9246,N_9372);
and U9443 (N_9443,N_9260,N_9228);
nand U9444 (N_9444,N_9344,N_9307);
nor U9445 (N_9445,N_9244,N_9252);
or U9446 (N_9446,N_9220,N_9219);
nor U9447 (N_9447,N_9208,N_9230);
nand U9448 (N_9448,N_9301,N_9304);
or U9449 (N_9449,N_9204,N_9264);
nand U9450 (N_9450,N_9207,N_9343);
or U9451 (N_9451,N_9399,N_9235);
xnor U9452 (N_9452,N_9239,N_9280);
nor U9453 (N_9453,N_9261,N_9202);
nor U9454 (N_9454,N_9266,N_9345);
and U9455 (N_9455,N_9321,N_9267);
or U9456 (N_9456,N_9376,N_9350);
and U9457 (N_9457,N_9365,N_9293);
and U9458 (N_9458,N_9245,N_9250);
and U9459 (N_9459,N_9368,N_9358);
and U9460 (N_9460,N_9346,N_9277);
nand U9461 (N_9461,N_9319,N_9395);
or U9462 (N_9462,N_9396,N_9271);
and U9463 (N_9463,N_9322,N_9291);
xnor U9464 (N_9464,N_9276,N_9287);
or U9465 (N_9465,N_9265,N_9237);
and U9466 (N_9466,N_9354,N_9379);
nor U9467 (N_9467,N_9242,N_9231);
and U9468 (N_9468,N_9296,N_9316);
xnor U9469 (N_9469,N_9281,N_9341);
nand U9470 (N_9470,N_9240,N_9355);
and U9471 (N_9471,N_9318,N_9369);
xnor U9472 (N_9472,N_9236,N_9390);
nor U9473 (N_9473,N_9325,N_9361);
and U9474 (N_9474,N_9206,N_9398);
and U9475 (N_9475,N_9222,N_9373);
nand U9476 (N_9476,N_9339,N_9270);
or U9477 (N_9477,N_9364,N_9255);
nor U9478 (N_9478,N_9248,N_9352);
or U9479 (N_9479,N_9303,N_9285);
nand U9480 (N_9480,N_9382,N_9253);
nand U9481 (N_9481,N_9397,N_9234);
and U9482 (N_9482,N_9326,N_9383);
xor U9483 (N_9483,N_9375,N_9328);
xnor U9484 (N_9484,N_9347,N_9309);
and U9485 (N_9485,N_9229,N_9226);
or U9486 (N_9486,N_9257,N_9359);
nor U9487 (N_9487,N_9334,N_9269);
nor U9488 (N_9488,N_9290,N_9210);
and U9489 (N_9489,N_9311,N_9335);
nor U9490 (N_9490,N_9360,N_9391);
xnor U9491 (N_9491,N_9380,N_9223);
nand U9492 (N_9492,N_9330,N_9357);
or U9493 (N_9493,N_9324,N_9249);
nand U9494 (N_9494,N_9392,N_9329);
or U9495 (N_9495,N_9232,N_9371);
and U9496 (N_9496,N_9200,N_9351);
nor U9497 (N_9497,N_9308,N_9297);
xnor U9498 (N_9498,N_9338,N_9320);
and U9499 (N_9499,N_9315,N_9314);
or U9500 (N_9500,N_9256,N_9281);
nor U9501 (N_9501,N_9320,N_9286);
nand U9502 (N_9502,N_9336,N_9237);
nor U9503 (N_9503,N_9358,N_9232);
or U9504 (N_9504,N_9256,N_9348);
nand U9505 (N_9505,N_9309,N_9325);
and U9506 (N_9506,N_9301,N_9387);
nand U9507 (N_9507,N_9350,N_9394);
or U9508 (N_9508,N_9292,N_9288);
nor U9509 (N_9509,N_9360,N_9273);
and U9510 (N_9510,N_9207,N_9200);
or U9511 (N_9511,N_9224,N_9228);
and U9512 (N_9512,N_9257,N_9237);
and U9513 (N_9513,N_9230,N_9264);
or U9514 (N_9514,N_9353,N_9228);
and U9515 (N_9515,N_9222,N_9340);
nand U9516 (N_9516,N_9245,N_9216);
and U9517 (N_9517,N_9217,N_9395);
nand U9518 (N_9518,N_9319,N_9254);
or U9519 (N_9519,N_9203,N_9287);
nor U9520 (N_9520,N_9398,N_9314);
nand U9521 (N_9521,N_9390,N_9284);
nor U9522 (N_9522,N_9236,N_9318);
xor U9523 (N_9523,N_9282,N_9369);
and U9524 (N_9524,N_9217,N_9214);
nand U9525 (N_9525,N_9239,N_9240);
nor U9526 (N_9526,N_9330,N_9230);
and U9527 (N_9527,N_9248,N_9313);
nand U9528 (N_9528,N_9315,N_9355);
or U9529 (N_9529,N_9294,N_9301);
nor U9530 (N_9530,N_9216,N_9214);
and U9531 (N_9531,N_9256,N_9393);
or U9532 (N_9532,N_9229,N_9363);
nor U9533 (N_9533,N_9310,N_9393);
nor U9534 (N_9534,N_9292,N_9315);
nor U9535 (N_9535,N_9291,N_9207);
nor U9536 (N_9536,N_9318,N_9294);
and U9537 (N_9537,N_9361,N_9200);
or U9538 (N_9538,N_9274,N_9397);
and U9539 (N_9539,N_9313,N_9357);
nand U9540 (N_9540,N_9382,N_9283);
nand U9541 (N_9541,N_9233,N_9359);
nand U9542 (N_9542,N_9358,N_9340);
or U9543 (N_9543,N_9321,N_9327);
nor U9544 (N_9544,N_9212,N_9201);
or U9545 (N_9545,N_9353,N_9220);
and U9546 (N_9546,N_9243,N_9261);
or U9547 (N_9547,N_9216,N_9264);
nand U9548 (N_9548,N_9212,N_9315);
and U9549 (N_9549,N_9284,N_9235);
nand U9550 (N_9550,N_9292,N_9289);
or U9551 (N_9551,N_9355,N_9399);
and U9552 (N_9552,N_9243,N_9359);
nor U9553 (N_9553,N_9201,N_9264);
and U9554 (N_9554,N_9287,N_9229);
xor U9555 (N_9555,N_9263,N_9306);
nor U9556 (N_9556,N_9337,N_9394);
or U9557 (N_9557,N_9222,N_9233);
nand U9558 (N_9558,N_9271,N_9326);
nor U9559 (N_9559,N_9356,N_9286);
nand U9560 (N_9560,N_9218,N_9275);
nand U9561 (N_9561,N_9272,N_9242);
or U9562 (N_9562,N_9237,N_9225);
nor U9563 (N_9563,N_9232,N_9298);
xnor U9564 (N_9564,N_9327,N_9223);
or U9565 (N_9565,N_9346,N_9224);
nor U9566 (N_9566,N_9243,N_9232);
nor U9567 (N_9567,N_9277,N_9358);
and U9568 (N_9568,N_9296,N_9308);
and U9569 (N_9569,N_9395,N_9248);
or U9570 (N_9570,N_9252,N_9323);
and U9571 (N_9571,N_9201,N_9339);
nor U9572 (N_9572,N_9371,N_9201);
and U9573 (N_9573,N_9341,N_9368);
or U9574 (N_9574,N_9347,N_9232);
xor U9575 (N_9575,N_9239,N_9253);
nand U9576 (N_9576,N_9258,N_9386);
nor U9577 (N_9577,N_9297,N_9292);
nand U9578 (N_9578,N_9386,N_9312);
and U9579 (N_9579,N_9260,N_9332);
and U9580 (N_9580,N_9385,N_9313);
and U9581 (N_9581,N_9368,N_9343);
nor U9582 (N_9582,N_9257,N_9275);
nor U9583 (N_9583,N_9341,N_9282);
or U9584 (N_9584,N_9268,N_9235);
nor U9585 (N_9585,N_9268,N_9325);
and U9586 (N_9586,N_9372,N_9253);
nand U9587 (N_9587,N_9351,N_9316);
nor U9588 (N_9588,N_9391,N_9202);
nor U9589 (N_9589,N_9303,N_9367);
or U9590 (N_9590,N_9359,N_9391);
nand U9591 (N_9591,N_9281,N_9296);
nor U9592 (N_9592,N_9395,N_9252);
nor U9593 (N_9593,N_9340,N_9350);
or U9594 (N_9594,N_9242,N_9301);
xor U9595 (N_9595,N_9289,N_9288);
nand U9596 (N_9596,N_9234,N_9219);
nor U9597 (N_9597,N_9229,N_9382);
xnor U9598 (N_9598,N_9348,N_9352);
or U9599 (N_9599,N_9216,N_9286);
nand U9600 (N_9600,N_9422,N_9462);
nand U9601 (N_9601,N_9464,N_9533);
and U9602 (N_9602,N_9472,N_9437);
and U9603 (N_9603,N_9402,N_9532);
and U9604 (N_9604,N_9482,N_9529);
and U9605 (N_9605,N_9404,N_9421);
nand U9606 (N_9606,N_9561,N_9587);
and U9607 (N_9607,N_9415,N_9526);
nor U9608 (N_9608,N_9591,N_9436);
or U9609 (N_9609,N_9584,N_9566);
nand U9610 (N_9610,N_9523,N_9494);
nor U9611 (N_9611,N_9595,N_9411);
and U9612 (N_9612,N_9508,N_9576);
nand U9613 (N_9613,N_9589,N_9454);
or U9614 (N_9614,N_9434,N_9567);
nor U9615 (N_9615,N_9516,N_9586);
nand U9616 (N_9616,N_9556,N_9548);
nand U9617 (N_9617,N_9480,N_9488);
or U9618 (N_9618,N_9418,N_9505);
nand U9619 (N_9619,N_9545,N_9475);
or U9620 (N_9620,N_9527,N_9493);
or U9621 (N_9621,N_9559,N_9440);
and U9622 (N_9622,N_9400,N_9552);
or U9623 (N_9623,N_9554,N_9524);
nor U9624 (N_9624,N_9507,N_9585);
nor U9625 (N_9625,N_9483,N_9445);
nand U9626 (N_9626,N_9401,N_9407);
and U9627 (N_9627,N_9514,N_9427);
and U9628 (N_9628,N_9497,N_9405);
nand U9629 (N_9629,N_9438,N_9502);
nand U9630 (N_9630,N_9571,N_9594);
xnor U9631 (N_9631,N_9429,N_9439);
or U9632 (N_9632,N_9562,N_9538);
or U9633 (N_9633,N_9456,N_9410);
and U9634 (N_9634,N_9459,N_9460);
or U9635 (N_9635,N_9453,N_9512);
and U9636 (N_9636,N_9536,N_9423);
nor U9637 (N_9637,N_9408,N_9424);
nand U9638 (N_9638,N_9578,N_9542);
and U9639 (N_9639,N_9504,N_9583);
nor U9640 (N_9640,N_9558,N_9458);
nand U9641 (N_9641,N_9485,N_9481);
or U9642 (N_9642,N_9468,N_9515);
or U9643 (N_9643,N_9503,N_9574);
xor U9644 (N_9644,N_9496,N_9581);
or U9645 (N_9645,N_9573,N_9553);
and U9646 (N_9646,N_9593,N_9461);
or U9647 (N_9647,N_9489,N_9565);
or U9648 (N_9648,N_9577,N_9441);
and U9649 (N_9649,N_9406,N_9544);
and U9650 (N_9650,N_9500,N_9549);
nor U9651 (N_9651,N_9444,N_9564);
nand U9652 (N_9652,N_9528,N_9465);
nand U9653 (N_9653,N_9572,N_9484);
or U9654 (N_9654,N_9579,N_9477);
or U9655 (N_9655,N_9448,N_9443);
nor U9656 (N_9656,N_9563,N_9580);
nand U9657 (N_9657,N_9522,N_9539);
nor U9658 (N_9658,N_9520,N_9449);
xnor U9659 (N_9659,N_9432,N_9547);
nor U9660 (N_9660,N_9519,N_9403);
or U9661 (N_9661,N_9499,N_9476);
or U9662 (N_9662,N_9435,N_9451);
nor U9663 (N_9663,N_9555,N_9492);
or U9664 (N_9664,N_9419,N_9551);
and U9665 (N_9665,N_9428,N_9446);
nor U9666 (N_9666,N_9506,N_9412);
nor U9667 (N_9667,N_9513,N_9469);
xor U9668 (N_9668,N_9431,N_9531);
and U9669 (N_9669,N_9582,N_9537);
nand U9670 (N_9670,N_9409,N_9592);
and U9671 (N_9671,N_9479,N_9541);
and U9672 (N_9672,N_9425,N_9597);
and U9673 (N_9673,N_9546,N_9510);
nand U9674 (N_9674,N_9495,N_9534);
or U9675 (N_9675,N_9568,N_9442);
nor U9676 (N_9676,N_9470,N_9414);
nor U9677 (N_9677,N_9413,N_9509);
or U9678 (N_9678,N_9550,N_9457);
or U9679 (N_9679,N_9420,N_9474);
and U9680 (N_9680,N_9569,N_9467);
nor U9681 (N_9681,N_9590,N_9433);
or U9682 (N_9682,N_9540,N_9560);
nor U9683 (N_9683,N_9473,N_9491);
and U9684 (N_9684,N_9530,N_9417);
and U9685 (N_9685,N_9430,N_9450);
or U9686 (N_9686,N_9598,N_9525);
xnor U9687 (N_9687,N_9455,N_9486);
nand U9688 (N_9688,N_9511,N_9487);
and U9689 (N_9689,N_9426,N_9471);
and U9690 (N_9690,N_9521,N_9575);
and U9691 (N_9691,N_9570,N_9557);
nor U9692 (N_9692,N_9501,N_9478);
and U9693 (N_9693,N_9463,N_9588);
nor U9694 (N_9694,N_9517,N_9596);
nand U9695 (N_9695,N_9466,N_9447);
or U9696 (N_9696,N_9452,N_9543);
nor U9697 (N_9697,N_9490,N_9498);
and U9698 (N_9698,N_9518,N_9535);
nand U9699 (N_9699,N_9599,N_9416);
and U9700 (N_9700,N_9567,N_9444);
xnor U9701 (N_9701,N_9578,N_9517);
nor U9702 (N_9702,N_9529,N_9553);
and U9703 (N_9703,N_9589,N_9530);
xor U9704 (N_9704,N_9575,N_9551);
and U9705 (N_9705,N_9587,N_9593);
or U9706 (N_9706,N_9440,N_9460);
nor U9707 (N_9707,N_9451,N_9592);
nor U9708 (N_9708,N_9422,N_9576);
nand U9709 (N_9709,N_9504,N_9490);
nor U9710 (N_9710,N_9596,N_9472);
xnor U9711 (N_9711,N_9581,N_9408);
nand U9712 (N_9712,N_9553,N_9490);
nand U9713 (N_9713,N_9492,N_9414);
and U9714 (N_9714,N_9556,N_9414);
or U9715 (N_9715,N_9486,N_9467);
nand U9716 (N_9716,N_9430,N_9477);
or U9717 (N_9717,N_9582,N_9572);
or U9718 (N_9718,N_9403,N_9524);
or U9719 (N_9719,N_9496,N_9556);
nand U9720 (N_9720,N_9466,N_9510);
xnor U9721 (N_9721,N_9539,N_9574);
nand U9722 (N_9722,N_9426,N_9513);
nor U9723 (N_9723,N_9404,N_9463);
and U9724 (N_9724,N_9422,N_9400);
or U9725 (N_9725,N_9522,N_9496);
nand U9726 (N_9726,N_9460,N_9489);
or U9727 (N_9727,N_9512,N_9432);
and U9728 (N_9728,N_9587,N_9574);
and U9729 (N_9729,N_9482,N_9438);
nor U9730 (N_9730,N_9572,N_9507);
nor U9731 (N_9731,N_9472,N_9466);
nand U9732 (N_9732,N_9551,N_9429);
or U9733 (N_9733,N_9402,N_9514);
or U9734 (N_9734,N_9457,N_9499);
or U9735 (N_9735,N_9539,N_9452);
nor U9736 (N_9736,N_9467,N_9487);
nand U9737 (N_9737,N_9564,N_9449);
and U9738 (N_9738,N_9487,N_9586);
nor U9739 (N_9739,N_9567,N_9497);
xnor U9740 (N_9740,N_9420,N_9595);
or U9741 (N_9741,N_9455,N_9443);
or U9742 (N_9742,N_9443,N_9428);
nand U9743 (N_9743,N_9426,N_9521);
and U9744 (N_9744,N_9586,N_9517);
nand U9745 (N_9745,N_9456,N_9428);
nor U9746 (N_9746,N_9540,N_9442);
and U9747 (N_9747,N_9500,N_9498);
xnor U9748 (N_9748,N_9514,N_9503);
nand U9749 (N_9749,N_9510,N_9513);
nor U9750 (N_9750,N_9437,N_9592);
or U9751 (N_9751,N_9585,N_9573);
and U9752 (N_9752,N_9450,N_9592);
nor U9753 (N_9753,N_9557,N_9430);
xnor U9754 (N_9754,N_9545,N_9435);
xor U9755 (N_9755,N_9588,N_9529);
nand U9756 (N_9756,N_9552,N_9483);
nor U9757 (N_9757,N_9402,N_9430);
and U9758 (N_9758,N_9566,N_9415);
xor U9759 (N_9759,N_9597,N_9591);
nand U9760 (N_9760,N_9459,N_9534);
and U9761 (N_9761,N_9478,N_9521);
and U9762 (N_9762,N_9553,N_9559);
nor U9763 (N_9763,N_9595,N_9509);
nor U9764 (N_9764,N_9488,N_9585);
or U9765 (N_9765,N_9514,N_9517);
or U9766 (N_9766,N_9439,N_9458);
nor U9767 (N_9767,N_9454,N_9438);
and U9768 (N_9768,N_9568,N_9411);
nor U9769 (N_9769,N_9501,N_9465);
nand U9770 (N_9770,N_9538,N_9484);
and U9771 (N_9771,N_9469,N_9531);
xor U9772 (N_9772,N_9426,N_9488);
xor U9773 (N_9773,N_9508,N_9556);
nand U9774 (N_9774,N_9441,N_9437);
or U9775 (N_9775,N_9468,N_9433);
nand U9776 (N_9776,N_9406,N_9472);
and U9777 (N_9777,N_9587,N_9438);
nor U9778 (N_9778,N_9482,N_9587);
xor U9779 (N_9779,N_9477,N_9514);
and U9780 (N_9780,N_9530,N_9519);
nand U9781 (N_9781,N_9423,N_9520);
xnor U9782 (N_9782,N_9579,N_9493);
or U9783 (N_9783,N_9509,N_9440);
nor U9784 (N_9784,N_9425,N_9524);
xor U9785 (N_9785,N_9481,N_9483);
or U9786 (N_9786,N_9400,N_9478);
nand U9787 (N_9787,N_9409,N_9449);
and U9788 (N_9788,N_9450,N_9571);
or U9789 (N_9789,N_9592,N_9414);
nor U9790 (N_9790,N_9556,N_9553);
nor U9791 (N_9791,N_9455,N_9448);
nand U9792 (N_9792,N_9540,N_9429);
nor U9793 (N_9793,N_9433,N_9461);
xor U9794 (N_9794,N_9442,N_9482);
and U9795 (N_9795,N_9452,N_9494);
nor U9796 (N_9796,N_9540,N_9427);
nor U9797 (N_9797,N_9454,N_9582);
xnor U9798 (N_9798,N_9502,N_9558);
or U9799 (N_9799,N_9569,N_9451);
nand U9800 (N_9800,N_9667,N_9760);
and U9801 (N_9801,N_9665,N_9650);
and U9802 (N_9802,N_9682,N_9721);
nor U9803 (N_9803,N_9684,N_9778);
and U9804 (N_9804,N_9748,N_9630);
and U9805 (N_9805,N_9746,N_9625);
or U9806 (N_9806,N_9668,N_9636);
nand U9807 (N_9807,N_9756,N_9716);
nand U9808 (N_9808,N_9754,N_9632);
or U9809 (N_9809,N_9727,N_9734);
and U9810 (N_9810,N_9705,N_9641);
nand U9811 (N_9811,N_9779,N_9612);
nor U9812 (N_9812,N_9611,N_9653);
or U9813 (N_9813,N_9613,N_9732);
nor U9814 (N_9814,N_9792,N_9643);
or U9815 (N_9815,N_9693,N_9725);
or U9816 (N_9816,N_9736,N_9622);
nand U9817 (N_9817,N_9680,N_9752);
xor U9818 (N_9818,N_9769,N_9749);
nand U9819 (N_9819,N_9758,N_9768);
nand U9820 (N_9820,N_9739,N_9678);
and U9821 (N_9821,N_9671,N_9713);
xnor U9822 (N_9822,N_9793,N_9794);
or U9823 (N_9823,N_9652,N_9781);
and U9824 (N_9824,N_9697,N_9692);
and U9825 (N_9825,N_9610,N_9743);
and U9826 (N_9826,N_9762,N_9644);
nand U9827 (N_9827,N_9617,N_9730);
xnor U9828 (N_9828,N_9712,N_9742);
or U9829 (N_9829,N_9688,N_9602);
nor U9830 (N_9830,N_9626,N_9783);
nor U9831 (N_9831,N_9631,N_9658);
nor U9832 (N_9832,N_9745,N_9790);
nor U9833 (N_9833,N_9656,N_9606);
nor U9834 (N_9834,N_9789,N_9798);
and U9835 (N_9835,N_9603,N_9791);
nand U9836 (N_9836,N_9757,N_9700);
nor U9837 (N_9837,N_9696,N_9640);
nand U9838 (N_9838,N_9735,N_9660);
nor U9839 (N_9839,N_9775,N_9724);
and U9840 (N_9840,N_9699,N_9620);
xnor U9841 (N_9841,N_9642,N_9799);
or U9842 (N_9842,N_9689,N_9717);
nor U9843 (N_9843,N_9767,N_9619);
nor U9844 (N_9844,N_9672,N_9635);
nor U9845 (N_9845,N_9627,N_9751);
or U9846 (N_9846,N_9675,N_9659);
nand U9847 (N_9847,N_9608,N_9703);
or U9848 (N_9848,N_9679,N_9629);
nand U9849 (N_9849,N_9763,N_9664);
nor U9850 (N_9850,N_9733,N_9686);
nor U9851 (N_9851,N_9738,N_9681);
nand U9852 (N_9852,N_9764,N_9774);
and U9853 (N_9853,N_9714,N_9655);
and U9854 (N_9854,N_9720,N_9722);
nand U9855 (N_9855,N_9723,N_9624);
and U9856 (N_9856,N_9674,N_9651);
nand U9857 (N_9857,N_9765,N_9607);
nand U9858 (N_9858,N_9601,N_9691);
nand U9859 (N_9859,N_9657,N_9761);
and U9860 (N_9860,N_9729,N_9604);
and U9861 (N_9861,N_9795,N_9628);
nor U9862 (N_9862,N_9662,N_9649);
and U9863 (N_9863,N_9711,N_9605);
and U9864 (N_9864,N_9615,N_9786);
nand U9865 (N_9865,N_9609,N_9646);
xnor U9866 (N_9866,N_9770,N_9747);
nand U9867 (N_9867,N_9788,N_9785);
nor U9868 (N_9868,N_9633,N_9755);
nor U9869 (N_9869,N_9637,N_9704);
nand U9870 (N_9870,N_9673,N_9685);
and U9871 (N_9871,N_9616,N_9690);
nand U9872 (N_9872,N_9740,N_9614);
or U9873 (N_9873,N_9796,N_9787);
nand U9874 (N_9874,N_9694,N_9731);
xor U9875 (N_9875,N_9687,N_9772);
and U9876 (N_9876,N_9695,N_9645);
and U9877 (N_9877,N_9623,N_9710);
or U9878 (N_9878,N_9726,N_9702);
nand U9879 (N_9879,N_9701,N_9737);
nand U9880 (N_9880,N_9719,N_9750);
nand U9881 (N_9881,N_9661,N_9647);
or U9882 (N_9882,N_9654,N_9776);
nand U9883 (N_9883,N_9669,N_9784);
nor U9884 (N_9884,N_9666,N_9663);
xor U9885 (N_9885,N_9759,N_9780);
nand U9886 (N_9886,N_9634,N_9741);
or U9887 (N_9887,N_9708,N_9773);
or U9888 (N_9888,N_9766,N_9777);
or U9889 (N_9889,N_9744,N_9753);
nor U9890 (N_9890,N_9677,N_9706);
xnor U9891 (N_9891,N_9600,N_9715);
or U9892 (N_9892,N_9728,N_9707);
and U9893 (N_9893,N_9698,N_9683);
nand U9894 (N_9894,N_9676,N_9618);
nor U9895 (N_9895,N_9709,N_9621);
or U9896 (N_9896,N_9797,N_9771);
or U9897 (N_9897,N_9648,N_9670);
nand U9898 (N_9898,N_9639,N_9638);
nand U9899 (N_9899,N_9718,N_9782);
nor U9900 (N_9900,N_9749,N_9659);
or U9901 (N_9901,N_9774,N_9762);
xor U9902 (N_9902,N_9621,N_9799);
and U9903 (N_9903,N_9605,N_9780);
and U9904 (N_9904,N_9766,N_9658);
xor U9905 (N_9905,N_9640,N_9772);
xor U9906 (N_9906,N_9775,N_9776);
and U9907 (N_9907,N_9685,N_9710);
or U9908 (N_9908,N_9745,N_9714);
nor U9909 (N_9909,N_9674,N_9655);
or U9910 (N_9910,N_9697,N_9614);
and U9911 (N_9911,N_9750,N_9646);
nand U9912 (N_9912,N_9705,N_9701);
and U9913 (N_9913,N_9622,N_9611);
nand U9914 (N_9914,N_9787,N_9661);
nor U9915 (N_9915,N_9716,N_9702);
or U9916 (N_9916,N_9719,N_9692);
nor U9917 (N_9917,N_9711,N_9652);
or U9918 (N_9918,N_9760,N_9720);
nor U9919 (N_9919,N_9726,N_9787);
and U9920 (N_9920,N_9735,N_9608);
or U9921 (N_9921,N_9753,N_9788);
and U9922 (N_9922,N_9602,N_9752);
and U9923 (N_9923,N_9688,N_9652);
and U9924 (N_9924,N_9720,N_9645);
and U9925 (N_9925,N_9665,N_9628);
and U9926 (N_9926,N_9798,N_9700);
nor U9927 (N_9927,N_9747,N_9736);
or U9928 (N_9928,N_9709,N_9686);
nand U9929 (N_9929,N_9780,N_9648);
and U9930 (N_9930,N_9775,N_9712);
nor U9931 (N_9931,N_9739,N_9636);
and U9932 (N_9932,N_9621,N_9633);
or U9933 (N_9933,N_9769,N_9670);
and U9934 (N_9934,N_9707,N_9775);
nand U9935 (N_9935,N_9779,N_9767);
xor U9936 (N_9936,N_9651,N_9726);
or U9937 (N_9937,N_9796,N_9771);
nand U9938 (N_9938,N_9637,N_9772);
nand U9939 (N_9939,N_9782,N_9673);
nor U9940 (N_9940,N_9702,N_9749);
or U9941 (N_9941,N_9669,N_9741);
and U9942 (N_9942,N_9780,N_9630);
nand U9943 (N_9943,N_9768,N_9689);
or U9944 (N_9944,N_9651,N_9714);
nand U9945 (N_9945,N_9615,N_9666);
nor U9946 (N_9946,N_9657,N_9658);
nand U9947 (N_9947,N_9710,N_9695);
and U9948 (N_9948,N_9627,N_9623);
or U9949 (N_9949,N_9671,N_9614);
nand U9950 (N_9950,N_9794,N_9654);
or U9951 (N_9951,N_9644,N_9741);
nand U9952 (N_9952,N_9718,N_9604);
nor U9953 (N_9953,N_9775,N_9700);
xnor U9954 (N_9954,N_9621,N_9742);
nor U9955 (N_9955,N_9621,N_9720);
xnor U9956 (N_9956,N_9704,N_9661);
nand U9957 (N_9957,N_9643,N_9755);
or U9958 (N_9958,N_9702,N_9689);
nor U9959 (N_9959,N_9634,N_9611);
nand U9960 (N_9960,N_9641,N_9659);
nand U9961 (N_9961,N_9613,N_9660);
xnor U9962 (N_9962,N_9788,N_9645);
nor U9963 (N_9963,N_9610,N_9668);
nand U9964 (N_9964,N_9776,N_9788);
nor U9965 (N_9965,N_9706,N_9616);
xnor U9966 (N_9966,N_9701,N_9627);
and U9967 (N_9967,N_9730,N_9677);
nor U9968 (N_9968,N_9735,N_9705);
nor U9969 (N_9969,N_9601,N_9694);
nor U9970 (N_9970,N_9760,N_9737);
xor U9971 (N_9971,N_9637,N_9621);
xor U9972 (N_9972,N_9797,N_9633);
and U9973 (N_9973,N_9772,N_9716);
nor U9974 (N_9974,N_9693,N_9757);
nor U9975 (N_9975,N_9735,N_9625);
nand U9976 (N_9976,N_9749,N_9670);
or U9977 (N_9977,N_9796,N_9723);
or U9978 (N_9978,N_9640,N_9606);
nor U9979 (N_9979,N_9717,N_9795);
nor U9980 (N_9980,N_9679,N_9644);
xor U9981 (N_9981,N_9696,N_9768);
nor U9982 (N_9982,N_9799,N_9628);
nor U9983 (N_9983,N_9656,N_9609);
nor U9984 (N_9984,N_9762,N_9740);
and U9985 (N_9985,N_9606,N_9770);
xor U9986 (N_9986,N_9706,N_9667);
nor U9987 (N_9987,N_9677,N_9685);
nand U9988 (N_9988,N_9640,N_9685);
nor U9989 (N_9989,N_9608,N_9778);
xnor U9990 (N_9990,N_9715,N_9601);
nor U9991 (N_9991,N_9672,N_9750);
nand U9992 (N_9992,N_9696,N_9684);
or U9993 (N_9993,N_9793,N_9792);
nand U9994 (N_9994,N_9639,N_9652);
nand U9995 (N_9995,N_9731,N_9749);
nor U9996 (N_9996,N_9763,N_9608);
and U9997 (N_9997,N_9744,N_9781);
nand U9998 (N_9998,N_9740,N_9603);
and U9999 (N_9999,N_9675,N_9671);
or UO_0 (O_0,N_9958,N_9995);
xnor UO_1 (O_1,N_9936,N_9887);
and UO_2 (O_2,N_9976,N_9952);
and UO_3 (O_3,N_9909,N_9908);
nand UO_4 (O_4,N_9962,N_9959);
nand UO_5 (O_5,N_9918,N_9928);
nand UO_6 (O_6,N_9849,N_9913);
or UO_7 (O_7,N_9807,N_9864);
and UO_8 (O_8,N_9815,N_9964);
and UO_9 (O_9,N_9945,N_9892);
and UO_10 (O_10,N_9949,N_9927);
nand UO_11 (O_11,N_9824,N_9810);
nor UO_12 (O_12,N_9953,N_9894);
and UO_13 (O_13,N_9867,N_9893);
xor UO_14 (O_14,N_9983,N_9970);
nor UO_15 (O_15,N_9941,N_9873);
nor UO_16 (O_16,N_9984,N_9842);
or UO_17 (O_17,N_9989,N_9811);
and UO_18 (O_18,N_9866,N_9858);
nand UO_19 (O_19,N_9971,N_9847);
xnor UO_20 (O_20,N_9802,N_9939);
and UO_21 (O_21,N_9933,N_9967);
or UO_22 (O_22,N_9957,N_9820);
xor UO_23 (O_23,N_9818,N_9865);
or UO_24 (O_24,N_9803,N_9999);
nand UO_25 (O_25,N_9910,N_9934);
or UO_26 (O_26,N_9924,N_9821);
nor UO_27 (O_27,N_9833,N_9950);
nor UO_28 (O_28,N_9823,N_9863);
nand UO_29 (O_29,N_9854,N_9940);
nand UO_30 (O_30,N_9897,N_9828);
nor UO_31 (O_31,N_9961,N_9981);
nand UO_32 (O_32,N_9878,N_9982);
and UO_33 (O_33,N_9882,N_9948);
nor UO_34 (O_34,N_9923,N_9980);
nand UO_35 (O_35,N_9972,N_9921);
nor UO_36 (O_36,N_9840,N_9917);
and UO_37 (O_37,N_9951,N_9969);
and UO_38 (O_38,N_9929,N_9914);
or UO_39 (O_39,N_9920,N_9903);
nor UO_40 (O_40,N_9975,N_9832);
or UO_41 (O_41,N_9905,N_9956);
or UO_42 (O_42,N_9819,N_9896);
and UO_43 (O_43,N_9937,N_9907);
xor UO_44 (O_44,N_9871,N_9835);
nand UO_45 (O_45,N_9987,N_9986);
and UO_46 (O_46,N_9895,N_9862);
nand UO_47 (O_47,N_9966,N_9998);
and UO_48 (O_48,N_9960,N_9991);
and UO_49 (O_49,N_9801,N_9898);
or UO_50 (O_50,N_9834,N_9845);
and UO_51 (O_51,N_9841,N_9994);
nor UO_52 (O_52,N_9804,N_9944);
and UO_53 (O_53,N_9859,N_9968);
or UO_54 (O_54,N_9925,N_9861);
xor UO_55 (O_55,N_9906,N_9880);
nand UO_56 (O_56,N_9839,N_9800);
and UO_57 (O_57,N_9851,N_9881);
and UO_58 (O_58,N_9872,N_9963);
or UO_59 (O_59,N_9827,N_9926);
and UO_60 (O_60,N_9808,N_9837);
or UO_61 (O_61,N_9901,N_9955);
nand UO_62 (O_62,N_9855,N_9974);
nand UO_63 (O_63,N_9805,N_9826);
and UO_64 (O_64,N_9992,N_9943);
nor UO_65 (O_65,N_9813,N_9990);
nand UO_66 (O_66,N_9922,N_9935);
nor UO_67 (O_67,N_9916,N_9877);
or UO_68 (O_68,N_9988,N_9996);
xor UO_69 (O_69,N_9942,N_9930);
nor UO_70 (O_70,N_9822,N_9856);
and UO_71 (O_71,N_9812,N_9890);
or UO_72 (O_72,N_9829,N_9904);
or UO_73 (O_73,N_9836,N_9997);
nor UO_74 (O_74,N_9912,N_9915);
or UO_75 (O_75,N_9938,N_9838);
nand UO_76 (O_76,N_9993,N_9816);
or UO_77 (O_77,N_9900,N_9830);
nand UO_78 (O_78,N_9883,N_9831);
nand UO_79 (O_79,N_9853,N_9884);
and UO_80 (O_80,N_9985,N_9846);
or UO_81 (O_81,N_9844,N_9879);
and UO_82 (O_82,N_9806,N_9911);
xnor UO_83 (O_83,N_9978,N_9874);
nor UO_84 (O_84,N_9886,N_9852);
nand UO_85 (O_85,N_9848,N_9947);
xor UO_86 (O_86,N_9979,N_9977);
nand UO_87 (O_87,N_9965,N_9932);
and UO_88 (O_88,N_9902,N_9857);
nand UO_89 (O_89,N_9899,N_9868);
or UO_90 (O_90,N_9825,N_9869);
and UO_91 (O_91,N_9889,N_9891);
nand UO_92 (O_92,N_9843,N_9885);
xor UO_93 (O_93,N_9870,N_9814);
nor UO_94 (O_94,N_9931,N_9973);
nor UO_95 (O_95,N_9860,N_9809);
and UO_96 (O_96,N_9919,N_9888);
nor UO_97 (O_97,N_9876,N_9875);
nand UO_98 (O_98,N_9946,N_9954);
or UO_99 (O_99,N_9817,N_9850);
nor UO_100 (O_100,N_9912,N_9866);
nor UO_101 (O_101,N_9870,N_9830);
nand UO_102 (O_102,N_9974,N_9859);
nor UO_103 (O_103,N_9894,N_9970);
xnor UO_104 (O_104,N_9901,N_9959);
or UO_105 (O_105,N_9997,N_9931);
nand UO_106 (O_106,N_9984,N_9859);
nor UO_107 (O_107,N_9991,N_9881);
and UO_108 (O_108,N_9857,N_9948);
nand UO_109 (O_109,N_9911,N_9809);
nand UO_110 (O_110,N_9854,N_9911);
nor UO_111 (O_111,N_9915,N_9883);
nor UO_112 (O_112,N_9917,N_9962);
and UO_113 (O_113,N_9957,N_9818);
nor UO_114 (O_114,N_9860,N_9828);
and UO_115 (O_115,N_9800,N_9917);
nor UO_116 (O_116,N_9845,N_9824);
nand UO_117 (O_117,N_9980,N_9884);
or UO_118 (O_118,N_9878,N_9943);
nor UO_119 (O_119,N_9908,N_9977);
nor UO_120 (O_120,N_9905,N_9874);
xor UO_121 (O_121,N_9895,N_9855);
nor UO_122 (O_122,N_9983,N_9944);
nand UO_123 (O_123,N_9818,N_9929);
nand UO_124 (O_124,N_9833,N_9936);
nand UO_125 (O_125,N_9803,N_9965);
nand UO_126 (O_126,N_9826,N_9994);
or UO_127 (O_127,N_9971,N_9978);
or UO_128 (O_128,N_9964,N_9886);
nor UO_129 (O_129,N_9966,N_9869);
nand UO_130 (O_130,N_9983,N_9921);
nand UO_131 (O_131,N_9961,N_9878);
nand UO_132 (O_132,N_9805,N_9950);
nor UO_133 (O_133,N_9909,N_9826);
nand UO_134 (O_134,N_9859,N_9950);
nand UO_135 (O_135,N_9818,N_9943);
nor UO_136 (O_136,N_9989,N_9925);
or UO_137 (O_137,N_9842,N_9849);
or UO_138 (O_138,N_9932,N_9917);
xnor UO_139 (O_139,N_9964,N_9996);
or UO_140 (O_140,N_9896,N_9926);
xnor UO_141 (O_141,N_9815,N_9922);
or UO_142 (O_142,N_9840,N_9982);
and UO_143 (O_143,N_9960,N_9913);
nor UO_144 (O_144,N_9869,N_9868);
nand UO_145 (O_145,N_9927,N_9974);
or UO_146 (O_146,N_9854,N_9873);
or UO_147 (O_147,N_9818,N_9857);
nor UO_148 (O_148,N_9908,N_9969);
nor UO_149 (O_149,N_9937,N_9961);
nor UO_150 (O_150,N_9976,N_9902);
nand UO_151 (O_151,N_9918,N_9914);
and UO_152 (O_152,N_9843,N_9911);
nand UO_153 (O_153,N_9917,N_9877);
and UO_154 (O_154,N_9925,N_9809);
and UO_155 (O_155,N_9964,N_9948);
and UO_156 (O_156,N_9924,N_9885);
and UO_157 (O_157,N_9963,N_9933);
and UO_158 (O_158,N_9971,N_9816);
nand UO_159 (O_159,N_9827,N_9825);
nand UO_160 (O_160,N_9918,N_9937);
nand UO_161 (O_161,N_9872,N_9930);
nand UO_162 (O_162,N_9830,N_9808);
nand UO_163 (O_163,N_9850,N_9932);
or UO_164 (O_164,N_9973,N_9980);
nand UO_165 (O_165,N_9817,N_9873);
and UO_166 (O_166,N_9924,N_9947);
nand UO_167 (O_167,N_9836,N_9995);
and UO_168 (O_168,N_9981,N_9979);
nand UO_169 (O_169,N_9828,N_9976);
and UO_170 (O_170,N_9915,N_9932);
nor UO_171 (O_171,N_9840,N_9905);
or UO_172 (O_172,N_9947,N_9802);
and UO_173 (O_173,N_9855,N_9896);
and UO_174 (O_174,N_9914,N_9955);
or UO_175 (O_175,N_9851,N_9999);
or UO_176 (O_176,N_9997,N_9809);
and UO_177 (O_177,N_9998,N_9993);
xnor UO_178 (O_178,N_9891,N_9928);
or UO_179 (O_179,N_9968,N_9836);
nand UO_180 (O_180,N_9815,N_9810);
and UO_181 (O_181,N_9823,N_9913);
nand UO_182 (O_182,N_9904,N_9997);
xor UO_183 (O_183,N_9997,N_9803);
or UO_184 (O_184,N_9865,N_9912);
xor UO_185 (O_185,N_9877,N_9915);
or UO_186 (O_186,N_9861,N_9807);
or UO_187 (O_187,N_9863,N_9926);
and UO_188 (O_188,N_9883,N_9862);
or UO_189 (O_189,N_9844,N_9860);
or UO_190 (O_190,N_9951,N_9882);
nand UO_191 (O_191,N_9936,N_9963);
or UO_192 (O_192,N_9946,N_9840);
nand UO_193 (O_193,N_9830,N_9965);
xnor UO_194 (O_194,N_9843,N_9825);
and UO_195 (O_195,N_9893,N_9976);
nand UO_196 (O_196,N_9956,N_9839);
nand UO_197 (O_197,N_9856,N_9940);
nand UO_198 (O_198,N_9934,N_9884);
or UO_199 (O_199,N_9952,N_9957);
nand UO_200 (O_200,N_9803,N_9842);
nand UO_201 (O_201,N_9954,N_9904);
or UO_202 (O_202,N_9805,N_9855);
nor UO_203 (O_203,N_9951,N_9956);
xor UO_204 (O_204,N_9974,N_9835);
or UO_205 (O_205,N_9892,N_9870);
or UO_206 (O_206,N_9982,N_9913);
and UO_207 (O_207,N_9937,N_9965);
nand UO_208 (O_208,N_9987,N_9993);
nor UO_209 (O_209,N_9806,N_9970);
nand UO_210 (O_210,N_9935,N_9855);
nor UO_211 (O_211,N_9916,N_9801);
or UO_212 (O_212,N_9909,N_9885);
and UO_213 (O_213,N_9926,N_9879);
nand UO_214 (O_214,N_9924,N_9984);
nor UO_215 (O_215,N_9912,N_9804);
nor UO_216 (O_216,N_9855,N_9948);
nor UO_217 (O_217,N_9904,N_9811);
or UO_218 (O_218,N_9866,N_9997);
nand UO_219 (O_219,N_9829,N_9963);
nor UO_220 (O_220,N_9840,N_9993);
nand UO_221 (O_221,N_9832,N_9815);
nand UO_222 (O_222,N_9882,N_9945);
or UO_223 (O_223,N_9918,N_9929);
nand UO_224 (O_224,N_9876,N_9834);
nand UO_225 (O_225,N_9857,N_9909);
xor UO_226 (O_226,N_9834,N_9963);
or UO_227 (O_227,N_9810,N_9866);
or UO_228 (O_228,N_9990,N_9865);
or UO_229 (O_229,N_9951,N_9947);
nand UO_230 (O_230,N_9829,N_9876);
and UO_231 (O_231,N_9884,N_9987);
nor UO_232 (O_232,N_9827,N_9953);
xnor UO_233 (O_233,N_9887,N_9830);
xnor UO_234 (O_234,N_9917,N_9976);
nand UO_235 (O_235,N_9982,N_9911);
nand UO_236 (O_236,N_9831,N_9937);
and UO_237 (O_237,N_9874,N_9989);
nand UO_238 (O_238,N_9988,N_9876);
nand UO_239 (O_239,N_9890,N_9991);
nand UO_240 (O_240,N_9875,N_9938);
nand UO_241 (O_241,N_9955,N_9879);
xor UO_242 (O_242,N_9887,N_9875);
xnor UO_243 (O_243,N_9905,N_9842);
nor UO_244 (O_244,N_9941,N_9993);
xnor UO_245 (O_245,N_9994,N_9925);
nand UO_246 (O_246,N_9884,N_9993);
xnor UO_247 (O_247,N_9802,N_9804);
xor UO_248 (O_248,N_9947,N_9827);
nand UO_249 (O_249,N_9891,N_9882);
nor UO_250 (O_250,N_9993,N_9838);
nor UO_251 (O_251,N_9977,N_9809);
xor UO_252 (O_252,N_9983,N_9818);
nor UO_253 (O_253,N_9930,N_9845);
and UO_254 (O_254,N_9897,N_9896);
nand UO_255 (O_255,N_9924,N_9868);
or UO_256 (O_256,N_9999,N_9974);
nand UO_257 (O_257,N_9899,N_9957);
and UO_258 (O_258,N_9844,N_9958);
nand UO_259 (O_259,N_9860,N_9811);
nor UO_260 (O_260,N_9876,N_9893);
nor UO_261 (O_261,N_9997,N_9817);
nor UO_262 (O_262,N_9812,N_9982);
nand UO_263 (O_263,N_9912,N_9859);
nor UO_264 (O_264,N_9983,N_9883);
nand UO_265 (O_265,N_9903,N_9939);
nand UO_266 (O_266,N_9858,N_9814);
and UO_267 (O_267,N_9952,N_9934);
nand UO_268 (O_268,N_9860,N_9868);
nor UO_269 (O_269,N_9951,N_9817);
xor UO_270 (O_270,N_9968,N_9801);
nor UO_271 (O_271,N_9815,N_9862);
and UO_272 (O_272,N_9835,N_9886);
xnor UO_273 (O_273,N_9926,N_9885);
nor UO_274 (O_274,N_9878,N_9956);
and UO_275 (O_275,N_9918,N_9838);
nand UO_276 (O_276,N_9948,N_9837);
xnor UO_277 (O_277,N_9865,N_9951);
and UO_278 (O_278,N_9901,N_9892);
nor UO_279 (O_279,N_9864,N_9948);
and UO_280 (O_280,N_9902,N_9850);
xnor UO_281 (O_281,N_9812,N_9903);
or UO_282 (O_282,N_9889,N_9944);
nand UO_283 (O_283,N_9912,N_9843);
nand UO_284 (O_284,N_9929,N_9948);
or UO_285 (O_285,N_9903,N_9886);
or UO_286 (O_286,N_9914,N_9931);
nor UO_287 (O_287,N_9874,N_9820);
xor UO_288 (O_288,N_9810,N_9835);
nor UO_289 (O_289,N_9968,N_9991);
or UO_290 (O_290,N_9864,N_9945);
and UO_291 (O_291,N_9829,N_9931);
nor UO_292 (O_292,N_9850,N_9875);
or UO_293 (O_293,N_9917,N_9834);
and UO_294 (O_294,N_9853,N_9911);
nand UO_295 (O_295,N_9966,N_9856);
or UO_296 (O_296,N_9870,N_9924);
nand UO_297 (O_297,N_9908,N_9919);
nand UO_298 (O_298,N_9818,N_9836);
xnor UO_299 (O_299,N_9907,N_9880);
or UO_300 (O_300,N_9821,N_9954);
or UO_301 (O_301,N_9921,N_9994);
xnor UO_302 (O_302,N_9824,N_9840);
or UO_303 (O_303,N_9902,N_9822);
and UO_304 (O_304,N_9842,N_9854);
nor UO_305 (O_305,N_9894,N_9900);
nand UO_306 (O_306,N_9839,N_9892);
or UO_307 (O_307,N_9928,N_9889);
nor UO_308 (O_308,N_9944,N_9980);
and UO_309 (O_309,N_9961,N_9955);
or UO_310 (O_310,N_9873,N_9861);
nand UO_311 (O_311,N_9900,N_9969);
and UO_312 (O_312,N_9804,N_9838);
and UO_313 (O_313,N_9854,N_9933);
or UO_314 (O_314,N_9801,N_9985);
xnor UO_315 (O_315,N_9926,N_9929);
nor UO_316 (O_316,N_9836,N_9876);
xnor UO_317 (O_317,N_9863,N_9900);
xor UO_318 (O_318,N_9879,N_9936);
xnor UO_319 (O_319,N_9938,N_9837);
or UO_320 (O_320,N_9878,N_9978);
nor UO_321 (O_321,N_9974,N_9893);
or UO_322 (O_322,N_9979,N_9920);
nand UO_323 (O_323,N_9808,N_9910);
or UO_324 (O_324,N_9922,N_9873);
nor UO_325 (O_325,N_9855,N_9883);
xnor UO_326 (O_326,N_9925,N_9884);
or UO_327 (O_327,N_9902,N_9999);
nand UO_328 (O_328,N_9933,N_9943);
and UO_329 (O_329,N_9961,N_9949);
nor UO_330 (O_330,N_9943,N_9863);
xor UO_331 (O_331,N_9802,N_9893);
or UO_332 (O_332,N_9918,N_9921);
nand UO_333 (O_333,N_9912,N_9809);
nand UO_334 (O_334,N_9928,N_9897);
or UO_335 (O_335,N_9991,N_9822);
nand UO_336 (O_336,N_9915,N_9802);
nand UO_337 (O_337,N_9923,N_9842);
or UO_338 (O_338,N_9831,N_9986);
and UO_339 (O_339,N_9847,N_9915);
and UO_340 (O_340,N_9811,N_9805);
or UO_341 (O_341,N_9932,N_9994);
nand UO_342 (O_342,N_9930,N_9868);
or UO_343 (O_343,N_9998,N_9985);
and UO_344 (O_344,N_9978,N_9923);
nor UO_345 (O_345,N_9846,N_9958);
or UO_346 (O_346,N_9907,N_9890);
or UO_347 (O_347,N_9969,N_9882);
nor UO_348 (O_348,N_9811,N_9849);
and UO_349 (O_349,N_9954,N_9800);
and UO_350 (O_350,N_9910,N_9829);
or UO_351 (O_351,N_9937,N_9852);
and UO_352 (O_352,N_9899,N_9839);
or UO_353 (O_353,N_9826,N_9942);
or UO_354 (O_354,N_9957,N_9867);
or UO_355 (O_355,N_9955,N_9986);
nand UO_356 (O_356,N_9821,N_9971);
nor UO_357 (O_357,N_9805,N_9880);
or UO_358 (O_358,N_9930,N_9807);
and UO_359 (O_359,N_9814,N_9842);
nor UO_360 (O_360,N_9976,N_9938);
nand UO_361 (O_361,N_9845,N_9837);
or UO_362 (O_362,N_9810,N_9944);
nor UO_363 (O_363,N_9874,N_9960);
nor UO_364 (O_364,N_9926,N_9882);
and UO_365 (O_365,N_9994,N_9970);
or UO_366 (O_366,N_9924,N_9943);
and UO_367 (O_367,N_9833,N_9994);
nor UO_368 (O_368,N_9800,N_9976);
xnor UO_369 (O_369,N_9966,N_9805);
nand UO_370 (O_370,N_9843,N_9823);
and UO_371 (O_371,N_9875,N_9960);
and UO_372 (O_372,N_9844,N_9851);
nand UO_373 (O_373,N_9960,N_9881);
nand UO_374 (O_374,N_9948,N_9945);
nor UO_375 (O_375,N_9816,N_9803);
nor UO_376 (O_376,N_9862,N_9971);
or UO_377 (O_377,N_9864,N_9824);
nor UO_378 (O_378,N_9916,N_9976);
nand UO_379 (O_379,N_9971,N_9898);
or UO_380 (O_380,N_9969,N_9873);
or UO_381 (O_381,N_9886,N_9805);
nand UO_382 (O_382,N_9954,N_9829);
and UO_383 (O_383,N_9989,N_9982);
and UO_384 (O_384,N_9809,N_9906);
or UO_385 (O_385,N_9859,N_9807);
and UO_386 (O_386,N_9899,N_9844);
nor UO_387 (O_387,N_9902,N_9938);
or UO_388 (O_388,N_9993,N_9947);
xnor UO_389 (O_389,N_9933,N_9924);
and UO_390 (O_390,N_9849,N_9869);
nor UO_391 (O_391,N_9900,N_9901);
or UO_392 (O_392,N_9852,N_9933);
and UO_393 (O_393,N_9900,N_9959);
nor UO_394 (O_394,N_9998,N_9927);
nand UO_395 (O_395,N_9872,N_9849);
nand UO_396 (O_396,N_9873,N_9822);
and UO_397 (O_397,N_9880,N_9888);
or UO_398 (O_398,N_9839,N_9882);
or UO_399 (O_399,N_9811,N_9978);
or UO_400 (O_400,N_9847,N_9998);
nor UO_401 (O_401,N_9967,N_9931);
or UO_402 (O_402,N_9825,N_9902);
nor UO_403 (O_403,N_9902,N_9833);
or UO_404 (O_404,N_9978,N_9935);
xor UO_405 (O_405,N_9919,N_9836);
nor UO_406 (O_406,N_9813,N_9867);
xor UO_407 (O_407,N_9922,N_9944);
xnor UO_408 (O_408,N_9832,N_9986);
or UO_409 (O_409,N_9845,N_9874);
and UO_410 (O_410,N_9850,N_9947);
or UO_411 (O_411,N_9959,N_9910);
or UO_412 (O_412,N_9868,N_9914);
xor UO_413 (O_413,N_9848,N_9863);
nand UO_414 (O_414,N_9809,N_9966);
or UO_415 (O_415,N_9854,N_9979);
nand UO_416 (O_416,N_9934,N_9936);
nor UO_417 (O_417,N_9828,N_9896);
nand UO_418 (O_418,N_9801,N_9952);
xnor UO_419 (O_419,N_9937,N_9807);
nor UO_420 (O_420,N_9815,N_9989);
and UO_421 (O_421,N_9867,N_9969);
nor UO_422 (O_422,N_9908,N_9957);
or UO_423 (O_423,N_9841,N_9873);
or UO_424 (O_424,N_9854,N_9994);
xor UO_425 (O_425,N_9929,N_9901);
nand UO_426 (O_426,N_9819,N_9807);
and UO_427 (O_427,N_9862,N_9995);
and UO_428 (O_428,N_9980,N_9948);
nand UO_429 (O_429,N_9925,N_9857);
or UO_430 (O_430,N_9808,N_9918);
nor UO_431 (O_431,N_9992,N_9886);
and UO_432 (O_432,N_9810,N_9890);
and UO_433 (O_433,N_9826,N_9827);
or UO_434 (O_434,N_9977,N_9964);
or UO_435 (O_435,N_9914,N_9840);
xor UO_436 (O_436,N_9977,N_9993);
nand UO_437 (O_437,N_9919,N_9951);
or UO_438 (O_438,N_9958,N_9990);
nand UO_439 (O_439,N_9838,N_9989);
nor UO_440 (O_440,N_9963,N_9889);
nand UO_441 (O_441,N_9850,N_9901);
xnor UO_442 (O_442,N_9891,N_9826);
nand UO_443 (O_443,N_9818,N_9918);
or UO_444 (O_444,N_9934,N_9924);
nor UO_445 (O_445,N_9987,N_9943);
nand UO_446 (O_446,N_9953,N_9876);
or UO_447 (O_447,N_9807,N_9831);
xnor UO_448 (O_448,N_9982,N_9803);
nand UO_449 (O_449,N_9959,N_9899);
nand UO_450 (O_450,N_9974,N_9875);
nand UO_451 (O_451,N_9985,N_9964);
or UO_452 (O_452,N_9867,N_9973);
and UO_453 (O_453,N_9891,N_9807);
and UO_454 (O_454,N_9901,N_9823);
nor UO_455 (O_455,N_9910,N_9880);
or UO_456 (O_456,N_9955,N_9939);
nand UO_457 (O_457,N_9994,N_9918);
nand UO_458 (O_458,N_9890,N_9845);
nor UO_459 (O_459,N_9804,N_9911);
or UO_460 (O_460,N_9998,N_9968);
nand UO_461 (O_461,N_9806,N_9965);
nand UO_462 (O_462,N_9955,N_9847);
xnor UO_463 (O_463,N_9832,N_9829);
nand UO_464 (O_464,N_9957,N_9993);
nor UO_465 (O_465,N_9914,N_9870);
or UO_466 (O_466,N_9801,N_9943);
nand UO_467 (O_467,N_9921,N_9880);
or UO_468 (O_468,N_9992,N_9980);
or UO_469 (O_469,N_9929,N_9861);
or UO_470 (O_470,N_9847,N_9966);
nand UO_471 (O_471,N_9934,N_9811);
and UO_472 (O_472,N_9847,N_9912);
xor UO_473 (O_473,N_9884,N_9843);
or UO_474 (O_474,N_9857,N_9954);
nand UO_475 (O_475,N_9804,N_9817);
or UO_476 (O_476,N_9921,N_9911);
nand UO_477 (O_477,N_9804,N_9833);
nand UO_478 (O_478,N_9890,N_9962);
or UO_479 (O_479,N_9857,N_9974);
and UO_480 (O_480,N_9869,N_9986);
xnor UO_481 (O_481,N_9839,N_9971);
and UO_482 (O_482,N_9811,N_9896);
or UO_483 (O_483,N_9805,N_9931);
or UO_484 (O_484,N_9943,N_9997);
nor UO_485 (O_485,N_9982,N_9859);
nand UO_486 (O_486,N_9871,N_9919);
or UO_487 (O_487,N_9949,N_9924);
and UO_488 (O_488,N_9959,N_9929);
nor UO_489 (O_489,N_9913,N_9818);
nand UO_490 (O_490,N_9955,N_9877);
or UO_491 (O_491,N_9853,N_9878);
nand UO_492 (O_492,N_9965,N_9986);
and UO_493 (O_493,N_9862,N_9913);
and UO_494 (O_494,N_9844,N_9908);
nand UO_495 (O_495,N_9866,N_9971);
or UO_496 (O_496,N_9919,N_9966);
nor UO_497 (O_497,N_9845,N_9913);
nor UO_498 (O_498,N_9983,N_9950);
and UO_499 (O_499,N_9826,N_9936);
nand UO_500 (O_500,N_9806,N_9982);
or UO_501 (O_501,N_9822,N_9803);
or UO_502 (O_502,N_9925,N_9998);
and UO_503 (O_503,N_9931,N_9959);
nand UO_504 (O_504,N_9946,N_9998);
xnor UO_505 (O_505,N_9992,N_9897);
or UO_506 (O_506,N_9994,N_9979);
nor UO_507 (O_507,N_9868,N_9873);
and UO_508 (O_508,N_9970,N_9984);
nand UO_509 (O_509,N_9850,N_9893);
nand UO_510 (O_510,N_9887,N_9962);
and UO_511 (O_511,N_9915,N_9923);
xnor UO_512 (O_512,N_9980,N_9905);
and UO_513 (O_513,N_9922,N_9983);
and UO_514 (O_514,N_9914,N_9959);
or UO_515 (O_515,N_9948,N_9973);
nor UO_516 (O_516,N_9960,N_9832);
xor UO_517 (O_517,N_9984,N_9979);
or UO_518 (O_518,N_9839,N_9939);
nor UO_519 (O_519,N_9903,N_9839);
nor UO_520 (O_520,N_9861,N_9958);
and UO_521 (O_521,N_9846,N_9929);
xnor UO_522 (O_522,N_9991,N_9895);
nand UO_523 (O_523,N_9886,N_9997);
nand UO_524 (O_524,N_9887,N_9837);
or UO_525 (O_525,N_9819,N_9881);
nand UO_526 (O_526,N_9880,N_9803);
nor UO_527 (O_527,N_9990,N_9942);
nor UO_528 (O_528,N_9809,N_9998);
or UO_529 (O_529,N_9905,N_9810);
and UO_530 (O_530,N_9981,N_9964);
and UO_531 (O_531,N_9863,N_9833);
or UO_532 (O_532,N_9996,N_9829);
nand UO_533 (O_533,N_9958,N_9874);
or UO_534 (O_534,N_9875,N_9970);
and UO_535 (O_535,N_9845,N_9826);
and UO_536 (O_536,N_9807,N_9824);
xor UO_537 (O_537,N_9983,N_9962);
nand UO_538 (O_538,N_9840,N_9830);
and UO_539 (O_539,N_9847,N_9911);
xnor UO_540 (O_540,N_9971,N_9991);
nor UO_541 (O_541,N_9851,N_9835);
and UO_542 (O_542,N_9828,N_9955);
nor UO_543 (O_543,N_9918,N_9872);
or UO_544 (O_544,N_9892,N_9916);
nor UO_545 (O_545,N_9990,N_9841);
xnor UO_546 (O_546,N_9845,N_9879);
nor UO_547 (O_547,N_9966,N_9987);
nor UO_548 (O_548,N_9988,N_9831);
nand UO_549 (O_549,N_9954,N_9932);
and UO_550 (O_550,N_9819,N_9959);
nand UO_551 (O_551,N_9982,N_9829);
nor UO_552 (O_552,N_9948,N_9868);
nand UO_553 (O_553,N_9851,N_9910);
nand UO_554 (O_554,N_9852,N_9916);
nand UO_555 (O_555,N_9850,N_9976);
nor UO_556 (O_556,N_9944,N_9989);
or UO_557 (O_557,N_9859,N_9921);
and UO_558 (O_558,N_9858,N_9839);
and UO_559 (O_559,N_9912,N_9852);
and UO_560 (O_560,N_9826,N_9816);
and UO_561 (O_561,N_9897,N_9831);
nand UO_562 (O_562,N_9999,N_9987);
nand UO_563 (O_563,N_9878,N_9929);
nor UO_564 (O_564,N_9964,N_9801);
or UO_565 (O_565,N_9807,N_9813);
or UO_566 (O_566,N_9819,N_9908);
nand UO_567 (O_567,N_9990,N_9957);
nand UO_568 (O_568,N_9901,N_9876);
nor UO_569 (O_569,N_9924,N_9925);
nor UO_570 (O_570,N_9962,N_9804);
nor UO_571 (O_571,N_9914,N_9800);
nand UO_572 (O_572,N_9994,N_9956);
nand UO_573 (O_573,N_9832,N_9811);
or UO_574 (O_574,N_9852,N_9851);
xnor UO_575 (O_575,N_9867,N_9942);
xnor UO_576 (O_576,N_9948,N_9800);
and UO_577 (O_577,N_9900,N_9914);
or UO_578 (O_578,N_9833,N_9890);
and UO_579 (O_579,N_9878,N_9971);
or UO_580 (O_580,N_9839,N_9880);
nor UO_581 (O_581,N_9981,N_9995);
nor UO_582 (O_582,N_9999,N_9892);
nand UO_583 (O_583,N_9858,N_9908);
nor UO_584 (O_584,N_9944,N_9883);
nor UO_585 (O_585,N_9979,N_9937);
nand UO_586 (O_586,N_9977,N_9948);
or UO_587 (O_587,N_9996,N_9807);
and UO_588 (O_588,N_9931,N_9971);
xnor UO_589 (O_589,N_9977,N_9985);
and UO_590 (O_590,N_9829,N_9883);
and UO_591 (O_591,N_9880,N_9868);
and UO_592 (O_592,N_9829,N_9944);
xor UO_593 (O_593,N_9980,N_9855);
nor UO_594 (O_594,N_9800,N_9804);
nor UO_595 (O_595,N_9957,N_9915);
or UO_596 (O_596,N_9818,N_9854);
xor UO_597 (O_597,N_9826,N_9954);
or UO_598 (O_598,N_9943,N_9830);
nor UO_599 (O_599,N_9813,N_9944);
nand UO_600 (O_600,N_9980,N_9886);
nand UO_601 (O_601,N_9878,N_9807);
and UO_602 (O_602,N_9932,N_9859);
nand UO_603 (O_603,N_9829,N_9862);
and UO_604 (O_604,N_9938,N_9811);
nand UO_605 (O_605,N_9850,N_9811);
nand UO_606 (O_606,N_9904,N_9933);
xnor UO_607 (O_607,N_9975,N_9997);
and UO_608 (O_608,N_9894,N_9975);
or UO_609 (O_609,N_9922,N_9970);
or UO_610 (O_610,N_9953,N_9815);
xnor UO_611 (O_611,N_9975,N_9956);
nand UO_612 (O_612,N_9929,N_9933);
nor UO_613 (O_613,N_9843,N_9866);
or UO_614 (O_614,N_9911,N_9916);
or UO_615 (O_615,N_9971,N_9967);
nor UO_616 (O_616,N_9828,N_9869);
or UO_617 (O_617,N_9829,N_9866);
xnor UO_618 (O_618,N_9973,N_9840);
nand UO_619 (O_619,N_9846,N_9893);
or UO_620 (O_620,N_9899,N_9832);
or UO_621 (O_621,N_9947,N_9948);
xor UO_622 (O_622,N_9932,N_9832);
nand UO_623 (O_623,N_9915,N_9853);
or UO_624 (O_624,N_9998,N_9857);
or UO_625 (O_625,N_9936,N_9955);
nor UO_626 (O_626,N_9928,N_9852);
nor UO_627 (O_627,N_9992,N_9917);
nor UO_628 (O_628,N_9868,N_9954);
xnor UO_629 (O_629,N_9946,N_9829);
nand UO_630 (O_630,N_9954,N_9896);
nor UO_631 (O_631,N_9961,N_9867);
nand UO_632 (O_632,N_9958,N_9902);
nor UO_633 (O_633,N_9818,N_9838);
and UO_634 (O_634,N_9971,N_9879);
nand UO_635 (O_635,N_9950,N_9809);
xnor UO_636 (O_636,N_9942,N_9825);
and UO_637 (O_637,N_9865,N_9891);
nand UO_638 (O_638,N_9834,N_9841);
and UO_639 (O_639,N_9988,N_9841);
or UO_640 (O_640,N_9933,N_9871);
nand UO_641 (O_641,N_9909,N_9950);
nor UO_642 (O_642,N_9838,N_9982);
and UO_643 (O_643,N_9965,N_9955);
or UO_644 (O_644,N_9929,N_9979);
or UO_645 (O_645,N_9806,N_9864);
and UO_646 (O_646,N_9923,N_9907);
or UO_647 (O_647,N_9877,N_9897);
or UO_648 (O_648,N_9915,N_9899);
nor UO_649 (O_649,N_9925,N_9835);
xor UO_650 (O_650,N_9816,N_9847);
xor UO_651 (O_651,N_9805,N_9871);
nand UO_652 (O_652,N_9844,N_9994);
and UO_653 (O_653,N_9963,N_9848);
nand UO_654 (O_654,N_9989,N_9880);
nand UO_655 (O_655,N_9913,N_9856);
nand UO_656 (O_656,N_9876,N_9848);
nor UO_657 (O_657,N_9914,N_9899);
nor UO_658 (O_658,N_9804,N_9835);
nor UO_659 (O_659,N_9941,N_9827);
nor UO_660 (O_660,N_9988,N_9943);
nor UO_661 (O_661,N_9978,N_9942);
nand UO_662 (O_662,N_9877,N_9921);
nor UO_663 (O_663,N_9839,N_9873);
or UO_664 (O_664,N_9826,N_9806);
xor UO_665 (O_665,N_9838,N_9831);
nor UO_666 (O_666,N_9896,N_9938);
and UO_667 (O_667,N_9930,N_9946);
and UO_668 (O_668,N_9984,N_9846);
nand UO_669 (O_669,N_9840,N_9951);
or UO_670 (O_670,N_9924,N_9812);
or UO_671 (O_671,N_9950,N_9893);
nand UO_672 (O_672,N_9873,N_9897);
nor UO_673 (O_673,N_9866,N_9803);
nor UO_674 (O_674,N_9884,N_9836);
nand UO_675 (O_675,N_9819,N_9998);
nand UO_676 (O_676,N_9945,N_9819);
and UO_677 (O_677,N_9851,N_9994);
or UO_678 (O_678,N_9872,N_9856);
nand UO_679 (O_679,N_9980,N_9926);
and UO_680 (O_680,N_9948,N_9900);
nand UO_681 (O_681,N_9804,N_9950);
or UO_682 (O_682,N_9997,N_9974);
and UO_683 (O_683,N_9917,N_9889);
and UO_684 (O_684,N_9943,N_9876);
nor UO_685 (O_685,N_9858,N_9848);
nor UO_686 (O_686,N_9929,N_9883);
xnor UO_687 (O_687,N_9915,N_9843);
nor UO_688 (O_688,N_9993,N_9946);
and UO_689 (O_689,N_9827,N_9883);
nand UO_690 (O_690,N_9973,N_9841);
nand UO_691 (O_691,N_9986,N_9829);
nor UO_692 (O_692,N_9901,N_9898);
and UO_693 (O_693,N_9943,N_9824);
and UO_694 (O_694,N_9843,N_9859);
or UO_695 (O_695,N_9989,N_9976);
xnor UO_696 (O_696,N_9835,N_9812);
nor UO_697 (O_697,N_9852,N_9940);
nor UO_698 (O_698,N_9997,N_9938);
nand UO_699 (O_699,N_9850,N_9937);
nor UO_700 (O_700,N_9874,N_9895);
nand UO_701 (O_701,N_9946,N_9911);
or UO_702 (O_702,N_9850,N_9845);
and UO_703 (O_703,N_9854,N_9890);
or UO_704 (O_704,N_9957,N_9987);
and UO_705 (O_705,N_9896,N_9919);
nand UO_706 (O_706,N_9982,N_9868);
or UO_707 (O_707,N_9875,N_9803);
and UO_708 (O_708,N_9850,N_9961);
nand UO_709 (O_709,N_9950,N_9977);
or UO_710 (O_710,N_9966,N_9854);
xnor UO_711 (O_711,N_9873,N_9905);
nand UO_712 (O_712,N_9918,N_9896);
or UO_713 (O_713,N_9968,N_9803);
nand UO_714 (O_714,N_9990,N_9848);
and UO_715 (O_715,N_9905,N_9996);
nand UO_716 (O_716,N_9983,N_9808);
nor UO_717 (O_717,N_9987,N_9831);
nor UO_718 (O_718,N_9954,N_9980);
nor UO_719 (O_719,N_9986,N_9812);
and UO_720 (O_720,N_9924,N_9844);
nor UO_721 (O_721,N_9904,N_9887);
and UO_722 (O_722,N_9996,N_9947);
or UO_723 (O_723,N_9870,N_9963);
or UO_724 (O_724,N_9803,N_9885);
nand UO_725 (O_725,N_9942,N_9856);
or UO_726 (O_726,N_9903,N_9976);
nand UO_727 (O_727,N_9985,N_9910);
nor UO_728 (O_728,N_9915,N_9902);
nor UO_729 (O_729,N_9846,N_9996);
nor UO_730 (O_730,N_9921,N_9943);
or UO_731 (O_731,N_9969,N_9914);
nor UO_732 (O_732,N_9898,N_9851);
nor UO_733 (O_733,N_9850,N_9956);
or UO_734 (O_734,N_9847,N_9965);
nand UO_735 (O_735,N_9947,N_9884);
nand UO_736 (O_736,N_9866,N_9823);
nor UO_737 (O_737,N_9958,N_9971);
and UO_738 (O_738,N_9870,N_9833);
nor UO_739 (O_739,N_9936,N_9880);
nor UO_740 (O_740,N_9891,N_9823);
or UO_741 (O_741,N_9888,N_9957);
and UO_742 (O_742,N_9883,N_9865);
nor UO_743 (O_743,N_9835,N_9856);
and UO_744 (O_744,N_9909,N_9951);
nor UO_745 (O_745,N_9826,N_9898);
nand UO_746 (O_746,N_9826,N_9965);
and UO_747 (O_747,N_9806,N_9912);
nand UO_748 (O_748,N_9888,N_9978);
xor UO_749 (O_749,N_9830,N_9985);
nand UO_750 (O_750,N_9902,N_9957);
nor UO_751 (O_751,N_9811,N_9959);
nor UO_752 (O_752,N_9805,N_9896);
and UO_753 (O_753,N_9826,N_9875);
or UO_754 (O_754,N_9874,N_9844);
and UO_755 (O_755,N_9899,N_9958);
nand UO_756 (O_756,N_9808,N_9819);
or UO_757 (O_757,N_9915,N_9819);
or UO_758 (O_758,N_9808,N_9855);
nand UO_759 (O_759,N_9801,N_9906);
or UO_760 (O_760,N_9863,N_9911);
or UO_761 (O_761,N_9976,N_9821);
or UO_762 (O_762,N_9894,N_9918);
and UO_763 (O_763,N_9898,N_9937);
nor UO_764 (O_764,N_9804,N_9940);
and UO_765 (O_765,N_9817,N_9958);
xor UO_766 (O_766,N_9910,N_9937);
nand UO_767 (O_767,N_9822,N_9819);
and UO_768 (O_768,N_9869,N_9954);
nor UO_769 (O_769,N_9838,N_9859);
nand UO_770 (O_770,N_9805,N_9850);
or UO_771 (O_771,N_9905,N_9900);
nand UO_772 (O_772,N_9816,N_9806);
nand UO_773 (O_773,N_9990,N_9810);
nor UO_774 (O_774,N_9868,N_9915);
nand UO_775 (O_775,N_9982,N_9824);
nor UO_776 (O_776,N_9853,N_9820);
or UO_777 (O_777,N_9977,N_9875);
nor UO_778 (O_778,N_9861,N_9848);
nor UO_779 (O_779,N_9994,N_9968);
or UO_780 (O_780,N_9986,N_9895);
and UO_781 (O_781,N_9809,N_9870);
or UO_782 (O_782,N_9914,N_9980);
and UO_783 (O_783,N_9836,N_9969);
or UO_784 (O_784,N_9996,N_9987);
nand UO_785 (O_785,N_9961,N_9960);
and UO_786 (O_786,N_9859,N_9947);
or UO_787 (O_787,N_9986,N_9904);
and UO_788 (O_788,N_9915,N_9921);
and UO_789 (O_789,N_9844,N_9882);
nand UO_790 (O_790,N_9860,N_9925);
or UO_791 (O_791,N_9880,N_9984);
nand UO_792 (O_792,N_9837,N_9869);
nor UO_793 (O_793,N_9824,N_9940);
and UO_794 (O_794,N_9819,N_9928);
nand UO_795 (O_795,N_9940,N_9946);
nor UO_796 (O_796,N_9829,N_9998);
nor UO_797 (O_797,N_9889,N_9916);
nor UO_798 (O_798,N_9880,N_9899);
and UO_799 (O_799,N_9975,N_9820);
xnor UO_800 (O_800,N_9917,N_9905);
or UO_801 (O_801,N_9832,N_9922);
and UO_802 (O_802,N_9930,N_9920);
nand UO_803 (O_803,N_9988,N_9990);
or UO_804 (O_804,N_9822,N_9940);
or UO_805 (O_805,N_9940,N_9976);
nand UO_806 (O_806,N_9826,N_9910);
and UO_807 (O_807,N_9889,N_9835);
nor UO_808 (O_808,N_9935,N_9836);
nor UO_809 (O_809,N_9928,N_9965);
or UO_810 (O_810,N_9909,N_9993);
nor UO_811 (O_811,N_9823,N_9919);
and UO_812 (O_812,N_9897,N_9946);
nor UO_813 (O_813,N_9893,N_9955);
nor UO_814 (O_814,N_9897,N_9871);
or UO_815 (O_815,N_9858,N_9928);
or UO_816 (O_816,N_9974,N_9920);
or UO_817 (O_817,N_9993,N_9959);
or UO_818 (O_818,N_9862,N_9898);
and UO_819 (O_819,N_9821,N_9833);
and UO_820 (O_820,N_9999,N_9986);
nor UO_821 (O_821,N_9977,N_9804);
and UO_822 (O_822,N_9957,N_9976);
or UO_823 (O_823,N_9816,N_9924);
nand UO_824 (O_824,N_9978,N_9823);
nand UO_825 (O_825,N_9936,N_9976);
nand UO_826 (O_826,N_9962,N_9858);
and UO_827 (O_827,N_9953,N_9999);
nand UO_828 (O_828,N_9816,N_9840);
or UO_829 (O_829,N_9906,N_9847);
and UO_830 (O_830,N_9843,N_9801);
nor UO_831 (O_831,N_9826,N_9973);
or UO_832 (O_832,N_9896,N_9904);
nor UO_833 (O_833,N_9959,N_9906);
or UO_834 (O_834,N_9915,N_9983);
or UO_835 (O_835,N_9916,N_9827);
nand UO_836 (O_836,N_9975,N_9835);
or UO_837 (O_837,N_9882,N_9849);
or UO_838 (O_838,N_9923,N_9847);
nor UO_839 (O_839,N_9926,N_9987);
xor UO_840 (O_840,N_9892,N_9904);
and UO_841 (O_841,N_9955,N_9967);
and UO_842 (O_842,N_9844,N_9986);
nor UO_843 (O_843,N_9804,N_9865);
nand UO_844 (O_844,N_9994,N_9998);
nand UO_845 (O_845,N_9945,N_9908);
xnor UO_846 (O_846,N_9948,N_9839);
xor UO_847 (O_847,N_9915,N_9825);
nor UO_848 (O_848,N_9816,N_9891);
or UO_849 (O_849,N_9948,N_9862);
or UO_850 (O_850,N_9947,N_9923);
or UO_851 (O_851,N_9867,N_9812);
nand UO_852 (O_852,N_9839,N_9872);
or UO_853 (O_853,N_9820,N_9937);
and UO_854 (O_854,N_9838,N_9801);
or UO_855 (O_855,N_9814,N_9840);
xnor UO_856 (O_856,N_9997,N_9810);
nand UO_857 (O_857,N_9864,N_9819);
nand UO_858 (O_858,N_9982,N_9917);
nand UO_859 (O_859,N_9839,N_9994);
nand UO_860 (O_860,N_9928,N_9832);
and UO_861 (O_861,N_9944,N_9984);
or UO_862 (O_862,N_9940,N_9975);
xor UO_863 (O_863,N_9822,N_9942);
or UO_864 (O_864,N_9845,N_9811);
or UO_865 (O_865,N_9868,N_9974);
or UO_866 (O_866,N_9908,N_9911);
or UO_867 (O_867,N_9901,N_9815);
and UO_868 (O_868,N_9947,N_9818);
or UO_869 (O_869,N_9974,N_9941);
or UO_870 (O_870,N_9816,N_9872);
or UO_871 (O_871,N_9881,N_9888);
or UO_872 (O_872,N_9845,N_9968);
and UO_873 (O_873,N_9845,N_9801);
nor UO_874 (O_874,N_9890,N_9939);
nand UO_875 (O_875,N_9826,N_9867);
xnor UO_876 (O_876,N_9930,N_9833);
or UO_877 (O_877,N_9958,N_9937);
or UO_878 (O_878,N_9950,N_9838);
nand UO_879 (O_879,N_9885,N_9904);
xnor UO_880 (O_880,N_9859,N_9919);
nand UO_881 (O_881,N_9854,N_9895);
nor UO_882 (O_882,N_9984,N_9997);
or UO_883 (O_883,N_9913,N_9807);
and UO_884 (O_884,N_9893,N_9827);
nor UO_885 (O_885,N_9939,N_9800);
nand UO_886 (O_886,N_9930,N_9881);
or UO_887 (O_887,N_9885,N_9965);
nand UO_888 (O_888,N_9993,N_9949);
or UO_889 (O_889,N_9933,N_9993);
nand UO_890 (O_890,N_9841,N_9968);
and UO_891 (O_891,N_9916,N_9860);
and UO_892 (O_892,N_9817,N_9998);
nand UO_893 (O_893,N_9905,N_9865);
or UO_894 (O_894,N_9995,N_9803);
and UO_895 (O_895,N_9804,N_9973);
nor UO_896 (O_896,N_9981,N_9974);
or UO_897 (O_897,N_9813,N_9902);
or UO_898 (O_898,N_9886,N_9957);
or UO_899 (O_899,N_9997,N_9844);
or UO_900 (O_900,N_9856,N_9808);
nand UO_901 (O_901,N_9999,N_9903);
or UO_902 (O_902,N_9959,N_9824);
and UO_903 (O_903,N_9899,N_9801);
nand UO_904 (O_904,N_9850,N_9898);
nor UO_905 (O_905,N_9959,N_9930);
nand UO_906 (O_906,N_9966,N_9889);
nor UO_907 (O_907,N_9914,N_9869);
or UO_908 (O_908,N_9888,N_9940);
or UO_909 (O_909,N_9877,N_9882);
or UO_910 (O_910,N_9911,N_9977);
nand UO_911 (O_911,N_9809,N_9974);
or UO_912 (O_912,N_9867,N_9903);
nand UO_913 (O_913,N_9897,N_9851);
and UO_914 (O_914,N_9853,N_9800);
or UO_915 (O_915,N_9940,N_9929);
nor UO_916 (O_916,N_9839,N_9990);
nor UO_917 (O_917,N_9988,N_9847);
and UO_918 (O_918,N_9939,N_9805);
or UO_919 (O_919,N_9886,N_9812);
nand UO_920 (O_920,N_9809,N_9947);
nor UO_921 (O_921,N_9991,N_9891);
nor UO_922 (O_922,N_9851,N_9939);
nor UO_923 (O_923,N_9937,N_9884);
nor UO_924 (O_924,N_9879,N_9972);
xor UO_925 (O_925,N_9806,N_9827);
nor UO_926 (O_926,N_9914,N_9942);
and UO_927 (O_927,N_9887,N_9817);
nor UO_928 (O_928,N_9828,N_9992);
nand UO_929 (O_929,N_9812,N_9948);
and UO_930 (O_930,N_9928,N_9931);
nor UO_931 (O_931,N_9821,N_9875);
or UO_932 (O_932,N_9895,N_9816);
or UO_933 (O_933,N_9968,N_9832);
xnor UO_934 (O_934,N_9830,N_9958);
xor UO_935 (O_935,N_9889,N_9837);
or UO_936 (O_936,N_9966,N_9807);
and UO_937 (O_937,N_9982,N_9800);
and UO_938 (O_938,N_9819,N_9838);
or UO_939 (O_939,N_9819,N_9974);
xnor UO_940 (O_940,N_9956,N_9908);
or UO_941 (O_941,N_9946,N_9906);
nor UO_942 (O_942,N_9872,N_9905);
xor UO_943 (O_943,N_9947,N_9978);
and UO_944 (O_944,N_9825,N_9985);
and UO_945 (O_945,N_9915,N_9834);
nand UO_946 (O_946,N_9915,N_9916);
and UO_947 (O_947,N_9965,N_9933);
or UO_948 (O_948,N_9853,N_9862);
nor UO_949 (O_949,N_9887,N_9874);
or UO_950 (O_950,N_9991,N_9864);
nor UO_951 (O_951,N_9912,N_9903);
nand UO_952 (O_952,N_9992,N_9812);
or UO_953 (O_953,N_9906,N_9971);
or UO_954 (O_954,N_9988,N_9845);
nor UO_955 (O_955,N_9958,N_9951);
and UO_956 (O_956,N_9890,N_9924);
nand UO_957 (O_957,N_9865,N_9801);
or UO_958 (O_958,N_9863,N_9901);
nor UO_959 (O_959,N_9867,N_9923);
or UO_960 (O_960,N_9851,N_9923);
and UO_961 (O_961,N_9827,N_9959);
and UO_962 (O_962,N_9898,N_9993);
or UO_963 (O_963,N_9881,N_9948);
or UO_964 (O_964,N_9854,N_9865);
nand UO_965 (O_965,N_9824,N_9878);
nand UO_966 (O_966,N_9860,N_9935);
or UO_967 (O_967,N_9830,N_9866);
xnor UO_968 (O_968,N_9800,N_9814);
nand UO_969 (O_969,N_9952,N_9840);
nand UO_970 (O_970,N_9844,N_9839);
or UO_971 (O_971,N_9985,N_9975);
nand UO_972 (O_972,N_9988,N_9986);
or UO_973 (O_973,N_9846,N_9804);
or UO_974 (O_974,N_9920,N_9918);
nor UO_975 (O_975,N_9815,N_9995);
and UO_976 (O_976,N_9922,N_9811);
and UO_977 (O_977,N_9901,N_9998);
nand UO_978 (O_978,N_9996,N_9967);
and UO_979 (O_979,N_9856,N_9824);
or UO_980 (O_980,N_9934,N_9856);
nor UO_981 (O_981,N_9851,N_9966);
and UO_982 (O_982,N_9808,N_9893);
or UO_983 (O_983,N_9938,N_9810);
or UO_984 (O_984,N_9981,N_9911);
and UO_985 (O_985,N_9990,N_9884);
nand UO_986 (O_986,N_9877,N_9806);
nor UO_987 (O_987,N_9812,N_9841);
nor UO_988 (O_988,N_9990,N_9991);
nor UO_989 (O_989,N_9979,N_9833);
nor UO_990 (O_990,N_9962,N_9899);
or UO_991 (O_991,N_9914,N_9807);
and UO_992 (O_992,N_9958,N_9845);
and UO_993 (O_993,N_9947,N_9939);
nand UO_994 (O_994,N_9839,N_9973);
nand UO_995 (O_995,N_9983,N_9975);
and UO_996 (O_996,N_9813,N_9851);
nand UO_997 (O_997,N_9967,N_9974);
nand UO_998 (O_998,N_9917,N_9864);
and UO_999 (O_999,N_9907,N_9993);
and UO_1000 (O_1000,N_9885,N_9934);
or UO_1001 (O_1001,N_9974,N_9973);
nand UO_1002 (O_1002,N_9800,N_9871);
and UO_1003 (O_1003,N_9981,N_9876);
and UO_1004 (O_1004,N_9876,N_9880);
nand UO_1005 (O_1005,N_9974,N_9990);
or UO_1006 (O_1006,N_9963,N_9900);
nand UO_1007 (O_1007,N_9843,N_9807);
and UO_1008 (O_1008,N_9915,N_9946);
nor UO_1009 (O_1009,N_9894,N_9973);
nand UO_1010 (O_1010,N_9963,N_9927);
and UO_1011 (O_1011,N_9888,N_9954);
and UO_1012 (O_1012,N_9851,N_9906);
nand UO_1013 (O_1013,N_9822,N_9835);
and UO_1014 (O_1014,N_9998,N_9916);
or UO_1015 (O_1015,N_9836,N_9941);
nand UO_1016 (O_1016,N_9974,N_9980);
nand UO_1017 (O_1017,N_9937,N_9976);
and UO_1018 (O_1018,N_9912,N_9976);
nand UO_1019 (O_1019,N_9914,N_9961);
nor UO_1020 (O_1020,N_9958,N_9972);
nor UO_1021 (O_1021,N_9957,N_9861);
and UO_1022 (O_1022,N_9930,N_9961);
or UO_1023 (O_1023,N_9939,N_9968);
nor UO_1024 (O_1024,N_9988,N_9836);
nand UO_1025 (O_1025,N_9833,N_9907);
nand UO_1026 (O_1026,N_9910,N_9911);
xor UO_1027 (O_1027,N_9973,N_9986);
xor UO_1028 (O_1028,N_9936,N_9914);
and UO_1029 (O_1029,N_9967,N_9821);
or UO_1030 (O_1030,N_9863,N_9872);
and UO_1031 (O_1031,N_9940,N_9910);
and UO_1032 (O_1032,N_9816,N_9810);
and UO_1033 (O_1033,N_9910,N_9885);
nor UO_1034 (O_1034,N_9942,N_9926);
and UO_1035 (O_1035,N_9885,N_9848);
or UO_1036 (O_1036,N_9949,N_9862);
nor UO_1037 (O_1037,N_9886,N_9838);
and UO_1038 (O_1038,N_9914,N_9975);
nand UO_1039 (O_1039,N_9848,N_9921);
nand UO_1040 (O_1040,N_9818,N_9994);
nand UO_1041 (O_1041,N_9802,N_9844);
and UO_1042 (O_1042,N_9897,N_9952);
and UO_1043 (O_1043,N_9815,N_9905);
or UO_1044 (O_1044,N_9985,N_9852);
xor UO_1045 (O_1045,N_9803,N_9996);
nor UO_1046 (O_1046,N_9812,N_9915);
or UO_1047 (O_1047,N_9885,N_9831);
nor UO_1048 (O_1048,N_9829,N_9856);
and UO_1049 (O_1049,N_9971,N_9920);
and UO_1050 (O_1050,N_9861,N_9845);
or UO_1051 (O_1051,N_9845,N_9840);
nand UO_1052 (O_1052,N_9992,N_9951);
nor UO_1053 (O_1053,N_9813,N_9907);
nor UO_1054 (O_1054,N_9976,N_9891);
or UO_1055 (O_1055,N_9858,N_9947);
nand UO_1056 (O_1056,N_9843,N_9857);
and UO_1057 (O_1057,N_9813,N_9884);
nand UO_1058 (O_1058,N_9812,N_9958);
nor UO_1059 (O_1059,N_9991,N_9899);
and UO_1060 (O_1060,N_9933,N_9991);
or UO_1061 (O_1061,N_9936,N_9893);
nor UO_1062 (O_1062,N_9939,N_9893);
nor UO_1063 (O_1063,N_9804,N_9819);
nor UO_1064 (O_1064,N_9809,N_9992);
and UO_1065 (O_1065,N_9861,N_9931);
and UO_1066 (O_1066,N_9837,N_9888);
and UO_1067 (O_1067,N_9869,N_9805);
xor UO_1068 (O_1068,N_9968,N_9812);
or UO_1069 (O_1069,N_9989,N_9846);
and UO_1070 (O_1070,N_9869,N_9826);
and UO_1071 (O_1071,N_9882,N_9857);
nand UO_1072 (O_1072,N_9856,N_9848);
nand UO_1073 (O_1073,N_9951,N_9859);
xor UO_1074 (O_1074,N_9986,N_9821);
or UO_1075 (O_1075,N_9936,N_9984);
or UO_1076 (O_1076,N_9802,N_9849);
nand UO_1077 (O_1077,N_9822,N_9906);
xor UO_1078 (O_1078,N_9868,N_9996);
nor UO_1079 (O_1079,N_9979,N_9866);
nor UO_1080 (O_1080,N_9920,N_9895);
nor UO_1081 (O_1081,N_9894,N_9804);
nor UO_1082 (O_1082,N_9863,N_9861);
nand UO_1083 (O_1083,N_9895,N_9961);
nand UO_1084 (O_1084,N_9945,N_9884);
and UO_1085 (O_1085,N_9936,N_9863);
nand UO_1086 (O_1086,N_9919,N_9931);
nor UO_1087 (O_1087,N_9994,N_9904);
nor UO_1088 (O_1088,N_9912,N_9923);
xor UO_1089 (O_1089,N_9827,N_9831);
or UO_1090 (O_1090,N_9889,N_9964);
or UO_1091 (O_1091,N_9996,N_9994);
nor UO_1092 (O_1092,N_9911,N_9924);
and UO_1093 (O_1093,N_9955,N_9863);
or UO_1094 (O_1094,N_9872,N_9967);
nand UO_1095 (O_1095,N_9912,N_9938);
or UO_1096 (O_1096,N_9957,N_9905);
nor UO_1097 (O_1097,N_9825,N_9817);
nand UO_1098 (O_1098,N_9921,N_9927);
nor UO_1099 (O_1099,N_9890,N_9904);
and UO_1100 (O_1100,N_9819,N_9809);
and UO_1101 (O_1101,N_9905,N_9809);
xnor UO_1102 (O_1102,N_9814,N_9856);
nor UO_1103 (O_1103,N_9931,N_9836);
nor UO_1104 (O_1104,N_9880,N_9981);
and UO_1105 (O_1105,N_9872,N_9871);
or UO_1106 (O_1106,N_9991,N_9977);
xnor UO_1107 (O_1107,N_9924,N_9818);
and UO_1108 (O_1108,N_9945,N_9885);
and UO_1109 (O_1109,N_9906,N_9824);
nor UO_1110 (O_1110,N_9814,N_9926);
nor UO_1111 (O_1111,N_9919,N_9862);
nand UO_1112 (O_1112,N_9927,N_9826);
and UO_1113 (O_1113,N_9964,N_9879);
nand UO_1114 (O_1114,N_9983,N_9925);
and UO_1115 (O_1115,N_9839,N_9867);
or UO_1116 (O_1116,N_9944,N_9848);
and UO_1117 (O_1117,N_9850,N_9934);
nor UO_1118 (O_1118,N_9918,N_9835);
or UO_1119 (O_1119,N_9910,N_9939);
nand UO_1120 (O_1120,N_9941,N_9816);
or UO_1121 (O_1121,N_9867,N_9998);
nor UO_1122 (O_1122,N_9979,N_9830);
and UO_1123 (O_1123,N_9854,N_9919);
and UO_1124 (O_1124,N_9919,N_9952);
nor UO_1125 (O_1125,N_9990,N_9921);
and UO_1126 (O_1126,N_9918,N_9941);
nand UO_1127 (O_1127,N_9843,N_9999);
nand UO_1128 (O_1128,N_9950,N_9981);
or UO_1129 (O_1129,N_9906,N_9894);
xnor UO_1130 (O_1130,N_9904,N_9822);
or UO_1131 (O_1131,N_9972,N_9979);
or UO_1132 (O_1132,N_9885,N_9816);
and UO_1133 (O_1133,N_9830,N_9983);
and UO_1134 (O_1134,N_9953,N_9983);
and UO_1135 (O_1135,N_9815,N_9944);
nor UO_1136 (O_1136,N_9896,N_9845);
or UO_1137 (O_1137,N_9919,N_9847);
and UO_1138 (O_1138,N_9820,N_9842);
and UO_1139 (O_1139,N_9986,N_9956);
nor UO_1140 (O_1140,N_9924,N_9854);
or UO_1141 (O_1141,N_9870,N_9920);
and UO_1142 (O_1142,N_9999,N_9801);
or UO_1143 (O_1143,N_9974,N_9838);
and UO_1144 (O_1144,N_9838,N_9961);
nor UO_1145 (O_1145,N_9824,N_9800);
or UO_1146 (O_1146,N_9805,N_9944);
and UO_1147 (O_1147,N_9984,N_9948);
nand UO_1148 (O_1148,N_9837,N_9910);
nand UO_1149 (O_1149,N_9860,N_9900);
and UO_1150 (O_1150,N_9903,N_9990);
nor UO_1151 (O_1151,N_9864,N_9809);
nand UO_1152 (O_1152,N_9820,N_9996);
xnor UO_1153 (O_1153,N_9852,N_9867);
or UO_1154 (O_1154,N_9825,N_9874);
nand UO_1155 (O_1155,N_9921,N_9907);
nand UO_1156 (O_1156,N_9858,N_9817);
and UO_1157 (O_1157,N_9981,N_9877);
or UO_1158 (O_1158,N_9828,N_9933);
and UO_1159 (O_1159,N_9990,N_9868);
or UO_1160 (O_1160,N_9820,N_9931);
and UO_1161 (O_1161,N_9825,N_9979);
and UO_1162 (O_1162,N_9822,N_9817);
nand UO_1163 (O_1163,N_9868,N_9825);
and UO_1164 (O_1164,N_9986,N_9860);
nand UO_1165 (O_1165,N_9989,N_9827);
nor UO_1166 (O_1166,N_9846,N_9994);
nor UO_1167 (O_1167,N_9860,N_9866);
and UO_1168 (O_1168,N_9815,N_9970);
and UO_1169 (O_1169,N_9823,N_9809);
nand UO_1170 (O_1170,N_9936,N_9803);
nand UO_1171 (O_1171,N_9835,N_9947);
nor UO_1172 (O_1172,N_9998,N_9954);
nor UO_1173 (O_1173,N_9976,N_9947);
nand UO_1174 (O_1174,N_9877,N_9870);
or UO_1175 (O_1175,N_9823,N_9837);
xor UO_1176 (O_1176,N_9844,N_9957);
nand UO_1177 (O_1177,N_9983,N_9999);
and UO_1178 (O_1178,N_9932,N_9934);
nor UO_1179 (O_1179,N_9822,N_9900);
nand UO_1180 (O_1180,N_9822,N_9874);
nor UO_1181 (O_1181,N_9952,N_9962);
and UO_1182 (O_1182,N_9926,N_9847);
nand UO_1183 (O_1183,N_9970,N_9953);
xnor UO_1184 (O_1184,N_9810,N_9987);
nand UO_1185 (O_1185,N_9831,N_9940);
nor UO_1186 (O_1186,N_9809,N_9982);
and UO_1187 (O_1187,N_9912,N_9951);
nand UO_1188 (O_1188,N_9823,N_9968);
or UO_1189 (O_1189,N_9896,N_9800);
and UO_1190 (O_1190,N_9873,N_9958);
nand UO_1191 (O_1191,N_9916,N_9867);
nor UO_1192 (O_1192,N_9979,N_9809);
and UO_1193 (O_1193,N_9939,N_9902);
nor UO_1194 (O_1194,N_9832,N_9892);
and UO_1195 (O_1195,N_9981,N_9943);
nor UO_1196 (O_1196,N_9914,N_9885);
and UO_1197 (O_1197,N_9955,N_9890);
or UO_1198 (O_1198,N_9885,N_9829);
nand UO_1199 (O_1199,N_9985,N_9894);
nor UO_1200 (O_1200,N_9869,N_9862);
and UO_1201 (O_1201,N_9948,N_9893);
nand UO_1202 (O_1202,N_9927,N_9848);
nor UO_1203 (O_1203,N_9975,N_9935);
nor UO_1204 (O_1204,N_9880,N_9812);
or UO_1205 (O_1205,N_9801,N_9872);
and UO_1206 (O_1206,N_9870,N_9932);
nor UO_1207 (O_1207,N_9864,N_9951);
and UO_1208 (O_1208,N_9820,N_9912);
nor UO_1209 (O_1209,N_9905,N_9801);
nand UO_1210 (O_1210,N_9888,N_9859);
nand UO_1211 (O_1211,N_9916,N_9977);
xor UO_1212 (O_1212,N_9912,N_9880);
nor UO_1213 (O_1213,N_9980,N_9870);
xnor UO_1214 (O_1214,N_9934,N_9875);
or UO_1215 (O_1215,N_9814,N_9880);
and UO_1216 (O_1216,N_9967,N_9977);
nor UO_1217 (O_1217,N_9918,N_9891);
nor UO_1218 (O_1218,N_9837,N_9849);
nand UO_1219 (O_1219,N_9946,N_9837);
xnor UO_1220 (O_1220,N_9953,N_9928);
or UO_1221 (O_1221,N_9828,N_9945);
xnor UO_1222 (O_1222,N_9878,N_9902);
nand UO_1223 (O_1223,N_9908,N_9893);
and UO_1224 (O_1224,N_9986,N_9816);
xnor UO_1225 (O_1225,N_9914,N_9919);
and UO_1226 (O_1226,N_9913,N_9961);
and UO_1227 (O_1227,N_9929,N_9957);
xnor UO_1228 (O_1228,N_9949,N_9883);
xnor UO_1229 (O_1229,N_9909,N_9892);
xor UO_1230 (O_1230,N_9958,N_9838);
xnor UO_1231 (O_1231,N_9920,N_9995);
or UO_1232 (O_1232,N_9874,N_9906);
nor UO_1233 (O_1233,N_9902,N_9929);
xnor UO_1234 (O_1234,N_9873,N_9843);
and UO_1235 (O_1235,N_9877,N_9841);
xor UO_1236 (O_1236,N_9860,N_9895);
or UO_1237 (O_1237,N_9901,N_9996);
nor UO_1238 (O_1238,N_9904,N_9824);
nor UO_1239 (O_1239,N_9974,N_9987);
nand UO_1240 (O_1240,N_9800,N_9822);
nand UO_1241 (O_1241,N_9881,N_9961);
nand UO_1242 (O_1242,N_9950,N_9801);
and UO_1243 (O_1243,N_9865,N_9908);
or UO_1244 (O_1244,N_9873,N_9877);
or UO_1245 (O_1245,N_9840,N_9864);
nor UO_1246 (O_1246,N_9998,N_9987);
nor UO_1247 (O_1247,N_9817,N_9901);
nor UO_1248 (O_1248,N_9976,N_9851);
and UO_1249 (O_1249,N_9924,N_9961);
and UO_1250 (O_1250,N_9800,N_9846);
and UO_1251 (O_1251,N_9952,N_9859);
or UO_1252 (O_1252,N_9819,N_9982);
and UO_1253 (O_1253,N_9935,N_9902);
xor UO_1254 (O_1254,N_9921,N_9819);
nor UO_1255 (O_1255,N_9833,N_9816);
nand UO_1256 (O_1256,N_9985,N_9984);
nand UO_1257 (O_1257,N_9972,N_9863);
or UO_1258 (O_1258,N_9842,N_9841);
nor UO_1259 (O_1259,N_9933,N_9834);
nand UO_1260 (O_1260,N_9978,N_9938);
nor UO_1261 (O_1261,N_9925,N_9837);
and UO_1262 (O_1262,N_9936,N_9964);
and UO_1263 (O_1263,N_9940,N_9957);
or UO_1264 (O_1264,N_9976,N_9888);
nor UO_1265 (O_1265,N_9870,N_9801);
nor UO_1266 (O_1266,N_9851,N_9981);
nand UO_1267 (O_1267,N_9912,N_9810);
or UO_1268 (O_1268,N_9842,N_9918);
and UO_1269 (O_1269,N_9851,N_9937);
nor UO_1270 (O_1270,N_9821,N_9882);
nor UO_1271 (O_1271,N_9837,N_9838);
and UO_1272 (O_1272,N_9943,N_9805);
and UO_1273 (O_1273,N_9966,N_9820);
and UO_1274 (O_1274,N_9933,N_9928);
or UO_1275 (O_1275,N_9821,N_9939);
or UO_1276 (O_1276,N_9867,N_9888);
nand UO_1277 (O_1277,N_9951,N_9803);
nor UO_1278 (O_1278,N_9897,N_9804);
nand UO_1279 (O_1279,N_9915,N_9960);
xor UO_1280 (O_1280,N_9808,N_9982);
and UO_1281 (O_1281,N_9875,N_9872);
nand UO_1282 (O_1282,N_9983,N_9821);
nand UO_1283 (O_1283,N_9819,N_9961);
nand UO_1284 (O_1284,N_9961,N_9912);
nor UO_1285 (O_1285,N_9904,N_9889);
nor UO_1286 (O_1286,N_9961,N_9824);
nor UO_1287 (O_1287,N_9844,N_9834);
or UO_1288 (O_1288,N_9818,N_9954);
or UO_1289 (O_1289,N_9818,N_9830);
nor UO_1290 (O_1290,N_9940,N_9802);
and UO_1291 (O_1291,N_9849,N_9848);
nand UO_1292 (O_1292,N_9819,N_9906);
and UO_1293 (O_1293,N_9817,N_9947);
nor UO_1294 (O_1294,N_9950,N_9836);
or UO_1295 (O_1295,N_9956,N_9987);
nand UO_1296 (O_1296,N_9975,N_9928);
nand UO_1297 (O_1297,N_9955,N_9911);
or UO_1298 (O_1298,N_9924,N_9823);
and UO_1299 (O_1299,N_9883,N_9942);
nand UO_1300 (O_1300,N_9852,N_9843);
nand UO_1301 (O_1301,N_9848,N_9838);
and UO_1302 (O_1302,N_9978,N_9977);
or UO_1303 (O_1303,N_9986,N_9879);
or UO_1304 (O_1304,N_9973,N_9935);
xnor UO_1305 (O_1305,N_9885,N_9928);
nor UO_1306 (O_1306,N_9894,N_9855);
xor UO_1307 (O_1307,N_9960,N_9868);
and UO_1308 (O_1308,N_9856,N_9827);
xor UO_1309 (O_1309,N_9833,N_9943);
and UO_1310 (O_1310,N_9909,N_9831);
and UO_1311 (O_1311,N_9929,N_9894);
or UO_1312 (O_1312,N_9846,N_9990);
nand UO_1313 (O_1313,N_9832,N_9824);
nand UO_1314 (O_1314,N_9970,N_9872);
nor UO_1315 (O_1315,N_9992,N_9956);
and UO_1316 (O_1316,N_9871,N_9943);
nor UO_1317 (O_1317,N_9866,N_9952);
or UO_1318 (O_1318,N_9873,N_9923);
xor UO_1319 (O_1319,N_9826,N_9818);
or UO_1320 (O_1320,N_9912,N_9908);
xnor UO_1321 (O_1321,N_9955,N_9878);
nand UO_1322 (O_1322,N_9902,N_9995);
xnor UO_1323 (O_1323,N_9961,N_9966);
nor UO_1324 (O_1324,N_9842,N_9967);
nor UO_1325 (O_1325,N_9860,N_9832);
nor UO_1326 (O_1326,N_9837,N_9915);
nor UO_1327 (O_1327,N_9807,N_9918);
and UO_1328 (O_1328,N_9805,N_9843);
nand UO_1329 (O_1329,N_9839,N_9831);
nand UO_1330 (O_1330,N_9830,N_9876);
nand UO_1331 (O_1331,N_9809,N_9993);
nand UO_1332 (O_1332,N_9926,N_9985);
nor UO_1333 (O_1333,N_9809,N_9946);
or UO_1334 (O_1334,N_9881,N_9917);
nand UO_1335 (O_1335,N_9951,N_9807);
xnor UO_1336 (O_1336,N_9961,N_9812);
and UO_1337 (O_1337,N_9926,N_9849);
nand UO_1338 (O_1338,N_9983,N_9887);
and UO_1339 (O_1339,N_9834,N_9875);
and UO_1340 (O_1340,N_9992,N_9869);
nor UO_1341 (O_1341,N_9909,N_9834);
and UO_1342 (O_1342,N_9835,N_9828);
nor UO_1343 (O_1343,N_9958,N_9826);
xnor UO_1344 (O_1344,N_9825,N_9990);
and UO_1345 (O_1345,N_9819,N_9966);
and UO_1346 (O_1346,N_9808,N_9884);
nand UO_1347 (O_1347,N_9921,N_9999);
or UO_1348 (O_1348,N_9873,N_9808);
and UO_1349 (O_1349,N_9969,N_9891);
nand UO_1350 (O_1350,N_9876,N_9842);
xnor UO_1351 (O_1351,N_9853,N_9877);
nor UO_1352 (O_1352,N_9837,N_9880);
or UO_1353 (O_1353,N_9865,N_9921);
or UO_1354 (O_1354,N_9979,N_9967);
or UO_1355 (O_1355,N_9862,N_9994);
and UO_1356 (O_1356,N_9880,N_9924);
or UO_1357 (O_1357,N_9942,N_9985);
or UO_1358 (O_1358,N_9816,N_9851);
xor UO_1359 (O_1359,N_9922,N_9816);
or UO_1360 (O_1360,N_9850,N_9864);
nor UO_1361 (O_1361,N_9840,N_9910);
nand UO_1362 (O_1362,N_9844,N_9825);
or UO_1363 (O_1363,N_9902,N_9816);
and UO_1364 (O_1364,N_9969,N_9964);
and UO_1365 (O_1365,N_9856,N_9810);
or UO_1366 (O_1366,N_9810,N_9928);
nor UO_1367 (O_1367,N_9810,N_9847);
nand UO_1368 (O_1368,N_9996,N_9854);
nor UO_1369 (O_1369,N_9998,N_9996);
nand UO_1370 (O_1370,N_9816,N_9888);
nor UO_1371 (O_1371,N_9870,N_9893);
and UO_1372 (O_1372,N_9914,N_9864);
xnor UO_1373 (O_1373,N_9985,N_9868);
and UO_1374 (O_1374,N_9817,N_9834);
nor UO_1375 (O_1375,N_9861,N_9800);
nand UO_1376 (O_1376,N_9908,N_9954);
nor UO_1377 (O_1377,N_9908,N_9910);
and UO_1378 (O_1378,N_9995,N_9911);
or UO_1379 (O_1379,N_9987,N_9877);
nor UO_1380 (O_1380,N_9807,N_9960);
nand UO_1381 (O_1381,N_9815,N_9917);
nand UO_1382 (O_1382,N_9840,N_9995);
and UO_1383 (O_1383,N_9992,N_9806);
nand UO_1384 (O_1384,N_9826,N_9830);
nand UO_1385 (O_1385,N_9870,N_9816);
xnor UO_1386 (O_1386,N_9966,N_9936);
nor UO_1387 (O_1387,N_9876,N_9939);
and UO_1388 (O_1388,N_9982,N_9882);
or UO_1389 (O_1389,N_9815,N_9833);
or UO_1390 (O_1390,N_9901,N_9803);
or UO_1391 (O_1391,N_9969,N_9972);
or UO_1392 (O_1392,N_9890,N_9808);
nand UO_1393 (O_1393,N_9990,N_9930);
and UO_1394 (O_1394,N_9817,N_9862);
and UO_1395 (O_1395,N_9979,N_9839);
and UO_1396 (O_1396,N_9870,N_9983);
nand UO_1397 (O_1397,N_9824,N_9908);
nand UO_1398 (O_1398,N_9878,N_9869);
nand UO_1399 (O_1399,N_9872,N_9853);
or UO_1400 (O_1400,N_9896,N_9830);
nand UO_1401 (O_1401,N_9916,N_9891);
or UO_1402 (O_1402,N_9958,N_9931);
and UO_1403 (O_1403,N_9950,N_9843);
and UO_1404 (O_1404,N_9837,N_9947);
nand UO_1405 (O_1405,N_9999,N_9992);
nor UO_1406 (O_1406,N_9866,N_9837);
nor UO_1407 (O_1407,N_9860,N_9906);
nor UO_1408 (O_1408,N_9905,N_9978);
nor UO_1409 (O_1409,N_9921,N_9818);
nor UO_1410 (O_1410,N_9898,N_9804);
nor UO_1411 (O_1411,N_9944,N_9996);
or UO_1412 (O_1412,N_9980,N_9803);
or UO_1413 (O_1413,N_9880,N_9995);
nor UO_1414 (O_1414,N_9825,N_9898);
nor UO_1415 (O_1415,N_9972,N_9851);
nand UO_1416 (O_1416,N_9808,N_9977);
nor UO_1417 (O_1417,N_9810,N_9817);
nor UO_1418 (O_1418,N_9860,N_9857);
or UO_1419 (O_1419,N_9905,N_9947);
nand UO_1420 (O_1420,N_9889,N_9857);
nor UO_1421 (O_1421,N_9843,N_9846);
nand UO_1422 (O_1422,N_9840,N_9932);
xnor UO_1423 (O_1423,N_9975,N_9848);
nand UO_1424 (O_1424,N_9925,N_9934);
and UO_1425 (O_1425,N_9963,N_9854);
xor UO_1426 (O_1426,N_9983,N_9935);
or UO_1427 (O_1427,N_9976,N_9948);
nor UO_1428 (O_1428,N_9823,N_9965);
and UO_1429 (O_1429,N_9923,N_9862);
or UO_1430 (O_1430,N_9912,N_9885);
nand UO_1431 (O_1431,N_9852,N_9963);
nand UO_1432 (O_1432,N_9893,N_9945);
nand UO_1433 (O_1433,N_9828,N_9898);
or UO_1434 (O_1434,N_9999,N_9993);
nand UO_1435 (O_1435,N_9827,N_9942);
nor UO_1436 (O_1436,N_9815,N_9900);
xnor UO_1437 (O_1437,N_9858,N_9815);
nand UO_1438 (O_1438,N_9966,N_9950);
and UO_1439 (O_1439,N_9958,N_9872);
and UO_1440 (O_1440,N_9811,N_9897);
and UO_1441 (O_1441,N_9943,N_9976);
or UO_1442 (O_1442,N_9824,N_9886);
xnor UO_1443 (O_1443,N_9983,N_9938);
nand UO_1444 (O_1444,N_9949,N_9906);
nand UO_1445 (O_1445,N_9804,N_9946);
nor UO_1446 (O_1446,N_9929,N_9892);
nand UO_1447 (O_1447,N_9946,N_9957);
nand UO_1448 (O_1448,N_9841,N_9978);
and UO_1449 (O_1449,N_9993,N_9915);
xor UO_1450 (O_1450,N_9963,N_9901);
and UO_1451 (O_1451,N_9854,N_9889);
xnor UO_1452 (O_1452,N_9873,N_9942);
nand UO_1453 (O_1453,N_9857,N_9945);
and UO_1454 (O_1454,N_9876,N_9895);
and UO_1455 (O_1455,N_9896,N_9899);
nand UO_1456 (O_1456,N_9982,N_9953);
nand UO_1457 (O_1457,N_9836,N_9934);
or UO_1458 (O_1458,N_9841,N_9906);
or UO_1459 (O_1459,N_9955,N_9860);
and UO_1460 (O_1460,N_9855,N_9967);
nand UO_1461 (O_1461,N_9848,N_9859);
and UO_1462 (O_1462,N_9987,N_9846);
nand UO_1463 (O_1463,N_9900,N_9980);
nand UO_1464 (O_1464,N_9958,N_9852);
xnor UO_1465 (O_1465,N_9971,N_9819);
and UO_1466 (O_1466,N_9975,N_9850);
or UO_1467 (O_1467,N_9832,N_9896);
and UO_1468 (O_1468,N_9941,N_9923);
nand UO_1469 (O_1469,N_9836,N_9829);
or UO_1470 (O_1470,N_9839,N_9935);
and UO_1471 (O_1471,N_9972,N_9963);
nor UO_1472 (O_1472,N_9873,N_9837);
and UO_1473 (O_1473,N_9934,N_9975);
nor UO_1474 (O_1474,N_9814,N_9998);
and UO_1475 (O_1475,N_9964,N_9863);
nor UO_1476 (O_1476,N_9984,N_9857);
and UO_1477 (O_1477,N_9990,N_9820);
nor UO_1478 (O_1478,N_9987,N_9963);
and UO_1479 (O_1479,N_9985,N_9849);
nor UO_1480 (O_1480,N_9953,N_9985);
nor UO_1481 (O_1481,N_9925,N_9829);
and UO_1482 (O_1482,N_9947,N_9820);
and UO_1483 (O_1483,N_9954,N_9880);
and UO_1484 (O_1484,N_9984,N_9823);
nand UO_1485 (O_1485,N_9921,N_9905);
nor UO_1486 (O_1486,N_9990,N_9873);
and UO_1487 (O_1487,N_9952,N_9904);
nand UO_1488 (O_1488,N_9856,N_9838);
or UO_1489 (O_1489,N_9857,N_9999);
nand UO_1490 (O_1490,N_9854,N_9869);
nor UO_1491 (O_1491,N_9809,N_9956);
or UO_1492 (O_1492,N_9802,N_9908);
or UO_1493 (O_1493,N_9916,N_9822);
or UO_1494 (O_1494,N_9963,N_9830);
nand UO_1495 (O_1495,N_9956,N_9805);
xnor UO_1496 (O_1496,N_9988,N_9910);
xor UO_1497 (O_1497,N_9832,N_9835);
and UO_1498 (O_1498,N_9935,N_9865);
or UO_1499 (O_1499,N_9846,N_9802);
endmodule