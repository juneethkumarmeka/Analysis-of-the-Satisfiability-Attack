module basic_1500_15000_2000_5_levels_5xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
or U0 (N_0,In_729,In_1395);
and U1 (N_1,In_382,In_1385);
nor U2 (N_2,In_59,In_261);
nor U3 (N_3,In_749,In_832);
nand U4 (N_4,In_398,In_430);
nor U5 (N_5,In_172,In_1336);
and U6 (N_6,In_131,In_1489);
nand U7 (N_7,In_1217,In_1309);
or U8 (N_8,In_544,In_1152);
nand U9 (N_9,In_90,In_46);
or U10 (N_10,In_1208,In_459);
or U11 (N_11,In_1308,In_677);
nor U12 (N_12,In_244,In_1268);
or U13 (N_13,In_1014,In_306);
nor U14 (N_14,In_684,In_1212);
nand U15 (N_15,In_356,In_840);
nand U16 (N_16,In_825,In_1434);
or U17 (N_17,In_942,In_1391);
or U18 (N_18,In_753,In_693);
or U19 (N_19,In_708,In_334);
or U20 (N_20,In_110,In_581);
nand U21 (N_21,In_1098,In_1362);
and U22 (N_22,In_401,In_643);
nand U23 (N_23,In_1174,In_432);
nand U24 (N_24,In_641,In_1115);
nand U25 (N_25,In_1079,In_169);
or U26 (N_26,In_828,In_966);
nand U27 (N_27,In_1193,In_409);
and U28 (N_28,In_1435,In_849);
or U29 (N_29,In_1335,In_454);
or U30 (N_30,In_616,In_488);
nor U31 (N_31,In_592,In_983);
nor U32 (N_32,In_1339,In_122);
nor U33 (N_33,In_13,In_501);
nand U34 (N_34,In_967,In_293);
and U35 (N_35,In_1191,In_628);
nand U36 (N_36,In_972,In_1293);
or U37 (N_37,In_1388,In_882);
nand U38 (N_38,In_299,In_1457);
nor U39 (N_39,In_580,In_253);
nor U40 (N_40,In_880,In_337);
and U41 (N_41,In_878,In_396);
or U42 (N_42,In_328,In_1414);
nor U43 (N_43,In_370,In_745);
nand U44 (N_44,In_309,In_1478);
or U45 (N_45,In_417,In_153);
nand U46 (N_46,In_720,In_702);
nor U47 (N_47,In_130,In_518);
nor U48 (N_48,In_197,In_671);
or U49 (N_49,In_1473,In_1360);
or U50 (N_50,In_1342,In_845);
nor U51 (N_51,In_158,In_167);
nor U52 (N_52,In_460,In_248);
nand U53 (N_53,In_272,In_848);
nand U54 (N_54,In_111,In_116);
nor U55 (N_55,In_1400,In_723);
nand U56 (N_56,In_857,In_60);
xnor U57 (N_57,In_1348,In_388);
nand U58 (N_58,In_807,In_639);
nor U59 (N_59,In_1330,In_215);
and U60 (N_60,In_1428,In_222);
or U61 (N_61,In_95,In_1124);
or U62 (N_62,In_1323,In_319);
nand U63 (N_63,In_1498,In_1034);
and U64 (N_64,In_593,In_70);
and U65 (N_65,In_663,In_1017);
and U66 (N_66,In_860,In_66);
or U67 (N_67,In_1039,In_19);
or U68 (N_68,In_511,In_1470);
nand U69 (N_69,In_203,In_837);
nand U70 (N_70,In_1029,In_785);
or U71 (N_71,In_926,In_870);
xor U72 (N_72,In_771,In_1369);
and U73 (N_73,In_662,In_107);
nand U74 (N_74,In_1190,In_202);
nor U75 (N_75,In_850,In_41);
or U76 (N_76,In_188,In_455);
or U77 (N_77,In_665,In_226);
and U78 (N_78,In_548,In_1256);
and U79 (N_79,In_352,In_638);
and U80 (N_80,In_77,In_1363);
nand U81 (N_81,In_143,In_569);
xor U82 (N_82,In_264,In_217);
xor U83 (N_83,In_599,In_447);
nand U84 (N_84,In_1021,In_1444);
nand U85 (N_85,In_1225,In_1067);
or U86 (N_86,In_446,In_1317);
nor U87 (N_87,In_590,In_200);
and U88 (N_88,In_170,In_79);
and U89 (N_89,In_26,In_1277);
and U90 (N_90,In_386,In_274);
nand U91 (N_91,In_1340,In_100);
nand U92 (N_92,In_586,In_791);
nand U93 (N_93,In_414,In_265);
nor U94 (N_94,In_740,In_193);
nand U95 (N_95,In_783,In_698);
and U96 (N_96,In_1126,In_814);
nand U97 (N_97,In_890,In_1450);
nand U98 (N_98,In_503,In_44);
or U99 (N_99,In_1022,In_139);
or U100 (N_100,In_751,In_685);
nor U101 (N_101,In_50,In_1147);
and U102 (N_102,In_573,In_379);
and U103 (N_103,In_959,In_10);
nand U104 (N_104,In_423,In_1390);
and U105 (N_105,In_1297,In_376);
xnor U106 (N_106,In_320,In_52);
nand U107 (N_107,In_559,In_689);
or U108 (N_108,In_636,In_498);
nor U109 (N_109,In_822,In_1490);
or U110 (N_110,In_1194,In_457);
or U111 (N_111,In_1266,In_24);
and U112 (N_112,In_211,In_739);
and U113 (N_113,In_875,In_129);
or U114 (N_114,In_144,In_1180);
nor U115 (N_115,In_1040,In_932);
and U116 (N_116,In_87,In_1267);
xnor U117 (N_117,In_801,In_1387);
and U118 (N_118,In_325,In_735);
or U119 (N_119,In_919,In_744);
xor U120 (N_120,In_1084,In_1221);
nand U121 (N_121,In_1461,In_1062);
and U122 (N_122,In_1135,In_402);
nand U123 (N_123,In_1047,In_1337);
and U124 (N_124,In_895,In_658);
nor U125 (N_125,In_476,In_434);
and U126 (N_126,In_914,In_764);
and U127 (N_127,In_615,In_618);
xor U128 (N_128,In_726,In_1386);
xnor U129 (N_129,In_601,In_540);
nor U130 (N_130,In_61,In_271);
nand U131 (N_131,In_1006,In_977);
nand U132 (N_132,In_113,In_637);
nand U133 (N_133,In_1379,In_28);
and U134 (N_134,In_176,In_427);
and U135 (N_135,In_683,In_206);
xnor U136 (N_136,In_561,In_1364);
and U137 (N_137,In_1482,In_492);
and U138 (N_138,In_1455,In_329);
nor U139 (N_139,In_247,In_268);
nor U140 (N_140,In_1168,In_763);
and U141 (N_141,In_437,In_1321);
and U142 (N_142,In_408,In_886);
nor U143 (N_143,In_1198,In_709);
xor U144 (N_144,In_536,In_236);
or U145 (N_145,In_691,In_201);
nand U146 (N_146,In_1311,In_350);
nor U147 (N_147,In_1465,In_951);
or U148 (N_148,In_1245,In_54);
or U149 (N_149,In_1258,In_1100);
nor U150 (N_150,In_1015,In_1052);
and U151 (N_151,In_1413,In_1378);
and U152 (N_152,In_578,In_574);
nand U153 (N_153,In_8,In_1081);
nor U154 (N_154,In_1296,In_101);
nand U155 (N_155,In_1496,In_1218);
nand U156 (N_156,In_522,In_1398);
nor U157 (N_157,In_515,In_1043);
or U158 (N_158,In_589,In_1046);
nor U159 (N_159,In_1058,In_642);
xor U160 (N_160,In_1246,In_1053);
nand U161 (N_161,In_1204,In_680);
nand U162 (N_162,In_533,In_703);
or U163 (N_163,In_542,In_302);
nand U164 (N_164,In_757,In_519);
and U165 (N_165,In_975,In_1289);
nor U166 (N_166,In_1487,In_1264);
nand U167 (N_167,In_96,In_15);
or U168 (N_168,In_734,In_1403);
or U169 (N_169,In_1109,In_1236);
nor U170 (N_170,In_109,In_681);
and U171 (N_171,In_997,In_464);
nor U172 (N_172,In_1005,In_190);
and U173 (N_173,In_961,In_1057);
nor U174 (N_174,In_32,In_338);
and U175 (N_175,In_797,In_1442);
nand U176 (N_176,In_450,In_1026);
nand U177 (N_177,In_300,In_1083);
and U178 (N_178,In_173,In_847);
or U179 (N_179,In_1300,In_512);
or U180 (N_180,In_359,In_1430);
or U181 (N_181,In_864,In_214);
or U182 (N_182,In_944,In_965);
or U183 (N_183,In_583,In_1106);
xnor U184 (N_184,In_678,In_92);
nand U185 (N_185,In_867,In_768);
or U186 (N_186,In_56,In_1088);
xnor U187 (N_187,In_1423,In_1054);
xnor U188 (N_188,In_1214,In_1304);
nand U189 (N_189,In_899,In_547);
nand U190 (N_190,In_1351,In_315);
nand U191 (N_191,In_587,In_968);
or U192 (N_192,In_818,In_1234);
nor U193 (N_193,In_378,In_1485);
nand U194 (N_194,In_1161,In_842);
and U195 (N_195,In_1279,In_62);
or U196 (N_196,In_324,In_1071);
or U197 (N_197,In_999,In_1154);
or U198 (N_198,In_520,In_808);
nand U199 (N_199,In_854,In_1238);
and U200 (N_200,In_456,In_1068);
nor U201 (N_201,In_963,In_4);
nand U202 (N_202,In_413,In_876);
and U203 (N_203,In_83,In_672);
xor U204 (N_204,In_91,In_1099);
and U205 (N_205,In_1497,In_149);
and U206 (N_206,In_635,In_1272);
and U207 (N_207,In_12,In_531);
nor U208 (N_208,In_1024,In_357);
nand U209 (N_209,In_955,In_1305);
nor U210 (N_210,In_369,In_481);
nor U211 (N_211,In_1260,In_1032);
nor U212 (N_212,In_688,In_551);
nand U213 (N_213,In_534,In_1295);
and U214 (N_214,In_935,In_567);
nand U215 (N_215,In_1185,In_1493);
or U216 (N_216,In_1073,In_910);
nand U217 (N_217,In_1326,In_1105);
nor U218 (N_218,In_68,In_995);
and U219 (N_219,In_1050,In_354);
and U220 (N_220,In_556,In_1247);
nor U221 (N_221,In_1449,In_1285);
and U222 (N_222,In_243,In_873);
nand U223 (N_223,In_1231,In_404);
nor U224 (N_224,In_106,In_348);
or U225 (N_225,In_51,In_855);
or U226 (N_226,In_1254,In_554);
or U227 (N_227,In_1086,In_1404);
nor U228 (N_228,In_523,In_988);
nand U229 (N_229,In_1411,In_546);
nand U230 (N_230,In_562,In_349);
and U231 (N_231,In_532,In_762);
or U232 (N_232,In_970,In_1156);
nor U233 (N_233,In_1440,In_998);
xor U234 (N_234,In_861,In_993);
nand U235 (N_235,In_1199,In_1007);
and U236 (N_236,In_1298,In_537);
and U237 (N_237,In_513,In_841);
or U238 (N_238,In_543,In_1359);
and U239 (N_239,In_45,In_697);
and U240 (N_240,In_669,In_1275);
nand U241 (N_241,In_256,In_507);
and U242 (N_242,In_1060,In_727);
nor U243 (N_243,In_1325,In_1002);
xor U244 (N_244,In_482,In_1331);
and U245 (N_245,In_1276,In_145);
xor U246 (N_246,In_1028,In_622);
or U247 (N_247,In_812,In_1251);
xnor U248 (N_248,In_1358,In_911);
nor U249 (N_249,In_939,In_1460);
and U250 (N_250,In_508,In_715);
nand U251 (N_251,In_1157,In_953);
xnor U252 (N_252,In_152,In_535);
and U253 (N_253,In_168,In_528);
nand U254 (N_254,In_1091,In_679);
nand U255 (N_255,In_58,In_611);
nand U256 (N_256,In_851,In_1352);
or U257 (N_257,In_314,In_815);
nor U258 (N_258,In_1408,In_405);
nor U259 (N_259,In_776,In_391);
nor U260 (N_260,In_1023,In_1063);
nand U261 (N_261,In_392,In_1030);
or U262 (N_262,In_245,In_853);
nand U263 (N_263,In_1409,In_1322);
nand U264 (N_264,In_332,In_1243);
nor U265 (N_265,In_541,In_1294);
nor U266 (N_266,In_42,In_7);
and U267 (N_267,In_1436,In_1255);
nand U268 (N_268,In_141,In_1009);
xor U269 (N_269,In_631,In_529);
or U270 (N_270,In_1468,In_666);
nand U271 (N_271,In_65,In_277);
nor U272 (N_272,In_18,In_1376);
nand U273 (N_273,In_805,In_279);
and U274 (N_274,In_1103,In_948);
and U275 (N_275,In_571,In_108);
nor U276 (N_276,In_155,In_725);
and U277 (N_277,In_322,In_1159);
and U278 (N_278,In_603,In_453);
and U279 (N_279,In_916,In_1175);
and U280 (N_280,In_557,In_228);
and U281 (N_281,In_136,In_227);
and U282 (N_282,In_287,In_1224);
nand U283 (N_283,In_1426,In_1158);
and U284 (N_284,In_598,In_1119);
and U285 (N_285,In_467,In_1282);
nand U286 (N_286,In_124,In_1371);
nor U287 (N_287,In_675,In_1059);
or U288 (N_288,In_1278,In_941);
nor U289 (N_289,In_539,In_755);
or U290 (N_290,In_112,In_1116);
nor U291 (N_291,In_1472,In_84);
nor U292 (N_292,In_415,In_572);
or U293 (N_293,In_527,In_1265);
or U294 (N_294,In_651,In_275);
or U295 (N_295,In_728,In_255);
nor U296 (N_296,In_353,In_400);
nor U297 (N_297,In_1458,In_1469);
and U298 (N_298,In_1447,In_741);
or U299 (N_299,In_1270,In_399);
and U300 (N_300,In_1454,In_746);
xor U301 (N_301,In_135,In_421);
xnor U302 (N_302,In_1149,In_907);
nor U303 (N_303,In_1417,In_146);
or U304 (N_304,In_700,In_496);
nor U305 (N_305,In_1405,In_291);
and U306 (N_306,In_385,In_260);
xor U307 (N_307,In_920,In_609);
nor U308 (N_308,In_1120,In_1075);
nand U309 (N_309,In_1074,In_270);
nand U310 (N_310,In_711,In_162);
and U311 (N_311,In_1499,In_219);
or U312 (N_312,In_1368,In_710);
or U313 (N_313,In_984,In_986);
xnor U314 (N_314,In_37,In_1025);
and U315 (N_315,In_363,In_1000);
and U316 (N_316,In_411,In_819);
nor U317 (N_317,In_1488,In_1222);
nand U318 (N_318,In_246,In_171);
or U319 (N_319,In_1087,In_80);
nor U320 (N_320,In_436,In_1189);
xor U321 (N_321,In_1286,In_67);
and U322 (N_322,In_184,In_954);
xor U323 (N_323,In_316,In_502);
and U324 (N_324,In_281,In_121);
or U325 (N_325,In_833,In_505);
nand U326 (N_326,In_748,In_1200);
or U327 (N_327,In_1483,In_1301);
nand U328 (N_328,In_462,In_1082);
nand U329 (N_329,In_294,In_150);
nor U330 (N_330,In_1128,In_1365);
nand U331 (N_331,In_483,In_1357);
and U332 (N_332,In_806,In_105);
and U333 (N_333,In_1010,In_1101);
nand U334 (N_334,In_667,In_93);
nand U335 (N_335,In_766,In_553);
nand U336 (N_336,In_835,In_389);
nor U337 (N_337,In_1142,In_1065);
and U338 (N_338,In_1038,In_923);
nand U339 (N_339,In_441,In_394);
nand U340 (N_340,In_1345,In_577);
or U341 (N_341,In_278,In_1077);
nor U342 (N_342,In_254,In_1003);
nand U343 (N_343,In_290,In_39);
or U344 (N_344,In_1441,In_591);
nand U345 (N_345,In_22,In_191);
nor U346 (N_346,In_1166,In_310);
or U347 (N_347,In_269,In_321);
xor U348 (N_348,In_1382,In_27);
xnor U349 (N_349,In_1179,In_686);
nor U350 (N_350,In_412,In_629);
nand U351 (N_351,In_366,In_355);
nand U352 (N_352,In_645,In_1480);
and U353 (N_353,In_584,In_836);
or U354 (N_354,In_605,In_881);
and U355 (N_355,In_904,In_1355);
nor U356 (N_356,In_1031,In_985);
or U357 (N_357,In_444,In_1096);
nand U358 (N_358,In_119,In_733);
or U359 (N_359,In_474,In_1452);
and U360 (N_360,In_208,In_132);
and U361 (N_361,In_403,In_380);
and U362 (N_362,In_1089,In_885);
or U363 (N_363,In_38,In_1133);
or U364 (N_364,In_829,In_189);
xor U365 (N_365,In_594,In_371);
or U366 (N_366,In_844,In_1292);
xnor U367 (N_367,In_339,In_1249);
or U368 (N_368,In_1377,In_266);
nor U369 (N_369,In_1397,In_687);
nor U370 (N_370,In_494,In_524);
or U371 (N_371,In_1248,In_81);
nand U372 (N_372,In_660,In_1134);
nand U373 (N_373,In_134,In_267);
nor U374 (N_374,In_1299,In_1216);
or U375 (N_375,In_296,In_486);
nand U376 (N_376,In_921,In_1011);
nor U377 (N_377,In_1284,In_231);
nand U378 (N_378,In_47,In_318);
or U379 (N_379,In_994,In_1164);
nand U380 (N_380,In_929,In_1240);
xor U381 (N_381,In_902,In_989);
nor U382 (N_382,In_1412,In_458);
and U383 (N_383,In_160,In_699);
nand U384 (N_384,In_649,In_1195);
and U385 (N_385,In_1192,In_416);
nand U386 (N_386,In_239,In_1132);
nor U387 (N_387,In_1257,In_816);
or U388 (N_388,In_722,In_1232);
nor U389 (N_389,In_351,In_1016);
and U390 (N_390,In_1250,In_826);
or U391 (N_391,In_862,In_30);
or U392 (N_392,In_730,In_117);
nor U393 (N_393,In_621,In_179);
and U394 (N_394,In_1113,In_510);
xnor U395 (N_395,In_140,In_1437);
nor U396 (N_396,In_509,In_104);
or U397 (N_397,In_644,In_646);
and U398 (N_398,In_283,In_786);
xnor U399 (N_399,In_465,In_971);
xor U400 (N_400,In_956,In_804);
nand U401 (N_401,In_387,In_1112);
xnor U402 (N_402,In_282,In_126);
or U403 (N_403,In_1061,In_1035);
xnor U404 (N_404,In_295,In_1463);
and U405 (N_405,In_1415,In_1269);
or U406 (N_406,In_964,In_1211);
nor U407 (N_407,In_33,In_1080);
xor U408 (N_408,In_1045,In_1181);
nor U409 (N_409,In_341,In_224);
and U410 (N_410,In_262,In_1036);
nand U411 (N_411,In_940,In_345);
or U412 (N_412,In_1271,In_1140);
or U413 (N_413,In_1280,In_1102);
nor U414 (N_414,In_996,In_1219);
nor U415 (N_415,In_887,In_297);
nand U416 (N_416,In_682,In_336);
nor U417 (N_417,In_588,In_617);
and U418 (N_418,In_1316,In_207);
nor U419 (N_419,In_506,In_990);
nand U420 (N_420,In_410,In_1392);
nor U421 (N_421,In_1462,In_795);
or U422 (N_422,In_1464,In_1055);
and U423 (N_423,In_154,In_470);
or U424 (N_424,In_924,In_273);
and U425 (N_425,In_576,In_419);
and U426 (N_426,In_186,In_128);
and U427 (N_427,In_1259,In_491);
nor U428 (N_428,In_824,In_690);
or U429 (N_429,In_118,In_838);
nor U430 (N_430,In_305,In_73);
and U431 (N_431,In_619,In_326);
xnor U432 (N_432,In_487,In_289);
and U433 (N_433,In_1303,In_1121);
and U434 (N_434,In_1475,In_1018);
nor U435 (N_435,In_1420,In_868);
and U436 (N_436,In_1173,In_1427);
nand U437 (N_437,In_1076,In_323);
and U438 (N_438,In_650,In_1093);
nor U439 (N_439,In_72,In_792);
and U440 (N_440,In_312,In_909);
or U441 (N_441,In_1008,In_879);
nor U442 (N_442,In_36,In_659);
nor U443 (N_443,In_374,In_1373);
nor U444 (N_444,In_525,In_1261);
nor U445 (N_445,In_1123,In_846);
and U446 (N_446,In_767,In_630);
or U447 (N_447,In_859,In_774);
nand U448 (N_448,In_183,In_946);
or U449 (N_449,In_57,In_159);
or U450 (N_450,In_793,In_865);
or U451 (N_451,In_1451,In_428);
xnor U452 (N_452,In_794,In_1162);
nor U453 (N_453,In_1394,In_1453);
or U454 (N_454,In_1027,In_839);
nor U455 (N_455,In_229,In_375);
nand U456 (N_456,In_195,In_976);
and U457 (N_457,In_1235,In_1407);
xor U458 (N_458,In_1344,In_969);
xnor U459 (N_459,In_898,In_1228);
xor U460 (N_460,In_877,In_1206);
nor U461 (N_461,In_234,In_1481);
and U462 (N_462,In_552,In_180);
or U463 (N_463,In_1477,In_1033);
nand U464 (N_464,In_1446,In_182);
and U465 (N_465,In_1237,In_913);
nand U466 (N_466,In_790,In_397);
and U467 (N_467,In_1486,In_406);
nor U468 (N_468,In_485,In_298);
or U469 (N_469,In_1341,In_435);
nor U470 (N_470,In_1374,In_575);
nand U471 (N_471,In_704,In_775);
and U472 (N_472,In_670,In_811);
and U473 (N_473,In_668,In_938);
nand U474 (N_474,In_1107,In_1252);
and U475 (N_475,In_438,In_1474);
or U476 (N_476,In_933,In_1416);
nor U477 (N_477,In_779,In_550);
or U478 (N_478,In_987,In_164);
nor U479 (N_479,In_657,In_76);
nor U480 (N_480,In_1090,In_908);
nand U481 (N_481,In_1419,In_177);
nand U482 (N_482,In_736,In_1233);
xnor U483 (N_483,In_614,In_521);
or U484 (N_484,In_1092,In_241);
or U485 (N_485,In_1160,In_1445);
or U486 (N_486,In_311,In_213);
nor U487 (N_487,In_205,In_1406);
and U488 (N_488,In_174,In_1318);
nand U489 (N_489,In_1306,In_252);
and U490 (N_490,In_468,In_196);
or U491 (N_491,In_1494,In_915);
nand U492 (N_492,In_1184,In_1422);
nor U493 (N_493,In_156,In_752);
and U494 (N_494,In_218,In_1383);
and U495 (N_495,In_640,In_706);
or U496 (N_496,In_69,In_1145);
xnor U497 (N_497,In_14,In_495);
nand U498 (N_498,In_1049,In_820);
nor U499 (N_499,In_654,In_1001);
nor U500 (N_500,In_934,In_1202);
nand U501 (N_501,In_1085,In_479);
nor U502 (N_502,In_308,In_1114);
and U503 (N_503,In_478,In_897);
and U504 (N_504,In_451,In_759);
and U505 (N_505,In_232,In_1226);
nor U506 (N_506,In_1431,In_16);
nand U507 (N_507,In_365,In_664);
or U508 (N_508,In_418,In_760);
nand U509 (N_509,In_157,In_673);
nand U510 (N_510,In_676,In_204);
or U511 (N_511,In_1197,In_891);
and U512 (N_512,In_11,In_390);
xor U513 (N_513,In_1108,In_43);
xnor U514 (N_514,In_743,In_55);
and U515 (N_515,In_1349,In_1401);
and U516 (N_516,In_863,In_1424);
xnor U517 (N_517,In_883,In_463);
nand U518 (N_518,In_777,In_49);
and U519 (N_519,In_943,In_992);
or U520 (N_520,In_1223,In_781);
xor U521 (N_521,In_185,In_737);
or U522 (N_522,In_624,In_221);
nor U523 (N_523,In_595,In_978);
nor U524 (N_524,In_330,In_788);
or U525 (N_525,In_303,In_716);
nand U526 (N_526,In_71,In_1467);
and U527 (N_527,In_425,In_344);
and U528 (N_528,In_99,In_1095);
or U529 (N_529,In_517,In_475);
xnor U530 (N_530,In_1312,In_1253);
xnor U531 (N_531,In_653,In_1069);
or U532 (N_532,In_123,In_94);
xor U533 (N_533,In_362,In_1361);
or U534 (N_534,In_545,In_979);
and U535 (N_535,In_165,In_604);
nor U536 (N_536,In_340,In_596);
nand U537 (N_537,In_560,In_17);
and U538 (N_538,In_166,In_821);
nor U539 (N_539,In_23,In_1443);
nand U540 (N_540,In_500,In_1334);
or U541 (N_541,In_216,In_623);
or U542 (N_542,In_1118,In_866);
nor U543 (N_543,In_613,In_1429);
and U544 (N_544,In_284,In_1110);
or U545 (N_545,In_442,In_490);
or U546 (N_546,In_1186,In_610);
nor U547 (N_547,In_1170,In_1042);
nor U548 (N_548,In_242,In_1315);
nor U549 (N_549,In_1210,In_960);
xnor U550 (N_550,In_1072,In_114);
xnor U551 (N_551,In_803,In_360);
xnor U552 (N_552,In_125,In_431);
nor U553 (N_553,In_884,In_335);
nand U554 (N_554,In_754,In_74);
nor U555 (N_555,In_1310,In_694);
nand U556 (N_556,In_980,In_634);
and U557 (N_557,In_381,In_912);
and U558 (N_558,In_1122,In_1290);
nor U559 (N_559,In_420,In_1418);
or U560 (N_560,In_872,In_1182);
nand U561 (N_561,In_473,In_1262);
or U562 (N_562,In_6,In_1187);
and U563 (N_563,In_1239,In_656);
and U564 (N_564,In_1287,In_288);
and U565 (N_565,In_1350,In_1343);
nand U566 (N_566,In_280,In_452);
xnor U567 (N_567,In_151,In_1155);
or U568 (N_568,In_220,In_1476);
and U569 (N_569,In_276,In_770);
and U570 (N_570,In_719,In_212);
and U571 (N_571,In_422,In_199);
nand U572 (N_572,In_750,In_830);
nand U573 (N_573,In_652,In_780);
nor U574 (N_574,In_343,In_597);
and U575 (N_575,In_1425,In_765);
and U576 (N_576,In_707,In_789);
and U577 (N_577,In_800,In_1066);
nor U578 (N_578,In_831,In_633);
or U579 (N_579,In_233,In_1130);
xnor U580 (N_580,In_307,In_133);
nor U581 (N_581,In_250,In_1205);
nor U582 (N_582,In_973,In_1051);
nand U583 (N_583,In_148,In_1203);
xnor U584 (N_584,In_249,In_1274);
nor U585 (N_585,In_1136,In_950);
nor U586 (N_586,In_692,In_936);
or U587 (N_587,In_439,In_1353);
xnor U588 (N_588,In_1144,In_856);
xnor U589 (N_589,In_982,In_802);
and U590 (N_590,In_1048,In_1078);
or U591 (N_591,In_477,In_187);
or U592 (N_592,In_1167,In_799);
nor U593 (N_593,In_620,In_424);
or U594 (N_594,In_1020,In_103);
nor U595 (N_595,In_1139,In_88);
nor U596 (N_596,In_1433,In_705);
nor U597 (N_597,In_563,In_957);
or U598 (N_598,In_1484,In_1196);
nor U599 (N_599,In_471,In_1380);
xor U600 (N_600,In_796,In_896);
and U601 (N_601,In_1125,In_1176);
nand U602 (N_602,In_632,In_695);
nand U603 (N_603,In_772,In_1273);
nand U604 (N_604,In_555,In_1177);
nor U605 (N_605,In_1056,In_1456);
nor U606 (N_606,In_1044,In_773);
or U607 (N_607,In_346,In_958);
or U608 (N_608,In_263,In_558);
and U609 (N_609,In_301,In_1438);
or U610 (N_610,In_5,In_426);
or U611 (N_611,In_1004,In_1207);
or U612 (N_612,In_1319,In_1466);
nor U613 (N_613,In_1372,In_327);
and U614 (N_614,In_1313,In_1384);
nand U615 (N_615,In_869,In_504);
nor U616 (N_616,In_0,In_383);
nor U617 (N_617,In_102,In_949);
nand U618 (N_618,In_1097,In_1104);
or U619 (N_619,In_433,In_1399);
xor U620 (N_620,In_29,In_251);
nand U621 (N_621,In_358,In_717);
nor U622 (N_622,In_484,In_1242);
or U623 (N_623,In_1183,In_568);
xnor U624 (N_624,In_384,In_372);
nor U625 (N_625,In_930,In_1129);
or U626 (N_626,In_1479,In_443);
nand U627 (N_627,In_718,In_361);
nor U628 (N_628,In_564,In_1410);
nor U629 (N_629,In_445,In_1327);
nand U630 (N_630,In_86,In_21);
nand U631 (N_631,In_917,In_778);
nor U632 (N_632,In_209,In_655);
nor U633 (N_633,In_858,In_210);
xor U634 (N_634,In_1230,In_991);
nor U635 (N_635,In_585,In_1459);
nor U636 (N_636,In_1421,In_701);
and U637 (N_637,In_514,In_1320);
nand U638 (N_638,In_1138,In_285);
nand U639 (N_639,In_674,In_175);
nor U640 (N_640,In_461,In_448);
nor U641 (N_641,In_64,In_600);
nand U642 (N_642,In_1070,In_35);
nor U643 (N_643,In_538,In_48);
or U644 (N_644,In_1111,In_782);
nand U645 (N_645,In_570,In_25);
nand U646 (N_646,In_1302,In_813);
nor U647 (N_647,In_1178,In_627);
nand U648 (N_648,In_901,In_810);
xor U649 (N_649,In_1151,In_178);
or U650 (N_650,In_952,In_1165);
and U651 (N_651,In_1019,In_922);
nor U652 (N_652,In_1143,In_1495);
nand U653 (N_653,In_1281,In_142);
nand U654 (N_654,In_97,In_713);
or U655 (N_655,In_286,In_1329);
nor U656 (N_656,In_1324,In_1171);
and U657 (N_657,In_2,In_1094);
nand U658 (N_658,In_1064,In_918);
nand U659 (N_659,In_225,In_1354);
or U660 (N_660,In_1153,In_1215);
nand U661 (N_661,In_1169,In_1491);
nand U662 (N_662,In_115,In_602);
nor U663 (N_663,In_1,In_606);
xor U664 (N_664,In_647,In_894);
xor U665 (N_665,In_787,In_742);
nand U666 (N_666,In_756,In_1241);
nand U667 (N_667,In_937,In_259);
and U668 (N_668,In_1213,In_900);
nand U669 (N_669,In_127,In_364);
xnor U670 (N_670,In_138,In_395);
nand U671 (N_671,In_852,In_827);
nor U672 (N_672,In_738,In_347);
nor U673 (N_673,In_549,In_721);
nor U674 (N_674,In_1188,In_469);
xnor U675 (N_675,In_1381,In_342);
or U676 (N_676,In_89,In_198);
xnor U677 (N_677,In_834,In_784);
nand U678 (N_678,In_731,In_1141);
nand U679 (N_679,In_85,In_161);
xnor U680 (N_680,In_1263,In_892);
nand U681 (N_681,In_927,In_931);
and U682 (N_682,In_1492,In_1037);
nand U683 (N_683,In_75,In_1471);
nand U684 (N_684,In_947,In_317);
nor U685 (N_685,In_1288,In_1146);
nor U686 (N_686,In_607,In_579);
xnor U687 (N_687,In_1346,In_903);
nand U688 (N_688,In_1338,In_1375);
xor U689 (N_689,In_817,In_237);
and U690 (N_690,In_292,In_1117);
or U691 (N_691,In_696,In_712);
or U692 (N_692,In_429,In_472);
or U693 (N_693,In_230,In_3);
or U694 (N_694,In_769,In_809);
nor U695 (N_695,In_1356,In_373);
or U696 (N_696,In_1367,In_1013);
nand U697 (N_697,In_313,In_1332);
nor U698 (N_698,In_1201,In_9);
nor U699 (N_699,In_1366,In_1291);
or U700 (N_700,In_530,In_1396);
or U701 (N_701,In_449,In_1333);
or U702 (N_702,In_874,In_238);
nor U703 (N_703,In_928,In_888);
and U704 (N_704,In_889,In_1172);
and U705 (N_705,In_582,In_377);
nand U706 (N_706,In_724,In_526);
or U707 (N_707,In_63,In_1012);
xor U708 (N_708,In_565,In_823);
nor U709 (N_709,In_714,In_1127);
or U710 (N_710,In_1328,In_1148);
or U711 (N_711,In_747,In_905);
nand U712 (N_712,In_367,In_368);
nand U713 (N_713,In_925,In_192);
xor U714 (N_714,In_906,In_1163);
nor U715 (N_715,In_1307,In_333);
nor U716 (N_716,In_1209,In_78);
and U717 (N_717,In_407,In_147);
nand U718 (N_718,In_732,In_1389);
and U719 (N_719,In_608,In_1314);
nand U720 (N_720,In_493,In_120);
or U721 (N_721,In_1229,In_626);
and U722 (N_722,In_258,In_1131);
xnor U723 (N_723,In_945,In_1439);
and U724 (N_724,In_981,In_34);
nor U725 (N_725,In_1220,In_758);
nor U726 (N_726,In_1432,In_194);
nor U727 (N_727,In_1393,In_1448);
nand U728 (N_728,In_1137,In_798);
and U729 (N_729,In_466,In_962);
nand U730 (N_730,In_1283,In_648);
or U731 (N_731,In_181,In_1041);
or U732 (N_732,In_1150,In_843);
or U733 (N_733,In_499,In_516);
and U734 (N_734,In_235,In_1227);
and U735 (N_735,In_1347,In_1244);
or U736 (N_736,In_53,In_440);
nor U737 (N_737,In_257,In_223);
xnor U738 (N_738,In_612,In_893);
nand U739 (N_739,In_40,In_240);
or U740 (N_740,In_625,In_871);
and U741 (N_741,In_82,In_98);
nor U742 (N_742,In_661,In_31);
nor U743 (N_743,In_761,In_331);
nand U744 (N_744,In_974,In_489);
or U745 (N_745,In_20,In_1370);
nand U746 (N_746,In_163,In_566);
nor U747 (N_747,In_137,In_304);
nor U748 (N_748,In_393,In_1402);
or U749 (N_749,In_480,In_497);
xor U750 (N_750,In_190,In_1252);
and U751 (N_751,In_471,In_358);
nor U752 (N_752,In_319,In_8);
or U753 (N_753,In_566,In_1277);
nand U754 (N_754,In_871,In_598);
nor U755 (N_755,In_1296,In_1120);
or U756 (N_756,In_537,In_1398);
nor U757 (N_757,In_1283,In_189);
or U758 (N_758,In_580,In_742);
nand U759 (N_759,In_285,In_1471);
and U760 (N_760,In_644,In_492);
nand U761 (N_761,In_1374,In_725);
nor U762 (N_762,In_902,In_965);
xnor U763 (N_763,In_525,In_1014);
or U764 (N_764,In_545,In_91);
xor U765 (N_765,In_398,In_312);
nand U766 (N_766,In_994,In_1291);
and U767 (N_767,In_257,In_381);
and U768 (N_768,In_1352,In_145);
nor U769 (N_769,In_940,In_271);
nand U770 (N_770,In_787,In_1075);
or U771 (N_771,In_292,In_1277);
nand U772 (N_772,In_487,In_448);
and U773 (N_773,In_416,In_389);
nor U774 (N_774,In_1372,In_1207);
or U775 (N_775,In_676,In_183);
xnor U776 (N_776,In_1374,In_1170);
nor U777 (N_777,In_963,In_15);
xnor U778 (N_778,In_754,In_1319);
nand U779 (N_779,In_1486,In_1257);
and U780 (N_780,In_167,In_416);
xor U781 (N_781,In_373,In_200);
nand U782 (N_782,In_553,In_300);
nor U783 (N_783,In_1036,In_1396);
nand U784 (N_784,In_575,In_881);
nand U785 (N_785,In_296,In_998);
nor U786 (N_786,In_995,In_737);
nand U787 (N_787,In_1455,In_760);
and U788 (N_788,In_529,In_634);
nor U789 (N_789,In_484,In_1425);
nor U790 (N_790,In_1446,In_173);
nor U791 (N_791,In_1020,In_1289);
and U792 (N_792,In_702,In_594);
xnor U793 (N_793,In_24,In_480);
or U794 (N_794,In_88,In_134);
nor U795 (N_795,In_1334,In_278);
nand U796 (N_796,In_332,In_1312);
or U797 (N_797,In_1361,In_461);
nand U798 (N_798,In_613,In_1477);
nand U799 (N_799,In_806,In_1398);
nor U800 (N_800,In_366,In_533);
nor U801 (N_801,In_552,In_422);
xnor U802 (N_802,In_1387,In_980);
or U803 (N_803,In_366,In_901);
nand U804 (N_804,In_899,In_128);
and U805 (N_805,In_816,In_93);
and U806 (N_806,In_40,In_839);
nand U807 (N_807,In_132,In_1163);
and U808 (N_808,In_858,In_266);
and U809 (N_809,In_1006,In_1499);
nand U810 (N_810,In_1156,In_1165);
nor U811 (N_811,In_146,In_1478);
nor U812 (N_812,In_67,In_161);
nand U813 (N_813,In_647,In_952);
or U814 (N_814,In_910,In_387);
nor U815 (N_815,In_745,In_402);
nand U816 (N_816,In_8,In_1430);
and U817 (N_817,In_246,In_772);
xor U818 (N_818,In_923,In_1189);
nand U819 (N_819,In_592,In_1206);
xor U820 (N_820,In_3,In_1116);
or U821 (N_821,In_185,In_172);
or U822 (N_822,In_643,In_316);
or U823 (N_823,In_426,In_734);
nand U824 (N_824,In_442,In_627);
and U825 (N_825,In_560,In_1083);
xnor U826 (N_826,In_1041,In_566);
xor U827 (N_827,In_911,In_1480);
nand U828 (N_828,In_1497,In_1114);
and U829 (N_829,In_1318,In_1482);
xnor U830 (N_830,In_905,In_938);
or U831 (N_831,In_950,In_514);
or U832 (N_832,In_794,In_337);
nand U833 (N_833,In_1256,In_594);
nand U834 (N_834,In_422,In_1027);
or U835 (N_835,In_1217,In_60);
or U836 (N_836,In_146,In_1493);
xnor U837 (N_837,In_980,In_582);
or U838 (N_838,In_1169,In_1330);
and U839 (N_839,In_33,In_1411);
nor U840 (N_840,In_365,In_1463);
nand U841 (N_841,In_109,In_498);
or U842 (N_842,In_893,In_412);
nor U843 (N_843,In_238,In_26);
and U844 (N_844,In_480,In_1358);
nand U845 (N_845,In_877,In_96);
and U846 (N_846,In_534,In_453);
and U847 (N_847,In_870,In_11);
nand U848 (N_848,In_468,In_757);
nor U849 (N_849,In_1343,In_896);
nand U850 (N_850,In_972,In_1330);
nor U851 (N_851,In_1010,In_1294);
xor U852 (N_852,In_659,In_211);
nand U853 (N_853,In_914,In_1353);
xnor U854 (N_854,In_236,In_353);
nor U855 (N_855,In_1189,In_969);
xor U856 (N_856,In_475,In_152);
nand U857 (N_857,In_265,In_1172);
nor U858 (N_858,In_1245,In_716);
nand U859 (N_859,In_760,In_405);
nand U860 (N_860,In_1125,In_423);
or U861 (N_861,In_238,In_647);
and U862 (N_862,In_547,In_1003);
nor U863 (N_863,In_609,In_938);
nor U864 (N_864,In_933,In_145);
nor U865 (N_865,In_941,In_934);
nor U866 (N_866,In_1216,In_561);
and U867 (N_867,In_1159,In_1346);
and U868 (N_868,In_1468,In_1493);
and U869 (N_869,In_1243,In_1192);
or U870 (N_870,In_1485,In_201);
and U871 (N_871,In_556,In_1126);
and U872 (N_872,In_1138,In_1441);
nand U873 (N_873,In_1129,In_1361);
nand U874 (N_874,In_599,In_1147);
or U875 (N_875,In_1253,In_1470);
or U876 (N_876,In_412,In_935);
xnor U877 (N_877,In_356,In_564);
nor U878 (N_878,In_700,In_1277);
and U879 (N_879,In_1416,In_746);
or U880 (N_880,In_1267,In_453);
and U881 (N_881,In_801,In_1322);
nand U882 (N_882,In_1427,In_434);
nor U883 (N_883,In_1093,In_1337);
nand U884 (N_884,In_584,In_269);
nor U885 (N_885,In_958,In_508);
nand U886 (N_886,In_1020,In_135);
and U887 (N_887,In_418,In_594);
nand U888 (N_888,In_82,In_1433);
and U889 (N_889,In_1281,In_640);
nand U890 (N_890,In_274,In_270);
nand U891 (N_891,In_1381,In_303);
or U892 (N_892,In_347,In_378);
nor U893 (N_893,In_119,In_1424);
or U894 (N_894,In_375,In_1301);
nor U895 (N_895,In_943,In_1227);
nand U896 (N_896,In_572,In_1200);
nor U897 (N_897,In_25,In_1399);
nand U898 (N_898,In_1369,In_972);
nor U899 (N_899,In_878,In_1445);
or U900 (N_900,In_538,In_648);
nand U901 (N_901,In_1470,In_531);
nand U902 (N_902,In_775,In_1336);
or U903 (N_903,In_1027,In_969);
or U904 (N_904,In_238,In_32);
and U905 (N_905,In_95,In_131);
nand U906 (N_906,In_446,In_1342);
or U907 (N_907,In_534,In_42);
nand U908 (N_908,In_326,In_788);
nor U909 (N_909,In_1469,In_165);
and U910 (N_910,In_713,In_853);
or U911 (N_911,In_90,In_1314);
nand U912 (N_912,In_378,In_7);
nor U913 (N_913,In_1499,In_481);
or U914 (N_914,In_1288,In_1374);
nand U915 (N_915,In_572,In_916);
nand U916 (N_916,In_514,In_228);
or U917 (N_917,In_1336,In_428);
and U918 (N_918,In_779,In_1245);
or U919 (N_919,In_418,In_407);
and U920 (N_920,In_855,In_1322);
or U921 (N_921,In_479,In_967);
or U922 (N_922,In_777,In_248);
and U923 (N_923,In_1427,In_1009);
nand U924 (N_924,In_709,In_584);
or U925 (N_925,In_641,In_554);
nand U926 (N_926,In_453,In_234);
nor U927 (N_927,In_1267,In_564);
nand U928 (N_928,In_127,In_1027);
nand U929 (N_929,In_1360,In_1021);
nand U930 (N_930,In_1399,In_1024);
xnor U931 (N_931,In_794,In_1281);
or U932 (N_932,In_674,In_207);
or U933 (N_933,In_762,In_143);
xor U934 (N_934,In_1308,In_207);
and U935 (N_935,In_772,In_83);
and U936 (N_936,In_1371,In_846);
nor U937 (N_937,In_1485,In_67);
and U938 (N_938,In_909,In_953);
or U939 (N_939,In_952,In_113);
and U940 (N_940,In_1113,In_1455);
and U941 (N_941,In_963,In_525);
nand U942 (N_942,In_1338,In_1368);
and U943 (N_943,In_162,In_1156);
and U944 (N_944,In_1080,In_946);
or U945 (N_945,In_736,In_916);
and U946 (N_946,In_482,In_537);
and U947 (N_947,In_603,In_1060);
and U948 (N_948,In_1358,In_59);
and U949 (N_949,In_915,In_564);
nand U950 (N_950,In_143,In_1010);
nand U951 (N_951,In_1063,In_5);
and U952 (N_952,In_872,In_935);
nor U953 (N_953,In_13,In_789);
nor U954 (N_954,In_780,In_1242);
nor U955 (N_955,In_594,In_390);
and U956 (N_956,In_440,In_886);
nand U957 (N_957,In_767,In_865);
and U958 (N_958,In_603,In_431);
nand U959 (N_959,In_1299,In_1482);
nand U960 (N_960,In_1421,In_205);
or U961 (N_961,In_122,In_412);
or U962 (N_962,In_510,In_156);
nor U963 (N_963,In_119,In_666);
nor U964 (N_964,In_1021,In_1079);
nor U965 (N_965,In_125,In_1256);
and U966 (N_966,In_500,In_21);
nor U967 (N_967,In_65,In_145);
xnor U968 (N_968,In_991,In_678);
and U969 (N_969,In_13,In_1410);
xor U970 (N_970,In_371,In_280);
nor U971 (N_971,In_1081,In_1190);
nor U972 (N_972,In_1214,In_711);
nor U973 (N_973,In_1344,In_114);
nor U974 (N_974,In_1428,In_520);
nand U975 (N_975,In_1340,In_694);
nand U976 (N_976,In_346,In_19);
nand U977 (N_977,In_959,In_849);
nor U978 (N_978,In_1441,In_398);
or U979 (N_979,In_474,In_1454);
and U980 (N_980,In_217,In_356);
nor U981 (N_981,In_1357,In_1146);
nand U982 (N_982,In_542,In_490);
nor U983 (N_983,In_1235,In_1200);
nand U984 (N_984,In_1399,In_1248);
xor U985 (N_985,In_980,In_1325);
or U986 (N_986,In_776,In_367);
or U987 (N_987,In_780,In_758);
and U988 (N_988,In_608,In_1222);
nand U989 (N_989,In_196,In_237);
nand U990 (N_990,In_1106,In_1492);
xor U991 (N_991,In_956,In_1101);
nand U992 (N_992,In_203,In_420);
nor U993 (N_993,In_561,In_715);
xnor U994 (N_994,In_491,In_920);
and U995 (N_995,In_367,In_122);
and U996 (N_996,In_1069,In_795);
or U997 (N_997,In_231,In_566);
nand U998 (N_998,In_519,In_1466);
nor U999 (N_999,In_290,In_760);
and U1000 (N_1000,In_60,In_999);
xor U1001 (N_1001,In_1445,In_1347);
and U1002 (N_1002,In_853,In_1467);
or U1003 (N_1003,In_245,In_1276);
and U1004 (N_1004,In_840,In_695);
nand U1005 (N_1005,In_761,In_1053);
nand U1006 (N_1006,In_401,In_325);
nor U1007 (N_1007,In_1234,In_1164);
and U1008 (N_1008,In_452,In_899);
nand U1009 (N_1009,In_1393,In_1013);
or U1010 (N_1010,In_240,In_32);
xnor U1011 (N_1011,In_448,In_1442);
and U1012 (N_1012,In_1200,In_701);
nand U1013 (N_1013,In_951,In_454);
and U1014 (N_1014,In_229,In_29);
nor U1015 (N_1015,In_1287,In_692);
nand U1016 (N_1016,In_1484,In_1245);
and U1017 (N_1017,In_1293,In_615);
nand U1018 (N_1018,In_352,In_164);
nand U1019 (N_1019,In_254,In_619);
xnor U1020 (N_1020,In_939,In_277);
xnor U1021 (N_1021,In_664,In_707);
nand U1022 (N_1022,In_750,In_28);
or U1023 (N_1023,In_133,In_1270);
or U1024 (N_1024,In_1473,In_557);
xnor U1025 (N_1025,In_1260,In_943);
and U1026 (N_1026,In_196,In_692);
nor U1027 (N_1027,In_1145,In_796);
nor U1028 (N_1028,In_284,In_8);
or U1029 (N_1029,In_939,In_545);
nor U1030 (N_1030,In_1438,In_720);
and U1031 (N_1031,In_1362,In_327);
nand U1032 (N_1032,In_1085,In_384);
nand U1033 (N_1033,In_1267,In_1229);
or U1034 (N_1034,In_212,In_1486);
nand U1035 (N_1035,In_644,In_868);
and U1036 (N_1036,In_1185,In_470);
or U1037 (N_1037,In_430,In_1125);
nor U1038 (N_1038,In_708,In_273);
nor U1039 (N_1039,In_324,In_282);
nor U1040 (N_1040,In_130,In_1335);
nor U1041 (N_1041,In_184,In_751);
nor U1042 (N_1042,In_1255,In_1294);
nor U1043 (N_1043,In_26,In_60);
nand U1044 (N_1044,In_1048,In_1166);
or U1045 (N_1045,In_825,In_934);
and U1046 (N_1046,In_51,In_1126);
nor U1047 (N_1047,In_702,In_761);
and U1048 (N_1048,In_664,In_1331);
or U1049 (N_1049,In_934,In_787);
nand U1050 (N_1050,In_814,In_101);
xnor U1051 (N_1051,In_914,In_1049);
or U1052 (N_1052,In_811,In_184);
nor U1053 (N_1053,In_799,In_1071);
or U1054 (N_1054,In_4,In_799);
nand U1055 (N_1055,In_1380,In_1268);
or U1056 (N_1056,In_200,In_1388);
and U1057 (N_1057,In_117,In_1476);
nand U1058 (N_1058,In_1468,In_1254);
and U1059 (N_1059,In_258,In_72);
nor U1060 (N_1060,In_684,In_633);
or U1061 (N_1061,In_767,In_1459);
or U1062 (N_1062,In_1359,In_479);
and U1063 (N_1063,In_240,In_732);
nand U1064 (N_1064,In_54,In_270);
nand U1065 (N_1065,In_846,In_480);
nor U1066 (N_1066,In_167,In_1242);
nor U1067 (N_1067,In_348,In_609);
xnor U1068 (N_1068,In_497,In_531);
and U1069 (N_1069,In_468,In_993);
or U1070 (N_1070,In_987,In_657);
nor U1071 (N_1071,In_1137,In_426);
and U1072 (N_1072,In_1317,In_448);
and U1073 (N_1073,In_1228,In_161);
and U1074 (N_1074,In_911,In_810);
nand U1075 (N_1075,In_128,In_316);
nand U1076 (N_1076,In_1220,In_1151);
nand U1077 (N_1077,In_1215,In_995);
nor U1078 (N_1078,In_123,In_322);
or U1079 (N_1079,In_1310,In_711);
nand U1080 (N_1080,In_1126,In_650);
nand U1081 (N_1081,In_1047,In_355);
nand U1082 (N_1082,In_140,In_149);
xor U1083 (N_1083,In_404,In_1000);
nor U1084 (N_1084,In_66,In_1192);
nor U1085 (N_1085,In_509,In_1106);
nor U1086 (N_1086,In_767,In_1238);
and U1087 (N_1087,In_536,In_769);
nand U1088 (N_1088,In_705,In_1480);
and U1089 (N_1089,In_680,In_788);
nor U1090 (N_1090,In_411,In_1090);
nor U1091 (N_1091,In_133,In_927);
or U1092 (N_1092,In_1111,In_748);
or U1093 (N_1093,In_1276,In_939);
or U1094 (N_1094,In_325,In_264);
or U1095 (N_1095,In_1054,In_1388);
nor U1096 (N_1096,In_1008,In_1447);
nor U1097 (N_1097,In_195,In_637);
or U1098 (N_1098,In_280,In_1324);
and U1099 (N_1099,In_1265,In_621);
or U1100 (N_1100,In_1054,In_1278);
and U1101 (N_1101,In_173,In_1351);
nand U1102 (N_1102,In_1178,In_205);
or U1103 (N_1103,In_660,In_1066);
xor U1104 (N_1104,In_939,In_913);
nand U1105 (N_1105,In_1387,In_30);
nand U1106 (N_1106,In_204,In_1488);
or U1107 (N_1107,In_386,In_285);
or U1108 (N_1108,In_906,In_446);
nor U1109 (N_1109,In_653,In_37);
xnor U1110 (N_1110,In_1014,In_731);
and U1111 (N_1111,In_1110,In_1193);
nand U1112 (N_1112,In_1338,In_0);
nor U1113 (N_1113,In_1319,In_1041);
nor U1114 (N_1114,In_84,In_267);
and U1115 (N_1115,In_293,In_1411);
and U1116 (N_1116,In_773,In_794);
nor U1117 (N_1117,In_597,In_243);
and U1118 (N_1118,In_859,In_22);
nand U1119 (N_1119,In_1198,In_1050);
and U1120 (N_1120,In_205,In_851);
and U1121 (N_1121,In_559,In_13);
and U1122 (N_1122,In_537,In_204);
nand U1123 (N_1123,In_148,In_697);
nor U1124 (N_1124,In_840,In_999);
nor U1125 (N_1125,In_287,In_1237);
nor U1126 (N_1126,In_751,In_1376);
nor U1127 (N_1127,In_1085,In_114);
nand U1128 (N_1128,In_543,In_964);
nand U1129 (N_1129,In_263,In_540);
and U1130 (N_1130,In_274,In_496);
nand U1131 (N_1131,In_1465,In_994);
xnor U1132 (N_1132,In_1121,In_992);
nor U1133 (N_1133,In_919,In_163);
or U1134 (N_1134,In_1129,In_160);
and U1135 (N_1135,In_601,In_700);
nor U1136 (N_1136,In_1295,In_978);
nand U1137 (N_1137,In_975,In_83);
and U1138 (N_1138,In_255,In_679);
or U1139 (N_1139,In_462,In_204);
xor U1140 (N_1140,In_1077,In_792);
or U1141 (N_1141,In_25,In_1339);
or U1142 (N_1142,In_281,In_835);
nor U1143 (N_1143,In_790,In_149);
nand U1144 (N_1144,In_157,In_302);
and U1145 (N_1145,In_478,In_115);
nand U1146 (N_1146,In_1015,In_830);
or U1147 (N_1147,In_686,In_1037);
nor U1148 (N_1148,In_1398,In_321);
or U1149 (N_1149,In_222,In_1483);
or U1150 (N_1150,In_453,In_1439);
and U1151 (N_1151,In_884,In_1417);
nand U1152 (N_1152,In_1015,In_19);
or U1153 (N_1153,In_547,In_201);
nand U1154 (N_1154,In_517,In_600);
or U1155 (N_1155,In_451,In_514);
and U1156 (N_1156,In_360,In_988);
or U1157 (N_1157,In_662,In_540);
nor U1158 (N_1158,In_1432,In_1010);
or U1159 (N_1159,In_847,In_463);
and U1160 (N_1160,In_971,In_1161);
or U1161 (N_1161,In_1182,In_630);
nand U1162 (N_1162,In_187,In_1252);
or U1163 (N_1163,In_907,In_506);
nand U1164 (N_1164,In_1477,In_1239);
or U1165 (N_1165,In_408,In_651);
nor U1166 (N_1166,In_174,In_891);
nor U1167 (N_1167,In_887,In_803);
nand U1168 (N_1168,In_1445,In_77);
xor U1169 (N_1169,In_494,In_1040);
nor U1170 (N_1170,In_479,In_543);
xor U1171 (N_1171,In_661,In_946);
nand U1172 (N_1172,In_592,In_780);
nor U1173 (N_1173,In_673,In_725);
xor U1174 (N_1174,In_64,In_918);
nand U1175 (N_1175,In_261,In_702);
and U1176 (N_1176,In_482,In_1088);
and U1177 (N_1177,In_1253,In_1434);
nand U1178 (N_1178,In_92,In_141);
nand U1179 (N_1179,In_1454,In_833);
and U1180 (N_1180,In_529,In_369);
nor U1181 (N_1181,In_1276,In_806);
or U1182 (N_1182,In_1074,In_1125);
and U1183 (N_1183,In_6,In_724);
nor U1184 (N_1184,In_1012,In_1114);
and U1185 (N_1185,In_500,In_36);
nor U1186 (N_1186,In_713,In_1153);
and U1187 (N_1187,In_160,In_1264);
nand U1188 (N_1188,In_771,In_552);
xnor U1189 (N_1189,In_275,In_245);
xor U1190 (N_1190,In_672,In_998);
or U1191 (N_1191,In_75,In_943);
or U1192 (N_1192,In_1064,In_4);
and U1193 (N_1193,In_697,In_1051);
and U1194 (N_1194,In_1125,In_217);
or U1195 (N_1195,In_898,In_1282);
xor U1196 (N_1196,In_671,In_539);
or U1197 (N_1197,In_698,In_1222);
and U1198 (N_1198,In_1146,In_1091);
and U1199 (N_1199,In_700,In_19);
nand U1200 (N_1200,In_301,In_1014);
or U1201 (N_1201,In_824,In_560);
nor U1202 (N_1202,In_1123,In_486);
xnor U1203 (N_1203,In_1186,In_241);
or U1204 (N_1204,In_826,In_958);
xor U1205 (N_1205,In_5,In_447);
and U1206 (N_1206,In_802,In_474);
xor U1207 (N_1207,In_346,In_935);
and U1208 (N_1208,In_151,In_1349);
nand U1209 (N_1209,In_1364,In_1470);
nand U1210 (N_1210,In_1407,In_86);
nor U1211 (N_1211,In_759,In_1409);
nand U1212 (N_1212,In_420,In_627);
and U1213 (N_1213,In_1063,In_1327);
nand U1214 (N_1214,In_1357,In_90);
nand U1215 (N_1215,In_456,In_424);
nor U1216 (N_1216,In_340,In_83);
nor U1217 (N_1217,In_1264,In_680);
or U1218 (N_1218,In_1305,In_482);
nand U1219 (N_1219,In_1100,In_1196);
and U1220 (N_1220,In_1048,In_158);
and U1221 (N_1221,In_1075,In_562);
and U1222 (N_1222,In_62,In_1064);
or U1223 (N_1223,In_1430,In_221);
nor U1224 (N_1224,In_33,In_385);
nand U1225 (N_1225,In_648,In_557);
and U1226 (N_1226,In_715,In_756);
or U1227 (N_1227,In_810,In_914);
and U1228 (N_1228,In_118,In_775);
nor U1229 (N_1229,In_1329,In_169);
and U1230 (N_1230,In_916,In_589);
or U1231 (N_1231,In_960,In_584);
nand U1232 (N_1232,In_1122,In_809);
nor U1233 (N_1233,In_515,In_407);
nor U1234 (N_1234,In_329,In_883);
or U1235 (N_1235,In_880,In_641);
nand U1236 (N_1236,In_1319,In_1254);
or U1237 (N_1237,In_363,In_1447);
nand U1238 (N_1238,In_269,In_1408);
nor U1239 (N_1239,In_1022,In_395);
nor U1240 (N_1240,In_1182,In_975);
nor U1241 (N_1241,In_267,In_1107);
and U1242 (N_1242,In_707,In_1273);
nor U1243 (N_1243,In_58,In_574);
nand U1244 (N_1244,In_307,In_462);
or U1245 (N_1245,In_1278,In_1001);
nand U1246 (N_1246,In_108,In_20);
nor U1247 (N_1247,In_1151,In_833);
nor U1248 (N_1248,In_664,In_690);
nor U1249 (N_1249,In_162,In_566);
or U1250 (N_1250,In_879,In_685);
and U1251 (N_1251,In_1122,In_1177);
and U1252 (N_1252,In_1359,In_878);
and U1253 (N_1253,In_137,In_1296);
and U1254 (N_1254,In_1020,In_1455);
and U1255 (N_1255,In_895,In_883);
xor U1256 (N_1256,In_1162,In_186);
or U1257 (N_1257,In_881,In_715);
or U1258 (N_1258,In_1464,In_115);
and U1259 (N_1259,In_749,In_646);
and U1260 (N_1260,In_755,In_171);
nand U1261 (N_1261,In_1414,In_64);
nor U1262 (N_1262,In_580,In_307);
or U1263 (N_1263,In_970,In_163);
or U1264 (N_1264,In_709,In_1350);
nor U1265 (N_1265,In_464,In_1246);
nand U1266 (N_1266,In_191,In_354);
and U1267 (N_1267,In_1417,In_4);
or U1268 (N_1268,In_742,In_963);
and U1269 (N_1269,In_926,In_430);
nor U1270 (N_1270,In_1038,In_100);
nor U1271 (N_1271,In_988,In_342);
nand U1272 (N_1272,In_327,In_497);
or U1273 (N_1273,In_465,In_1350);
and U1274 (N_1274,In_390,In_46);
xnor U1275 (N_1275,In_722,In_238);
nand U1276 (N_1276,In_1097,In_878);
or U1277 (N_1277,In_304,In_1493);
and U1278 (N_1278,In_536,In_1026);
nor U1279 (N_1279,In_67,In_404);
nand U1280 (N_1280,In_1476,In_498);
or U1281 (N_1281,In_1161,In_1236);
and U1282 (N_1282,In_681,In_641);
nand U1283 (N_1283,In_901,In_144);
nor U1284 (N_1284,In_1413,In_1482);
and U1285 (N_1285,In_182,In_1357);
or U1286 (N_1286,In_1082,In_309);
nand U1287 (N_1287,In_241,In_1474);
and U1288 (N_1288,In_802,In_34);
or U1289 (N_1289,In_463,In_1067);
nor U1290 (N_1290,In_381,In_1162);
nand U1291 (N_1291,In_1267,In_1219);
and U1292 (N_1292,In_885,In_609);
nor U1293 (N_1293,In_1297,In_370);
and U1294 (N_1294,In_429,In_519);
or U1295 (N_1295,In_413,In_468);
nand U1296 (N_1296,In_1293,In_970);
and U1297 (N_1297,In_449,In_1370);
nand U1298 (N_1298,In_944,In_714);
and U1299 (N_1299,In_66,In_1187);
or U1300 (N_1300,In_1441,In_1403);
or U1301 (N_1301,In_44,In_84);
and U1302 (N_1302,In_868,In_354);
and U1303 (N_1303,In_1061,In_6);
nand U1304 (N_1304,In_1214,In_1124);
nor U1305 (N_1305,In_859,In_832);
and U1306 (N_1306,In_551,In_490);
nand U1307 (N_1307,In_1029,In_935);
or U1308 (N_1308,In_856,In_12);
or U1309 (N_1309,In_1327,In_369);
nor U1310 (N_1310,In_1488,In_1071);
nor U1311 (N_1311,In_1316,In_455);
and U1312 (N_1312,In_624,In_664);
or U1313 (N_1313,In_1468,In_186);
and U1314 (N_1314,In_840,In_1178);
or U1315 (N_1315,In_207,In_80);
nand U1316 (N_1316,In_795,In_1328);
nor U1317 (N_1317,In_886,In_842);
or U1318 (N_1318,In_1,In_306);
or U1319 (N_1319,In_1044,In_814);
nand U1320 (N_1320,In_1063,In_1289);
and U1321 (N_1321,In_1284,In_890);
nand U1322 (N_1322,In_597,In_1230);
nor U1323 (N_1323,In_1124,In_1133);
and U1324 (N_1324,In_128,In_8);
xor U1325 (N_1325,In_482,In_989);
or U1326 (N_1326,In_183,In_456);
or U1327 (N_1327,In_136,In_1146);
nand U1328 (N_1328,In_628,In_152);
nand U1329 (N_1329,In_308,In_1326);
nand U1330 (N_1330,In_1413,In_780);
and U1331 (N_1331,In_1129,In_1412);
or U1332 (N_1332,In_912,In_1093);
nor U1333 (N_1333,In_850,In_680);
nand U1334 (N_1334,In_261,In_1177);
nand U1335 (N_1335,In_682,In_35);
nand U1336 (N_1336,In_1030,In_1225);
nor U1337 (N_1337,In_380,In_763);
or U1338 (N_1338,In_2,In_376);
and U1339 (N_1339,In_331,In_399);
nand U1340 (N_1340,In_447,In_1374);
nand U1341 (N_1341,In_971,In_562);
or U1342 (N_1342,In_707,In_538);
and U1343 (N_1343,In_689,In_54);
and U1344 (N_1344,In_1135,In_1158);
xor U1345 (N_1345,In_698,In_599);
and U1346 (N_1346,In_1004,In_1087);
xnor U1347 (N_1347,In_287,In_1013);
or U1348 (N_1348,In_864,In_481);
or U1349 (N_1349,In_1142,In_156);
or U1350 (N_1350,In_73,In_9);
or U1351 (N_1351,In_1375,In_271);
nand U1352 (N_1352,In_1487,In_101);
and U1353 (N_1353,In_1109,In_1240);
or U1354 (N_1354,In_1366,In_933);
nand U1355 (N_1355,In_147,In_112);
or U1356 (N_1356,In_572,In_1420);
xnor U1357 (N_1357,In_418,In_367);
nand U1358 (N_1358,In_1141,In_311);
nand U1359 (N_1359,In_1313,In_1478);
or U1360 (N_1360,In_490,In_23);
nor U1361 (N_1361,In_902,In_488);
xor U1362 (N_1362,In_1050,In_115);
nor U1363 (N_1363,In_1028,In_214);
nand U1364 (N_1364,In_530,In_746);
xor U1365 (N_1365,In_896,In_464);
and U1366 (N_1366,In_1440,In_1124);
nor U1367 (N_1367,In_1172,In_1139);
and U1368 (N_1368,In_1103,In_321);
and U1369 (N_1369,In_1346,In_702);
or U1370 (N_1370,In_1218,In_1419);
nand U1371 (N_1371,In_965,In_1132);
or U1372 (N_1372,In_1035,In_554);
nand U1373 (N_1373,In_628,In_1288);
and U1374 (N_1374,In_581,In_711);
and U1375 (N_1375,In_808,In_1345);
nor U1376 (N_1376,In_945,In_1332);
xor U1377 (N_1377,In_469,In_394);
nand U1378 (N_1378,In_98,In_9);
and U1379 (N_1379,In_888,In_1016);
or U1380 (N_1380,In_677,In_986);
or U1381 (N_1381,In_1331,In_1398);
nand U1382 (N_1382,In_1391,In_730);
and U1383 (N_1383,In_10,In_1153);
nor U1384 (N_1384,In_552,In_912);
nor U1385 (N_1385,In_556,In_1236);
or U1386 (N_1386,In_280,In_1026);
nand U1387 (N_1387,In_1184,In_842);
nor U1388 (N_1388,In_1124,In_708);
nor U1389 (N_1389,In_506,In_189);
or U1390 (N_1390,In_980,In_281);
nand U1391 (N_1391,In_1003,In_1186);
or U1392 (N_1392,In_1489,In_556);
and U1393 (N_1393,In_1035,In_929);
or U1394 (N_1394,In_718,In_339);
nor U1395 (N_1395,In_1333,In_470);
or U1396 (N_1396,In_53,In_1126);
nor U1397 (N_1397,In_815,In_309);
nand U1398 (N_1398,In_1443,In_1296);
nor U1399 (N_1399,In_507,In_81);
nand U1400 (N_1400,In_691,In_1421);
and U1401 (N_1401,In_1284,In_414);
and U1402 (N_1402,In_84,In_1011);
nand U1403 (N_1403,In_1342,In_841);
or U1404 (N_1404,In_1185,In_783);
nor U1405 (N_1405,In_1452,In_171);
and U1406 (N_1406,In_1361,In_235);
nor U1407 (N_1407,In_383,In_844);
nand U1408 (N_1408,In_952,In_833);
nand U1409 (N_1409,In_696,In_160);
or U1410 (N_1410,In_78,In_788);
and U1411 (N_1411,In_86,In_434);
and U1412 (N_1412,In_189,In_510);
and U1413 (N_1413,In_1335,In_807);
nand U1414 (N_1414,In_229,In_152);
nand U1415 (N_1415,In_723,In_1286);
and U1416 (N_1416,In_541,In_172);
and U1417 (N_1417,In_155,In_897);
nor U1418 (N_1418,In_300,In_67);
nor U1419 (N_1419,In_1453,In_1494);
and U1420 (N_1420,In_929,In_1220);
nand U1421 (N_1421,In_763,In_567);
nand U1422 (N_1422,In_1272,In_170);
nand U1423 (N_1423,In_70,In_54);
nor U1424 (N_1424,In_508,In_7);
or U1425 (N_1425,In_22,In_1309);
nand U1426 (N_1426,In_300,In_1138);
and U1427 (N_1427,In_713,In_939);
and U1428 (N_1428,In_1230,In_1185);
nor U1429 (N_1429,In_860,In_803);
or U1430 (N_1430,In_298,In_680);
nand U1431 (N_1431,In_170,In_1010);
and U1432 (N_1432,In_122,In_888);
or U1433 (N_1433,In_1066,In_1368);
or U1434 (N_1434,In_1222,In_489);
and U1435 (N_1435,In_235,In_1000);
or U1436 (N_1436,In_1332,In_190);
and U1437 (N_1437,In_1227,In_136);
nor U1438 (N_1438,In_1153,In_621);
nor U1439 (N_1439,In_132,In_176);
nor U1440 (N_1440,In_319,In_814);
nor U1441 (N_1441,In_1366,In_464);
xnor U1442 (N_1442,In_1124,In_786);
xor U1443 (N_1443,In_1169,In_264);
nor U1444 (N_1444,In_1377,In_1253);
nand U1445 (N_1445,In_1330,In_271);
xnor U1446 (N_1446,In_1291,In_460);
nand U1447 (N_1447,In_258,In_648);
nand U1448 (N_1448,In_695,In_810);
nand U1449 (N_1449,In_901,In_1451);
or U1450 (N_1450,In_1034,In_898);
and U1451 (N_1451,In_759,In_125);
or U1452 (N_1452,In_580,In_920);
or U1453 (N_1453,In_1151,In_243);
nor U1454 (N_1454,In_1496,In_1021);
and U1455 (N_1455,In_418,In_1013);
and U1456 (N_1456,In_335,In_600);
and U1457 (N_1457,In_505,In_846);
or U1458 (N_1458,In_989,In_1051);
or U1459 (N_1459,In_988,In_100);
or U1460 (N_1460,In_252,In_1470);
or U1461 (N_1461,In_875,In_1200);
and U1462 (N_1462,In_1107,In_1008);
nand U1463 (N_1463,In_526,In_14);
xor U1464 (N_1464,In_878,In_1462);
nand U1465 (N_1465,In_23,In_1201);
nor U1466 (N_1466,In_1467,In_232);
or U1467 (N_1467,In_1402,In_1297);
or U1468 (N_1468,In_862,In_1232);
and U1469 (N_1469,In_447,In_1013);
nand U1470 (N_1470,In_1180,In_368);
nand U1471 (N_1471,In_1428,In_311);
xnor U1472 (N_1472,In_273,In_1071);
nand U1473 (N_1473,In_1080,In_903);
nand U1474 (N_1474,In_636,In_156);
nor U1475 (N_1475,In_1459,In_839);
xnor U1476 (N_1476,In_919,In_35);
or U1477 (N_1477,In_1133,In_310);
nor U1478 (N_1478,In_155,In_435);
and U1479 (N_1479,In_571,In_1244);
nand U1480 (N_1480,In_336,In_643);
nand U1481 (N_1481,In_1100,In_1454);
nor U1482 (N_1482,In_140,In_1225);
nand U1483 (N_1483,In_9,In_354);
nand U1484 (N_1484,In_1148,In_121);
nand U1485 (N_1485,In_1487,In_562);
nand U1486 (N_1486,In_1445,In_1429);
and U1487 (N_1487,In_100,In_1349);
nor U1488 (N_1488,In_182,In_1252);
nor U1489 (N_1489,In_474,In_927);
nand U1490 (N_1490,In_118,In_1303);
nand U1491 (N_1491,In_1,In_256);
nand U1492 (N_1492,In_1042,In_832);
xor U1493 (N_1493,In_1338,In_985);
or U1494 (N_1494,In_650,In_906);
or U1495 (N_1495,In_892,In_285);
xnor U1496 (N_1496,In_240,In_497);
or U1497 (N_1497,In_11,In_701);
nor U1498 (N_1498,In_1186,In_209);
nor U1499 (N_1499,In_394,In_1112);
nand U1500 (N_1500,In_244,In_97);
and U1501 (N_1501,In_441,In_646);
nor U1502 (N_1502,In_1007,In_1496);
and U1503 (N_1503,In_793,In_711);
and U1504 (N_1504,In_997,In_261);
nor U1505 (N_1505,In_146,In_262);
nor U1506 (N_1506,In_1370,In_131);
nand U1507 (N_1507,In_166,In_1031);
and U1508 (N_1508,In_1466,In_444);
and U1509 (N_1509,In_564,In_756);
and U1510 (N_1510,In_902,In_555);
and U1511 (N_1511,In_807,In_1373);
and U1512 (N_1512,In_66,In_368);
and U1513 (N_1513,In_1374,In_1241);
and U1514 (N_1514,In_628,In_1379);
or U1515 (N_1515,In_821,In_1271);
nor U1516 (N_1516,In_623,In_772);
or U1517 (N_1517,In_1354,In_1050);
nor U1518 (N_1518,In_264,In_1232);
and U1519 (N_1519,In_477,In_84);
and U1520 (N_1520,In_1302,In_198);
or U1521 (N_1521,In_1006,In_1205);
and U1522 (N_1522,In_1202,In_1395);
or U1523 (N_1523,In_546,In_493);
nand U1524 (N_1524,In_440,In_1062);
nand U1525 (N_1525,In_742,In_453);
and U1526 (N_1526,In_739,In_1085);
nor U1527 (N_1527,In_920,In_533);
nand U1528 (N_1528,In_437,In_415);
nand U1529 (N_1529,In_474,In_23);
xnor U1530 (N_1530,In_1240,In_190);
nand U1531 (N_1531,In_1046,In_878);
nor U1532 (N_1532,In_180,In_583);
or U1533 (N_1533,In_819,In_414);
nor U1534 (N_1534,In_519,In_146);
nand U1535 (N_1535,In_673,In_830);
nand U1536 (N_1536,In_123,In_279);
and U1537 (N_1537,In_178,In_495);
xor U1538 (N_1538,In_903,In_194);
and U1539 (N_1539,In_1067,In_353);
xnor U1540 (N_1540,In_138,In_282);
nor U1541 (N_1541,In_1191,In_668);
and U1542 (N_1542,In_1226,In_985);
and U1543 (N_1543,In_603,In_1431);
and U1544 (N_1544,In_1352,In_1285);
or U1545 (N_1545,In_1022,In_116);
nor U1546 (N_1546,In_17,In_648);
nand U1547 (N_1547,In_1036,In_874);
or U1548 (N_1548,In_1140,In_1494);
nor U1549 (N_1549,In_1404,In_255);
nand U1550 (N_1550,In_133,In_297);
and U1551 (N_1551,In_153,In_919);
nor U1552 (N_1552,In_1311,In_1090);
or U1553 (N_1553,In_895,In_958);
and U1554 (N_1554,In_102,In_697);
or U1555 (N_1555,In_634,In_1466);
and U1556 (N_1556,In_1117,In_1216);
nand U1557 (N_1557,In_522,In_622);
and U1558 (N_1558,In_539,In_1269);
nand U1559 (N_1559,In_316,In_273);
xnor U1560 (N_1560,In_46,In_170);
xnor U1561 (N_1561,In_1254,In_1292);
nor U1562 (N_1562,In_442,In_679);
nand U1563 (N_1563,In_1445,In_1110);
nand U1564 (N_1564,In_815,In_646);
or U1565 (N_1565,In_1360,In_613);
and U1566 (N_1566,In_195,In_712);
or U1567 (N_1567,In_326,In_789);
nand U1568 (N_1568,In_958,In_930);
and U1569 (N_1569,In_1427,In_133);
or U1570 (N_1570,In_297,In_1040);
xnor U1571 (N_1571,In_1175,In_148);
nor U1572 (N_1572,In_964,In_1130);
nand U1573 (N_1573,In_1127,In_889);
or U1574 (N_1574,In_554,In_399);
or U1575 (N_1575,In_46,In_254);
or U1576 (N_1576,In_217,In_1064);
or U1577 (N_1577,In_774,In_767);
nand U1578 (N_1578,In_1181,In_1333);
and U1579 (N_1579,In_895,In_1138);
nand U1580 (N_1580,In_52,In_917);
nor U1581 (N_1581,In_1215,In_250);
nand U1582 (N_1582,In_417,In_1055);
nand U1583 (N_1583,In_1385,In_245);
nor U1584 (N_1584,In_230,In_779);
nand U1585 (N_1585,In_1015,In_597);
or U1586 (N_1586,In_340,In_667);
nor U1587 (N_1587,In_1069,In_1423);
and U1588 (N_1588,In_1016,In_1161);
nand U1589 (N_1589,In_998,In_639);
xor U1590 (N_1590,In_417,In_1061);
or U1591 (N_1591,In_886,In_736);
or U1592 (N_1592,In_720,In_61);
nor U1593 (N_1593,In_1199,In_532);
and U1594 (N_1594,In_306,In_388);
nor U1595 (N_1595,In_1410,In_1329);
or U1596 (N_1596,In_241,In_220);
or U1597 (N_1597,In_730,In_1376);
nor U1598 (N_1598,In_1197,In_764);
nor U1599 (N_1599,In_740,In_1212);
nor U1600 (N_1600,In_1043,In_193);
and U1601 (N_1601,In_1035,In_1431);
nor U1602 (N_1602,In_904,In_1239);
and U1603 (N_1603,In_1315,In_873);
xor U1604 (N_1604,In_507,In_1041);
nor U1605 (N_1605,In_814,In_1374);
and U1606 (N_1606,In_922,In_1056);
nor U1607 (N_1607,In_976,In_84);
nand U1608 (N_1608,In_1329,In_774);
nand U1609 (N_1609,In_261,In_1070);
or U1610 (N_1610,In_655,In_709);
and U1611 (N_1611,In_1411,In_1466);
xnor U1612 (N_1612,In_342,In_1000);
and U1613 (N_1613,In_275,In_827);
or U1614 (N_1614,In_1010,In_774);
or U1615 (N_1615,In_752,In_824);
and U1616 (N_1616,In_1471,In_74);
nand U1617 (N_1617,In_778,In_1490);
or U1618 (N_1618,In_1279,In_997);
nand U1619 (N_1619,In_738,In_62);
nor U1620 (N_1620,In_1225,In_964);
or U1621 (N_1621,In_693,In_1203);
or U1622 (N_1622,In_510,In_237);
nor U1623 (N_1623,In_1168,In_1436);
or U1624 (N_1624,In_138,In_513);
xor U1625 (N_1625,In_405,In_1254);
nor U1626 (N_1626,In_200,In_1143);
and U1627 (N_1627,In_489,In_451);
or U1628 (N_1628,In_1064,In_29);
or U1629 (N_1629,In_957,In_571);
nor U1630 (N_1630,In_924,In_348);
or U1631 (N_1631,In_810,In_669);
nand U1632 (N_1632,In_666,In_820);
xor U1633 (N_1633,In_963,In_578);
nor U1634 (N_1634,In_311,In_123);
and U1635 (N_1635,In_1021,In_226);
or U1636 (N_1636,In_282,In_1162);
nand U1637 (N_1637,In_401,In_670);
nand U1638 (N_1638,In_1302,In_1123);
or U1639 (N_1639,In_1416,In_167);
nor U1640 (N_1640,In_975,In_553);
nor U1641 (N_1641,In_664,In_682);
nor U1642 (N_1642,In_1267,In_1409);
or U1643 (N_1643,In_1064,In_150);
nor U1644 (N_1644,In_862,In_311);
and U1645 (N_1645,In_1420,In_365);
nand U1646 (N_1646,In_1241,In_733);
nand U1647 (N_1647,In_231,In_857);
nand U1648 (N_1648,In_1387,In_759);
and U1649 (N_1649,In_1447,In_690);
nand U1650 (N_1650,In_908,In_1054);
and U1651 (N_1651,In_329,In_1482);
nand U1652 (N_1652,In_17,In_1185);
and U1653 (N_1653,In_169,In_845);
nand U1654 (N_1654,In_1295,In_185);
or U1655 (N_1655,In_1457,In_1203);
or U1656 (N_1656,In_40,In_899);
and U1657 (N_1657,In_1105,In_59);
nand U1658 (N_1658,In_661,In_1186);
nand U1659 (N_1659,In_1222,In_509);
and U1660 (N_1660,In_664,In_955);
and U1661 (N_1661,In_43,In_987);
or U1662 (N_1662,In_1274,In_623);
nor U1663 (N_1663,In_287,In_1448);
or U1664 (N_1664,In_808,In_1417);
and U1665 (N_1665,In_871,In_1358);
nor U1666 (N_1666,In_1422,In_1210);
and U1667 (N_1667,In_251,In_1110);
or U1668 (N_1668,In_1378,In_1202);
nor U1669 (N_1669,In_992,In_173);
nor U1670 (N_1670,In_1306,In_1488);
nor U1671 (N_1671,In_1133,In_616);
and U1672 (N_1672,In_75,In_157);
nand U1673 (N_1673,In_289,In_133);
or U1674 (N_1674,In_1269,In_740);
or U1675 (N_1675,In_252,In_765);
or U1676 (N_1676,In_528,In_1457);
nor U1677 (N_1677,In_1089,In_1350);
nand U1678 (N_1678,In_186,In_480);
and U1679 (N_1679,In_563,In_1332);
or U1680 (N_1680,In_1225,In_1074);
or U1681 (N_1681,In_414,In_506);
or U1682 (N_1682,In_671,In_885);
nor U1683 (N_1683,In_570,In_885);
or U1684 (N_1684,In_1178,In_119);
nand U1685 (N_1685,In_1002,In_456);
and U1686 (N_1686,In_704,In_1474);
nor U1687 (N_1687,In_275,In_1072);
nand U1688 (N_1688,In_1203,In_210);
and U1689 (N_1689,In_1003,In_369);
and U1690 (N_1690,In_1061,In_615);
nand U1691 (N_1691,In_1439,In_653);
and U1692 (N_1692,In_101,In_1099);
nor U1693 (N_1693,In_884,In_1149);
and U1694 (N_1694,In_220,In_303);
and U1695 (N_1695,In_469,In_1436);
or U1696 (N_1696,In_886,In_93);
or U1697 (N_1697,In_925,In_1487);
nor U1698 (N_1698,In_533,In_13);
xnor U1699 (N_1699,In_451,In_563);
or U1700 (N_1700,In_815,In_257);
or U1701 (N_1701,In_985,In_1211);
nor U1702 (N_1702,In_703,In_1190);
and U1703 (N_1703,In_376,In_139);
nor U1704 (N_1704,In_534,In_176);
or U1705 (N_1705,In_216,In_1034);
and U1706 (N_1706,In_35,In_1204);
nand U1707 (N_1707,In_1494,In_1132);
or U1708 (N_1708,In_561,In_1297);
nand U1709 (N_1709,In_496,In_818);
nor U1710 (N_1710,In_1494,In_1255);
nor U1711 (N_1711,In_1030,In_1029);
and U1712 (N_1712,In_174,In_599);
or U1713 (N_1713,In_672,In_1269);
nand U1714 (N_1714,In_1374,In_466);
and U1715 (N_1715,In_112,In_386);
nand U1716 (N_1716,In_957,In_280);
nand U1717 (N_1717,In_120,In_1490);
nand U1718 (N_1718,In_162,In_765);
xor U1719 (N_1719,In_422,In_29);
nand U1720 (N_1720,In_820,In_1423);
xor U1721 (N_1721,In_429,In_1255);
or U1722 (N_1722,In_763,In_1226);
or U1723 (N_1723,In_604,In_1132);
nor U1724 (N_1724,In_456,In_1036);
nand U1725 (N_1725,In_605,In_130);
nor U1726 (N_1726,In_1116,In_1415);
nand U1727 (N_1727,In_1391,In_204);
and U1728 (N_1728,In_1010,In_570);
nor U1729 (N_1729,In_1319,In_951);
or U1730 (N_1730,In_1367,In_692);
nor U1731 (N_1731,In_858,In_1064);
nand U1732 (N_1732,In_1455,In_554);
nand U1733 (N_1733,In_56,In_721);
nand U1734 (N_1734,In_330,In_1223);
and U1735 (N_1735,In_737,In_270);
nor U1736 (N_1736,In_1419,In_327);
nor U1737 (N_1737,In_801,In_1307);
and U1738 (N_1738,In_280,In_1369);
nand U1739 (N_1739,In_318,In_471);
xnor U1740 (N_1740,In_40,In_30);
xnor U1741 (N_1741,In_73,In_1414);
or U1742 (N_1742,In_242,In_587);
or U1743 (N_1743,In_739,In_129);
nor U1744 (N_1744,In_1430,In_1468);
and U1745 (N_1745,In_759,In_334);
nor U1746 (N_1746,In_1164,In_1250);
nor U1747 (N_1747,In_551,In_1493);
nor U1748 (N_1748,In_879,In_247);
or U1749 (N_1749,In_319,In_1135);
nor U1750 (N_1750,In_1033,In_274);
nand U1751 (N_1751,In_1246,In_225);
nor U1752 (N_1752,In_491,In_412);
nand U1753 (N_1753,In_860,In_9);
nand U1754 (N_1754,In_1039,In_818);
or U1755 (N_1755,In_1384,In_927);
and U1756 (N_1756,In_199,In_1155);
or U1757 (N_1757,In_650,In_374);
or U1758 (N_1758,In_52,In_441);
nand U1759 (N_1759,In_774,In_149);
xnor U1760 (N_1760,In_1455,In_143);
xnor U1761 (N_1761,In_1354,In_322);
or U1762 (N_1762,In_1233,In_1334);
or U1763 (N_1763,In_836,In_273);
xnor U1764 (N_1764,In_1050,In_564);
or U1765 (N_1765,In_287,In_1034);
xor U1766 (N_1766,In_1330,In_341);
nor U1767 (N_1767,In_634,In_1397);
nand U1768 (N_1768,In_135,In_1334);
nor U1769 (N_1769,In_167,In_279);
nand U1770 (N_1770,In_391,In_1060);
xnor U1771 (N_1771,In_200,In_1040);
nand U1772 (N_1772,In_365,In_545);
nor U1773 (N_1773,In_345,In_913);
or U1774 (N_1774,In_1301,In_139);
nor U1775 (N_1775,In_398,In_234);
and U1776 (N_1776,In_1129,In_920);
nand U1777 (N_1777,In_269,In_1369);
and U1778 (N_1778,In_1453,In_1369);
nand U1779 (N_1779,In_604,In_613);
and U1780 (N_1780,In_355,In_690);
and U1781 (N_1781,In_434,In_717);
and U1782 (N_1782,In_508,In_662);
nor U1783 (N_1783,In_455,In_1152);
and U1784 (N_1784,In_235,In_597);
or U1785 (N_1785,In_1007,In_1030);
or U1786 (N_1786,In_389,In_124);
nand U1787 (N_1787,In_1169,In_1304);
or U1788 (N_1788,In_123,In_304);
or U1789 (N_1789,In_1454,In_1347);
nor U1790 (N_1790,In_37,In_630);
nor U1791 (N_1791,In_181,In_1432);
or U1792 (N_1792,In_1301,In_1036);
xnor U1793 (N_1793,In_896,In_650);
or U1794 (N_1794,In_886,In_228);
nor U1795 (N_1795,In_224,In_1473);
and U1796 (N_1796,In_772,In_35);
nand U1797 (N_1797,In_1219,In_869);
and U1798 (N_1798,In_19,In_60);
nor U1799 (N_1799,In_1424,In_399);
xnor U1800 (N_1800,In_1225,In_836);
nand U1801 (N_1801,In_1278,In_737);
nor U1802 (N_1802,In_680,In_297);
nand U1803 (N_1803,In_145,In_204);
and U1804 (N_1804,In_309,In_1395);
or U1805 (N_1805,In_689,In_1384);
and U1806 (N_1806,In_1145,In_1495);
nor U1807 (N_1807,In_62,In_609);
nand U1808 (N_1808,In_762,In_696);
nand U1809 (N_1809,In_659,In_742);
or U1810 (N_1810,In_514,In_699);
nand U1811 (N_1811,In_649,In_850);
and U1812 (N_1812,In_292,In_985);
nor U1813 (N_1813,In_182,In_844);
and U1814 (N_1814,In_1036,In_1379);
nand U1815 (N_1815,In_1021,In_570);
and U1816 (N_1816,In_1338,In_825);
or U1817 (N_1817,In_248,In_870);
xor U1818 (N_1818,In_395,In_1316);
nor U1819 (N_1819,In_354,In_426);
and U1820 (N_1820,In_688,In_1218);
nor U1821 (N_1821,In_127,In_1226);
or U1822 (N_1822,In_1075,In_850);
nor U1823 (N_1823,In_529,In_240);
nand U1824 (N_1824,In_497,In_389);
nor U1825 (N_1825,In_575,In_227);
nand U1826 (N_1826,In_60,In_454);
nand U1827 (N_1827,In_540,In_178);
or U1828 (N_1828,In_91,In_1229);
nand U1829 (N_1829,In_912,In_889);
xnor U1830 (N_1830,In_594,In_261);
or U1831 (N_1831,In_43,In_888);
or U1832 (N_1832,In_287,In_1378);
nor U1833 (N_1833,In_278,In_656);
and U1834 (N_1834,In_747,In_297);
nor U1835 (N_1835,In_67,In_1169);
xnor U1836 (N_1836,In_549,In_152);
nor U1837 (N_1837,In_856,In_444);
nor U1838 (N_1838,In_1267,In_701);
and U1839 (N_1839,In_1471,In_1042);
nor U1840 (N_1840,In_1099,In_1290);
or U1841 (N_1841,In_1408,In_326);
nor U1842 (N_1842,In_1482,In_1464);
nand U1843 (N_1843,In_306,In_1064);
and U1844 (N_1844,In_531,In_1236);
nor U1845 (N_1845,In_812,In_1085);
nor U1846 (N_1846,In_989,In_1316);
nor U1847 (N_1847,In_1151,In_107);
nor U1848 (N_1848,In_68,In_80);
nor U1849 (N_1849,In_1047,In_782);
nor U1850 (N_1850,In_848,In_1405);
and U1851 (N_1851,In_806,In_174);
nand U1852 (N_1852,In_103,In_1221);
and U1853 (N_1853,In_1301,In_386);
and U1854 (N_1854,In_1266,In_1309);
nor U1855 (N_1855,In_475,In_998);
nand U1856 (N_1856,In_32,In_103);
nand U1857 (N_1857,In_1440,In_296);
or U1858 (N_1858,In_405,In_784);
nor U1859 (N_1859,In_136,In_905);
nor U1860 (N_1860,In_650,In_328);
or U1861 (N_1861,In_545,In_497);
nor U1862 (N_1862,In_333,In_1005);
nand U1863 (N_1863,In_373,In_1079);
or U1864 (N_1864,In_116,In_500);
or U1865 (N_1865,In_1397,In_441);
nand U1866 (N_1866,In_543,In_567);
nor U1867 (N_1867,In_993,In_1006);
nand U1868 (N_1868,In_931,In_1039);
or U1869 (N_1869,In_1180,In_85);
or U1870 (N_1870,In_1251,In_942);
nor U1871 (N_1871,In_750,In_1162);
nand U1872 (N_1872,In_1215,In_35);
or U1873 (N_1873,In_711,In_39);
and U1874 (N_1874,In_1446,In_1226);
or U1875 (N_1875,In_621,In_296);
and U1876 (N_1876,In_1189,In_95);
or U1877 (N_1877,In_1474,In_799);
xor U1878 (N_1878,In_1003,In_1017);
nor U1879 (N_1879,In_1396,In_836);
and U1880 (N_1880,In_1035,In_411);
nor U1881 (N_1881,In_173,In_709);
nand U1882 (N_1882,In_643,In_534);
xnor U1883 (N_1883,In_73,In_192);
nor U1884 (N_1884,In_351,In_602);
and U1885 (N_1885,In_84,In_790);
and U1886 (N_1886,In_221,In_1259);
or U1887 (N_1887,In_1413,In_1132);
or U1888 (N_1888,In_126,In_389);
and U1889 (N_1889,In_41,In_1415);
nand U1890 (N_1890,In_1381,In_58);
and U1891 (N_1891,In_65,In_573);
and U1892 (N_1892,In_1191,In_1453);
nand U1893 (N_1893,In_768,In_647);
or U1894 (N_1894,In_1044,In_630);
nand U1895 (N_1895,In_295,In_1146);
nand U1896 (N_1896,In_515,In_1108);
and U1897 (N_1897,In_718,In_341);
nor U1898 (N_1898,In_534,In_391);
nand U1899 (N_1899,In_458,In_1278);
nor U1900 (N_1900,In_766,In_602);
nand U1901 (N_1901,In_914,In_591);
and U1902 (N_1902,In_645,In_1117);
nor U1903 (N_1903,In_655,In_682);
or U1904 (N_1904,In_32,In_713);
or U1905 (N_1905,In_825,In_122);
nor U1906 (N_1906,In_730,In_861);
or U1907 (N_1907,In_735,In_725);
and U1908 (N_1908,In_1462,In_1126);
xor U1909 (N_1909,In_1180,In_1121);
and U1910 (N_1910,In_370,In_227);
and U1911 (N_1911,In_350,In_1195);
nor U1912 (N_1912,In_488,In_627);
and U1913 (N_1913,In_578,In_14);
nor U1914 (N_1914,In_1404,In_844);
or U1915 (N_1915,In_1276,In_117);
nand U1916 (N_1916,In_1169,In_1149);
or U1917 (N_1917,In_924,In_929);
xor U1918 (N_1918,In_176,In_59);
nand U1919 (N_1919,In_98,In_30);
nor U1920 (N_1920,In_1152,In_306);
nand U1921 (N_1921,In_1156,In_1046);
or U1922 (N_1922,In_441,In_354);
nand U1923 (N_1923,In_1141,In_1156);
and U1924 (N_1924,In_258,In_1221);
xor U1925 (N_1925,In_23,In_797);
nand U1926 (N_1926,In_1438,In_608);
and U1927 (N_1927,In_458,In_328);
or U1928 (N_1928,In_369,In_1415);
and U1929 (N_1929,In_428,In_107);
nor U1930 (N_1930,In_993,In_1216);
nand U1931 (N_1931,In_704,In_1066);
and U1932 (N_1932,In_1255,In_797);
or U1933 (N_1933,In_1331,In_1064);
and U1934 (N_1934,In_247,In_80);
and U1935 (N_1935,In_668,In_802);
or U1936 (N_1936,In_668,In_4);
nor U1937 (N_1937,In_1283,In_54);
xnor U1938 (N_1938,In_702,In_945);
nand U1939 (N_1939,In_974,In_288);
or U1940 (N_1940,In_857,In_936);
nand U1941 (N_1941,In_1131,In_922);
nor U1942 (N_1942,In_1322,In_1493);
or U1943 (N_1943,In_619,In_860);
nand U1944 (N_1944,In_127,In_14);
nand U1945 (N_1945,In_384,In_283);
nand U1946 (N_1946,In_1382,In_264);
nand U1947 (N_1947,In_814,In_1049);
and U1948 (N_1948,In_201,In_586);
nand U1949 (N_1949,In_777,In_796);
nand U1950 (N_1950,In_1122,In_51);
and U1951 (N_1951,In_809,In_222);
nor U1952 (N_1952,In_1366,In_433);
nand U1953 (N_1953,In_916,In_349);
and U1954 (N_1954,In_1292,In_606);
nor U1955 (N_1955,In_1434,In_330);
nor U1956 (N_1956,In_1034,In_1003);
nor U1957 (N_1957,In_744,In_1253);
nor U1958 (N_1958,In_344,In_263);
nor U1959 (N_1959,In_578,In_669);
and U1960 (N_1960,In_458,In_766);
nor U1961 (N_1961,In_1054,In_722);
and U1962 (N_1962,In_392,In_977);
nand U1963 (N_1963,In_409,In_699);
xor U1964 (N_1964,In_1460,In_937);
or U1965 (N_1965,In_335,In_578);
nand U1966 (N_1966,In_71,In_1036);
or U1967 (N_1967,In_1269,In_1290);
nand U1968 (N_1968,In_906,In_396);
nand U1969 (N_1969,In_588,In_34);
and U1970 (N_1970,In_1125,In_45);
or U1971 (N_1971,In_365,In_549);
nand U1972 (N_1972,In_60,In_1062);
nor U1973 (N_1973,In_122,In_637);
xnor U1974 (N_1974,In_1160,In_504);
xnor U1975 (N_1975,In_1149,In_1198);
xor U1976 (N_1976,In_586,In_1037);
or U1977 (N_1977,In_346,In_285);
nor U1978 (N_1978,In_510,In_365);
xor U1979 (N_1979,In_442,In_288);
and U1980 (N_1980,In_287,In_802);
nand U1981 (N_1981,In_541,In_283);
nor U1982 (N_1982,In_41,In_909);
and U1983 (N_1983,In_686,In_1356);
xor U1984 (N_1984,In_1033,In_137);
nor U1985 (N_1985,In_885,In_478);
nor U1986 (N_1986,In_158,In_1441);
or U1987 (N_1987,In_97,In_1312);
nor U1988 (N_1988,In_658,In_871);
or U1989 (N_1989,In_938,In_1136);
and U1990 (N_1990,In_961,In_82);
nor U1991 (N_1991,In_688,In_762);
nor U1992 (N_1992,In_298,In_904);
nand U1993 (N_1993,In_1151,In_1246);
or U1994 (N_1994,In_1362,In_632);
and U1995 (N_1995,In_137,In_280);
xor U1996 (N_1996,In_803,In_1173);
xnor U1997 (N_1997,In_943,In_409);
nand U1998 (N_1998,In_1340,In_462);
xor U1999 (N_1999,In_1093,In_989);
or U2000 (N_2000,In_512,In_874);
nor U2001 (N_2001,In_1165,In_1355);
and U2002 (N_2002,In_569,In_162);
nor U2003 (N_2003,In_1454,In_1019);
nor U2004 (N_2004,In_56,In_860);
and U2005 (N_2005,In_218,In_453);
xnor U2006 (N_2006,In_1122,In_1049);
and U2007 (N_2007,In_904,In_52);
and U2008 (N_2008,In_281,In_1433);
or U2009 (N_2009,In_512,In_188);
nand U2010 (N_2010,In_39,In_147);
or U2011 (N_2011,In_1146,In_1272);
or U2012 (N_2012,In_393,In_1042);
or U2013 (N_2013,In_1381,In_1408);
or U2014 (N_2014,In_1345,In_632);
and U2015 (N_2015,In_1029,In_314);
xor U2016 (N_2016,In_768,In_791);
nor U2017 (N_2017,In_1391,In_701);
nor U2018 (N_2018,In_253,In_323);
nand U2019 (N_2019,In_1232,In_1199);
or U2020 (N_2020,In_411,In_829);
nand U2021 (N_2021,In_1263,In_718);
and U2022 (N_2022,In_49,In_71);
nand U2023 (N_2023,In_596,In_658);
and U2024 (N_2024,In_182,In_111);
or U2025 (N_2025,In_36,In_138);
nor U2026 (N_2026,In_144,In_1435);
and U2027 (N_2027,In_1047,In_76);
or U2028 (N_2028,In_816,In_73);
nand U2029 (N_2029,In_1313,In_465);
nor U2030 (N_2030,In_10,In_1326);
xor U2031 (N_2031,In_515,In_862);
xnor U2032 (N_2032,In_1252,In_118);
nor U2033 (N_2033,In_708,In_252);
nor U2034 (N_2034,In_1367,In_1323);
or U2035 (N_2035,In_172,In_432);
and U2036 (N_2036,In_988,In_187);
nand U2037 (N_2037,In_152,In_383);
and U2038 (N_2038,In_1388,In_785);
or U2039 (N_2039,In_1157,In_1212);
and U2040 (N_2040,In_826,In_985);
xor U2041 (N_2041,In_1059,In_155);
nor U2042 (N_2042,In_248,In_603);
and U2043 (N_2043,In_83,In_1023);
nor U2044 (N_2044,In_1280,In_531);
xor U2045 (N_2045,In_106,In_1018);
xor U2046 (N_2046,In_419,In_237);
or U2047 (N_2047,In_982,In_470);
and U2048 (N_2048,In_1479,In_1202);
nand U2049 (N_2049,In_872,In_674);
xor U2050 (N_2050,In_944,In_147);
or U2051 (N_2051,In_1165,In_616);
nand U2052 (N_2052,In_555,In_698);
and U2053 (N_2053,In_619,In_92);
nand U2054 (N_2054,In_1137,In_772);
or U2055 (N_2055,In_1452,In_0);
and U2056 (N_2056,In_1114,In_1375);
nor U2057 (N_2057,In_1346,In_744);
and U2058 (N_2058,In_409,In_1229);
nor U2059 (N_2059,In_875,In_1329);
or U2060 (N_2060,In_801,In_595);
nand U2061 (N_2061,In_238,In_1173);
or U2062 (N_2062,In_1163,In_893);
nand U2063 (N_2063,In_567,In_113);
or U2064 (N_2064,In_966,In_590);
and U2065 (N_2065,In_894,In_651);
or U2066 (N_2066,In_1378,In_1300);
or U2067 (N_2067,In_615,In_1177);
or U2068 (N_2068,In_35,In_371);
and U2069 (N_2069,In_1165,In_1015);
and U2070 (N_2070,In_82,In_1020);
nand U2071 (N_2071,In_1486,In_1207);
nand U2072 (N_2072,In_1014,In_1202);
or U2073 (N_2073,In_134,In_1343);
and U2074 (N_2074,In_318,In_1077);
or U2075 (N_2075,In_239,In_1240);
nand U2076 (N_2076,In_1157,In_338);
and U2077 (N_2077,In_593,In_1479);
nand U2078 (N_2078,In_1141,In_1361);
and U2079 (N_2079,In_1478,In_756);
and U2080 (N_2080,In_182,In_872);
or U2081 (N_2081,In_1049,In_891);
and U2082 (N_2082,In_60,In_572);
and U2083 (N_2083,In_1059,In_994);
nor U2084 (N_2084,In_746,In_1460);
or U2085 (N_2085,In_274,In_545);
xnor U2086 (N_2086,In_341,In_1283);
nor U2087 (N_2087,In_1408,In_558);
or U2088 (N_2088,In_314,In_347);
or U2089 (N_2089,In_723,In_399);
and U2090 (N_2090,In_890,In_734);
or U2091 (N_2091,In_194,In_1419);
and U2092 (N_2092,In_705,In_272);
and U2093 (N_2093,In_1087,In_1489);
nor U2094 (N_2094,In_740,In_158);
nor U2095 (N_2095,In_159,In_628);
nand U2096 (N_2096,In_43,In_1440);
and U2097 (N_2097,In_935,In_1442);
or U2098 (N_2098,In_884,In_1213);
and U2099 (N_2099,In_853,In_78);
or U2100 (N_2100,In_624,In_1157);
nor U2101 (N_2101,In_342,In_948);
xor U2102 (N_2102,In_956,In_1370);
nand U2103 (N_2103,In_150,In_110);
or U2104 (N_2104,In_825,In_160);
and U2105 (N_2105,In_331,In_597);
or U2106 (N_2106,In_964,In_1245);
xnor U2107 (N_2107,In_574,In_930);
or U2108 (N_2108,In_1490,In_975);
xnor U2109 (N_2109,In_1215,In_1079);
nor U2110 (N_2110,In_257,In_927);
nor U2111 (N_2111,In_780,In_452);
xor U2112 (N_2112,In_993,In_214);
nand U2113 (N_2113,In_277,In_214);
and U2114 (N_2114,In_27,In_1311);
and U2115 (N_2115,In_1204,In_666);
nand U2116 (N_2116,In_799,In_1451);
nand U2117 (N_2117,In_494,In_665);
xnor U2118 (N_2118,In_1186,In_874);
nor U2119 (N_2119,In_561,In_1405);
or U2120 (N_2120,In_917,In_892);
or U2121 (N_2121,In_1484,In_1329);
and U2122 (N_2122,In_315,In_47);
nand U2123 (N_2123,In_116,In_1077);
nor U2124 (N_2124,In_716,In_71);
nor U2125 (N_2125,In_1061,In_1379);
nor U2126 (N_2126,In_185,In_893);
or U2127 (N_2127,In_635,In_356);
and U2128 (N_2128,In_1260,In_183);
nand U2129 (N_2129,In_1314,In_1494);
or U2130 (N_2130,In_711,In_666);
nor U2131 (N_2131,In_1070,In_139);
nor U2132 (N_2132,In_357,In_68);
and U2133 (N_2133,In_692,In_1342);
nand U2134 (N_2134,In_138,In_26);
and U2135 (N_2135,In_606,In_576);
and U2136 (N_2136,In_814,In_423);
nand U2137 (N_2137,In_190,In_1319);
xor U2138 (N_2138,In_867,In_1491);
and U2139 (N_2139,In_647,In_731);
or U2140 (N_2140,In_754,In_1080);
nor U2141 (N_2141,In_673,In_1287);
nor U2142 (N_2142,In_899,In_1348);
nand U2143 (N_2143,In_1195,In_1299);
nand U2144 (N_2144,In_1378,In_462);
nand U2145 (N_2145,In_1457,In_1106);
xor U2146 (N_2146,In_587,In_1140);
nor U2147 (N_2147,In_190,In_457);
nor U2148 (N_2148,In_963,In_822);
xnor U2149 (N_2149,In_1131,In_1295);
or U2150 (N_2150,In_1411,In_1100);
and U2151 (N_2151,In_183,In_412);
xnor U2152 (N_2152,In_519,In_884);
nor U2153 (N_2153,In_851,In_292);
xnor U2154 (N_2154,In_1464,In_289);
nand U2155 (N_2155,In_984,In_1141);
xnor U2156 (N_2156,In_1098,In_1055);
nand U2157 (N_2157,In_1374,In_769);
nand U2158 (N_2158,In_522,In_283);
nor U2159 (N_2159,In_441,In_1019);
nand U2160 (N_2160,In_184,In_108);
and U2161 (N_2161,In_617,In_1246);
and U2162 (N_2162,In_1108,In_1403);
xnor U2163 (N_2163,In_172,In_206);
or U2164 (N_2164,In_585,In_728);
nand U2165 (N_2165,In_304,In_756);
nand U2166 (N_2166,In_221,In_353);
nand U2167 (N_2167,In_546,In_833);
or U2168 (N_2168,In_552,In_835);
xor U2169 (N_2169,In_1282,In_11);
and U2170 (N_2170,In_622,In_1214);
or U2171 (N_2171,In_715,In_661);
or U2172 (N_2172,In_1139,In_1141);
and U2173 (N_2173,In_1279,In_1400);
nand U2174 (N_2174,In_1046,In_1221);
xor U2175 (N_2175,In_48,In_401);
and U2176 (N_2176,In_1203,In_594);
nor U2177 (N_2177,In_1135,In_1366);
nor U2178 (N_2178,In_28,In_850);
or U2179 (N_2179,In_1304,In_584);
nor U2180 (N_2180,In_975,In_180);
nor U2181 (N_2181,In_1494,In_187);
or U2182 (N_2182,In_65,In_1238);
xnor U2183 (N_2183,In_1233,In_441);
nor U2184 (N_2184,In_12,In_193);
and U2185 (N_2185,In_1317,In_1244);
or U2186 (N_2186,In_327,In_48);
and U2187 (N_2187,In_1353,In_1472);
and U2188 (N_2188,In_1317,In_560);
or U2189 (N_2189,In_126,In_649);
and U2190 (N_2190,In_1182,In_785);
or U2191 (N_2191,In_193,In_107);
and U2192 (N_2192,In_146,In_470);
nor U2193 (N_2193,In_1307,In_847);
xnor U2194 (N_2194,In_1452,In_675);
nand U2195 (N_2195,In_454,In_158);
or U2196 (N_2196,In_284,In_1252);
xnor U2197 (N_2197,In_948,In_1006);
and U2198 (N_2198,In_1471,In_1422);
or U2199 (N_2199,In_1422,In_1106);
nor U2200 (N_2200,In_1271,In_610);
or U2201 (N_2201,In_96,In_987);
and U2202 (N_2202,In_1001,In_1285);
or U2203 (N_2203,In_963,In_312);
or U2204 (N_2204,In_1271,In_1104);
xor U2205 (N_2205,In_722,In_1024);
nand U2206 (N_2206,In_228,In_32);
nand U2207 (N_2207,In_179,In_1498);
nand U2208 (N_2208,In_966,In_855);
xor U2209 (N_2209,In_782,In_885);
or U2210 (N_2210,In_613,In_892);
nor U2211 (N_2211,In_705,In_115);
nor U2212 (N_2212,In_136,In_919);
or U2213 (N_2213,In_689,In_1001);
xor U2214 (N_2214,In_104,In_390);
nand U2215 (N_2215,In_1226,In_516);
or U2216 (N_2216,In_1415,In_958);
nor U2217 (N_2217,In_1286,In_136);
nand U2218 (N_2218,In_531,In_870);
or U2219 (N_2219,In_1072,In_464);
nand U2220 (N_2220,In_907,In_828);
or U2221 (N_2221,In_83,In_1418);
or U2222 (N_2222,In_1468,In_413);
and U2223 (N_2223,In_664,In_990);
nor U2224 (N_2224,In_878,In_628);
nor U2225 (N_2225,In_659,In_59);
or U2226 (N_2226,In_1174,In_32);
or U2227 (N_2227,In_1305,In_74);
nor U2228 (N_2228,In_421,In_365);
nand U2229 (N_2229,In_1172,In_1363);
nor U2230 (N_2230,In_1174,In_131);
and U2231 (N_2231,In_1470,In_1194);
nand U2232 (N_2232,In_1289,In_572);
or U2233 (N_2233,In_1306,In_724);
and U2234 (N_2234,In_724,In_775);
and U2235 (N_2235,In_722,In_1213);
nor U2236 (N_2236,In_219,In_1113);
nor U2237 (N_2237,In_16,In_155);
and U2238 (N_2238,In_1041,In_647);
nand U2239 (N_2239,In_1264,In_76);
and U2240 (N_2240,In_191,In_374);
xor U2241 (N_2241,In_962,In_595);
nor U2242 (N_2242,In_305,In_426);
nand U2243 (N_2243,In_1449,In_311);
or U2244 (N_2244,In_1149,In_1374);
or U2245 (N_2245,In_436,In_1422);
nor U2246 (N_2246,In_846,In_821);
and U2247 (N_2247,In_921,In_390);
or U2248 (N_2248,In_707,In_826);
or U2249 (N_2249,In_1177,In_671);
nor U2250 (N_2250,In_1024,In_160);
nor U2251 (N_2251,In_387,In_78);
nand U2252 (N_2252,In_900,In_402);
or U2253 (N_2253,In_393,In_1090);
nand U2254 (N_2254,In_1432,In_1229);
or U2255 (N_2255,In_946,In_528);
nand U2256 (N_2256,In_71,In_1123);
nor U2257 (N_2257,In_718,In_430);
nor U2258 (N_2258,In_625,In_653);
xnor U2259 (N_2259,In_1023,In_289);
or U2260 (N_2260,In_1166,In_1103);
or U2261 (N_2261,In_1154,In_1197);
or U2262 (N_2262,In_547,In_929);
nand U2263 (N_2263,In_1025,In_767);
nand U2264 (N_2264,In_179,In_72);
and U2265 (N_2265,In_416,In_53);
nor U2266 (N_2266,In_23,In_1256);
and U2267 (N_2267,In_1106,In_1252);
and U2268 (N_2268,In_4,In_425);
or U2269 (N_2269,In_481,In_1129);
or U2270 (N_2270,In_67,In_364);
and U2271 (N_2271,In_831,In_782);
nor U2272 (N_2272,In_1472,In_1327);
or U2273 (N_2273,In_78,In_436);
nor U2274 (N_2274,In_1308,In_223);
nor U2275 (N_2275,In_880,In_259);
nor U2276 (N_2276,In_859,In_1358);
or U2277 (N_2277,In_808,In_830);
nor U2278 (N_2278,In_16,In_828);
or U2279 (N_2279,In_1445,In_1349);
or U2280 (N_2280,In_349,In_46);
or U2281 (N_2281,In_563,In_74);
nand U2282 (N_2282,In_262,In_1337);
or U2283 (N_2283,In_1235,In_975);
nand U2284 (N_2284,In_299,In_91);
or U2285 (N_2285,In_1042,In_853);
xor U2286 (N_2286,In_370,In_254);
nor U2287 (N_2287,In_1359,In_514);
and U2288 (N_2288,In_84,In_464);
or U2289 (N_2289,In_883,In_496);
and U2290 (N_2290,In_1223,In_620);
or U2291 (N_2291,In_16,In_518);
nor U2292 (N_2292,In_481,In_507);
nor U2293 (N_2293,In_616,In_1032);
xor U2294 (N_2294,In_395,In_1333);
nand U2295 (N_2295,In_851,In_1189);
and U2296 (N_2296,In_195,In_272);
xor U2297 (N_2297,In_731,In_987);
nor U2298 (N_2298,In_624,In_578);
or U2299 (N_2299,In_631,In_1272);
nand U2300 (N_2300,In_1346,In_1194);
or U2301 (N_2301,In_797,In_28);
nand U2302 (N_2302,In_58,In_35);
nor U2303 (N_2303,In_169,In_650);
nor U2304 (N_2304,In_1055,In_787);
nor U2305 (N_2305,In_582,In_93);
nor U2306 (N_2306,In_1125,In_1352);
nand U2307 (N_2307,In_262,In_1428);
nand U2308 (N_2308,In_1453,In_905);
nand U2309 (N_2309,In_391,In_129);
or U2310 (N_2310,In_477,In_336);
nor U2311 (N_2311,In_559,In_1277);
nand U2312 (N_2312,In_1348,In_467);
nand U2313 (N_2313,In_165,In_293);
nor U2314 (N_2314,In_1048,In_420);
and U2315 (N_2315,In_491,In_454);
or U2316 (N_2316,In_688,In_1147);
nand U2317 (N_2317,In_285,In_839);
or U2318 (N_2318,In_664,In_909);
and U2319 (N_2319,In_1101,In_1210);
nor U2320 (N_2320,In_555,In_840);
or U2321 (N_2321,In_782,In_304);
nor U2322 (N_2322,In_679,In_362);
xnor U2323 (N_2323,In_1006,In_524);
nor U2324 (N_2324,In_393,In_111);
and U2325 (N_2325,In_854,In_158);
xnor U2326 (N_2326,In_63,In_1071);
nand U2327 (N_2327,In_214,In_1088);
nor U2328 (N_2328,In_1440,In_442);
xnor U2329 (N_2329,In_917,In_368);
or U2330 (N_2330,In_655,In_1238);
or U2331 (N_2331,In_819,In_738);
nand U2332 (N_2332,In_923,In_1044);
nor U2333 (N_2333,In_799,In_1415);
or U2334 (N_2334,In_1097,In_946);
xnor U2335 (N_2335,In_1320,In_1254);
nor U2336 (N_2336,In_130,In_805);
or U2337 (N_2337,In_963,In_1469);
nor U2338 (N_2338,In_461,In_105);
nor U2339 (N_2339,In_45,In_1248);
and U2340 (N_2340,In_1325,In_1090);
and U2341 (N_2341,In_1143,In_356);
and U2342 (N_2342,In_879,In_320);
xor U2343 (N_2343,In_40,In_1296);
nor U2344 (N_2344,In_136,In_712);
xor U2345 (N_2345,In_856,In_622);
or U2346 (N_2346,In_1425,In_840);
nand U2347 (N_2347,In_1297,In_1299);
nand U2348 (N_2348,In_355,In_410);
and U2349 (N_2349,In_727,In_98);
nand U2350 (N_2350,In_959,In_1283);
or U2351 (N_2351,In_1024,In_510);
and U2352 (N_2352,In_579,In_1067);
nand U2353 (N_2353,In_142,In_1221);
nor U2354 (N_2354,In_669,In_72);
nor U2355 (N_2355,In_628,In_181);
and U2356 (N_2356,In_266,In_853);
nand U2357 (N_2357,In_147,In_335);
and U2358 (N_2358,In_178,In_1223);
and U2359 (N_2359,In_1490,In_800);
nor U2360 (N_2360,In_856,In_298);
nor U2361 (N_2361,In_91,In_603);
xnor U2362 (N_2362,In_599,In_785);
nor U2363 (N_2363,In_1133,In_1394);
and U2364 (N_2364,In_419,In_271);
nand U2365 (N_2365,In_282,In_242);
nor U2366 (N_2366,In_212,In_622);
or U2367 (N_2367,In_1118,In_1449);
nand U2368 (N_2368,In_863,In_175);
nor U2369 (N_2369,In_177,In_392);
nor U2370 (N_2370,In_378,In_207);
and U2371 (N_2371,In_1170,In_481);
and U2372 (N_2372,In_367,In_120);
or U2373 (N_2373,In_776,In_1432);
and U2374 (N_2374,In_1411,In_1456);
or U2375 (N_2375,In_893,In_283);
nor U2376 (N_2376,In_839,In_845);
or U2377 (N_2377,In_19,In_891);
xor U2378 (N_2378,In_94,In_545);
nor U2379 (N_2379,In_553,In_995);
nor U2380 (N_2380,In_1247,In_1273);
or U2381 (N_2381,In_338,In_1481);
nand U2382 (N_2382,In_959,In_251);
nand U2383 (N_2383,In_1375,In_338);
or U2384 (N_2384,In_437,In_662);
xor U2385 (N_2385,In_10,In_1292);
nor U2386 (N_2386,In_60,In_1122);
xnor U2387 (N_2387,In_110,In_550);
nand U2388 (N_2388,In_1370,In_1071);
nor U2389 (N_2389,In_61,In_982);
nor U2390 (N_2390,In_928,In_1235);
or U2391 (N_2391,In_966,In_766);
or U2392 (N_2392,In_440,In_9);
nor U2393 (N_2393,In_625,In_1057);
nand U2394 (N_2394,In_1464,In_817);
nor U2395 (N_2395,In_891,In_358);
nor U2396 (N_2396,In_1243,In_1286);
nand U2397 (N_2397,In_878,In_1412);
or U2398 (N_2398,In_1261,In_271);
nand U2399 (N_2399,In_1354,In_138);
nor U2400 (N_2400,In_610,In_666);
nor U2401 (N_2401,In_1423,In_801);
and U2402 (N_2402,In_1012,In_445);
and U2403 (N_2403,In_1150,In_80);
nor U2404 (N_2404,In_973,In_66);
nor U2405 (N_2405,In_591,In_405);
or U2406 (N_2406,In_260,In_1483);
and U2407 (N_2407,In_773,In_1040);
nand U2408 (N_2408,In_1290,In_1201);
or U2409 (N_2409,In_895,In_1120);
or U2410 (N_2410,In_879,In_337);
or U2411 (N_2411,In_962,In_126);
or U2412 (N_2412,In_109,In_1173);
and U2413 (N_2413,In_57,In_891);
nor U2414 (N_2414,In_302,In_631);
nand U2415 (N_2415,In_1130,In_1417);
nor U2416 (N_2416,In_251,In_995);
xnor U2417 (N_2417,In_712,In_1273);
or U2418 (N_2418,In_150,In_148);
nand U2419 (N_2419,In_1087,In_1491);
or U2420 (N_2420,In_466,In_814);
xnor U2421 (N_2421,In_1026,In_624);
or U2422 (N_2422,In_728,In_1377);
nor U2423 (N_2423,In_911,In_704);
xnor U2424 (N_2424,In_949,In_992);
or U2425 (N_2425,In_1312,In_640);
nand U2426 (N_2426,In_522,In_382);
and U2427 (N_2427,In_869,In_660);
nor U2428 (N_2428,In_1258,In_425);
nor U2429 (N_2429,In_210,In_582);
or U2430 (N_2430,In_1125,In_1106);
nor U2431 (N_2431,In_1156,In_371);
xnor U2432 (N_2432,In_1131,In_1292);
and U2433 (N_2433,In_407,In_71);
or U2434 (N_2434,In_1354,In_860);
and U2435 (N_2435,In_27,In_21);
nor U2436 (N_2436,In_530,In_1390);
nor U2437 (N_2437,In_822,In_148);
nand U2438 (N_2438,In_1254,In_1023);
and U2439 (N_2439,In_691,In_1200);
nand U2440 (N_2440,In_1326,In_1152);
nand U2441 (N_2441,In_1418,In_742);
and U2442 (N_2442,In_999,In_871);
and U2443 (N_2443,In_220,In_1033);
or U2444 (N_2444,In_1374,In_1371);
xnor U2445 (N_2445,In_854,In_960);
xnor U2446 (N_2446,In_1435,In_1182);
nand U2447 (N_2447,In_890,In_1127);
nor U2448 (N_2448,In_1241,In_873);
and U2449 (N_2449,In_1223,In_278);
or U2450 (N_2450,In_613,In_743);
and U2451 (N_2451,In_1342,In_80);
xnor U2452 (N_2452,In_1403,In_62);
nor U2453 (N_2453,In_1079,In_1170);
nor U2454 (N_2454,In_1249,In_751);
or U2455 (N_2455,In_1234,In_276);
and U2456 (N_2456,In_398,In_1118);
or U2457 (N_2457,In_1063,In_24);
and U2458 (N_2458,In_1220,In_1290);
or U2459 (N_2459,In_164,In_1476);
or U2460 (N_2460,In_520,In_1180);
or U2461 (N_2461,In_44,In_1023);
nand U2462 (N_2462,In_1021,In_674);
nor U2463 (N_2463,In_508,In_754);
and U2464 (N_2464,In_1001,In_927);
nor U2465 (N_2465,In_1176,In_603);
nor U2466 (N_2466,In_1000,In_1224);
and U2467 (N_2467,In_13,In_1134);
or U2468 (N_2468,In_178,In_292);
nor U2469 (N_2469,In_1166,In_353);
nand U2470 (N_2470,In_601,In_1136);
or U2471 (N_2471,In_317,In_1359);
or U2472 (N_2472,In_415,In_1396);
or U2473 (N_2473,In_0,In_1134);
and U2474 (N_2474,In_1362,In_827);
or U2475 (N_2475,In_796,In_889);
nor U2476 (N_2476,In_1161,In_986);
xnor U2477 (N_2477,In_725,In_976);
nor U2478 (N_2478,In_380,In_648);
or U2479 (N_2479,In_522,In_488);
nor U2480 (N_2480,In_806,In_357);
xnor U2481 (N_2481,In_598,In_666);
nor U2482 (N_2482,In_742,In_847);
nor U2483 (N_2483,In_1426,In_164);
or U2484 (N_2484,In_399,In_1127);
nand U2485 (N_2485,In_303,In_78);
nand U2486 (N_2486,In_130,In_1252);
nand U2487 (N_2487,In_549,In_1012);
nand U2488 (N_2488,In_174,In_1406);
nor U2489 (N_2489,In_1140,In_905);
nand U2490 (N_2490,In_420,In_570);
nand U2491 (N_2491,In_298,In_1149);
or U2492 (N_2492,In_226,In_433);
or U2493 (N_2493,In_1000,In_691);
nand U2494 (N_2494,In_1186,In_1418);
or U2495 (N_2495,In_1032,In_1345);
nand U2496 (N_2496,In_44,In_739);
and U2497 (N_2497,In_191,In_722);
xnor U2498 (N_2498,In_791,In_604);
nor U2499 (N_2499,In_1228,In_739);
nor U2500 (N_2500,In_814,In_923);
or U2501 (N_2501,In_1070,In_1423);
nor U2502 (N_2502,In_755,In_1216);
or U2503 (N_2503,In_643,In_986);
xor U2504 (N_2504,In_845,In_28);
or U2505 (N_2505,In_974,In_382);
or U2506 (N_2506,In_1026,In_1010);
nor U2507 (N_2507,In_82,In_840);
and U2508 (N_2508,In_1015,In_1202);
and U2509 (N_2509,In_1215,In_89);
nor U2510 (N_2510,In_382,In_977);
or U2511 (N_2511,In_283,In_615);
or U2512 (N_2512,In_477,In_676);
and U2513 (N_2513,In_443,In_377);
nor U2514 (N_2514,In_56,In_1398);
and U2515 (N_2515,In_633,In_843);
nand U2516 (N_2516,In_873,In_628);
and U2517 (N_2517,In_1194,In_141);
nand U2518 (N_2518,In_948,In_165);
or U2519 (N_2519,In_1316,In_230);
nand U2520 (N_2520,In_446,In_709);
nand U2521 (N_2521,In_296,In_549);
xor U2522 (N_2522,In_761,In_353);
nor U2523 (N_2523,In_575,In_951);
or U2524 (N_2524,In_696,In_327);
nand U2525 (N_2525,In_725,In_42);
nand U2526 (N_2526,In_37,In_681);
nand U2527 (N_2527,In_568,In_1003);
and U2528 (N_2528,In_290,In_927);
nor U2529 (N_2529,In_857,In_1461);
xnor U2530 (N_2530,In_102,In_1211);
nand U2531 (N_2531,In_1245,In_1362);
nand U2532 (N_2532,In_1420,In_1367);
nand U2533 (N_2533,In_514,In_349);
nand U2534 (N_2534,In_625,In_534);
xnor U2535 (N_2535,In_1356,In_492);
nand U2536 (N_2536,In_404,In_439);
or U2537 (N_2537,In_762,In_565);
nor U2538 (N_2538,In_58,In_692);
xnor U2539 (N_2539,In_1307,In_461);
and U2540 (N_2540,In_1183,In_433);
nor U2541 (N_2541,In_379,In_729);
or U2542 (N_2542,In_48,In_740);
or U2543 (N_2543,In_1195,In_284);
nor U2544 (N_2544,In_1312,In_1275);
nand U2545 (N_2545,In_563,In_71);
nor U2546 (N_2546,In_1485,In_682);
and U2547 (N_2547,In_420,In_1076);
nand U2548 (N_2548,In_147,In_1442);
and U2549 (N_2549,In_844,In_762);
and U2550 (N_2550,In_376,In_107);
nand U2551 (N_2551,In_646,In_1196);
nand U2552 (N_2552,In_297,In_888);
and U2553 (N_2553,In_1203,In_1042);
nor U2554 (N_2554,In_1379,In_950);
or U2555 (N_2555,In_1408,In_159);
nand U2556 (N_2556,In_965,In_73);
and U2557 (N_2557,In_719,In_917);
nand U2558 (N_2558,In_555,In_554);
xnor U2559 (N_2559,In_439,In_1030);
and U2560 (N_2560,In_216,In_357);
xnor U2561 (N_2561,In_1396,In_1216);
nor U2562 (N_2562,In_1435,In_343);
nor U2563 (N_2563,In_1499,In_250);
xnor U2564 (N_2564,In_280,In_601);
nor U2565 (N_2565,In_1443,In_1158);
nand U2566 (N_2566,In_671,In_499);
nor U2567 (N_2567,In_626,In_222);
nor U2568 (N_2568,In_399,In_90);
xor U2569 (N_2569,In_499,In_510);
or U2570 (N_2570,In_603,In_572);
and U2571 (N_2571,In_318,In_1393);
nor U2572 (N_2572,In_9,In_1406);
xnor U2573 (N_2573,In_993,In_1453);
nor U2574 (N_2574,In_1085,In_1018);
nor U2575 (N_2575,In_769,In_77);
nand U2576 (N_2576,In_1042,In_981);
xor U2577 (N_2577,In_1244,In_1336);
and U2578 (N_2578,In_234,In_1198);
nor U2579 (N_2579,In_645,In_1061);
nand U2580 (N_2580,In_673,In_109);
xnor U2581 (N_2581,In_152,In_1248);
xor U2582 (N_2582,In_55,In_617);
nand U2583 (N_2583,In_757,In_864);
and U2584 (N_2584,In_1160,In_848);
or U2585 (N_2585,In_555,In_21);
or U2586 (N_2586,In_47,In_708);
xor U2587 (N_2587,In_2,In_887);
or U2588 (N_2588,In_750,In_257);
or U2589 (N_2589,In_1490,In_1451);
xnor U2590 (N_2590,In_1081,In_147);
nor U2591 (N_2591,In_756,In_1098);
nand U2592 (N_2592,In_1392,In_36);
nand U2593 (N_2593,In_885,In_1499);
nor U2594 (N_2594,In_241,In_311);
and U2595 (N_2595,In_58,In_290);
and U2596 (N_2596,In_1493,In_853);
and U2597 (N_2597,In_3,In_209);
nor U2598 (N_2598,In_1453,In_971);
nor U2599 (N_2599,In_714,In_955);
nand U2600 (N_2600,In_1228,In_1339);
nand U2601 (N_2601,In_366,In_26);
nor U2602 (N_2602,In_700,In_371);
nand U2603 (N_2603,In_1209,In_319);
nor U2604 (N_2604,In_621,In_1405);
and U2605 (N_2605,In_586,In_721);
nor U2606 (N_2606,In_38,In_272);
nor U2607 (N_2607,In_420,In_1214);
nor U2608 (N_2608,In_356,In_1387);
nand U2609 (N_2609,In_544,In_1010);
and U2610 (N_2610,In_1495,In_1055);
nand U2611 (N_2611,In_1009,In_1178);
nand U2612 (N_2612,In_76,In_308);
or U2613 (N_2613,In_760,In_924);
and U2614 (N_2614,In_859,In_1170);
or U2615 (N_2615,In_140,In_12);
nor U2616 (N_2616,In_827,In_245);
nor U2617 (N_2617,In_1463,In_907);
and U2618 (N_2618,In_331,In_484);
nand U2619 (N_2619,In_317,In_1331);
or U2620 (N_2620,In_1339,In_1307);
and U2621 (N_2621,In_424,In_471);
nand U2622 (N_2622,In_714,In_153);
or U2623 (N_2623,In_651,In_363);
and U2624 (N_2624,In_1362,In_1326);
and U2625 (N_2625,In_1422,In_685);
and U2626 (N_2626,In_914,In_1216);
or U2627 (N_2627,In_746,In_181);
and U2628 (N_2628,In_854,In_1002);
nor U2629 (N_2629,In_1396,In_806);
or U2630 (N_2630,In_236,In_245);
nand U2631 (N_2631,In_1294,In_80);
and U2632 (N_2632,In_4,In_71);
and U2633 (N_2633,In_1090,In_1331);
nand U2634 (N_2634,In_790,In_691);
and U2635 (N_2635,In_1261,In_248);
nor U2636 (N_2636,In_145,In_1397);
or U2637 (N_2637,In_49,In_240);
nand U2638 (N_2638,In_347,In_1299);
and U2639 (N_2639,In_973,In_114);
and U2640 (N_2640,In_63,In_551);
nand U2641 (N_2641,In_676,In_1325);
and U2642 (N_2642,In_534,In_1303);
and U2643 (N_2643,In_257,In_822);
nor U2644 (N_2644,In_375,In_634);
or U2645 (N_2645,In_516,In_162);
and U2646 (N_2646,In_742,In_191);
nor U2647 (N_2647,In_1107,In_793);
nor U2648 (N_2648,In_118,In_1088);
nor U2649 (N_2649,In_942,In_562);
or U2650 (N_2650,In_91,In_957);
or U2651 (N_2651,In_158,In_1320);
xor U2652 (N_2652,In_1346,In_1178);
or U2653 (N_2653,In_158,In_1298);
and U2654 (N_2654,In_1345,In_613);
and U2655 (N_2655,In_972,In_300);
xnor U2656 (N_2656,In_1018,In_291);
or U2657 (N_2657,In_184,In_742);
xor U2658 (N_2658,In_649,In_458);
and U2659 (N_2659,In_1485,In_758);
nand U2660 (N_2660,In_942,In_493);
nor U2661 (N_2661,In_1240,In_1223);
and U2662 (N_2662,In_1188,In_757);
nor U2663 (N_2663,In_542,In_679);
nor U2664 (N_2664,In_1158,In_1456);
nand U2665 (N_2665,In_468,In_0);
nand U2666 (N_2666,In_282,In_608);
nor U2667 (N_2667,In_813,In_544);
nand U2668 (N_2668,In_627,In_1123);
and U2669 (N_2669,In_1015,In_1351);
or U2670 (N_2670,In_761,In_1281);
and U2671 (N_2671,In_156,In_566);
or U2672 (N_2672,In_188,In_313);
and U2673 (N_2673,In_4,In_934);
or U2674 (N_2674,In_1165,In_1455);
nand U2675 (N_2675,In_639,In_790);
and U2676 (N_2676,In_1395,In_1167);
and U2677 (N_2677,In_180,In_443);
or U2678 (N_2678,In_1222,In_820);
nand U2679 (N_2679,In_586,In_325);
and U2680 (N_2680,In_159,In_1185);
or U2681 (N_2681,In_855,In_419);
nor U2682 (N_2682,In_1327,In_831);
and U2683 (N_2683,In_1343,In_152);
nand U2684 (N_2684,In_1469,In_375);
nand U2685 (N_2685,In_157,In_1033);
nand U2686 (N_2686,In_1287,In_92);
xnor U2687 (N_2687,In_855,In_1226);
and U2688 (N_2688,In_1280,In_247);
nor U2689 (N_2689,In_569,In_451);
and U2690 (N_2690,In_727,In_305);
and U2691 (N_2691,In_1241,In_1259);
nor U2692 (N_2692,In_182,In_1339);
nor U2693 (N_2693,In_868,In_647);
xor U2694 (N_2694,In_628,In_1215);
nand U2695 (N_2695,In_560,In_399);
nand U2696 (N_2696,In_67,In_696);
nand U2697 (N_2697,In_1293,In_175);
nand U2698 (N_2698,In_1410,In_80);
and U2699 (N_2699,In_1112,In_699);
and U2700 (N_2700,In_991,In_42);
nand U2701 (N_2701,In_1475,In_985);
nand U2702 (N_2702,In_125,In_1178);
nor U2703 (N_2703,In_25,In_1037);
nand U2704 (N_2704,In_250,In_1069);
or U2705 (N_2705,In_429,In_264);
and U2706 (N_2706,In_836,In_1284);
and U2707 (N_2707,In_67,In_1070);
and U2708 (N_2708,In_708,In_406);
nand U2709 (N_2709,In_706,In_1397);
and U2710 (N_2710,In_1175,In_584);
or U2711 (N_2711,In_1427,In_608);
nor U2712 (N_2712,In_694,In_913);
and U2713 (N_2713,In_436,In_1418);
nand U2714 (N_2714,In_657,In_1372);
nand U2715 (N_2715,In_205,In_1362);
nor U2716 (N_2716,In_1472,In_712);
nor U2717 (N_2717,In_1457,In_1260);
and U2718 (N_2718,In_1325,In_1049);
nand U2719 (N_2719,In_90,In_893);
nand U2720 (N_2720,In_857,In_947);
and U2721 (N_2721,In_1312,In_689);
nor U2722 (N_2722,In_417,In_1499);
and U2723 (N_2723,In_917,In_1211);
nand U2724 (N_2724,In_1465,In_208);
xor U2725 (N_2725,In_923,In_922);
nand U2726 (N_2726,In_486,In_744);
and U2727 (N_2727,In_234,In_163);
nand U2728 (N_2728,In_1450,In_1167);
or U2729 (N_2729,In_425,In_1406);
nor U2730 (N_2730,In_246,In_37);
nor U2731 (N_2731,In_1340,In_862);
and U2732 (N_2732,In_464,In_528);
nor U2733 (N_2733,In_1049,In_1409);
and U2734 (N_2734,In_1164,In_915);
and U2735 (N_2735,In_39,In_383);
and U2736 (N_2736,In_608,In_451);
nor U2737 (N_2737,In_529,In_279);
and U2738 (N_2738,In_24,In_786);
nor U2739 (N_2739,In_1374,In_824);
nor U2740 (N_2740,In_1087,In_1047);
and U2741 (N_2741,In_47,In_773);
xnor U2742 (N_2742,In_912,In_557);
nor U2743 (N_2743,In_541,In_771);
nand U2744 (N_2744,In_529,In_775);
and U2745 (N_2745,In_41,In_1418);
nor U2746 (N_2746,In_193,In_805);
and U2747 (N_2747,In_1191,In_886);
xor U2748 (N_2748,In_1223,In_322);
nor U2749 (N_2749,In_994,In_1283);
nor U2750 (N_2750,In_472,In_1488);
nor U2751 (N_2751,In_878,In_265);
xor U2752 (N_2752,In_546,In_307);
and U2753 (N_2753,In_1033,In_1267);
and U2754 (N_2754,In_519,In_1145);
or U2755 (N_2755,In_433,In_1278);
and U2756 (N_2756,In_1263,In_1320);
or U2757 (N_2757,In_834,In_1046);
xor U2758 (N_2758,In_491,In_886);
nand U2759 (N_2759,In_861,In_1074);
nand U2760 (N_2760,In_1110,In_211);
nand U2761 (N_2761,In_614,In_1110);
or U2762 (N_2762,In_1132,In_327);
nand U2763 (N_2763,In_1027,In_40);
and U2764 (N_2764,In_1094,In_687);
nor U2765 (N_2765,In_77,In_845);
and U2766 (N_2766,In_798,In_926);
and U2767 (N_2767,In_848,In_1352);
and U2768 (N_2768,In_1324,In_119);
xnor U2769 (N_2769,In_525,In_706);
and U2770 (N_2770,In_64,In_288);
and U2771 (N_2771,In_1366,In_359);
nand U2772 (N_2772,In_421,In_49);
nor U2773 (N_2773,In_1076,In_606);
and U2774 (N_2774,In_900,In_1031);
nor U2775 (N_2775,In_1128,In_1288);
nand U2776 (N_2776,In_913,In_607);
nand U2777 (N_2777,In_1212,In_1491);
or U2778 (N_2778,In_620,In_1326);
nand U2779 (N_2779,In_1241,In_1239);
nand U2780 (N_2780,In_296,In_418);
or U2781 (N_2781,In_954,In_633);
xor U2782 (N_2782,In_631,In_1421);
nor U2783 (N_2783,In_1209,In_757);
or U2784 (N_2784,In_1457,In_1293);
nor U2785 (N_2785,In_396,In_750);
nand U2786 (N_2786,In_1157,In_1340);
nor U2787 (N_2787,In_1362,In_985);
or U2788 (N_2788,In_606,In_447);
or U2789 (N_2789,In_113,In_446);
xnor U2790 (N_2790,In_598,In_1477);
xor U2791 (N_2791,In_1369,In_1013);
or U2792 (N_2792,In_637,In_1122);
nand U2793 (N_2793,In_882,In_970);
nor U2794 (N_2794,In_74,In_128);
and U2795 (N_2795,In_1059,In_1492);
nand U2796 (N_2796,In_1433,In_809);
nand U2797 (N_2797,In_491,In_990);
nand U2798 (N_2798,In_1079,In_1347);
nand U2799 (N_2799,In_915,In_509);
nand U2800 (N_2800,In_1212,In_358);
or U2801 (N_2801,In_1087,In_1233);
and U2802 (N_2802,In_387,In_373);
nand U2803 (N_2803,In_439,In_36);
nand U2804 (N_2804,In_732,In_720);
nand U2805 (N_2805,In_394,In_215);
nor U2806 (N_2806,In_836,In_1266);
or U2807 (N_2807,In_950,In_200);
and U2808 (N_2808,In_490,In_425);
or U2809 (N_2809,In_1259,In_1390);
and U2810 (N_2810,In_1234,In_1156);
nor U2811 (N_2811,In_1493,In_459);
nand U2812 (N_2812,In_152,In_956);
nand U2813 (N_2813,In_1477,In_877);
nor U2814 (N_2814,In_1139,In_1181);
and U2815 (N_2815,In_87,In_824);
and U2816 (N_2816,In_333,In_1258);
and U2817 (N_2817,In_646,In_1055);
and U2818 (N_2818,In_1091,In_1412);
and U2819 (N_2819,In_1436,In_119);
or U2820 (N_2820,In_173,In_827);
or U2821 (N_2821,In_1242,In_210);
and U2822 (N_2822,In_1107,In_277);
nand U2823 (N_2823,In_145,In_209);
nand U2824 (N_2824,In_1142,In_471);
nor U2825 (N_2825,In_1244,In_424);
and U2826 (N_2826,In_119,In_782);
or U2827 (N_2827,In_1461,In_1398);
or U2828 (N_2828,In_1144,In_1306);
or U2829 (N_2829,In_1211,In_202);
and U2830 (N_2830,In_1044,In_855);
and U2831 (N_2831,In_168,In_190);
or U2832 (N_2832,In_1079,In_74);
xor U2833 (N_2833,In_1352,In_948);
nor U2834 (N_2834,In_1412,In_1093);
and U2835 (N_2835,In_508,In_911);
and U2836 (N_2836,In_1224,In_812);
or U2837 (N_2837,In_531,In_883);
xnor U2838 (N_2838,In_429,In_1045);
nand U2839 (N_2839,In_350,In_1128);
nand U2840 (N_2840,In_541,In_112);
and U2841 (N_2841,In_213,In_1032);
nand U2842 (N_2842,In_966,In_1292);
nand U2843 (N_2843,In_188,In_1164);
nand U2844 (N_2844,In_576,In_424);
nand U2845 (N_2845,In_445,In_652);
or U2846 (N_2846,In_1153,In_181);
and U2847 (N_2847,In_116,In_1183);
or U2848 (N_2848,In_743,In_377);
and U2849 (N_2849,In_64,In_485);
or U2850 (N_2850,In_247,In_1017);
or U2851 (N_2851,In_1439,In_705);
and U2852 (N_2852,In_405,In_883);
and U2853 (N_2853,In_499,In_34);
and U2854 (N_2854,In_545,In_1232);
and U2855 (N_2855,In_357,In_175);
nand U2856 (N_2856,In_878,In_1466);
nor U2857 (N_2857,In_508,In_513);
nor U2858 (N_2858,In_224,In_1189);
and U2859 (N_2859,In_938,In_745);
nand U2860 (N_2860,In_1088,In_1410);
or U2861 (N_2861,In_1204,In_1305);
or U2862 (N_2862,In_1278,In_1434);
xor U2863 (N_2863,In_28,In_1357);
and U2864 (N_2864,In_1378,In_381);
nand U2865 (N_2865,In_146,In_650);
or U2866 (N_2866,In_238,In_91);
nor U2867 (N_2867,In_695,In_1199);
nor U2868 (N_2868,In_1416,In_125);
and U2869 (N_2869,In_158,In_750);
and U2870 (N_2870,In_962,In_427);
or U2871 (N_2871,In_962,In_250);
and U2872 (N_2872,In_1376,In_798);
nand U2873 (N_2873,In_745,In_478);
or U2874 (N_2874,In_1291,In_450);
nand U2875 (N_2875,In_334,In_85);
xor U2876 (N_2876,In_788,In_1035);
nand U2877 (N_2877,In_124,In_719);
and U2878 (N_2878,In_562,In_140);
and U2879 (N_2879,In_914,In_927);
nor U2880 (N_2880,In_254,In_284);
or U2881 (N_2881,In_756,In_1041);
nand U2882 (N_2882,In_857,In_873);
and U2883 (N_2883,In_751,In_636);
nand U2884 (N_2884,In_703,In_1059);
nand U2885 (N_2885,In_647,In_307);
nand U2886 (N_2886,In_983,In_1175);
nand U2887 (N_2887,In_132,In_533);
and U2888 (N_2888,In_714,In_958);
nand U2889 (N_2889,In_121,In_1114);
nor U2890 (N_2890,In_996,In_906);
or U2891 (N_2891,In_55,In_716);
or U2892 (N_2892,In_1271,In_1273);
nor U2893 (N_2893,In_167,In_194);
nor U2894 (N_2894,In_944,In_908);
nand U2895 (N_2895,In_826,In_721);
or U2896 (N_2896,In_448,In_1475);
nor U2897 (N_2897,In_1456,In_958);
or U2898 (N_2898,In_849,In_1377);
and U2899 (N_2899,In_959,In_617);
xnor U2900 (N_2900,In_773,In_1244);
xor U2901 (N_2901,In_446,In_1018);
nor U2902 (N_2902,In_1190,In_270);
and U2903 (N_2903,In_460,In_1128);
nand U2904 (N_2904,In_617,In_38);
nand U2905 (N_2905,In_98,In_60);
xnor U2906 (N_2906,In_1055,In_876);
nor U2907 (N_2907,In_1208,In_314);
nor U2908 (N_2908,In_1239,In_1353);
nor U2909 (N_2909,In_399,In_661);
and U2910 (N_2910,In_358,In_1404);
and U2911 (N_2911,In_991,In_547);
xnor U2912 (N_2912,In_1225,In_287);
or U2913 (N_2913,In_87,In_1085);
nand U2914 (N_2914,In_1093,In_376);
nand U2915 (N_2915,In_1115,In_1005);
and U2916 (N_2916,In_878,In_1188);
nand U2917 (N_2917,In_541,In_580);
and U2918 (N_2918,In_982,In_1260);
nand U2919 (N_2919,In_1182,In_470);
nand U2920 (N_2920,In_1372,In_1223);
or U2921 (N_2921,In_849,In_968);
xnor U2922 (N_2922,In_914,In_920);
nand U2923 (N_2923,In_405,In_353);
nor U2924 (N_2924,In_4,In_548);
nor U2925 (N_2925,In_482,In_1067);
nand U2926 (N_2926,In_608,In_838);
xnor U2927 (N_2927,In_619,In_522);
nand U2928 (N_2928,In_1146,In_931);
nand U2929 (N_2929,In_1366,In_1242);
xnor U2930 (N_2930,In_1106,In_402);
and U2931 (N_2931,In_888,In_456);
and U2932 (N_2932,In_1381,In_1474);
nor U2933 (N_2933,In_1408,In_374);
nor U2934 (N_2934,In_347,In_45);
nand U2935 (N_2935,In_1036,In_715);
or U2936 (N_2936,In_13,In_1469);
or U2937 (N_2937,In_466,In_1154);
or U2938 (N_2938,In_1348,In_244);
nand U2939 (N_2939,In_678,In_248);
nor U2940 (N_2940,In_767,In_248);
or U2941 (N_2941,In_634,In_369);
or U2942 (N_2942,In_1120,In_512);
nand U2943 (N_2943,In_893,In_62);
nor U2944 (N_2944,In_737,In_566);
and U2945 (N_2945,In_929,In_720);
and U2946 (N_2946,In_143,In_895);
and U2947 (N_2947,In_1242,In_852);
and U2948 (N_2948,In_1379,In_926);
and U2949 (N_2949,In_323,In_608);
nor U2950 (N_2950,In_507,In_213);
nor U2951 (N_2951,In_166,In_890);
and U2952 (N_2952,In_793,In_41);
nand U2953 (N_2953,In_202,In_64);
nor U2954 (N_2954,In_299,In_878);
or U2955 (N_2955,In_311,In_1451);
and U2956 (N_2956,In_684,In_234);
nand U2957 (N_2957,In_1268,In_1015);
nand U2958 (N_2958,In_1177,In_1321);
or U2959 (N_2959,In_860,In_723);
nor U2960 (N_2960,In_1446,In_479);
and U2961 (N_2961,In_1302,In_1249);
nor U2962 (N_2962,In_27,In_184);
or U2963 (N_2963,In_923,In_100);
xnor U2964 (N_2964,In_155,In_117);
or U2965 (N_2965,In_553,In_1360);
or U2966 (N_2966,In_1149,In_1300);
xor U2967 (N_2967,In_1425,In_712);
and U2968 (N_2968,In_1259,In_160);
xor U2969 (N_2969,In_864,In_844);
xnor U2970 (N_2970,In_1156,In_653);
nand U2971 (N_2971,In_994,In_1403);
xnor U2972 (N_2972,In_1261,In_1197);
xnor U2973 (N_2973,In_696,In_523);
nor U2974 (N_2974,In_914,In_970);
xnor U2975 (N_2975,In_926,In_613);
nor U2976 (N_2976,In_979,In_1171);
xor U2977 (N_2977,In_1360,In_1419);
xnor U2978 (N_2978,In_568,In_582);
nor U2979 (N_2979,In_687,In_1332);
nor U2980 (N_2980,In_653,In_614);
and U2981 (N_2981,In_428,In_1419);
xor U2982 (N_2982,In_1175,In_457);
nand U2983 (N_2983,In_1119,In_1423);
xnor U2984 (N_2984,In_145,In_177);
and U2985 (N_2985,In_1154,In_1188);
and U2986 (N_2986,In_1331,In_1155);
xor U2987 (N_2987,In_171,In_624);
nand U2988 (N_2988,In_963,In_1325);
nor U2989 (N_2989,In_1427,In_327);
or U2990 (N_2990,In_1036,In_388);
or U2991 (N_2991,In_556,In_1060);
nand U2992 (N_2992,In_49,In_164);
or U2993 (N_2993,In_1482,In_978);
and U2994 (N_2994,In_1042,In_228);
and U2995 (N_2995,In_976,In_1348);
or U2996 (N_2996,In_606,In_71);
xnor U2997 (N_2997,In_1364,In_1195);
and U2998 (N_2998,In_1297,In_1458);
nor U2999 (N_2999,In_882,In_1424);
and U3000 (N_3000,N_2792,N_1913);
or U3001 (N_3001,N_2776,N_1077);
nor U3002 (N_3002,N_1761,N_2213);
and U3003 (N_3003,N_975,N_463);
or U3004 (N_3004,N_2192,N_88);
nand U3005 (N_3005,N_2468,N_667);
nand U3006 (N_3006,N_1401,N_2483);
nor U3007 (N_3007,N_2104,N_1237);
or U3008 (N_3008,N_404,N_1208);
nor U3009 (N_3009,N_379,N_1267);
or U3010 (N_3010,N_1117,N_2357);
nand U3011 (N_3011,N_201,N_2867);
and U3012 (N_3012,N_1550,N_43);
and U3013 (N_3013,N_729,N_1317);
nand U3014 (N_3014,N_1386,N_1191);
nor U3015 (N_3015,N_550,N_1694);
nand U3016 (N_3016,N_693,N_332);
or U3017 (N_3017,N_1094,N_2131);
xnor U3018 (N_3018,N_1434,N_10);
nor U3019 (N_3019,N_1882,N_245);
nor U3020 (N_3020,N_1,N_665);
or U3021 (N_3021,N_1491,N_310);
nand U3022 (N_3022,N_103,N_2020);
nor U3023 (N_3023,N_584,N_1081);
nand U3024 (N_3024,N_1044,N_1345);
or U3025 (N_3025,N_1417,N_2610);
nand U3026 (N_3026,N_779,N_1514);
nand U3027 (N_3027,N_2177,N_2287);
nor U3028 (N_3028,N_1259,N_2616);
nor U3029 (N_3029,N_2773,N_1742);
nand U3030 (N_3030,N_396,N_2607);
xor U3031 (N_3031,N_2377,N_373);
nand U3032 (N_3032,N_1214,N_152);
and U3033 (N_3033,N_2390,N_980);
nand U3034 (N_3034,N_48,N_1126);
nor U3035 (N_3035,N_978,N_1704);
or U3036 (N_3036,N_1226,N_1034);
or U3037 (N_3037,N_2032,N_326);
xnor U3038 (N_3038,N_2319,N_41);
xnor U3039 (N_3039,N_520,N_1458);
or U3040 (N_3040,N_9,N_1294);
or U3041 (N_3041,N_1529,N_1561);
or U3042 (N_3042,N_1552,N_987);
nand U3043 (N_3043,N_1978,N_1653);
or U3044 (N_3044,N_151,N_2623);
or U3045 (N_3045,N_1860,N_1925);
nand U3046 (N_3046,N_1994,N_2183);
nor U3047 (N_3047,N_1114,N_1996);
nand U3048 (N_3048,N_2138,N_1712);
nor U3049 (N_3049,N_285,N_2642);
xor U3050 (N_3050,N_75,N_652);
or U3051 (N_3051,N_514,N_715);
nor U3052 (N_3052,N_2026,N_2393);
or U3053 (N_3053,N_2612,N_2304);
and U3054 (N_3054,N_440,N_2105);
nand U3055 (N_3055,N_25,N_1227);
nor U3056 (N_3056,N_1961,N_1176);
nand U3057 (N_3057,N_2807,N_2202);
and U3058 (N_3058,N_1505,N_734);
nor U3059 (N_3059,N_2939,N_1954);
nand U3060 (N_3060,N_231,N_624);
or U3061 (N_3061,N_637,N_2808);
nor U3062 (N_3062,N_1406,N_216);
or U3063 (N_3063,N_568,N_607);
nand U3064 (N_3064,N_117,N_498);
nand U3065 (N_3065,N_650,N_1664);
nor U3066 (N_3066,N_2200,N_1749);
or U3067 (N_3067,N_757,N_2651);
xor U3068 (N_3068,N_1698,N_1384);
xor U3069 (N_3069,N_2122,N_179);
and U3070 (N_3070,N_710,N_2386);
nor U3071 (N_3071,N_2566,N_2619);
nor U3072 (N_3072,N_909,N_2660);
nand U3073 (N_3073,N_2342,N_2333);
and U3074 (N_3074,N_2235,N_730);
nor U3075 (N_3075,N_1970,N_130);
nor U3076 (N_3076,N_1883,N_1006);
or U3077 (N_3077,N_1171,N_1919);
xor U3078 (N_3078,N_1839,N_673);
nor U3079 (N_3079,N_1437,N_496);
and U3080 (N_3080,N_712,N_1671);
nor U3081 (N_3081,N_106,N_572);
or U3082 (N_3082,N_2355,N_2910);
nor U3083 (N_3083,N_907,N_165);
nor U3084 (N_3084,N_1893,N_1484);
and U3085 (N_3085,N_811,N_132);
and U3086 (N_3086,N_1667,N_2930);
or U3087 (N_3087,N_686,N_586);
and U3088 (N_3088,N_588,N_2023);
nand U3089 (N_3089,N_721,N_1692);
and U3090 (N_3090,N_603,N_1197);
nand U3091 (N_3091,N_2258,N_806);
or U3092 (N_3092,N_2132,N_1119);
nor U3093 (N_3093,N_2313,N_1974);
nor U3094 (N_3094,N_1891,N_2339);
nor U3095 (N_3095,N_597,N_2749);
or U3096 (N_3096,N_2549,N_1292);
and U3097 (N_3097,N_388,N_324);
and U3098 (N_3098,N_1270,N_2753);
nor U3099 (N_3099,N_1503,N_731);
and U3100 (N_3100,N_1788,N_803);
and U3101 (N_3101,N_325,N_1181);
and U3102 (N_3102,N_834,N_1307);
and U3103 (N_3103,N_2031,N_574);
and U3104 (N_3104,N_489,N_1390);
nor U3105 (N_3105,N_782,N_1768);
and U3106 (N_3106,N_206,N_1516);
nand U3107 (N_3107,N_2362,N_552);
nor U3108 (N_3108,N_1313,N_1474);
and U3109 (N_3109,N_2412,N_1282);
or U3110 (N_3110,N_415,N_1007);
or U3111 (N_3111,N_2346,N_1449);
nand U3112 (N_3112,N_794,N_2530);
nand U3113 (N_3113,N_456,N_2556);
nand U3114 (N_3114,N_2949,N_27);
nor U3115 (N_3115,N_649,N_2225);
and U3116 (N_3116,N_738,N_73);
nand U3117 (N_3117,N_1154,N_292);
or U3118 (N_3118,N_128,N_2863);
nand U3119 (N_3119,N_2107,N_1859);
nor U3120 (N_3120,N_242,N_2300);
nor U3121 (N_3121,N_2990,N_911);
xnor U3122 (N_3122,N_2812,N_1563);
or U3123 (N_3123,N_2065,N_2272);
xor U3124 (N_3124,N_2006,N_1492);
or U3125 (N_3125,N_2028,N_958);
nand U3126 (N_3126,N_2312,N_833);
and U3127 (N_3127,N_2019,N_1543);
and U3128 (N_3128,N_2204,N_977);
nor U3129 (N_3129,N_2986,N_2325);
nor U3130 (N_3130,N_2034,N_1689);
and U3131 (N_3131,N_348,N_1151);
and U3132 (N_3132,N_1220,N_2963);
nand U3133 (N_3133,N_1235,N_2680);
and U3134 (N_3134,N_1400,N_2975);
or U3135 (N_3135,N_2080,N_695);
and U3136 (N_3136,N_1097,N_1857);
or U3137 (N_3137,N_2926,N_1337);
nor U3138 (N_3138,N_2781,N_2292);
and U3139 (N_3139,N_390,N_2759);
or U3140 (N_3140,N_995,N_1146);
nand U3141 (N_3141,N_1990,N_2653);
nor U3142 (N_3142,N_2274,N_976);
or U3143 (N_3143,N_2622,N_2162);
xnor U3144 (N_3144,N_2182,N_2500);
or U3145 (N_3145,N_2538,N_2259);
nand U3146 (N_3146,N_1129,N_294);
nand U3147 (N_3147,N_799,N_2700);
xor U3148 (N_3148,N_688,N_792);
or U3149 (N_3149,N_470,N_1187);
xnor U3150 (N_3150,N_2324,N_1914);
xnor U3151 (N_3151,N_2314,N_2553);
nand U3152 (N_3152,N_2550,N_110);
nor U3153 (N_3153,N_2181,N_426);
xnor U3154 (N_3154,N_2253,N_1054);
xnor U3155 (N_3155,N_2209,N_964);
nor U3156 (N_3156,N_1037,N_2852);
and U3157 (N_3157,N_596,N_2659);
or U3158 (N_3158,N_1777,N_696);
and U3159 (N_3159,N_1311,N_1479);
and U3160 (N_3160,N_662,N_1904);
and U3161 (N_3161,N_2371,N_1623);
nand U3162 (N_3162,N_2465,N_2826);
nor U3163 (N_3163,N_272,N_2726);
or U3164 (N_3164,N_2137,N_2351);
nor U3165 (N_3165,N_1085,N_114);
xor U3166 (N_3166,N_532,N_1161);
and U3167 (N_3167,N_232,N_2350);
and U3168 (N_3168,N_2343,N_756);
or U3169 (N_3169,N_1240,N_1295);
or U3170 (N_3170,N_2721,N_98);
nand U3171 (N_3171,N_1971,N_2109);
nor U3172 (N_3172,N_579,N_626);
nand U3173 (N_3173,N_2524,N_1116);
and U3174 (N_3174,N_716,N_1879);
nor U3175 (N_3175,N_248,N_2017);
or U3176 (N_3176,N_1663,N_2279);
or U3177 (N_3177,N_663,N_2890);
and U3178 (N_3178,N_931,N_990);
xor U3179 (N_3179,N_1786,N_1394);
xnor U3180 (N_3180,N_1473,N_2282);
nor U3181 (N_3181,N_253,N_1293);
xor U3182 (N_3182,N_1759,N_2447);
and U3183 (N_3183,N_1269,N_2521);
and U3184 (N_3184,N_68,N_1876);
and U3185 (N_3185,N_2811,N_764);
and U3186 (N_3186,N_2143,N_1321);
nor U3187 (N_3187,N_2932,N_2048);
xnor U3188 (N_3188,N_2563,N_2203);
nand U3189 (N_3189,N_1784,N_1090);
nor U3190 (N_3190,N_2909,N_1275);
or U3191 (N_3191,N_2806,N_2148);
nand U3192 (N_3192,N_2389,N_303);
or U3193 (N_3193,N_1011,N_2264);
or U3194 (N_3194,N_2596,N_2384);
xnor U3195 (N_3195,N_2038,N_955);
nand U3196 (N_3196,N_2636,N_1066);
or U3197 (N_3197,N_647,N_2505);
or U3198 (N_3198,N_1620,N_2845);
xor U3199 (N_3199,N_869,N_807);
or U3200 (N_3200,N_2956,N_462);
or U3201 (N_3201,N_1682,N_518);
xnor U3202 (N_3202,N_2410,N_2309);
and U3203 (N_3203,N_2617,N_2071);
nand U3204 (N_3204,N_2102,N_2268);
nand U3205 (N_3205,N_2373,N_1602);
nand U3206 (N_3206,N_815,N_2914);
or U3207 (N_3207,N_276,N_2905);
nand U3208 (N_3208,N_741,N_1842);
and U3209 (N_3209,N_356,N_1091);
and U3210 (N_3210,N_944,N_2992);
or U3211 (N_3211,N_2560,N_1053);
and U3212 (N_3212,N_670,N_849);
nand U3213 (N_3213,N_1840,N_1725);
or U3214 (N_3214,N_2180,N_1245);
nor U3215 (N_3215,N_1523,N_494);
or U3216 (N_3216,N_2385,N_347);
and U3217 (N_3217,N_4,N_1142);
and U3218 (N_3218,N_761,N_2398);
xnor U3219 (N_3219,N_954,N_2174);
and U3220 (N_3220,N_2545,N_2403);
and U3221 (N_3221,N_30,N_77);
or U3222 (N_3222,N_2778,N_2451);
nand U3223 (N_3223,N_2087,N_2882);
nor U3224 (N_3224,N_2218,N_2561);
or U3225 (N_3225,N_2825,N_2349);
nor U3226 (N_3226,N_1265,N_578);
nand U3227 (N_3227,N_1506,N_1729);
nor U3228 (N_3228,N_2654,N_541);
nor U3229 (N_3229,N_2823,N_2720);
or U3230 (N_3230,N_2564,N_1170);
nor U3231 (N_3231,N_2190,N_21);
nor U3232 (N_3232,N_602,N_1822);
and U3233 (N_3233,N_2918,N_992);
nor U3234 (N_3234,N_1192,N_1388);
nand U3235 (N_3235,N_1419,N_1195);
and U3236 (N_3236,N_2511,N_2704);
and U3237 (N_3237,N_2070,N_1120);
nand U3238 (N_3238,N_2775,N_2069);
or U3239 (N_3239,N_832,N_927);
and U3240 (N_3240,N_2924,N_1019);
nand U3241 (N_3241,N_858,N_2537);
or U3242 (N_3242,N_1105,N_1530);
and U3243 (N_3243,N_170,N_2730);
nand U3244 (N_3244,N_448,N_923);
and U3245 (N_3245,N_1708,N_824);
or U3246 (N_3246,N_1180,N_2499);
nand U3247 (N_3247,N_1456,N_1363);
and U3248 (N_3248,N_2944,N_280);
and U3249 (N_3249,N_2941,N_508);
nand U3250 (N_3250,N_1643,N_2551);
and U3251 (N_3251,N_372,N_2922);
or U3252 (N_3252,N_723,N_559);
and U3253 (N_3253,N_1415,N_1014);
and U3254 (N_3254,N_1222,N_1832);
nand U3255 (N_3255,N_1215,N_2599);
nor U3256 (N_3256,N_1249,N_1209);
nor U3257 (N_3257,N_2121,N_1817);
or U3258 (N_3258,N_2779,N_2078);
xnor U3259 (N_3259,N_826,N_2671);
nor U3260 (N_3260,N_478,N_589);
and U3261 (N_3261,N_2645,N_2630);
and U3262 (N_3262,N_2488,N_2237);
nor U3263 (N_3263,N_1442,N_1763);
and U3264 (N_3264,N_2340,N_1507);
and U3265 (N_3265,N_1823,N_1398);
and U3266 (N_3266,N_2461,N_742);
nor U3267 (N_3267,N_1816,N_1113);
or U3268 (N_3268,N_29,N_2581);
nor U3269 (N_3269,N_2687,N_1421);
nor U3270 (N_3270,N_862,N_1397);
nor U3271 (N_3271,N_1695,N_1225);
nand U3272 (N_3272,N_2146,N_1795);
or U3273 (N_3273,N_2883,N_989);
or U3274 (N_3274,N_235,N_91);
nor U3275 (N_3275,N_2358,N_264);
and U3276 (N_3276,N_2788,N_2802);
nand U3277 (N_3277,N_1940,N_2576);
nand U3278 (N_3278,N_1894,N_1939);
and U3279 (N_3279,N_2853,N_1646);
and U3280 (N_3280,N_59,N_1610);
xor U3281 (N_3281,N_984,N_13);
and U3282 (N_3282,N_1067,N_904);
xor U3283 (N_3283,N_1128,N_1869);
nand U3284 (N_3284,N_2529,N_367);
and U3285 (N_3285,N_1622,N_2647);
nand U3286 (N_3286,N_2372,N_2805);
nand U3287 (N_3287,N_1338,N_2929);
nor U3288 (N_3288,N_1736,N_2232);
nand U3289 (N_3289,N_1501,N_2027);
nor U3290 (N_3290,N_429,N_2846);
and U3291 (N_3291,N_2409,N_2419);
nor U3292 (N_3292,N_2803,N_770);
nand U3293 (N_3293,N_2793,N_2089);
nand U3294 (N_3294,N_1319,N_1892);
or U3295 (N_3295,N_1774,N_47);
nand U3296 (N_3296,N_1821,N_1329);
and U3297 (N_3297,N_2436,N_1854);
nand U3298 (N_3298,N_2794,N_2029);
or U3299 (N_3299,N_79,N_296);
or U3300 (N_3300,N_107,N_2201);
nor U3301 (N_3301,N_2620,N_1030);
or U3302 (N_3302,N_2049,N_1253);
xor U3303 (N_3303,N_1548,N_610);
nand U3304 (N_3304,N_871,N_570);
nand U3305 (N_3305,N_630,N_172);
or U3306 (N_3306,N_1280,N_320);
or U3307 (N_3307,N_772,N_786);
xnor U3308 (N_3308,N_1613,N_1581);
and U3309 (N_3309,N_2081,N_1322);
nor U3310 (N_3310,N_2597,N_2248);
and U3311 (N_3311,N_1848,N_1304);
nand U3312 (N_3312,N_1800,N_156);
nand U3313 (N_3313,N_1865,N_1193);
nand U3314 (N_3314,N_2719,N_2379);
and U3315 (N_3315,N_671,N_1660);
nor U3316 (N_3316,N_2809,N_2227);
or U3317 (N_3317,N_1027,N_554);
and U3318 (N_3318,N_479,N_875);
or U3319 (N_3319,N_1685,N_1934);
nand U3320 (N_3320,N_471,N_386);
nor U3321 (N_3321,N_2217,N_1109);
nor U3322 (N_3322,N_1219,N_2943);
or U3323 (N_3323,N_2439,N_1099);
nand U3324 (N_3324,N_979,N_1794);
nand U3325 (N_3325,N_2051,N_654);
and U3326 (N_3326,N_2737,N_2934);
or U3327 (N_3327,N_2578,N_2067);
or U3328 (N_3328,N_328,N_1179);
xnor U3329 (N_3329,N_2959,N_1462);
and U3330 (N_3330,N_2763,N_1864);
or U3331 (N_3331,N_873,N_2250);
nand U3332 (N_3332,N_2835,N_19);
nand U3333 (N_3333,N_2681,N_1573);
nand U3334 (N_3334,N_583,N_2176);
and U3335 (N_3335,N_382,N_896);
and U3336 (N_3336,N_135,N_22);
and U3337 (N_3337,N_2902,N_1058);
nor U3338 (N_3338,N_1976,N_1315);
or U3339 (N_3339,N_1031,N_1804);
xor U3340 (N_3340,N_115,N_736);
nor U3341 (N_3341,N_436,N_171);
and U3342 (N_3342,N_1785,N_1519);
or U3343 (N_3343,N_1787,N_1050);
nand U3344 (N_3344,N_2613,N_1183);
nor U3345 (N_3345,N_1103,N_116);
or U3346 (N_3346,N_141,N_2718);
nor U3347 (N_3347,N_1178,N_2432);
nor U3348 (N_3348,N_606,N_427);
nand U3349 (N_3349,N_2236,N_1448);
nand U3350 (N_3350,N_655,N_2459);
nor U3351 (N_3351,N_1165,N_1847);
and U3352 (N_3352,N_1201,N_2593);
nand U3353 (N_3353,N_2600,N_2090);
nor U3354 (N_3354,N_1782,N_898);
nor U3355 (N_3355,N_1837,N_2856);
nor U3356 (N_3356,N_2205,N_2366);
or U3357 (N_3357,N_2869,N_2925);
and U3358 (N_3358,N_881,N_2050);
or U3359 (N_3359,N_2820,N_2762);
nor U3360 (N_3360,N_1895,N_1347);
nor U3361 (N_3361,N_2044,N_1436);
nand U3362 (N_3362,N_2285,N_1039);
nand U3363 (N_3363,N_2053,N_785);
nand U3364 (N_3364,N_2037,N_2711);
nand U3365 (N_3365,N_2828,N_938);
or U3366 (N_3366,N_380,N_2668);
nor U3367 (N_3367,N_1086,N_1843);
and U3368 (N_3368,N_2927,N_1808);
nand U3369 (N_3369,N_2106,N_2618);
or U3370 (N_3370,N_1987,N_1182);
nand U3371 (N_3371,N_2969,N_2117);
nand U3372 (N_3372,N_1164,N_2850);
nand U3373 (N_3373,N_2077,N_2627);
or U3374 (N_3374,N_2662,N_947);
nor U3375 (N_3375,N_2145,N_309);
nor U3376 (N_3376,N_525,N_1809);
xnor U3377 (N_3377,N_67,N_1983);
xor U3378 (N_3378,N_771,N_316);
and U3379 (N_3379,N_2494,N_594);
and U3380 (N_3380,N_194,N_651);
or U3381 (N_3381,N_2994,N_2197);
and U3382 (N_3382,N_2518,N_2637);
and U3383 (N_3383,N_2507,N_1029);
nor U3384 (N_3384,N_2004,N_1403);
and U3385 (N_3385,N_1268,N_2900);
and U3386 (N_3386,N_1657,N_55);
and U3387 (N_3387,N_965,N_1829);
nor U3388 (N_3388,N_2097,N_2516);
nand U3389 (N_3389,N_474,N_523);
nand U3390 (N_3390,N_1377,N_717);
nor U3391 (N_3391,N_2405,N_1078);
or U3392 (N_3392,N_368,N_277);
nor U3393 (N_3393,N_2689,N_1416);
xnor U3394 (N_3394,N_2378,N_1494);
nand U3395 (N_3395,N_677,N_1977);
and U3396 (N_3396,N_2207,N_2359);
or U3397 (N_3397,N_691,N_1022);
and U3398 (N_3398,N_2764,N_2303);
and U3399 (N_3399,N_2723,N_725);
xor U3400 (N_3400,N_1323,N_2634);
nand U3401 (N_3401,N_2635,N_1867);
nor U3402 (N_3402,N_119,N_244);
or U3403 (N_3403,N_51,N_1720);
nor U3404 (N_3404,N_2508,N_713);
nor U3405 (N_3405,N_2532,N_1647);
and U3406 (N_3406,N_2515,N_1825);
and U3407 (N_3407,N_2134,N_374);
nor U3408 (N_3408,N_839,N_2254);
and U3409 (N_3409,N_70,N_816);
nor U3410 (N_3410,N_2785,N_391);
xor U3411 (N_3411,N_1609,N_1049);
nand U3412 (N_3412,N_378,N_1851);
nand U3413 (N_3413,N_1359,N_2387);
and U3414 (N_3414,N_1827,N_1969);
and U3415 (N_3415,N_24,N_790);
xnor U3416 (N_3416,N_1630,N_1818);
nor U3417 (N_3417,N_519,N_2194);
or U3418 (N_3418,N_2942,N_780);
or U3419 (N_3419,N_2684,N_1953);
xnor U3420 (N_3420,N_351,N_1365);
and U3421 (N_3421,N_2040,N_1607);
or U3422 (N_3422,N_1508,N_416);
nand U3423 (N_3423,N_2230,N_1688);
or U3424 (N_3424,N_1157,N_1497);
nor U3425 (N_3425,N_561,N_2945);
or U3426 (N_3426,N_377,N_533);
and U3427 (N_3427,N_2454,N_1735);
xnor U3428 (N_3428,N_184,N_345);
nand U3429 (N_3429,N_1341,N_167);
nor U3430 (N_3430,N_961,N_1637);
or U3431 (N_3431,N_823,N_2256);
and U3432 (N_3432,N_611,N_1551);
xnor U3433 (N_3433,N_953,N_181);
and U3434 (N_3434,N_551,N_2961);
xnor U3435 (N_3435,N_2695,N_1465);
and U3436 (N_3436,N_2283,N_2045);
or U3437 (N_3437,N_2527,N_361);
or U3438 (N_3438,N_2736,N_92);
nor U3439 (N_3439,N_2712,N_1445);
nand U3440 (N_3440,N_732,N_2897);
or U3441 (N_3441,N_1706,N_83);
and U3442 (N_3442,N_1412,N_510);
and U3443 (N_3443,N_720,N_2703);
or U3444 (N_3444,N_1264,N_2673);
nand U3445 (N_3445,N_1528,N_2815);
or U3446 (N_3446,N_2471,N_1095);
or U3447 (N_3447,N_2861,N_1263);
nor U3448 (N_3448,N_1746,N_497);
or U3449 (N_3449,N_452,N_2173);
and U3450 (N_3450,N_1107,N_183);
nor U3451 (N_3451,N_2495,N_1999);
nor U3452 (N_3452,N_1927,N_219);
xor U3453 (N_3453,N_2790,N_1950);
or U3454 (N_3454,N_1233,N_2172);
or U3455 (N_3455,N_1443,N_1881);
and U3456 (N_3456,N_2933,N_2091);
or U3457 (N_3457,N_1318,N_1525);
and U3458 (N_3458,N_1918,N_690);
and U3459 (N_3459,N_2082,N_2166);
nor U3460 (N_3460,N_2000,N_2898);
or U3461 (N_3461,N_1967,N_701);
and U3462 (N_3462,N_121,N_1320);
nor U3463 (N_3463,N_1510,N_1680);
nand U3464 (N_3464,N_445,N_53);
or U3465 (N_3465,N_461,N_2559);
nand U3466 (N_3466,N_2033,N_1877);
nor U3467 (N_3467,N_1335,N_421);
nor U3468 (N_3468,N_922,N_100);
xnor U3469 (N_3469,N_1130,N_1177);
nand U3470 (N_3470,N_2851,N_2874);
or U3471 (N_3471,N_1162,N_405);
nand U3472 (N_3472,N_1100,N_1684);
xnor U3473 (N_3473,N_1721,N_1303);
nor U3474 (N_3474,N_2998,N_2601);
and U3475 (N_3475,N_1061,N_2609);
or U3476 (N_3476,N_2239,N_1943);
nor U3477 (N_3477,N_143,N_2421);
nand U3478 (N_3478,N_1174,N_1762);
nand U3479 (N_3479,N_2155,N_1046);
nor U3480 (N_3480,N_1679,N_1228);
nand U3481 (N_3481,N_2725,N_861);
nand U3482 (N_3482,N_2936,N_414);
or U3483 (N_3483,N_1727,N_2984);
nor U3484 (N_3484,N_2976,N_2114);
nor U3485 (N_3485,N_2799,N_2135);
nand U3486 (N_3486,N_2140,N_1380);
nor U3487 (N_3487,N_1973,N_2126);
and U3488 (N_3488,N_1717,N_941);
nand U3489 (N_3489,N_1702,N_1642);
nand U3490 (N_3490,N_65,N_2679);
and U3491 (N_3491,N_166,N_2887);
or U3492 (N_3492,N_164,N_2179);
and U3493 (N_3493,N_2442,N_2013);
and U3494 (N_3494,N_1661,N_1141);
nand U3495 (N_3495,N_548,N_895);
nor U3496 (N_3496,N_180,N_1739);
and U3497 (N_3497,N_370,N_1210);
nand U3498 (N_3498,N_1570,N_2093);
nor U3499 (N_3499,N_521,N_215);
and U3500 (N_3500,N_534,N_318);
and U3501 (N_3501,N_15,N_666);
and U3502 (N_3502,N_2294,N_962);
nor U3503 (N_3503,N_2025,N_221);
and U3504 (N_3504,N_1554,N_854);
and U3505 (N_3505,N_2548,N_1744);
nand U3506 (N_3506,N_2813,N_199);
nand U3507 (N_3507,N_2257,N_2568);
or U3508 (N_3508,N_1715,N_581);
and U3509 (N_3509,N_2643,N_2913);
nor U3510 (N_3510,N_1101,N_2535);
nand U3511 (N_3511,N_754,N_789);
nor U3512 (N_3512,N_2231,N_2780);
nand U3513 (N_3513,N_1896,N_261);
xnor U3514 (N_3514,N_2587,N_1687);
nor U3515 (N_3515,N_2021,N_2487);
nor U3516 (N_3516,N_1047,N_2450);
nand U3517 (N_3517,N_336,N_1989);
or U3518 (N_3518,N_360,N_1025);
xnor U3519 (N_3519,N_40,N_887);
nor U3520 (N_3520,N_1344,N_457);
nand U3521 (N_3521,N_1781,N_2249);
or U3522 (N_3522,N_2472,N_2347);
and U3523 (N_3523,N_2269,N_2191);
and U3524 (N_3524,N_2769,N_84);
and U3525 (N_3525,N_491,N_2407);
or U3526 (N_3526,N_266,N_2088);
and U3527 (N_3527,N_1797,N_2640);
xor U3528 (N_3528,N_1542,N_999);
nor U3529 (N_3529,N_255,N_997);
and U3530 (N_3530,N_870,N_442);
xnor U3531 (N_3531,N_1104,N_1083);
and U3532 (N_3532,N_2397,N_56);
and U3533 (N_3533,N_2591,N_2115);
and U3534 (N_3534,N_250,N_1522);
nand U3535 (N_3535,N_1668,N_2540);
and U3536 (N_3536,N_233,N_1121);
xnor U3537 (N_3537,N_446,N_1982);
and U3538 (N_3538,N_1862,N_1284);
or U3539 (N_3539,N_1490,N_1743);
xor U3540 (N_3540,N_1756,N_643);
and U3541 (N_3541,N_2076,N_1080);
xnor U3542 (N_3542,N_94,N_1964);
nor U3543 (N_3543,N_2360,N_1908);
and U3544 (N_3544,N_2818,N_1051);
nand U3545 (N_3545,N_1790,N_565);
nor U3546 (N_3546,N_350,N_105);
or U3547 (N_3547,N_1952,N_2188);
nand U3548 (N_3548,N_2784,N_1957);
nor U3549 (N_3549,N_1231,N_2127);
nand U3550 (N_3550,N_575,N_7);
and U3551 (N_3551,N_1984,N_2655);
nand U3552 (N_3552,N_2894,N_2699);
and U3553 (N_3553,N_2101,N_126);
and U3554 (N_3554,N_1381,N_1457);
nor U3555 (N_3555,N_2767,N_1951);
xor U3556 (N_3556,N_459,N_587);
nand U3557 (N_3557,N_993,N_591);
nand U3558 (N_3558,N_1980,N_1873);
nor U3559 (N_3559,N_297,N_2951);
xnor U3560 (N_3560,N_2672,N_1127);
nand U3561 (N_3561,N_797,N_127);
or U3562 (N_3562,N_1909,N_2099);
and U3563 (N_3563,N_2880,N_852);
xnor U3564 (N_3564,N_749,N_983);
nand U3565 (N_3565,N_1468,N_1169);
and U3566 (N_3566,N_1159,N_1758);
xnor U3567 (N_3567,N_443,N_507);
nand U3568 (N_3568,N_2460,N_1733);
and U3569 (N_3569,N_886,N_423);
or U3570 (N_3570,N_835,N_1470);
nor U3571 (N_3571,N_252,N_719);
nand U3572 (N_3572,N_2042,N_1301);
nand U3573 (N_3573,N_675,N_813);
xnor U3574 (N_3574,N_1572,N_2931);
xor U3575 (N_3575,N_1418,N_2834);
nor U3576 (N_3576,N_134,N_218);
xnor U3577 (N_3577,N_1813,N_1929);
nand U3578 (N_3578,N_441,N_1238);
or U3579 (N_3579,N_1619,N_1897);
or U3580 (N_3580,N_466,N_2585);
and U3581 (N_3581,N_744,N_2878);
nor U3582 (N_3582,N_915,N_564);
or U3583 (N_3583,N_1521,N_1057);
and U3584 (N_3584,N_1544,N_16);
or U3585 (N_3585,N_631,N_737);
nand U3586 (N_3586,N_475,N_2960);
and U3587 (N_3587,N_2810,N_1453);
xnor U3588 (N_3588,N_1844,N_275);
or U3589 (N_3589,N_473,N_113);
nand U3590 (N_3590,N_817,N_1439);
or U3591 (N_3591,N_2710,N_2586);
nor U3592 (N_3592,N_1132,N_2382);
xor U3593 (N_3593,N_808,N_1093);
nand U3594 (N_3594,N_1331,N_411);
and U3595 (N_3595,N_1584,N_1524);
and U3596 (N_3596,N_2353,N_480);
nand U3597 (N_3597,N_2525,N_2433);
nand U3598 (N_3598,N_1975,N_949);
xor U3599 (N_3599,N_573,N_2638);
and U3600 (N_3600,N_364,N_1615);
nand U3601 (N_3601,N_1010,N_851);
or U3602 (N_3602,N_1965,N_1515);
and U3603 (N_3603,N_2891,N_299);
nor U3604 (N_3604,N_2463,N_2571);
or U3605 (N_3605,N_2443,N_2404);
or U3606 (N_3606,N_2141,N_211);
or U3607 (N_3607,N_1750,N_2693);
nor U3608 (N_3608,N_281,N_1599);
nor U3609 (N_3609,N_493,N_971);
nand U3610 (N_3610,N_2701,N_967);
or U3611 (N_3611,N_659,N_1591);
or U3612 (N_3612,N_1367,N_1310);
nor U3613 (N_3613,N_900,N_2946);
or U3614 (N_3614,N_136,N_538);
nand U3615 (N_3615,N_270,N_2838);
and U3616 (N_3616,N_2787,N_504);
nor U3617 (N_3617,N_1741,N_1811);
nand U3618 (N_3618,N_767,N_2302);
or U3619 (N_3619,N_2244,N_1020);
nor U3620 (N_3620,N_1636,N_1261);
xnor U3621 (N_3621,N_2993,N_2967);
and U3622 (N_3622,N_1947,N_490);
nor U3623 (N_3623,N_502,N_1446);
nand U3624 (N_3624,N_842,N_334);
nand U3625 (N_3625,N_506,N_1213);
or U3626 (N_3626,N_1922,N_728);
nor U3627 (N_3627,N_481,N_1728);
nor U3628 (N_3628,N_524,N_674);
and U3629 (N_3629,N_108,N_2697);
nor U3630 (N_3630,N_1305,N_2458);
nor U3631 (N_3631,N_1773,N_2241);
nand U3632 (N_3632,N_2667,N_2770);
or U3633 (N_3633,N_1353,N_61);
and U3634 (N_3634,N_1730,N_894);
and U3635 (N_3635,N_1370,N_2896);
nand U3636 (N_3636,N_535,N_424);
and U3637 (N_3637,N_542,N_668);
or U3638 (N_3638,N_801,N_1273);
nand U3639 (N_3639,N_760,N_672);
or U3640 (N_3640,N_2683,N_1537);
or U3641 (N_3641,N_403,N_1407);
and U3642 (N_3642,N_2706,N_2441);
or U3643 (N_3643,N_286,N_1194);
or U3644 (N_3644,N_1500,N_1472);
nand U3645 (N_3645,N_981,N_289);
xnor U3646 (N_3646,N_2830,N_2819);
nor U3647 (N_3647,N_1941,N_890);
or U3648 (N_3648,N_1845,N_2058);
and U3649 (N_3649,N_766,N_2394);
xnor U3650 (N_3650,N_145,N_1082);
and U3651 (N_3651,N_1221,N_513);
and U3652 (N_3652,N_2344,N_2821);
nor U3653 (N_3653,N_2656,N_1834);
nand U3654 (N_3654,N_36,N_2452);
nor U3655 (N_3655,N_638,N_102);
nor U3656 (N_3656,N_985,N_2663);
xor U3657 (N_3657,N_2743,N_37);
or U3658 (N_3658,N_1673,N_1942);
or U3659 (N_3659,N_1766,N_1923);
nand U3660 (N_3660,N_2766,N_2957);
nor U3661 (N_3661,N_933,N_1131);
or U3662 (N_3662,N_1422,N_910);
nand U3663 (N_3663,N_2624,N_1198);
and U3664 (N_3664,N_148,N_1455);
and U3665 (N_3665,N_1569,N_2381);
nand U3666 (N_3666,N_1705,N_1556);
xor U3667 (N_3667,N_1004,N_109);
or U3668 (N_3668,N_2255,N_2334);
and U3669 (N_3669,N_2416,N_2427);
nand U3670 (N_3670,N_943,N_2513);
or U3671 (N_3671,N_1830,N_511);
xnor U3672 (N_3672,N_2187,N_2395);
nor U3673 (N_3673,N_889,N_2243);
nor U3674 (N_3674,N_762,N_2108);
and U3675 (N_3675,N_1791,N_1358);
xor U3676 (N_3676,N_1339,N_2708);
nand U3677 (N_3677,N_2455,N_1772);
and U3678 (N_3678,N_2073,N_1361);
or U3679 (N_3679,N_338,N_1475);
and U3680 (N_3680,N_1013,N_1651);
nor U3681 (N_3681,N_2167,N_2338);
nor U3682 (N_3682,N_454,N_422);
or U3683 (N_3683,N_841,N_139);
or U3684 (N_3684,N_2112,N_1134);
or U3685 (N_3685,N_2870,N_613);
nor U3686 (N_3686,N_1748,N_305);
and U3687 (N_3687,N_1924,N_614);
and U3688 (N_3688,N_419,N_2474);
or U3689 (N_3689,N_1775,N_2682);
and U3690 (N_3690,N_2030,N_1296);
or U3691 (N_3691,N_387,N_1861);
xor U3692 (N_3692,N_395,N_2804);
xor U3693 (N_3693,N_1932,N_1063);
nand U3694 (N_3694,N_257,N_2296);
or U3695 (N_3695,N_2440,N_138);
nand U3696 (N_3696,N_916,N_2356);
nand U3697 (N_3697,N_893,N_777);
nor U3698 (N_3698,N_2445,N_182);
or U3699 (N_3699,N_2128,N_540);
or U3700 (N_3700,N_2670,N_2731);
or U3701 (N_3701,N_62,N_74);
and U3702 (N_3702,N_2466,N_2657);
and U3703 (N_3703,N_246,N_884);
and U3704 (N_3704,N_2311,N_146);
and U3705 (N_3705,N_2839,N_1431);
and U3706 (N_3706,N_2506,N_1440);
nor U3707 (N_3707,N_2981,N_1652);
and U3708 (N_3708,N_1250,N_465);
nor U3709 (N_3709,N_2156,N_1122);
or U3710 (N_3710,N_1644,N_1435);
nand U3711 (N_3711,N_1517,N_2317);
xnor U3712 (N_3712,N_2310,N_2210);
or U3713 (N_3713,N_430,N_1481);
nand U3714 (N_3714,N_195,N_1287);
nand U3715 (N_3715,N_228,N_485);
nor U3716 (N_3716,N_1184,N_1806);
nor U3717 (N_3717,N_2795,N_2526);
and U3718 (N_3718,N_2648,N_2018);
xnor U3719 (N_3719,N_2938,N_1633);
xor U3720 (N_3720,N_1627,N_1017);
and U3721 (N_3721,N_2423,N_190);
nand U3722 (N_3722,N_2849,N_2417);
nor U3723 (N_3723,N_577,N_301);
or U3724 (N_3724,N_1731,N_2486);
nor U3725 (N_3725,N_1153,N_879);
nor U3726 (N_3726,N_1575,N_616);
nor U3727 (N_3727,N_2868,N_2367);
nor U3728 (N_3728,N_919,N_2276);
nor U3729 (N_3729,N_2301,N_2277);
or U3730 (N_3730,N_1541,N_63);
and U3731 (N_3731,N_827,N_1639);
nor U3732 (N_3732,N_72,N_2522);
and U3733 (N_3733,N_1598,N_1945);
nor U3734 (N_3734,N_776,N_2954);
or U3735 (N_3735,N_1369,N_2047);
nor U3736 (N_3736,N_271,N_1498);
nand U3737 (N_3737,N_365,N_1539);
nand U3738 (N_3738,N_49,N_1272);
nand U3739 (N_3739,N_1374,N_2980);
and U3740 (N_3740,N_45,N_394);
or U3741 (N_3741,N_447,N_2429);
and U3742 (N_3742,N_2165,N_1395);
and U3743 (N_3743,N_2212,N_708);
and U3744 (N_3744,N_1713,N_751);
or U3745 (N_3745,N_2872,N_2836);
nand U3746 (N_3746,N_1055,N_1589);
or U3747 (N_3747,N_288,N_393);
xor U3748 (N_3748,N_1678,N_2968);
and U3749 (N_3749,N_2614,N_1805);
xnor U3750 (N_3750,N_1223,N_580);
and U3751 (N_3751,N_623,N_1482);
nand U3752 (N_3752,N_1577,N_1110);
or U3753 (N_3753,N_435,N_1764);
and U3754 (N_3754,N_1357,N_1408);
xor U3755 (N_3755,N_408,N_1625);
or U3756 (N_3756,N_1340,N_2696);
or U3757 (N_3757,N_1349,N_2479);
nor U3758 (N_3758,N_35,N_204);
xnor U3759 (N_3759,N_2448,N_2265);
and U3760 (N_3760,N_1555,N_1710);
nor U3761 (N_3761,N_5,N_1681);
nor U3762 (N_3762,N_2641,N_2252);
nor U3763 (N_3763,N_645,N_2116);
or U3764 (N_3764,N_2374,N_2039);
nor U3765 (N_3765,N_2075,N_1216);
and U3766 (N_3766,N_2987,N_1944);
or U3767 (N_3767,N_304,N_2130);
xnor U3768 (N_3768,N_1535,N_2833);
nand U3769 (N_3769,N_337,N_400);
or U3770 (N_3770,N_2860,N_1696);
nand U3771 (N_3771,N_290,N_874);
nand U3772 (N_3772,N_1963,N_1059);
and U3773 (N_3773,N_28,N_223);
nand U3774 (N_3774,N_64,N_2698);
nand U3775 (N_3775,N_2298,N_1065);
xor U3776 (N_3776,N_2966,N_2273);
nand U3777 (N_3777,N_698,N_0);
nand U3778 (N_3778,N_2119,N_747);
nand U3779 (N_3779,N_2575,N_262);
nand U3780 (N_3780,N_2582,N_2685);
or U3781 (N_3781,N_627,N_208);
and U3782 (N_3782,N_1549,N_656);
or U3783 (N_3783,N_590,N_2555);
or U3784 (N_3784,N_2709,N_2903);
or U3785 (N_3785,N_1796,N_635);
nor U3786 (N_3786,N_1557,N_2741);
or U3787 (N_3787,N_973,N_1593);
and U3788 (N_3788,N_557,N_2573);
and U3789 (N_3789,N_484,N_558);
and U3790 (N_3790,N_1855,N_2798);
or U3791 (N_3791,N_144,N_1486);
nand U3792 (N_3792,N_2473,N_2580);
nand U3793 (N_3793,N_2206,N_389);
or U3794 (N_3794,N_2271,N_2251);
and U3795 (N_3795,N_371,N_85);
nor U3796 (N_3796,N_908,N_207);
nor U3797 (N_3797,N_1958,N_1385);
nand U3798 (N_3798,N_1425,N_302);
and U3799 (N_3799,N_2594,N_2738);
and U3800 (N_3800,N_1092,N_1424);
and U3801 (N_3801,N_2444,N_1089);
nor U3802 (N_3802,N_592,N_585);
and U3803 (N_3803,N_1592,N_86);
xnor U3804 (N_3804,N_185,N_1248);
and U3805 (N_3805,N_1670,N_2229);
or U3806 (N_3806,N_1376,N_1354);
nor U3807 (N_3807,N_1608,N_1450);
nand U3808 (N_3808,N_2746,N_791);
or U3809 (N_3809,N_1009,N_2777);
nor U3810 (N_3810,N_2536,N_2133);
and U3811 (N_3811,N_1789,N_2983);
nor U3812 (N_3812,N_3,N_2791);
or U3813 (N_3813,N_2392,N_694);
nor U3814 (N_3814,N_2348,N_169);
nand U3815 (N_3815,N_899,N_240);
and U3816 (N_3816,N_147,N_1564);
and U3817 (N_3817,N_2185,N_2036);
or U3818 (N_3818,N_1246,N_1915);
nor U3819 (N_3819,N_2608,N_2974);
nand U3820 (N_3820,N_308,N_1629);
and U3821 (N_3821,N_2418,N_1907);
nor U3822 (N_3822,N_154,N_1509);
and U3823 (N_3823,N_798,N_355);
or U3824 (N_3824,N_2060,N_1459);
nand U3825 (N_3825,N_176,N_2003);
nor U3826 (N_3826,N_2625,N_1931);
nor U3827 (N_3827,N_1167,N_1665);
or U3828 (N_3828,N_625,N_247);
or U3829 (N_3829,N_545,N_1447);
nand U3830 (N_3830,N_2503,N_549);
and U3831 (N_3831,N_2430,N_819);
nor U3832 (N_3832,N_1718,N_1278);
nor U3833 (N_3833,N_287,N_1526);
xor U3834 (N_3834,N_1068,N_1426);
nor U3835 (N_3835,N_2046,N_2965);
nand U3836 (N_3836,N_1124,N_2496);
nand U3837 (N_3837,N_291,N_788);
nand U3838 (N_3838,N_1106,N_937);
and U3839 (N_3839,N_640,N_1520);
nor U3840 (N_3840,N_998,N_2661);
and U3841 (N_3841,N_2072,N_986);
xnor U3842 (N_3842,N_8,N_2928);
and U3843 (N_3843,N_1737,N_2873);
nor U3844 (N_3844,N_2492,N_227);
nand U3845 (N_3845,N_256,N_1298);
and U3846 (N_3846,N_859,N_1023);
nor U3847 (N_3847,N_857,N_1738);
or U3848 (N_3848,N_243,N_2669);
or U3849 (N_3849,N_2329,N_970);
or U3850 (N_3850,N_563,N_1392);
nor U3851 (N_3851,N_1460,N_2912);
and U3852 (N_3852,N_1186,N_648);
and U3853 (N_3853,N_2074,N_709);
and U3854 (N_3854,N_1163,N_265);
or U3855 (N_3855,N_2125,N_1655);
xnor U3856 (N_3856,N_129,N_417);
nor U3857 (N_3857,N_1771,N_1088);
and U3858 (N_3858,N_1488,N_2602);
nor U3859 (N_3859,N_50,N_2011);
or U3860 (N_3860,N_409,N_2948);
and U3861 (N_3861,N_1512,N_2841);
and U3862 (N_3862,N_2514,N_1546);
or U3863 (N_3863,N_1326,N_2383);
nor U3864 (N_3864,N_925,N_2633);
nor U3865 (N_3865,N_339,N_1874);
and U3866 (N_3866,N_956,N_1991);
nor U3867 (N_3867,N_1560,N_653);
xor U3868 (N_3868,N_1346,N_1277);
nand U3869 (N_3869,N_178,N_1202);
nand U3870 (N_3870,N_1826,N_1658);
or U3871 (N_3871,N_865,N_768);
nand U3872 (N_3872,N_2562,N_936);
and U3873 (N_3873,N_2307,N_335);
nor U3874 (N_3874,N_173,N_89);
or U3875 (N_3875,N_2062,N_2691);
nand U3876 (N_3876,N_840,N_2152);
and U3877 (N_3877,N_547,N_2485);
nor U3878 (N_3878,N_526,N_2705);
nor U3879 (N_3879,N_2855,N_2840);
xnor U3880 (N_3880,N_1634,N_1478);
and U3881 (N_3881,N_658,N_2014);
xor U3882 (N_3882,N_1466,N_57);
nand U3883 (N_3883,N_1810,N_349);
nor U3884 (N_3884,N_2111,N_2884);
nand U3885 (N_3885,N_773,N_26);
and U3886 (N_3886,N_2985,N_2437);
and U3887 (N_3887,N_878,N_2895);
and U3888 (N_3888,N_2539,N_2323);
or U3889 (N_3889,N_1399,N_1314);
nor U3890 (N_3890,N_2677,N_1531);
nor U3891 (N_3891,N_500,N_2247);
nand U3892 (N_3892,N_926,N_2431);
xor U3893 (N_3893,N_76,N_901);
nor U3894 (N_3894,N_2541,N_112);
xnor U3895 (N_3895,N_2151,N_1594);
nor U3896 (N_3896,N_2915,N_1211);
and U3897 (N_3897,N_2426,N_1428);
xnor U3898 (N_3898,N_2543,N_2260);
or U3899 (N_3899,N_726,N_1880);
xor U3900 (N_3900,N_1906,N_876);
nand U3901 (N_3901,N_1477,N_2827);
nor U3902 (N_3902,N_2901,N_38);
nand U3903 (N_3903,N_1239,N_1714);
and U3904 (N_3904,N_2198,N_897);
and U3905 (N_3905,N_401,N_1645);
nor U3906 (N_3906,N_810,N_2354);
and U3907 (N_3907,N_1217,N_2714);
xor U3908 (N_3908,N_467,N_1898);
nand U3909 (N_3909,N_704,N_196);
and U3910 (N_3910,N_2646,N_2064);
or U3911 (N_3911,N_2226,N_2579);
and U3912 (N_3912,N_2401,N_1143);
and U3913 (N_3913,N_2605,N_1545);
nand U3914 (N_3914,N_1032,N_957);
and U3915 (N_3915,N_2920,N_2908);
nor U3916 (N_3916,N_14,N_1578);
or U3917 (N_3917,N_2246,N_537);
nor U3918 (N_3918,N_1621,N_1271);
or U3919 (N_3919,N_644,N_945);
nor U3920 (N_3920,N_1917,N_920);
and U3921 (N_3921,N_2475,N_2768);
nand U3922 (N_3922,N_2305,N_458);
xnor U3923 (N_3923,N_263,N_402);
nor U3924 (N_3924,N_198,N_2124);
nor U3925 (N_3925,N_2098,N_2824);
nand U3926 (N_3926,N_2278,N_793);
nand U3927 (N_3927,N_2085,N_2345);
and U3928 (N_3928,N_1356,N_1297);
and U3929 (N_3929,N_2024,N_2907);
nand U3930 (N_3930,N_137,N_2857);
nand U3931 (N_3931,N_2110,N_2295);
nor U3932 (N_3932,N_1875,N_913);
nor U3933 (N_3933,N_2100,N_855);
nor U3934 (N_3934,N_2005,N_1172);
and U3935 (N_3935,N_2724,N_1260);
or U3936 (N_3936,N_2223,N_2606);
xor U3937 (N_3937,N_353,N_2096);
xnor U3938 (N_3938,N_598,N_2542);
nand U3939 (N_3939,N_1045,N_2228);
or U3940 (N_3940,N_2158,N_2504);
nand U3941 (N_3941,N_399,N_2084);
or U3942 (N_3942,N_1935,N_492);
nor U3943 (N_3943,N_1224,N_118);
and U3944 (N_3944,N_1815,N_1624);
or U3945 (N_3945,N_2438,N_376);
nand U3946 (N_3946,N_646,N_2747);
nor U3947 (N_3947,N_2800,N_268);
nor U3948 (N_3948,N_1995,N_1538);
and U3949 (N_3949,N_18,N_1383);
and U3950 (N_3950,N_1015,N_1409);
or U3951 (N_3951,N_1518,N_1368);
xnor U3952 (N_3952,N_682,N_877);
and U3953 (N_3953,N_1595,N_2715);
nand U3954 (N_3954,N_2318,N_2859);
nand U3955 (N_3955,N_2888,N_571);
nand U3956 (N_3956,N_2001,N_1160);
or U3957 (N_3957,N_2364,N_2893);
nor U3958 (N_3958,N_1396,N_2196);
nand U3959 (N_3959,N_846,N_642);
nand U3960 (N_3960,N_2567,N_1948);
xnor U3961 (N_3961,N_505,N_634);
or U3962 (N_3962,N_727,N_2569);
or U3963 (N_3963,N_2388,N_2322);
and U3964 (N_3964,N_2484,N_2263);
nand U3965 (N_3965,N_450,N_2848);
and U3966 (N_3966,N_2510,N_1886);
or U3967 (N_3967,N_2881,N_1697);
and U3968 (N_3968,N_1342,N_2315);
or U3969 (N_3969,N_2876,N_197);
xor U3970 (N_3970,N_17,N_1812);
or U3971 (N_3971,N_914,N_1632);
nor U3972 (N_3972,N_2631,N_1753);
xor U3973 (N_3973,N_123,N_2588);
nand U3974 (N_3974,N_2370,N_412);
or U3975 (N_3975,N_1200,N_1930);
nand U3976 (N_3976,N_1254,N_362);
or U3977 (N_3977,N_1654,N_2414);
and U3978 (N_3978,N_1274,N_2215);
xor U3979 (N_3979,N_1612,N_2978);
nor U3980 (N_3980,N_2275,N_1140);
nand U3981 (N_3981,N_1890,N_2877);
or U3982 (N_3982,N_237,N_2220);
or U3983 (N_3983,N_569,N_1496);
nor U3984 (N_3984,N_2299,N_2999);
nand U3985 (N_3985,N_2086,N_282);
xor U3986 (N_3986,N_556,N_2899);
xor U3987 (N_3987,N_2995,N_1133);
nor U3988 (N_3988,N_831,N_2222);
nor U3989 (N_3989,N_1487,N_968);
nand U3990 (N_3990,N_315,N_2163);
xor U3991 (N_3991,N_2950,N_476);
xnor U3992 (N_3992,N_1203,N_1324);
and U3993 (N_3993,N_1152,N_2733);
nand U3994 (N_3994,N_1352,N_825);
nor U3995 (N_3995,N_718,N_488);
nand U3996 (N_3996,N_66,N_848);
nor U3997 (N_3997,N_2854,N_203);
nand U3998 (N_3998,N_2341,N_1722);
nor U3999 (N_3999,N_940,N_2261);
and U4000 (N_4000,N_1123,N_142);
and U4001 (N_4001,N_2055,N_2664);
nand U4002 (N_4002,N_2509,N_392);
or U4003 (N_4003,N_2686,N_660);
nor U4004 (N_4004,N_1145,N_341);
nand U4005 (N_4005,N_2702,N_2604);
and U4006 (N_4006,N_847,N_177);
xor U4007 (N_4007,N_1196,N_236);
or U4008 (N_4008,N_2234,N_1933);
nor U4009 (N_4009,N_2061,N_1108);
nor U4010 (N_4010,N_1778,N_1547);
nand U4011 (N_4011,N_1776,N_1606);
nand U4012 (N_4012,N_1204,N_1638);
nor U4013 (N_4013,N_2722,N_2519);
nand U4014 (N_4014,N_1574,N_605);
xnor U4015 (N_4015,N_1420,N_1042);
and U4016 (N_4016,N_1286,N_150);
xnor U4017 (N_4017,N_330,N_2940);
nor U4018 (N_4018,N_42,N_2989);
or U4019 (N_4019,N_2751,N_885);
nand U4020 (N_4020,N_209,N_2979);
nand U4021 (N_4021,N_2284,N_342);
nand U4022 (N_4022,N_1981,N_1666);
and U4023 (N_4023,N_1016,N_1648);
and U4024 (N_4024,N_515,N_314);
and U4025 (N_4025,N_1946,N_1709);
or U4026 (N_4026,N_2727,N_1640);
or U4027 (N_4027,N_912,N_1601);
xor U4028 (N_4028,N_1888,N_331);
and U4029 (N_4029,N_1711,N_1256);
or U4030 (N_4030,N_80,N_1389);
and U4031 (N_4031,N_2184,N_1910);
nor U4032 (N_4032,N_2750,N_1828);
nor U4033 (N_4033,N_2063,N_2470);
nor U4034 (N_4034,N_1461,N_413);
and U4035 (N_4035,N_1012,N_1683);
and U4036 (N_4036,N_707,N_1959);
or U4037 (N_4037,N_251,N_352);
or U4038 (N_4038,N_2570,N_939);
and U4039 (N_4039,N_428,N_333);
and U4040 (N_4040,N_1617,N_1327);
nand U4041 (N_4041,N_1579,N_921);
and U4042 (N_4042,N_781,N_1288);
nor U4043 (N_4043,N_702,N_33);
nand U4044 (N_4044,N_1056,N_104);
or U4045 (N_4045,N_1566,N_2219);
or U4046 (N_4046,N_410,N_2368);
xnor U4047 (N_4047,N_163,N_2238);
and U4048 (N_4048,N_1281,N_1576);
nor U4049 (N_4049,N_2467,N_755);
and U4050 (N_4050,N_2572,N_2864);
xor U4051 (N_4051,N_1700,N_2842);
nand U4052 (N_4052,N_1835,N_745);
or U4053 (N_4053,N_1325,N_230);
and U4054 (N_4054,N_1597,N_928);
nor U4055 (N_4055,N_1769,N_1190);
or U4056 (N_4056,N_1021,N_398);
or U4057 (N_4057,N_866,N_906);
xnor U4058 (N_4058,N_189,N_2729);
and U4059 (N_4059,N_2161,N_1631);
or U4060 (N_4060,N_1949,N_81);
nand U4061 (N_4061,N_522,N_1205);
or U4062 (N_4062,N_1734,N_2422);
nand U4063 (N_4063,N_1962,N_93);
or U4064 (N_4064,N_1111,N_1427);
nand U4065 (N_4065,N_175,N_639);
or U4066 (N_4066,N_633,N_1382);
nor U4067 (N_4067,N_375,N_2958);
nor U4068 (N_4068,N_95,N_1429);
nand U4069 (N_4069,N_2189,N_636);
nand U4070 (N_4070,N_2639,N_2658);
xor U4071 (N_4071,N_1905,N_2611);
or U4072 (N_4072,N_2652,N_2290);
nor U4073 (N_4073,N_531,N_2009);
or U4074 (N_4074,N_567,N_2739);
nor U4075 (N_4075,N_124,N_241);
nand U4076 (N_4076,N_929,N_1144);
nand U4077 (N_4077,N_2650,N_1656);
xnor U4078 (N_4078,N_853,N_1798);
xnor U4079 (N_4079,N_162,N_1614);
and U4080 (N_4080,N_2449,N_1156);
nor U4081 (N_4081,N_758,N_1073);
nor U4082 (N_4082,N_157,N_284);
nor U4083 (N_4083,N_689,N_357);
and U4084 (N_4084,N_1866,N_1955);
nand U4085 (N_4085,N_1173,N_2817);
nor U4086 (N_4086,N_1098,N_2953);
or U4087 (N_4087,N_2434,N_2171);
or U4088 (N_4088,N_300,N_608);
or U4089 (N_4089,N_2728,N_2649);
or U4090 (N_4090,N_1532,N_1052);
nor U4091 (N_4091,N_274,N_1604);
nor U4092 (N_4092,N_1343,N_158);
and U4093 (N_4093,N_2583,N_1540);
nor U4094 (N_4094,N_863,N_1582);
nand U4095 (N_4095,N_460,N_60);
or U4096 (N_4096,N_210,N_1956);
nand U4097 (N_4097,N_434,N_845);
nor U4098 (N_4098,N_2280,N_2420);
nor U4099 (N_4099,N_239,N_796);
nor U4100 (N_4100,N_1504,N_1603);
or U4101 (N_4101,N_2498,N_2997);
nor U4102 (N_4102,N_903,N_684);
nor U4103 (N_4103,N_2531,N_1087);
nor U4104 (N_4104,N_1701,N_1819);
or U4105 (N_4105,N_1364,N_200);
and U4106 (N_4106,N_1062,N_319);
and U4107 (N_4107,N_2632,N_714);
nor U4108 (N_4108,N_2035,N_752);
xor U4109 (N_4109,N_1285,N_1451);
or U4110 (N_4110,N_225,N_311);
or U4111 (N_4111,N_1283,N_2916);
nor U4112 (N_4112,N_2546,N_1553);
nand U4113 (N_4113,N_517,N_2921);
nor U4114 (N_4114,N_891,N_2786);
nand U4115 (N_4115,N_966,N_2068);
and U4116 (N_4116,N_1493,N_733);
xor U4117 (N_4117,N_750,N_1001);
or U4118 (N_4118,N_1628,N_2892);
and U4119 (N_4119,N_2758,N_2266);
nor U4120 (N_4120,N_2829,N_1889);
nand U4121 (N_4121,N_278,N_2690);
and U4122 (N_4122,N_2408,N_369);
or U4123 (N_4123,N_681,N_830);
and U4124 (N_4124,N_381,N_2554);
xnor U4125 (N_4125,N_2862,N_2552);
and U4126 (N_4126,N_234,N_868);
or U4127 (N_4127,N_2796,N_293);
nor U4128 (N_4128,N_1626,N_1102);
nand U4129 (N_4129,N_1831,N_2335);
or U4130 (N_4130,N_2937,N_2010);
or U4131 (N_4131,N_140,N_2707);
or U4132 (N_4132,N_2129,N_1780);
or U4133 (N_4133,N_560,N_2752);
xnor U4134 (N_4134,N_2435,N_451);
xnor U4135 (N_4135,N_1137,N_153);
and U4136 (N_4136,N_438,N_1350);
nand U4137 (N_4137,N_2159,N_2481);
xor U4138 (N_4138,N_1926,N_872);
and U4139 (N_4139,N_528,N_867);
and U4140 (N_4140,N_2982,N_483);
and U4141 (N_4141,N_425,N_1188);
nor U4142 (N_4142,N_620,N_1635);
nand U4143 (N_4143,N_2754,N_1489);
and U4144 (N_4144,N_111,N_58);
or U4145 (N_4145,N_963,N_566);
or U4146 (N_4146,N_2716,N_213);
and U4147 (N_4147,N_1212,N_1414);
or U4148 (N_4148,N_1410,N_1236);
xor U4149 (N_4149,N_1779,N_12);
and U4150 (N_4150,N_1070,N_951);
or U4151 (N_4151,N_1043,N_2665);
nor U4152 (N_4152,N_298,N_2457);
nor U4153 (N_4153,N_2480,N_1571);
xor U4154 (N_4154,N_2413,N_661);
or U4155 (N_4155,N_249,N_1674);
nand U4156 (N_4156,N_1040,N_1585);
or U4157 (N_4157,N_628,N_2923);
nand U4158 (N_4158,N_787,N_321);
xor U4159 (N_4159,N_527,N_1334);
nor U4160 (N_4160,N_543,N_1041);
and U4161 (N_4161,N_604,N_1075);
and U4162 (N_4162,N_205,N_621);
nand U4163 (N_4163,N_2331,N_1960);
or U4164 (N_4164,N_1002,N_1803);
nand U4165 (N_4165,N_2875,N_229);
and U4166 (N_4166,N_2195,N_1266);
nand U4167 (N_4167,N_1218,N_902);
or U4168 (N_4168,N_384,N_385);
and U4169 (N_4169,N_1243,N_1801);
nand U4170 (N_4170,N_2904,N_2306);
or U4171 (N_4171,N_358,N_1586);
nand U4172 (N_4172,N_2782,N_1112);
nor U4173 (N_4173,N_1887,N_1005);
nor U4174 (N_4174,N_1096,N_477);
nor U4175 (N_4175,N_2822,N_1675);
and U4176 (N_4176,N_1916,N_2092);
xnor U4177 (N_4177,N_1719,N_1911);
nor U4178 (N_4178,N_2054,N_1747);
and U4179 (N_4179,N_2771,N_1048);
or U4180 (N_4180,N_2149,N_860);
and U4181 (N_4181,N_2022,N_705);
nor U4182 (N_4182,N_2316,N_1251);
or U4183 (N_4183,N_2512,N_2866);
nor U4184 (N_4184,N_2369,N_2847);
nand U4185 (N_4185,N_2988,N_191);
or U4186 (N_4186,N_2120,N_2528);
and U4187 (N_4187,N_2558,N_546);
and U4188 (N_4188,N_1767,N_2320);
nor U4189 (N_4189,N_934,N_991);
or U4190 (N_4190,N_340,N_1336);
and U4191 (N_4191,N_1792,N_2744);
and U4192 (N_4192,N_2186,N_706);
nor U4193 (N_4193,N_383,N_1902);
and U4194 (N_4194,N_2885,N_763);
or U4195 (N_4195,N_1850,N_23);
nor U4196 (N_4196,N_617,N_2490);
nand U4197 (N_4197,N_472,N_313);
and U4198 (N_4198,N_2879,N_1366);
xor U4199 (N_4199,N_622,N_1846);
or U4200 (N_4200,N_783,N_131);
nand U4201 (N_4201,N_2692,N_942);
and U4202 (N_4202,N_743,N_193);
nand U4203 (N_4203,N_1467,N_220);
or U4204 (N_4204,N_2094,N_809);
or U4205 (N_4205,N_168,N_1993);
nor U4206 (N_4206,N_883,N_2734);
and U4207 (N_4207,N_1858,N_888);
xnor U4208 (N_4208,N_2501,N_1378);
nor U4209 (N_4209,N_1770,N_1559);
nand U4210 (N_4210,N_748,N_1565);
and U4211 (N_4211,N_2400,N_700);
and U4212 (N_4212,N_2837,N_2365);
nor U4213 (N_4213,N_2224,N_125);
or U4214 (N_4214,N_44,N_1807);
and U4215 (N_4215,N_1175,N_267);
or U4216 (N_4216,N_407,N_2411);
nand U4217 (N_4217,N_1799,N_1471);
or U4218 (N_4218,N_1920,N_323);
nor U4219 (N_4219,N_1241,N_2772);
nand U4220 (N_4220,N_2144,N_1242);
nand U4221 (N_4221,N_1536,N_553);
and U4222 (N_4222,N_160,N_1755);
or U4223 (N_4223,N_2380,N_836);
and U4224 (N_4224,N_2952,N_2415);
and U4225 (N_4225,N_905,N_1008);
and U4226 (N_4226,N_1672,N_2955);
and U4227 (N_4227,N_2917,N_2760);
nor U4228 (N_4228,N_722,N_437);
and U4229 (N_4229,N_1912,N_155);
nor U4230 (N_4230,N_1411,N_669);
or U4231 (N_4231,N_159,N_2352);
and U4232 (N_4232,N_2621,N_601);
and U4233 (N_4233,N_2139,N_1199);
or U4234 (N_4234,N_439,N_735);
and U4235 (N_4235,N_599,N_683);
xnor U4236 (N_4236,N_1814,N_2168);
nor U4237 (N_4237,N_482,N_530);
nand U4238 (N_4238,N_1998,N_1360);
and U4239 (N_4239,N_2644,N_259);
and U4240 (N_4240,N_1699,N_312);
and U4241 (N_4241,N_1469,N_2012);
and U4242 (N_4242,N_1618,N_1391);
or U4243 (N_4243,N_2399,N_2592);
nor U4244 (N_4244,N_238,N_822);
nand U4245 (N_4245,N_1611,N_2493);
or U4246 (N_4246,N_202,N_2391);
or U4247 (N_4247,N_1348,N_1884);
nor U4248 (N_4248,N_2233,N_254);
or U4249 (N_4249,N_2732,N_2628);
xor U4250 (N_4250,N_2886,N_2002);
and U4251 (N_4251,N_2208,N_1138);
or U4252 (N_4252,N_664,N_829);
nand U4253 (N_4253,N_1676,N_2142);
or U4254 (N_4254,N_2565,N_1028);
or U4255 (N_4255,N_1135,N_69);
or U4256 (N_4256,N_509,N_1076);
nor U4257 (N_4257,N_187,N_2147);
nor U4258 (N_4258,N_2008,N_1404);
nand U4259 (N_4259,N_1452,N_562);
nor U4260 (N_4260,N_1309,N_2424);
xnor U4261 (N_4261,N_499,N_31);
nor U4262 (N_4262,N_1583,N_2476);
and U4263 (N_4263,N_2688,N_692);
nor U4264 (N_4264,N_1558,N_279);
and U4265 (N_4265,N_329,N_1838);
or U4266 (N_4266,N_1972,N_363);
nand U4267 (N_4267,N_1444,N_2103);
or U4268 (N_4268,N_2871,N_1863);
nand U4269 (N_4269,N_536,N_317);
and U4270 (N_4270,N_2590,N_765);
and U4271 (N_4271,N_1262,N_1247);
nand U4272 (N_4272,N_2262,N_2544);
or U4273 (N_4273,N_2136,N_1229);
or U4274 (N_4274,N_2095,N_87);
nor U4275 (N_4275,N_1856,N_837);
xor U4276 (N_4276,N_354,N_1372);
nor U4277 (N_4277,N_2547,N_632);
or U4278 (N_4278,N_39,N_346);
and U4279 (N_4279,N_1605,N_1513);
and U4280 (N_4280,N_1903,N_2293);
nand U4281 (N_4281,N_1760,N_2534);
or U4282 (N_4282,N_2375,N_1289);
or U4283 (N_4283,N_420,N_2336);
or U4284 (N_4284,N_343,N_20);
or U4285 (N_4285,N_212,N_2843);
or U4286 (N_4286,N_1596,N_283);
nor U4287 (N_4287,N_2178,N_1997);
and U4288 (N_4288,N_678,N_2757);
nand U4289 (N_4289,N_1485,N_1502);
or U4290 (N_4290,N_1148,N_2761);
nor U4291 (N_4291,N_1115,N_1441);
and U4292 (N_4292,N_90,N_1690);
xor U4293 (N_4293,N_699,N_680);
nor U4294 (N_4294,N_1463,N_2396);
or U4295 (N_4295,N_800,N_1533);
nor U4296 (N_4296,N_174,N_724);
xor U4297 (N_4297,N_2153,N_1038);
nand U4298 (N_4298,N_2245,N_2797);
nor U4299 (N_4299,N_2169,N_1072);
and U4300 (N_4300,N_948,N_1745);
nand U4301 (N_4301,N_1732,N_2603);
nand U4302 (N_4302,N_2211,N_1430);
nand U4303 (N_4303,N_1258,N_1662);
nand U4304 (N_4304,N_1707,N_1641);
or U4305 (N_4305,N_576,N_1024);
and U4306 (N_4306,N_2477,N_1168);
or U4307 (N_4307,N_1252,N_96);
nand U4308 (N_4308,N_406,N_2584);
nor U4309 (N_4309,N_1754,N_805);
and U4310 (N_4310,N_99,N_295);
xor U4311 (N_4311,N_703,N_1432);
xnor U4312 (N_4312,N_1255,N_1824);
nor U4313 (N_4313,N_544,N_988);
or U4314 (N_4314,N_269,N_2453);
and U4315 (N_4315,N_600,N_1740);
nand U4316 (N_4316,N_54,N_1464);
or U4317 (N_4317,N_1616,N_2240);
nor U4318 (N_4318,N_1649,N_2497);
or U4319 (N_4319,N_2742,N_1158);
and U4320 (N_4320,N_516,N_192);
nor U4321 (N_4321,N_2150,N_950);
and U4322 (N_4322,N_1333,N_1026);
or U4323 (N_4323,N_52,N_2717);
or U4324 (N_4324,N_2858,N_6);
nor U4325 (N_4325,N_2043,N_2675);
nand U4326 (N_4326,N_1580,N_1438);
nand U4327 (N_4327,N_2783,N_1290);
nand U4328 (N_4328,N_1300,N_1483);
nand U4329 (N_4329,N_1562,N_1820);
nor U4330 (N_4330,N_273,N_2291);
nand U4331 (N_4331,N_1312,N_697);
nand U4332 (N_4332,N_2844,N_2491);
xnor U4333 (N_4333,N_1330,N_994);
and U4334 (N_4334,N_469,N_2308);
or U4335 (N_4335,N_1495,N_1985);
and U4336 (N_4336,N_1587,N_746);
nand U4337 (N_4337,N_433,N_1979);
and U4338 (N_4338,N_982,N_1003);
or U4339 (N_4339,N_679,N_2059);
nor U4340 (N_4340,N_1992,N_1677);
or U4341 (N_4341,N_34,N_2911);
or U4342 (N_4342,N_850,N_612);
or U4343 (N_4343,N_1118,N_2972);
nor U4344 (N_4344,N_1185,N_1402);
or U4345 (N_4345,N_2199,N_753);
and U4346 (N_4346,N_327,N_97);
xor U4347 (N_4347,N_2666,N_918);
nand U4348 (N_4348,N_2865,N_2216);
xor U4349 (N_4349,N_1511,N_2406);
nor U4350 (N_4350,N_2079,N_101);
or U4351 (N_4351,N_880,N_1405);
or U4352 (N_4352,N_2326,N_1074);
nand U4353 (N_4353,N_1064,N_2971);
nor U4354 (N_4354,N_1669,N_432);
nand U4355 (N_4355,N_2330,N_2517);
nor U4356 (N_4356,N_2462,N_2523);
and U4357 (N_4357,N_2626,N_739);
nand U4358 (N_4358,N_820,N_224);
nand U4359 (N_4359,N_1166,N_1355);
nand U4360 (N_4360,N_1299,N_464);
xnor U4361 (N_4361,N_595,N_1302);
and U4362 (N_4362,N_1150,N_2991);
or U4363 (N_4363,N_1139,N_1279);
and U4364 (N_4364,N_974,N_784);
nand U4365 (N_4365,N_924,N_1033);
nor U4366 (N_4366,N_1588,N_2973);
nand U4367 (N_4367,N_804,N_740);
or U4368 (N_4368,N_2170,N_1018);
nor U4369 (N_4369,N_2482,N_1079);
and U4370 (N_4370,N_2425,N_1534);
and U4371 (N_4371,N_1071,N_186);
or U4372 (N_4372,N_844,N_2469);
or U4373 (N_4373,N_759,N_307);
or U4374 (N_4374,N_618,N_2289);
and U4375 (N_4375,N_1868,N_2801);
nor U4376 (N_4376,N_512,N_2889);
nor U4377 (N_4377,N_1841,N_2056);
nand U4378 (N_4378,N_2,N_1726);
nand U4379 (N_4379,N_2052,N_2598);
or U4380 (N_4380,N_1852,N_1362);
nand U4381 (N_4381,N_711,N_1793);
and U4382 (N_4382,N_322,N_2221);
nand U4383 (N_4383,N_2748,N_1232);
xnor U4384 (N_4384,N_2332,N_1783);
xor U4385 (N_4385,N_1499,N_1328);
nor U4386 (N_4386,N_2674,N_258);
or U4387 (N_4387,N_1069,N_214);
or U4388 (N_4388,N_2520,N_418);
nand U4389 (N_4389,N_946,N_1351);
nand U4390 (N_4390,N_449,N_1035);
nor U4391 (N_4391,N_2154,N_2118);
or U4392 (N_4392,N_1870,N_2083);
and U4393 (N_4393,N_2676,N_2713);
nand U4394 (N_4394,N_2789,N_2574);
and U4395 (N_4395,N_2765,N_2557);
nor U4396 (N_4396,N_882,N_2774);
nor U4397 (N_4397,N_1928,N_1189);
nand U4398 (N_4398,N_892,N_960);
or U4399 (N_4399,N_1433,N_2970);
and U4400 (N_4400,N_2446,N_444);
and U4401 (N_4401,N_2113,N_1833);
or U4402 (N_4402,N_2464,N_2328);
and U4403 (N_4403,N_2595,N_1393);
nor U4404 (N_4404,N_2164,N_2935);
and U4405 (N_4405,N_593,N_1147);
nand U4406 (N_4406,N_1650,N_1716);
or U4407 (N_4407,N_2286,N_2281);
nor U4408 (N_4408,N_1527,N_2814);
xnor U4409 (N_4409,N_641,N_1723);
or U4410 (N_4410,N_812,N_2502);
nor U4411 (N_4411,N_1936,N_1454);
and U4412 (N_4412,N_487,N_344);
nand U4413 (N_4413,N_306,N_222);
or U4414 (N_4414,N_2015,N_2041);
nor U4415 (N_4415,N_1413,N_1724);
xnor U4416 (N_4416,N_775,N_2906);
nor U4417 (N_4417,N_2756,N_2745);
and U4418 (N_4418,N_657,N_778);
or U4419 (N_4419,N_503,N_2066);
and U4420 (N_4420,N_1276,N_1423);
and U4421 (N_4421,N_2577,N_2016);
or U4422 (N_4422,N_188,N_1872);
nand U4423 (N_4423,N_1000,N_802);
and U4424 (N_4424,N_774,N_2816);
nor U4425 (N_4425,N_996,N_1476);
xnor U4426 (N_4426,N_120,N_1155);
xor U4427 (N_4427,N_397,N_453);
nor U4428 (N_4428,N_969,N_838);
and U4429 (N_4429,N_1316,N_2678);
xor U4430 (N_4430,N_818,N_2297);
nand U4431 (N_4431,N_217,N_1921);
nand U4432 (N_4432,N_2694,N_2123);
nand U4433 (N_4433,N_431,N_2214);
nor U4434 (N_4434,N_2428,N_82);
or U4435 (N_4435,N_2456,N_1308);
or U4436 (N_4436,N_1149,N_685);
and U4437 (N_4437,N_1036,N_1590);
and U4438 (N_4438,N_2996,N_1306);
nand U4439 (N_4439,N_2376,N_1600);
xnor U4440 (N_4440,N_2919,N_930);
nand U4441 (N_4441,N_2740,N_133);
nor U4442 (N_4442,N_46,N_1901);
and U4443 (N_4443,N_2964,N_529);
or U4444 (N_4444,N_539,N_2735);
nand U4445 (N_4445,N_226,N_629);
nor U4446 (N_4446,N_1937,N_149);
nor U4447 (N_4447,N_687,N_260);
and U4448 (N_4448,N_2361,N_2962);
nand U4449 (N_4449,N_78,N_1802);
and U4450 (N_4450,N_1568,N_795);
nor U4451 (N_4451,N_1885,N_1899);
nor U4452 (N_4452,N_2615,N_769);
or U4453 (N_4453,N_32,N_972);
or U4454 (N_4454,N_1084,N_122);
and U4455 (N_4455,N_2160,N_959);
xor U4456 (N_4456,N_2489,N_1230);
or U4457 (N_4457,N_2831,N_1757);
nand U4458 (N_4458,N_1332,N_2363);
and U4459 (N_4459,N_1567,N_1938);
nand U4460 (N_4460,N_1988,N_1693);
and U4461 (N_4461,N_2832,N_856);
nor U4462 (N_4462,N_2175,N_2977);
nor U4463 (N_4463,N_814,N_2755);
nand U4464 (N_4464,N_1752,N_932);
or U4465 (N_4465,N_582,N_1968);
nor U4466 (N_4466,N_843,N_1966);
and U4467 (N_4467,N_2533,N_486);
xnor U4468 (N_4468,N_1291,N_2288);
nor U4469 (N_4469,N_1986,N_1379);
nand U4470 (N_4470,N_1060,N_821);
or U4471 (N_4471,N_2242,N_1257);
and U4472 (N_4472,N_609,N_2057);
nand U4473 (N_4473,N_1765,N_864);
and U4474 (N_4474,N_917,N_2270);
or U4475 (N_4475,N_1751,N_1853);
nand U4476 (N_4476,N_619,N_1480);
or U4477 (N_4477,N_1206,N_2947);
xor U4478 (N_4478,N_11,N_1387);
nor U4479 (N_4479,N_2478,N_2629);
or U4480 (N_4480,N_2402,N_935);
nand U4481 (N_4481,N_1207,N_1703);
and U4482 (N_4482,N_1836,N_2321);
or U4483 (N_4483,N_1849,N_71);
nand U4484 (N_4484,N_1125,N_676);
nand U4485 (N_4485,N_366,N_2327);
nand U4486 (N_4486,N_1691,N_2007);
nor U4487 (N_4487,N_161,N_1375);
nor U4488 (N_4488,N_1371,N_828);
nor U4489 (N_4489,N_1686,N_501);
xnor U4490 (N_4490,N_2337,N_495);
nand U4491 (N_4491,N_1244,N_1373);
and U4492 (N_4492,N_2267,N_2193);
or U4493 (N_4493,N_1871,N_1659);
and U4494 (N_4494,N_615,N_2157);
nand U4495 (N_4495,N_2589,N_1878);
nor U4496 (N_4496,N_359,N_1234);
xor U4497 (N_4497,N_952,N_455);
and U4498 (N_4498,N_468,N_555);
nor U4499 (N_4499,N_1136,N_1900);
and U4500 (N_4500,N_816,N_1310);
nor U4501 (N_4501,N_1247,N_2157);
nor U4502 (N_4502,N_1676,N_204);
nand U4503 (N_4503,N_2913,N_374);
and U4504 (N_4504,N_1216,N_557);
nand U4505 (N_4505,N_2445,N_369);
nor U4506 (N_4506,N_2259,N_192);
xnor U4507 (N_4507,N_1809,N_2324);
nor U4508 (N_4508,N_1662,N_903);
nand U4509 (N_4509,N_1445,N_630);
nor U4510 (N_4510,N_1481,N_879);
and U4511 (N_4511,N_2489,N_611);
nor U4512 (N_4512,N_91,N_605);
nand U4513 (N_4513,N_457,N_172);
or U4514 (N_4514,N_9,N_1957);
or U4515 (N_4515,N_749,N_1547);
or U4516 (N_4516,N_1339,N_220);
or U4517 (N_4517,N_2684,N_170);
and U4518 (N_4518,N_1061,N_1590);
or U4519 (N_4519,N_2726,N_2111);
nand U4520 (N_4520,N_1591,N_1443);
nor U4521 (N_4521,N_164,N_2005);
nand U4522 (N_4522,N_2498,N_1737);
or U4523 (N_4523,N_153,N_2085);
xnor U4524 (N_4524,N_37,N_1531);
nor U4525 (N_4525,N_2810,N_1658);
or U4526 (N_4526,N_1120,N_1854);
or U4527 (N_4527,N_433,N_1326);
nand U4528 (N_4528,N_2884,N_34);
nor U4529 (N_4529,N_1428,N_1185);
nor U4530 (N_4530,N_2337,N_1151);
and U4531 (N_4531,N_1506,N_146);
nand U4532 (N_4532,N_2999,N_276);
nand U4533 (N_4533,N_1353,N_2578);
nor U4534 (N_4534,N_1511,N_281);
or U4535 (N_4535,N_42,N_1323);
or U4536 (N_4536,N_1107,N_1260);
nor U4537 (N_4537,N_2908,N_691);
nand U4538 (N_4538,N_65,N_406);
or U4539 (N_4539,N_1603,N_44);
nor U4540 (N_4540,N_2072,N_2887);
and U4541 (N_4541,N_1805,N_1622);
nor U4542 (N_4542,N_2670,N_2125);
nand U4543 (N_4543,N_1629,N_2491);
xnor U4544 (N_4544,N_632,N_2624);
nand U4545 (N_4545,N_1777,N_1264);
nor U4546 (N_4546,N_2890,N_1850);
nor U4547 (N_4547,N_851,N_635);
xor U4548 (N_4548,N_2886,N_973);
and U4549 (N_4549,N_1673,N_1183);
or U4550 (N_4550,N_1603,N_447);
or U4551 (N_4551,N_50,N_1206);
nand U4552 (N_4552,N_1590,N_1407);
or U4553 (N_4553,N_2974,N_1345);
or U4554 (N_4554,N_2037,N_2416);
nor U4555 (N_4555,N_2222,N_215);
or U4556 (N_4556,N_552,N_2484);
nand U4557 (N_4557,N_1431,N_2351);
and U4558 (N_4558,N_729,N_94);
nand U4559 (N_4559,N_2434,N_827);
or U4560 (N_4560,N_765,N_1874);
nand U4561 (N_4561,N_1053,N_1830);
or U4562 (N_4562,N_235,N_2345);
and U4563 (N_4563,N_2837,N_1998);
nand U4564 (N_4564,N_2398,N_840);
nand U4565 (N_4565,N_950,N_1059);
and U4566 (N_4566,N_926,N_2393);
or U4567 (N_4567,N_1002,N_101);
or U4568 (N_4568,N_1359,N_1955);
and U4569 (N_4569,N_356,N_2191);
nor U4570 (N_4570,N_2063,N_125);
nor U4571 (N_4571,N_1515,N_977);
nand U4572 (N_4572,N_1630,N_297);
nand U4573 (N_4573,N_227,N_1122);
nor U4574 (N_4574,N_2172,N_2848);
xnor U4575 (N_4575,N_1769,N_134);
or U4576 (N_4576,N_1328,N_1145);
xor U4577 (N_4577,N_1442,N_938);
and U4578 (N_4578,N_2835,N_57);
nand U4579 (N_4579,N_436,N_950);
nor U4580 (N_4580,N_2834,N_1337);
and U4581 (N_4581,N_1533,N_2076);
or U4582 (N_4582,N_2478,N_1661);
or U4583 (N_4583,N_578,N_1366);
and U4584 (N_4584,N_2052,N_1194);
nor U4585 (N_4585,N_1181,N_2755);
or U4586 (N_4586,N_2343,N_489);
or U4587 (N_4587,N_1886,N_2894);
or U4588 (N_4588,N_561,N_2424);
xnor U4589 (N_4589,N_2098,N_2094);
or U4590 (N_4590,N_1195,N_1520);
or U4591 (N_4591,N_1016,N_957);
xor U4592 (N_4592,N_341,N_1258);
nor U4593 (N_4593,N_1795,N_2038);
xnor U4594 (N_4594,N_2411,N_2237);
nor U4595 (N_4595,N_2545,N_1297);
and U4596 (N_4596,N_2283,N_2381);
nand U4597 (N_4597,N_1462,N_1541);
or U4598 (N_4598,N_584,N_2075);
or U4599 (N_4599,N_825,N_917);
nand U4600 (N_4600,N_2064,N_556);
nor U4601 (N_4601,N_543,N_2203);
or U4602 (N_4602,N_513,N_2023);
or U4603 (N_4603,N_1508,N_2458);
or U4604 (N_4604,N_2457,N_2298);
nand U4605 (N_4605,N_2044,N_2645);
or U4606 (N_4606,N_1667,N_1799);
or U4607 (N_4607,N_2366,N_623);
and U4608 (N_4608,N_612,N_2794);
xnor U4609 (N_4609,N_618,N_1595);
and U4610 (N_4610,N_1854,N_2134);
nor U4611 (N_4611,N_982,N_1113);
nand U4612 (N_4612,N_787,N_2526);
nor U4613 (N_4613,N_1342,N_1942);
xor U4614 (N_4614,N_2050,N_308);
and U4615 (N_4615,N_141,N_2304);
nand U4616 (N_4616,N_1061,N_1546);
nor U4617 (N_4617,N_2002,N_1981);
nand U4618 (N_4618,N_2897,N_1960);
xnor U4619 (N_4619,N_2216,N_1636);
or U4620 (N_4620,N_2425,N_252);
nor U4621 (N_4621,N_2781,N_816);
nor U4622 (N_4622,N_2472,N_1580);
nor U4623 (N_4623,N_1887,N_1216);
or U4624 (N_4624,N_56,N_2591);
nor U4625 (N_4625,N_1390,N_646);
nand U4626 (N_4626,N_556,N_316);
and U4627 (N_4627,N_1528,N_1679);
or U4628 (N_4628,N_756,N_290);
nand U4629 (N_4629,N_2418,N_1523);
or U4630 (N_4630,N_1677,N_480);
or U4631 (N_4631,N_334,N_1778);
or U4632 (N_4632,N_1191,N_1639);
xnor U4633 (N_4633,N_1771,N_1330);
or U4634 (N_4634,N_2385,N_653);
nor U4635 (N_4635,N_839,N_1828);
or U4636 (N_4636,N_2982,N_615);
or U4637 (N_4637,N_2314,N_303);
or U4638 (N_4638,N_2673,N_381);
or U4639 (N_4639,N_276,N_2465);
nor U4640 (N_4640,N_2973,N_611);
nor U4641 (N_4641,N_972,N_68);
and U4642 (N_4642,N_2049,N_2151);
nor U4643 (N_4643,N_2066,N_1919);
nand U4644 (N_4644,N_899,N_2618);
and U4645 (N_4645,N_1851,N_1288);
nor U4646 (N_4646,N_2209,N_1925);
nand U4647 (N_4647,N_1694,N_2181);
xor U4648 (N_4648,N_2719,N_1992);
nor U4649 (N_4649,N_2652,N_2759);
nor U4650 (N_4650,N_1431,N_2114);
and U4651 (N_4651,N_1264,N_558);
nand U4652 (N_4652,N_1259,N_1840);
nand U4653 (N_4653,N_234,N_1971);
nor U4654 (N_4654,N_2564,N_2191);
and U4655 (N_4655,N_2490,N_449);
and U4656 (N_4656,N_2969,N_159);
and U4657 (N_4657,N_1164,N_937);
nor U4658 (N_4658,N_1535,N_1848);
or U4659 (N_4659,N_758,N_1196);
nor U4660 (N_4660,N_1809,N_1655);
or U4661 (N_4661,N_264,N_2173);
nand U4662 (N_4662,N_2021,N_1873);
or U4663 (N_4663,N_68,N_1063);
or U4664 (N_4664,N_2504,N_1218);
or U4665 (N_4665,N_1740,N_2526);
and U4666 (N_4666,N_453,N_1710);
or U4667 (N_4667,N_1439,N_2402);
or U4668 (N_4668,N_168,N_916);
nand U4669 (N_4669,N_1628,N_455);
and U4670 (N_4670,N_1436,N_1264);
xor U4671 (N_4671,N_1863,N_2880);
or U4672 (N_4672,N_1262,N_1623);
and U4673 (N_4673,N_1539,N_2590);
and U4674 (N_4674,N_2799,N_150);
nand U4675 (N_4675,N_2747,N_1535);
or U4676 (N_4676,N_387,N_2695);
and U4677 (N_4677,N_2556,N_1266);
or U4678 (N_4678,N_127,N_59);
or U4679 (N_4679,N_2873,N_48);
and U4680 (N_4680,N_1240,N_2171);
or U4681 (N_4681,N_2406,N_1692);
nand U4682 (N_4682,N_584,N_2168);
nor U4683 (N_4683,N_2225,N_2799);
nor U4684 (N_4684,N_1656,N_2347);
or U4685 (N_4685,N_2860,N_796);
or U4686 (N_4686,N_2860,N_2684);
nor U4687 (N_4687,N_1309,N_1487);
or U4688 (N_4688,N_227,N_1116);
nor U4689 (N_4689,N_1560,N_2329);
or U4690 (N_4690,N_2496,N_2452);
and U4691 (N_4691,N_1003,N_2796);
nand U4692 (N_4692,N_2051,N_525);
nand U4693 (N_4693,N_2874,N_1150);
nand U4694 (N_4694,N_355,N_1843);
nor U4695 (N_4695,N_2194,N_2184);
nand U4696 (N_4696,N_189,N_1899);
nand U4697 (N_4697,N_210,N_650);
or U4698 (N_4698,N_2520,N_2995);
and U4699 (N_4699,N_2280,N_1086);
nand U4700 (N_4700,N_2484,N_3);
or U4701 (N_4701,N_2440,N_2771);
and U4702 (N_4702,N_717,N_909);
and U4703 (N_4703,N_1780,N_2411);
and U4704 (N_4704,N_333,N_2053);
and U4705 (N_4705,N_2266,N_1928);
and U4706 (N_4706,N_674,N_2902);
and U4707 (N_4707,N_2147,N_2227);
and U4708 (N_4708,N_589,N_1177);
nor U4709 (N_4709,N_928,N_490);
and U4710 (N_4710,N_747,N_461);
nor U4711 (N_4711,N_1282,N_2860);
nand U4712 (N_4712,N_2063,N_1809);
or U4713 (N_4713,N_1457,N_260);
nor U4714 (N_4714,N_2450,N_20);
nand U4715 (N_4715,N_2673,N_1358);
nand U4716 (N_4716,N_202,N_1040);
nand U4717 (N_4717,N_1678,N_1136);
nand U4718 (N_4718,N_28,N_351);
nor U4719 (N_4719,N_1888,N_1365);
nand U4720 (N_4720,N_1621,N_88);
nand U4721 (N_4721,N_363,N_2233);
or U4722 (N_4722,N_1928,N_2017);
and U4723 (N_4723,N_1281,N_1802);
and U4724 (N_4724,N_65,N_1610);
or U4725 (N_4725,N_2450,N_772);
or U4726 (N_4726,N_2097,N_1190);
nand U4727 (N_4727,N_1753,N_151);
nor U4728 (N_4728,N_2186,N_1561);
nand U4729 (N_4729,N_320,N_1732);
and U4730 (N_4730,N_2849,N_2552);
xor U4731 (N_4731,N_1865,N_1107);
and U4732 (N_4732,N_2444,N_1499);
nor U4733 (N_4733,N_2812,N_2699);
or U4734 (N_4734,N_1742,N_27);
nor U4735 (N_4735,N_233,N_1695);
and U4736 (N_4736,N_2254,N_1236);
nand U4737 (N_4737,N_2683,N_2127);
nor U4738 (N_4738,N_2414,N_1022);
and U4739 (N_4739,N_1036,N_371);
nand U4740 (N_4740,N_1077,N_765);
xor U4741 (N_4741,N_1197,N_2702);
xor U4742 (N_4742,N_2410,N_203);
nor U4743 (N_4743,N_885,N_261);
nand U4744 (N_4744,N_483,N_2753);
xnor U4745 (N_4745,N_1578,N_1614);
or U4746 (N_4746,N_577,N_779);
nand U4747 (N_4747,N_1406,N_1068);
nand U4748 (N_4748,N_1615,N_2158);
nor U4749 (N_4749,N_1581,N_1464);
nand U4750 (N_4750,N_1603,N_1629);
nor U4751 (N_4751,N_476,N_2273);
nand U4752 (N_4752,N_2215,N_929);
nor U4753 (N_4753,N_2041,N_2867);
xnor U4754 (N_4754,N_1999,N_1882);
or U4755 (N_4755,N_723,N_1807);
or U4756 (N_4756,N_2509,N_1324);
and U4757 (N_4757,N_2972,N_1004);
and U4758 (N_4758,N_694,N_280);
nor U4759 (N_4759,N_1605,N_1113);
nor U4760 (N_4760,N_2953,N_2343);
or U4761 (N_4761,N_504,N_1256);
and U4762 (N_4762,N_843,N_955);
or U4763 (N_4763,N_763,N_1906);
or U4764 (N_4764,N_2820,N_2801);
or U4765 (N_4765,N_2003,N_546);
or U4766 (N_4766,N_1402,N_1817);
nor U4767 (N_4767,N_883,N_711);
or U4768 (N_4768,N_1831,N_1141);
nor U4769 (N_4769,N_2913,N_773);
nand U4770 (N_4770,N_114,N_2165);
nor U4771 (N_4771,N_150,N_1679);
nor U4772 (N_4772,N_1910,N_2632);
nand U4773 (N_4773,N_772,N_581);
nand U4774 (N_4774,N_324,N_455);
and U4775 (N_4775,N_852,N_2969);
nand U4776 (N_4776,N_516,N_315);
nor U4777 (N_4777,N_530,N_1983);
nand U4778 (N_4778,N_776,N_856);
or U4779 (N_4779,N_999,N_1300);
or U4780 (N_4780,N_581,N_309);
and U4781 (N_4781,N_100,N_1931);
nand U4782 (N_4782,N_2014,N_1628);
or U4783 (N_4783,N_1273,N_742);
nand U4784 (N_4784,N_767,N_594);
or U4785 (N_4785,N_2847,N_798);
nand U4786 (N_4786,N_2769,N_1409);
nor U4787 (N_4787,N_812,N_1937);
nand U4788 (N_4788,N_561,N_1261);
nand U4789 (N_4789,N_967,N_954);
xnor U4790 (N_4790,N_2568,N_1499);
and U4791 (N_4791,N_606,N_354);
or U4792 (N_4792,N_2168,N_1245);
or U4793 (N_4793,N_1888,N_2650);
nor U4794 (N_4794,N_1143,N_1450);
and U4795 (N_4795,N_2161,N_1639);
nand U4796 (N_4796,N_2848,N_589);
nor U4797 (N_4797,N_385,N_132);
nand U4798 (N_4798,N_1633,N_1046);
or U4799 (N_4799,N_2717,N_1229);
nand U4800 (N_4800,N_1907,N_1554);
nand U4801 (N_4801,N_576,N_2445);
nor U4802 (N_4802,N_1250,N_2320);
nor U4803 (N_4803,N_66,N_2302);
or U4804 (N_4804,N_2751,N_691);
nor U4805 (N_4805,N_657,N_1765);
nand U4806 (N_4806,N_981,N_1942);
and U4807 (N_4807,N_688,N_929);
nand U4808 (N_4808,N_1822,N_860);
and U4809 (N_4809,N_918,N_2341);
or U4810 (N_4810,N_2305,N_541);
nor U4811 (N_4811,N_2200,N_315);
and U4812 (N_4812,N_1469,N_1382);
nor U4813 (N_4813,N_27,N_396);
nor U4814 (N_4814,N_1593,N_2626);
or U4815 (N_4815,N_2865,N_821);
or U4816 (N_4816,N_737,N_862);
nor U4817 (N_4817,N_1693,N_2641);
nor U4818 (N_4818,N_71,N_625);
and U4819 (N_4819,N_1256,N_453);
and U4820 (N_4820,N_1883,N_423);
nand U4821 (N_4821,N_985,N_759);
nor U4822 (N_4822,N_2307,N_569);
nor U4823 (N_4823,N_734,N_818);
or U4824 (N_4824,N_2842,N_2695);
or U4825 (N_4825,N_829,N_2850);
and U4826 (N_4826,N_2058,N_2963);
or U4827 (N_4827,N_1973,N_1968);
xnor U4828 (N_4828,N_303,N_1148);
nor U4829 (N_4829,N_1637,N_1281);
nor U4830 (N_4830,N_705,N_905);
or U4831 (N_4831,N_1243,N_2830);
nand U4832 (N_4832,N_281,N_714);
nor U4833 (N_4833,N_705,N_2136);
or U4834 (N_4834,N_1323,N_1786);
nand U4835 (N_4835,N_2895,N_1311);
xnor U4836 (N_4836,N_335,N_1320);
and U4837 (N_4837,N_138,N_1165);
nand U4838 (N_4838,N_2516,N_1468);
or U4839 (N_4839,N_1819,N_2391);
nand U4840 (N_4840,N_2689,N_2515);
nor U4841 (N_4841,N_156,N_2199);
nor U4842 (N_4842,N_2940,N_567);
or U4843 (N_4843,N_179,N_266);
xor U4844 (N_4844,N_1015,N_387);
and U4845 (N_4845,N_2510,N_595);
nand U4846 (N_4846,N_2585,N_2841);
nand U4847 (N_4847,N_2507,N_1168);
nor U4848 (N_4848,N_1126,N_237);
and U4849 (N_4849,N_866,N_1181);
or U4850 (N_4850,N_1440,N_388);
nor U4851 (N_4851,N_231,N_521);
xor U4852 (N_4852,N_83,N_1384);
and U4853 (N_4853,N_1180,N_2179);
and U4854 (N_4854,N_1986,N_1517);
or U4855 (N_4855,N_2704,N_1364);
or U4856 (N_4856,N_1573,N_1464);
nor U4857 (N_4857,N_1852,N_442);
nor U4858 (N_4858,N_1680,N_1037);
nor U4859 (N_4859,N_1354,N_2990);
and U4860 (N_4860,N_2742,N_2686);
nor U4861 (N_4861,N_1982,N_550);
xor U4862 (N_4862,N_2249,N_1702);
nor U4863 (N_4863,N_1658,N_538);
or U4864 (N_4864,N_766,N_2794);
or U4865 (N_4865,N_2491,N_2570);
nor U4866 (N_4866,N_21,N_1574);
or U4867 (N_4867,N_10,N_2127);
or U4868 (N_4868,N_973,N_1329);
nand U4869 (N_4869,N_2525,N_1033);
or U4870 (N_4870,N_1843,N_1717);
nand U4871 (N_4871,N_2314,N_2889);
nor U4872 (N_4872,N_2266,N_870);
nor U4873 (N_4873,N_2755,N_1365);
nand U4874 (N_4874,N_1083,N_1493);
nand U4875 (N_4875,N_1924,N_2455);
nor U4876 (N_4876,N_1610,N_1591);
and U4877 (N_4877,N_370,N_961);
nand U4878 (N_4878,N_194,N_2205);
and U4879 (N_4879,N_2725,N_873);
and U4880 (N_4880,N_820,N_2837);
or U4881 (N_4881,N_2519,N_1408);
nor U4882 (N_4882,N_1305,N_1801);
and U4883 (N_4883,N_905,N_1585);
or U4884 (N_4884,N_2658,N_1930);
nor U4885 (N_4885,N_753,N_834);
and U4886 (N_4886,N_2978,N_1301);
nand U4887 (N_4887,N_2380,N_2359);
xnor U4888 (N_4888,N_2066,N_729);
nand U4889 (N_4889,N_523,N_476);
nand U4890 (N_4890,N_2813,N_865);
nand U4891 (N_4891,N_2049,N_2814);
nand U4892 (N_4892,N_2866,N_2730);
nor U4893 (N_4893,N_2028,N_2412);
and U4894 (N_4894,N_2184,N_1214);
and U4895 (N_4895,N_2604,N_2550);
xor U4896 (N_4896,N_593,N_760);
xnor U4897 (N_4897,N_1462,N_1549);
or U4898 (N_4898,N_1680,N_2851);
nand U4899 (N_4899,N_687,N_1751);
nor U4900 (N_4900,N_797,N_1725);
and U4901 (N_4901,N_1697,N_1815);
nand U4902 (N_4902,N_1453,N_2842);
nor U4903 (N_4903,N_2302,N_1146);
and U4904 (N_4904,N_917,N_1475);
and U4905 (N_4905,N_375,N_2927);
or U4906 (N_4906,N_832,N_1173);
nor U4907 (N_4907,N_1755,N_2742);
nor U4908 (N_4908,N_2273,N_1710);
nand U4909 (N_4909,N_1756,N_261);
xor U4910 (N_4910,N_1787,N_1743);
nor U4911 (N_4911,N_2403,N_116);
or U4912 (N_4912,N_2634,N_69);
xor U4913 (N_4913,N_1220,N_719);
xor U4914 (N_4914,N_2329,N_2548);
and U4915 (N_4915,N_2001,N_2618);
or U4916 (N_4916,N_1340,N_2602);
nor U4917 (N_4917,N_1575,N_1263);
nand U4918 (N_4918,N_103,N_141);
nand U4919 (N_4919,N_2729,N_1139);
nand U4920 (N_4920,N_1804,N_1043);
nand U4921 (N_4921,N_878,N_1632);
nand U4922 (N_4922,N_2226,N_965);
xnor U4923 (N_4923,N_1832,N_2874);
or U4924 (N_4924,N_1396,N_2847);
nor U4925 (N_4925,N_729,N_1805);
nor U4926 (N_4926,N_713,N_1457);
nand U4927 (N_4927,N_2160,N_2348);
nor U4928 (N_4928,N_1299,N_2539);
nor U4929 (N_4929,N_586,N_2186);
xnor U4930 (N_4930,N_1666,N_1889);
and U4931 (N_4931,N_2784,N_161);
nor U4932 (N_4932,N_2681,N_2898);
or U4933 (N_4933,N_520,N_1886);
nand U4934 (N_4934,N_1088,N_888);
and U4935 (N_4935,N_2396,N_740);
nand U4936 (N_4936,N_1809,N_1065);
nor U4937 (N_4937,N_1359,N_694);
nand U4938 (N_4938,N_291,N_1069);
and U4939 (N_4939,N_206,N_1770);
and U4940 (N_4940,N_1004,N_1239);
or U4941 (N_4941,N_2516,N_2184);
nand U4942 (N_4942,N_708,N_2528);
and U4943 (N_4943,N_1002,N_1224);
and U4944 (N_4944,N_1243,N_189);
nand U4945 (N_4945,N_1810,N_392);
and U4946 (N_4946,N_2068,N_922);
xnor U4947 (N_4947,N_1027,N_2494);
xor U4948 (N_4948,N_1537,N_2531);
and U4949 (N_4949,N_1565,N_368);
xnor U4950 (N_4950,N_1398,N_135);
nand U4951 (N_4951,N_772,N_2800);
nor U4952 (N_4952,N_1592,N_2348);
nor U4953 (N_4953,N_2579,N_1846);
nand U4954 (N_4954,N_2500,N_307);
xnor U4955 (N_4955,N_610,N_2585);
and U4956 (N_4956,N_447,N_661);
or U4957 (N_4957,N_2820,N_2214);
and U4958 (N_4958,N_1266,N_1903);
and U4959 (N_4959,N_650,N_2231);
or U4960 (N_4960,N_2454,N_2125);
and U4961 (N_4961,N_2391,N_982);
nor U4962 (N_4962,N_400,N_367);
or U4963 (N_4963,N_1758,N_2861);
and U4964 (N_4964,N_2028,N_1066);
or U4965 (N_4965,N_2248,N_1407);
nor U4966 (N_4966,N_170,N_268);
xnor U4967 (N_4967,N_1661,N_805);
and U4968 (N_4968,N_254,N_776);
nor U4969 (N_4969,N_2601,N_1172);
or U4970 (N_4970,N_1919,N_1050);
nor U4971 (N_4971,N_905,N_2202);
nand U4972 (N_4972,N_1868,N_1257);
and U4973 (N_4973,N_171,N_256);
or U4974 (N_4974,N_2932,N_1360);
or U4975 (N_4975,N_2905,N_248);
and U4976 (N_4976,N_1568,N_2855);
xnor U4977 (N_4977,N_75,N_169);
nor U4978 (N_4978,N_1619,N_1343);
nor U4979 (N_4979,N_1402,N_1974);
xnor U4980 (N_4980,N_2215,N_2720);
or U4981 (N_4981,N_694,N_2209);
or U4982 (N_4982,N_1336,N_718);
nand U4983 (N_4983,N_2997,N_2946);
or U4984 (N_4984,N_1082,N_1523);
nor U4985 (N_4985,N_1116,N_1396);
nand U4986 (N_4986,N_2353,N_2510);
nand U4987 (N_4987,N_894,N_2107);
nand U4988 (N_4988,N_996,N_919);
xnor U4989 (N_4989,N_763,N_51);
nand U4990 (N_4990,N_1767,N_1486);
and U4991 (N_4991,N_2958,N_2597);
nand U4992 (N_4992,N_59,N_892);
nor U4993 (N_4993,N_306,N_2401);
and U4994 (N_4994,N_1263,N_1830);
xnor U4995 (N_4995,N_780,N_2180);
nor U4996 (N_4996,N_1752,N_873);
xor U4997 (N_4997,N_7,N_2004);
nor U4998 (N_4998,N_1744,N_1152);
nor U4999 (N_4999,N_545,N_2571);
xor U5000 (N_5000,N_2502,N_1179);
nor U5001 (N_5001,N_1471,N_2405);
or U5002 (N_5002,N_2675,N_1931);
and U5003 (N_5003,N_2372,N_1241);
nor U5004 (N_5004,N_683,N_841);
and U5005 (N_5005,N_428,N_908);
xnor U5006 (N_5006,N_1008,N_2449);
nand U5007 (N_5007,N_2332,N_861);
or U5008 (N_5008,N_228,N_1330);
or U5009 (N_5009,N_1165,N_1613);
nand U5010 (N_5010,N_67,N_2261);
and U5011 (N_5011,N_413,N_696);
and U5012 (N_5012,N_782,N_2961);
or U5013 (N_5013,N_377,N_2236);
and U5014 (N_5014,N_961,N_1767);
nor U5015 (N_5015,N_495,N_2883);
nor U5016 (N_5016,N_1023,N_2693);
and U5017 (N_5017,N_715,N_342);
nor U5018 (N_5018,N_734,N_2392);
or U5019 (N_5019,N_2409,N_450);
or U5020 (N_5020,N_2545,N_1014);
or U5021 (N_5021,N_2118,N_1717);
and U5022 (N_5022,N_57,N_1442);
or U5023 (N_5023,N_884,N_2794);
nand U5024 (N_5024,N_664,N_776);
and U5025 (N_5025,N_960,N_1619);
or U5026 (N_5026,N_125,N_2965);
xor U5027 (N_5027,N_2728,N_156);
nand U5028 (N_5028,N_1921,N_2859);
nor U5029 (N_5029,N_10,N_1490);
or U5030 (N_5030,N_2396,N_1776);
nand U5031 (N_5031,N_2119,N_2941);
nand U5032 (N_5032,N_1024,N_58);
nand U5033 (N_5033,N_804,N_2625);
or U5034 (N_5034,N_1532,N_715);
nand U5035 (N_5035,N_537,N_1729);
nand U5036 (N_5036,N_2960,N_1696);
nand U5037 (N_5037,N_743,N_2483);
and U5038 (N_5038,N_799,N_641);
nor U5039 (N_5039,N_1460,N_774);
or U5040 (N_5040,N_2386,N_1736);
nand U5041 (N_5041,N_1128,N_1095);
nor U5042 (N_5042,N_2691,N_1326);
and U5043 (N_5043,N_1575,N_1774);
nor U5044 (N_5044,N_1359,N_110);
or U5045 (N_5045,N_2468,N_2466);
nor U5046 (N_5046,N_28,N_52);
and U5047 (N_5047,N_1501,N_2786);
or U5048 (N_5048,N_1288,N_1977);
nand U5049 (N_5049,N_428,N_12);
and U5050 (N_5050,N_1667,N_1991);
nor U5051 (N_5051,N_742,N_1849);
nor U5052 (N_5052,N_1774,N_297);
nor U5053 (N_5053,N_384,N_251);
xor U5054 (N_5054,N_70,N_760);
nor U5055 (N_5055,N_2049,N_2828);
nor U5056 (N_5056,N_681,N_1045);
nand U5057 (N_5057,N_2420,N_880);
nand U5058 (N_5058,N_1818,N_2641);
and U5059 (N_5059,N_2106,N_2444);
and U5060 (N_5060,N_30,N_275);
and U5061 (N_5061,N_972,N_1104);
and U5062 (N_5062,N_329,N_1932);
or U5063 (N_5063,N_2446,N_1331);
or U5064 (N_5064,N_1163,N_2848);
or U5065 (N_5065,N_369,N_1917);
and U5066 (N_5066,N_2044,N_2290);
and U5067 (N_5067,N_1854,N_1536);
nor U5068 (N_5068,N_1800,N_2077);
nor U5069 (N_5069,N_2612,N_994);
or U5070 (N_5070,N_1321,N_2614);
nor U5071 (N_5071,N_799,N_231);
or U5072 (N_5072,N_1468,N_2953);
nand U5073 (N_5073,N_2406,N_799);
nand U5074 (N_5074,N_1086,N_1873);
nand U5075 (N_5075,N_1529,N_2727);
nor U5076 (N_5076,N_174,N_589);
and U5077 (N_5077,N_2779,N_1128);
and U5078 (N_5078,N_790,N_2790);
and U5079 (N_5079,N_844,N_2919);
nand U5080 (N_5080,N_1879,N_1683);
xnor U5081 (N_5081,N_1698,N_1540);
and U5082 (N_5082,N_2924,N_2504);
or U5083 (N_5083,N_1952,N_632);
nand U5084 (N_5084,N_2428,N_32);
nand U5085 (N_5085,N_2942,N_326);
nand U5086 (N_5086,N_2359,N_1862);
nor U5087 (N_5087,N_2190,N_2035);
nor U5088 (N_5088,N_2751,N_2713);
nand U5089 (N_5089,N_1600,N_1636);
nand U5090 (N_5090,N_170,N_2412);
xnor U5091 (N_5091,N_1536,N_2617);
or U5092 (N_5092,N_1870,N_1250);
or U5093 (N_5093,N_2996,N_2031);
nor U5094 (N_5094,N_600,N_551);
or U5095 (N_5095,N_396,N_883);
nor U5096 (N_5096,N_1612,N_786);
nor U5097 (N_5097,N_2597,N_2313);
xnor U5098 (N_5098,N_1267,N_1550);
or U5099 (N_5099,N_13,N_2834);
nor U5100 (N_5100,N_2049,N_1427);
xnor U5101 (N_5101,N_1286,N_252);
and U5102 (N_5102,N_981,N_1764);
nand U5103 (N_5103,N_654,N_2867);
and U5104 (N_5104,N_858,N_1816);
nor U5105 (N_5105,N_606,N_1058);
or U5106 (N_5106,N_1839,N_2198);
nor U5107 (N_5107,N_1226,N_1987);
and U5108 (N_5108,N_1345,N_2882);
or U5109 (N_5109,N_2037,N_701);
and U5110 (N_5110,N_2905,N_1391);
nor U5111 (N_5111,N_2813,N_1581);
and U5112 (N_5112,N_233,N_653);
and U5113 (N_5113,N_2736,N_1457);
or U5114 (N_5114,N_2252,N_445);
or U5115 (N_5115,N_447,N_2736);
xnor U5116 (N_5116,N_2961,N_1403);
xor U5117 (N_5117,N_508,N_744);
or U5118 (N_5118,N_381,N_483);
nor U5119 (N_5119,N_2801,N_2955);
and U5120 (N_5120,N_1094,N_75);
nor U5121 (N_5121,N_1699,N_2689);
and U5122 (N_5122,N_558,N_447);
or U5123 (N_5123,N_2164,N_2197);
or U5124 (N_5124,N_1821,N_638);
nand U5125 (N_5125,N_1750,N_1227);
nand U5126 (N_5126,N_2491,N_2746);
nor U5127 (N_5127,N_1819,N_2762);
nor U5128 (N_5128,N_2370,N_176);
nor U5129 (N_5129,N_2102,N_1061);
and U5130 (N_5130,N_831,N_2550);
and U5131 (N_5131,N_1458,N_1530);
nand U5132 (N_5132,N_917,N_1649);
and U5133 (N_5133,N_1002,N_2899);
nor U5134 (N_5134,N_1425,N_2054);
nand U5135 (N_5135,N_1007,N_1003);
nand U5136 (N_5136,N_1904,N_2941);
and U5137 (N_5137,N_2760,N_6);
nand U5138 (N_5138,N_692,N_2758);
nor U5139 (N_5139,N_1302,N_2303);
nor U5140 (N_5140,N_2170,N_1247);
xnor U5141 (N_5141,N_2,N_304);
nand U5142 (N_5142,N_1538,N_2431);
nor U5143 (N_5143,N_2843,N_118);
and U5144 (N_5144,N_1868,N_320);
or U5145 (N_5145,N_2339,N_2695);
nor U5146 (N_5146,N_1730,N_1837);
and U5147 (N_5147,N_2537,N_407);
and U5148 (N_5148,N_2175,N_664);
xnor U5149 (N_5149,N_2051,N_1065);
and U5150 (N_5150,N_2848,N_1507);
nand U5151 (N_5151,N_2813,N_927);
nor U5152 (N_5152,N_708,N_337);
nand U5153 (N_5153,N_2542,N_2110);
nand U5154 (N_5154,N_2778,N_675);
nor U5155 (N_5155,N_2003,N_2237);
or U5156 (N_5156,N_2486,N_861);
nand U5157 (N_5157,N_2449,N_1539);
and U5158 (N_5158,N_2866,N_2673);
or U5159 (N_5159,N_706,N_2820);
and U5160 (N_5160,N_1534,N_1264);
nor U5161 (N_5161,N_1989,N_847);
nand U5162 (N_5162,N_1379,N_170);
or U5163 (N_5163,N_1702,N_1871);
nand U5164 (N_5164,N_1628,N_294);
or U5165 (N_5165,N_1024,N_1917);
and U5166 (N_5166,N_2043,N_1299);
nor U5167 (N_5167,N_1570,N_287);
nor U5168 (N_5168,N_992,N_1366);
and U5169 (N_5169,N_2783,N_2099);
nand U5170 (N_5170,N_184,N_1837);
nand U5171 (N_5171,N_2653,N_1829);
nor U5172 (N_5172,N_1028,N_379);
nand U5173 (N_5173,N_2174,N_2824);
nand U5174 (N_5174,N_2175,N_852);
and U5175 (N_5175,N_2928,N_2534);
or U5176 (N_5176,N_2612,N_2950);
nor U5177 (N_5177,N_2110,N_48);
or U5178 (N_5178,N_289,N_92);
nand U5179 (N_5179,N_49,N_324);
nand U5180 (N_5180,N_357,N_916);
nor U5181 (N_5181,N_612,N_548);
or U5182 (N_5182,N_1099,N_919);
xor U5183 (N_5183,N_1269,N_962);
xnor U5184 (N_5184,N_929,N_2610);
xnor U5185 (N_5185,N_2219,N_50);
and U5186 (N_5186,N_2424,N_2757);
and U5187 (N_5187,N_2847,N_1871);
or U5188 (N_5188,N_2739,N_1717);
and U5189 (N_5189,N_1578,N_1326);
nor U5190 (N_5190,N_2251,N_102);
nand U5191 (N_5191,N_2683,N_2385);
xor U5192 (N_5192,N_645,N_2329);
nor U5193 (N_5193,N_1206,N_357);
nand U5194 (N_5194,N_1606,N_2426);
nand U5195 (N_5195,N_607,N_1984);
and U5196 (N_5196,N_1273,N_2778);
or U5197 (N_5197,N_459,N_1247);
nand U5198 (N_5198,N_2965,N_1212);
or U5199 (N_5199,N_650,N_2997);
nor U5200 (N_5200,N_1971,N_20);
nor U5201 (N_5201,N_215,N_2112);
and U5202 (N_5202,N_2795,N_1733);
nand U5203 (N_5203,N_437,N_330);
and U5204 (N_5204,N_2446,N_2094);
and U5205 (N_5205,N_66,N_1492);
nor U5206 (N_5206,N_2234,N_1623);
nor U5207 (N_5207,N_520,N_2990);
and U5208 (N_5208,N_1616,N_2221);
or U5209 (N_5209,N_2185,N_1742);
or U5210 (N_5210,N_1034,N_812);
nor U5211 (N_5211,N_1225,N_392);
nand U5212 (N_5212,N_841,N_316);
nand U5213 (N_5213,N_2605,N_937);
and U5214 (N_5214,N_2100,N_87);
or U5215 (N_5215,N_1336,N_1794);
nand U5216 (N_5216,N_929,N_935);
xor U5217 (N_5217,N_1053,N_2381);
nand U5218 (N_5218,N_1903,N_1846);
or U5219 (N_5219,N_1404,N_459);
xnor U5220 (N_5220,N_1501,N_1293);
or U5221 (N_5221,N_2521,N_621);
nor U5222 (N_5222,N_1154,N_2402);
and U5223 (N_5223,N_2542,N_122);
nand U5224 (N_5224,N_2087,N_348);
or U5225 (N_5225,N_2691,N_1084);
xor U5226 (N_5226,N_2669,N_1506);
xnor U5227 (N_5227,N_2179,N_2007);
and U5228 (N_5228,N_1755,N_2213);
and U5229 (N_5229,N_2050,N_181);
or U5230 (N_5230,N_1145,N_1067);
nor U5231 (N_5231,N_596,N_2316);
nor U5232 (N_5232,N_2423,N_314);
nand U5233 (N_5233,N_2118,N_2618);
nand U5234 (N_5234,N_1074,N_617);
nand U5235 (N_5235,N_1091,N_813);
xnor U5236 (N_5236,N_1979,N_2999);
or U5237 (N_5237,N_1624,N_701);
and U5238 (N_5238,N_2667,N_245);
and U5239 (N_5239,N_2645,N_497);
xnor U5240 (N_5240,N_2529,N_273);
nor U5241 (N_5241,N_689,N_1466);
nand U5242 (N_5242,N_2699,N_1485);
or U5243 (N_5243,N_1101,N_42);
nand U5244 (N_5244,N_1849,N_2437);
and U5245 (N_5245,N_1714,N_100);
and U5246 (N_5246,N_565,N_1003);
and U5247 (N_5247,N_1887,N_2517);
and U5248 (N_5248,N_518,N_2661);
and U5249 (N_5249,N_1750,N_2140);
nor U5250 (N_5250,N_516,N_501);
xor U5251 (N_5251,N_376,N_2893);
and U5252 (N_5252,N_2243,N_1599);
and U5253 (N_5253,N_2090,N_708);
or U5254 (N_5254,N_118,N_489);
nor U5255 (N_5255,N_193,N_2198);
nand U5256 (N_5256,N_477,N_185);
nand U5257 (N_5257,N_1501,N_2229);
or U5258 (N_5258,N_2549,N_1632);
xnor U5259 (N_5259,N_1380,N_145);
nor U5260 (N_5260,N_1793,N_1276);
nand U5261 (N_5261,N_2934,N_1263);
nand U5262 (N_5262,N_1581,N_1005);
and U5263 (N_5263,N_695,N_170);
or U5264 (N_5264,N_2610,N_1419);
nor U5265 (N_5265,N_2683,N_1488);
and U5266 (N_5266,N_2253,N_2282);
or U5267 (N_5267,N_1110,N_2535);
nor U5268 (N_5268,N_80,N_1191);
xnor U5269 (N_5269,N_785,N_1235);
and U5270 (N_5270,N_1521,N_2561);
nor U5271 (N_5271,N_533,N_31);
xor U5272 (N_5272,N_197,N_650);
and U5273 (N_5273,N_1803,N_4);
nand U5274 (N_5274,N_959,N_1311);
nor U5275 (N_5275,N_1146,N_1987);
and U5276 (N_5276,N_1698,N_757);
nor U5277 (N_5277,N_708,N_2132);
and U5278 (N_5278,N_1504,N_627);
nor U5279 (N_5279,N_1796,N_1719);
nand U5280 (N_5280,N_1447,N_1529);
and U5281 (N_5281,N_1107,N_869);
nor U5282 (N_5282,N_845,N_2689);
nor U5283 (N_5283,N_1992,N_538);
or U5284 (N_5284,N_2325,N_2157);
nand U5285 (N_5285,N_1456,N_1384);
or U5286 (N_5286,N_426,N_1273);
nand U5287 (N_5287,N_882,N_1391);
xor U5288 (N_5288,N_2765,N_2222);
or U5289 (N_5289,N_1838,N_62);
or U5290 (N_5290,N_1933,N_877);
nand U5291 (N_5291,N_2889,N_1726);
and U5292 (N_5292,N_2936,N_996);
xor U5293 (N_5293,N_1152,N_808);
or U5294 (N_5294,N_937,N_1384);
and U5295 (N_5295,N_1371,N_1533);
nor U5296 (N_5296,N_1542,N_2120);
and U5297 (N_5297,N_1522,N_2264);
nand U5298 (N_5298,N_2002,N_1065);
or U5299 (N_5299,N_1015,N_2004);
and U5300 (N_5300,N_2953,N_662);
and U5301 (N_5301,N_2855,N_228);
or U5302 (N_5302,N_2889,N_1998);
xnor U5303 (N_5303,N_1686,N_2237);
nor U5304 (N_5304,N_187,N_1244);
nor U5305 (N_5305,N_2117,N_894);
nand U5306 (N_5306,N_2559,N_1457);
or U5307 (N_5307,N_2251,N_2057);
nor U5308 (N_5308,N_1431,N_1165);
nand U5309 (N_5309,N_1263,N_936);
nand U5310 (N_5310,N_1901,N_2654);
or U5311 (N_5311,N_1550,N_1437);
nor U5312 (N_5312,N_1827,N_1600);
nor U5313 (N_5313,N_1795,N_1303);
or U5314 (N_5314,N_1793,N_2123);
nor U5315 (N_5315,N_1461,N_1066);
nand U5316 (N_5316,N_2244,N_818);
and U5317 (N_5317,N_1496,N_2275);
and U5318 (N_5318,N_2233,N_1960);
and U5319 (N_5319,N_345,N_1942);
nor U5320 (N_5320,N_75,N_1231);
or U5321 (N_5321,N_2744,N_1098);
and U5322 (N_5322,N_2246,N_1300);
and U5323 (N_5323,N_1459,N_2621);
nor U5324 (N_5324,N_2760,N_1152);
or U5325 (N_5325,N_1080,N_1409);
nor U5326 (N_5326,N_805,N_416);
or U5327 (N_5327,N_170,N_2321);
or U5328 (N_5328,N_2638,N_547);
or U5329 (N_5329,N_405,N_1276);
or U5330 (N_5330,N_465,N_1307);
and U5331 (N_5331,N_2712,N_763);
and U5332 (N_5332,N_1549,N_2084);
or U5333 (N_5333,N_67,N_717);
or U5334 (N_5334,N_2463,N_1145);
and U5335 (N_5335,N_2849,N_549);
nor U5336 (N_5336,N_2116,N_2998);
or U5337 (N_5337,N_3,N_2307);
nand U5338 (N_5338,N_2187,N_2385);
and U5339 (N_5339,N_271,N_1488);
nor U5340 (N_5340,N_1484,N_2063);
nor U5341 (N_5341,N_1832,N_2447);
and U5342 (N_5342,N_98,N_2206);
nor U5343 (N_5343,N_1740,N_1666);
and U5344 (N_5344,N_1813,N_330);
or U5345 (N_5345,N_1563,N_643);
and U5346 (N_5346,N_925,N_2533);
or U5347 (N_5347,N_2718,N_1168);
and U5348 (N_5348,N_1403,N_1374);
nand U5349 (N_5349,N_1647,N_2222);
and U5350 (N_5350,N_1832,N_620);
and U5351 (N_5351,N_1902,N_1459);
nor U5352 (N_5352,N_2772,N_481);
nand U5353 (N_5353,N_1795,N_2899);
nand U5354 (N_5354,N_2296,N_2714);
and U5355 (N_5355,N_186,N_2494);
nor U5356 (N_5356,N_802,N_7);
xnor U5357 (N_5357,N_2236,N_568);
and U5358 (N_5358,N_1721,N_2071);
nand U5359 (N_5359,N_2906,N_2928);
nor U5360 (N_5360,N_2481,N_530);
nand U5361 (N_5361,N_487,N_1395);
or U5362 (N_5362,N_2829,N_1468);
or U5363 (N_5363,N_2992,N_2890);
or U5364 (N_5364,N_405,N_260);
nor U5365 (N_5365,N_2558,N_2128);
nor U5366 (N_5366,N_2849,N_482);
nor U5367 (N_5367,N_2858,N_2360);
nor U5368 (N_5368,N_890,N_181);
or U5369 (N_5369,N_498,N_348);
nor U5370 (N_5370,N_603,N_1882);
and U5371 (N_5371,N_2236,N_512);
and U5372 (N_5372,N_110,N_1830);
nand U5373 (N_5373,N_329,N_2030);
or U5374 (N_5374,N_619,N_1147);
and U5375 (N_5375,N_2240,N_1934);
nor U5376 (N_5376,N_831,N_131);
or U5377 (N_5377,N_1455,N_1192);
and U5378 (N_5378,N_411,N_3);
and U5379 (N_5379,N_1112,N_2805);
or U5380 (N_5380,N_19,N_2347);
and U5381 (N_5381,N_2401,N_1642);
nor U5382 (N_5382,N_987,N_1287);
nand U5383 (N_5383,N_343,N_2093);
or U5384 (N_5384,N_1982,N_1905);
xor U5385 (N_5385,N_2971,N_296);
xor U5386 (N_5386,N_559,N_2459);
nand U5387 (N_5387,N_975,N_1337);
nand U5388 (N_5388,N_955,N_112);
nand U5389 (N_5389,N_2816,N_2444);
or U5390 (N_5390,N_2428,N_846);
and U5391 (N_5391,N_2261,N_2601);
nor U5392 (N_5392,N_2706,N_510);
xor U5393 (N_5393,N_1995,N_981);
and U5394 (N_5394,N_1748,N_656);
nor U5395 (N_5395,N_1473,N_1911);
and U5396 (N_5396,N_1953,N_1443);
nor U5397 (N_5397,N_2498,N_2236);
or U5398 (N_5398,N_2006,N_1151);
nor U5399 (N_5399,N_634,N_1734);
nor U5400 (N_5400,N_986,N_1682);
and U5401 (N_5401,N_2028,N_2787);
nor U5402 (N_5402,N_2159,N_2431);
or U5403 (N_5403,N_2386,N_2776);
xor U5404 (N_5404,N_1257,N_510);
nor U5405 (N_5405,N_2553,N_1884);
nor U5406 (N_5406,N_194,N_207);
or U5407 (N_5407,N_2396,N_2154);
nand U5408 (N_5408,N_419,N_1553);
xor U5409 (N_5409,N_2182,N_775);
nand U5410 (N_5410,N_692,N_2136);
nand U5411 (N_5411,N_1903,N_1795);
nand U5412 (N_5412,N_1705,N_2116);
nor U5413 (N_5413,N_187,N_1701);
or U5414 (N_5414,N_55,N_1023);
nor U5415 (N_5415,N_1872,N_110);
and U5416 (N_5416,N_1180,N_2036);
nor U5417 (N_5417,N_1142,N_366);
or U5418 (N_5418,N_887,N_2674);
xor U5419 (N_5419,N_1645,N_1333);
nor U5420 (N_5420,N_2156,N_195);
nor U5421 (N_5421,N_2621,N_75);
nor U5422 (N_5422,N_2045,N_2635);
and U5423 (N_5423,N_901,N_1962);
nor U5424 (N_5424,N_1377,N_2446);
and U5425 (N_5425,N_1320,N_886);
nand U5426 (N_5426,N_582,N_2449);
nor U5427 (N_5427,N_1418,N_1053);
or U5428 (N_5428,N_1441,N_1226);
and U5429 (N_5429,N_925,N_1737);
or U5430 (N_5430,N_2163,N_2888);
nor U5431 (N_5431,N_471,N_2547);
xor U5432 (N_5432,N_1707,N_762);
or U5433 (N_5433,N_1714,N_2074);
or U5434 (N_5434,N_1829,N_577);
xor U5435 (N_5435,N_1611,N_85);
xnor U5436 (N_5436,N_112,N_2926);
or U5437 (N_5437,N_2851,N_1709);
or U5438 (N_5438,N_1404,N_2532);
nor U5439 (N_5439,N_2157,N_2006);
nor U5440 (N_5440,N_1642,N_493);
nand U5441 (N_5441,N_793,N_2454);
nand U5442 (N_5442,N_636,N_2403);
or U5443 (N_5443,N_2001,N_2253);
and U5444 (N_5444,N_2541,N_1206);
nor U5445 (N_5445,N_455,N_1847);
nor U5446 (N_5446,N_2454,N_1233);
nand U5447 (N_5447,N_250,N_237);
nor U5448 (N_5448,N_244,N_867);
and U5449 (N_5449,N_1113,N_1825);
or U5450 (N_5450,N_1259,N_1641);
xor U5451 (N_5451,N_2500,N_1544);
or U5452 (N_5452,N_2153,N_1180);
or U5453 (N_5453,N_2575,N_1942);
and U5454 (N_5454,N_37,N_1485);
or U5455 (N_5455,N_374,N_468);
and U5456 (N_5456,N_1640,N_2569);
or U5457 (N_5457,N_1409,N_460);
or U5458 (N_5458,N_2413,N_1074);
and U5459 (N_5459,N_45,N_1518);
and U5460 (N_5460,N_2715,N_2884);
or U5461 (N_5461,N_1928,N_478);
or U5462 (N_5462,N_1888,N_927);
xor U5463 (N_5463,N_594,N_1769);
nor U5464 (N_5464,N_2691,N_1678);
and U5465 (N_5465,N_2280,N_1839);
and U5466 (N_5466,N_2121,N_2230);
or U5467 (N_5467,N_1972,N_1298);
or U5468 (N_5468,N_573,N_1258);
xnor U5469 (N_5469,N_871,N_2724);
nand U5470 (N_5470,N_2328,N_2063);
nand U5471 (N_5471,N_2822,N_2086);
and U5472 (N_5472,N_1231,N_378);
xor U5473 (N_5473,N_802,N_219);
nor U5474 (N_5474,N_2008,N_1938);
nor U5475 (N_5475,N_234,N_1283);
or U5476 (N_5476,N_2045,N_1821);
and U5477 (N_5477,N_1392,N_2153);
or U5478 (N_5478,N_612,N_1005);
xnor U5479 (N_5479,N_457,N_929);
nand U5480 (N_5480,N_841,N_1669);
or U5481 (N_5481,N_1923,N_2972);
or U5482 (N_5482,N_2618,N_399);
or U5483 (N_5483,N_2109,N_758);
nand U5484 (N_5484,N_1082,N_590);
or U5485 (N_5485,N_2531,N_1707);
and U5486 (N_5486,N_2486,N_2699);
nor U5487 (N_5487,N_1860,N_2862);
and U5488 (N_5488,N_1199,N_350);
and U5489 (N_5489,N_1764,N_2168);
or U5490 (N_5490,N_48,N_874);
nor U5491 (N_5491,N_2173,N_1991);
nor U5492 (N_5492,N_1589,N_540);
nor U5493 (N_5493,N_896,N_1362);
nand U5494 (N_5494,N_410,N_1149);
nand U5495 (N_5495,N_1032,N_1736);
nand U5496 (N_5496,N_404,N_2268);
nand U5497 (N_5497,N_769,N_2841);
and U5498 (N_5498,N_1618,N_30);
xnor U5499 (N_5499,N_409,N_2595);
nand U5500 (N_5500,N_1331,N_2979);
nand U5501 (N_5501,N_1653,N_1042);
nor U5502 (N_5502,N_1132,N_946);
nand U5503 (N_5503,N_324,N_2042);
or U5504 (N_5504,N_1374,N_2668);
or U5505 (N_5505,N_1967,N_1179);
or U5506 (N_5506,N_2366,N_1714);
nor U5507 (N_5507,N_796,N_428);
nand U5508 (N_5508,N_2325,N_323);
nand U5509 (N_5509,N_2199,N_536);
nor U5510 (N_5510,N_1501,N_1409);
or U5511 (N_5511,N_1204,N_1159);
or U5512 (N_5512,N_2230,N_186);
xor U5513 (N_5513,N_860,N_175);
and U5514 (N_5514,N_62,N_859);
and U5515 (N_5515,N_843,N_319);
xnor U5516 (N_5516,N_1007,N_1100);
and U5517 (N_5517,N_998,N_1406);
and U5518 (N_5518,N_669,N_14);
nand U5519 (N_5519,N_271,N_1302);
nand U5520 (N_5520,N_2952,N_2696);
and U5521 (N_5521,N_2045,N_2567);
or U5522 (N_5522,N_99,N_89);
and U5523 (N_5523,N_1382,N_522);
nor U5524 (N_5524,N_339,N_958);
and U5525 (N_5525,N_2123,N_2690);
nand U5526 (N_5526,N_1753,N_2870);
and U5527 (N_5527,N_1748,N_417);
and U5528 (N_5528,N_389,N_1036);
nand U5529 (N_5529,N_1029,N_1066);
nor U5530 (N_5530,N_1426,N_2667);
nand U5531 (N_5531,N_1938,N_2704);
or U5532 (N_5532,N_1933,N_477);
and U5533 (N_5533,N_388,N_1457);
nand U5534 (N_5534,N_2112,N_458);
and U5535 (N_5535,N_311,N_1468);
nand U5536 (N_5536,N_2742,N_1308);
nand U5537 (N_5537,N_1945,N_1752);
or U5538 (N_5538,N_1534,N_635);
nand U5539 (N_5539,N_999,N_100);
or U5540 (N_5540,N_2366,N_806);
xor U5541 (N_5541,N_72,N_1492);
nor U5542 (N_5542,N_2391,N_1401);
nor U5543 (N_5543,N_794,N_915);
nand U5544 (N_5544,N_1961,N_246);
nand U5545 (N_5545,N_1588,N_100);
nor U5546 (N_5546,N_2832,N_1644);
nor U5547 (N_5547,N_1650,N_1639);
and U5548 (N_5548,N_1680,N_155);
xnor U5549 (N_5549,N_1716,N_2831);
and U5550 (N_5550,N_440,N_718);
nand U5551 (N_5551,N_2759,N_804);
nor U5552 (N_5552,N_314,N_1613);
or U5553 (N_5553,N_1160,N_953);
xor U5554 (N_5554,N_2383,N_159);
nor U5555 (N_5555,N_516,N_1861);
nand U5556 (N_5556,N_698,N_1547);
and U5557 (N_5557,N_1838,N_1409);
xor U5558 (N_5558,N_1537,N_2356);
and U5559 (N_5559,N_2847,N_907);
nand U5560 (N_5560,N_906,N_1810);
nand U5561 (N_5561,N_416,N_2258);
and U5562 (N_5562,N_1634,N_1088);
and U5563 (N_5563,N_2261,N_2172);
nor U5564 (N_5564,N_2173,N_2873);
and U5565 (N_5565,N_2881,N_2095);
xnor U5566 (N_5566,N_401,N_867);
and U5567 (N_5567,N_1687,N_95);
xnor U5568 (N_5568,N_89,N_2989);
and U5569 (N_5569,N_0,N_1422);
or U5570 (N_5570,N_2276,N_1956);
or U5571 (N_5571,N_595,N_2270);
nand U5572 (N_5572,N_2799,N_1409);
nand U5573 (N_5573,N_2508,N_95);
and U5574 (N_5574,N_723,N_240);
xor U5575 (N_5575,N_2581,N_32);
nor U5576 (N_5576,N_2259,N_1417);
or U5577 (N_5577,N_1015,N_237);
or U5578 (N_5578,N_231,N_451);
and U5579 (N_5579,N_1135,N_496);
nor U5580 (N_5580,N_2903,N_351);
or U5581 (N_5581,N_64,N_912);
or U5582 (N_5582,N_902,N_254);
and U5583 (N_5583,N_1435,N_2433);
or U5584 (N_5584,N_2610,N_2090);
and U5585 (N_5585,N_2118,N_582);
nor U5586 (N_5586,N_2706,N_1520);
and U5587 (N_5587,N_53,N_1316);
nor U5588 (N_5588,N_983,N_1766);
nand U5589 (N_5589,N_1335,N_168);
or U5590 (N_5590,N_2408,N_2043);
or U5591 (N_5591,N_250,N_316);
nand U5592 (N_5592,N_1227,N_2252);
nor U5593 (N_5593,N_2444,N_871);
nor U5594 (N_5594,N_443,N_1468);
nand U5595 (N_5595,N_238,N_2246);
xor U5596 (N_5596,N_45,N_1513);
and U5597 (N_5597,N_2914,N_2903);
and U5598 (N_5598,N_2797,N_1287);
nand U5599 (N_5599,N_225,N_2059);
or U5600 (N_5600,N_2504,N_2136);
xnor U5601 (N_5601,N_2827,N_1604);
or U5602 (N_5602,N_1731,N_653);
or U5603 (N_5603,N_175,N_1159);
and U5604 (N_5604,N_467,N_92);
and U5605 (N_5605,N_1908,N_1204);
or U5606 (N_5606,N_992,N_2997);
nor U5607 (N_5607,N_1891,N_1848);
and U5608 (N_5608,N_216,N_239);
nor U5609 (N_5609,N_2543,N_1708);
nand U5610 (N_5610,N_654,N_2416);
nand U5611 (N_5611,N_1640,N_272);
and U5612 (N_5612,N_2378,N_2458);
nor U5613 (N_5613,N_2516,N_777);
nand U5614 (N_5614,N_647,N_2626);
nand U5615 (N_5615,N_58,N_289);
nand U5616 (N_5616,N_533,N_2701);
xnor U5617 (N_5617,N_1409,N_494);
nor U5618 (N_5618,N_2285,N_1255);
nor U5619 (N_5619,N_1336,N_2254);
xnor U5620 (N_5620,N_18,N_2208);
nand U5621 (N_5621,N_642,N_1359);
nor U5622 (N_5622,N_369,N_2300);
nand U5623 (N_5623,N_334,N_2118);
nand U5624 (N_5624,N_1200,N_2559);
xnor U5625 (N_5625,N_2099,N_1459);
and U5626 (N_5626,N_1331,N_1685);
or U5627 (N_5627,N_2169,N_470);
and U5628 (N_5628,N_1172,N_345);
or U5629 (N_5629,N_281,N_254);
nor U5630 (N_5630,N_2167,N_1516);
nand U5631 (N_5631,N_1501,N_2721);
and U5632 (N_5632,N_2543,N_1719);
nand U5633 (N_5633,N_2537,N_2242);
or U5634 (N_5634,N_1105,N_594);
nand U5635 (N_5635,N_222,N_1412);
nor U5636 (N_5636,N_2814,N_1854);
and U5637 (N_5637,N_2543,N_2769);
or U5638 (N_5638,N_492,N_930);
and U5639 (N_5639,N_1050,N_268);
nand U5640 (N_5640,N_1699,N_2371);
and U5641 (N_5641,N_2144,N_203);
nand U5642 (N_5642,N_1070,N_26);
nor U5643 (N_5643,N_2230,N_1082);
nor U5644 (N_5644,N_2687,N_288);
and U5645 (N_5645,N_451,N_1761);
nand U5646 (N_5646,N_2235,N_1635);
or U5647 (N_5647,N_86,N_68);
nor U5648 (N_5648,N_2970,N_374);
nor U5649 (N_5649,N_1212,N_520);
nand U5650 (N_5650,N_2672,N_254);
or U5651 (N_5651,N_411,N_2737);
nand U5652 (N_5652,N_259,N_2079);
nand U5653 (N_5653,N_1767,N_2175);
nor U5654 (N_5654,N_969,N_1086);
nor U5655 (N_5655,N_2076,N_1386);
or U5656 (N_5656,N_2012,N_2649);
nor U5657 (N_5657,N_538,N_1517);
or U5658 (N_5658,N_45,N_852);
and U5659 (N_5659,N_113,N_1361);
or U5660 (N_5660,N_2138,N_1694);
nand U5661 (N_5661,N_1345,N_1180);
xor U5662 (N_5662,N_2356,N_942);
nor U5663 (N_5663,N_1420,N_2809);
or U5664 (N_5664,N_660,N_1225);
or U5665 (N_5665,N_2372,N_2825);
nand U5666 (N_5666,N_669,N_2903);
and U5667 (N_5667,N_310,N_470);
nor U5668 (N_5668,N_1940,N_2033);
or U5669 (N_5669,N_1577,N_2942);
and U5670 (N_5670,N_534,N_628);
xnor U5671 (N_5671,N_1746,N_90);
nor U5672 (N_5672,N_2151,N_1242);
nand U5673 (N_5673,N_31,N_1397);
and U5674 (N_5674,N_2524,N_1647);
and U5675 (N_5675,N_1102,N_2070);
nand U5676 (N_5676,N_572,N_2771);
and U5677 (N_5677,N_2978,N_2352);
nand U5678 (N_5678,N_2505,N_1229);
or U5679 (N_5679,N_2388,N_299);
xor U5680 (N_5680,N_833,N_672);
or U5681 (N_5681,N_470,N_862);
or U5682 (N_5682,N_2813,N_1061);
nand U5683 (N_5683,N_1203,N_143);
or U5684 (N_5684,N_820,N_267);
nor U5685 (N_5685,N_1009,N_1581);
and U5686 (N_5686,N_1881,N_2594);
nor U5687 (N_5687,N_2051,N_2325);
nand U5688 (N_5688,N_2887,N_137);
nor U5689 (N_5689,N_381,N_2316);
and U5690 (N_5690,N_82,N_871);
or U5691 (N_5691,N_132,N_1389);
nand U5692 (N_5692,N_1926,N_1018);
nor U5693 (N_5693,N_1377,N_885);
or U5694 (N_5694,N_1821,N_1190);
and U5695 (N_5695,N_1634,N_2090);
and U5696 (N_5696,N_455,N_1828);
xor U5697 (N_5697,N_180,N_1463);
nor U5698 (N_5698,N_1539,N_2458);
nand U5699 (N_5699,N_754,N_1415);
nor U5700 (N_5700,N_1259,N_1104);
nand U5701 (N_5701,N_1941,N_414);
nand U5702 (N_5702,N_2169,N_2640);
and U5703 (N_5703,N_2906,N_1910);
nor U5704 (N_5704,N_2890,N_1022);
and U5705 (N_5705,N_598,N_646);
nor U5706 (N_5706,N_1239,N_1139);
or U5707 (N_5707,N_1901,N_2577);
and U5708 (N_5708,N_1131,N_1117);
xor U5709 (N_5709,N_2086,N_1226);
nor U5710 (N_5710,N_2585,N_472);
nor U5711 (N_5711,N_2863,N_2551);
nor U5712 (N_5712,N_2846,N_1964);
and U5713 (N_5713,N_1534,N_1323);
or U5714 (N_5714,N_313,N_2266);
or U5715 (N_5715,N_380,N_477);
nor U5716 (N_5716,N_866,N_81);
nor U5717 (N_5717,N_138,N_1875);
and U5718 (N_5718,N_1176,N_343);
and U5719 (N_5719,N_2010,N_790);
or U5720 (N_5720,N_1472,N_2166);
nand U5721 (N_5721,N_1069,N_394);
xnor U5722 (N_5722,N_683,N_247);
nand U5723 (N_5723,N_768,N_356);
or U5724 (N_5724,N_1094,N_2157);
nor U5725 (N_5725,N_2082,N_1267);
nor U5726 (N_5726,N_1542,N_2594);
nand U5727 (N_5727,N_2777,N_252);
or U5728 (N_5728,N_267,N_1881);
and U5729 (N_5729,N_976,N_2492);
or U5730 (N_5730,N_911,N_338);
xor U5731 (N_5731,N_2787,N_1818);
nand U5732 (N_5732,N_1556,N_1068);
nor U5733 (N_5733,N_2103,N_115);
or U5734 (N_5734,N_1318,N_1277);
nor U5735 (N_5735,N_1921,N_2834);
or U5736 (N_5736,N_1639,N_444);
nor U5737 (N_5737,N_2059,N_678);
or U5738 (N_5738,N_2391,N_241);
or U5739 (N_5739,N_1580,N_794);
and U5740 (N_5740,N_47,N_2957);
nand U5741 (N_5741,N_2197,N_1568);
nand U5742 (N_5742,N_2661,N_1032);
nand U5743 (N_5743,N_1572,N_2972);
nand U5744 (N_5744,N_290,N_2047);
nor U5745 (N_5745,N_2064,N_1239);
nor U5746 (N_5746,N_2098,N_560);
xnor U5747 (N_5747,N_139,N_653);
or U5748 (N_5748,N_846,N_1465);
and U5749 (N_5749,N_710,N_883);
and U5750 (N_5750,N_748,N_506);
and U5751 (N_5751,N_1819,N_1291);
and U5752 (N_5752,N_773,N_128);
xor U5753 (N_5753,N_1923,N_1793);
or U5754 (N_5754,N_55,N_499);
or U5755 (N_5755,N_334,N_1185);
or U5756 (N_5756,N_826,N_1010);
and U5757 (N_5757,N_576,N_2094);
and U5758 (N_5758,N_2196,N_2183);
nand U5759 (N_5759,N_1286,N_1349);
nand U5760 (N_5760,N_1657,N_16);
or U5761 (N_5761,N_494,N_1335);
and U5762 (N_5762,N_1836,N_806);
and U5763 (N_5763,N_2864,N_1383);
nor U5764 (N_5764,N_300,N_146);
nand U5765 (N_5765,N_1698,N_963);
xnor U5766 (N_5766,N_2191,N_2474);
or U5767 (N_5767,N_422,N_1858);
and U5768 (N_5768,N_1577,N_381);
or U5769 (N_5769,N_476,N_401);
nor U5770 (N_5770,N_2751,N_1203);
nor U5771 (N_5771,N_2707,N_2837);
nor U5772 (N_5772,N_997,N_2870);
or U5773 (N_5773,N_2522,N_653);
nor U5774 (N_5774,N_794,N_1298);
and U5775 (N_5775,N_2835,N_1502);
nor U5776 (N_5776,N_950,N_1700);
nand U5777 (N_5777,N_1870,N_2406);
nor U5778 (N_5778,N_867,N_1727);
nand U5779 (N_5779,N_2384,N_1837);
xor U5780 (N_5780,N_1480,N_1197);
nand U5781 (N_5781,N_1975,N_1015);
and U5782 (N_5782,N_7,N_1490);
xnor U5783 (N_5783,N_2483,N_752);
nand U5784 (N_5784,N_2408,N_2666);
or U5785 (N_5785,N_1812,N_1544);
or U5786 (N_5786,N_661,N_43);
nand U5787 (N_5787,N_2678,N_1489);
and U5788 (N_5788,N_364,N_2795);
nand U5789 (N_5789,N_1557,N_1155);
xor U5790 (N_5790,N_1497,N_1121);
xor U5791 (N_5791,N_163,N_189);
and U5792 (N_5792,N_2,N_1031);
nor U5793 (N_5793,N_1512,N_1623);
or U5794 (N_5794,N_586,N_271);
nor U5795 (N_5795,N_605,N_367);
nor U5796 (N_5796,N_1870,N_2067);
xnor U5797 (N_5797,N_2598,N_2614);
and U5798 (N_5798,N_1138,N_1982);
nand U5799 (N_5799,N_24,N_733);
or U5800 (N_5800,N_2724,N_1325);
nand U5801 (N_5801,N_2020,N_979);
nor U5802 (N_5802,N_663,N_1600);
nor U5803 (N_5803,N_2332,N_2577);
nor U5804 (N_5804,N_696,N_2224);
nor U5805 (N_5805,N_2390,N_758);
nor U5806 (N_5806,N_533,N_2897);
nor U5807 (N_5807,N_2079,N_2864);
or U5808 (N_5808,N_1493,N_2436);
and U5809 (N_5809,N_1199,N_2155);
or U5810 (N_5810,N_1716,N_811);
nand U5811 (N_5811,N_174,N_1822);
nand U5812 (N_5812,N_261,N_1082);
nor U5813 (N_5813,N_2697,N_1642);
and U5814 (N_5814,N_2324,N_161);
or U5815 (N_5815,N_1552,N_1277);
and U5816 (N_5816,N_634,N_2858);
xnor U5817 (N_5817,N_1598,N_2958);
or U5818 (N_5818,N_14,N_2666);
and U5819 (N_5819,N_1688,N_2144);
nand U5820 (N_5820,N_1682,N_1013);
or U5821 (N_5821,N_2064,N_2849);
nand U5822 (N_5822,N_184,N_1805);
and U5823 (N_5823,N_1827,N_1268);
or U5824 (N_5824,N_607,N_478);
or U5825 (N_5825,N_2467,N_55);
and U5826 (N_5826,N_1789,N_219);
and U5827 (N_5827,N_178,N_2281);
and U5828 (N_5828,N_1947,N_2261);
xor U5829 (N_5829,N_480,N_2691);
xor U5830 (N_5830,N_1959,N_1813);
nor U5831 (N_5831,N_2912,N_1866);
and U5832 (N_5832,N_685,N_1984);
or U5833 (N_5833,N_2474,N_1880);
and U5834 (N_5834,N_2474,N_1335);
nand U5835 (N_5835,N_880,N_2472);
nor U5836 (N_5836,N_1630,N_2761);
nor U5837 (N_5837,N_888,N_462);
nor U5838 (N_5838,N_2540,N_1341);
and U5839 (N_5839,N_2434,N_2928);
xor U5840 (N_5840,N_862,N_941);
or U5841 (N_5841,N_600,N_1134);
nor U5842 (N_5842,N_2426,N_2263);
and U5843 (N_5843,N_2995,N_1497);
nor U5844 (N_5844,N_2689,N_1848);
nor U5845 (N_5845,N_2744,N_1258);
nor U5846 (N_5846,N_2673,N_417);
nand U5847 (N_5847,N_52,N_1413);
nand U5848 (N_5848,N_1733,N_1369);
and U5849 (N_5849,N_2126,N_258);
nand U5850 (N_5850,N_216,N_2708);
nor U5851 (N_5851,N_355,N_371);
or U5852 (N_5852,N_23,N_2449);
or U5853 (N_5853,N_938,N_636);
or U5854 (N_5854,N_191,N_279);
or U5855 (N_5855,N_2450,N_2580);
nor U5856 (N_5856,N_1836,N_1508);
nor U5857 (N_5857,N_2139,N_2168);
nor U5858 (N_5858,N_2257,N_2578);
nor U5859 (N_5859,N_1242,N_1642);
nand U5860 (N_5860,N_1815,N_2923);
xor U5861 (N_5861,N_111,N_2981);
nor U5862 (N_5862,N_2798,N_433);
or U5863 (N_5863,N_2215,N_1085);
nor U5864 (N_5864,N_2895,N_2877);
or U5865 (N_5865,N_1107,N_1292);
nand U5866 (N_5866,N_1059,N_2162);
or U5867 (N_5867,N_435,N_907);
nand U5868 (N_5868,N_1110,N_1163);
nand U5869 (N_5869,N_2996,N_1522);
xnor U5870 (N_5870,N_2444,N_1331);
nand U5871 (N_5871,N_145,N_1528);
nand U5872 (N_5872,N_804,N_201);
nor U5873 (N_5873,N_1397,N_2843);
or U5874 (N_5874,N_2986,N_2261);
or U5875 (N_5875,N_692,N_2268);
nand U5876 (N_5876,N_180,N_1594);
and U5877 (N_5877,N_1317,N_2439);
xor U5878 (N_5878,N_1308,N_2978);
nor U5879 (N_5879,N_6,N_1745);
xor U5880 (N_5880,N_2506,N_998);
or U5881 (N_5881,N_122,N_1021);
or U5882 (N_5882,N_1899,N_2701);
nor U5883 (N_5883,N_2334,N_1897);
or U5884 (N_5884,N_2632,N_1453);
nand U5885 (N_5885,N_567,N_2105);
or U5886 (N_5886,N_82,N_119);
and U5887 (N_5887,N_1183,N_1819);
and U5888 (N_5888,N_568,N_1943);
nand U5889 (N_5889,N_2297,N_2813);
xor U5890 (N_5890,N_1223,N_2052);
or U5891 (N_5891,N_1755,N_814);
or U5892 (N_5892,N_1337,N_790);
and U5893 (N_5893,N_2986,N_1321);
nor U5894 (N_5894,N_2040,N_1900);
and U5895 (N_5895,N_435,N_2251);
and U5896 (N_5896,N_2553,N_1803);
nand U5897 (N_5897,N_1888,N_1867);
and U5898 (N_5898,N_253,N_1096);
nand U5899 (N_5899,N_533,N_2730);
nor U5900 (N_5900,N_2086,N_122);
and U5901 (N_5901,N_2573,N_2963);
nor U5902 (N_5902,N_1709,N_1032);
or U5903 (N_5903,N_610,N_611);
and U5904 (N_5904,N_817,N_826);
or U5905 (N_5905,N_881,N_2043);
nor U5906 (N_5906,N_2449,N_350);
nand U5907 (N_5907,N_1503,N_380);
xor U5908 (N_5908,N_283,N_2093);
nand U5909 (N_5909,N_24,N_1091);
and U5910 (N_5910,N_1463,N_1679);
xor U5911 (N_5911,N_1389,N_2479);
xor U5912 (N_5912,N_2387,N_2041);
nand U5913 (N_5913,N_1141,N_627);
and U5914 (N_5914,N_1695,N_1344);
nand U5915 (N_5915,N_1668,N_2097);
and U5916 (N_5916,N_2073,N_2727);
or U5917 (N_5917,N_2878,N_1688);
nor U5918 (N_5918,N_2748,N_1659);
or U5919 (N_5919,N_2161,N_120);
and U5920 (N_5920,N_1615,N_1206);
nand U5921 (N_5921,N_2258,N_973);
or U5922 (N_5922,N_2565,N_1191);
and U5923 (N_5923,N_680,N_483);
nor U5924 (N_5924,N_1683,N_306);
and U5925 (N_5925,N_2338,N_1366);
or U5926 (N_5926,N_1062,N_2666);
nor U5927 (N_5927,N_582,N_349);
nand U5928 (N_5928,N_42,N_2542);
xnor U5929 (N_5929,N_427,N_1487);
xor U5930 (N_5930,N_2919,N_1699);
nor U5931 (N_5931,N_1063,N_2570);
nor U5932 (N_5932,N_2447,N_1363);
xor U5933 (N_5933,N_1491,N_1627);
nand U5934 (N_5934,N_1145,N_2834);
and U5935 (N_5935,N_2834,N_2933);
nand U5936 (N_5936,N_2583,N_1881);
nor U5937 (N_5937,N_2098,N_2117);
nor U5938 (N_5938,N_897,N_2214);
nor U5939 (N_5939,N_2233,N_1737);
or U5940 (N_5940,N_976,N_575);
nand U5941 (N_5941,N_555,N_2215);
nor U5942 (N_5942,N_1072,N_1688);
nor U5943 (N_5943,N_2394,N_2244);
xor U5944 (N_5944,N_1212,N_2544);
and U5945 (N_5945,N_2699,N_2828);
nand U5946 (N_5946,N_1412,N_1960);
nand U5947 (N_5947,N_1278,N_2824);
nor U5948 (N_5948,N_1321,N_2730);
or U5949 (N_5949,N_734,N_988);
or U5950 (N_5950,N_1278,N_528);
nand U5951 (N_5951,N_2745,N_46);
nand U5952 (N_5952,N_893,N_2304);
nand U5953 (N_5953,N_344,N_2947);
nor U5954 (N_5954,N_2627,N_2082);
or U5955 (N_5955,N_2765,N_2294);
nor U5956 (N_5956,N_2306,N_2910);
nor U5957 (N_5957,N_2691,N_2264);
or U5958 (N_5958,N_187,N_2884);
nand U5959 (N_5959,N_1707,N_890);
xnor U5960 (N_5960,N_781,N_583);
nor U5961 (N_5961,N_1293,N_2715);
and U5962 (N_5962,N_1000,N_627);
nor U5963 (N_5963,N_2309,N_1502);
nand U5964 (N_5964,N_738,N_1660);
or U5965 (N_5965,N_1372,N_2639);
nor U5966 (N_5966,N_1355,N_191);
or U5967 (N_5967,N_852,N_1900);
or U5968 (N_5968,N_963,N_685);
or U5969 (N_5969,N_2229,N_218);
and U5970 (N_5970,N_2333,N_1688);
or U5971 (N_5971,N_921,N_2767);
and U5972 (N_5972,N_626,N_162);
or U5973 (N_5973,N_2379,N_2842);
or U5974 (N_5974,N_124,N_1243);
nor U5975 (N_5975,N_1227,N_1372);
or U5976 (N_5976,N_9,N_2098);
nor U5977 (N_5977,N_868,N_1853);
or U5978 (N_5978,N_638,N_504);
nand U5979 (N_5979,N_475,N_1543);
and U5980 (N_5980,N_1891,N_2885);
nand U5981 (N_5981,N_900,N_434);
or U5982 (N_5982,N_2531,N_1116);
nor U5983 (N_5983,N_2116,N_2739);
and U5984 (N_5984,N_300,N_551);
nor U5985 (N_5985,N_741,N_875);
and U5986 (N_5986,N_1672,N_781);
nand U5987 (N_5987,N_353,N_1762);
or U5988 (N_5988,N_1027,N_2015);
nand U5989 (N_5989,N_1644,N_987);
xnor U5990 (N_5990,N_1876,N_483);
and U5991 (N_5991,N_2516,N_1914);
nand U5992 (N_5992,N_737,N_2771);
nor U5993 (N_5993,N_1611,N_422);
xnor U5994 (N_5994,N_2790,N_2747);
or U5995 (N_5995,N_1689,N_452);
and U5996 (N_5996,N_1912,N_2511);
xnor U5997 (N_5997,N_105,N_2140);
nand U5998 (N_5998,N_2454,N_1664);
xnor U5999 (N_5999,N_2512,N_2989);
nand U6000 (N_6000,N_5233,N_4402);
and U6001 (N_6001,N_5528,N_4260);
nor U6002 (N_6002,N_4337,N_3292);
or U6003 (N_6003,N_5683,N_5368);
nor U6004 (N_6004,N_4426,N_3851);
xnor U6005 (N_6005,N_5302,N_3414);
nand U6006 (N_6006,N_5345,N_4517);
or U6007 (N_6007,N_4524,N_3108);
or U6008 (N_6008,N_4803,N_3690);
or U6009 (N_6009,N_4725,N_5309);
and U6010 (N_6010,N_3712,N_3918);
nor U6011 (N_6011,N_5121,N_4492);
nor U6012 (N_6012,N_4660,N_5997);
or U6013 (N_6013,N_4903,N_4757);
nor U6014 (N_6014,N_4844,N_4230);
nand U6015 (N_6015,N_5999,N_3044);
or U6016 (N_6016,N_3728,N_4646);
xor U6017 (N_6017,N_3177,N_5787);
or U6018 (N_6018,N_3556,N_4314);
xnor U6019 (N_6019,N_5743,N_3087);
nand U6020 (N_6020,N_3542,N_4630);
or U6021 (N_6021,N_4760,N_5391);
nor U6022 (N_6022,N_5372,N_3833);
xnor U6023 (N_6023,N_5001,N_3760);
and U6024 (N_6024,N_5585,N_3591);
nand U6025 (N_6025,N_4752,N_5559);
nand U6026 (N_6026,N_3269,N_4419);
and U6027 (N_6027,N_4380,N_5489);
nand U6028 (N_6028,N_3603,N_3408);
nand U6029 (N_6029,N_4296,N_5061);
nand U6030 (N_6030,N_3447,N_5106);
or U6031 (N_6031,N_5171,N_4931);
xnor U6032 (N_6032,N_3321,N_3919);
or U6033 (N_6033,N_3621,N_3175);
or U6034 (N_6034,N_4675,N_5190);
and U6035 (N_6035,N_3140,N_3187);
nor U6036 (N_6036,N_3575,N_3901);
and U6037 (N_6037,N_3758,N_4773);
or U6038 (N_6038,N_3407,N_5782);
nand U6039 (N_6039,N_5568,N_3642);
and U6040 (N_6040,N_3295,N_5055);
and U6041 (N_6041,N_3643,N_5367);
and U6042 (N_6042,N_4043,N_3331);
and U6043 (N_6043,N_4800,N_3368);
and U6044 (N_6044,N_3171,N_3877);
and U6045 (N_6045,N_3644,N_4326);
nand U6046 (N_6046,N_3845,N_3344);
nand U6047 (N_6047,N_4627,N_4123);
nand U6048 (N_6048,N_3191,N_5826);
xor U6049 (N_6049,N_3064,N_4245);
nand U6050 (N_6050,N_5040,N_3155);
and U6051 (N_6051,N_3325,N_3518);
or U6052 (N_6052,N_3464,N_5948);
or U6053 (N_6053,N_5729,N_5886);
nor U6054 (N_6054,N_4420,N_3489);
or U6055 (N_6055,N_3415,N_4160);
and U6056 (N_6056,N_3126,N_3821);
and U6057 (N_6057,N_5242,N_5870);
xnor U6058 (N_6058,N_5664,N_4862);
nand U6059 (N_6059,N_4078,N_4340);
nor U6060 (N_6060,N_4716,N_3737);
nand U6061 (N_6061,N_5764,N_4632);
and U6062 (N_6062,N_5910,N_4553);
nand U6063 (N_6063,N_5103,N_3498);
nor U6064 (N_6064,N_5926,N_5861);
or U6065 (N_6065,N_4051,N_4892);
or U6066 (N_6066,N_5735,N_5689);
and U6067 (N_6067,N_4568,N_4379);
nand U6068 (N_6068,N_3239,N_3079);
xor U6069 (N_6069,N_3638,N_5370);
and U6070 (N_6070,N_4277,N_4201);
nor U6071 (N_6071,N_3063,N_3990);
and U6072 (N_6072,N_4073,N_4166);
nand U6073 (N_6073,N_4698,N_5941);
nand U6074 (N_6074,N_4182,N_3858);
nand U6075 (N_6075,N_4343,N_5324);
nor U6076 (N_6076,N_5537,N_4584);
or U6077 (N_6077,N_5621,N_3396);
and U6078 (N_6078,N_5165,N_4672);
and U6079 (N_6079,N_5726,N_4055);
xnor U6080 (N_6080,N_4975,N_3127);
xnor U6081 (N_6081,N_5730,N_3247);
and U6082 (N_6082,N_5600,N_4830);
and U6083 (N_6083,N_5665,N_5245);
nand U6084 (N_6084,N_4465,N_3099);
xnor U6085 (N_6085,N_4651,N_4662);
and U6086 (N_6086,N_5771,N_5047);
nand U6087 (N_6087,N_5656,N_5339);
and U6088 (N_6088,N_4572,N_5202);
and U6089 (N_6089,N_3262,N_4585);
and U6090 (N_6090,N_5393,N_3328);
or U6091 (N_6091,N_3049,N_3101);
nor U6092 (N_6092,N_5752,N_3549);
nor U6093 (N_6093,N_4140,N_4767);
nand U6094 (N_6094,N_4994,N_5863);
or U6095 (N_6095,N_3592,N_3504);
nor U6096 (N_6096,N_5108,N_4816);
or U6097 (N_6097,N_3873,N_3445);
nand U6098 (N_6098,N_4555,N_4566);
and U6099 (N_6099,N_3452,N_4837);
nor U6100 (N_6100,N_4839,N_4152);
nor U6101 (N_6101,N_3991,N_3503);
or U6102 (N_6102,N_4414,N_3154);
xnor U6103 (N_6103,N_3293,N_3037);
nand U6104 (N_6104,N_5150,N_5510);
nand U6105 (N_6105,N_3029,N_4557);
nor U6106 (N_6106,N_3531,N_5456);
or U6107 (N_6107,N_4470,N_3691);
nor U6108 (N_6108,N_3680,N_5298);
or U6109 (N_6109,N_5535,N_5359);
xor U6110 (N_6110,N_3189,N_5971);
or U6111 (N_6111,N_3032,N_3455);
nor U6112 (N_6112,N_3273,N_4149);
nor U6113 (N_6113,N_5919,N_4597);
or U6114 (N_6114,N_4375,N_4915);
or U6115 (N_6115,N_3750,N_5337);
and U6116 (N_6116,N_4951,N_3905);
nor U6117 (N_6117,N_4439,N_3280);
and U6118 (N_6118,N_5360,N_5855);
xnor U6119 (N_6119,N_4818,N_4466);
nand U6120 (N_6120,N_5525,N_3228);
xnor U6121 (N_6121,N_3499,N_5966);
nand U6122 (N_6122,N_5675,N_5566);
nor U6123 (N_6123,N_4449,N_4594);
xor U6124 (N_6124,N_4516,N_4993);
or U6125 (N_6125,N_5305,N_3904);
and U6126 (N_6126,N_4367,N_3791);
nor U6127 (N_6127,N_3539,N_3852);
or U6128 (N_6128,N_5868,N_5482);
or U6129 (N_6129,N_4709,N_3220);
or U6130 (N_6130,N_3875,N_4985);
nand U6131 (N_6131,N_4522,N_3304);
and U6132 (N_6132,N_5728,N_3115);
and U6133 (N_6133,N_3254,N_4718);
nor U6134 (N_6134,N_3695,N_4612);
nor U6135 (N_6135,N_4741,N_3561);
xnor U6136 (N_6136,N_3011,N_5292);
nor U6137 (N_6137,N_3552,N_4783);
nor U6138 (N_6138,N_3959,N_4219);
xor U6139 (N_6139,N_3129,N_3743);
nor U6140 (N_6140,N_3672,N_5802);
xnor U6141 (N_6141,N_5267,N_5043);
and U6142 (N_6142,N_3020,N_3217);
xnor U6143 (N_6143,N_3496,N_5934);
nand U6144 (N_6144,N_3299,N_3401);
and U6145 (N_6145,N_3738,N_5832);
or U6146 (N_6146,N_5662,N_4722);
xnor U6147 (N_6147,N_5167,N_4657);
nand U6148 (N_6148,N_4527,N_4387);
nor U6149 (N_6149,N_5085,N_5490);
or U6150 (N_6150,N_4050,N_4864);
or U6151 (N_6151,N_5046,N_4826);
nand U6152 (N_6152,N_3306,N_4059);
nor U6153 (N_6153,N_5842,N_5457);
nor U6154 (N_6154,N_5590,N_5024);
nand U6155 (N_6155,N_3416,N_5307);
nand U6156 (N_6156,N_5288,N_3409);
nor U6157 (N_6157,N_4040,N_4445);
or U6158 (N_6158,N_5351,N_5386);
nand U6159 (N_6159,N_4952,N_5443);
nand U6160 (N_6160,N_4537,N_4444);
and U6161 (N_6161,N_3437,N_3716);
nand U6162 (N_6162,N_3628,N_5821);
xnor U6163 (N_6163,N_5991,N_3656);
and U6164 (N_6164,N_4007,N_3137);
or U6165 (N_6165,N_4857,N_4834);
nor U6166 (N_6166,N_3072,N_4887);
nor U6167 (N_6167,N_3080,N_4755);
nor U6168 (N_6168,N_5979,N_3448);
nand U6169 (N_6169,N_5349,N_5059);
nand U6170 (N_6170,N_3967,N_5952);
and U6171 (N_6171,N_3000,N_5033);
nand U6172 (N_6172,N_4960,N_3847);
nand U6173 (N_6173,N_3505,N_3146);
or U6174 (N_6174,N_5994,N_4796);
nor U6175 (N_6175,N_5446,N_5332);
and U6176 (N_6176,N_3889,N_3138);
xor U6177 (N_6177,N_4883,N_3418);
xor U6178 (N_6178,N_5240,N_4141);
or U6179 (N_6179,N_4401,N_3966);
nor U6180 (N_6180,N_4407,N_5776);
or U6181 (N_6181,N_4114,N_5481);
and U6182 (N_6182,N_4649,N_5811);
nand U6183 (N_6183,N_4884,N_4103);
or U6184 (N_6184,N_5008,N_3491);
or U6185 (N_6185,N_5834,N_4167);
nand U6186 (N_6186,N_4028,N_5485);
or U6187 (N_6187,N_5904,N_4731);
and U6188 (N_6188,N_5617,N_3082);
and U6189 (N_6189,N_4045,N_4094);
nand U6190 (N_6190,N_3669,N_3679);
or U6191 (N_6191,N_4569,N_5875);
xnor U6192 (N_6192,N_3394,N_5714);
and U6193 (N_6193,N_3349,N_3604);
nor U6194 (N_6194,N_3693,N_3593);
nand U6195 (N_6195,N_5918,N_3182);
nand U6196 (N_6196,N_5101,N_3620);
nor U6197 (N_6197,N_5291,N_3653);
and U6198 (N_6198,N_3783,N_3970);
nand U6199 (N_6199,N_5218,N_5563);
and U6200 (N_6200,N_3098,N_5711);
or U6201 (N_6201,N_4986,N_3454);
or U6202 (N_6202,N_3497,N_3666);
nor U6203 (N_6203,N_4183,N_5287);
and U6204 (N_6204,N_3759,N_5756);
and U6205 (N_6205,N_3757,N_5416);
nand U6206 (N_6206,N_4575,N_4270);
nand U6207 (N_6207,N_5417,N_3264);
or U6208 (N_6208,N_5920,N_4408);
and U6209 (N_6209,N_4081,N_4500);
nand U6210 (N_6210,N_4604,N_4618);
nand U6211 (N_6211,N_3864,N_5791);
or U6212 (N_6212,N_3219,N_4482);
nand U6213 (N_6213,N_5399,N_3085);
and U6214 (N_6214,N_5118,N_3937);
and U6215 (N_6215,N_3869,N_4392);
nor U6216 (N_6216,N_4274,N_5125);
and U6217 (N_6217,N_5956,N_3233);
nand U6218 (N_6218,N_5885,N_3198);
and U6219 (N_6219,N_5820,N_3086);
nand U6220 (N_6220,N_4089,N_5573);
and U6221 (N_6221,N_3244,N_3466);
or U6222 (N_6222,N_3152,N_5951);
nand U6223 (N_6223,N_4002,N_4224);
nor U6224 (N_6224,N_5471,N_3962);
nor U6225 (N_6225,N_5463,N_5676);
nor U6226 (N_6226,N_3008,N_3661);
and U6227 (N_6227,N_5915,N_4308);
and U6228 (N_6228,N_5965,N_3957);
and U6229 (N_6229,N_4368,N_4806);
or U6230 (N_6230,N_4652,N_4980);
and U6231 (N_6231,N_5803,N_3659);
or U6232 (N_6232,N_3793,N_3381);
or U6233 (N_6233,N_3494,N_3482);
or U6234 (N_6234,N_4708,N_3402);
nand U6235 (N_6235,N_3802,N_5807);
nand U6236 (N_6236,N_5587,N_5320);
or U6237 (N_6237,N_4240,N_5769);
and U6238 (N_6238,N_4582,N_4679);
nand U6239 (N_6239,N_5284,N_4345);
or U6240 (N_6240,N_5459,N_3316);
nor U6241 (N_6241,N_5111,N_4513);
nor U6242 (N_6242,N_4289,N_3799);
and U6243 (N_6243,N_4782,N_3151);
or U6244 (N_6244,N_4588,N_3610);
nand U6245 (N_6245,N_5051,N_5686);
xnor U6246 (N_6246,N_4925,N_5840);
and U6247 (N_6247,N_4893,N_5565);
or U6248 (N_6248,N_3781,N_4619);
and U6249 (N_6249,N_5596,N_3710);
nand U6250 (N_6250,N_3551,N_3277);
nand U6251 (N_6251,N_5308,N_5330);
xor U6252 (N_6252,N_5524,N_3065);
nor U6253 (N_6253,N_3472,N_3136);
or U6254 (N_6254,N_3023,N_5445);
xor U6255 (N_6255,N_4822,N_5015);
and U6256 (N_6256,N_5819,N_3289);
and U6257 (N_6257,N_4727,N_5846);
and U6258 (N_6258,N_3536,N_3211);
or U6259 (N_6259,N_3600,N_5458);
nand U6260 (N_6260,N_4906,N_3492);
or U6261 (N_6261,N_5251,N_4199);
nor U6262 (N_6262,N_5579,N_3263);
nor U6263 (N_6263,N_4019,N_4876);
nor U6264 (N_6264,N_5488,N_5042);
and U6265 (N_6265,N_4587,N_5311);
nand U6266 (N_6266,N_5206,N_3131);
nand U6267 (N_6267,N_3083,N_3203);
nor U6268 (N_6268,N_3558,N_3458);
nor U6269 (N_6269,N_4010,N_4840);
and U6270 (N_6270,N_5060,N_3382);
nor U6271 (N_6271,N_3365,N_3446);
nand U6272 (N_6272,N_5243,N_4335);
or U6273 (N_6273,N_4736,N_3726);
nand U6274 (N_6274,N_4694,N_4236);
or U6275 (N_6275,N_4382,N_5007);
and U6276 (N_6276,N_4153,N_4281);
nor U6277 (N_6277,N_3166,N_3846);
nand U6278 (N_6278,N_5020,N_3808);
or U6279 (N_6279,N_5583,N_4902);
nor U6280 (N_6280,N_4677,N_3804);
nand U6281 (N_6281,N_3910,N_4968);
or U6282 (N_6282,N_3976,N_5938);
nor U6283 (N_6283,N_3606,N_4285);
and U6284 (N_6284,N_5631,N_4122);
nand U6285 (N_6285,N_3145,N_5606);
nor U6286 (N_6286,N_4520,N_5589);
and U6287 (N_6287,N_3731,N_3839);
nor U6288 (N_6288,N_5452,N_5312);
xor U6289 (N_6289,N_3607,N_4080);
and U6290 (N_6290,N_4739,N_4601);
or U6291 (N_6291,N_3256,N_4771);
xor U6292 (N_6292,N_3216,N_4640);
nand U6293 (N_6293,N_5653,N_4944);
xor U6294 (N_6294,N_4713,N_4777);
and U6295 (N_6295,N_3309,N_5197);
and U6296 (N_6296,N_4135,N_5173);
nor U6297 (N_6297,N_4415,N_3983);
nand U6298 (N_6298,N_5031,N_5232);
and U6299 (N_6299,N_3865,N_4854);
and U6300 (N_6300,N_5113,N_5790);
nor U6301 (N_6301,N_5502,N_3942);
nand U6302 (N_6302,N_4674,N_3232);
or U6303 (N_6303,N_5044,N_4247);
and U6304 (N_6304,N_5361,N_3279);
or U6305 (N_6305,N_4064,N_5858);
or U6306 (N_6306,N_3426,N_3487);
or U6307 (N_6307,N_3729,N_4728);
and U6308 (N_6308,N_4702,N_3794);
nand U6309 (N_6309,N_5102,N_5911);
and U6310 (N_6310,N_4033,N_5239);
nand U6311 (N_6311,N_5380,N_3378);
xnor U6312 (N_6312,N_3436,N_4364);
nor U6313 (N_6313,N_3837,N_4507);
nand U6314 (N_6314,N_3350,N_3343);
and U6315 (N_6315,N_5430,N_4614);
nand U6316 (N_6316,N_5246,N_5969);
nor U6317 (N_6317,N_3868,N_4106);
and U6318 (N_6318,N_5112,N_4879);
or U6319 (N_6319,N_3921,N_3719);
nand U6320 (N_6320,N_5747,N_5972);
and U6321 (N_6321,N_4999,N_4726);
nand U6322 (N_6322,N_3158,N_3281);
and U6323 (N_6323,N_4363,N_5141);
nand U6324 (N_6324,N_3897,N_3894);
xor U6325 (N_6325,N_5555,N_5140);
or U6326 (N_6326,N_4433,N_3595);
and U6327 (N_6327,N_4406,N_5947);
nand U6328 (N_6328,N_5304,N_4961);
and U6329 (N_6329,N_4813,N_5572);
and U6330 (N_6330,N_5758,N_4100);
and U6331 (N_6331,N_5654,N_3334);
and U6332 (N_6332,N_3355,N_5013);
nand U6333 (N_6333,N_4720,N_4996);
xor U6334 (N_6334,N_4548,N_4322);
xnor U6335 (N_6335,N_3625,N_4061);
and U6336 (N_6336,N_5827,N_3134);
nor U6337 (N_6337,N_4328,N_3914);
and U6338 (N_6338,N_4788,N_3611);
xor U6339 (N_6339,N_3547,N_5815);
and U6340 (N_6340,N_4290,N_4983);
nor U6341 (N_6341,N_5757,N_5741);
nor U6342 (N_6342,N_4859,N_5878);
and U6343 (N_6343,N_5666,N_4888);
nand U6344 (N_6344,N_5039,N_5017);
nor U6345 (N_6345,N_5301,N_3576);
or U6346 (N_6346,N_4110,N_4339);
and U6347 (N_6347,N_5179,N_3697);
nor U6348 (N_6348,N_4850,N_5494);
and U6349 (N_6349,N_5375,N_5453);
and U6350 (N_6350,N_4044,N_5745);
nor U6351 (N_6351,N_5196,N_3261);
and U6352 (N_6352,N_4855,N_3946);
nor U6353 (N_6353,N_4742,N_4596);
or U6354 (N_6354,N_4734,N_4173);
or U6355 (N_6355,N_5696,N_5483);
xor U6356 (N_6356,N_3753,N_3582);
nand U6357 (N_6357,N_3734,N_3874);
xnor U6358 (N_6358,N_5241,N_3500);
nor U6359 (N_6359,N_4851,N_3057);
nand U6360 (N_6360,N_4391,N_3287);
xnor U6361 (N_6361,N_5469,N_3112);
or U6362 (N_6362,N_3391,N_5219);
nor U6363 (N_6363,N_5867,N_3773);
nand U6364 (N_6364,N_5774,N_4307);
or U6365 (N_6365,N_3276,N_5503);
or U6366 (N_6366,N_5329,N_5333);
or U6367 (N_6367,N_5680,N_4286);
or U6368 (N_6368,N_4827,N_3641);
nand U6369 (N_6369,N_3372,N_4536);
nand U6370 (N_6370,N_3824,N_5522);
nand U6371 (N_6371,N_3570,N_5176);
nor U6372 (N_6372,N_4292,N_5006);
or U6373 (N_6373,N_5424,N_5500);
nand U6374 (N_6374,N_4443,N_5152);
or U6375 (N_6375,N_4399,N_4676);
nor U6376 (N_6376,N_5561,N_5772);
xnor U6377 (N_6377,N_3811,N_4222);
and U6378 (N_6378,N_5069,N_5900);
nand U6379 (N_6379,N_3163,N_5130);
nor U6380 (N_6380,N_3985,N_5210);
and U6381 (N_6381,N_3143,N_5721);
nor U6382 (N_6382,N_5005,N_3473);
and U6383 (N_6383,N_4977,N_5449);
nand U6384 (N_6384,N_4478,N_3827);
nor U6385 (N_6385,N_4769,N_5843);
and U6386 (N_6386,N_3483,N_5408);
nor U6387 (N_6387,N_5731,N_3825);
nand U6388 (N_6388,N_3968,N_5135);
xor U6389 (N_6389,N_3829,N_3853);
or U6390 (N_6390,N_4098,N_4776);
or U6391 (N_6391,N_3924,N_3311);
xor U6392 (N_6392,N_4795,N_5259);
nand U6393 (N_6393,N_5922,N_4559);
nor U6394 (N_6394,N_5086,N_4268);
nand U6395 (N_6395,N_5993,N_4016);
and U6396 (N_6396,N_4001,N_4483);
nand U6397 (N_6397,N_4144,N_4271);
nor U6398 (N_6398,N_4000,N_4504);
and U6399 (N_6399,N_5973,N_5073);
nand U6400 (N_6400,N_3400,N_5497);
nand U6401 (N_6401,N_4872,N_4609);
nor U6402 (N_6402,N_5250,N_4987);
nor U6403 (N_6403,N_4086,N_5157);
xnor U6404 (N_6404,N_4519,N_4819);
or U6405 (N_6405,N_5213,N_5340);
nor U6406 (N_6406,N_3980,N_4869);
or U6407 (N_6407,N_5521,N_4197);
or U6408 (N_6408,N_5174,N_3260);
nor U6409 (N_6409,N_3928,N_4206);
and U6410 (N_6410,N_3945,N_4956);
and U6411 (N_6411,N_4486,N_5134);
and U6412 (N_6412,N_3297,N_5464);
nand U6413 (N_6413,N_5890,N_4969);
nor U6414 (N_6414,N_3231,N_4785);
and U6415 (N_6415,N_4416,N_3623);
and U6416 (N_6416,N_4057,N_5831);
or U6417 (N_6417,N_5607,N_3673);
nor U6418 (N_6418,N_5306,N_4860);
and U6419 (N_6419,N_5433,N_4914);
nand U6420 (N_6420,N_5734,N_4992);
or U6421 (N_6421,N_5530,N_4095);
xor U6422 (N_6422,N_4654,N_4309);
and U6423 (N_6423,N_3885,N_4272);
or U6424 (N_6424,N_3006,N_5688);
xor U6425 (N_6425,N_3883,N_4658);
xnor U6426 (N_6426,N_5860,N_3373);
and U6427 (N_6427,N_4828,N_4241);
or U6428 (N_6428,N_4802,N_5836);
nand U6429 (N_6429,N_3950,N_3823);
and U6430 (N_6430,N_3649,N_3588);
or U6431 (N_6431,N_4984,N_4801);
or U6432 (N_6432,N_4125,N_4038);
and U6433 (N_6433,N_5877,N_5071);
nor U6434 (N_6434,N_3067,N_4495);
nand U6435 (N_6435,N_3568,N_5859);
xnor U6436 (N_6436,N_3480,N_5833);
or U6437 (N_6437,N_4683,N_5949);
or U6438 (N_6438,N_3174,N_5358);
and U6439 (N_6439,N_5623,N_4120);
and U6440 (N_6440,N_3490,N_5271);
and U6441 (N_6441,N_4323,N_3526);
and U6442 (N_6442,N_5207,N_4283);
xor U6443 (N_6443,N_5545,N_3453);
xor U6444 (N_6444,N_5062,N_4481);
nand U6445 (N_6445,N_3954,N_5401);
xnor U6446 (N_6446,N_3535,N_4901);
or U6447 (N_6447,N_4128,N_4409);
and U6448 (N_6448,N_3417,N_5549);
and U6449 (N_6449,N_3486,N_3544);
nor U6450 (N_6450,N_4162,N_5099);
xor U6451 (N_6451,N_4253,N_5603);
xnor U6452 (N_6452,N_5512,N_4468);
or U6453 (N_6453,N_3806,N_3363);
nor U6454 (N_6454,N_5074,N_4209);
or U6455 (N_6455,N_4824,N_4200);
nand U6456 (N_6456,N_3943,N_3813);
nor U6457 (N_6457,N_5737,N_5775);
nand U6458 (N_6458,N_3533,N_5850);
and U6459 (N_6459,N_4633,N_3675);
or U6460 (N_6460,N_4347,N_5905);
nand U6461 (N_6461,N_3699,N_4234);
nand U6462 (N_6462,N_3249,N_5880);
nand U6463 (N_6463,N_5170,N_4320);
and U6464 (N_6464,N_4306,N_5188);
nand U6465 (N_6465,N_3925,N_4330);
nor U6466 (N_6466,N_5397,N_5199);
and U6467 (N_6467,N_5933,N_4910);
nand U6468 (N_6468,N_4325,N_3303);
or U6469 (N_6469,N_5209,N_5705);
nand U6470 (N_6470,N_4208,N_5322);
nand U6471 (N_6471,N_3988,N_5857);
nor U6472 (N_6472,N_3347,N_3613);
or U6473 (N_6473,N_4025,N_5493);
nor U6474 (N_6474,N_4212,N_4079);
or U6475 (N_6475,N_4539,N_5194);
or U6476 (N_6476,N_5009,N_4266);
nor U6477 (N_6477,N_5873,N_4087);
nor U6478 (N_6478,N_3708,N_4052);
nand U6479 (N_6479,N_3936,N_4461);
or U6480 (N_6480,N_5420,N_3393);
nand U6481 (N_6481,N_5781,N_4549);
and U6482 (N_6482,N_4229,N_3040);
and U6483 (N_6483,N_4273,N_3428);
nand U6484 (N_6484,N_5768,N_3161);
nor U6485 (N_6485,N_4502,N_3411);
and U6486 (N_6486,N_4484,N_4838);
nor U6487 (N_6487,N_5988,N_4175);
nand U6488 (N_6488,N_3056,N_4610);
and U6489 (N_6489,N_5618,N_5917);
nor U6490 (N_6490,N_3388,N_5200);
nand U6491 (N_6491,N_4579,N_4397);
and U6492 (N_6492,N_3252,N_3369);
or U6493 (N_6493,N_4946,N_5037);
nor U6494 (N_6494,N_4678,N_3308);
and U6495 (N_6495,N_3749,N_5182);
and U6496 (N_6496,N_3527,N_5789);
and U6497 (N_6497,N_3207,N_4003);
nand U6498 (N_6498,N_4378,N_4832);
nor U6499 (N_6499,N_3070,N_3036);
nor U6500 (N_6500,N_5110,N_3450);
nor U6501 (N_6501,N_5404,N_3682);
nand U6502 (N_6502,N_3961,N_3090);
or U6503 (N_6503,N_5395,N_5431);
and U6504 (N_6504,N_5338,N_4070);
nand U6505 (N_6505,N_4259,N_5817);
and U6506 (N_6506,N_5963,N_5169);
nor U6507 (N_6507,N_3340,N_4265);
nor U6508 (N_6508,N_4552,N_3844);
nor U6509 (N_6509,N_3412,N_5475);
or U6510 (N_6510,N_5981,N_5315);
or U6511 (N_6511,N_4279,N_4185);
or U6512 (N_6512,N_3553,N_3550);
or U6513 (N_6513,N_3474,N_5082);
nor U6514 (N_6514,N_4192,N_5185);
xnor U6515 (N_6515,N_5263,N_3030);
nor U6516 (N_6516,N_5432,N_3380);
and U6517 (N_6517,N_5793,N_4267);
nor U6518 (N_6518,N_5286,N_5189);
nand U6519 (N_6519,N_5848,N_4176);
nand U6520 (N_6520,N_5706,N_3270);
and U6521 (N_6521,N_5844,N_5788);
nor U6522 (N_6522,N_5898,N_4905);
nand U6523 (N_6523,N_4023,N_3345);
nand U6524 (N_6524,N_3451,N_3332);
nand U6525 (N_6525,N_3713,N_5129);
and U6526 (N_6526,N_3658,N_3971);
and U6527 (N_6527,N_4794,N_4493);
and U6528 (N_6528,N_3314,N_5578);
nand U6529 (N_6529,N_5983,N_3055);
nor U6530 (N_6530,N_5912,N_5203);
or U6531 (N_6531,N_5746,N_4327);
or U6532 (N_6532,N_4623,N_4474);
and U6533 (N_6533,N_5365,N_3088);
xor U6534 (N_6534,N_4900,N_4227);
and U6535 (N_6535,N_5183,N_5719);
nand U6536 (N_6536,N_3986,N_5580);
nand U6537 (N_6537,N_5541,N_3654);
or U6538 (N_6538,N_4765,N_5508);
or U6539 (N_6539,N_3430,N_3769);
and U6540 (N_6540,N_3236,N_4317);
nand U6541 (N_6541,N_5694,N_5363);
or U6542 (N_6542,N_5570,N_4665);
and U6543 (N_6543,N_5950,N_5342);
xor U6544 (N_6544,N_5028,N_3935);
nand U6545 (N_6545,N_3178,N_3275);
nand U6546 (N_6546,N_4858,N_4315);
and U6547 (N_6547,N_5426,N_3460);
nor U6548 (N_6548,N_3810,N_5633);
nor U6549 (N_6549,N_3167,N_5216);
nor U6550 (N_6550,N_5253,N_3123);
nor U6551 (N_6551,N_5531,N_5154);
or U6552 (N_6552,N_3139,N_3515);
or U6553 (N_6553,N_4853,N_4429);
and U6554 (N_6554,N_4751,N_4362);
nand U6555 (N_6555,N_3389,N_5285);
or U6556 (N_6556,N_3060,N_4875);
or U6557 (N_6557,N_3929,N_4021);
and U6558 (N_6558,N_3424,N_3698);
nand U6559 (N_6559,N_3714,N_5710);
nor U6560 (N_6560,N_5136,N_4446);
nand U6561 (N_6561,N_4644,N_4600);
nor U6562 (N_6562,N_5916,N_3909);
and U6563 (N_6563,N_5423,N_5862);
and U6564 (N_6564,N_5649,N_4374);
or U6565 (N_6565,N_5635,N_4116);
nand U6566 (N_6566,N_5582,N_3190);
and U6567 (N_6567,N_5468,N_3886);
nor U6568 (N_6568,N_5884,N_4974);
nand U6569 (N_6569,N_4015,N_5155);
nand U6570 (N_6570,N_5874,N_5352);
or U6571 (N_6571,N_3838,N_3462);
xor U6572 (N_6572,N_3371,N_5742);
or U6573 (N_6573,N_3756,N_4196);
or U6574 (N_6574,N_5383,N_3342);
or U6575 (N_6575,N_3686,N_5639);
or U6576 (N_6576,N_3665,N_4570);
nor U6577 (N_6577,N_4215,N_5000);
and U6578 (N_6578,N_4898,N_3495);
and U6579 (N_6579,N_3059,N_4811);
and U6580 (N_6580,N_3021,N_4430);
nand U6581 (N_6581,N_4046,N_3237);
or U6582 (N_6582,N_3078,N_3329);
nor U6583 (N_6583,N_4510,N_4447);
and U6584 (N_6584,N_3639,N_5229);
xnor U6585 (N_6585,N_5014,N_5838);
or U6586 (N_6586,N_4589,N_4105);
and U6587 (N_6587,N_5513,N_3353);
nor U6588 (N_6588,N_5795,N_4431);
nand U6589 (N_6589,N_3274,N_3307);
nand U6590 (N_6590,N_4223,N_5036);
nand U6591 (N_6591,N_3465,N_3807);
nor U6592 (N_6592,N_5738,N_4041);
or U6593 (N_6593,N_3053,N_4508);
xor U6594 (N_6594,N_3227,N_4761);
nand U6595 (N_6595,N_3951,N_5181);
or U6596 (N_6596,N_3948,N_5685);
nor U6597 (N_6597,N_4607,N_4203);
xnor U6598 (N_6598,N_4972,N_4096);
or U6599 (N_6599,N_3449,N_5975);
nand U6600 (N_6600,N_3404,N_5474);
and U6601 (N_6601,N_3045,N_5670);
or U6602 (N_6602,N_3141,N_5252);
nor U6603 (N_6603,N_4693,N_4284);
nand U6604 (N_6604,N_5230,N_5237);
or U6605 (N_6605,N_3938,N_4124);
xor U6606 (N_6606,N_3917,N_5684);
nor U6607 (N_6607,N_5382,N_4560);
and U6608 (N_6608,N_4631,N_5906);
and U6609 (N_6609,N_3379,N_4711);
or U6610 (N_6610,N_4542,N_4954);
nor U6611 (N_6611,N_3003,N_5515);
nor U6612 (N_6612,N_5214,N_4967);
nor U6613 (N_6613,N_5148,N_3041);
nor U6614 (N_6614,N_3696,N_4554);
xor U6615 (N_6615,N_4926,N_4184);
nand U6616 (N_6616,N_3626,N_4263);
and U6617 (N_6617,N_5678,N_4072);
or U6618 (N_6618,N_5586,N_4613);
and U6619 (N_6619,N_5057,N_5818);
or U6620 (N_6620,N_4376,N_3169);
nand U6621 (N_6621,N_3322,N_4042);
nor U6622 (N_6622,N_4068,N_5364);
or U6623 (N_6623,N_3004,N_3048);
nor U6624 (N_6624,N_3506,N_3912);
or U6625 (N_6625,N_5265,N_3820);
and U6626 (N_6626,N_3106,N_5652);
nand U6627 (N_6627,N_5837,N_3803);
and U6628 (N_6628,N_4084,N_3667);
nand U6629 (N_6629,N_5816,N_3801);
nand U6630 (N_6630,N_3047,N_5097);
or U6631 (N_6631,N_4528,N_3636);
nand U6632 (N_6632,N_3121,N_5740);
nor U6633 (N_6633,N_4459,N_5577);
xnor U6634 (N_6634,N_3615,N_5220);
and U6635 (N_6635,N_3730,N_5650);
nand U6636 (N_6636,N_3164,N_5343);
and U6637 (N_6637,N_3024,N_4849);
xor U6638 (N_6638,N_3577,N_3157);
and U6639 (N_6639,N_5996,N_5891);
nand U6640 (N_6640,N_5192,N_4424);
nor U6641 (N_6641,N_4808,N_5435);
nor U6642 (N_6642,N_4435,N_4438);
and U6643 (N_6643,N_4538,N_5132);
nand U6644 (N_6644,N_4047,N_5098);
nor U6645 (N_6645,N_4514,N_3459);
and U6646 (N_6646,N_4372,N_4365);
or U6647 (N_6647,N_3602,N_3815);
nand U6648 (N_6648,N_4498,N_3242);
and U6649 (N_6649,N_5866,N_3984);
or U6650 (N_6650,N_4170,N_4958);
nand U6651 (N_6651,N_4299,N_3857);
nand U6652 (N_6652,N_5278,N_3633);
and U6653 (N_6653,N_5895,N_5492);
nand U6654 (N_6654,N_3782,N_4942);
nand U6655 (N_6655,N_3688,N_3856);
and U6656 (N_6656,N_5479,N_5403);
nor U6657 (N_6657,N_5270,N_5256);
and U6658 (N_6658,N_4930,N_4256);
xor U6659 (N_6659,N_3964,N_3835);
nor U6660 (N_6660,N_4147,N_5574);
and U6661 (N_6661,N_3354,N_3130);
and U6662 (N_6662,N_5133,N_3681);
nor U6663 (N_6663,N_5461,N_4798);
or U6664 (N_6664,N_5357,N_3240);
and U6665 (N_6665,N_3095,N_4714);
nor U6666 (N_6666,N_5773,N_4448);
or U6667 (N_6667,N_4112,N_5280);
or U6668 (N_6668,N_5520,N_3025);
and U6669 (N_6669,N_5767,N_4163);
nor U6670 (N_6670,N_3327,N_4186);
or U6671 (N_6671,N_3922,N_3955);
or U6672 (N_6672,N_4143,N_3257);
xnor U6673 (N_6673,N_3438,N_3206);
or U6674 (N_6674,N_3170,N_5581);
nand U6675 (N_6675,N_4950,N_4371);
or U6676 (N_6676,N_3370,N_5959);
or U6677 (N_6677,N_4641,N_4035);
and U6678 (N_6678,N_3479,N_3818);
or U6679 (N_6679,N_5323,N_4799);
and U6680 (N_6680,N_4331,N_4829);
nand U6681 (N_6681,N_4216,N_4562);
nand U6682 (N_6682,N_5460,N_5019);
or U6683 (N_6683,N_5939,N_4011);
or U6684 (N_6684,N_5822,N_5638);
and U6685 (N_6685,N_5551,N_4436);
nand U6686 (N_6686,N_3301,N_3635);
and U6687 (N_6687,N_3421,N_4598);
and U6688 (N_6688,N_5478,N_3870);
xor U6689 (N_6689,N_5925,N_4990);
nor U6690 (N_6690,N_4896,N_5927);
nand U6691 (N_6691,N_4704,N_4935);
and U6692 (N_6692,N_5557,N_3194);
nor U6693 (N_6693,N_3432,N_3819);
nor U6694 (N_6694,N_4479,N_5034);
nor U6695 (N_6695,N_3764,N_4118);
or U6696 (N_6696,N_4356,N_3881);
or U6697 (N_6697,N_5109,N_5505);
or U6698 (N_6698,N_5398,N_5976);
and U6699 (N_6699,N_5384,N_5576);
nor U6700 (N_6700,N_3397,N_3554);
and U6701 (N_6701,N_4812,N_4738);
and U6702 (N_6702,N_5908,N_3077);
nor U6703 (N_6703,N_5454,N_4164);
nor U6704 (N_6704,N_4366,N_4158);
and U6705 (N_6705,N_4242,N_5698);
and U6706 (N_6706,N_3100,N_4899);
nor U6707 (N_6707,N_3627,N_4823);
xor U6708 (N_6708,N_4031,N_4871);
nor U6709 (N_6709,N_5727,N_5663);
and U6710 (N_6710,N_3230,N_5065);
nor U6711 (N_6711,N_3184,N_4101);
nor U6712 (N_6712,N_3336,N_4344);
or U6713 (N_6713,N_5318,N_4724);
nand U6714 (N_6714,N_5396,N_5903);
nand U6715 (N_6715,N_4130,N_4807);
nor U6716 (N_6716,N_5716,N_5887);
xor U6717 (N_6717,N_5986,N_5327);
nand U6718 (N_6718,N_3195,N_5902);
nor U6719 (N_6719,N_3594,N_4970);
or U6720 (N_6720,N_4686,N_3213);
nor U6721 (N_6721,N_4207,N_4874);
nor U6722 (N_6722,N_3054,N_3014);
or U6723 (N_6723,N_4938,N_3579);
nor U6724 (N_6724,N_3118,N_4355);
nor U6725 (N_6725,N_5257,N_4913);
and U6726 (N_6726,N_5946,N_4546);
nand U6727 (N_6727,N_3488,N_4411);
nand U6728 (N_6728,N_5119,N_5068);
and U6729 (N_6729,N_4302,N_4395);
and U6730 (N_6730,N_3359,N_3923);
or U6731 (N_6731,N_4150,N_4890);
and U6732 (N_6732,N_4567,N_4661);
xnor U6733 (N_6733,N_4998,N_3291);
xnor U6734 (N_6734,N_3916,N_5314);
nor U6735 (N_6735,N_5629,N_4564);
or U6736 (N_6736,N_3933,N_3584);
and U6737 (N_6737,N_4940,N_5564);
nand U6738 (N_6738,N_3433,N_3563);
nand U6739 (N_6739,N_5377,N_5143);
and U6740 (N_6740,N_4404,N_4833);
nand U6741 (N_6741,N_5932,N_5297);
nand U6742 (N_6742,N_5808,N_5063);
or U6743 (N_6743,N_5149,N_4809);
xor U6744 (N_6744,N_3517,N_5496);
nand U6745 (N_6745,N_4503,N_3915);
or U6746 (N_6746,N_5717,N_5592);
nand U6747 (N_6747,N_4959,N_5995);
and U6748 (N_6748,N_3094,N_5931);
and U6749 (N_6749,N_4687,N_4148);
and U6750 (N_6750,N_4922,N_4586);
xnor U6751 (N_6751,N_5894,N_4670);
or U6752 (N_6752,N_3463,N_3907);
and U6753 (N_6753,N_4790,N_5978);
nor U6754 (N_6754,N_3892,N_5249);
nand U6755 (N_6755,N_4036,N_5980);
xor U6756 (N_6756,N_3012,N_3772);
nand U6757 (N_6757,N_5759,N_3253);
or U6758 (N_6758,N_3830,N_3573);
xnor U6759 (N_6759,N_3895,N_3200);
nand U6760 (N_6760,N_3703,N_3313);
nor U6761 (N_6761,N_3880,N_5548);
nand U6762 (N_6762,N_4831,N_5796);
and U6763 (N_6763,N_3205,N_5107);
and U6764 (N_6764,N_4014,N_3443);
and U6765 (N_6765,N_5163,N_5374);
nor U6766 (N_6766,N_3548,N_5347);
nand U6767 (N_6767,N_3511,N_3617);
and U6768 (N_6768,N_3392,N_4174);
xnor U6769 (N_6769,N_3987,N_4065);
nand U6770 (N_6770,N_4880,N_4642);
and U6771 (N_6771,N_3160,N_5083);
nand U6772 (N_6772,N_5484,N_5849);
and U6773 (N_6773,N_3634,N_4360);
nor U6774 (N_6774,N_3180,N_5187);
or U6775 (N_6775,N_4434,N_5854);
nor U6776 (N_6776,N_4238,N_4316);
and U6777 (N_6777,N_3223,N_5624);
nand U6778 (N_6778,N_4168,N_4060);
and U6779 (N_6779,N_5501,N_3578);
nand U6780 (N_6780,N_4533,N_3748);
nand U6781 (N_6781,N_4868,N_3050);
nor U6782 (N_6782,N_5543,N_5695);
nand U6783 (N_6783,N_4556,N_4962);
nor U6784 (N_6784,N_4291,N_4156);
xor U6785 (N_6785,N_4121,N_5715);
and U6786 (N_6786,N_3201,N_4300);
nand U6787 (N_6787,N_3522,N_5387);
or U6788 (N_6788,N_3771,N_5224);
or U6789 (N_6789,N_4936,N_4246);
nor U6790 (N_6790,N_5462,N_3192);
nor U6791 (N_6791,N_3662,N_3181);
or U6792 (N_6792,N_3585,N_5114);
nor U6793 (N_6793,N_5779,N_4437);
nor U6794 (N_6794,N_4932,N_3685);
and U6795 (N_6795,N_4454,N_3061);
xor U6796 (N_6796,N_4877,N_3493);
nor U6797 (N_6797,N_4695,N_4301);
nor U6798 (N_6798,N_4772,N_3972);
and U6799 (N_6799,N_5647,N_4233);
nor U6800 (N_6800,N_4480,N_4963);
xnor U6801 (N_6801,N_4723,N_5599);
nor U6802 (N_6802,N_3668,N_5010);
nor U6803 (N_6803,N_3564,N_3540);
and U6804 (N_6804,N_3677,N_4171);
or U6805 (N_6805,N_4428,N_3367);
nand U6806 (N_6806,N_5100,N_3395);
nand U6807 (N_6807,N_3022,N_5212);
and U6808 (N_6808,N_3507,N_5117);
or U6809 (N_6809,N_4574,N_5553);
xnor U6810 (N_6810,N_5244,N_4947);
and U6811 (N_6811,N_5296,N_3442);
nor U6812 (N_6812,N_4460,N_5215);
or U6813 (N_6813,N_5744,N_3016);
xnor U6814 (N_6814,N_4097,N_3420);
nor U6815 (N_6815,N_4523,N_3193);
nor U6816 (N_6816,N_5142,N_4298);
and U6817 (N_6817,N_5041,N_3978);
nor U6818 (N_6818,N_5703,N_3305);
and U6819 (N_6819,N_3709,N_4471);
nor U6820 (N_6820,N_5506,N_5087);
nand U6821 (N_6821,N_4009,N_3559);
or U6822 (N_6822,N_3102,N_5799);
or U6823 (N_6823,N_4845,N_5276);
or U6824 (N_6824,N_3009,N_5778);
nor U6825 (N_6825,N_3241,N_3429);
and U6826 (N_6826,N_3569,N_3104);
and U6827 (N_6827,N_3779,N_4988);
xnor U6828 (N_6828,N_3614,N_4076);
or U6829 (N_6829,N_3776,N_3560);
nand U6830 (N_6830,N_3210,N_4787);
nand U6831 (N_6831,N_4634,N_4264);
xor U6832 (N_6832,N_5081,N_5335);
xnor U6833 (N_6833,N_3467,N_4740);
nor U6834 (N_6834,N_4099,N_5186);
nor U6835 (N_6835,N_5137,N_3754);
nand U6836 (N_6836,N_5211,N_5567);
nor U6837 (N_6837,N_4842,N_4018);
and U6838 (N_6838,N_3931,N_3413);
nor U6839 (N_6839,N_3234,N_3530);
and U6840 (N_6840,N_3557,N_4310);
or U6841 (N_6841,N_3196,N_5828);
xnor U6842 (N_6842,N_4544,N_5466);
xor U6843 (N_6843,N_3005,N_5720);
xor U6844 (N_6844,N_3425,N_5954);
or U6845 (N_6845,N_5354,N_5414);
and U6846 (N_6846,N_5876,N_5645);
nor U6847 (N_6847,N_5693,N_3792);
and U6848 (N_6848,N_3704,N_5984);
and U6849 (N_6849,N_4805,N_3650);
nor U6850 (N_6850,N_4225,N_5258);
nor U6851 (N_6851,N_4006,N_4863);
or U6852 (N_6852,N_5105,N_5222);
nand U6853 (N_6853,N_4108,N_4119);
or U6854 (N_6854,N_4891,N_4700);
and U6855 (N_6855,N_4172,N_4452);
xor U6856 (N_6856,N_3596,N_3566);
nor U6857 (N_6857,N_5845,N_3186);
nand U6858 (N_6858,N_5091,N_3376);
nand U6859 (N_6859,N_4417,N_5371);
nand U6860 (N_6860,N_3683,N_5362);
or U6861 (N_6861,N_5937,N_4852);
nand U6862 (N_6862,N_5096,N_4762);
or U6863 (N_6863,N_4717,N_4187);
nand U6864 (N_6864,N_5381,N_5733);
or U6865 (N_6865,N_4442,N_5072);
nand U6866 (N_6866,N_5023,N_3013);
nand U6867 (N_6867,N_5538,N_4177);
nor U6868 (N_6868,N_3994,N_4039);
nand U6869 (N_6869,N_5798,N_3197);
nor U6870 (N_6870,N_3965,N_5943);
xor U6871 (N_6871,N_5536,N_4137);
and U6872 (N_6872,N_3386,N_4786);
xnor U6873 (N_6873,N_3651,N_4294);
and U6874 (N_6874,N_5070,N_3629);
nand U6875 (N_6875,N_5473,N_3612);
xnor U6876 (N_6876,N_5713,N_5871);
or U6877 (N_6877,N_3255,N_5615);
or U6878 (N_6878,N_3786,N_4753);
nor U6879 (N_6879,N_3142,N_5272);
nand U6880 (N_6880,N_4359,N_3456);
or U6881 (N_6881,N_5533,N_3534);
nor U6882 (N_6882,N_4075,N_4024);
nand U6883 (N_6883,N_3538,N_4304);
or U6884 (N_6884,N_4334,N_5765);
or U6885 (N_6885,N_5657,N_3028);
nand U6886 (N_6886,N_3903,N_5162);
or U6887 (N_6887,N_3785,N_4463);
nor U6888 (N_6888,N_4781,N_3832);
nand U6889 (N_6889,N_5411,N_3218);
and U6890 (N_6890,N_3828,N_4836);
nor U6891 (N_6891,N_4385,N_4004);
and U6892 (N_6892,N_4691,N_5709);
and U6893 (N_6893,N_4629,N_4591);
or U6894 (N_6894,N_5011,N_4991);
and U6895 (N_6895,N_5770,N_3732);
nand U6896 (N_6896,N_3120,N_3927);
and U6897 (N_6897,N_5668,N_3026);
nor U6898 (N_6898,N_5499,N_5282);
or U6899 (N_6899,N_3648,N_5622);
xor U6900 (N_6900,N_4013,N_3018);
xnor U6901 (N_6901,N_4943,N_4934);
and U6902 (N_6902,N_3834,N_5455);
xor U6903 (N_6903,N_5144,N_5053);
nand U6904 (N_6904,N_4211,N_4293);
and U6905 (N_6905,N_3884,N_5217);
and U6906 (N_6906,N_4981,N_4353);
or U6907 (N_6907,N_4973,N_3720);
nor U6908 (N_6908,N_4329,N_5438);
and U6909 (N_6909,N_4102,N_3599);
nor U6910 (N_6910,N_5123,N_5498);
or U6911 (N_6911,N_3374,N_3093);
or U6912 (N_6912,N_3958,N_3660);
or U6913 (N_6913,N_4697,N_3543);
nand U6914 (N_6914,N_3066,N_3670);
nand U6915 (N_6915,N_3148,N_5184);
and U6916 (N_6916,N_3105,N_5090);
xor U6917 (N_6917,N_5389,N_5131);
or U6918 (N_6918,N_5608,N_3069);
or U6919 (N_6919,N_3657,N_4791);
and U6920 (N_6920,N_5275,N_5050);
nor U6921 (N_6921,N_3089,N_5400);
nor U6922 (N_6922,N_3073,N_5127);
and U6923 (N_6923,N_5514,N_4303);
nand U6924 (N_6924,N_4706,N_5027);
nor U6925 (N_6925,N_3410,N_3859);
and U6926 (N_6926,N_4455,N_3243);
nand U6927 (N_6927,N_5089,N_4179);
nor U6928 (N_6928,N_4531,N_3589);
or U6929 (N_6929,N_4142,N_5052);
and U6930 (N_6930,N_4526,N_3290);
and U6931 (N_6931,N_5547,N_5341);
or U6932 (N_6932,N_5554,N_4134);
or U6933 (N_6933,N_4667,N_5883);
and U6934 (N_6934,N_3780,N_4593);
nor U6935 (N_6935,N_3477,N_3229);
and U6936 (N_6936,N_3039,N_5355);
or U6937 (N_6937,N_4577,N_4349);
xnor U6938 (N_6938,N_4194,N_5467);
and U6939 (N_6939,N_4841,N_3908);
nor U6940 (N_6940,N_5511,N_5124);
nand U6941 (N_6941,N_5690,N_3899);
nand U6942 (N_6942,N_5429,N_4421);
or U6943 (N_6943,N_3684,N_4477);
and U6944 (N_6944,N_5268,N_5783);
nand U6945 (N_6945,N_5021,N_5095);
or U6946 (N_6946,N_5896,N_5552);
nor U6947 (N_6947,N_4835,N_3323);
nor U6948 (N_6948,N_5936,N_5823);
nand U6949 (N_6949,N_5839,N_4688);
or U6950 (N_6950,N_5385,N_5228);
nand U6951 (N_6951,N_3647,N_3215);
or U6952 (N_6952,N_4161,N_4690);
or U6953 (N_6953,N_4729,N_5266);
or U6954 (N_6954,N_3528,N_3624);
and U6955 (N_6955,N_5841,N_4756);
nand U6956 (N_6956,N_4351,N_4846);
nand U6957 (N_6957,N_3546,N_3226);
and U6958 (N_6958,N_3212,N_5760);
nand U6959 (N_6959,N_4026,N_4949);
or U6960 (N_6960,N_5872,N_3179);
nand U6961 (N_6961,N_5739,N_5421);
and U6962 (N_6962,N_4617,N_5487);
and U6963 (N_6963,N_4626,N_5235);
and U6964 (N_6964,N_5982,N_4886);
xnor U6965 (N_6965,N_5178,N_5625);
nor U6966 (N_6966,N_5195,N_5804);
nor U6967 (N_6967,N_4090,N_4067);
or U6968 (N_6968,N_4131,N_3002);
or U6969 (N_6969,N_4602,N_5985);
or U6970 (N_6970,N_4093,N_4037);
nor U6971 (N_6971,N_4948,N_3711);
and U6972 (N_6972,N_3854,N_4336);
and U6973 (N_6973,N_4029,N_5594);
nand U6974 (N_6974,N_4746,N_5378);
xor U6975 (N_6975,N_5509,N_3718);
xor U6976 (N_6976,N_4132,N_4370);
or U6977 (N_6977,N_5677,N_3678);
nand U6978 (N_6978,N_3019,N_5968);
nor U6979 (N_6979,N_3324,N_3572);
nor U6980 (N_6980,N_5177,N_4020);
or U6981 (N_6981,N_5970,N_4792);
nor U6982 (N_6982,N_3387,N_5526);
nand U6983 (N_6983,N_4354,N_5532);
nand U6984 (N_6984,N_4113,N_4754);
nor U6985 (N_6985,N_3422,N_5407);
nand U6986 (N_6986,N_3468,N_4425);
and U6987 (N_6987,N_3356,N_3202);
xnor U6988 (N_6988,N_3081,N_3516);
nor U6989 (N_6989,N_3645,N_3841);
nor U6990 (N_6990,N_5045,N_5627);
or U6991 (N_6991,N_5436,N_4400);
nand U6992 (N_6992,N_4603,N_5504);
xnor U6993 (N_6993,N_3117,N_4377);
or U6994 (N_6994,N_3977,N_5998);
xnor U6995 (N_6995,N_4275,N_3068);
or U6996 (N_6996,N_5786,N_3366);
nand U6997 (N_6997,N_4664,N_5987);
and U6998 (N_6998,N_4920,N_4157);
xnor U6999 (N_6999,N_5613,N_5723);
nor U7000 (N_7000,N_5558,N_5390);
nor U7001 (N_7001,N_4648,N_4671);
and U7002 (N_7002,N_4251,N_4847);
nor U7003 (N_7003,N_5026,N_3076);
or U7004 (N_7004,N_3071,N_4169);
or U7005 (N_7005,N_3476,N_5415);
nor U7006 (N_7006,N_4333,N_3116);
and U7007 (N_7007,N_4472,N_4737);
nor U7008 (N_7008,N_4573,N_3993);
nor U7009 (N_7009,N_4205,N_3035);
nor U7010 (N_7010,N_5321,N_4311);
or U7011 (N_7011,N_4027,N_3632);
nand U7012 (N_7012,N_3222,N_3934);
nand U7013 (N_7013,N_4635,N_4394);
xnor U7014 (N_7014,N_5289,N_4653);
nand U7015 (N_7015,N_3891,N_4904);
or U7016 (N_7016,N_3567,N_3135);
and U7017 (N_7017,N_5595,N_5472);
or U7018 (N_7018,N_5465,N_3555);
nand U7019 (N_7019,N_3736,N_4744);
xnor U7020 (N_7020,N_4535,N_3882);
or U7021 (N_7021,N_5785,N_5921);
xnor U7022 (N_7022,N_3383,N_4747);
nor U7023 (N_7023,N_4743,N_4221);
or U7024 (N_7024,N_3842,N_3246);
nand U7025 (N_7025,N_4927,N_5598);
and U7026 (N_7026,N_4159,N_4338);
and U7027 (N_7027,N_3423,N_5761);
nor U7028 (N_7028,N_3896,N_3911);
nand U7029 (N_7029,N_3062,N_3941);
xnor U7030 (N_7030,N_3752,N_3822);
nor U7031 (N_7031,N_3587,N_4685);
and U7032 (N_7032,N_5907,N_5753);
nand U7033 (N_7033,N_3110,N_4450);
nand U7034 (N_7034,N_3015,N_3944);
nor U7035 (N_7035,N_3705,N_5529);
nor U7036 (N_7036,N_3214,N_4109);
and U7037 (N_7037,N_4082,N_3150);
or U7038 (N_7038,N_4989,N_4820);
nor U7039 (N_7039,N_5223,N_4348);
or U7040 (N_7040,N_3597,N_3778);
or U7041 (N_7041,N_3125,N_3521);
xnor U7042 (N_7042,N_4669,N_5439);
or U7043 (N_7043,N_4692,N_4497);
nor U7044 (N_7044,N_3902,N_5591);
xnor U7045 (N_7045,N_5422,N_3268);
xor U7046 (N_7046,N_5290,N_3789);
nand U7047 (N_7047,N_4346,N_4997);
and U7048 (N_7048,N_3352,N_5748);
nand U7049 (N_7049,N_3840,N_3655);
and U7050 (N_7050,N_3618,N_4624);
or U7051 (N_7051,N_4237,N_5093);
nand U7052 (N_7052,N_3440,N_5924);
nor U7053 (N_7053,N_5300,N_4133);
or U7054 (N_7054,N_3485,N_5671);
nand U7055 (N_7055,N_3524,N_5794);
or U7056 (N_7056,N_3956,N_3952);
and U7057 (N_7057,N_3689,N_3622);
or U7058 (N_7058,N_3630,N_3999);
and U7059 (N_7059,N_4202,N_3315);
nor U7060 (N_7060,N_4476,N_4262);
nand U7061 (N_7061,N_3700,N_5527);
or U7062 (N_7062,N_4361,N_3097);
nand U7063 (N_7063,N_5205,N_4590);
or U7064 (N_7064,N_3153,N_3601);
nor U7065 (N_7065,N_4254,N_4917);
nand U7066 (N_7066,N_4699,N_3727);
nor U7067 (N_7067,N_3096,N_5612);
xor U7068 (N_7068,N_5231,N_3508);
nor U7069 (N_7069,N_3435,N_4441);
xnor U7070 (N_7070,N_3746,N_4261);
nand U7071 (N_7071,N_5636,N_5168);
and U7072 (N_7072,N_4881,N_4136);
nor U7073 (N_7073,N_3399,N_4878);
and U7074 (N_7074,N_3360,N_5145);
nand U7075 (N_7075,N_4908,N_3745);
nand U7076 (N_7076,N_5571,N_4885);
and U7077 (N_7077,N_4592,N_3706);
nand U7078 (N_7078,N_5732,N_5792);
nand U7079 (N_7079,N_4797,N_5164);
and U7080 (N_7080,N_3831,N_4063);
or U7081 (N_7081,N_4005,N_3284);
nor U7082 (N_7082,N_4017,N_3805);
nor U7083 (N_7083,N_5674,N_5658);
xnor U7084 (N_7084,N_5632,N_3441);
and U7085 (N_7085,N_3939,N_3017);
and U7086 (N_7086,N_4576,N_3898);
or U7087 (N_7087,N_4719,N_4139);
nand U7088 (N_7088,N_3119,N_4978);
and U7089 (N_7089,N_3209,N_3310);
and U7090 (N_7090,N_3346,N_4022);
nand U7091 (N_7091,N_5022,N_3541);
and U7092 (N_7092,N_5814,N_4280);
xor U7093 (N_7093,N_5958,N_3337);
and U7094 (N_7094,N_4066,N_4909);
nor U7095 (N_7095,N_5977,N_4104);
and U7096 (N_7096,N_5616,N_4193);
nand U7097 (N_7097,N_3788,N_4912);
nor U7098 (N_7098,N_4696,N_3850);
nor U7099 (N_7099,N_3149,N_3333);
and U7100 (N_7100,N_4324,N_4595);
or U7101 (N_7101,N_5810,N_5402);
nand U7102 (N_7102,N_5281,N_4712);
or U7103 (N_7103,N_3809,N_3949);
and U7104 (N_7104,N_5540,N_4843);
or U7105 (N_7105,N_3107,N_4894);
nand U7106 (N_7106,N_4563,N_5078);
and U7107 (N_7107,N_5248,N_5923);
or U7108 (N_7108,N_3860,N_5444);
or U7109 (N_7109,N_5437,N_5491);
nor U7110 (N_7110,N_3162,N_5692);
and U7111 (N_7111,N_5856,N_4115);
nand U7112 (N_7112,N_4181,N_5388);
and U7113 (N_7113,N_3795,N_3406);
or U7114 (N_7114,N_5961,N_4410);
or U7115 (N_7115,N_3133,N_3652);
nor U7116 (N_7116,N_5754,N_3814);
xnor U7117 (N_7117,N_4218,N_5620);
nand U7118 (N_7118,N_5780,N_5126);
and U7119 (N_7119,N_5766,N_5325);
xor U7120 (N_7120,N_3812,N_4412);
or U7121 (N_7121,N_4530,N_4971);
or U7122 (N_7122,N_5546,N_5234);
nand U7123 (N_7123,N_3740,N_3871);
or U7124 (N_7124,N_3608,N_5762);
nor U7125 (N_7125,N_3027,N_3478);
xnor U7126 (N_7126,N_3995,N_4509);
xor U7127 (N_7127,N_5048,N_5882);
and U7128 (N_7128,N_4318,N_5777);
or U7129 (N_7129,N_5405,N_3364);
and U7130 (N_7130,N_4636,N_3733);
nand U7131 (N_7131,N_4313,N_5519);
or U7132 (N_7132,N_5626,N_5273);
nor U7133 (N_7133,N_5990,N_4239);
nor U7134 (N_7134,N_5076,N_4295);
or U7135 (N_7135,N_3319,N_5470);
nor U7136 (N_7136,N_3997,N_3724);
nor U7137 (N_7137,N_5784,N_3341);
and U7138 (N_7138,N_3266,N_4505);
nand U7139 (N_7139,N_5350,N_3168);
and U7140 (N_7140,N_4543,N_5348);
nor U7141 (N_7141,N_3890,N_4580);
nor U7142 (N_7142,N_5601,N_5702);
and U7143 (N_7143,N_4583,N_4599);
nand U7144 (N_7144,N_4750,N_5630);
xnor U7145 (N_7145,N_3960,N_4784);
nor U7146 (N_7146,N_3529,N_3565);
and U7147 (N_7147,N_4226,N_5914);
nor U7148 (N_7148,N_5609,N_4848);
nand U7149 (N_7149,N_5225,N_4117);
or U7150 (N_7150,N_5830,N_3475);
or U7151 (N_7151,N_4965,N_5295);
nand U7152 (N_7152,N_4384,N_3583);
and U7153 (N_7153,N_4561,N_5945);
nor U7154 (N_7154,N_5824,N_4897);
nand U7155 (N_7155,N_3361,N_5156);
xor U7156 (N_7156,N_4232,N_4427);
nand U7157 (N_7157,N_5942,N_5992);
or U7158 (N_7158,N_5974,N_4774);
and U7159 (N_7159,N_4475,N_3405);
and U7160 (N_7160,N_4707,N_4451);
and U7161 (N_7161,N_4608,N_4403);
or U7162 (N_7162,N_4515,N_3221);
nand U7163 (N_7163,N_4255,N_3282);
nand U7164 (N_7164,N_3766,N_3790);
nand U7165 (N_7165,N_4715,N_3590);
nand U7166 (N_7166,N_4861,N_4107);
nand U7167 (N_7167,N_3481,N_4214);
and U7168 (N_7168,N_3513,N_5316);
nor U7169 (N_7169,N_3042,N_4034);
and U7170 (N_7170,N_3052,N_5441);
nor U7171 (N_7171,N_5147,N_5569);
or U7172 (N_7172,N_4129,N_4189);
and U7173 (N_7173,N_3051,N_4705);
nand U7174 (N_7174,N_3768,N_4518);
nor U7175 (N_7175,N_4964,N_4735);
nand U7176 (N_7176,N_5193,N_5394);
xnor U7177 (N_7177,N_4957,N_3330);
and U7178 (N_7178,N_4058,N_3701);
nand U7179 (N_7179,N_5064,N_5161);
nor U7180 (N_7180,N_3797,N_4680);
nand U7181 (N_7181,N_5602,N_4198);
nor U7182 (N_7182,N_3878,N_3953);
nor U7183 (N_7183,N_4341,N_5725);
and U7184 (N_7184,N_3586,N_4210);
nor U7185 (N_7185,N_4381,N_3598);
or U7186 (N_7186,N_4248,N_4405);
nand U7187 (N_7187,N_5030,N_3176);
and U7188 (N_7188,N_4453,N_4710);
and U7189 (N_7189,N_3742,N_3723);
nand U7190 (N_7190,N_5025,N_3235);
and U7191 (N_7191,N_4231,N_5687);
xnor U7192 (N_7192,N_3519,N_4645);
or U7193 (N_7193,N_5763,N_4487);
and U7194 (N_7194,N_3384,N_5660);
xnor U7195 (N_7195,N_5889,N_4369);
or U7196 (N_7196,N_4650,N_5523);
or U7197 (N_7197,N_3338,N_3103);
or U7198 (N_7198,N_3523,N_3692);
nor U7199 (N_7199,N_3982,N_4733);
nand U7200 (N_7200,N_3046,N_3739);
or U7201 (N_7201,N_4923,N_5556);
and U7202 (N_7202,N_3251,N_5749);
xor U7203 (N_7203,N_4673,N_5637);
or U7204 (N_7204,N_4911,N_5226);
or U7205 (N_7205,N_3817,N_4491);
nor U7206 (N_7206,N_3185,N_5447);
nand U7207 (N_7207,N_3755,N_5701);
nor U7208 (N_7208,N_5813,N_3113);
nand U7209 (N_7209,N_3265,N_4305);
xor U7210 (N_7210,N_3156,N_3775);
nand U7211 (N_7211,N_3767,N_4464);
or U7212 (N_7212,N_5094,N_5619);
xor U7213 (N_7213,N_4953,N_4473);
and U7214 (N_7214,N_4440,N_5138);
nor U7215 (N_7215,N_4145,N_4496);
xor U7216 (N_7216,N_5442,N_4764);
nand U7217 (N_7217,N_5755,N_3283);
and U7218 (N_7218,N_4390,N_4540);
nor U7219 (N_7219,N_4867,N_3717);
xnor U7220 (N_7220,N_4321,N_3248);
and U7221 (N_7221,N_5913,N_3687);
or U7222 (N_7222,N_3312,N_5369);
nor U7223 (N_7223,N_5293,N_4154);
nand U7224 (N_7224,N_3762,N_3637);
or U7225 (N_7225,N_4388,N_5628);
and U7226 (N_7226,N_5151,N_3258);
nor U7227 (N_7227,N_5641,N_3826);
xnor U7228 (N_7228,N_5899,N_4008);
nand U7229 (N_7229,N_3377,N_3715);
or U7230 (N_7230,N_5944,N_4918);
nor U7231 (N_7231,N_4373,N_5651);
nor U7232 (N_7232,N_3619,N_5847);
nor U7233 (N_7233,N_3751,N_5964);
and U7234 (N_7234,N_5672,N_3674);
or U7235 (N_7235,N_5610,N_4547);
nor U7236 (N_7236,N_5865,N_3188);
and U7237 (N_7237,N_4319,N_5962);
nor U7238 (N_7238,N_4941,N_3514);
nand U7239 (N_7239,N_3444,N_3159);
and U7240 (N_7240,N_3001,N_3998);
xor U7241 (N_7241,N_3861,N_3286);
or U7242 (N_7242,N_5054,N_5035);
xor U7243 (N_7243,N_3979,N_3843);
nor U7244 (N_7244,N_3132,N_4668);
nor U7245 (N_7245,N_5336,N_5604);
nor U7246 (N_7246,N_3204,N_4814);
or U7247 (N_7247,N_5960,N_4982);
nor U7248 (N_7248,N_4616,N_4928);
or U7249 (N_7249,N_5379,N_5897);
or U7250 (N_7250,N_5801,N_3318);
nor U7251 (N_7251,N_3855,N_4195);
nand U7252 (N_7252,N_3357,N_5313);
nor U7253 (N_7253,N_4924,N_3326);
and U7254 (N_7254,N_5317,N_5575);
and U7255 (N_7255,N_3574,N_4085);
and U7256 (N_7256,N_3224,N_5092);
nand U7257 (N_7257,N_3427,N_5077);
and U7258 (N_7258,N_4581,N_5718);
nor U7259 (N_7259,N_5440,N_3031);
and U7260 (N_7260,N_5679,N_3663);
nand U7261 (N_7261,N_4288,N_5989);
or U7262 (N_7262,N_5476,N_5221);
nor U7263 (N_7263,N_5929,N_5331);
nand U7264 (N_7264,N_5418,N_3457);
xor U7265 (N_7265,N_5084,N_3532);
or U7266 (N_7266,N_3348,N_3913);
or U7267 (N_7267,N_3147,N_3510);
xnor U7268 (N_7268,N_4643,N_5704);
nor U7269 (N_7269,N_3007,N_4578);
nor U7270 (N_7270,N_3109,N_3562);
nand U7271 (N_7271,N_5279,N_5116);
nor U7272 (N_7272,N_5539,N_3777);
and U7273 (N_7273,N_4418,N_5667);
nor U7274 (N_7274,N_4506,N_4269);
and U7275 (N_7275,N_4220,N_4146);
and U7276 (N_7276,N_4467,N_3571);
and U7277 (N_7277,N_4779,N_3183);
and U7278 (N_7278,N_3509,N_4088);
xnor U7279 (N_7279,N_3996,N_4155);
and U7280 (N_7280,N_3862,N_5328);
nor U7281 (N_7281,N_3969,N_3537);
nor U7282 (N_7282,N_3358,N_5413);
and U7283 (N_7283,N_5012,N_5038);
nor U7284 (N_7284,N_4249,N_4870);
or U7285 (N_7285,N_5032,N_5376);
nand U7286 (N_7286,N_5056,N_4976);
nand U7287 (N_7287,N_4789,N_3091);
or U7288 (N_7288,N_5016,N_4655);
or U7289 (N_7289,N_3784,N_4937);
xor U7290 (N_7290,N_4666,N_5691);
nand U7291 (N_7291,N_4682,N_4745);
or U7292 (N_7292,N_4606,N_5851);
nand U7293 (N_7293,N_5673,N_5366);
nor U7294 (N_7294,N_3580,N_5428);
nand U7295 (N_7295,N_3631,N_5283);
or U7296 (N_7296,N_3887,N_4778);
nand U7297 (N_7297,N_3520,N_3403);
or U7298 (N_7298,N_4625,N_3043);
nand U7299 (N_7299,N_3075,N_5644);
and U7300 (N_7300,N_4213,N_3581);
nand U7301 (N_7301,N_3974,N_5425);
and U7302 (N_7302,N_5825,N_5419);
or U7303 (N_7303,N_4929,N_5344);
nor U7304 (N_7304,N_4663,N_5392);
xor U7305 (N_7305,N_5261,N_3385);
or U7306 (N_7306,N_4541,N_3434);
or U7307 (N_7307,N_4352,N_5262);
or U7308 (N_7308,N_5274,N_3272);
or U7309 (N_7309,N_5326,N_4681);
or U7310 (N_7310,N_3989,N_4916);
nor U7311 (N_7311,N_4550,N_4866);
nand U7312 (N_7312,N_4485,N_5708);
nand U7313 (N_7313,N_4032,N_5208);
or U7314 (N_7314,N_4638,N_5955);
nor U7315 (N_7315,N_5139,N_5269);
or U7316 (N_7316,N_4810,N_4297);
xor U7317 (N_7317,N_3849,N_5852);
nand U7318 (N_7318,N_4933,N_4423);
nor U7319 (N_7319,N_4758,N_5700);
or U7320 (N_7320,N_4628,N_3774);
nor U7321 (N_7321,N_3390,N_5080);
nand U7322 (N_7322,N_4621,N_4287);
nor U7323 (N_7323,N_4939,N_4701);
nor U7324 (N_7324,N_5901,N_3339);
xnor U7325 (N_7325,N_5642,N_4462);
or U7326 (N_7326,N_5236,N_5930);
nand U7327 (N_7327,N_3800,N_5797);
or U7328 (N_7328,N_3058,N_5669);
nor U7329 (N_7329,N_3302,N_4865);
and U7330 (N_7330,N_5448,N_5517);
nand U7331 (N_7331,N_5655,N_4815);
nand U7332 (N_7332,N_5227,N_3525);
and U7333 (N_7333,N_4499,N_5605);
or U7334 (N_7334,N_4180,N_4342);
or U7335 (N_7335,N_4083,N_4565);
or U7336 (N_7336,N_3320,N_4995);
nor U7337 (N_7337,N_4532,N_3640);
nand U7338 (N_7338,N_5661,N_5648);
nand U7339 (N_7339,N_3128,N_4357);
or U7340 (N_7340,N_5507,N_5412);
nor U7341 (N_7341,N_5560,N_5634);
nor U7342 (N_7342,N_5614,N_3787);
nor U7343 (N_7343,N_3975,N_4804);
nand U7344 (N_7344,N_3298,N_3114);
nand U7345 (N_7345,N_4637,N_5319);
nand U7346 (N_7346,N_5806,N_4749);
or U7347 (N_7347,N_4571,N_3502);
xnor U7348 (N_7348,N_3866,N_3144);
or U7349 (N_7349,N_3278,N_4456);
or U7350 (N_7350,N_4204,N_5334);
nor U7351 (N_7351,N_4257,N_5940);
nand U7352 (N_7352,N_5682,N_3848);
or U7353 (N_7353,N_5953,N_4766);
xnor U7354 (N_7354,N_5058,N_4622);
nor U7355 (N_7355,N_4689,N_5079);
nor U7356 (N_7356,N_4235,N_4979);
and U7357 (N_7357,N_4069,N_5255);
nand U7358 (N_7358,N_3267,N_4821);
nor U7359 (N_7359,N_4469,N_4490);
or U7360 (N_7360,N_3735,N_5434);
nand U7361 (N_7361,N_4525,N_4620);
and U7362 (N_7362,N_5829,N_5247);
nand U7363 (N_7363,N_5004,N_5597);
or U7364 (N_7364,N_3770,N_5310);
nor U7365 (N_7365,N_4656,N_5104);
nor U7366 (N_7366,N_4244,N_4488);
or U7367 (N_7367,N_4558,N_3694);
nor U7368 (N_7368,N_3285,N_5750);
and U7369 (N_7369,N_4458,N_5805);
and U7370 (N_7370,N_4413,N_5303);
xnor U7371 (N_7371,N_3722,N_4457);
nand U7372 (N_7372,N_4126,N_4775);
nor U7373 (N_7373,N_5736,N_5128);
nor U7374 (N_7374,N_5049,N_3033);
or U7375 (N_7375,N_3879,N_3092);
or U7376 (N_7376,N_3038,N_5640);
or U7377 (N_7377,N_4611,N_4012);
or U7378 (N_7378,N_4358,N_4071);
and U7379 (N_7379,N_4529,N_3419);
and U7380 (N_7380,N_4048,N_4252);
nand U7381 (N_7381,N_5201,N_3245);
or U7382 (N_7382,N_4647,N_3836);
nand U7383 (N_7383,N_4282,N_3034);
and U7384 (N_7384,N_4312,N_5067);
nand U7385 (N_7385,N_5018,N_4825);
nand U7386 (N_7386,N_4511,N_4780);
nand U7387 (N_7387,N_3702,N_3296);
nand U7388 (N_7388,N_5120,N_4684);
xor U7389 (N_7389,N_4258,N_5722);
xnor U7390 (N_7390,N_5294,N_4398);
or U7391 (N_7391,N_5002,N_4332);
and U7392 (N_7392,N_5542,N_3398);
nor U7393 (N_7393,N_5495,N_5115);
and U7394 (N_7394,N_4178,N_4276);
and U7395 (N_7395,N_4389,N_4030);
nor U7396 (N_7396,N_3351,N_3876);
nand U7397 (N_7397,N_4730,N_4393);
and U7398 (N_7398,N_3111,N_3867);
or U7399 (N_7399,N_4703,N_5800);
and U7400 (N_7400,N_4422,N_3512);
or U7401 (N_7401,N_4889,N_4659);
and U7402 (N_7402,N_5888,N_5277);
and U7403 (N_7403,N_3765,N_5928);
nor U7404 (N_7404,N_5659,N_4350);
nand U7405 (N_7405,N_4732,N_5158);
xnor U7406 (N_7406,N_4605,N_5477);
xor U7407 (N_7407,N_3900,N_5707);
nand U7408 (N_7408,N_3761,N_5146);
or U7409 (N_7409,N_5172,N_4817);
and U7410 (N_7410,N_5238,N_3671);
nand U7411 (N_7411,N_3469,N_5957);
nand U7412 (N_7412,N_5409,N_5853);
or U7413 (N_7413,N_5198,N_5681);
nor U7414 (N_7414,N_3816,N_3173);
xnor U7415 (N_7415,N_4768,N_4165);
or U7416 (N_7416,N_4386,N_3947);
nor U7417 (N_7417,N_5066,N_4895);
nand U7418 (N_7418,N_4188,N_3940);
and U7419 (N_7419,N_3470,N_5593);
nand U7420 (N_7420,N_3926,N_5869);
nand U7421 (N_7421,N_3199,N_3250);
or U7422 (N_7422,N_3074,N_5712);
or U7423 (N_7423,N_5450,N_4921);
and U7424 (N_7424,N_4054,N_3707);
nor U7425 (N_7425,N_5260,N_4053);
or U7426 (N_7426,N_4138,N_4191);
or U7427 (N_7427,N_3294,N_4074);
or U7428 (N_7428,N_3259,N_4945);
nand U7429 (N_7429,N_3124,N_5588);
nand U7430 (N_7430,N_5180,N_5518);
xnor U7431 (N_7431,N_3238,N_3744);
nor U7432 (N_7432,N_3172,N_5909);
or U7433 (N_7433,N_4615,N_5204);
or U7434 (N_7434,N_5881,N_5893);
nand U7435 (N_7435,N_5153,N_3208);
xor U7436 (N_7436,N_4049,N_5486);
nand U7437 (N_7437,N_3335,N_3501);
and U7438 (N_7438,N_3930,N_4873);
nor U7439 (N_7439,N_5697,N_5029);
and U7440 (N_7440,N_4092,N_4190);
nor U7441 (N_7441,N_5427,N_4494);
or U7442 (N_7442,N_4383,N_3888);
nand U7443 (N_7443,N_4062,N_3664);
xor U7444 (N_7444,N_4489,N_4919);
nand U7445 (N_7445,N_3605,N_3122);
or U7446 (N_7446,N_5935,N_3288);
nor U7447 (N_7447,N_5809,N_3920);
nor U7448 (N_7448,N_4056,N_5160);
or U7449 (N_7449,N_3646,N_3992);
nor U7450 (N_7450,N_4907,N_3616);
nand U7451 (N_7451,N_5480,N_5544);
and U7452 (N_7452,N_4217,N_3725);
nor U7453 (N_7453,N_3721,N_4432);
xor U7454 (N_7454,N_4551,N_5550);
xor U7455 (N_7455,N_5835,N_4955);
or U7456 (N_7456,N_5346,N_3893);
and U7457 (N_7457,N_5643,N_4151);
nor U7458 (N_7458,N_5088,N_3471);
or U7459 (N_7459,N_4111,N_5584);
and U7460 (N_7460,N_4721,N_5254);
nand U7461 (N_7461,N_4091,N_3165);
xnor U7462 (N_7462,N_4748,N_5159);
nor U7463 (N_7463,N_5562,N_5356);
xnor U7464 (N_7464,N_4793,N_3431);
nor U7465 (N_7465,N_5724,N_3863);
nand U7466 (N_7466,N_5967,N_5646);
and U7467 (N_7467,N_3271,N_4521);
and U7468 (N_7468,N_4501,N_3741);
nor U7469 (N_7469,N_3484,N_3676);
and U7470 (N_7470,N_4243,N_3981);
or U7471 (N_7471,N_5299,N_3796);
and U7472 (N_7472,N_5879,N_3763);
and U7473 (N_7473,N_4966,N_3010);
or U7474 (N_7474,N_5264,N_3932);
and U7475 (N_7475,N_5373,N_5534);
nor U7476 (N_7476,N_3609,N_4770);
nor U7477 (N_7477,N_4077,N_5406);
nand U7478 (N_7478,N_3461,N_5410);
nand U7479 (N_7479,N_4856,N_4127);
or U7480 (N_7480,N_3963,N_5699);
or U7481 (N_7481,N_5166,N_4759);
nor U7482 (N_7482,N_3439,N_5191);
or U7483 (N_7483,N_3872,N_4512);
nor U7484 (N_7484,N_4250,N_3375);
and U7485 (N_7485,N_3906,N_5122);
and U7486 (N_7486,N_5175,N_5864);
nand U7487 (N_7487,N_3300,N_5812);
and U7488 (N_7488,N_4639,N_4396);
xor U7489 (N_7489,N_3545,N_3084);
nand U7490 (N_7490,N_3317,N_4278);
or U7491 (N_7491,N_5611,N_4545);
or U7492 (N_7492,N_5075,N_3362);
nand U7493 (N_7493,N_4763,N_4882);
nor U7494 (N_7494,N_3973,N_3225);
and U7495 (N_7495,N_5003,N_3747);
and U7496 (N_7496,N_5353,N_4534);
nand U7497 (N_7497,N_3798,N_5892);
and U7498 (N_7498,N_5751,N_5451);
nand U7499 (N_7499,N_4228,N_5516);
and U7500 (N_7500,N_5120,N_4740);
and U7501 (N_7501,N_3877,N_4633);
nand U7502 (N_7502,N_3845,N_3608);
nor U7503 (N_7503,N_5068,N_3911);
nand U7504 (N_7504,N_5289,N_5842);
nand U7505 (N_7505,N_3279,N_5244);
and U7506 (N_7506,N_3985,N_4042);
nor U7507 (N_7507,N_4162,N_3981);
nand U7508 (N_7508,N_5187,N_3611);
nand U7509 (N_7509,N_3869,N_4543);
nand U7510 (N_7510,N_4553,N_5463);
and U7511 (N_7511,N_3432,N_5121);
or U7512 (N_7512,N_3696,N_5760);
nand U7513 (N_7513,N_5629,N_3459);
or U7514 (N_7514,N_3108,N_3726);
nand U7515 (N_7515,N_4133,N_4038);
xnor U7516 (N_7516,N_3940,N_4842);
nand U7517 (N_7517,N_5228,N_3113);
and U7518 (N_7518,N_3328,N_5451);
and U7519 (N_7519,N_4597,N_5946);
xor U7520 (N_7520,N_4024,N_4666);
nand U7521 (N_7521,N_3607,N_5327);
nor U7522 (N_7522,N_4922,N_5603);
xnor U7523 (N_7523,N_4286,N_3682);
xnor U7524 (N_7524,N_5394,N_5261);
xnor U7525 (N_7525,N_3162,N_4642);
nor U7526 (N_7526,N_5514,N_5527);
nor U7527 (N_7527,N_3182,N_5006);
nand U7528 (N_7528,N_4312,N_3222);
nor U7529 (N_7529,N_5852,N_5043);
and U7530 (N_7530,N_4738,N_3586);
or U7531 (N_7531,N_3024,N_3835);
nor U7532 (N_7532,N_5272,N_4079);
or U7533 (N_7533,N_5142,N_3305);
xnor U7534 (N_7534,N_4853,N_5329);
and U7535 (N_7535,N_4804,N_5076);
nor U7536 (N_7536,N_4765,N_3715);
or U7537 (N_7537,N_5953,N_3252);
nor U7538 (N_7538,N_5773,N_3676);
nor U7539 (N_7539,N_5955,N_3429);
or U7540 (N_7540,N_4305,N_4350);
nand U7541 (N_7541,N_5676,N_4839);
and U7542 (N_7542,N_3107,N_3532);
nor U7543 (N_7543,N_3341,N_3433);
nand U7544 (N_7544,N_4305,N_3917);
and U7545 (N_7545,N_3110,N_5226);
or U7546 (N_7546,N_4576,N_4141);
xor U7547 (N_7547,N_5525,N_3853);
and U7548 (N_7548,N_5144,N_5949);
nor U7549 (N_7549,N_3896,N_3676);
nand U7550 (N_7550,N_4256,N_5776);
nor U7551 (N_7551,N_4985,N_5951);
xor U7552 (N_7552,N_5916,N_5014);
nand U7553 (N_7553,N_3491,N_3570);
nor U7554 (N_7554,N_5641,N_4294);
xnor U7555 (N_7555,N_5741,N_5942);
nand U7556 (N_7556,N_5878,N_4647);
and U7557 (N_7557,N_4327,N_4404);
nand U7558 (N_7558,N_3137,N_5896);
nand U7559 (N_7559,N_5696,N_5822);
and U7560 (N_7560,N_5406,N_4950);
and U7561 (N_7561,N_4405,N_4145);
or U7562 (N_7562,N_3773,N_5409);
nor U7563 (N_7563,N_3587,N_5428);
nand U7564 (N_7564,N_4053,N_5711);
xnor U7565 (N_7565,N_3683,N_3541);
nor U7566 (N_7566,N_4495,N_5621);
and U7567 (N_7567,N_3803,N_3603);
nor U7568 (N_7568,N_3639,N_3992);
nor U7569 (N_7569,N_5685,N_5269);
or U7570 (N_7570,N_4702,N_4777);
xnor U7571 (N_7571,N_3561,N_5839);
nand U7572 (N_7572,N_3106,N_3638);
xor U7573 (N_7573,N_5838,N_5065);
nor U7574 (N_7574,N_3399,N_4617);
nand U7575 (N_7575,N_3590,N_4659);
nor U7576 (N_7576,N_4637,N_3774);
and U7577 (N_7577,N_4604,N_4112);
xor U7578 (N_7578,N_4086,N_3336);
nor U7579 (N_7579,N_3434,N_3185);
and U7580 (N_7580,N_5709,N_5749);
nand U7581 (N_7581,N_4666,N_5340);
nand U7582 (N_7582,N_5837,N_5860);
and U7583 (N_7583,N_5482,N_3524);
xnor U7584 (N_7584,N_4116,N_5770);
or U7585 (N_7585,N_5423,N_5860);
or U7586 (N_7586,N_4395,N_3875);
and U7587 (N_7587,N_5787,N_4291);
and U7588 (N_7588,N_4033,N_4126);
xor U7589 (N_7589,N_5025,N_3649);
nand U7590 (N_7590,N_3326,N_5145);
and U7591 (N_7591,N_4161,N_5725);
or U7592 (N_7592,N_3551,N_5747);
nand U7593 (N_7593,N_3840,N_3166);
nor U7594 (N_7594,N_4733,N_4564);
nand U7595 (N_7595,N_3633,N_4691);
or U7596 (N_7596,N_5745,N_4476);
nor U7597 (N_7597,N_5125,N_3717);
nand U7598 (N_7598,N_4077,N_5332);
or U7599 (N_7599,N_3738,N_5228);
nand U7600 (N_7600,N_3200,N_5820);
or U7601 (N_7601,N_3385,N_3787);
and U7602 (N_7602,N_5258,N_4009);
xnor U7603 (N_7603,N_5292,N_4838);
nor U7604 (N_7604,N_3137,N_4705);
or U7605 (N_7605,N_4012,N_4375);
nand U7606 (N_7606,N_5902,N_3082);
or U7607 (N_7607,N_5164,N_4145);
nand U7608 (N_7608,N_5044,N_4539);
and U7609 (N_7609,N_3415,N_4382);
nand U7610 (N_7610,N_4328,N_3065);
nor U7611 (N_7611,N_5041,N_4828);
nand U7612 (N_7612,N_4218,N_5551);
nor U7613 (N_7613,N_5142,N_3791);
nand U7614 (N_7614,N_3382,N_4003);
nor U7615 (N_7615,N_4693,N_3911);
or U7616 (N_7616,N_3393,N_5708);
nor U7617 (N_7617,N_4607,N_4210);
nand U7618 (N_7618,N_4662,N_4244);
and U7619 (N_7619,N_3802,N_4245);
nand U7620 (N_7620,N_3240,N_4946);
and U7621 (N_7621,N_3952,N_4724);
or U7622 (N_7622,N_4218,N_3701);
nand U7623 (N_7623,N_3877,N_3205);
and U7624 (N_7624,N_3071,N_5337);
nand U7625 (N_7625,N_3577,N_5338);
and U7626 (N_7626,N_3547,N_5708);
and U7627 (N_7627,N_5701,N_3724);
nor U7628 (N_7628,N_4910,N_3106);
or U7629 (N_7629,N_3586,N_4885);
xnor U7630 (N_7630,N_5695,N_4394);
or U7631 (N_7631,N_5727,N_3097);
or U7632 (N_7632,N_3829,N_4116);
nand U7633 (N_7633,N_5597,N_3145);
and U7634 (N_7634,N_5714,N_5067);
and U7635 (N_7635,N_5530,N_4837);
and U7636 (N_7636,N_3785,N_4461);
nor U7637 (N_7637,N_5366,N_5982);
or U7638 (N_7638,N_3209,N_4278);
nor U7639 (N_7639,N_3226,N_5723);
xor U7640 (N_7640,N_4261,N_3247);
and U7641 (N_7641,N_4645,N_5480);
and U7642 (N_7642,N_4721,N_3677);
nand U7643 (N_7643,N_3906,N_3938);
xor U7644 (N_7644,N_4126,N_4341);
or U7645 (N_7645,N_3313,N_5178);
xnor U7646 (N_7646,N_4470,N_5507);
and U7647 (N_7647,N_5910,N_5885);
nor U7648 (N_7648,N_4642,N_3043);
nor U7649 (N_7649,N_3757,N_5402);
nand U7650 (N_7650,N_4605,N_4882);
or U7651 (N_7651,N_3759,N_4722);
nor U7652 (N_7652,N_3273,N_5274);
xnor U7653 (N_7653,N_5273,N_4025);
nor U7654 (N_7654,N_5714,N_5434);
xnor U7655 (N_7655,N_5856,N_3865);
nor U7656 (N_7656,N_4862,N_3214);
nor U7657 (N_7657,N_3686,N_5506);
xor U7658 (N_7658,N_5167,N_5776);
nor U7659 (N_7659,N_3479,N_4158);
and U7660 (N_7660,N_5737,N_4260);
nor U7661 (N_7661,N_5446,N_5920);
nor U7662 (N_7662,N_5679,N_5422);
and U7663 (N_7663,N_4104,N_4281);
nand U7664 (N_7664,N_3950,N_4648);
nor U7665 (N_7665,N_5069,N_3935);
or U7666 (N_7666,N_5407,N_5530);
nand U7667 (N_7667,N_5475,N_4879);
nor U7668 (N_7668,N_4863,N_4188);
or U7669 (N_7669,N_3893,N_4100);
nand U7670 (N_7670,N_5003,N_5913);
and U7671 (N_7671,N_4954,N_3266);
nor U7672 (N_7672,N_5576,N_4944);
and U7673 (N_7673,N_3259,N_5868);
and U7674 (N_7674,N_4477,N_3742);
or U7675 (N_7675,N_4852,N_4109);
xnor U7676 (N_7676,N_5065,N_3526);
and U7677 (N_7677,N_5889,N_4564);
or U7678 (N_7678,N_3853,N_3762);
nand U7679 (N_7679,N_3541,N_4965);
and U7680 (N_7680,N_5421,N_5345);
or U7681 (N_7681,N_3011,N_5179);
xnor U7682 (N_7682,N_5626,N_4863);
xor U7683 (N_7683,N_3218,N_3935);
xor U7684 (N_7684,N_4454,N_5439);
nand U7685 (N_7685,N_4256,N_3917);
or U7686 (N_7686,N_5384,N_5748);
nand U7687 (N_7687,N_3496,N_4528);
and U7688 (N_7688,N_5120,N_4295);
or U7689 (N_7689,N_3366,N_4900);
and U7690 (N_7690,N_5034,N_5035);
nand U7691 (N_7691,N_4327,N_4157);
and U7692 (N_7692,N_5977,N_4703);
nor U7693 (N_7693,N_4085,N_4290);
xnor U7694 (N_7694,N_3679,N_4730);
nand U7695 (N_7695,N_3085,N_5216);
nand U7696 (N_7696,N_3943,N_4216);
nand U7697 (N_7697,N_3532,N_5189);
or U7698 (N_7698,N_5324,N_5545);
nand U7699 (N_7699,N_5481,N_4141);
nor U7700 (N_7700,N_3157,N_4381);
nand U7701 (N_7701,N_3188,N_4934);
and U7702 (N_7702,N_4432,N_3930);
and U7703 (N_7703,N_5783,N_3765);
nand U7704 (N_7704,N_3418,N_3858);
nor U7705 (N_7705,N_5665,N_5494);
xnor U7706 (N_7706,N_4917,N_4265);
and U7707 (N_7707,N_5336,N_3198);
nor U7708 (N_7708,N_4053,N_3141);
nor U7709 (N_7709,N_3912,N_3352);
nand U7710 (N_7710,N_4419,N_4334);
or U7711 (N_7711,N_5452,N_5648);
nand U7712 (N_7712,N_5333,N_3880);
or U7713 (N_7713,N_4634,N_4207);
xnor U7714 (N_7714,N_4845,N_3117);
and U7715 (N_7715,N_5000,N_4950);
nand U7716 (N_7716,N_3098,N_3409);
and U7717 (N_7717,N_3534,N_3684);
and U7718 (N_7718,N_5273,N_3839);
xnor U7719 (N_7719,N_4249,N_5820);
or U7720 (N_7720,N_3282,N_4805);
nand U7721 (N_7721,N_3125,N_3067);
nor U7722 (N_7722,N_4061,N_5855);
or U7723 (N_7723,N_4058,N_3896);
or U7724 (N_7724,N_4756,N_3661);
xnor U7725 (N_7725,N_3880,N_5232);
nor U7726 (N_7726,N_5452,N_5000);
and U7727 (N_7727,N_5374,N_5352);
and U7728 (N_7728,N_4842,N_4243);
nor U7729 (N_7729,N_5131,N_4778);
nand U7730 (N_7730,N_3151,N_4150);
and U7731 (N_7731,N_5505,N_4708);
and U7732 (N_7732,N_5304,N_4054);
nand U7733 (N_7733,N_5499,N_5659);
nand U7734 (N_7734,N_3873,N_5379);
or U7735 (N_7735,N_3225,N_3441);
or U7736 (N_7736,N_4557,N_3432);
nor U7737 (N_7737,N_5174,N_3351);
and U7738 (N_7738,N_3853,N_3332);
nor U7739 (N_7739,N_5449,N_4546);
nand U7740 (N_7740,N_5508,N_5780);
and U7741 (N_7741,N_3211,N_3084);
and U7742 (N_7742,N_3365,N_4597);
and U7743 (N_7743,N_4057,N_5675);
xor U7744 (N_7744,N_4788,N_5393);
and U7745 (N_7745,N_5770,N_5022);
nand U7746 (N_7746,N_4134,N_4809);
and U7747 (N_7747,N_3216,N_3945);
or U7748 (N_7748,N_4776,N_4487);
nor U7749 (N_7749,N_3690,N_5610);
nand U7750 (N_7750,N_4469,N_4936);
nor U7751 (N_7751,N_4055,N_5417);
or U7752 (N_7752,N_5293,N_4215);
or U7753 (N_7753,N_3233,N_5264);
nand U7754 (N_7754,N_4798,N_3895);
nor U7755 (N_7755,N_4302,N_5600);
nand U7756 (N_7756,N_3984,N_5139);
or U7757 (N_7757,N_5081,N_5444);
xor U7758 (N_7758,N_5976,N_3019);
nand U7759 (N_7759,N_4376,N_5682);
and U7760 (N_7760,N_3558,N_3519);
nand U7761 (N_7761,N_4154,N_5807);
and U7762 (N_7762,N_5598,N_3757);
nor U7763 (N_7763,N_3688,N_5050);
nor U7764 (N_7764,N_4970,N_3389);
xnor U7765 (N_7765,N_3409,N_5689);
nor U7766 (N_7766,N_4584,N_3531);
and U7767 (N_7767,N_4211,N_5024);
nor U7768 (N_7768,N_3167,N_5768);
nor U7769 (N_7769,N_4725,N_3639);
or U7770 (N_7770,N_4492,N_4336);
and U7771 (N_7771,N_3824,N_5607);
nor U7772 (N_7772,N_5247,N_3441);
or U7773 (N_7773,N_3735,N_3055);
nor U7774 (N_7774,N_4349,N_5149);
nand U7775 (N_7775,N_4426,N_5253);
nand U7776 (N_7776,N_5384,N_5681);
xnor U7777 (N_7777,N_4002,N_5213);
nand U7778 (N_7778,N_3566,N_3243);
or U7779 (N_7779,N_5703,N_3112);
and U7780 (N_7780,N_4340,N_4601);
or U7781 (N_7781,N_3208,N_3942);
and U7782 (N_7782,N_5430,N_4207);
nand U7783 (N_7783,N_3764,N_5289);
or U7784 (N_7784,N_3367,N_4608);
nor U7785 (N_7785,N_3945,N_5823);
nand U7786 (N_7786,N_4672,N_5630);
nand U7787 (N_7787,N_5634,N_3680);
nand U7788 (N_7788,N_3484,N_5899);
nor U7789 (N_7789,N_5823,N_4739);
or U7790 (N_7790,N_4082,N_5354);
or U7791 (N_7791,N_4958,N_3384);
nor U7792 (N_7792,N_4728,N_3803);
or U7793 (N_7793,N_3422,N_4222);
or U7794 (N_7794,N_3054,N_4255);
nand U7795 (N_7795,N_4854,N_3112);
nor U7796 (N_7796,N_4719,N_5967);
nor U7797 (N_7797,N_4285,N_5443);
or U7798 (N_7798,N_5232,N_3426);
nand U7799 (N_7799,N_3173,N_5834);
nor U7800 (N_7800,N_3190,N_3842);
or U7801 (N_7801,N_4602,N_5909);
or U7802 (N_7802,N_3192,N_3011);
nor U7803 (N_7803,N_4499,N_4943);
nor U7804 (N_7804,N_5374,N_4023);
and U7805 (N_7805,N_4442,N_3195);
or U7806 (N_7806,N_4824,N_3912);
nand U7807 (N_7807,N_4580,N_3843);
or U7808 (N_7808,N_5435,N_4232);
and U7809 (N_7809,N_3195,N_4821);
and U7810 (N_7810,N_4812,N_3256);
nand U7811 (N_7811,N_3019,N_5573);
and U7812 (N_7812,N_5983,N_4653);
nand U7813 (N_7813,N_4265,N_3259);
xor U7814 (N_7814,N_4047,N_3688);
nand U7815 (N_7815,N_5876,N_5110);
and U7816 (N_7816,N_4340,N_5421);
nor U7817 (N_7817,N_3470,N_5950);
nor U7818 (N_7818,N_3443,N_5724);
nor U7819 (N_7819,N_5085,N_5834);
xor U7820 (N_7820,N_5058,N_5502);
nor U7821 (N_7821,N_5480,N_4217);
or U7822 (N_7822,N_4253,N_5246);
nor U7823 (N_7823,N_4928,N_5944);
nand U7824 (N_7824,N_5293,N_5784);
xnor U7825 (N_7825,N_3702,N_4022);
nand U7826 (N_7826,N_5072,N_3202);
nand U7827 (N_7827,N_5640,N_5222);
or U7828 (N_7828,N_5218,N_3354);
and U7829 (N_7829,N_4145,N_4540);
nand U7830 (N_7830,N_4124,N_5841);
or U7831 (N_7831,N_4242,N_4708);
and U7832 (N_7832,N_4449,N_3700);
or U7833 (N_7833,N_3307,N_5346);
or U7834 (N_7834,N_3281,N_3197);
nor U7835 (N_7835,N_4958,N_3524);
and U7836 (N_7836,N_4510,N_4988);
nor U7837 (N_7837,N_4340,N_5264);
nand U7838 (N_7838,N_5342,N_5748);
xnor U7839 (N_7839,N_3591,N_3726);
and U7840 (N_7840,N_3707,N_5373);
nor U7841 (N_7841,N_5349,N_4943);
nor U7842 (N_7842,N_5016,N_4407);
nor U7843 (N_7843,N_4285,N_5015);
or U7844 (N_7844,N_5061,N_4978);
nor U7845 (N_7845,N_3245,N_3907);
and U7846 (N_7846,N_4257,N_3108);
and U7847 (N_7847,N_3861,N_4560);
xnor U7848 (N_7848,N_4937,N_5540);
nor U7849 (N_7849,N_5273,N_3793);
and U7850 (N_7850,N_4120,N_3911);
nor U7851 (N_7851,N_3971,N_5111);
and U7852 (N_7852,N_5868,N_3088);
xor U7853 (N_7853,N_3649,N_5386);
nand U7854 (N_7854,N_5697,N_4041);
and U7855 (N_7855,N_3678,N_3221);
and U7856 (N_7856,N_5233,N_5441);
nor U7857 (N_7857,N_5903,N_3182);
or U7858 (N_7858,N_5201,N_3377);
or U7859 (N_7859,N_3324,N_5653);
and U7860 (N_7860,N_3558,N_3152);
nor U7861 (N_7861,N_5956,N_3330);
or U7862 (N_7862,N_3364,N_4743);
nor U7863 (N_7863,N_3369,N_5979);
nand U7864 (N_7864,N_4725,N_3042);
nor U7865 (N_7865,N_3809,N_3367);
nand U7866 (N_7866,N_4178,N_5778);
nor U7867 (N_7867,N_4127,N_5397);
and U7868 (N_7868,N_3449,N_3101);
and U7869 (N_7869,N_3457,N_4580);
or U7870 (N_7870,N_3961,N_5463);
and U7871 (N_7871,N_5050,N_4347);
nor U7872 (N_7872,N_5240,N_4379);
or U7873 (N_7873,N_5003,N_5230);
xor U7874 (N_7874,N_3293,N_4475);
and U7875 (N_7875,N_3403,N_5631);
or U7876 (N_7876,N_5335,N_5675);
xor U7877 (N_7877,N_5994,N_3541);
nand U7878 (N_7878,N_5560,N_5265);
or U7879 (N_7879,N_4734,N_3628);
nor U7880 (N_7880,N_3347,N_3208);
nand U7881 (N_7881,N_4755,N_3054);
nand U7882 (N_7882,N_5625,N_3628);
or U7883 (N_7883,N_4840,N_4830);
and U7884 (N_7884,N_5946,N_5512);
nand U7885 (N_7885,N_4030,N_4198);
or U7886 (N_7886,N_4109,N_5215);
nor U7887 (N_7887,N_5431,N_3550);
and U7888 (N_7888,N_5418,N_3842);
xor U7889 (N_7889,N_5627,N_3310);
or U7890 (N_7890,N_3156,N_4883);
and U7891 (N_7891,N_4972,N_4491);
nor U7892 (N_7892,N_4435,N_4960);
and U7893 (N_7893,N_3148,N_4782);
and U7894 (N_7894,N_3650,N_5880);
xnor U7895 (N_7895,N_5271,N_4688);
nand U7896 (N_7896,N_3257,N_4786);
xor U7897 (N_7897,N_3982,N_3799);
nand U7898 (N_7898,N_4812,N_5512);
nor U7899 (N_7899,N_5341,N_4544);
nor U7900 (N_7900,N_3649,N_3392);
and U7901 (N_7901,N_4890,N_4814);
nor U7902 (N_7902,N_4715,N_3899);
nor U7903 (N_7903,N_3740,N_5249);
nor U7904 (N_7904,N_3085,N_5346);
and U7905 (N_7905,N_4422,N_3380);
xnor U7906 (N_7906,N_3973,N_5674);
nor U7907 (N_7907,N_4542,N_4505);
nand U7908 (N_7908,N_4829,N_3043);
nand U7909 (N_7909,N_4672,N_5151);
or U7910 (N_7910,N_5901,N_5948);
nand U7911 (N_7911,N_3919,N_4063);
or U7912 (N_7912,N_5051,N_4176);
nand U7913 (N_7913,N_3400,N_3429);
xor U7914 (N_7914,N_3381,N_4645);
or U7915 (N_7915,N_4051,N_3179);
or U7916 (N_7916,N_4622,N_3620);
or U7917 (N_7917,N_4816,N_5922);
or U7918 (N_7918,N_4818,N_3176);
nand U7919 (N_7919,N_5096,N_5769);
or U7920 (N_7920,N_4961,N_4456);
and U7921 (N_7921,N_5836,N_4784);
nor U7922 (N_7922,N_3062,N_4176);
and U7923 (N_7923,N_4048,N_4500);
nand U7924 (N_7924,N_3121,N_5319);
xor U7925 (N_7925,N_4386,N_4286);
and U7926 (N_7926,N_3989,N_3325);
nor U7927 (N_7927,N_4852,N_4142);
or U7928 (N_7928,N_4235,N_5251);
nor U7929 (N_7929,N_4130,N_4833);
or U7930 (N_7930,N_5386,N_4427);
and U7931 (N_7931,N_4659,N_5165);
nand U7932 (N_7932,N_4947,N_5729);
nand U7933 (N_7933,N_5330,N_4397);
or U7934 (N_7934,N_4633,N_5147);
nor U7935 (N_7935,N_4868,N_4778);
and U7936 (N_7936,N_3467,N_5829);
nand U7937 (N_7937,N_5498,N_4461);
or U7938 (N_7938,N_5697,N_3220);
or U7939 (N_7939,N_3709,N_5618);
nand U7940 (N_7940,N_3221,N_5992);
or U7941 (N_7941,N_5943,N_4019);
nor U7942 (N_7942,N_5800,N_4744);
nand U7943 (N_7943,N_4927,N_3039);
xor U7944 (N_7944,N_5973,N_4247);
nand U7945 (N_7945,N_3110,N_5371);
nand U7946 (N_7946,N_3966,N_3280);
and U7947 (N_7947,N_5133,N_5120);
nand U7948 (N_7948,N_5176,N_5893);
or U7949 (N_7949,N_4742,N_3685);
xor U7950 (N_7950,N_4512,N_5804);
nand U7951 (N_7951,N_4665,N_3619);
nand U7952 (N_7952,N_3613,N_3129);
and U7953 (N_7953,N_5057,N_3528);
nor U7954 (N_7954,N_4100,N_5694);
or U7955 (N_7955,N_5381,N_4777);
nand U7956 (N_7956,N_3966,N_4503);
or U7957 (N_7957,N_4407,N_4352);
nand U7958 (N_7958,N_3148,N_4512);
nand U7959 (N_7959,N_4049,N_3879);
nor U7960 (N_7960,N_4629,N_4006);
xnor U7961 (N_7961,N_5213,N_3952);
xnor U7962 (N_7962,N_5716,N_5337);
and U7963 (N_7963,N_5488,N_5516);
nand U7964 (N_7964,N_4483,N_4195);
nor U7965 (N_7965,N_4936,N_5840);
nand U7966 (N_7966,N_4657,N_3462);
xor U7967 (N_7967,N_5645,N_3237);
nor U7968 (N_7968,N_4053,N_3945);
and U7969 (N_7969,N_4526,N_5430);
and U7970 (N_7970,N_5495,N_4828);
nand U7971 (N_7971,N_4034,N_5816);
nor U7972 (N_7972,N_5233,N_5874);
xor U7973 (N_7973,N_4689,N_5255);
xnor U7974 (N_7974,N_4126,N_5718);
and U7975 (N_7975,N_3761,N_4301);
nor U7976 (N_7976,N_3624,N_4375);
and U7977 (N_7977,N_4836,N_4336);
nor U7978 (N_7978,N_5334,N_3397);
nand U7979 (N_7979,N_4156,N_3943);
or U7980 (N_7980,N_3150,N_4258);
nand U7981 (N_7981,N_3934,N_5288);
or U7982 (N_7982,N_5435,N_3507);
nand U7983 (N_7983,N_3721,N_3691);
or U7984 (N_7984,N_3303,N_3258);
nor U7985 (N_7985,N_3842,N_4862);
and U7986 (N_7986,N_4672,N_4305);
or U7987 (N_7987,N_4842,N_4976);
nor U7988 (N_7988,N_4345,N_3343);
nor U7989 (N_7989,N_5650,N_4387);
nand U7990 (N_7990,N_4751,N_4078);
nor U7991 (N_7991,N_5286,N_5686);
nor U7992 (N_7992,N_5327,N_5409);
nand U7993 (N_7993,N_3723,N_5153);
and U7994 (N_7994,N_3573,N_5896);
or U7995 (N_7995,N_5936,N_5935);
and U7996 (N_7996,N_3383,N_3110);
nor U7997 (N_7997,N_5123,N_5502);
xor U7998 (N_7998,N_4778,N_3344);
and U7999 (N_7999,N_5034,N_4915);
nand U8000 (N_8000,N_5972,N_3349);
or U8001 (N_8001,N_3672,N_3271);
or U8002 (N_8002,N_3958,N_3713);
and U8003 (N_8003,N_5255,N_5556);
xnor U8004 (N_8004,N_4570,N_3755);
and U8005 (N_8005,N_3009,N_4975);
and U8006 (N_8006,N_4692,N_5875);
nor U8007 (N_8007,N_5072,N_3999);
and U8008 (N_8008,N_5366,N_5183);
nand U8009 (N_8009,N_4878,N_5371);
xor U8010 (N_8010,N_5808,N_3348);
xor U8011 (N_8011,N_5487,N_4132);
and U8012 (N_8012,N_4013,N_5146);
nor U8013 (N_8013,N_3681,N_3514);
xnor U8014 (N_8014,N_3530,N_3950);
nor U8015 (N_8015,N_4814,N_3233);
nor U8016 (N_8016,N_5415,N_4420);
nand U8017 (N_8017,N_5967,N_3727);
or U8018 (N_8018,N_4248,N_3450);
or U8019 (N_8019,N_4966,N_3274);
and U8020 (N_8020,N_3189,N_3651);
nor U8021 (N_8021,N_5616,N_5913);
xor U8022 (N_8022,N_3230,N_4172);
xnor U8023 (N_8023,N_4563,N_3654);
nand U8024 (N_8024,N_5332,N_4244);
nor U8025 (N_8025,N_5812,N_5505);
or U8026 (N_8026,N_3079,N_5069);
nand U8027 (N_8027,N_4729,N_5828);
nor U8028 (N_8028,N_3379,N_3364);
and U8029 (N_8029,N_4229,N_5210);
nor U8030 (N_8030,N_4144,N_4975);
xnor U8031 (N_8031,N_4229,N_3521);
or U8032 (N_8032,N_4824,N_4247);
nor U8033 (N_8033,N_4190,N_3614);
nand U8034 (N_8034,N_3209,N_3477);
nor U8035 (N_8035,N_4731,N_5963);
or U8036 (N_8036,N_4487,N_3021);
or U8037 (N_8037,N_5946,N_5999);
and U8038 (N_8038,N_5142,N_5003);
or U8039 (N_8039,N_5459,N_5242);
nor U8040 (N_8040,N_5295,N_5791);
nand U8041 (N_8041,N_5983,N_4335);
or U8042 (N_8042,N_3710,N_4492);
or U8043 (N_8043,N_5599,N_4580);
and U8044 (N_8044,N_5076,N_4351);
or U8045 (N_8045,N_3137,N_5583);
and U8046 (N_8046,N_3651,N_3830);
and U8047 (N_8047,N_5730,N_3455);
nor U8048 (N_8048,N_3600,N_4289);
xor U8049 (N_8049,N_3619,N_4084);
nand U8050 (N_8050,N_5461,N_5975);
and U8051 (N_8051,N_5198,N_3225);
nand U8052 (N_8052,N_4345,N_3497);
nor U8053 (N_8053,N_5177,N_3712);
nand U8054 (N_8054,N_4169,N_3422);
nor U8055 (N_8055,N_5731,N_5210);
and U8056 (N_8056,N_4900,N_4331);
or U8057 (N_8057,N_5410,N_4373);
and U8058 (N_8058,N_4957,N_3425);
nand U8059 (N_8059,N_4376,N_3868);
or U8060 (N_8060,N_4113,N_3315);
nor U8061 (N_8061,N_4231,N_3334);
xor U8062 (N_8062,N_5302,N_4968);
or U8063 (N_8063,N_4057,N_5570);
or U8064 (N_8064,N_5928,N_3776);
nand U8065 (N_8065,N_4626,N_4661);
or U8066 (N_8066,N_5073,N_5137);
nor U8067 (N_8067,N_5213,N_4253);
nand U8068 (N_8068,N_5468,N_3564);
nand U8069 (N_8069,N_4885,N_3731);
and U8070 (N_8070,N_5032,N_4652);
nor U8071 (N_8071,N_4195,N_5423);
nand U8072 (N_8072,N_4001,N_4450);
nor U8073 (N_8073,N_5193,N_5041);
nor U8074 (N_8074,N_5870,N_5003);
and U8075 (N_8075,N_4568,N_5229);
or U8076 (N_8076,N_5249,N_3041);
nand U8077 (N_8077,N_5336,N_5716);
xnor U8078 (N_8078,N_5708,N_3352);
and U8079 (N_8079,N_5164,N_5731);
nor U8080 (N_8080,N_5776,N_3604);
nand U8081 (N_8081,N_4308,N_4003);
xor U8082 (N_8082,N_4704,N_5435);
nor U8083 (N_8083,N_5132,N_4828);
nand U8084 (N_8084,N_3047,N_4983);
and U8085 (N_8085,N_5094,N_5104);
nor U8086 (N_8086,N_5900,N_4499);
or U8087 (N_8087,N_3697,N_5433);
and U8088 (N_8088,N_3259,N_3733);
or U8089 (N_8089,N_4847,N_3705);
nor U8090 (N_8090,N_3794,N_4022);
or U8091 (N_8091,N_4772,N_4491);
nand U8092 (N_8092,N_3057,N_4422);
nor U8093 (N_8093,N_3611,N_5709);
nand U8094 (N_8094,N_3051,N_4816);
and U8095 (N_8095,N_4931,N_5294);
or U8096 (N_8096,N_5179,N_4154);
nand U8097 (N_8097,N_5015,N_4827);
or U8098 (N_8098,N_4069,N_5970);
nand U8099 (N_8099,N_5508,N_5375);
nor U8100 (N_8100,N_3057,N_3385);
nand U8101 (N_8101,N_3437,N_4936);
and U8102 (N_8102,N_4773,N_4377);
nor U8103 (N_8103,N_5531,N_5308);
nor U8104 (N_8104,N_3723,N_4387);
nor U8105 (N_8105,N_5874,N_4254);
xor U8106 (N_8106,N_3168,N_3850);
nor U8107 (N_8107,N_3681,N_3481);
nor U8108 (N_8108,N_3507,N_4837);
or U8109 (N_8109,N_3619,N_5312);
nand U8110 (N_8110,N_5614,N_4167);
nor U8111 (N_8111,N_4901,N_4974);
nand U8112 (N_8112,N_5141,N_4260);
or U8113 (N_8113,N_3033,N_4957);
xnor U8114 (N_8114,N_4011,N_4499);
or U8115 (N_8115,N_3828,N_4325);
and U8116 (N_8116,N_5824,N_5968);
or U8117 (N_8117,N_5897,N_5125);
or U8118 (N_8118,N_5371,N_5832);
and U8119 (N_8119,N_4135,N_5380);
nand U8120 (N_8120,N_4102,N_4321);
nor U8121 (N_8121,N_4843,N_4250);
nor U8122 (N_8122,N_3894,N_5845);
nand U8123 (N_8123,N_5203,N_5951);
nor U8124 (N_8124,N_4004,N_3532);
nor U8125 (N_8125,N_4595,N_5178);
or U8126 (N_8126,N_4749,N_4761);
and U8127 (N_8127,N_4529,N_5515);
nand U8128 (N_8128,N_3597,N_4065);
and U8129 (N_8129,N_5158,N_5266);
or U8130 (N_8130,N_5915,N_4502);
xnor U8131 (N_8131,N_4386,N_3328);
xnor U8132 (N_8132,N_3731,N_5811);
nor U8133 (N_8133,N_3075,N_4639);
nor U8134 (N_8134,N_5951,N_4134);
or U8135 (N_8135,N_5692,N_5404);
nand U8136 (N_8136,N_3648,N_3727);
or U8137 (N_8137,N_5622,N_5568);
and U8138 (N_8138,N_4544,N_5383);
nor U8139 (N_8139,N_4578,N_5103);
nand U8140 (N_8140,N_5020,N_3646);
and U8141 (N_8141,N_5815,N_3173);
or U8142 (N_8142,N_4899,N_5470);
or U8143 (N_8143,N_4565,N_3472);
nand U8144 (N_8144,N_4957,N_4357);
or U8145 (N_8145,N_4593,N_4460);
xor U8146 (N_8146,N_4825,N_5680);
nand U8147 (N_8147,N_5371,N_4900);
and U8148 (N_8148,N_3167,N_3658);
nand U8149 (N_8149,N_4748,N_5596);
and U8150 (N_8150,N_4572,N_4579);
or U8151 (N_8151,N_4863,N_5904);
xnor U8152 (N_8152,N_3792,N_3018);
and U8153 (N_8153,N_5290,N_3939);
nand U8154 (N_8154,N_5601,N_4722);
and U8155 (N_8155,N_5963,N_4917);
or U8156 (N_8156,N_4050,N_5816);
and U8157 (N_8157,N_4835,N_5860);
or U8158 (N_8158,N_3735,N_5703);
or U8159 (N_8159,N_4149,N_3341);
and U8160 (N_8160,N_3338,N_3831);
nand U8161 (N_8161,N_5919,N_3050);
and U8162 (N_8162,N_3762,N_4351);
or U8163 (N_8163,N_4813,N_5576);
nand U8164 (N_8164,N_3212,N_3198);
nand U8165 (N_8165,N_3045,N_5200);
nor U8166 (N_8166,N_5524,N_4043);
nor U8167 (N_8167,N_5749,N_3294);
or U8168 (N_8168,N_3499,N_5893);
or U8169 (N_8169,N_5634,N_4868);
nand U8170 (N_8170,N_5142,N_4183);
xor U8171 (N_8171,N_5851,N_5942);
or U8172 (N_8172,N_4850,N_4600);
nor U8173 (N_8173,N_5768,N_5358);
and U8174 (N_8174,N_4061,N_5402);
or U8175 (N_8175,N_3727,N_5423);
and U8176 (N_8176,N_5994,N_4480);
and U8177 (N_8177,N_4486,N_3224);
or U8178 (N_8178,N_5277,N_5820);
nand U8179 (N_8179,N_5556,N_5701);
and U8180 (N_8180,N_5935,N_4478);
nand U8181 (N_8181,N_4734,N_4657);
or U8182 (N_8182,N_3398,N_3926);
nor U8183 (N_8183,N_5371,N_4450);
nor U8184 (N_8184,N_3445,N_3955);
nor U8185 (N_8185,N_4665,N_3132);
and U8186 (N_8186,N_5191,N_3392);
xnor U8187 (N_8187,N_3303,N_3509);
and U8188 (N_8188,N_3135,N_4939);
and U8189 (N_8189,N_4245,N_5410);
or U8190 (N_8190,N_4936,N_4603);
nor U8191 (N_8191,N_3624,N_5235);
nand U8192 (N_8192,N_4916,N_3348);
nand U8193 (N_8193,N_3256,N_3768);
nand U8194 (N_8194,N_5958,N_5894);
nor U8195 (N_8195,N_3546,N_4039);
nand U8196 (N_8196,N_3841,N_5714);
or U8197 (N_8197,N_3524,N_3865);
nand U8198 (N_8198,N_3072,N_5845);
or U8199 (N_8199,N_4866,N_4408);
and U8200 (N_8200,N_3305,N_4457);
and U8201 (N_8201,N_4886,N_4285);
and U8202 (N_8202,N_5550,N_5509);
xor U8203 (N_8203,N_3612,N_5272);
or U8204 (N_8204,N_3999,N_5885);
and U8205 (N_8205,N_4571,N_3137);
or U8206 (N_8206,N_4954,N_4167);
nand U8207 (N_8207,N_4324,N_4468);
and U8208 (N_8208,N_3919,N_5642);
nand U8209 (N_8209,N_4802,N_5367);
xnor U8210 (N_8210,N_3791,N_3131);
nand U8211 (N_8211,N_4653,N_4006);
nor U8212 (N_8212,N_3873,N_5535);
xor U8213 (N_8213,N_5533,N_5480);
and U8214 (N_8214,N_4079,N_4685);
and U8215 (N_8215,N_3920,N_4117);
xnor U8216 (N_8216,N_3987,N_4864);
nor U8217 (N_8217,N_4664,N_5902);
nor U8218 (N_8218,N_5097,N_5524);
nand U8219 (N_8219,N_5125,N_5457);
nor U8220 (N_8220,N_3981,N_5456);
xor U8221 (N_8221,N_4045,N_3732);
nor U8222 (N_8222,N_3619,N_3788);
or U8223 (N_8223,N_5269,N_5213);
nand U8224 (N_8224,N_5192,N_4655);
and U8225 (N_8225,N_4389,N_3341);
nand U8226 (N_8226,N_4302,N_4462);
nand U8227 (N_8227,N_3470,N_3189);
and U8228 (N_8228,N_3784,N_3356);
nand U8229 (N_8229,N_4444,N_4160);
nor U8230 (N_8230,N_4443,N_5740);
or U8231 (N_8231,N_3101,N_4599);
nor U8232 (N_8232,N_4962,N_3894);
or U8233 (N_8233,N_3245,N_3289);
nor U8234 (N_8234,N_5971,N_4262);
and U8235 (N_8235,N_5077,N_5443);
nand U8236 (N_8236,N_4080,N_3515);
or U8237 (N_8237,N_5995,N_5550);
nor U8238 (N_8238,N_4189,N_4840);
or U8239 (N_8239,N_4117,N_4127);
xor U8240 (N_8240,N_5198,N_3109);
and U8241 (N_8241,N_5372,N_4260);
or U8242 (N_8242,N_4263,N_5126);
or U8243 (N_8243,N_5285,N_5882);
or U8244 (N_8244,N_3563,N_5287);
or U8245 (N_8245,N_5741,N_5353);
or U8246 (N_8246,N_5013,N_3071);
nor U8247 (N_8247,N_4526,N_5481);
and U8248 (N_8248,N_4716,N_3794);
nor U8249 (N_8249,N_4828,N_4895);
or U8250 (N_8250,N_5883,N_5217);
and U8251 (N_8251,N_3852,N_3122);
nand U8252 (N_8252,N_3325,N_3913);
or U8253 (N_8253,N_4619,N_3031);
xor U8254 (N_8254,N_5960,N_5281);
or U8255 (N_8255,N_5883,N_4365);
or U8256 (N_8256,N_4168,N_3737);
nand U8257 (N_8257,N_3765,N_5877);
nor U8258 (N_8258,N_3281,N_3297);
nand U8259 (N_8259,N_3995,N_4098);
or U8260 (N_8260,N_4820,N_4652);
nand U8261 (N_8261,N_4968,N_4127);
or U8262 (N_8262,N_3155,N_5665);
and U8263 (N_8263,N_5682,N_4222);
nand U8264 (N_8264,N_3147,N_3277);
nand U8265 (N_8265,N_4363,N_3163);
and U8266 (N_8266,N_3115,N_3322);
or U8267 (N_8267,N_4752,N_3525);
and U8268 (N_8268,N_5988,N_3624);
and U8269 (N_8269,N_5502,N_5724);
or U8270 (N_8270,N_3510,N_5341);
xnor U8271 (N_8271,N_4158,N_3761);
or U8272 (N_8272,N_4772,N_5194);
or U8273 (N_8273,N_5698,N_4794);
nand U8274 (N_8274,N_4449,N_4103);
nand U8275 (N_8275,N_4608,N_5736);
nor U8276 (N_8276,N_4794,N_5482);
xnor U8277 (N_8277,N_4354,N_3539);
or U8278 (N_8278,N_3433,N_3501);
and U8279 (N_8279,N_5813,N_4454);
or U8280 (N_8280,N_4299,N_5858);
nand U8281 (N_8281,N_3667,N_4389);
or U8282 (N_8282,N_3091,N_5851);
and U8283 (N_8283,N_4857,N_4117);
or U8284 (N_8284,N_4575,N_5260);
and U8285 (N_8285,N_3696,N_4982);
or U8286 (N_8286,N_4530,N_4751);
nor U8287 (N_8287,N_4866,N_3352);
or U8288 (N_8288,N_5948,N_4339);
or U8289 (N_8289,N_4727,N_3087);
and U8290 (N_8290,N_4583,N_3144);
or U8291 (N_8291,N_4929,N_5036);
nor U8292 (N_8292,N_5507,N_3284);
xor U8293 (N_8293,N_4477,N_5903);
xor U8294 (N_8294,N_5304,N_3403);
nand U8295 (N_8295,N_5934,N_4902);
nand U8296 (N_8296,N_3345,N_5219);
or U8297 (N_8297,N_3894,N_5471);
xor U8298 (N_8298,N_5935,N_4449);
nand U8299 (N_8299,N_5464,N_4933);
or U8300 (N_8300,N_5268,N_3311);
xor U8301 (N_8301,N_4103,N_4819);
and U8302 (N_8302,N_3090,N_5768);
xor U8303 (N_8303,N_3605,N_4715);
nand U8304 (N_8304,N_5933,N_5401);
and U8305 (N_8305,N_3300,N_5286);
xor U8306 (N_8306,N_4098,N_3703);
nand U8307 (N_8307,N_3908,N_4478);
and U8308 (N_8308,N_3997,N_4187);
xnor U8309 (N_8309,N_3960,N_4511);
or U8310 (N_8310,N_3693,N_5244);
nor U8311 (N_8311,N_3125,N_4380);
or U8312 (N_8312,N_3068,N_3238);
nor U8313 (N_8313,N_5993,N_4575);
or U8314 (N_8314,N_4882,N_4366);
nand U8315 (N_8315,N_5791,N_3717);
nor U8316 (N_8316,N_5266,N_3563);
nor U8317 (N_8317,N_4451,N_4562);
nand U8318 (N_8318,N_5303,N_4736);
or U8319 (N_8319,N_4233,N_4935);
or U8320 (N_8320,N_4750,N_4994);
nor U8321 (N_8321,N_4942,N_3788);
nand U8322 (N_8322,N_4727,N_4916);
nand U8323 (N_8323,N_4787,N_5009);
or U8324 (N_8324,N_4042,N_5193);
or U8325 (N_8325,N_4282,N_3698);
nand U8326 (N_8326,N_4725,N_3429);
nand U8327 (N_8327,N_3710,N_5801);
and U8328 (N_8328,N_5142,N_4603);
and U8329 (N_8329,N_3901,N_5308);
and U8330 (N_8330,N_5769,N_3753);
nor U8331 (N_8331,N_5806,N_4985);
nand U8332 (N_8332,N_3799,N_5762);
nor U8333 (N_8333,N_4683,N_5049);
nor U8334 (N_8334,N_4610,N_3026);
nor U8335 (N_8335,N_5224,N_3264);
and U8336 (N_8336,N_5464,N_3984);
or U8337 (N_8337,N_4779,N_3472);
and U8338 (N_8338,N_4305,N_5439);
and U8339 (N_8339,N_4867,N_3386);
nand U8340 (N_8340,N_5410,N_4382);
nand U8341 (N_8341,N_4695,N_5062);
and U8342 (N_8342,N_3278,N_4112);
xnor U8343 (N_8343,N_3364,N_5803);
nor U8344 (N_8344,N_5382,N_4060);
and U8345 (N_8345,N_4002,N_3998);
and U8346 (N_8346,N_4890,N_3692);
or U8347 (N_8347,N_4838,N_5302);
nand U8348 (N_8348,N_3931,N_3210);
nor U8349 (N_8349,N_3605,N_4592);
nor U8350 (N_8350,N_3960,N_4127);
or U8351 (N_8351,N_5793,N_5183);
nand U8352 (N_8352,N_4858,N_4849);
and U8353 (N_8353,N_4807,N_5460);
and U8354 (N_8354,N_3627,N_5813);
nand U8355 (N_8355,N_3948,N_5941);
nor U8356 (N_8356,N_4589,N_4283);
and U8357 (N_8357,N_4330,N_5554);
or U8358 (N_8358,N_3548,N_5931);
nand U8359 (N_8359,N_4823,N_4851);
nor U8360 (N_8360,N_5220,N_3345);
nor U8361 (N_8361,N_4975,N_3790);
nand U8362 (N_8362,N_4853,N_3844);
nand U8363 (N_8363,N_4278,N_5852);
or U8364 (N_8364,N_4821,N_3600);
and U8365 (N_8365,N_3653,N_5140);
or U8366 (N_8366,N_3879,N_3336);
nand U8367 (N_8367,N_5829,N_5710);
and U8368 (N_8368,N_3279,N_5208);
nor U8369 (N_8369,N_3609,N_5520);
and U8370 (N_8370,N_4309,N_4088);
nor U8371 (N_8371,N_3400,N_3841);
or U8372 (N_8372,N_3944,N_5279);
nand U8373 (N_8373,N_5278,N_5770);
nor U8374 (N_8374,N_3027,N_5893);
xnor U8375 (N_8375,N_3320,N_4221);
nor U8376 (N_8376,N_4053,N_4073);
nand U8377 (N_8377,N_4311,N_4809);
nor U8378 (N_8378,N_5427,N_4669);
or U8379 (N_8379,N_5698,N_3706);
and U8380 (N_8380,N_5656,N_4072);
nand U8381 (N_8381,N_5624,N_5499);
nor U8382 (N_8382,N_3040,N_4939);
and U8383 (N_8383,N_3101,N_4353);
nor U8384 (N_8384,N_5214,N_5931);
nor U8385 (N_8385,N_4301,N_5359);
and U8386 (N_8386,N_4107,N_3470);
or U8387 (N_8387,N_4044,N_5938);
nand U8388 (N_8388,N_5407,N_5313);
nand U8389 (N_8389,N_3520,N_5509);
or U8390 (N_8390,N_3628,N_4771);
and U8391 (N_8391,N_5304,N_4920);
or U8392 (N_8392,N_5529,N_3126);
xor U8393 (N_8393,N_5560,N_4028);
or U8394 (N_8394,N_4905,N_3227);
xnor U8395 (N_8395,N_4261,N_5395);
nor U8396 (N_8396,N_3974,N_4221);
or U8397 (N_8397,N_4137,N_4067);
nor U8398 (N_8398,N_5306,N_5403);
and U8399 (N_8399,N_5652,N_5334);
and U8400 (N_8400,N_4468,N_4268);
or U8401 (N_8401,N_4664,N_4120);
nor U8402 (N_8402,N_4957,N_3119);
and U8403 (N_8403,N_4577,N_3950);
and U8404 (N_8404,N_4241,N_5521);
xnor U8405 (N_8405,N_4917,N_5771);
nand U8406 (N_8406,N_4814,N_3822);
nand U8407 (N_8407,N_5607,N_3506);
and U8408 (N_8408,N_3537,N_3611);
or U8409 (N_8409,N_3777,N_4059);
or U8410 (N_8410,N_4238,N_3357);
nor U8411 (N_8411,N_3559,N_5337);
or U8412 (N_8412,N_5422,N_5873);
or U8413 (N_8413,N_5280,N_5212);
nand U8414 (N_8414,N_3629,N_4420);
nand U8415 (N_8415,N_5704,N_3182);
nand U8416 (N_8416,N_4395,N_4600);
xor U8417 (N_8417,N_4600,N_4720);
nand U8418 (N_8418,N_3185,N_3190);
nand U8419 (N_8419,N_3579,N_3593);
and U8420 (N_8420,N_3951,N_4681);
or U8421 (N_8421,N_3693,N_5953);
or U8422 (N_8422,N_4593,N_4606);
or U8423 (N_8423,N_5724,N_3200);
or U8424 (N_8424,N_5994,N_3371);
xnor U8425 (N_8425,N_4889,N_4958);
nor U8426 (N_8426,N_4377,N_5991);
nand U8427 (N_8427,N_5363,N_4363);
or U8428 (N_8428,N_5517,N_3721);
and U8429 (N_8429,N_3106,N_5616);
nor U8430 (N_8430,N_5656,N_3635);
and U8431 (N_8431,N_3664,N_5305);
xnor U8432 (N_8432,N_3626,N_5186);
xnor U8433 (N_8433,N_4047,N_5341);
nor U8434 (N_8434,N_4267,N_5804);
nor U8435 (N_8435,N_4148,N_4216);
and U8436 (N_8436,N_5957,N_4241);
nand U8437 (N_8437,N_5731,N_4674);
nor U8438 (N_8438,N_4702,N_3327);
nor U8439 (N_8439,N_5891,N_5139);
nor U8440 (N_8440,N_3729,N_5442);
and U8441 (N_8441,N_3346,N_3774);
or U8442 (N_8442,N_5409,N_5982);
or U8443 (N_8443,N_4720,N_5778);
nand U8444 (N_8444,N_4571,N_4622);
nor U8445 (N_8445,N_5612,N_4083);
nor U8446 (N_8446,N_4750,N_4431);
nor U8447 (N_8447,N_3253,N_5776);
or U8448 (N_8448,N_4794,N_3962);
or U8449 (N_8449,N_3071,N_4039);
nand U8450 (N_8450,N_5820,N_5432);
and U8451 (N_8451,N_3113,N_4472);
nor U8452 (N_8452,N_3890,N_3964);
xnor U8453 (N_8453,N_4673,N_4457);
and U8454 (N_8454,N_4618,N_3818);
or U8455 (N_8455,N_4520,N_3234);
nor U8456 (N_8456,N_5816,N_4821);
or U8457 (N_8457,N_4551,N_3183);
or U8458 (N_8458,N_4211,N_4774);
and U8459 (N_8459,N_5632,N_5432);
nor U8460 (N_8460,N_4540,N_3462);
or U8461 (N_8461,N_5121,N_5993);
xnor U8462 (N_8462,N_4867,N_5990);
or U8463 (N_8463,N_3505,N_4936);
nor U8464 (N_8464,N_3640,N_5195);
and U8465 (N_8465,N_3499,N_3183);
or U8466 (N_8466,N_3590,N_3730);
nand U8467 (N_8467,N_3923,N_3989);
or U8468 (N_8468,N_5662,N_3879);
nand U8469 (N_8469,N_3410,N_4125);
and U8470 (N_8470,N_4863,N_5105);
or U8471 (N_8471,N_3976,N_4680);
xor U8472 (N_8472,N_4256,N_5605);
and U8473 (N_8473,N_5670,N_3474);
nor U8474 (N_8474,N_4095,N_4471);
and U8475 (N_8475,N_3014,N_5446);
or U8476 (N_8476,N_4859,N_3138);
nand U8477 (N_8477,N_4699,N_5318);
nor U8478 (N_8478,N_4842,N_4321);
nand U8479 (N_8479,N_5507,N_4291);
or U8480 (N_8480,N_4684,N_4839);
or U8481 (N_8481,N_3269,N_3467);
nand U8482 (N_8482,N_3850,N_5763);
nand U8483 (N_8483,N_3813,N_3138);
and U8484 (N_8484,N_3645,N_3586);
nand U8485 (N_8485,N_5741,N_5344);
nand U8486 (N_8486,N_4913,N_3740);
and U8487 (N_8487,N_5160,N_5116);
or U8488 (N_8488,N_5824,N_4431);
and U8489 (N_8489,N_4963,N_3617);
nand U8490 (N_8490,N_4904,N_3098);
xor U8491 (N_8491,N_3316,N_4133);
nand U8492 (N_8492,N_5365,N_3600);
and U8493 (N_8493,N_3306,N_4651);
nand U8494 (N_8494,N_4540,N_5991);
nor U8495 (N_8495,N_4423,N_4767);
and U8496 (N_8496,N_5182,N_5344);
xnor U8497 (N_8497,N_5497,N_3399);
or U8498 (N_8498,N_4247,N_4335);
nand U8499 (N_8499,N_4004,N_4628);
or U8500 (N_8500,N_5345,N_4748);
xor U8501 (N_8501,N_3930,N_3337);
nor U8502 (N_8502,N_4111,N_4904);
or U8503 (N_8503,N_4002,N_4749);
or U8504 (N_8504,N_5329,N_3420);
or U8505 (N_8505,N_5366,N_3312);
and U8506 (N_8506,N_3213,N_5342);
or U8507 (N_8507,N_4092,N_5689);
and U8508 (N_8508,N_3324,N_4528);
xnor U8509 (N_8509,N_5951,N_4661);
nand U8510 (N_8510,N_5029,N_4581);
and U8511 (N_8511,N_3902,N_5183);
and U8512 (N_8512,N_3375,N_3125);
and U8513 (N_8513,N_3173,N_4204);
nor U8514 (N_8514,N_3813,N_4145);
and U8515 (N_8515,N_4519,N_5667);
nor U8516 (N_8516,N_4059,N_5029);
nor U8517 (N_8517,N_3060,N_5374);
nand U8518 (N_8518,N_4078,N_4315);
nand U8519 (N_8519,N_5812,N_3278);
and U8520 (N_8520,N_3703,N_3208);
xnor U8521 (N_8521,N_4668,N_3637);
and U8522 (N_8522,N_3281,N_5100);
nand U8523 (N_8523,N_5867,N_4536);
and U8524 (N_8524,N_4781,N_5453);
or U8525 (N_8525,N_4957,N_5713);
or U8526 (N_8526,N_5563,N_4583);
or U8527 (N_8527,N_3416,N_3244);
nand U8528 (N_8528,N_4191,N_4453);
nor U8529 (N_8529,N_4180,N_4464);
nand U8530 (N_8530,N_4171,N_3527);
nor U8531 (N_8531,N_5678,N_4752);
xor U8532 (N_8532,N_5179,N_5976);
nor U8533 (N_8533,N_4275,N_4257);
or U8534 (N_8534,N_3081,N_5506);
and U8535 (N_8535,N_5775,N_3410);
nor U8536 (N_8536,N_5352,N_5117);
or U8537 (N_8537,N_5006,N_3940);
nand U8538 (N_8538,N_3406,N_3196);
or U8539 (N_8539,N_4047,N_4556);
or U8540 (N_8540,N_4665,N_4036);
and U8541 (N_8541,N_3715,N_4386);
nand U8542 (N_8542,N_5646,N_3581);
nor U8543 (N_8543,N_5093,N_4451);
nand U8544 (N_8544,N_5846,N_5702);
or U8545 (N_8545,N_3038,N_3903);
nor U8546 (N_8546,N_5918,N_5740);
nor U8547 (N_8547,N_5161,N_4120);
and U8548 (N_8548,N_3769,N_4143);
and U8549 (N_8549,N_5174,N_3816);
nand U8550 (N_8550,N_4174,N_4591);
nor U8551 (N_8551,N_3109,N_5211);
and U8552 (N_8552,N_4330,N_5678);
or U8553 (N_8553,N_3126,N_5196);
nor U8554 (N_8554,N_5152,N_4191);
nand U8555 (N_8555,N_3485,N_3604);
nand U8556 (N_8556,N_4821,N_4296);
or U8557 (N_8557,N_3461,N_5805);
nand U8558 (N_8558,N_5920,N_3618);
or U8559 (N_8559,N_5729,N_5288);
nand U8560 (N_8560,N_5784,N_4221);
and U8561 (N_8561,N_4848,N_3205);
and U8562 (N_8562,N_5128,N_5839);
nand U8563 (N_8563,N_4072,N_3644);
nand U8564 (N_8564,N_5645,N_5444);
and U8565 (N_8565,N_3884,N_5024);
and U8566 (N_8566,N_4896,N_4599);
and U8567 (N_8567,N_3467,N_3387);
or U8568 (N_8568,N_3832,N_3803);
and U8569 (N_8569,N_4705,N_4657);
or U8570 (N_8570,N_3211,N_3617);
or U8571 (N_8571,N_3532,N_5746);
and U8572 (N_8572,N_4199,N_5736);
or U8573 (N_8573,N_5157,N_3878);
nand U8574 (N_8574,N_3833,N_5530);
nand U8575 (N_8575,N_3127,N_3077);
or U8576 (N_8576,N_3321,N_3493);
or U8577 (N_8577,N_5434,N_3892);
nor U8578 (N_8578,N_5978,N_4705);
and U8579 (N_8579,N_5616,N_4914);
nor U8580 (N_8580,N_3061,N_4989);
or U8581 (N_8581,N_4011,N_5505);
nand U8582 (N_8582,N_4223,N_3487);
nor U8583 (N_8583,N_4997,N_4582);
nor U8584 (N_8584,N_5876,N_4102);
xnor U8585 (N_8585,N_5569,N_5286);
or U8586 (N_8586,N_3662,N_3587);
and U8587 (N_8587,N_4942,N_5288);
and U8588 (N_8588,N_4488,N_3290);
and U8589 (N_8589,N_3884,N_3544);
and U8590 (N_8590,N_5866,N_4940);
and U8591 (N_8591,N_3814,N_3350);
or U8592 (N_8592,N_4946,N_5292);
and U8593 (N_8593,N_3097,N_4206);
nand U8594 (N_8594,N_4797,N_4068);
or U8595 (N_8595,N_3640,N_4065);
nand U8596 (N_8596,N_4748,N_3878);
or U8597 (N_8597,N_4924,N_4805);
or U8598 (N_8598,N_3637,N_5608);
and U8599 (N_8599,N_4863,N_3511);
nor U8600 (N_8600,N_5316,N_4913);
and U8601 (N_8601,N_5099,N_4046);
nor U8602 (N_8602,N_4912,N_5640);
nand U8603 (N_8603,N_4997,N_4552);
and U8604 (N_8604,N_3341,N_5737);
xnor U8605 (N_8605,N_5840,N_3079);
nand U8606 (N_8606,N_4538,N_3761);
and U8607 (N_8607,N_3623,N_5811);
nand U8608 (N_8608,N_4796,N_3613);
xnor U8609 (N_8609,N_5712,N_4239);
or U8610 (N_8610,N_4515,N_4003);
and U8611 (N_8611,N_4787,N_5609);
nand U8612 (N_8612,N_4018,N_3582);
or U8613 (N_8613,N_3121,N_5188);
or U8614 (N_8614,N_5674,N_5423);
and U8615 (N_8615,N_3282,N_4452);
nand U8616 (N_8616,N_5361,N_5023);
and U8617 (N_8617,N_5117,N_4291);
or U8618 (N_8618,N_4769,N_3541);
and U8619 (N_8619,N_3336,N_4060);
nor U8620 (N_8620,N_5787,N_5141);
nand U8621 (N_8621,N_4402,N_3366);
nand U8622 (N_8622,N_4827,N_5730);
and U8623 (N_8623,N_4958,N_5507);
and U8624 (N_8624,N_5465,N_5933);
nor U8625 (N_8625,N_3251,N_3347);
nor U8626 (N_8626,N_3462,N_3768);
and U8627 (N_8627,N_3649,N_4626);
nor U8628 (N_8628,N_3128,N_4187);
or U8629 (N_8629,N_4882,N_3768);
nand U8630 (N_8630,N_4801,N_3504);
nor U8631 (N_8631,N_3945,N_4866);
nor U8632 (N_8632,N_5075,N_4896);
nand U8633 (N_8633,N_5822,N_5863);
or U8634 (N_8634,N_4635,N_5512);
nor U8635 (N_8635,N_5719,N_5366);
and U8636 (N_8636,N_3340,N_3035);
or U8637 (N_8637,N_4311,N_4661);
nand U8638 (N_8638,N_4840,N_4442);
nor U8639 (N_8639,N_3916,N_4685);
nand U8640 (N_8640,N_3722,N_5984);
and U8641 (N_8641,N_4279,N_4985);
nor U8642 (N_8642,N_5136,N_5246);
and U8643 (N_8643,N_3599,N_3113);
and U8644 (N_8644,N_5068,N_5005);
nor U8645 (N_8645,N_5930,N_4782);
nand U8646 (N_8646,N_5983,N_3700);
nor U8647 (N_8647,N_4929,N_5093);
nor U8648 (N_8648,N_3720,N_5430);
or U8649 (N_8649,N_4672,N_5634);
nand U8650 (N_8650,N_5116,N_3175);
nor U8651 (N_8651,N_5360,N_5819);
and U8652 (N_8652,N_3609,N_3911);
nand U8653 (N_8653,N_4348,N_4742);
nor U8654 (N_8654,N_5160,N_3429);
xor U8655 (N_8655,N_5429,N_4295);
and U8656 (N_8656,N_4628,N_4778);
or U8657 (N_8657,N_3196,N_5014);
and U8658 (N_8658,N_4503,N_3289);
nor U8659 (N_8659,N_3202,N_5759);
or U8660 (N_8660,N_5888,N_3146);
nand U8661 (N_8661,N_4129,N_4196);
and U8662 (N_8662,N_5678,N_5512);
and U8663 (N_8663,N_4531,N_4279);
nand U8664 (N_8664,N_3246,N_4445);
and U8665 (N_8665,N_3872,N_4383);
or U8666 (N_8666,N_3582,N_3362);
or U8667 (N_8667,N_3934,N_4803);
nor U8668 (N_8668,N_3492,N_3550);
or U8669 (N_8669,N_3790,N_5569);
or U8670 (N_8670,N_4079,N_3845);
nand U8671 (N_8671,N_5475,N_3360);
nor U8672 (N_8672,N_5339,N_3189);
and U8673 (N_8673,N_3974,N_5660);
nor U8674 (N_8674,N_3822,N_5457);
nor U8675 (N_8675,N_3846,N_5254);
xnor U8676 (N_8676,N_3392,N_5336);
and U8677 (N_8677,N_3178,N_3081);
nor U8678 (N_8678,N_4580,N_5989);
nand U8679 (N_8679,N_5473,N_5757);
nor U8680 (N_8680,N_5809,N_5247);
nand U8681 (N_8681,N_5145,N_5208);
nor U8682 (N_8682,N_3973,N_5026);
nand U8683 (N_8683,N_3514,N_5484);
or U8684 (N_8684,N_3149,N_5418);
xnor U8685 (N_8685,N_3551,N_4998);
and U8686 (N_8686,N_5266,N_5217);
or U8687 (N_8687,N_4053,N_4005);
xnor U8688 (N_8688,N_4352,N_4220);
nor U8689 (N_8689,N_5385,N_5692);
or U8690 (N_8690,N_3487,N_4715);
nor U8691 (N_8691,N_5438,N_4342);
or U8692 (N_8692,N_3162,N_3835);
nor U8693 (N_8693,N_3042,N_5874);
or U8694 (N_8694,N_5473,N_4260);
xor U8695 (N_8695,N_5711,N_3596);
nand U8696 (N_8696,N_5126,N_4481);
xnor U8697 (N_8697,N_5854,N_4652);
or U8698 (N_8698,N_5450,N_5475);
nand U8699 (N_8699,N_5447,N_4614);
or U8700 (N_8700,N_4300,N_4760);
or U8701 (N_8701,N_5452,N_3205);
and U8702 (N_8702,N_5866,N_3874);
nand U8703 (N_8703,N_4376,N_4937);
xor U8704 (N_8704,N_3270,N_3369);
nand U8705 (N_8705,N_5908,N_4820);
nand U8706 (N_8706,N_4252,N_4141);
or U8707 (N_8707,N_3234,N_5893);
and U8708 (N_8708,N_3883,N_5209);
nand U8709 (N_8709,N_4211,N_4422);
and U8710 (N_8710,N_5257,N_5396);
and U8711 (N_8711,N_3285,N_3317);
nand U8712 (N_8712,N_5139,N_5615);
xor U8713 (N_8713,N_3038,N_3271);
or U8714 (N_8714,N_3727,N_5840);
nor U8715 (N_8715,N_4778,N_3574);
or U8716 (N_8716,N_3700,N_5196);
or U8717 (N_8717,N_5688,N_4504);
nor U8718 (N_8718,N_5146,N_4650);
xor U8719 (N_8719,N_4972,N_4945);
nand U8720 (N_8720,N_5359,N_5624);
and U8721 (N_8721,N_4607,N_4928);
or U8722 (N_8722,N_3427,N_5795);
or U8723 (N_8723,N_3824,N_4747);
or U8724 (N_8724,N_5536,N_5868);
or U8725 (N_8725,N_4004,N_5573);
nand U8726 (N_8726,N_3485,N_4846);
and U8727 (N_8727,N_5451,N_3250);
xor U8728 (N_8728,N_5436,N_3540);
nor U8729 (N_8729,N_3110,N_5147);
nand U8730 (N_8730,N_4179,N_3466);
or U8731 (N_8731,N_5412,N_3955);
and U8732 (N_8732,N_3991,N_5207);
and U8733 (N_8733,N_3096,N_5116);
or U8734 (N_8734,N_5002,N_4725);
nor U8735 (N_8735,N_3891,N_3575);
and U8736 (N_8736,N_4365,N_3661);
and U8737 (N_8737,N_5037,N_4367);
nand U8738 (N_8738,N_5206,N_3900);
and U8739 (N_8739,N_5945,N_3938);
nand U8740 (N_8740,N_4803,N_4110);
nor U8741 (N_8741,N_4723,N_4292);
nand U8742 (N_8742,N_3547,N_5263);
or U8743 (N_8743,N_3852,N_5201);
or U8744 (N_8744,N_3101,N_3072);
nand U8745 (N_8745,N_4866,N_3095);
nor U8746 (N_8746,N_3014,N_4108);
xnor U8747 (N_8747,N_5089,N_4129);
and U8748 (N_8748,N_4818,N_5626);
nor U8749 (N_8749,N_3740,N_4141);
and U8750 (N_8750,N_3675,N_5075);
or U8751 (N_8751,N_4835,N_5889);
or U8752 (N_8752,N_4595,N_5120);
nand U8753 (N_8753,N_5187,N_3980);
or U8754 (N_8754,N_3336,N_4863);
xnor U8755 (N_8755,N_5380,N_5502);
or U8756 (N_8756,N_4960,N_3873);
nand U8757 (N_8757,N_4671,N_5998);
nand U8758 (N_8758,N_5614,N_3125);
nor U8759 (N_8759,N_3276,N_4129);
or U8760 (N_8760,N_4589,N_3255);
and U8761 (N_8761,N_5939,N_3823);
nand U8762 (N_8762,N_4202,N_5899);
nor U8763 (N_8763,N_4989,N_4277);
xnor U8764 (N_8764,N_4150,N_3752);
nand U8765 (N_8765,N_5521,N_5899);
nand U8766 (N_8766,N_4635,N_4162);
xnor U8767 (N_8767,N_5553,N_3923);
or U8768 (N_8768,N_5102,N_3656);
and U8769 (N_8769,N_4498,N_4749);
and U8770 (N_8770,N_4486,N_3651);
xnor U8771 (N_8771,N_3005,N_3521);
and U8772 (N_8772,N_3344,N_4257);
nor U8773 (N_8773,N_4998,N_3062);
and U8774 (N_8774,N_3025,N_4118);
nor U8775 (N_8775,N_5425,N_4950);
and U8776 (N_8776,N_5088,N_3327);
nor U8777 (N_8777,N_3245,N_5851);
or U8778 (N_8778,N_5305,N_3969);
xnor U8779 (N_8779,N_4685,N_5065);
xnor U8780 (N_8780,N_4466,N_3548);
nor U8781 (N_8781,N_4022,N_5119);
nand U8782 (N_8782,N_4723,N_3934);
nand U8783 (N_8783,N_3359,N_3389);
nor U8784 (N_8784,N_4991,N_5058);
nand U8785 (N_8785,N_4524,N_3925);
nand U8786 (N_8786,N_3534,N_5015);
xor U8787 (N_8787,N_4367,N_3519);
nand U8788 (N_8788,N_4986,N_3797);
nor U8789 (N_8789,N_3259,N_4414);
or U8790 (N_8790,N_5990,N_5437);
nor U8791 (N_8791,N_4686,N_3978);
and U8792 (N_8792,N_4486,N_5238);
nand U8793 (N_8793,N_4120,N_4270);
and U8794 (N_8794,N_5589,N_5962);
or U8795 (N_8795,N_4223,N_3360);
or U8796 (N_8796,N_5719,N_4355);
xor U8797 (N_8797,N_4263,N_4181);
nor U8798 (N_8798,N_3754,N_3279);
and U8799 (N_8799,N_5195,N_3984);
xor U8800 (N_8800,N_3466,N_5855);
nand U8801 (N_8801,N_3030,N_4254);
nand U8802 (N_8802,N_3486,N_5123);
nor U8803 (N_8803,N_5635,N_4061);
xor U8804 (N_8804,N_3140,N_5165);
nand U8805 (N_8805,N_4731,N_3777);
and U8806 (N_8806,N_4449,N_5247);
or U8807 (N_8807,N_4320,N_4019);
nand U8808 (N_8808,N_3410,N_4352);
and U8809 (N_8809,N_5857,N_4339);
nand U8810 (N_8810,N_4428,N_5608);
or U8811 (N_8811,N_4479,N_3298);
nand U8812 (N_8812,N_3488,N_5446);
and U8813 (N_8813,N_4017,N_4344);
nand U8814 (N_8814,N_5211,N_4615);
nor U8815 (N_8815,N_4457,N_5045);
and U8816 (N_8816,N_4665,N_3165);
or U8817 (N_8817,N_3957,N_3661);
nor U8818 (N_8818,N_5841,N_4754);
or U8819 (N_8819,N_4399,N_4050);
or U8820 (N_8820,N_4875,N_4067);
nor U8821 (N_8821,N_5073,N_5535);
and U8822 (N_8822,N_3168,N_5608);
nand U8823 (N_8823,N_4735,N_5576);
nand U8824 (N_8824,N_5704,N_4748);
or U8825 (N_8825,N_3832,N_3504);
and U8826 (N_8826,N_5871,N_3778);
xnor U8827 (N_8827,N_3530,N_5551);
xor U8828 (N_8828,N_4580,N_5275);
and U8829 (N_8829,N_3604,N_5562);
and U8830 (N_8830,N_3304,N_3687);
or U8831 (N_8831,N_5757,N_4898);
nand U8832 (N_8832,N_4132,N_4443);
nand U8833 (N_8833,N_5067,N_5563);
or U8834 (N_8834,N_4816,N_4355);
or U8835 (N_8835,N_4756,N_5430);
or U8836 (N_8836,N_3973,N_4062);
and U8837 (N_8837,N_4884,N_5631);
or U8838 (N_8838,N_4962,N_5836);
xnor U8839 (N_8839,N_3441,N_4155);
nor U8840 (N_8840,N_4830,N_5279);
nor U8841 (N_8841,N_5777,N_5430);
or U8842 (N_8842,N_5136,N_4574);
nand U8843 (N_8843,N_5997,N_3340);
or U8844 (N_8844,N_5276,N_3560);
or U8845 (N_8845,N_4177,N_3535);
nor U8846 (N_8846,N_3262,N_3668);
nand U8847 (N_8847,N_5966,N_3987);
nor U8848 (N_8848,N_5575,N_4441);
or U8849 (N_8849,N_5159,N_4478);
and U8850 (N_8850,N_3759,N_3831);
nor U8851 (N_8851,N_3565,N_5386);
xor U8852 (N_8852,N_4951,N_3608);
xnor U8853 (N_8853,N_3961,N_3534);
nor U8854 (N_8854,N_3910,N_3354);
nor U8855 (N_8855,N_3030,N_4279);
nand U8856 (N_8856,N_5820,N_5480);
nand U8857 (N_8857,N_3174,N_5625);
or U8858 (N_8858,N_3375,N_5338);
nand U8859 (N_8859,N_4654,N_4638);
and U8860 (N_8860,N_5678,N_5867);
xnor U8861 (N_8861,N_5898,N_3560);
or U8862 (N_8862,N_4173,N_4532);
nor U8863 (N_8863,N_3916,N_5316);
nand U8864 (N_8864,N_4966,N_3911);
xnor U8865 (N_8865,N_5361,N_5094);
nor U8866 (N_8866,N_5174,N_5497);
or U8867 (N_8867,N_5695,N_5974);
and U8868 (N_8868,N_5477,N_4282);
or U8869 (N_8869,N_3584,N_3075);
and U8870 (N_8870,N_5904,N_5398);
nor U8871 (N_8871,N_4743,N_3388);
nand U8872 (N_8872,N_3536,N_5152);
or U8873 (N_8873,N_5705,N_4356);
or U8874 (N_8874,N_5036,N_3169);
or U8875 (N_8875,N_4593,N_4926);
and U8876 (N_8876,N_5958,N_5092);
and U8877 (N_8877,N_3601,N_4307);
or U8878 (N_8878,N_4277,N_4516);
and U8879 (N_8879,N_4041,N_3986);
or U8880 (N_8880,N_4136,N_3879);
and U8881 (N_8881,N_4391,N_5369);
and U8882 (N_8882,N_3195,N_3066);
and U8883 (N_8883,N_3123,N_3284);
and U8884 (N_8884,N_4378,N_3928);
or U8885 (N_8885,N_3444,N_5377);
and U8886 (N_8886,N_5906,N_4902);
or U8887 (N_8887,N_4258,N_5876);
nand U8888 (N_8888,N_3809,N_3173);
xnor U8889 (N_8889,N_5167,N_4410);
xor U8890 (N_8890,N_3073,N_5291);
nand U8891 (N_8891,N_5714,N_3308);
or U8892 (N_8892,N_4665,N_4295);
or U8893 (N_8893,N_4377,N_3431);
nand U8894 (N_8894,N_3727,N_5348);
or U8895 (N_8895,N_5492,N_4169);
or U8896 (N_8896,N_3014,N_4895);
nand U8897 (N_8897,N_3393,N_3799);
xnor U8898 (N_8898,N_3032,N_3885);
nand U8899 (N_8899,N_5389,N_3981);
and U8900 (N_8900,N_5587,N_4160);
and U8901 (N_8901,N_3127,N_4720);
and U8902 (N_8902,N_4459,N_3878);
or U8903 (N_8903,N_4035,N_4225);
nand U8904 (N_8904,N_4393,N_4776);
and U8905 (N_8905,N_4945,N_5265);
nor U8906 (N_8906,N_5777,N_5991);
nor U8907 (N_8907,N_3691,N_4706);
nand U8908 (N_8908,N_5341,N_3205);
nor U8909 (N_8909,N_5672,N_3471);
or U8910 (N_8910,N_4519,N_3748);
or U8911 (N_8911,N_3625,N_4646);
or U8912 (N_8912,N_4333,N_4047);
and U8913 (N_8913,N_3788,N_3760);
xnor U8914 (N_8914,N_4559,N_4013);
xnor U8915 (N_8915,N_3629,N_5193);
or U8916 (N_8916,N_4900,N_3275);
nor U8917 (N_8917,N_5789,N_3530);
nor U8918 (N_8918,N_4075,N_4405);
and U8919 (N_8919,N_4502,N_3071);
or U8920 (N_8920,N_3684,N_3419);
nor U8921 (N_8921,N_3117,N_5952);
and U8922 (N_8922,N_4339,N_4315);
xnor U8923 (N_8923,N_5221,N_5054);
or U8924 (N_8924,N_3198,N_3557);
or U8925 (N_8925,N_4006,N_4024);
nand U8926 (N_8926,N_4297,N_5494);
and U8927 (N_8927,N_4899,N_4902);
nand U8928 (N_8928,N_4605,N_5668);
and U8929 (N_8929,N_3198,N_4984);
nand U8930 (N_8930,N_3849,N_5652);
and U8931 (N_8931,N_3706,N_4695);
or U8932 (N_8932,N_4677,N_4388);
and U8933 (N_8933,N_5344,N_4984);
nor U8934 (N_8934,N_5292,N_5503);
nand U8935 (N_8935,N_5955,N_5209);
and U8936 (N_8936,N_5915,N_5087);
and U8937 (N_8937,N_3631,N_5620);
nor U8938 (N_8938,N_5934,N_5451);
and U8939 (N_8939,N_5267,N_3461);
and U8940 (N_8940,N_3594,N_5856);
and U8941 (N_8941,N_4152,N_4345);
nand U8942 (N_8942,N_5658,N_4156);
or U8943 (N_8943,N_4236,N_4301);
or U8944 (N_8944,N_3069,N_3835);
nand U8945 (N_8945,N_3506,N_5832);
or U8946 (N_8946,N_4910,N_4499);
nand U8947 (N_8947,N_3452,N_4906);
or U8948 (N_8948,N_5138,N_3151);
and U8949 (N_8949,N_3633,N_5863);
or U8950 (N_8950,N_5958,N_4246);
nand U8951 (N_8951,N_4730,N_5117);
nor U8952 (N_8952,N_5857,N_5878);
or U8953 (N_8953,N_4588,N_3068);
or U8954 (N_8954,N_4892,N_4540);
or U8955 (N_8955,N_5244,N_5819);
nand U8956 (N_8956,N_4973,N_5761);
nand U8957 (N_8957,N_3561,N_5902);
nor U8958 (N_8958,N_3324,N_4689);
nand U8959 (N_8959,N_3215,N_4957);
or U8960 (N_8960,N_4174,N_5478);
or U8961 (N_8961,N_5349,N_4995);
nand U8962 (N_8962,N_4103,N_3694);
nor U8963 (N_8963,N_5392,N_5382);
or U8964 (N_8964,N_5115,N_3442);
and U8965 (N_8965,N_3644,N_3485);
nand U8966 (N_8966,N_3916,N_5463);
or U8967 (N_8967,N_3814,N_4093);
nor U8968 (N_8968,N_3674,N_5134);
or U8969 (N_8969,N_4090,N_4343);
and U8970 (N_8970,N_3796,N_3703);
nor U8971 (N_8971,N_4982,N_5793);
nand U8972 (N_8972,N_4323,N_3565);
nand U8973 (N_8973,N_4867,N_4733);
nand U8974 (N_8974,N_3865,N_3265);
nand U8975 (N_8975,N_4638,N_5492);
and U8976 (N_8976,N_4095,N_4592);
nand U8977 (N_8977,N_3697,N_5515);
nor U8978 (N_8978,N_5795,N_4945);
nand U8979 (N_8979,N_5414,N_3260);
nor U8980 (N_8980,N_3816,N_5087);
nand U8981 (N_8981,N_4586,N_3724);
and U8982 (N_8982,N_4563,N_5230);
or U8983 (N_8983,N_4452,N_5969);
or U8984 (N_8984,N_3055,N_3259);
or U8985 (N_8985,N_4971,N_4133);
nand U8986 (N_8986,N_5240,N_5183);
xor U8987 (N_8987,N_3110,N_4540);
and U8988 (N_8988,N_5645,N_3854);
and U8989 (N_8989,N_4650,N_3060);
nand U8990 (N_8990,N_4267,N_5425);
nor U8991 (N_8991,N_4434,N_3134);
or U8992 (N_8992,N_3724,N_3524);
xnor U8993 (N_8993,N_5776,N_5098);
and U8994 (N_8994,N_3057,N_4044);
and U8995 (N_8995,N_5693,N_5352);
nor U8996 (N_8996,N_3915,N_3587);
and U8997 (N_8997,N_3995,N_4766);
or U8998 (N_8998,N_5622,N_3334);
nor U8999 (N_8999,N_3945,N_3493);
or U9000 (N_9000,N_7229,N_8747);
nand U9001 (N_9001,N_6685,N_7687);
nand U9002 (N_9002,N_8820,N_8178);
and U9003 (N_9003,N_8794,N_6402);
nor U9004 (N_9004,N_7216,N_6470);
nand U9005 (N_9005,N_7039,N_7208);
and U9006 (N_9006,N_6842,N_7425);
xnor U9007 (N_9007,N_8310,N_7830);
xnor U9008 (N_9008,N_6110,N_8826);
or U9009 (N_9009,N_7214,N_6741);
xor U9010 (N_9010,N_8144,N_6139);
nor U9011 (N_9011,N_6515,N_7044);
or U9012 (N_9012,N_8743,N_7218);
nor U9013 (N_9013,N_7041,N_8807);
nand U9014 (N_9014,N_6076,N_7672);
and U9015 (N_9015,N_8946,N_6424);
nand U9016 (N_9016,N_8362,N_6814);
nor U9017 (N_9017,N_6581,N_8082);
nand U9018 (N_9018,N_8625,N_6479);
nand U9019 (N_9019,N_7501,N_8890);
and U9020 (N_9020,N_8430,N_8524);
nor U9021 (N_9021,N_7077,N_6882);
nand U9022 (N_9022,N_8428,N_6995);
nor U9023 (N_9023,N_6486,N_6901);
and U9024 (N_9024,N_6699,N_8356);
nor U9025 (N_9025,N_8843,N_6019);
or U9026 (N_9026,N_6744,N_8357);
and U9027 (N_9027,N_6442,N_7226);
nand U9028 (N_9028,N_6282,N_6360);
nor U9029 (N_9029,N_6841,N_7976);
nand U9030 (N_9030,N_6129,N_7197);
xor U9031 (N_9031,N_8053,N_8241);
nand U9032 (N_9032,N_6449,N_8790);
nor U9033 (N_9033,N_7099,N_8891);
and U9034 (N_9034,N_8019,N_6326);
xnor U9035 (N_9035,N_8847,N_7401);
or U9036 (N_9036,N_8793,N_8086);
xnor U9037 (N_9037,N_7428,N_8018);
nand U9038 (N_9038,N_7122,N_8186);
nand U9039 (N_9039,N_8766,N_8569);
or U9040 (N_9040,N_7967,N_8746);
or U9041 (N_9041,N_7613,N_6607);
or U9042 (N_9042,N_6567,N_7343);
nand U9043 (N_9043,N_8094,N_8051);
nand U9044 (N_9044,N_8325,N_7492);
and U9045 (N_9045,N_8870,N_7811);
nor U9046 (N_9046,N_8596,N_7138);
nand U9047 (N_9047,N_8618,N_8912);
nor U9048 (N_9048,N_6527,N_7600);
or U9049 (N_9049,N_7498,N_8373);
and U9050 (N_9050,N_6105,N_7421);
or U9051 (N_9051,N_6312,N_6565);
nand U9052 (N_9052,N_6276,N_8267);
and U9053 (N_9053,N_7506,N_6650);
or U9054 (N_9054,N_6031,N_8426);
nand U9055 (N_9055,N_6109,N_8063);
or U9056 (N_9056,N_8553,N_7992);
and U9057 (N_9057,N_7786,N_8175);
and U9058 (N_9058,N_6697,N_7043);
nand U9059 (N_9059,N_7815,N_6965);
nand U9060 (N_9060,N_7544,N_7223);
and U9061 (N_9061,N_8117,N_7693);
nor U9062 (N_9062,N_8719,N_8903);
nor U9063 (N_9063,N_7283,N_6497);
or U9064 (N_9064,N_7433,N_6473);
nand U9065 (N_9065,N_6827,N_6016);
or U9066 (N_9066,N_7861,N_8473);
and U9067 (N_9067,N_6376,N_7130);
xor U9068 (N_9068,N_7233,N_6906);
and U9069 (N_9069,N_8346,N_6379);
and U9070 (N_9070,N_8106,N_6730);
nor U9071 (N_9071,N_7256,N_8209);
and U9072 (N_9072,N_6093,N_6400);
or U9073 (N_9073,N_8338,N_8978);
and U9074 (N_9074,N_7641,N_7125);
nor U9075 (N_9075,N_7705,N_7002);
or U9076 (N_9076,N_7007,N_6026);
or U9077 (N_9077,N_7995,N_7943);
and U9078 (N_9078,N_6696,N_7543);
nand U9079 (N_9079,N_6949,N_6340);
and U9080 (N_9080,N_7537,N_6427);
nor U9081 (N_9081,N_8301,N_8035);
nand U9082 (N_9082,N_6252,N_8855);
or U9083 (N_9083,N_8535,N_8353);
xnor U9084 (N_9084,N_7795,N_6406);
nand U9085 (N_9085,N_7953,N_6418);
nand U9086 (N_9086,N_6186,N_6417);
or U9087 (N_9087,N_8312,N_6434);
nand U9088 (N_9088,N_6571,N_7610);
nand U9089 (N_9089,N_7594,N_6444);
or U9090 (N_9090,N_6035,N_6051);
or U9091 (N_9091,N_8690,N_7586);
or U9092 (N_9092,N_8940,N_6726);
and U9093 (N_9093,N_7465,N_6315);
and U9094 (N_9094,N_7652,N_7602);
xor U9095 (N_9095,N_7514,N_7758);
xnor U9096 (N_9096,N_7154,N_7726);
nor U9097 (N_9097,N_7413,N_7450);
and U9098 (N_9098,N_7496,N_6222);
nand U9099 (N_9099,N_7087,N_7552);
nor U9100 (N_9100,N_6407,N_7904);
and U9101 (N_9101,N_8152,N_7669);
or U9102 (N_9102,N_6301,N_6560);
nand U9103 (N_9103,N_7018,N_8273);
nor U9104 (N_9104,N_7101,N_6500);
and U9105 (N_9105,N_7117,N_8497);
nor U9106 (N_9106,N_7377,N_8114);
nand U9107 (N_9107,N_8882,N_8172);
or U9108 (N_9108,N_6523,N_8953);
or U9109 (N_9109,N_7707,N_7050);
nand U9110 (N_9110,N_7667,N_7031);
nor U9111 (N_9111,N_7604,N_7710);
and U9112 (N_9112,N_7239,N_7589);
nor U9113 (N_9113,N_6982,N_7362);
nor U9114 (N_9114,N_7615,N_8115);
nand U9115 (N_9115,N_7032,N_7668);
nor U9116 (N_9116,N_6123,N_6126);
or U9117 (N_9117,N_8071,N_6707);
and U9118 (N_9118,N_8307,N_8588);
nor U9119 (N_9119,N_8097,N_6154);
nand U9120 (N_9120,N_6671,N_8374);
or U9121 (N_9121,N_7415,N_8213);
nand U9122 (N_9122,N_8955,N_6270);
or U9123 (N_9123,N_7777,N_8815);
or U9124 (N_9124,N_7158,N_8600);
xnor U9125 (N_9125,N_6217,N_7079);
and U9126 (N_9126,N_7434,N_8122);
or U9127 (N_9127,N_7633,N_6094);
or U9128 (N_9128,N_8958,N_7689);
nand U9129 (N_9129,N_8701,N_7700);
and U9130 (N_9130,N_8523,N_8449);
or U9131 (N_9131,N_8693,N_6150);
or U9132 (N_9132,N_6724,N_8350);
or U9133 (N_9133,N_8567,N_7398);
and U9134 (N_9134,N_6463,N_7728);
nor U9135 (N_9135,N_6902,N_6678);
xor U9136 (N_9136,N_6302,N_8381);
or U9137 (N_9137,N_8004,N_7460);
xnor U9138 (N_9138,N_8399,N_6169);
and U9139 (N_9139,N_6398,N_8272);
nand U9140 (N_9140,N_7166,N_8914);
nand U9141 (N_9141,N_8661,N_8101);
nand U9142 (N_9142,N_7753,N_6433);
and U9143 (N_9143,N_8964,N_8364);
nor U9144 (N_9144,N_7356,N_8664);
nand U9145 (N_9145,N_8037,N_7912);
xor U9146 (N_9146,N_8601,N_7269);
and U9147 (N_9147,N_8005,N_8187);
and U9148 (N_9148,N_6192,N_7408);
and U9149 (N_9149,N_7301,N_6632);
xor U9150 (N_9150,N_8983,N_8311);
nand U9151 (N_9151,N_7782,N_6388);
or U9152 (N_9152,N_6119,N_6522);
or U9153 (N_9153,N_6610,N_7476);
or U9154 (N_9154,N_6365,N_7140);
nor U9155 (N_9155,N_8634,N_7332);
xor U9156 (N_9156,N_6116,N_7987);
xnor U9157 (N_9157,N_6494,N_7368);
nor U9158 (N_9158,N_6140,N_8676);
nor U9159 (N_9159,N_6163,N_8192);
and U9160 (N_9160,N_8735,N_7989);
and U9161 (N_9161,N_7837,N_6245);
and U9162 (N_9162,N_6847,N_7380);
and U9163 (N_9163,N_6448,N_8788);
nand U9164 (N_9164,N_7027,N_8653);
nand U9165 (N_9165,N_6115,N_8015);
nor U9166 (N_9166,N_8467,N_8910);
and U9167 (N_9167,N_8243,N_6719);
nand U9168 (N_9168,N_6443,N_8442);
or U9169 (N_9169,N_7581,N_7255);
nor U9170 (N_9170,N_6553,N_6499);
xor U9171 (N_9171,N_8262,N_8576);
nor U9172 (N_9172,N_6863,N_7926);
nor U9173 (N_9173,N_7824,N_7149);
and U9174 (N_9174,N_7504,N_7677);
or U9175 (N_9175,N_8002,N_8230);
or U9176 (N_9176,N_6808,N_7232);
or U9177 (N_9177,N_8227,N_6209);
and U9178 (N_9178,N_7126,N_8704);
and U9179 (N_9179,N_8103,N_8879);
nand U9180 (N_9180,N_7509,N_8096);
and U9181 (N_9181,N_7371,N_6042);
nor U9182 (N_9182,N_8067,N_7467);
and U9183 (N_9183,N_7073,N_8223);
or U9184 (N_9184,N_8972,N_8681);
nand U9185 (N_9185,N_8039,N_8771);
and U9186 (N_9186,N_6839,N_7253);
xnor U9187 (N_9187,N_6914,N_7142);
xnor U9188 (N_9188,N_6175,N_7175);
nand U9189 (N_9189,N_6688,N_8594);
nor U9190 (N_9190,N_7135,N_8516);
nand U9191 (N_9191,N_6904,N_6011);
nor U9192 (N_9192,N_8974,N_8684);
and U9193 (N_9193,N_7858,N_8526);
and U9194 (N_9194,N_8705,N_6722);
and U9195 (N_9195,N_8389,N_8702);
nor U9196 (N_9196,N_7778,N_8421);
nor U9197 (N_9197,N_8369,N_7273);
nor U9198 (N_9198,N_8176,N_8812);
nand U9199 (N_9199,N_7522,N_6201);
nor U9200 (N_9200,N_8395,N_8218);
or U9201 (N_9201,N_6819,N_7784);
and U9202 (N_9202,N_6555,N_8465);
or U9203 (N_9203,N_8518,N_6426);
nor U9204 (N_9204,N_7823,N_6060);
or U9205 (N_9205,N_7023,N_8583);
xnor U9206 (N_9206,N_7671,N_6968);
or U9207 (N_9207,N_6751,N_6259);
or U9208 (N_9208,N_8425,N_7213);
and U9209 (N_9209,N_6256,N_8451);
or U9210 (N_9210,N_6541,N_7097);
and U9211 (N_9211,N_6138,N_7405);
nor U9212 (N_9212,N_7850,N_6771);
nor U9213 (N_9213,N_8210,N_7436);
nand U9214 (N_9214,N_6912,N_6759);
and U9215 (N_9215,N_8132,N_8611);
or U9216 (N_9216,N_6155,N_8023);
nand U9217 (N_9217,N_8453,N_7691);
nand U9218 (N_9218,N_6728,N_7296);
and U9219 (N_9219,N_7058,N_6505);
nor U9220 (N_9220,N_6929,N_8249);
xnor U9221 (N_9221,N_8995,N_8058);
or U9222 (N_9222,N_8748,N_6304);
and U9223 (N_9223,N_7030,N_8251);
and U9224 (N_9224,N_8556,N_8171);
or U9225 (N_9225,N_8075,N_8087);
or U9226 (N_9226,N_6190,N_8226);
and U9227 (N_9227,N_8734,N_8936);
nand U9228 (N_9228,N_7185,N_6324);
or U9229 (N_9229,N_8976,N_8860);
nor U9230 (N_9230,N_7429,N_6215);
and U9231 (N_9231,N_8502,N_6600);
xnor U9232 (N_9232,N_6158,N_7596);
and U9233 (N_9233,N_6512,N_7284);
and U9234 (N_9234,N_6212,N_6768);
nand U9235 (N_9235,N_8375,N_7127);
nand U9236 (N_9236,N_8540,N_7095);
xor U9237 (N_9237,N_8479,N_7045);
nand U9238 (N_9238,N_8480,N_7748);
and U9239 (N_9239,N_7300,N_7374);
nand U9240 (N_9240,N_8763,N_6091);
xnor U9241 (N_9241,N_6062,N_7611);
nor U9242 (N_9242,N_7416,N_8396);
nor U9243 (N_9243,N_6219,N_6344);
nor U9244 (N_9244,N_8590,N_7660);
and U9245 (N_9245,N_8169,N_7462);
nand U9246 (N_9246,N_7915,N_8554);
or U9247 (N_9247,N_8143,N_6660);
nor U9248 (N_9248,N_7341,N_7055);
nor U9249 (N_9249,N_6227,N_7015);
nand U9250 (N_9250,N_6519,N_8149);
nor U9251 (N_9251,N_8351,N_7128);
or U9252 (N_9252,N_8306,N_8379);
and U9253 (N_9253,N_8507,N_6920);
and U9254 (N_9254,N_7983,N_7235);
or U9255 (N_9255,N_6080,N_8088);
or U9256 (N_9256,N_7732,N_7182);
nor U9257 (N_9257,N_7717,N_8089);
nand U9258 (N_9258,N_6576,N_6718);
or U9259 (N_9259,N_6288,N_7422);
nand U9260 (N_9260,N_8943,N_7205);
or U9261 (N_9261,N_7195,N_7712);
or U9262 (N_9262,N_8770,N_6936);
nor U9263 (N_9263,N_6992,N_7593);
or U9264 (N_9264,N_6220,N_6675);
and U9265 (N_9265,N_6225,N_7550);
nand U9266 (N_9266,N_8343,N_7005);
and U9267 (N_9267,N_6777,N_6280);
nor U9268 (N_9268,N_8626,N_6241);
or U9269 (N_9269,N_7231,N_7661);
and U9270 (N_9270,N_7694,N_6639);
nand U9271 (N_9271,N_6757,N_7692);
nor U9272 (N_9272,N_6531,N_6880);
nand U9273 (N_9273,N_7688,N_8040);
nand U9274 (N_9274,N_7209,N_7603);
and U9275 (N_9275,N_7647,N_8326);
xnor U9276 (N_9276,N_6795,N_7449);
and U9277 (N_9277,N_8737,N_6956);
and U9278 (N_9278,N_8427,N_7599);
or U9279 (N_9279,N_6414,N_8046);
or U9280 (N_9280,N_7165,N_8745);
xor U9281 (N_9281,N_8020,N_6638);
nor U9282 (N_9282,N_6058,N_7179);
nand U9283 (N_9283,N_8913,N_6642);
and U9284 (N_9284,N_6455,N_8068);
or U9285 (N_9285,N_7914,N_7156);
nor U9286 (N_9286,N_6916,N_6018);
nor U9287 (N_9287,N_6437,N_6788);
or U9288 (N_9288,N_6378,N_8566);
nor U9289 (N_9289,N_8283,N_7564);
nor U9290 (N_9290,N_6471,N_8100);
nor U9291 (N_9291,N_7086,N_7243);
nor U9292 (N_9292,N_7959,N_7892);
and U9293 (N_9293,N_7807,N_7665);
nor U9294 (N_9294,N_6859,N_6983);
nand U9295 (N_9295,N_6113,N_8560);
nand U9296 (N_9296,N_8334,N_7868);
nor U9297 (N_9297,N_7013,N_7630);
nor U9298 (N_9298,N_8081,N_7626);
or U9299 (N_9299,N_7240,N_8167);
nor U9300 (N_9300,N_8599,N_8304);
nor U9301 (N_9301,N_6763,N_8506);
or U9302 (N_9302,N_6202,N_7789);
nor U9303 (N_9303,N_8650,N_6749);
or U9304 (N_9304,N_8501,N_7458);
nand U9305 (N_9305,N_7533,N_7286);
or U9306 (N_9306,N_7894,N_7200);
or U9307 (N_9307,N_6391,N_6967);
or U9308 (N_9308,N_6164,N_6521);
xor U9309 (N_9309,N_7632,N_6203);
and U9310 (N_9310,N_7819,N_8722);
or U9311 (N_9311,N_8844,N_7891);
and U9312 (N_9312,N_6268,N_6242);
or U9313 (N_9313,N_8742,N_7112);
nand U9314 (N_9314,N_8973,N_6559);
and U9315 (N_9315,N_8145,N_7921);
nand U9316 (N_9316,N_8281,N_6258);
nand U9317 (N_9317,N_8199,N_7134);
xnor U9318 (N_9318,N_6142,N_8629);
nor U9319 (N_9319,N_8930,N_7975);
and U9320 (N_9320,N_8655,N_8545);
nand U9321 (N_9321,N_6752,N_6392);
or U9322 (N_9322,N_8092,N_7805);
and U9323 (N_9323,N_8392,N_8104);
nand U9324 (N_9324,N_7765,N_6474);
nor U9325 (N_9325,N_7771,N_8448);
nor U9326 (N_9326,N_7206,N_6145);
and U9327 (N_9327,N_8666,N_6529);
nor U9328 (N_9328,N_8027,N_8499);
nand U9329 (N_9329,N_8975,N_6740);
nand U9330 (N_9330,N_7250,N_8108);
or U9331 (N_9331,N_6940,N_6877);
and U9332 (N_9332,N_6782,N_7016);
nand U9333 (N_9333,N_6191,N_8007);
nor U9334 (N_9334,N_8464,N_7474);
nor U9335 (N_9335,N_6127,N_7574);
and U9336 (N_9336,N_8013,N_8048);
nor U9337 (N_9337,N_6261,N_7663);
and U9338 (N_9338,N_6193,N_7192);
and U9339 (N_9339,N_7012,N_7406);
or U9340 (N_9340,N_7257,N_8869);
or U9341 (N_9341,N_8572,N_7991);
or U9342 (N_9342,N_7836,N_6524);
and U9343 (N_9343,N_6794,N_8959);
or U9344 (N_9344,N_8069,N_7121);
nor U9345 (N_9345,N_6342,N_8091);
nor U9346 (N_9346,N_8967,N_6278);
xor U9347 (N_9347,N_6088,N_6933);
and U9348 (N_9348,N_8062,N_6980);
nor U9349 (N_9349,N_8827,N_8873);
nor U9350 (N_9350,N_7342,N_6770);
xor U9351 (N_9351,N_7350,N_7990);
and U9352 (N_9352,N_8387,N_8407);
and U9353 (N_9353,N_8452,N_7499);
and U9354 (N_9354,N_7106,N_7312);
nor U9355 (N_9355,N_7486,N_7322);
or U9356 (N_9356,N_6254,N_7737);
and U9357 (N_9357,N_7244,N_8488);
nand U9358 (N_9358,N_8876,N_6646);
or U9359 (N_9359,N_8587,N_7718);
nor U9360 (N_9360,N_6716,N_7484);
nand U9361 (N_9361,N_6265,N_8530);
nor U9362 (N_9362,N_8920,N_6305);
or U9363 (N_9363,N_7020,N_6626);
or U9364 (N_9364,N_8378,N_7102);
xnor U9365 (N_9365,N_7373,N_8120);
nor U9366 (N_9366,N_6753,N_8563);
nand U9367 (N_9367,N_8235,N_7011);
nor U9368 (N_9368,N_8168,N_8263);
or U9369 (N_9369,N_6159,N_7761);
xor U9370 (N_9370,N_8901,N_7996);
nand U9371 (N_9371,N_6403,N_7493);
nand U9372 (N_9372,N_6628,N_7224);
nor U9373 (N_9373,N_6167,N_8116);
nand U9374 (N_9374,N_8348,N_6825);
and U9375 (N_9375,N_6338,N_6336);
nand U9376 (N_9376,N_6787,N_7870);
nand U9377 (N_9377,N_6528,N_6755);
nand U9378 (N_9378,N_8549,N_6732);
and U9379 (N_9379,N_7567,N_6629);
nor U9380 (N_9380,N_6511,N_8997);
nor U9381 (N_9381,N_6985,N_7475);
xnor U9382 (N_9382,N_7616,N_6681);
nand U9383 (N_9383,N_8574,N_8993);
and U9384 (N_9384,N_8987,N_8950);
nor U9385 (N_9385,N_8225,N_6004);
nand U9386 (N_9386,N_8923,N_6335);
or U9387 (N_9387,N_7482,N_6900);
and U9388 (N_9388,N_8450,N_7290);
or U9389 (N_9389,N_7866,N_8400);
nor U9390 (N_9390,N_7749,N_8998);
nor U9391 (N_9391,N_6510,N_8544);
nor U9392 (N_9392,N_7129,N_8679);
and U9393 (N_9393,N_7793,N_8830);
nand U9394 (N_9394,N_6171,N_7885);
nor U9395 (N_9395,N_6068,N_6878);
and U9396 (N_9396,N_8277,N_6721);
nor U9397 (N_9397,N_8864,N_6014);
or U9398 (N_9398,N_6001,N_6492);
nand U9399 (N_9399,N_6144,N_8319);
nand U9400 (N_9400,N_7909,N_6101);
or U9401 (N_9401,N_7399,N_8254);
or U9402 (N_9402,N_7721,N_6811);
nand U9403 (N_9403,N_6246,N_7090);
nand U9404 (N_9404,N_7841,N_8849);
or U9405 (N_9405,N_6563,N_7924);
nor U9406 (N_9406,N_6941,N_7572);
or U9407 (N_9407,N_8577,N_7472);
and U9408 (N_9408,N_7560,N_6120);
or U9409 (N_9409,N_8819,N_8158);
and U9410 (N_9410,N_6578,N_7420);
or U9411 (N_9411,N_6468,N_8848);
xnor U9412 (N_9412,N_6824,N_8289);
nor U9413 (N_9413,N_7776,N_8372);
and U9414 (N_9414,N_7757,N_6691);
nor U9415 (N_9415,N_7770,N_8129);
and U9416 (N_9416,N_7958,N_8651);
and U9417 (N_9417,N_7755,N_7324);
nand U9418 (N_9418,N_8619,N_7093);
nand U9419 (N_9419,N_8347,N_7741);
nand U9420 (N_9420,N_8200,N_6490);
or U9421 (N_9421,N_6988,N_8469);
nand U9422 (N_9422,N_6346,N_8729);
and U9423 (N_9423,N_7968,N_8484);
xor U9424 (N_9424,N_6204,N_8712);
nand U9425 (N_9425,N_7723,N_7901);
and U9426 (N_9426,N_7558,N_8579);
or U9427 (N_9427,N_6489,N_8061);
xnor U9428 (N_9428,N_6273,N_6911);
and U9429 (N_9429,N_7237,N_6679);
nand U9430 (N_9430,N_8386,N_6244);
nand U9431 (N_9431,N_7781,N_7531);
and U9432 (N_9432,N_7536,N_7961);
and U9433 (N_9433,N_6290,N_7621);
nand U9434 (N_9434,N_8839,N_6274);
or U9435 (N_9435,N_8123,N_8905);
and U9436 (N_9436,N_8999,N_7625);
xnor U9437 (N_9437,N_7230,N_8580);
nand U9438 (N_9438,N_7877,N_7172);
xor U9439 (N_9439,N_7487,N_6613);
and U9440 (N_9440,N_8197,N_7766);
or U9441 (N_9441,N_6889,N_8439);
nor U9442 (N_9442,N_6399,N_6173);
and U9443 (N_9443,N_7542,N_6606);
or U9444 (N_9444,N_6739,N_6513);
xnor U9445 (N_9445,N_6189,N_8279);
nor U9446 (N_9446,N_8543,N_8720);
or U9447 (N_9447,N_7066,N_8529);
nor U9448 (N_9448,N_6837,N_7038);
nor U9449 (N_9449,N_8985,N_7553);
nand U9450 (N_9450,N_8355,N_7211);
nand U9451 (N_9451,N_6548,N_7820);
or U9452 (N_9452,N_8297,N_7973);
and U9453 (N_9453,N_8561,N_8202);
or U9454 (N_9454,N_7187,N_8979);
or U9455 (N_9455,N_7612,N_8107);
or U9456 (N_9456,N_7938,N_7869);
nand U9457 (N_9457,N_6790,N_8429);
nand U9458 (N_9458,N_7392,N_8754);
and U9459 (N_9459,N_6823,N_7335);
nor U9460 (N_9460,N_8969,N_8884);
or U9461 (N_9461,N_7816,N_6461);
xnor U9462 (N_9462,N_8942,N_8825);
nor U9463 (N_9463,N_6705,N_7287);
nand U9464 (N_9464,N_7540,N_6373);
and U9465 (N_9465,N_8183,N_6277);
nor U9466 (N_9466,N_8240,N_8617);
nor U9467 (N_9467,N_7261,N_8093);
nor U9468 (N_9468,N_7575,N_6922);
nand U9469 (N_9469,N_6785,N_6237);
nand U9470 (N_9470,N_8683,N_7167);
and U9471 (N_9471,N_6973,N_8787);
nand U9472 (N_9472,N_8242,N_6695);
nor U9473 (N_9473,N_7927,N_8189);
nor U9474 (N_9474,N_6892,N_7309);
and U9475 (N_9475,N_6341,N_6374);
or U9476 (N_9476,N_7974,N_7191);
or U9477 (N_9477,N_7517,N_6089);
and U9478 (N_9478,N_8723,N_8476);
nand U9479 (N_9479,N_6654,N_6797);
or U9480 (N_9480,N_8179,N_8687);
nor U9481 (N_9481,N_8932,N_8778);
nor U9482 (N_9482,N_8652,N_6251);
or U9483 (N_9483,N_6485,N_8917);
xor U9484 (N_9484,N_6767,N_8066);
or U9485 (N_9485,N_8986,N_6149);
nand U9486 (N_9486,N_6789,N_7662);
nand U9487 (N_9487,N_8836,N_7565);
and U9488 (N_9488,N_6836,N_8960);
and U9489 (N_9489,N_6224,N_6551);
nand U9490 (N_9490,N_6924,N_6715);
or U9491 (N_9491,N_8099,N_8494);
or U9492 (N_9492,N_6078,N_6676);
and U9493 (N_9493,N_6311,N_8916);
nand U9494 (N_9494,N_6432,N_6393);
nand U9495 (N_9495,N_6308,N_6776);
xor U9496 (N_9496,N_6855,N_8238);
nand U9497 (N_9497,N_8828,N_7893);
nor U9498 (N_9498,N_6319,N_8850);
or U9499 (N_9499,N_8454,N_7238);
nor U9500 (N_9500,N_7949,N_8382);
nand U9501 (N_9501,N_7289,N_7880);
nand U9502 (N_9502,N_8741,N_8475);
or U9503 (N_9503,N_8403,N_8065);
xnor U9504 (N_9504,N_7485,N_7908);
or U9505 (N_9505,N_7715,N_6938);
nor U9506 (N_9506,N_6955,N_8118);
or U9507 (N_9507,N_7886,N_7750);
or U9508 (N_9508,N_6591,N_8411);
nand U9509 (N_9509,N_8989,N_6153);
or U9510 (N_9510,N_8622,N_8604);
nand U9511 (N_9511,N_8121,N_7608);
xnor U9512 (N_9512,N_8383,N_7631);
nand U9513 (N_9513,N_7800,N_6598);
nor U9514 (N_9514,N_7124,N_6292);
and U9515 (N_9515,N_8490,N_6614);
and U9516 (N_9516,N_7078,N_6221);
or U9517 (N_9517,N_6896,N_6354);
or U9518 (N_9518,N_8962,N_6396);
nor U9519 (N_9519,N_8112,N_6864);
nand U9520 (N_9520,N_7787,N_6321);
nor U9521 (N_9521,N_8402,N_8725);
nand U9522 (N_9522,N_7176,N_6366);
or U9523 (N_9523,N_8533,N_6890);
nor U9524 (N_9524,N_6546,N_8889);
nor U9525 (N_9525,N_8662,N_6821);
and U9526 (N_9526,N_7477,N_6595);
nand U9527 (N_9527,N_6298,N_6543);
or U9528 (N_9528,N_7679,N_7942);
or U9529 (N_9529,N_7116,N_8956);
xnor U9530 (N_9530,N_8340,N_6930);
nand U9531 (N_9531,N_6872,N_6012);
xor U9532 (N_9532,N_6445,N_6389);
nor U9533 (N_9533,N_7411,N_8492);
nand U9534 (N_9534,N_6761,N_6637);
and U9535 (N_9535,N_8257,N_8074);
or U9536 (N_9536,N_7463,N_6059);
and U9537 (N_9537,N_8216,N_8816);
xnor U9538 (N_9538,N_7547,N_7490);
or U9539 (N_9539,N_6231,N_6736);
nor U9540 (N_9540,N_6625,N_7675);
and U9541 (N_9541,N_7650,N_7190);
nor U9542 (N_9542,N_8717,N_8416);
and U9543 (N_9543,N_8161,N_7272);
xor U9544 (N_9544,N_7383,N_6725);
or U9545 (N_9545,N_8482,N_8585);
nand U9546 (N_9546,N_7252,N_6990);
or U9547 (N_9547,N_8937,N_8696);
nand U9548 (N_9548,N_8649,N_6603);
and U9549 (N_9549,N_8548,N_7376);
nor U9550 (N_9550,N_6170,N_7977);
nand U9551 (N_9551,N_6826,N_6908);
xnor U9552 (N_9552,N_7897,N_8274);
nor U9553 (N_9553,N_8435,N_8491);
or U9554 (N_9554,N_7855,N_6333);
nor U9555 (N_9555,N_8924,N_8174);
nand U9556 (N_9556,N_8418,N_7948);
nor U9557 (N_9557,N_6128,N_8952);
nand U9558 (N_9558,N_6415,N_8011);
nand U9559 (N_9559,N_6670,N_6833);
or U9560 (N_9560,N_7196,N_8780);
nor U9561 (N_9561,N_6034,N_7447);
and U9562 (N_9562,N_7526,N_6200);
and U9563 (N_9563,N_8090,N_7113);
nand U9564 (N_9564,N_7678,N_6645);
and U9565 (N_9565,N_7189,N_6762);
or U9566 (N_9566,N_6425,N_7204);
or U9567 (N_9567,N_8538,N_7098);
or U9568 (N_9568,N_6238,N_7471);
and U9569 (N_9569,N_6409,N_6694);
nand U9570 (N_9570,N_8631,N_7386);
and U9571 (N_9571,N_8638,N_7561);
or U9572 (N_9572,N_8510,N_7790);
nor U9573 (N_9573,N_6480,N_8150);
and U9574 (N_9574,N_6537,N_6386);
or U9575 (N_9575,N_8159,N_7656);
xor U9576 (N_9576,N_7745,N_8485);
nor U9577 (N_9577,N_6049,N_6618);
nor U9578 (N_9578,N_7178,N_7375);
or U9579 (N_9579,N_6084,N_6194);
nor U9580 (N_9580,N_8211,N_6102);
nor U9581 (N_9581,N_8460,N_8207);
and U9582 (N_9582,N_6588,N_7676);
or U9583 (N_9583,N_7638,N_7336);
nor U9584 (N_9584,N_6413,N_6931);
nand U9585 (N_9585,N_7642,N_8783);
nand U9586 (N_9586,N_7871,N_7111);
nand U9587 (N_9587,N_7118,N_8517);
nand U9588 (N_9588,N_7110,N_8001);
nor U9589 (N_9589,N_7772,N_7248);
and U9590 (N_9590,N_6608,N_8750);
or U9591 (N_9591,N_8643,N_6351);
or U9592 (N_9592,N_7597,N_6452);
or U9593 (N_9593,N_6913,N_6714);
and U9594 (N_9594,N_6478,N_6156);
nor U9595 (N_9595,N_7956,N_6742);
nand U9596 (N_9596,N_6648,N_6495);
or U9597 (N_9597,N_7227,N_8341);
or U9598 (N_9598,N_7981,N_7792);
nor U9599 (N_9599,N_8208,N_8461);
xor U9600 (N_9600,N_6050,N_8694);
or U9601 (N_9601,N_8234,N_6283);
xor U9602 (N_9602,N_7972,N_7340);
and U9603 (N_9603,N_8468,N_6307);
xor U9604 (N_9604,N_7164,N_7941);
and U9605 (N_9605,N_8026,N_8434);
nand U9606 (N_9606,N_7937,N_8616);
or U9607 (N_9607,N_7370,N_8675);
xor U9608 (N_9608,N_8692,N_6520);
nor U9609 (N_9609,N_6350,N_6652);
or U9610 (N_9610,N_7695,N_6672);
nand U9611 (N_9611,N_7875,N_7282);
and U9612 (N_9612,N_6323,N_8330);
nand U9613 (N_9613,N_7666,N_8472);
and U9614 (N_9614,N_7354,N_7168);
nor U9615 (N_9615,N_8514,N_7169);
or U9616 (N_9616,N_6592,N_8797);
or U9617 (N_9617,N_8906,N_8513);
nand U9618 (N_9618,N_8044,N_6028);
xnor U9619 (N_9619,N_6743,N_6666);
nor U9620 (N_9620,N_6210,N_8291);
nor U9621 (N_9621,N_7329,N_6849);
nor U9622 (N_9622,N_6460,N_6939);
xnor U9623 (N_9623,N_8776,N_7225);
xor U9624 (N_9624,N_8636,N_8772);
nor U9625 (N_9625,N_8721,N_8852);
or U9626 (N_9626,N_7313,N_8799);
nor U9627 (N_9627,N_7655,N_7062);
or U9628 (N_9628,N_7404,N_6593);
nor U9629 (N_9629,N_8761,N_6651);
and U9630 (N_9630,N_8642,N_8470);
nand U9631 (N_9631,N_7285,N_6959);
and U9632 (N_9632,N_7391,N_8349);
nand U9633 (N_9633,N_7530,N_7864);
and U9634 (N_9634,N_8911,N_8981);
or U9635 (N_9635,N_8153,N_6005);
nand U9636 (N_9636,N_7507,N_7614);
and U9637 (N_9637,N_6907,N_8789);
or U9638 (N_9638,N_8802,N_6540);
nand U9639 (N_9639,N_8731,N_7683);
nor U9640 (N_9640,N_7969,N_6653);
and U9641 (N_9641,N_7451,N_6451);
or U9642 (N_9642,N_6343,N_6501);
nand U9643 (N_9643,N_7000,N_6700);
nand U9644 (N_9644,N_6419,N_8146);
and U9645 (N_9645,N_8031,N_6590);
and U9646 (N_9646,N_7320,N_8609);
nor U9647 (N_9647,N_8970,N_6781);
and U9648 (N_9648,N_8036,N_6584);
or U9649 (N_9649,N_6971,N_7727);
nor U9650 (N_9650,N_7262,N_8404);
or U9651 (N_9651,N_8393,N_7052);
nand U9652 (N_9652,N_6188,N_6053);
or U9653 (N_9653,N_7423,N_6435);
and U9654 (N_9654,N_7047,N_7277);
or U9655 (N_9655,N_6764,N_6066);
and U9656 (N_9656,N_6991,N_6615);
or U9657 (N_9657,N_6946,N_6619);
nand U9658 (N_9658,N_6803,N_6801);
nor U9659 (N_9659,N_6375,N_6972);
nor U9660 (N_9660,N_8148,N_8751);
and U9661 (N_9661,N_6038,N_6535);
and U9662 (N_9662,N_7220,N_6919);
nand U9663 (N_9663,N_6851,N_6786);
and U9664 (N_9664,N_8856,N_8857);
xor U9665 (N_9665,N_7072,N_8866);
or U9666 (N_9666,N_7264,N_6843);
nand U9667 (N_9667,N_6640,N_6387);
or U9668 (N_9668,N_6779,N_7234);
or U9669 (N_9669,N_6622,N_6944);
or U9670 (N_9670,N_6665,N_8264);
or U9671 (N_9671,N_6854,N_8245);
and U9672 (N_9672,N_8221,N_6196);
and U9673 (N_9673,N_6073,N_6405);
nand U9674 (N_9674,N_7080,N_6247);
xor U9675 (N_9675,N_8568,N_6586);
nand U9676 (N_9676,N_8621,N_8623);
and U9677 (N_9677,N_7555,N_8483);
nand U9678 (N_9678,N_7440,N_8440);
xnor U9679 (N_9679,N_6383,N_8368);
nor U9680 (N_9680,N_8907,N_8198);
xor U9681 (N_9681,N_8699,N_8041);
nor U9682 (N_9682,N_6172,N_6812);
and U9683 (N_9683,N_8134,N_7108);
or U9684 (N_9684,N_8496,N_8865);
nor U9685 (N_9685,N_8551,N_6055);
nand U9686 (N_9686,N_7985,N_8627);
nand U9687 (N_9687,N_8229,N_7068);
nor U9688 (N_9688,N_6765,N_7743);
and U9689 (N_9689,N_6964,N_7640);
xor U9690 (N_9690,N_8980,N_6580);
nand U9691 (N_9691,N_8961,N_8052);
nand U9692 (N_9692,N_7719,N_7997);
or U9693 (N_9693,N_7274,N_7573);
and U9694 (N_9694,N_6020,N_6353);
nand U9695 (N_9695,N_6573,N_8280);
or U9696 (N_9696,N_6680,N_8313);
and U9697 (N_9697,N_7545,N_6195);
and U9698 (N_9698,N_6162,N_6046);
or U9699 (N_9699,N_6888,N_7580);
and U9700 (N_9700,N_8079,N_8335);
and U9701 (N_9701,N_8656,N_7704);
nor U9702 (N_9702,N_7061,N_6813);
nand U9703 (N_9703,N_8409,N_6599);
nor U9704 (N_9704,N_8648,N_8925);
nor U9705 (N_9705,N_8072,N_6536);
nor U9706 (N_9706,N_7081,N_7605);
nand U9707 (N_9707,N_8547,N_6926);
or U9708 (N_9708,N_7598,N_7268);
or U9709 (N_9709,N_6517,N_6006);
nand U9710 (N_9710,N_8244,N_8823);
or U9711 (N_9711,N_8603,N_7978);
nor U9712 (N_9712,N_8321,N_6554);
nand U9713 (N_9713,N_7690,N_6630);
nand U9714 (N_9714,N_6064,N_7325);
nand U9715 (N_9715,N_7418,N_8824);
or U9716 (N_9716,N_6395,N_8559);
nor U9717 (N_9717,N_6289,N_6731);
nand U9718 (N_9718,N_6240,N_6429);
nand U9719 (N_9719,N_6545,N_6951);
nor U9720 (N_9720,N_8977,N_7188);
nor U9721 (N_9721,N_7637,N_7965);
nand U9722 (N_9722,N_7714,N_8206);
or U9723 (N_9723,N_6465,N_8302);
and U9724 (N_9724,N_6255,N_8542);
nand U9725 (N_9725,N_7107,N_6798);
xnor U9726 (N_9726,N_7353,N_6017);
and U9727 (N_9727,N_8336,N_6077);
xnor U9728 (N_9728,N_6228,N_8669);
nand U9729 (N_9729,N_6796,N_8345);
and U9730 (N_9730,N_8541,N_8711);
nand U9731 (N_9731,N_7385,N_7171);
nor U9732 (N_9732,N_6075,N_7270);
and U9733 (N_9733,N_7497,N_7940);
nor U9734 (N_9734,N_6928,N_8250);
xnor U9735 (N_9735,N_7303,N_7709);
nor U9736 (N_9736,N_7617,N_7177);
nand U9737 (N_9737,N_8420,N_7571);
nor U9738 (N_9738,N_7898,N_8110);
nand U9739 (N_9739,N_6623,N_6484);
xor U9740 (N_9740,N_7798,N_7735);
or U9741 (N_9741,N_8996,N_7065);
or U9742 (N_9742,N_6027,N_8632);
or U9743 (N_9743,N_8703,N_6178);
nand U9744 (N_9744,N_8680,N_6072);
nand U9745 (N_9745,N_8707,N_6689);
nor U9746 (N_9746,N_6181,N_8010);
or U9747 (N_9747,N_7999,N_8014);
nand U9748 (N_9748,N_8493,N_8320);
or U9749 (N_9749,N_8610,N_8728);
nand U9750 (N_9750,N_7217,N_7849);
and U9751 (N_9751,N_7518,N_8966);
or U9752 (N_9752,N_7944,N_7935);
or U9753 (N_9753,N_7194,N_8401);
xor U9754 (N_9754,N_8034,N_8762);
nor U9755 (N_9755,N_7535,N_8948);
xnor U9756 (N_9756,N_7524,N_8672);
nor U9757 (N_9757,N_6627,N_6087);
nor U9758 (N_9758,N_6516,N_8846);
and U9759 (N_9759,N_7584,N_6754);
or U9760 (N_9760,N_6656,N_7427);
nand U9761 (N_9761,N_7831,N_7933);
nor U9762 (N_9762,N_7900,N_7576);
and U9763 (N_9763,N_6248,N_6574);
and U9764 (N_9764,N_6430,N_7916);
xor U9765 (N_9765,N_6143,N_7180);
or U9766 (N_9766,N_7310,N_8798);
nor U9767 (N_9767,N_7856,N_6582);
or U9768 (N_9768,N_6356,N_8119);
and U9769 (N_9769,N_6966,N_7409);
or U9770 (N_9770,N_8342,N_8660);
nand U9771 (N_9771,N_7448,N_8266);
nand U9772 (N_9772,N_6157,N_7794);
and U9773 (N_9773,N_7828,N_6199);
xor U9774 (N_9774,N_8166,N_8073);
nor U9775 (N_9775,N_6683,N_8284);
and U9776 (N_9776,N_8539,N_6723);
or U9777 (N_9777,N_8060,N_7980);
nand U9778 (N_9778,N_6799,N_6828);
nand U9779 (N_9779,N_8445,N_7495);
nand U9780 (N_9780,N_8758,N_7843);
nand U9781 (N_9781,N_6698,N_7414);
or U9782 (N_9782,N_6860,N_8881);
and U9783 (N_9783,N_6483,N_7242);
nor U9784 (N_9784,N_8971,N_7412);
nand U9785 (N_9785,N_8287,N_7829);
or U9786 (N_9786,N_6997,N_7397);
and U9787 (N_9787,N_6693,N_8990);
nor U9788 (N_9788,N_7009,N_6791);
nor U9789 (N_9789,N_6447,N_8055);
nor U9790 (N_9790,N_7585,N_8628);
and U9791 (N_9791,N_6720,N_7534);
or U9792 (N_9792,N_6147,N_8562);
and U9793 (N_9793,N_8872,N_6207);
or U9794 (N_9794,N_6674,N_7738);
nand U9795 (N_9795,N_7696,N_7215);
nor U9796 (N_9796,N_8736,N_6706);
or U9797 (N_9797,N_8835,N_8139);
nor U9798 (N_9798,N_6577,N_8366);
nand U9799 (N_9799,N_6464,N_8391);
nand U9800 (N_9800,N_6213,N_8647);
nor U9801 (N_9801,N_7120,N_8458);
or U9802 (N_9802,N_8135,N_8412);
or U9803 (N_9803,N_6504,N_7473);
nand U9804 (N_9804,N_8935,N_6065);
nor U9805 (N_9805,N_8156,N_8337);
xnor U9806 (N_9806,N_8868,N_8582);
or U9807 (N_9807,N_6074,N_6125);
or U9808 (N_9808,N_7334,N_6040);
nor U9809 (N_9809,N_6838,N_6428);
xor U9810 (N_9810,N_8597,N_7527);
and U9811 (N_9811,N_6021,N_8740);
nand U9812 (N_9812,N_7082,N_8003);
nand U9813 (N_9813,N_6644,N_7291);
and U9814 (N_9814,N_8785,N_6587);
xnor U9815 (N_9815,N_6760,N_8354);
and U9816 (N_9816,N_6923,N_6439);
nor U9817 (N_9817,N_6416,N_6909);
xnor U9818 (N_9818,N_7145,N_7105);
or U9819 (N_9819,N_7161,N_6052);
nand U9820 (N_9820,N_6081,N_7838);
nand U9821 (N_9821,N_8000,N_6124);
or U9822 (N_9822,N_8550,N_8030);
nand U9823 (N_9823,N_6151,N_6408);
and U9824 (N_9824,N_6649,N_6861);
nor U9825 (N_9825,N_8775,N_7646);
and U9826 (N_9826,N_6953,N_6079);
nor U9827 (N_9827,N_8185,N_7133);
or U9828 (N_9828,N_7706,N_8755);
xnor U9829 (N_9829,N_6667,N_6205);
or U9830 (N_9830,N_7470,N_8154);
or U9831 (N_9831,N_7502,N_7146);
nand U9832 (N_9832,N_8813,N_8109);
or U9833 (N_9833,N_8504,N_8059);
and U9834 (N_9834,N_7578,N_6371);
nand U9835 (N_9835,N_6133,N_6000);
and U9836 (N_9836,N_8963,N_6310);
xor U9837 (N_9837,N_6815,N_6526);
and U9838 (N_9838,N_7042,N_7328);
and U9839 (N_9839,N_7263,N_8639);
nor U9840 (N_9840,N_8885,N_8671);
nor U9841 (N_9841,N_8405,N_6564);
nand U9842 (N_9842,N_7491,N_8805);
or U9843 (N_9843,N_7763,N_8481);
xor U9844 (N_9844,N_7478,N_8361);
nand U9845 (N_9845,N_6457,N_8436);
or U9846 (N_9846,N_6180,N_8028);
and U9847 (N_9847,N_7390,N_6487);
nor U9848 (N_9848,N_7326,N_8686);
and U9849 (N_9849,N_8593,N_8613);
nand U9850 (N_9850,N_8853,N_7801);
nand U9851 (N_9851,N_7582,N_6903);
xor U9852 (N_9852,N_8316,N_6266);
or U9853 (N_9853,N_7267,N_7004);
or U9854 (N_9854,N_8299,N_7210);
and U9855 (N_9855,N_6436,N_7089);
nor U9856 (N_9856,N_7174,N_6032);
and U9857 (N_9857,N_8443,N_8294);
nand U9858 (N_9858,N_6347,N_7664);
nand U9859 (N_9859,N_6974,N_7266);
or U9860 (N_9860,N_7314,N_7554);
nand U9861 (N_9861,N_6368,N_6663);
nand U9862 (N_9862,N_8017,N_6152);
nor U9863 (N_9863,N_8558,N_8644);
and U9864 (N_9864,N_6239,N_6249);
nor U9865 (N_9865,N_8247,N_7260);
and U9866 (N_9866,N_8730,N_6208);
and U9867 (N_9867,N_7541,N_6532);
nor U9868 (N_9868,N_7410,N_6579);
nand U9869 (N_9869,N_8915,N_7036);
or U9870 (N_9870,N_8259,N_6766);
or U9871 (N_9871,N_7457,N_7528);
nor U9872 (N_9872,N_6098,N_6122);
nor U9873 (N_9873,N_7859,N_6141);
nor U9874 (N_9874,N_8713,N_8578);
nand U9875 (N_9875,N_6918,N_6179);
nand U9876 (N_9876,N_8806,N_6260);
and U9877 (N_9877,N_6575,N_6275);
nor U9878 (N_9878,N_6748,N_7067);
nand U9879 (N_9879,N_8814,N_8248);
or U9880 (N_9880,N_6773,N_7890);
and U9881 (N_9881,N_6549,N_6267);
nor U9882 (N_9882,N_8575,N_8380);
nor U9883 (N_9883,N_7104,N_8724);
or U9884 (N_9884,N_6472,N_6817);
or U9885 (N_9885,N_6793,N_8665);
or U9886 (N_9886,N_7394,N_7512);
or U9887 (N_9887,N_6969,N_7783);
xor U9888 (N_9888,N_6876,N_7251);
and U9889 (N_9889,N_6894,N_6692);
nor U9890 (N_9890,N_8880,N_8818);
and U9891 (N_9891,N_8833,N_6476);
and U9892 (N_9892,N_7945,N_7330);
nor U9893 (N_9893,N_7670,N_7742);
or U9894 (N_9894,N_7920,N_6303);
and U9895 (N_9895,N_8367,N_6394);
and U9896 (N_9896,N_8670,N_7366);
nand U9897 (N_9897,N_8838,N_7590);
nand U9898 (N_9898,N_6250,N_6858);
nand U9899 (N_9899,N_8991,N_7017);
nor U9900 (N_9900,N_8256,N_7245);
nand U9901 (N_9901,N_7348,N_8260);
or U9902 (N_9902,N_7479,N_8515);
and U9903 (N_9903,N_8231,N_7629);
nor U9904 (N_9904,N_6611,N_7395);
and U9905 (N_9905,N_8678,N_8477);
or U9906 (N_9906,N_8760,N_7767);
and U9907 (N_9907,N_6708,N_8456);
nand U9908 (N_9908,N_8113,N_6082);
nor U9909 (N_9909,N_6879,N_8021);
and U9910 (N_9910,N_8716,N_7432);
nand U9911 (N_9911,N_7100,N_7588);
and U9912 (N_9912,N_6039,N_7481);
and U9913 (N_9913,N_7346,N_7923);
and U9914 (N_9914,N_8413,N_7620);
and U9915 (N_9915,N_6655,N_7323);
nand U9916 (N_9916,N_8050,N_8605);
or U9917 (N_9917,N_8875,N_7402);
nor U9918 (N_9918,N_6271,N_6104);
or U9919 (N_9919,N_6022,N_7559);
nor U9920 (N_9920,N_7096,N_6846);
or U9921 (N_9921,N_7644,N_6544);
or U9922 (N_9922,N_6910,N_6712);
nor U9923 (N_9923,N_7848,N_7056);
and U9924 (N_9924,N_6677,N_6100);
nor U9925 (N_9925,N_6045,N_6830);
or U9926 (N_9926,N_7957,N_8822);
or U9927 (N_9927,N_7292,N_7634);
nand U9928 (N_9928,N_6384,N_7835);
or U9929 (N_9929,N_8308,N_6174);
xnor U9930 (N_9930,N_6185,N_6296);
nor U9931 (N_9931,N_6263,N_8140);
nand U9932 (N_9932,N_6737,N_8796);
nor U9933 (N_9933,N_6934,N_6230);
nand U9934 (N_9934,N_6634,N_6806);
nor U9935 (N_9935,N_7109,N_6137);
nand U9936 (N_9936,N_7151,N_6961);
and U9937 (N_9937,N_6491,N_8607);
nor U9938 (N_9938,N_7747,N_7769);
xor U9939 (N_9939,N_6030,N_6331);
or U9940 (N_9940,N_6800,N_6557);
nor U9941 (N_9941,N_6160,N_7157);
and U9942 (N_9942,N_6359,N_7345);
nor U9943 (N_9943,N_7046,N_7780);
or U9944 (N_9944,N_8292,N_7201);
nand U9945 (N_9945,N_8804,N_8667);
nor U9946 (N_9946,N_6008,N_8173);
and U9947 (N_9947,N_7400,N_6558);
and U9948 (N_9948,N_7883,N_7337);
nand U9949 (N_9949,N_6071,N_7768);
or U9950 (N_9950,N_7682,N_7029);
nand U9951 (N_9951,N_8896,N_8471);
or U9952 (N_9952,N_8303,N_6015);
nand U9953 (N_9953,N_8682,N_7931);
and U9954 (N_9954,N_8965,N_6025);
or U9955 (N_9955,N_7925,N_6932);
or U9956 (N_9956,N_7899,N_7006);
nand U9957 (N_9957,N_8769,N_8941);
and U9958 (N_9958,N_8620,N_7833);
nor U9959 (N_9959,N_7703,N_7028);
and U9960 (N_9960,N_6117,N_7358);
nor U9961 (N_9961,N_6236,N_7932);
nor U9962 (N_9962,N_8275,N_7359);
or U9963 (N_9963,N_7302,N_8486);
nor U9964 (N_9964,N_8285,N_8363);
or U9965 (N_9965,N_8160,N_7381);
or U9966 (N_9966,N_8419,N_6056);
or U9967 (N_9967,N_8305,N_8726);
or U9968 (N_9968,N_6935,N_7456);
and U9969 (N_9969,N_6784,N_7884);
nor U9970 (N_9970,N_8332,N_8698);
and U9971 (N_9971,N_7003,N_7803);
and U9972 (N_9972,N_7021,N_7863);
or U9973 (N_9973,N_7327,N_8268);
nand U9974 (N_9974,N_8808,N_8663);
and U9975 (N_9975,N_6962,N_7929);
and U9976 (N_9976,N_8317,N_6482);
and U9977 (N_9977,N_6950,N_6314);
nor U9978 (N_9978,N_6589,N_7511);
or U9979 (N_9979,N_7186,N_6284);
nand U9980 (N_9980,N_8584,N_6539);
nand U9981 (N_9981,N_7606,N_7998);
xor U9982 (N_9982,N_6226,N_6320);
and U9983 (N_9983,N_7389,N_8024);
nand U9984 (N_9984,N_7279,N_6352);
or U9985 (N_9985,N_6317,N_7902);
or U9986 (N_9986,N_7071,N_8858);
or U9987 (N_9987,N_8992,N_7307);
nor U9988 (N_9988,N_6816,N_6507);
or U9989 (N_9989,N_7853,N_6041);
nand U9990 (N_9990,N_6963,N_7025);
nor U9991 (N_9991,N_8586,N_7839);
nor U9992 (N_9992,N_6947,N_8246);
and U9993 (N_9993,N_8927,N_7464);
nand U9994 (N_9994,N_8520,N_8898);
and U9995 (N_9995,N_7734,N_7865);
xor U9996 (N_9996,N_7114,N_8295);
and U9997 (N_9997,N_7821,N_7591);
or U9998 (N_9998,N_8111,N_8344);
or U9999 (N_9999,N_8459,N_8635);
or U10000 (N_10000,N_7494,N_7910);
or U10001 (N_10001,N_8801,N_6856);
nand U10002 (N_10002,N_7137,N_6214);
nor U10003 (N_10003,N_6996,N_8296);
nand U10004 (N_10004,N_8212,N_7722);
xnor U10005 (N_10005,N_8076,N_7281);
or U10006 (N_10006,N_7468,N_6747);
nand U10007 (N_10007,N_7051,N_8474);
or U10008 (N_10008,N_8298,N_6624);
nand U10009 (N_10009,N_6711,N_6362);
nor U10010 (N_10010,N_7752,N_8441);
or U10011 (N_10011,N_8293,N_7360);
or U10012 (N_10012,N_8938,N_6007);
nand U10013 (N_10013,N_6467,N_6704);
nor U10014 (N_10014,N_7579,N_7548);
xnor U10015 (N_10015,N_6318,N_8278);
or U10016 (N_10016,N_7019,N_7699);
or U10017 (N_10017,N_8239,N_8753);
nand U10018 (N_10018,N_6281,N_7453);
and U10019 (N_10019,N_8739,N_8700);
or U10020 (N_10020,N_8934,N_6313);
or U10021 (N_10021,N_7525,N_7529);
xor U10022 (N_10022,N_6852,N_8919);
nand U10023 (N_10023,N_7198,N_8323);
nor U10024 (N_10024,N_6994,N_6234);
or U10025 (N_10025,N_6509,N_8201);
nor U10026 (N_10026,N_8931,N_6477);
nor U10027 (N_10027,N_7040,N_7720);
nor U10028 (N_10028,N_8155,N_7254);
nor U10029 (N_10029,N_7813,N_8309);
xnor U10030 (N_10030,N_6867,N_8589);
and U10031 (N_10031,N_7466,N_8184);
xnor U10032 (N_10032,N_8033,N_8949);
nand U10033 (N_10033,N_8417,N_6818);
and U10034 (N_10034,N_6915,N_7150);
and U10035 (N_10035,N_6868,N_8191);
and U10036 (N_10036,N_6420,N_6099);
and U10037 (N_10037,N_7607,N_6945);
or U10038 (N_10038,N_7306,N_7685);
or U10039 (N_10039,N_7791,N_7026);
or U10040 (N_10040,N_7516,N_7369);
nor U10041 (N_10041,N_7488,N_8217);
nor U10042 (N_10042,N_8125,N_8641);
nand U10043 (N_10043,N_8265,N_7513);
and U10044 (N_10044,N_8674,N_7349);
nor U10045 (N_10045,N_8137,N_6112);
nor U10046 (N_10046,N_6746,N_6729);
nand U10047 (N_10047,N_6316,N_6253);
nor U10048 (N_10048,N_7814,N_7014);
or U10049 (N_10049,N_8862,N_6085);
and U10050 (N_10050,N_7636,N_8124);
nand U10051 (N_10051,N_7872,N_8360);
and U10052 (N_10052,N_8253,N_8181);
nand U10053 (N_10053,N_7317,N_6875);
nor U10054 (N_10054,N_6036,N_8083);
xor U10055 (N_10055,N_7053,N_6702);
nand U10056 (N_10056,N_6381,N_7653);
or U10057 (N_10057,N_7896,N_6954);
and U10058 (N_10058,N_7152,N_8781);
xor U10059 (N_10059,N_7459,N_7393);
nand U10060 (N_10060,N_8446,N_8495);
or U10061 (N_10061,N_8043,N_8795);
xor U10062 (N_10062,N_8749,N_8710);
and U10063 (N_10063,N_7070,N_8049);
nor U10064 (N_10064,N_7764,N_6211);
nand U10065 (N_10065,N_8455,N_6023);
xnor U10066 (N_10066,N_6897,N_7379);
and U10067 (N_10067,N_8141,N_8105);
nor U10068 (N_10068,N_7199,N_7551);
nor U10069 (N_10069,N_8602,N_7557);
xor U10070 (N_10070,N_8845,N_8791);
nand U10071 (N_10071,N_7539,N_8893);
and U10072 (N_10072,N_6533,N_8214);
or U10073 (N_10073,N_6009,N_6840);
and U10074 (N_10074,N_8673,N_7759);
nor U10075 (N_10075,N_8695,N_8232);
nand U10076 (N_10076,N_7984,N_8929);
and U10077 (N_10077,N_8064,N_7854);
or U10078 (N_10078,N_6132,N_6063);
and U10079 (N_10079,N_7775,N_8888);
nor U10080 (N_10080,N_7888,N_6090);
nand U10081 (N_10081,N_6502,N_8581);
xor U10082 (N_10082,N_7546,N_6197);
and U10083 (N_10083,N_8045,N_8331);
or U10084 (N_10084,N_8182,N_8433);
or U10085 (N_10085,N_7583,N_6493);
or U10086 (N_10086,N_8300,N_8933);
and U10087 (N_10087,N_7437,N_7054);
or U10088 (N_10088,N_8768,N_8552);
nor U10089 (N_10089,N_8689,N_8614);
nand U10090 (N_10090,N_7930,N_8084);
and U10091 (N_10091,N_6895,N_8921);
nor U10092 (N_10092,N_7619,N_6690);
nand U10093 (N_10093,N_6633,N_7873);
or U10094 (N_10094,N_7455,N_8038);
nor U10095 (N_10095,N_6168,N_7658);
nor U10096 (N_10096,N_6044,N_8237);
and U10097 (N_10097,N_6166,N_8358);
or U10098 (N_10098,N_6594,N_8633);
xnor U10099 (N_10099,N_8432,N_7860);
or U10100 (N_10100,N_7812,N_7103);
and U10101 (N_10101,N_6223,N_7063);
and U10102 (N_10102,N_6769,N_7818);
or U10103 (N_10103,N_6412,N_8854);
nor U10104 (N_10104,N_8505,N_7520);
nor U10105 (N_10105,N_8290,N_7278);
and U10106 (N_10106,N_6792,N_6309);
or U10107 (N_10107,N_6083,N_7889);
and U10108 (N_10108,N_6095,N_7384);
or U10109 (N_10109,N_8592,N_7876);
or U10110 (N_10110,N_6243,N_7806);
or U10111 (N_10111,N_8056,N_7170);
and U10112 (N_10112,N_6870,N_8657);
nor U10113 (N_10113,N_7887,N_6881);
nor U10114 (N_10114,N_8054,N_8258);
or U10115 (N_10115,N_8706,N_6111);
and U10116 (N_10116,N_7947,N_8668);
xor U10117 (N_10117,N_6561,N_6921);
nand U10118 (N_10118,N_7628,N_6886);
xor U10119 (N_10119,N_7173,N_6899);
xor U10120 (N_10120,N_8774,N_7515);
or U10121 (N_10121,N_7123,N_6423);
nand U10122 (N_10122,N_7438,N_7982);
or U10123 (N_10123,N_8398,N_7333);
nor U10124 (N_10124,N_6986,N_8489);
nand U10125 (N_10125,N_6874,N_7294);
or U10126 (N_10126,N_7963,N_6713);
xnor U10127 (N_10127,N_7378,N_6508);
nor U10128 (N_10128,N_7445,N_8784);
nand U10129 (N_10129,N_8193,N_6917);
nor U10130 (N_10130,N_6106,N_8047);
xor U10131 (N_10131,N_7131,N_8792);
nand U10132 (N_10132,N_8098,N_8764);
nor U10133 (N_10133,N_7913,N_7141);
nand U10134 (N_10134,N_7622,N_7736);
nor U10135 (N_10135,N_7955,N_6636);
nor U10136 (N_10136,N_8615,N_6306);
or U10137 (N_10137,N_6669,N_6361);
or U10138 (N_10138,N_6364,N_7075);
nand U10139 (N_10139,N_6829,N_7609);
nor U10140 (N_10140,N_7480,N_8511);
or U10141 (N_10141,N_7034,N_8654);
nor U10142 (N_10142,N_6330,N_6033);
nor U10143 (N_10143,N_6421,N_6440);
and U10144 (N_10144,N_6183,N_6329);
or U10145 (N_10145,N_6218,N_6538);
or U10146 (N_10146,N_6566,N_8016);
nand U10147 (N_10147,N_7729,N_8377);
nand U10148 (N_10148,N_8532,N_7132);
nor U10149 (N_10149,N_6658,N_6925);
nand U10150 (N_10150,N_8365,N_6738);
nand U10151 (N_10151,N_8951,N_6047);
nor U10152 (N_10152,N_7088,N_7259);
or U10153 (N_10153,N_7952,N_6993);
and U10154 (N_10154,N_6450,N_7731);
or U10155 (N_10155,N_7840,N_8840);
nor U10156 (N_10156,N_7788,N_7881);
nor U10157 (N_10157,N_7739,N_7834);
nor U10158 (N_10158,N_6475,N_7936);
or U10159 (N_10159,N_7648,N_7862);
and U10160 (N_10160,N_6322,N_7049);
nor U10161 (N_10161,N_8042,N_6411);
or U10162 (N_10162,N_6687,N_7338);
nor U10163 (N_10163,N_6369,N_7970);
or U10164 (N_10164,N_8859,N_6805);
nand U10165 (N_10165,N_6831,N_7510);
and U10166 (N_10166,N_7993,N_6756);
and U10167 (N_10167,N_6136,N_8236);
and U10168 (N_10168,N_6061,N_8288);
or U10169 (N_10169,N_6462,N_8900);
or U10170 (N_10170,N_6216,N_6998);
nand U10171 (N_10171,N_7852,N_7228);
and U10172 (N_10172,N_7315,N_7417);
nand U10173 (N_10173,N_8032,N_7532);
and U10174 (N_10174,N_7304,N_7971);
nor U10175 (N_10175,N_6958,N_8718);
nor U10176 (N_10176,N_7092,N_6750);
nor U10177 (N_10177,N_8829,N_8025);
and U10178 (N_10178,N_8194,N_8195);
and U10179 (N_10179,N_6807,N_7521);
nand U10180 (N_10180,N_6857,N_7519);
nor U10181 (N_10181,N_8557,N_8744);
or U10182 (N_10182,N_6337,N_8163);
nor U10183 (N_10183,N_8102,N_8645);
and U10184 (N_10184,N_8646,N_7779);
nor U10185 (N_10185,N_6135,N_7774);
and U10186 (N_10186,N_8525,N_6339);
or U10187 (N_10187,N_7686,N_7505);
nand U10188 (N_10188,N_8478,N_8130);
and U10189 (N_10189,N_8922,N_7994);
nor U10190 (N_10190,N_8624,N_8867);
nor U10191 (N_10191,N_8203,N_6161);
or U10192 (N_10192,N_7817,N_8928);
nand U10193 (N_10193,N_7033,N_6893);
nand U10194 (N_10194,N_7076,N_8127);
nor U10195 (N_10195,N_7297,N_6664);
and U10196 (N_10196,N_6869,N_6291);
and U10197 (N_10197,N_7698,N_6146);
and U10198 (N_10198,N_8945,N_8078);
and U10199 (N_10199,N_6334,N_7716);
or U10200 (N_10200,N_7439,N_7444);
nor U10201 (N_10201,N_8196,N_8410);
or U10202 (N_10202,N_7895,N_8384);
or U10203 (N_10203,N_7181,N_7355);
nor U10204 (N_10204,N_8837,N_6999);
and U10205 (N_10205,N_8984,N_7651);
nand U10206 (N_10206,N_8863,N_6182);
and U10207 (N_10207,N_8339,N_7740);
or U10208 (N_10208,N_8759,N_8534);
or U10209 (N_10209,N_8219,N_7212);
and U10210 (N_10210,N_7388,N_7483);
and U10211 (N_10211,N_8894,N_7500);
nand U10212 (N_10212,N_8841,N_8957);
or U10213 (N_10213,N_6684,N_6848);
and U10214 (N_10214,N_8188,N_7008);
or U10215 (N_10215,N_6662,N_6778);
or U10216 (N_10216,N_7645,N_7570);
and U10217 (N_10217,N_7059,N_8142);
nor U10218 (N_10218,N_7442,N_7842);
nand U10219 (N_10219,N_8954,N_6438);
and U10220 (N_10220,N_7351,N_8904);
and U10221 (N_10221,N_7946,N_6410);
xor U10222 (N_10222,N_7331,N_6735);
nand U10223 (N_10223,N_7162,N_6604);
nor U10224 (N_10224,N_7203,N_6187);
xor U10225 (N_10225,N_8487,N_8224);
xnor U10226 (N_10226,N_6397,N_7905);
nor U10227 (N_10227,N_7592,N_7879);
or U10228 (N_10228,N_6401,N_6905);
nor U10229 (N_10229,N_8630,N_6948);
or U10230 (N_10230,N_7751,N_8573);
nor U10231 (N_10231,N_8408,N_6121);
and U10232 (N_10232,N_7452,N_8803);
or U10233 (N_10233,N_6422,N_7867);
xor U10234 (N_10234,N_6446,N_8886);
and U10235 (N_10235,N_8757,N_7702);
nand U10236 (N_10236,N_8899,N_6232);
or U10237 (N_10237,N_8390,N_8371);
or U10238 (N_10238,N_6057,N_6377);
and U10239 (N_10239,N_6534,N_8765);
and U10240 (N_10240,N_7119,N_7010);
and U10241 (N_10241,N_8512,N_6286);
or U10242 (N_10242,N_6390,N_7733);
and U10243 (N_10243,N_6456,N_6177);
nor U10244 (N_10244,N_8423,N_6960);
nor U10245 (N_10245,N_6184,N_6070);
nor U10246 (N_10246,N_6506,N_8269);
or U10247 (N_10247,N_7265,N_8571);
and U10248 (N_10248,N_7060,N_7057);
or U10249 (N_10249,N_7911,N_6235);
xor U10250 (N_10250,N_7906,N_8394);
or U10251 (N_10251,N_8871,N_6984);
xnor U10252 (N_10252,N_8606,N_7595);
or U10253 (N_10253,N_7762,N_6404);
nand U10254 (N_10254,N_6372,N_6952);
nor U10255 (N_10255,N_6832,N_8286);
xor U10256 (N_10256,N_8897,N_6657);
and U10257 (N_10257,N_8909,N_8883);
or U10258 (N_10258,N_7280,N_8157);
and U10259 (N_10259,N_7299,N_6176);
or U10260 (N_10260,N_8531,N_6871);
or U10261 (N_10261,N_7461,N_7966);
and U10262 (N_10262,N_7419,N_8821);
nor U10263 (N_10263,N_6069,N_7568);
and U10264 (N_10264,N_7954,N_6363);
and U10265 (N_10265,N_8463,N_6572);
or U10266 (N_10266,N_7549,N_6454);
nand U10267 (N_10267,N_8528,N_7730);
nand U10268 (N_10268,N_6357,N_8677);
xor U10269 (N_10269,N_7247,N_7684);
or U10270 (N_10270,N_7643,N_7367);
nor U10271 (N_10271,N_7785,N_6585);
and U10272 (N_10272,N_6820,N_8190);
and U10273 (N_10273,N_8591,N_7344);
and U10274 (N_10274,N_6981,N_7960);
or U10275 (N_10275,N_8447,N_7725);
and U10276 (N_10276,N_7939,N_6975);
and U10277 (N_10277,N_8131,N_8503);
and U10278 (N_10278,N_8270,N_6873);
nand U10279 (N_10279,N_8640,N_6198);
and U10280 (N_10280,N_8834,N_7796);
and U10281 (N_10281,N_6272,N_6107);
or U10282 (N_10282,N_6067,N_6542);
xnor U10283 (N_10283,N_8508,N_6989);
nand U10284 (N_10284,N_7846,N_6556);
and U10285 (N_10285,N_8414,N_7627);
and U10286 (N_10286,N_7144,N_6293);
nor U10287 (N_10287,N_6029,N_7347);
nor U10288 (N_10288,N_6552,N_6727);
or U10289 (N_10289,N_8659,N_6458);
nand U10290 (N_10290,N_8555,N_7293);
xor U10291 (N_10291,N_6134,N_8077);
nor U10292 (N_10292,N_6010,N_6257);
or U10293 (N_10293,N_6024,N_8926);
nor U10294 (N_10294,N_7878,N_8982);
nand U10295 (N_10295,N_7951,N_7907);
nand U10296 (N_10296,N_7756,N_6772);
nand U10297 (N_10297,N_8328,N_7308);
and U10298 (N_10298,N_7275,N_8546);
and U10299 (N_10299,N_8817,N_7372);
or U10300 (N_10300,N_8939,N_6898);
and U10301 (N_10301,N_7316,N_7147);
nand U10302 (N_10302,N_6647,N_6300);
and U10303 (N_10303,N_6466,N_6596);
and U10304 (N_10304,N_7430,N_8902);
nand U10305 (N_10305,N_6348,N_7962);
and U10306 (N_10306,N_8738,N_6937);
and U10307 (N_10307,N_7064,N_7136);
xor U10308 (N_10308,N_6503,N_7799);
and U10309 (N_10309,N_6659,N_6294);
xor U10310 (N_10310,N_8715,N_6086);
nand U10311 (N_10311,N_8527,N_7903);
and U10312 (N_10312,N_7276,N_7917);
nand U10313 (N_10313,N_6612,N_6570);
and U10314 (N_10314,N_8595,N_7601);
nor U10315 (N_10315,N_6617,N_6853);
or U10316 (N_10316,N_6976,N_6148);
or U10317 (N_10317,N_6103,N_6597);
nand U10318 (N_10318,N_6733,N_8329);
or U10319 (N_10319,N_7382,N_7577);
xor U10320 (N_10320,N_6631,N_6978);
or U10321 (N_10321,N_6481,N_8352);
and U10322 (N_10322,N_7979,N_8851);
xnor U10323 (N_10323,N_6601,N_8832);
nand U10324 (N_10324,N_6459,N_7143);
xor U10325 (N_10325,N_7503,N_7826);
or U10326 (N_10326,N_7221,N_6609);
nand U10327 (N_10327,N_6710,N_8637);
or U10328 (N_10328,N_7115,N_7754);
nand U10329 (N_10329,N_7825,N_8126);
nor U10330 (N_10330,N_6345,N_7809);
nor U10331 (N_10331,N_8918,N_8878);
and U10332 (N_10332,N_7074,N_7035);
or U10333 (N_10333,N_6569,N_6380);
and U10334 (N_10334,N_8498,N_6605);
nor U10335 (N_10335,N_8138,N_6865);
or U10336 (N_10336,N_6295,N_6332);
xor U10337 (N_10337,N_6701,N_6979);
nand U10338 (N_10338,N_6043,N_7587);
nor U10339 (N_10339,N_8444,N_7711);
nor U10340 (N_10340,N_8767,N_6834);
nor U10341 (N_10341,N_8136,N_6498);
or U10342 (N_10342,N_6758,N_8006);
or U10343 (N_10343,N_6822,N_6002);
and U10344 (N_10344,N_7443,N_8947);
nor U10345 (N_10345,N_7339,N_6717);
nand U10346 (N_10346,N_8424,N_8861);
or U10347 (N_10347,N_6810,N_7827);
nor U10348 (N_10348,N_6097,N_7139);
xor U10349 (N_10349,N_7321,N_6530);
and U10350 (N_10350,N_7357,N_7964);
or U10351 (N_10351,N_7222,N_6118);
nand U10352 (N_10352,N_6927,N_7797);
and U10353 (N_10353,N_8388,N_7249);
nor U10354 (N_10354,N_8406,N_6382);
nor U10355 (N_10355,N_6328,N_8324);
nor U10356 (N_10356,N_8282,N_6108);
nand U10357 (N_10357,N_8874,N_8895);
or U10358 (N_10358,N_8220,N_8658);
xor U10359 (N_10359,N_8012,N_7808);
nand U10360 (N_10360,N_7298,N_8536);
or U10361 (N_10361,N_7562,N_8598);
nand U10362 (N_10362,N_6285,N_6550);
nor U10363 (N_10363,N_7928,N_6635);
nor U10364 (N_10364,N_8773,N_8688);
nand U10365 (N_10365,N_6431,N_8204);
and U10366 (N_10366,N_7851,N_7986);
or U10367 (N_10367,N_7918,N_8779);
xnor U10368 (N_10368,N_7288,N_6327);
and U10369 (N_10369,N_6547,N_8318);
nor U10370 (N_10370,N_8415,N_7713);
nor U10371 (N_10371,N_7922,N_8732);
xnor U10372 (N_10372,N_8887,N_7258);
nor U10373 (N_10373,N_7365,N_8147);
nor U10374 (N_10374,N_8177,N_6325);
nor U10375 (N_10375,N_6562,N_6131);
nor U10376 (N_10376,N_7844,N_6568);
nand U10377 (N_10377,N_7810,N_6745);
xor U10378 (N_10378,N_8521,N_7760);
nand U10379 (N_10379,N_8333,N_8810);
and U10380 (N_10380,N_7508,N_7649);
nand U10381 (N_10381,N_6054,N_8029);
and U10382 (N_10382,N_7569,N_8376);
nand U10383 (N_10383,N_7882,N_8057);
or U10384 (N_10384,N_7184,N_8522);
nor U10385 (N_10385,N_8359,N_8327);
nor U10386 (N_10386,N_7950,N_6514);
and U10387 (N_10387,N_6269,N_7657);
nand U10388 (N_10388,N_6165,N_7469);
nor U10389 (N_10389,N_7363,N_6206);
nand U10390 (N_10390,N_8968,N_8233);
xor U10391 (N_10391,N_7446,N_7246);
nand U10392 (N_10392,N_6661,N_8009);
and U10393 (N_10393,N_8437,N_8809);
xnor U10394 (N_10394,N_7364,N_6682);
xnor U10395 (N_10395,N_6525,N_7701);
and U10396 (N_10396,N_6703,N_8095);
or U10397 (N_10397,N_8714,N_6804);
xnor U10398 (N_10398,N_8205,N_7454);
nor U10399 (N_10399,N_6349,N_7048);
or U10400 (N_10400,N_6850,N_7207);
nor U10401 (N_10401,N_6287,N_8800);
nor U10402 (N_10402,N_6488,N_8151);
or U10403 (N_10403,N_7037,N_7523);
and U10404 (N_10404,N_6884,N_6013);
xor U10405 (N_10405,N_6942,N_7639);
or U10406 (N_10406,N_6686,N_7538);
and U10407 (N_10407,N_7426,N_6453);
and U10408 (N_10408,N_8519,N_6668);
nor U10409 (N_10409,N_8727,N_8908);
nand U10410 (N_10410,N_8842,N_8180);
nor U10411 (N_10411,N_6367,N_6780);
and U10412 (N_10412,N_7847,N_7219);
nor U10413 (N_10413,N_8228,N_7407);
or U10414 (N_10414,N_7563,N_6809);
and U10415 (N_10415,N_8438,N_7202);
and U10416 (N_10416,N_7822,N_6037);
or U10417 (N_10417,N_6620,N_6643);
and U10418 (N_10418,N_7319,N_8709);
or U10419 (N_10419,N_8608,N_7857);
or U10420 (N_10420,N_8892,N_6370);
or U10421 (N_10421,N_7435,N_7441);
and U10422 (N_10422,N_8988,N_7566);
nand U10423 (N_10423,N_7934,N_7424);
or U10424 (N_10424,N_7556,N_7271);
nor U10425 (N_10425,N_7654,N_7155);
and U10426 (N_10426,N_7624,N_7697);
or U10427 (N_10427,N_6775,N_6970);
and U10428 (N_10428,N_8276,N_6866);
nor U10429 (N_10429,N_8570,N_8315);
nand U10430 (N_10430,N_6673,N_8397);
or U10431 (N_10431,N_6385,N_7659);
nor U10432 (N_10432,N_8215,N_7680);
or U10433 (N_10433,N_8162,N_7084);
xnor U10434 (N_10434,N_8565,N_7802);
nand U10435 (N_10435,N_6092,N_6048);
or U10436 (N_10436,N_6774,N_7091);
or U10437 (N_10437,N_6262,N_6358);
xnor U10438 (N_10438,N_7159,N_6887);
nand U10439 (N_10439,N_8944,N_7919);
or U10440 (N_10440,N_7431,N_7396);
nor U10441 (N_10441,N_6885,N_6355);
or U10442 (N_10442,N_8500,N_6783);
nor U10443 (N_10443,N_7153,N_6229);
or U10444 (N_10444,N_7988,N_8085);
or U10445 (N_10445,N_8685,N_7148);
or U10446 (N_10446,N_7236,N_7094);
and U10447 (N_10447,N_6802,N_6943);
and U10448 (N_10448,N_7403,N_6297);
xnor U10449 (N_10449,N_8252,N_8752);
or U10450 (N_10450,N_8422,N_8133);
nor U10451 (N_10451,N_7744,N_7163);
nor U10452 (N_10452,N_7489,N_8691);
nor U10453 (N_10453,N_8255,N_6862);
xor U10454 (N_10454,N_7001,N_8733);
nand U10455 (N_10455,N_7773,N_7024);
or U10456 (N_10456,N_7387,N_7085);
nor U10457 (N_10457,N_8708,N_7635);
nand U10458 (N_10458,N_7623,N_8457);
and U10459 (N_10459,N_8782,N_6835);
and U10460 (N_10460,N_8994,N_6496);
nor U10461 (N_10461,N_7724,N_7311);
nor U10462 (N_10462,N_8697,N_6891);
nor U10463 (N_10463,N_6845,N_6518);
and U10464 (N_10464,N_8080,N_6844);
and U10465 (N_10465,N_6957,N_7160);
nand U10466 (N_10466,N_7352,N_8261);
xor U10467 (N_10467,N_7681,N_6003);
xnor U10468 (N_10468,N_8022,N_6130);
nand U10469 (N_10469,N_6616,N_6114);
nand U10470 (N_10470,N_6583,N_8811);
nand U10471 (N_10471,N_6469,N_7193);
nor U10472 (N_10472,N_8777,N_6233);
nand U10473 (N_10473,N_8385,N_7305);
or U10474 (N_10474,N_7295,N_7804);
nor U10475 (N_10475,N_7022,N_8008);
nor U10476 (N_10476,N_8831,N_8165);
nand U10477 (N_10477,N_8431,N_7069);
and U10478 (N_10478,N_8612,N_7673);
and U10479 (N_10479,N_7083,N_6977);
nor U10480 (N_10480,N_6096,N_7845);
and U10481 (N_10481,N_8537,N_7618);
or U10482 (N_10482,N_8322,N_8222);
and U10483 (N_10483,N_8314,N_6621);
or U10484 (N_10484,N_6883,N_6641);
nor U10485 (N_10485,N_7746,N_8271);
nor U10486 (N_10486,N_8128,N_7241);
and U10487 (N_10487,N_6709,N_7674);
or U10488 (N_10488,N_6279,N_7183);
nor U10489 (N_10489,N_8462,N_8164);
nand U10490 (N_10490,N_8877,N_8509);
nor U10491 (N_10491,N_8756,N_8466);
nand U10492 (N_10492,N_8170,N_7361);
or U10493 (N_10493,N_6987,N_8564);
nor U10494 (N_10494,N_8370,N_6299);
nand U10495 (N_10495,N_7708,N_6441);
or U10496 (N_10496,N_6602,N_6734);
nand U10497 (N_10497,N_7874,N_8786);
or U10498 (N_10498,N_7832,N_6264);
nand U10499 (N_10499,N_7318,N_8070);
xnor U10500 (N_10500,N_6833,N_7476);
or U10501 (N_10501,N_7025,N_8059);
nor U10502 (N_10502,N_7926,N_6658);
nor U10503 (N_10503,N_6751,N_7543);
nor U10504 (N_10504,N_8125,N_6839);
nor U10505 (N_10505,N_6093,N_8871);
or U10506 (N_10506,N_8542,N_7866);
nand U10507 (N_10507,N_8946,N_6132);
nor U10508 (N_10508,N_7697,N_8039);
or U10509 (N_10509,N_8349,N_8668);
and U10510 (N_10510,N_6280,N_8268);
xnor U10511 (N_10511,N_8806,N_8000);
or U10512 (N_10512,N_8356,N_6727);
and U10513 (N_10513,N_6337,N_7945);
or U10514 (N_10514,N_6195,N_7115);
or U10515 (N_10515,N_6355,N_6894);
or U10516 (N_10516,N_8845,N_8059);
xnor U10517 (N_10517,N_6224,N_6714);
nand U10518 (N_10518,N_7846,N_8977);
and U10519 (N_10519,N_7827,N_7863);
nor U10520 (N_10520,N_6193,N_7973);
or U10521 (N_10521,N_8460,N_8034);
nor U10522 (N_10522,N_8563,N_8458);
or U10523 (N_10523,N_6672,N_6350);
nand U10524 (N_10524,N_8129,N_7354);
nand U10525 (N_10525,N_6334,N_6682);
nor U10526 (N_10526,N_8565,N_6777);
nor U10527 (N_10527,N_8408,N_6536);
or U10528 (N_10528,N_7948,N_6020);
nand U10529 (N_10529,N_6950,N_8892);
or U10530 (N_10530,N_6942,N_7956);
nand U10531 (N_10531,N_7855,N_7006);
or U10532 (N_10532,N_6028,N_8779);
or U10533 (N_10533,N_7388,N_8807);
nor U10534 (N_10534,N_8583,N_8680);
or U10535 (N_10535,N_7497,N_8318);
or U10536 (N_10536,N_7933,N_7948);
nor U10537 (N_10537,N_8899,N_6334);
nand U10538 (N_10538,N_7738,N_6856);
nor U10539 (N_10539,N_7167,N_6030);
nor U10540 (N_10540,N_8014,N_8506);
or U10541 (N_10541,N_8168,N_7734);
nand U10542 (N_10542,N_8348,N_7264);
and U10543 (N_10543,N_7024,N_8114);
and U10544 (N_10544,N_7287,N_7537);
xnor U10545 (N_10545,N_8857,N_7071);
nand U10546 (N_10546,N_6181,N_7739);
nand U10547 (N_10547,N_6868,N_6298);
and U10548 (N_10548,N_8940,N_7027);
and U10549 (N_10549,N_7818,N_7985);
and U10550 (N_10550,N_7397,N_6309);
and U10551 (N_10551,N_6305,N_8334);
nor U10552 (N_10552,N_7139,N_6315);
and U10553 (N_10553,N_7248,N_8188);
nand U10554 (N_10554,N_6278,N_8153);
nand U10555 (N_10555,N_8208,N_6597);
or U10556 (N_10556,N_8721,N_8343);
and U10557 (N_10557,N_6924,N_6476);
xor U10558 (N_10558,N_8406,N_8039);
nor U10559 (N_10559,N_6077,N_6853);
nand U10560 (N_10560,N_8526,N_7552);
and U10561 (N_10561,N_6467,N_8419);
or U10562 (N_10562,N_7937,N_6636);
nand U10563 (N_10563,N_6580,N_6187);
and U10564 (N_10564,N_6312,N_8321);
nor U10565 (N_10565,N_8190,N_6676);
and U10566 (N_10566,N_6277,N_6056);
xnor U10567 (N_10567,N_8983,N_7929);
and U10568 (N_10568,N_6333,N_7536);
and U10569 (N_10569,N_7255,N_7092);
nand U10570 (N_10570,N_7581,N_6179);
nor U10571 (N_10571,N_7257,N_6589);
nor U10572 (N_10572,N_6564,N_8930);
and U10573 (N_10573,N_7647,N_6315);
nand U10574 (N_10574,N_8063,N_8526);
xor U10575 (N_10575,N_6272,N_8811);
nand U10576 (N_10576,N_7991,N_7442);
nor U10577 (N_10577,N_7129,N_8001);
or U10578 (N_10578,N_6443,N_8331);
nor U10579 (N_10579,N_7251,N_8492);
or U10580 (N_10580,N_7522,N_6037);
or U10581 (N_10581,N_8390,N_7906);
or U10582 (N_10582,N_8278,N_6029);
nor U10583 (N_10583,N_6641,N_8749);
and U10584 (N_10584,N_6669,N_6843);
or U10585 (N_10585,N_6371,N_7559);
and U10586 (N_10586,N_6957,N_8384);
nand U10587 (N_10587,N_7924,N_7516);
nor U10588 (N_10588,N_7893,N_7158);
xnor U10589 (N_10589,N_8210,N_7183);
nand U10590 (N_10590,N_7581,N_8933);
or U10591 (N_10591,N_6830,N_8110);
nor U10592 (N_10592,N_8566,N_6384);
nor U10593 (N_10593,N_7878,N_8716);
xnor U10594 (N_10594,N_7266,N_8687);
and U10595 (N_10595,N_6730,N_7716);
nand U10596 (N_10596,N_8157,N_8319);
nor U10597 (N_10597,N_7042,N_7023);
nor U10598 (N_10598,N_7372,N_6023);
nand U10599 (N_10599,N_8270,N_7404);
nor U10600 (N_10600,N_7296,N_7567);
or U10601 (N_10601,N_8980,N_7972);
xor U10602 (N_10602,N_7088,N_6686);
nand U10603 (N_10603,N_7378,N_6407);
nand U10604 (N_10604,N_6442,N_6738);
nand U10605 (N_10605,N_8803,N_7430);
nor U10606 (N_10606,N_6830,N_8486);
or U10607 (N_10607,N_8580,N_6469);
nand U10608 (N_10608,N_6995,N_7258);
xor U10609 (N_10609,N_8654,N_8445);
nor U10610 (N_10610,N_6977,N_6766);
and U10611 (N_10611,N_7362,N_8368);
nor U10612 (N_10612,N_7210,N_7600);
and U10613 (N_10613,N_7237,N_7809);
nand U10614 (N_10614,N_7165,N_8268);
xnor U10615 (N_10615,N_6870,N_7567);
nor U10616 (N_10616,N_6800,N_7975);
nor U10617 (N_10617,N_7411,N_8959);
nor U10618 (N_10618,N_8737,N_7790);
and U10619 (N_10619,N_8008,N_6000);
and U10620 (N_10620,N_8536,N_7915);
or U10621 (N_10621,N_8021,N_7076);
nor U10622 (N_10622,N_8529,N_6801);
and U10623 (N_10623,N_7342,N_6775);
nor U10624 (N_10624,N_8364,N_7751);
or U10625 (N_10625,N_6403,N_8966);
nor U10626 (N_10626,N_8021,N_6490);
xnor U10627 (N_10627,N_7757,N_7807);
and U10628 (N_10628,N_6820,N_8427);
nand U10629 (N_10629,N_7017,N_6068);
nand U10630 (N_10630,N_8773,N_6621);
nand U10631 (N_10631,N_7527,N_8944);
xnor U10632 (N_10632,N_8738,N_8410);
or U10633 (N_10633,N_8948,N_7470);
nor U10634 (N_10634,N_7529,N_7274);
nand U10635 (N_10635,N_6587,N_6631);
or U10636 (N_10636,N_8235,N_8259);
xnor U10637 (N_10637,N_6632,N_8435);
nor U10638 (N_10638,N_8617,N_8152);
nand U10639 (N_10639,N_7408,N_8719);
and U10640 (N_10640,N_7360,N_8062);
and U10641 (N_10641,N_8248,N_7109);
and U10642 (N_10642,N_8313,N_8860);
nand U10643 (N_10643,N_7407,N_8023);
or U10644 (N_10644,N_7782,N_7003);
or U10645 (N_10645,N_7368,N_7030);
nand U10646 (N_10646,N_8218,N_8147);
nand U10647 (N_10647,N_7175,N_6634);
nor U10648 (N_10648,N_8915,N_8094);
and U10649 (N_10649,N_8844,N_8476);
and U10650 (N_10650,N_8125,N_7553);
and U10651 (N_10651,N_8150,N_7817);
or U10652 (N_10652,N_6582,N_6787);
nand U10653 (N_10653,N_6434,N_7587);
and U10654 (N_10654,N_8170,N_6052);
and U10655 (N_10655,N_8242,N_6759);
xor U10656 (N_10656,N_8290,N_6999);
xor U10657 (N_10657,N_7242,N_8905);
or U10658 (N_10658,N_6180,N_7820);
nand U10659 (N_10659,N_7653,N_8641);
and U10660 (N_10660,N_8752,N_6492);
or U10661 (N_10661,N_6511,N_7125);
nor U10662 (N_10662,N_7807,N_8597);
nor U10663 (N_10663,N_8237,N_8846);
and U10664 (N_10664,N_6056,N_7278);
nand U10665 (N_10665,N_7192,N_7562);
nor U10666 (N_10666,N_8922,N_8039);
xor U10667 (N_10667,N_8183,N_8775);
or U10668 (N_10668,N_8504,N_7869);
nand U10669 (N_10669,N_7982,N_6191);
or U10670 (N_10670,N_7020,N_6669);
xnor U10671 (N_10671,N_8273,N_7727);
or U10672 (N_10672,N_7554,N_7661);
and U10673 (N_10673,N_7849,N_6844);
or U10674 (N_10674,N_6264,N_6225);
or U10675 (N_10675,N_7850,N_6240);
and U10676 (N_10676,N_8359,N_7855);
nand U10677 (N_10677,N_8235,N_6880);
nand U10678 (N_10678,N_6844,N_8653);
or U10679 (N_10679,N_8120,N_6122);
xnor U10680 (N_10680,N_7836,N_8978);
xnor U10681 (N_10681,N_8086,N_6038);
or U10682 (N_10682,N_7023,N_6683);
nand U10683 (N_10683,N_6163,N_7239);
xnor U10684 (N_10684,N_7514,N_7927);
and U10685 (N_10685,N_6304,N_6118);
nand U10686 (N_10686,N_8779,N_8299);
xnor U10687 (N_10687,N_8620,N_8855);
nand U10688 (N_10688,N_8882,N_7558);
nor U10689 (N_10689,N_7872,N_8520);
nand U10690 (N_10690,N_6223,N_7606);
or U10691 (N_10691,N_6256,N_7292);
nor U10692 (N_10692,N_6653,N_8021);
nor U10693 (N_10693,N_7403,N_6600);
or U10694 (N_10694,N_8218,N_7117);
nand U10695 (N_10695,N_8358,N_8436);
nor U10696 (N_10696,N_7582,N_6480);
nand U10697 (N_10697,N_8517,N_7451);
nor U10698 (N_10698,N_8676,N_6381);
xor U10699 (N_10699,N_6303,N_6242);
nor U10700 (N_10700,N_8738,N_8810);
nand U10701 (N_10701,N_6104,N_7681);
and U10702 (N_10702,N_7409,N_8425);
nor U10703 (N_10703,N_7244,N_7319);
nor U10704 (N_10704,N_6400,N_8110);
xnor U10705 (N_10705,N_6914,N_7633);
and U10706 (N_10706,N_8851,N_6854);
nand U10707 (N_10707,N_8861,N_8707);
nor U10708 (N_10708,N_7570,N_7611);
and U10709 (N_10709,N_8415,N_8695);
nor U10710 (N_10710,N_8497,N_6832);
nor U10711 (N_10711,N_7409,N_7429);
nand U10712 (N_10712,N_8628,N_6620);
xor U10713 (N_10713,N_6676,N_7116);
nand U10714 (N_10714,N_6143,N_8401);
nand U10715 (N_10715,N_7850,N_6364);
or U10716 (N_10716,N_7491,N_8268);
nor U10717 (N_10717,N_7670,N_8179);
nor U10718 (N_10718,N_6140,N_7371);
and U10719 (N_10719,N_6352,N_8233);
xor U10720 (N_10720,N_6041,N_8243);
or U10721 (N_10721,N_7196,N_7288);
nor U10722 (N_10722,N_6102,N_6122);
and U10723 (N_10723,N_8387,N_6822);
nand U10724 (N_10724,N_6501,N_8543);
and U10725 (N_10725,N_7913,N_6693);
nand U10726 (N_10726,N_7891,N_8837);
and U10727 (N_10727,N_8063,N_6746);
nand U10728 (N_10728,N_7950,N_8412);
nand U10729 (N_10729,N_7911,N_8826);
nor U10730 (N_10730,N_7396,N_6724);
or U10731 (N_10731,N_6121,N_7239);
and U10732 (N_10732,N_6284,N_8361);
and U10733 (N_10733,N_7534,N_7327);
nand U10734 (N_10734,N_7712,N_6764);
or U10735 (N_10735,N_8852,N_8508);
or U10736 (N_10736,N_8833,N_7309);
or U10737 (N_10737,N_6344,N_8611);
xnor U10738 (N_10738,N_7382,N_6296);
xor U10739 (N_10739,N_7524,N_8064);
or U10740 (N_10740,N_8689,N_7473);
and U10741 (N_10741,N_6800,N_8759);
nor U10742 (N_10742,N_8315,N_6505);
nand U10743 (N_10743,N_8810,N_8467);
nand U10744 (N_10744,N_7805,N_7309);
or U10745 (N_10745,N_8853,N_8252);
nand U10746 (N_10746,N_8686,N_6912);
and U10747 (N_10747,N_7770,N_7761);
nor U10748 (N_10748,N_8186,N_7839);
or U10749 (N_10749,N_7451,N_8934);
nand U10750 (N_10750,N_8813,N_8378);
nor U10751 (N_10751,N_6944,N_6798);
or U10752 (N_10752,N_8953,N_7909);
xnor U10753 (N_10753,N_6354,N_8800);
xor U10754 (N_10754,N_7801,N_6498);
xor U10755 (N_10755,N_8189,N_7808);
nor U10756 (N_10756,N_8761,N_8115);
nor U10757 (N_10757,N_8686,N_8988);
or U10758 (N_10758,N_6824,N_8822);
nand U10759 (N_10759,N_8681,N_6752);
nand U10760 (N_10760,N_6602,N_7130);
or U10761 (N_10761,N_7503,N_8788);
and U10762 (N_10762,N_7500,N_6237);
nor U10763 (N_10763,N_8444,N_6455);
nor U10764 (N_10764,N_7132,N_7240);
nand U10765 (N_10765,N_8162,N_8762);
or U10766 (N_10766,N_7089,N_7178);
xor U10767 (N_10767,N_8062,N_8361);
nor U10768 (N_10768,N_7836,N_6951);
and U10769 (N_10769,N_8975,N_8070);
and U10770 (N_10770,N_7378,N_8046);
xnor U10771 (N_10771,N_7250,N_8575);
nor U10772 (N_10772,N_6346,N_7708);
nor U10773 (N_10773,N_7310,N_8943);
nor U10774 (N_10774,N_8056,N_8089);
or U10775 (N_10775,N_8376,N_8766);
nand U10776 (N_10776,N_7865,N_7899);
nand U10777 (N_10777,N_7102,N_6734);
nand U10778 (N_10778,N_7160,N_7127);
nor U10779 (N_10779,N_8759,N_8052);
nor U10780 (N_10780,N_6664,N_7776);
nor U10781 (N_10781,N_8332,N_7458);
nand U10782 (N_10782,N_6723,N_6777);
nand U10783 (N_10783,N_6803,N_7710);
xnor U10784 (N_10784,N_6364,N_7875);
nand U10785 (N_10785,N_7576,N_7474);
nor U10786 (N_10786,N_6446,N_8720);
nand U10787 (N_10787,N_7928,N_7877);
nand U10788 (N_10788,N_8594,N_7078);
nor U10789 (N_10789,N_7293,N_7547);
or U10790 (N_10790,N_6964,N_6697);
or U10791 (N_10791,N_8106,N_8714);
nand U10792 (N_10792,N_7107,N_8684);
nor U10793 (N_10793,N_8330,N_7108);
nor U10794 (N_10794,N_6568,N_6241);
nor U10795 (N_10795,N_7170,N_8667);
nand U10796 (N_10796,N_7604,N_6240);
and U10797 (N_10797,N_6062,N_6235);
and U10798 (N_10798,N_8275,N_6706);
or U10799 (N_10799,N_7486,N_7840);
nor U10800 (N_10800,N_6108,N_6837);
nor U10801 (N_10801,N_8314,N_6182);
and U10802 (N_10802,N_8409,N_7798);
and U10803 (N_10803,N_8312,N_8771);
and U10804 (N_10804,N_7619,N_8889);
nand U10805 (N_10805,N_7912,N_6915);
or U10806 (N_10806,N_6829,N_6679);
nand U10807 (N_10807,N_7152,N_8341);
nand U10808 (N_10808,N_7253,N_8051);
or U10809 (N_10809,N_8876,N_8172);
xor U10810 (N_10810,N_7696,N_6270);
nor U10811 (N_10811,N_7013,N_6513);
or U10812 (N_10812,N_6892,N_6298);
and U10813 (N_10813,N_8800,N_8912);
nor U10814 (N_10814,N_7956,N_7022);
xnor U10815 (N_10815,N_7855,N_7439);
nor U10816 (N_10816,N_8654,N_6834);
or U10817 (N_10817,N_7065,N_6633);
nor U10818 (N_10818,N_8707,N_7903);
nor U10819 (N_10819,N_8937,N_8344);
and U10820 (N_10820,N_8883,N_8740);
or U10821 (N_10821,N_8927,N_6712);
and U10822 (N_10822,N_8074,N_7344);
nand U10823 (N_10823,N_6596,N_6933);
nand U10824 (N_10824,N_7124,N_7282);
nand U10825 (N_10825,N_6060,N_8804);
and U10826 (N_10826,N_6980,N_8825);
nand U10827 (N_10827,N_7902,N_7793);
or U10828 (N_10828,N_7162,N_6610);
and U10829 (N_10829,N_7709,N_8801);
and U10830 (N_10830,N_8927,N_7184);
nand U10831 (N_10831,N_6064,N_8460);
nand U10832 (N_10832,N_8690,N_8111);
and U10833 (N_10833,N_8568,N_6187);
nand U10834 (N_10834,N_6854,N_6649);
or U10835 (N_10835,N_7507,N_6214);
and U10836 (N_10836,N_6030,N_7969);
nand U10837 (N_10837,N_6183,N_8075);
or U10838 (N_10838,N_8367,N_8575);
nand U10839 (N_10839,N_8385,N_8377);
or U10840 (N_10840,N_8551,N_8406);
and U10841 (N_10841,N_7735,N_6076);
or U10842 (N_10842,N_6300,N_8674);
nor U10843 (N_10843,N_6725,N_6510);
or U10844 (N_10844,N_7343,N_7728);
nand U10845 (N_10845,N_7284,N_8368);
nor U10846 (N_10846,N_7880,N_8177);
nor U10847 (N_10847,N_8461,N_6779);
or U10848 (N_10848,N_7571,N_8549);
or U10849 (N_10849,N_7333,N_8509);
nand U10850 (N_10850,N_8631,N_6747);
nand U10851 (N_10851,N_8671,N_8834);
nand U10852 (N_10852,N_6509,N_8569);
or U10853 (N_10853,N_7994,N_6268);
and U10854 (N_10854,N_6759,N_6568);
or U10855 (N_10855,N_8995,N_6623);
xnor U10856 (N_10856,N_7052,N_7614);
or U10857 (N_10857,N_6650,N_6688);
and U10858 (N_10858,N_6437,N_6019);
nand U10859 (N_10859,N_7995,N_7186);
xnor U10860 (N_10860,N_8110,N_7107);
and U10861 (N_10861,N_6936,N_8571);
nor U10862 (N_10862,N_6231,N_6393);
nand U10863 (N_10863,N_8672,N_8292);
or U10864 (N_10864,N_6173,N_7768);
or U10865 (N_10865,N_7003,N_8234);
and U10866 (N_10866,N_7548,N_7092);
nand U10867 (N_10867,N_8011,N_7459);
xnor U10868 (N_10868,N_8660,N_8640);
and U10869 (N_10869,N_6254,N_7963);
nand U10870 (N_10870,N_8210,N_8255);
nand U10871 (N_10871,N_6588,N_6683);
or U10872 (N_10872,N_6717,N_6669);
nand U10873 (N_10873,N_6924,N_8007);
or U10874 (N_10874,N_6509,N_6958);
nand U10875 (N_10875,N_6527,N_8548);
and U10876 (N_10876,N_6637,N_6501);
and U10877 (N_10877,N_6601,N_8980);
or U10878 (N_10878,N_6120,N_6552);
or U10879 (N_10879,N_8174,N_7639);
or U10880 (N_10880,N_7813,N_8856);
and U10881 (N_10881,N_7428,N_8672);
nand U10882 (N_10882,N_8093,N_8048);
nand U10883 (N_10883,N_7256,N_6515);
xor U10884 (N_10884,N_8723,N_7941);
or U10885 (N_10885,N_8991,N_8185);
nor U10886 (N_10886,N_7910,N_7542);
nor U10887 (N_10887,N_8075,N_8426);
nand U10888 (N_10888,N_7367,N_7808);
or U10889 (N_10889,N_6228,N_6084);
nor U10890 (N_10890,N_6325,N_7478);
or U10891 (N_10891,N_6800,N_8012);
nor U10892 (N_10892,N_6495,N_7223);
nor U10893 (N_10893,N_8583,N_8318);
and U10894 (N_10894,N_6549,N_6177);
nand U10895 (N_10895,N_7314,N_8728);
nand U10896 (N_10896,N_8397,N_7931);
and U10897 (N_10897,N_7842,N_6639);
nor U10898 (N_10898,N_7280,N_6566);
nor U10899 (N_10899,N_6866,N_7145);
or U10900 (N_10900,N_6763,N_6624);
xnor U10901 (N_10901,N_6982,N_6592);
nand U10902 (N_10902,N_8241,N_8872);
or U10903 (N_10903,N_6557,N_7145);
nand U10904 (N_10904,N_6615,N_7762);
xor U10905 (N_10905,N_6790,N_7536);
nand U10906 (N_10906,N_7692,N_6141);
nand U10907 (N_10907,N_6574,N_8996);
nor U10908 (N_10908,N_8856,N_8903);
nor U10909 (N_10909,N_7832,N_7717);
or U10910 (N_10910,N_8373,N_8458);
nor U10911 (N_10911,N_6202,N_6950);
or U10912 (N_10912,N_7510,N_6421);
nor U10913 (N_10913,N_8889,N_6425);
nor U10914 (N_10914,N_7728,N_7925);
nand U10915 (N_10915,N_6200,N_6260);
nor U10916 (N_10916,N_7117,N_6446);
nand U10917 (N_10917,N_8551,N_7135);
or U10918 (N_10918,N_8892,N_7777);
or U10919 (N_10919,N_8514,N_7464);
or U10920 (N_10920,N_8145,N_7030);
nand U10921 (N_10921,N_7163,N_8175);
or U10922 (N_10922,N_8799,N_7699);
or U10923 (N_10923,N_8458,N_7831);
or U10924 (N_10924,N_8809,N_6725);
nor U10925 (N_10925,N_6865,N_8948);
and U10926 (N_10926,N_6694,N_7874);
nor U10927 (N_10927,N_7411,N_7729);
xnor U10928 (N_10928,N_7968,N_7488);
nor U10929 (N_10929,N_8713,N_8408);
and U10930 (N_10930,N_8701,N_8793);
and U10931 (N_10931,N_6630,N_6286);
nand U10932 (N_10932,N_7596,N_6047);
or U10933 (N_10933,N_6902,N_7657);
nand U10934 (N_10934,N_8866,N_7792);
nor U10935 (N_10935,N_8107,N_8832);
nand U10936 (N_10936,N_8139,N_7761);
or U10937 (N_10937,N_6765,N_6819);
nand U10938 (N_10938,N_6936,N_7403);
and U10939 (N_10939,N_6953,N_8116);
and U10940 (N_10940,N_8399,N_7333);
nor U10941 (N_10941,N_6654,N_7835);
and U10942 (N_10942,N_7668,N_6549);
nor U10943 (N_10943,N_8133,N_8434);
or U10944 (N_10944,N_7740,N_7938);
nand U10945 (N_10945,N_7298,N_6903);
or U10946 (N_10946,N_8229,N_6674);
nand U10947 (N_10947,N_6835,N_8370);
nor U10948 (N_10948,N_8101,N_7061);
nor U10949 (N_10949,N_6902,N_8571);
and U10950 (N_10950,N_8822,N_8229);
or U10951 (N_10951,N_6767,N_8966);
or U10952 (N_10952,N_6722,N_6979);
nand U10953 (N_10953,N_7699,N_7666);
and U10954 (N_10954,N_6626,N_8811);
and U10955 (N_10955,N_7174,N_7233);
or U10956 (N_10956,N_7590,N_8751);
and U10957 (N_10957,N_7419,N_8160);
nand U10958 (N_10958,N_6462,N_7753);
nor U10959 (N_10959,N_7922,N_8417);
xnor U10960 (N_10960,N_8480,N_7411);
and U10961 (N_10961,N_7313,N_7996);
and U10962 (N_10962,N_6712,N_8793);
or U10963 (N_10963,N_7799,N_7772);
and U10964 (N_10964,N_7257,N_6118);
nor U10965 (N_10965,N_7438,N_6519);
or U10966 (N_10966,N_7377,N_6607);
nand U10967 (N_10967,N_8711,N_8884);
xnor U10968 (N_10968,N_8272,N_7565);
nor U10969 (N_10969,N_6541,N_6444);
nor U10970 (N_10970,N_6380,N_6906);
and U10971 (N_10971,N_8563,N_6113);
and U10972 (N_10972,N_8523,N_7711);
nor U10973 (N_10973,N_6482,N_7938);
nand U10974 (N_10974,N_8970,N_8913);
nand U10975 (N_10975,N_7260,N_6857);
nor U10976 (N_10976,N_6715,N_7956);
nand U10977 (N_10977,N_7536,N_6386);
or U10978 (N_10978,N_6040,N_7018);
nand U10979 (N_10979,N_8759,N_8752);
nand U10980 (N_10980,N_6635,N_7487);
or U10981 (N_10981,N_8990,N_6931);
or U10982 (N_10982,N_7956,N_8651);
and U10983 (N_10983,N_6402,N_8126);
and U10984 (N_10984,N_7280,N_7837);
nor U10985 (N_10985,N_7245,N_6866);
nor U10986 (N_10986,N_6141,N_6370);
or U10987 (N_10987,N_6812,N_6607);
xnor U10988 (N_10988,N_8160,N_6652);
nor U10989 (N_10989,N_8315,N_8103);
and U10990 (N_10990,N_8614,N_6991);
nor U10991 (N_10991,N_8983,N_8590);
nor U10992 (N_10992,N_6124,N_8603);
nor U10993 (N_10993,N_8239,N_8191);
or U10994 (N_10994,N_6127,N_6294);
and U10995 (N_10995,N_8489,N_6724);
nor U10996 (N_10996,N_6168,N_8297);
and U10997 (N_10997,N_6379,N_7433);
nor U10998 (N_10998,N_8432,N_7415);
xor U10999 (N_10999,N_6761,N_7326);
or U11000 (N_11000,N_7487,N_6443);
nor U11001 (N_11001,N_8855,N_8061);
or U11002 (N_11002,N_7581,N_8225);
or U11003 (N_11003,N_8017,N_7084);
and U11004 (N_11004,N_6816,N_8956);
nand U11005 (N_11005,N_7196,N_6711);
and U11006 (N_11006,N_6294,N_7796);
nor U11007 (N_11007,N_7231,N_6236);
and U11008 (N_11008,N_6606,N_6688);
nand U11009 (N_11009,N_8806,N_7705);
and U11010 (N_11010,N_8286,N_8222);
or U11011 (N_11011,N_8618,N_7829);
and U11012 (N_11012,N_7169,N_6751);
or U11013 (N_11013,N_8986,N_8109);
and U11014 (N_11014,N_7654,N_7546);
nor U11015 (N_11015,N_8133,N_7276);
nor U11016 (N_11016,N_8297,N_7703);
nor U11017 (N_11017,N_8096,N_8151);
and U11018 (N_11018,N_8538,N_8680);
or U11019 (N_11019,N_6569,N_6959);
nand U11020 (N_11020,N_6256,N_7152);
and U11021 (N_11021,N_7747,N_6937);
or U11022 (N_11022,N_7563,N_6173);
nor U11023 (N_11023,N_7363,N_6344);
and U11024 (N_11024,N_6544,N_8944);
nand U11025 (N_11025,N_6126,N_6247);
nor U11026 (N_11026,N_7051,N_8321);
nor U11027 (N_11027,N_8097,N_6720);
or U11028 (N_11028,N_7136,N_7984);
nor U11029 (N_11029,N_7834,N_8411);
nor U11030 (N_11030,N_8259,N_8144);
and U11031 (N_11031,N_8007,N_6043);
or U11032 (N_11032,N_6105,N_7055);
nor U11033 (N_11033,N_6695,N_6715);
and U11034 (N_11034,N_6634,N_6320);
and U11035 (N_11035,N_8514,N_6879);
nand U11036 (N_11036,N_7792,N_8824);
nand U11037 (N_11037,N_6281,N_8828);
or U11038 (N_11038,N_6604,N_8306);
nor U11039 (N_11039,N_7015,N_6467);
or U11040 (N_11040,N_8618,N_7400);
nor U11041 (N_11041,N_8026,N_6549);
or U11042 (N_11042,N_7427,N_7777);
nand U11043 (N_11043,N_8764,N_7331);
nor U11044 (N_11044,N_7945,N_6043);
and U11045 (N_11045,N_7327,N_7727);
or U11046 (N_11046,N_6119,N_8591);
or U11047 (N_11047,N_8756,N_8788);
nor U11048 (N_11048,N_6641,N_6056);
nand U11049 (N_11049,N_6805,N_7142);
xor U11050 (N_11050,N_6460,N_7981);
or U11051 (N_11051,N_8671,N_6028);
or U11052 (N_11052,N_7968,N_8100);
and U11053 (N_11053,N_7786,N_6766);
nand U11054 (N_11054,N_8923,N_8265);
nor U11055 (N_11055,N_6660,N_6965);
or U11056 (N_11056,N_6013,N_6323);
nand U11057 (N_11057,N_7620,N_7920);
nand U11058 (N_11058,N_8463,N_6703);
and U11059 (N_11059,N_6454,N_8497);
or U11060 (N_11060,N_8002,N_7304);
xnor U11061 (N_11061,N_6252,N_7311);
nand U11062 (N_11062,N_6417,N_6378);
and U11063 (N_11063,N_7531,N_8493);
nand U11064 (N_11064,N_6796,N_8976);
and U11065 (N_11065,N_8695,N_6630);
nor U11066 (N_11066,N_8808,N_6465);
nor U11067 (N_11067,N_8120,N_7052);
nor U11068 (N_11068,N_8047,N_8727);
and U11069 (N_11069,N_8742,N_8366);
or U11070 (N_11070,N_7418,N_8004);
and U11071 (N_11071,N_6554,N_6076);
nor U11072 (N_11072,N_7154,N_6647);
nand U11073 (N_11073,N_6161,N_8312);
and U11074 (N_11074,N_8997,N_7436);
nand U11075 (N_11075,N_8032,N_6937);
nor U11076 (N_11076,N_6453,N_8279);
or U11077 (N_11077,N_6556,N_8727);
and U11078 (N_11078,N_8657,N_6829);
or U11079 (N_11079,N_7599,N_6546);
nor U11080 (N_11080,N_7211,N_6853);
nand U11081 (N_11081,N_6565,N_8846);
nor U11082 (N_11082,N_7036,N_8288);
and U11083 (N_11083,N_8185,N_7676);
nand U11084 (N_11084,N_8863,N_6333);
nor U11085 (N_11085,N_7467,N_6659);
and U11086 (N_11086,N_6088,N_7259);
and U11087 (N_11087,N_7675,N_7650);
or U11088 (N_11088,N_7720,N_8545);
nor U11089 (N_11089,N_6480,N_8994);
nand U11090 (N_11090,N_7591,N_6696);
nand U11091 (N_11091,N_6563,N_6327);
nand U11092 (N_11092,N_8606,N_6718);
xnor U11093 (N_11093,N_8807,N_8777);
nor U11094 (N_11094,N_6767,N_7577);
xor U11095 (N_11095,N_8373,N_6175);
nor U11096 (N_11096,N_8305,N_8736);
nand U11097 (N_11097,N_7731,N_7141);
nand U11098 (N_11098,N_8961,N_6679);
nand U11099 (N_11099,N_6637,N_8964);
or U11100 (N_11100,N_8491,N_8118);
and U11101 (N_11101,N_6125,N_6516);
nor U11102 (N_11102,N_8974,N_6654);
nand U11103 (N_11103,N_8923,N_8380);
nor U11104 (N_11104,N_6895,N_6627);
nor U11105 (N_11105,N_7855,N_6558);
and U11106 (N_11106,N_6323,N_8881);
and U11107 (N_11107,N_8121,N_6309);
and U11108 (N_11108,N_7817,N_8399);
nand U11109 (N_11109,N_8520,N_7023);
and U11110 (N_11110,N_6137,N_7107);
nor U11111 (N_11111,N_8909,N_7064);
or U11112 (N_11112,N_8877,N_7970);
nand U11113 (N_11113,N_7625,N_6949);
nand U11114 (N_11114,N_6804,N_6045);
nor U11115 (N_11115,N_7513,N_7220);
and U11116 (N_11116,N_8626,N_8511);
xnor U11117 (N_11117,N_8223,N_7220);
nor U11118 (N_11118,N_7751,N_7748);
or U11119 (N_11119,N_6346,N_6915);
and U11120 (N_11120,N_8557,N_7138);
nor U11121 (N_11121,N_7693,N_6648);
or U11122 (N_11122,N_6783,N_7050);
nand U11123 (N_11123,N_7766,N_8218);
nor U11124 (N_11124,N_6491,N_6972);
xnor U11125 (N_11125,N_8945,N_6935);
and U11126 (N_11126,N_6138,N_8752);
and U11127 (N_11127,N_8413,N_7740);
nor U11128 (N_11128,N_8267,N_6701);
nor U11129 (N_11129,N_7554,N_7343);
and U11130 (N_11130,N_6459,N_8618);
nor U11131 (N_11131,N_8583,N_7520);
or U11132 (N_11132,N_7235,N_8397);
nor U11133 (N_11133,N_6395,N_8360);
or U11134 (N_11134,N_7726,N_6537);
and U11135 (N_11135,N_6087,N_8722);
and U11136 (N_11136,N_7082,N_8675);
and U11137 (N_11137,N_6054,N_7115);
and U11138 (N_11138,N_8687,N_6103);
or U11139 (N_11139,N_7825,N_7759);
and U11140 (N_11140,N_7759,N_6354);
and U11141 (N_11141,N_7762,N_8697);
or U11142 (N_11142,N_7760,N_8955);
nor U11143 (N_11143,N_8032,N_6198);
nand U11144 (N_11144,N_6197,N_6406);
or U11145 (N_11145,N_8414,N_7784);
or U11146 (N_11146,N_6842,N_8271);
nor U11147 (N_11147,N_6305,N_6251);
or U11148 (N_11148,N_6314,N_6702);
or U11149 (N_11149,N_8826,N_8926);
nor U11150 (N_11150,N_6970,N_8620);
nand U11151 (N_11151,N_6486,N_7946);
and U11152 (N_11152,N_6892,N_6085);
nand U11153 (N_11153,N_8049,N_6864);
nor U11154 (N_11154,N_8157,N_7103);
and U11155 (N_11155,N_6253,N_8860);
or U11156 (N_11156,N_7117,N_7716);
or U11157 (N_11157,N_6321,N_6595);
and U11158 (N_11158,N_6103,N_7618);
and U11159 (N_11159,N_6263,N_8615);
xnor U11160 (N_11160,N_8915,N_8969);
nor U11161 (N_11161,N_6869,N_7759);
and U11162 (N_11162,N_6375,N_8693);
or U11163 (N_11163,N_6029,N_6329);
or U11164 (N_11164,N_7625,N_8338);
or U11165 (N_11165,N_8150,N_8456);
nor U11166 (N_11166,N_8183,N_6932);
xor U11167 (N_11167,N_6352,N_8201);
nand U11168 (N_11168,N_6575,N_8535);
nand U11169 (N_11169,N_8267,N_8536);
nor U11170 (N_11170,N_8033,N_8097);
and U11171 (N_11171,N_6438,N_8987);
nor U11172 (N_11172,N_7124,N_8836);
and U11173 (N_11173,N_8529,N_6397);
nand U11174 (N_11174,N_6243,N_8999);
or U11175 (N_11175,N_7713,N_8015);
and U11176 (N_11176,N_7850,N_6969);
or U11177 (N_11177,N_8286,N_7735);
or U11178 (N_11178,N_6582,N_7794);
nor U11179 (N_11179,N_8305,N_8235);
xnor U11180 (N_11180,N_8320,N_7140);
and U11181 (N_11181,N_7685,N_7274);
nand U11182 (N_11182,N_7288,N_8049);
nor U11183 (N_11183,N_8116,N_8956);
nor U11184 (N_11184,N_6540,N_7727);
nand U11185 (N_11185,N_7796,N_8302);
and U11186 (N_11186,N_8971,N_7966);
and U11187 (N_11187,N_7635,N_7413);
or U11188 (N_11188,N_6920,N_7030);
or U11189 (N_11189,N_6170,N_6575);
or U11190 (N_11190,N_6089,N_6003);
or U11191 (N_11191,N_6310,N_8591);
and U11192 (N_11192,N_8142,N_7940);
nand U11193 (N_11193,N_6007,N_7633);
or U11194 (N_11194,N_7174,N_6234);
nand U11195 (N_11195,N_7762,N_8400);
or U11196 (N_11196,N_8031,N_6572);
or U11197 (N_11197,N_6734,N_7592);
nor U11198 (N_11198,N_7904,N_6958);
or U11199 (N_11199,N_6564,N_7086);
or U11200 (N_11200,N_7412,N_8847);
nor U11201 (N_11201,N_8401,N_8649);
nor U11202 (N_11202,N_6948,N_6911);
or U11203 (N_11203,N_7892,N_7137);
xor U11204 (N_11204,N_7841,N_7132);
or U11205 (N_11205,N_8140,N_6228);
xor U11206 (N_11206,N_6300,N_7000);
and U11207 (N_11207,N_8313,N_6977);
and U11208 (N_11208,N_6985,N_8754);
or U11209 (N_11209,N_7330,N_6297);
nor U11210 (N_11210,N_8127,N_8274);
and U11211 (N_11211,N_8343,N_6561);
or U11212 (N_11212,N_7739,N_6959);
nand U11213 (N_11213,N_7468,N_6806);
nand U11214 (N_11214,N_7231,N_7855);
nand U11215 (N_11215,N_8813,N_7595);
and U11216 (N_11216,N_6280,N_6934);
nand U11217 (N_11217,N_7872,N_8799);
nor U11218 (N_11218,N_7548,N_6695);
nand U11219 (N_11219,N_8472,N_8649);
nor U11220 (N_11220,N_8367,N_8596);
nor U11221 (N_11221,N_8776,N_8108);
and U11222 (N_11222,N_6750,N_6293);
nand U11223 (N_11223,N_6278,N_6471);
xnor U11224 (N_11224,N_7661,N_6226);
nand U11225 (N_11225,N_8999,N_6335);
and U11226 (N_11226,N_6619,N_6841);
or U11227 (N_11227,N_7115,N_8748);
nor U11228 (N_11228,N_6204,N_7944);
and U11229 (N_11229,N_6265,N_6872);
nand U11230 (N_11230,N_6189,N_7080);
nor U11231 (N_11231,N_6016,N_8524);
or U11232 (N_11232,N_7172,N_8714);
and U11233 (N_11233,N_8876,N_6533);
or U11234 (N_11234,N_7090,N_8726);
or U11235 (N_11235,N_8053,N_7458);
nor U11236 (N_11236,N_7646,N_7975);
nor U11237 (N_11237,N_6360,N_8758);
nor U11238 (N_11238,N_8634,N_8735);
and U11239 (N_11239,N_8861,N_8517);
or U11240 (N_11240,N_7622,N_8732);
or U11241 (N_11241,N_7616,N_6360);
xnor U11242 (N_11242,N_7229,N_6578);
and U11243 (N_11243,N_7862,N_8779);
nand U11244 (N_11244,N_7688,N_6177);
or U11245 (N_11245,N_7802,N_8163);
and U11246 (N_11246,N_6787,N_7848);
nor U11247 (N_11247,N_8327,N_8654);
nor U11248 (N_11248,N_8549,N_7555);
nor U11249 (N_11249,N_7728,N_8359);
or U11250 (N_11250,N_7698,N_8279);
or U11251 (N_11251,N_6054,N_8808);
and U11252 (N_11252,N_6046,N_8099);
or U11253 (N_11253,N_8589,N_8007);
and U11254 (N_11254,N_8253,N_6908);
and U11255 (N_11255,N_6679,N_8663);
nor U11256 (N_11256,N_6716,N_7984);
and U11257 (N_11257,N_8352,N_7422);
and U11258 (N_11258,N_6160,N_8236);
or U11259 (N_11259,N_8816,N_8881);
or U11260 (N_11260,N_8266,N_7174);
and U11261 (N_11261,N_6054,N_7949);
and U11262 (N_11262,N_7999,N_7360);
and U11263 (N_11263,N_8469,N_8314);
and U11264 (N_11264,N_6163,N_7376);
xor U11265 (N_11265,N_6630,N_7331);
and U11266 (N_11266,N_8627,N_7703);
nand U11267 (N_11267,N_6126,N_8280);
and U11268 (N_11268,N_7287,N_7908);
nand U11269 (N_11269,N_6685,N_6715);
nand U11270 (N_11270,N_6104,N_6790);
nor U11271 (N_11271,N_6070,N_7443);
nand U11272 (N_11272,N_6953,N_8630);
nor U11273 (N_11273,N_8612,N_7870);
nand U11274 (N_11274,N_6006,N_8491);
or U11275 (N_11275,N_8824,N_6024);
xor U11276 (N_11276,N_7669,N_6849);
nand U11277 (N_11277,N_6333,N_8285);
or U11278 (N_11278,N_8038,N_6324);
nor U11279 (N_11279,N_8065,N_8559);
and U11280 (N_11280,N_7738,N_6474);
or U11281 (N_11281,N_7200,N_8105);
and U11282 (N_11282,N_6228,N_8812);
nor U11283 (N_11283,N_7519,N_6518);
nor U11284 (N_11284,N_6926,N_7467);
nand U11285 (N_11285,N_8130,N_6621);
xor U11286 (N_11286,N_8426,N_8458);
xnor U11287 (N_11287,N_8409,N_7139);
and U11288 (N_11288,N_8508,N_7791);
or U11289 (N_11289,N_6378,N_7417);
nor U11290 (N_11290,N_8482,N_6273);
xor U11291 (N_11291,N_8712,N_8923);
nand U11292 (N_11292,N_6588,N_7410);
and U11293 (N_11293,N_6217,N_7843);
nor U11294 (N_11294,N_8777,N_7877);
nor U11295 (N_11295,N_8880,N_8001);
xor U11296 (N_11296,N_6120,N_6309);
nor U11297 (N_11297,N_7856,N_7461);
or U11298 (N_11298,N_8186,N_7182);
or U11299 (N_11299,N_6983,N_7899);
nand U11300 (N_11300,N_8205,N_8516);
nor U11301 (N_11301,N_8562,N_6092);
or U11302 (N_11302,N_6629,N_8886);
nand U11303 (N_11303,N_7443,N_8406);
and U11304 (N_11304,N_8400,N_8843);
xor U11305 (N_11305,N_6551,N_6334);
or U11306 (N_11306,N_6769,N_8073);
and U11307 (N_11307,N_7316,N_7305);
and U11308 (N_11308,N_8269,N_8997);
and U11309 (N_11309,N_6067,N_7828);
nand U11310 (N_11310,N_8224,N_6515);
nand U11311 (N_11311,N_7574,N_8978);
or U11312 (N_11312,N_7060,N_8048);
xor U11313 (N_11313,N_6228,N_8151);
nand U11314 (N_11314,N_8448,N_7365);
and U11315 (N_11315,N_6641,N_6465);
and U11316 (N_11316,N_8475,N_6188);
nor U11317 (N_11317,N_8051,N_7082);
nand U11318 (N_11318,N_6441,N_6743);
or U11319 (N_11319,N_8791,N_7644);
and U11320 (N_11320,N_8936,N_7863);
or U11321 (N_11321,N_7334,N_7512);
and U11322 (N_11322,N_6024,N_7562);
xnor U11323 (N_11323,N_7939,N_6103);
and U11324 (N_11324,N_6708,N_6893);
nor U11325 (N_11325,N_6734,N_7912);
or U11326 (N_11326,N_7246,N_7461);
and U11327 (N_11327,N_6333,N_6034);
nand U11328 (N_11328,N_6754,N_6639);
nand U11329 (N_11329,N_8375,N_7491);
xnor U11330 (N_11330,N_7830,N_6192);
xor U11331 (N_11331,N_6816,N_7808);
nor U11332 (N_11332,N_7099,N_8614);
and U11333 (N_11333,N_8566,N_8760);
and U11334 (N_11334,N_6526,N_6527);
nand U11335 (N_11335,N_6323,N_7366);
and U11336 (N_11336,N_8012,N_8093);
or U11337 (N_11337,N_8753,N_7397);
and U11338 (N_11338,N_8259,N_7773);
nor U11339 (N_11339,N_7585,N_8143);
nand U11340 (N_11340,N_6337,N_7757);
and U11341 (N_11341,N_8038,N_8876);
or U11342 (N_11342,N_6608,N_6286);
nand U11343 (N_11343,N_8906,N_6618);
or U11344 (N_11344,N_6501,N_8350);
or U11345 (N_11345,N_7768,N_8555);
and U11346 (N_11346,N_7680,N_7326);
and U11347 (N_11347,N_6099,N_7435);
nor U11348 (N_11348,N_7165,N_7989);
and U11349 (N_11349,N_7101,N_7032);
nand U11350 (N_11350,N_6019,N_8872);
nor U11351 (N_11351,N_6116,N_6343);
nand U11352 (N_11352,N_6266,N_7296);
and U11353 (N_11353,N_7595,N_8175);
and U11354 (N_11354,N_6232,N_6153);
nor U11355 (N_11355,N_8550,N_8423);
or U11356 (N_11356,N_6609,N_7753);
nand U11357 (N_11357,N_7584,N_6788);
and U11358 (N_11358,N_6901,N_7186);
or U11359 (N_11359,N_6271,N_6876);
or U11360 (N_11360,N_6226,N_7411);
or U11361 (N_11361,N_8423,N_6774);
nand U11362 (N_11362,N_6965,N_7550);
nor U11363 (N_11363,N_8605,N_8516);
nor U11364 (N_11364,N_7773,N_8737);
or U11365 (N_11365,N_6370,N_7027);
nand U11366 (N_11366,N_7017,N_8101);
nand U11367 (N_11367,N_6872,N_6136);
xor U11368 (N_11368,N_7315,N_8313);
nand U11369 (N_11369,N_6080,N_6318);
nand U11370 (N_11370,N_8795,N_7294);
or U11371 (N_11371,N_8098,N_8848);
and U11372 (N_11372,N_6494,N_7847);
and U11373 (N_11373,N_8953,N_7538);
or U11374 (N_11374,N_8780,N_8534);
and U11375 (N_11375,N_6380,N_7319);
nand U11376 (N_11376,N_6667,N_6086);
nand U11377 (N_11377,N_7730,N_8918);
or U11378 (N_11378,N_8112,N_6612);
nand U11379 (N_11379,N_8160,N_8689);
and U11380 (N_11380,N_7936,N_7966);
nor U11381 (N_11381,N_7464,N_8498);
nand U11382 (N_11382,N_8709,N_6253);
or U11383 (N_11383,N_7747,N_6973);
or U11384 (N_11384,N_6161,N_6913);
nor U11385 (N_11385,N_6265,N_7235);
nor U11386 (N_11386,N_6754,N_6473);
or U11387 (N_11387,N_7191,N_6546);
or U11388 (N_11388,N_6944,N_6212);
or U11389 (N_11389,N_6734,N_7090);
nor U11390 (N_11390,N_7958,N_8462);
and U11391 (N_11391,N_8743,N_6784);
nand U11392 (N_11392,N_8068,N_8450);
nor U11393 (N_11393,N_7926,N_7228);
and U11394 (N_11394,N_8306,N_7525);
or U11395 (N_11395,N_8366,N_8854);
and U11396 (N_11396,N_7594,N_6261);
nand U11397 (N_11397,N_8064,N_8588);
or U11398 (N_11398,N_8122,N_7373);
nand U11399 (N_11399,N_7089,N_6483);
nand U11400 (N_11400,N_6533,N_7983);
xnor U11401 (N_11401,N_6753,N_6308);
or U11402 (N_11402,N_8120,N_6747);
nand U11403 (N_11403,N_6805,N_6437);
nor U11404 (N_11404,N_7377,N_6337);
and U11405 (N_11405,N_8394,N_7465);
and U11406 (N_11406,N_7579,N_7999);
xnor U11407 (N_11407,N_7726,N_8631);
nor U11408 (N_11408,N_7742,N_7547);
nor U11409 (N_11409,N_7987,N_6887);
or U11410 (N_11410,N_8540,N_7414);
nor U11411 (N_11411,N_6203,N_7279);
nor U11412 (N_11412,N_7714,N_6732);
and U11413 (N_11413,N_8585,N_8763);
nor U11414 (N_11414,N_8286,N_6044);
xnor U11415 (N_11415,N_7845,N_8588);
and U11416 (N_11416,N_6459,N_6698);
and U11417 (N_11417,N_6684,N_7627);
xnor U11418 (N_11418,N_8078,N_7193);
and U11419 (N_11419,N_8321,N_8757);
nor U11420 (N_11420,N_8211,N_6264);
nor U11421 (N_11421,N_7412,N_8624);
or U11422 (N_11422,N_7758,N_8927);
nand U11423 (N_11423,N_7837,N_8475);
and U11424 (N_11424,N_8325,N_6789);
nor U11425 (N_11425,N_7237,N_8290);
and U11426 (N_11426,N_7174,N_8639);
nor U11427 (N_11427,N_7077,N_6337);
nor U11428 (N_11428,N_8519,N_8310);
or U11429 (N_11429,N_6686,N_7914);
xnor U11430 (N_11430,N_8158,N_8661);
xor U11431 (N_11431,N_6568,N_8146);
or U11432 (N_11432,N_8586,N_6314);
nand U11433 (N_11433,N_8329,N_6775);
nand U11434 (N_11434,N_8906,N_8398);
nor U11435 (N_11435,N_7915,N_7157);
or U11436 (N_11436,N_8353,N_8758);
or U11437 (N_11437,N_8819,N_8736);
nand U11438 (N_11438,N_7482,N_8752);
and U11439 (N_11439,N_7574,N_8173);
or U11440 (N_11440,N_8843,N_8784);
nand U11441 (N_11441,N_6941,N_8202);
or U11442 (N_11442,N_7509,N_8695);
nor U11443 (N_11443,N_7459,N_6141);
or U11444 (N_11444,N_7863,N_6932);
or U11445 (N_11445,N_6844,N_7318);
nor U11446 (N_11446,N_8183,N_6864);
nand U11447 (N_11447,N_6587,N_8106);
and U11448 (N_11448,N_6612,N_6679);
nand U11449 (N_11449,N_8045,N_7123);
nand U11450 (N_11450,N_8885,N_7865);
nor U11451 (N_11451,N_6768,N_7140);
nand U11452 (N_11452,N_7112,N_6919);
nand U11453 (N_11453,N_6365,N_6798);
or U11454 (N_11454,N_6643,N_6982);
nor U11455 (N_11455,N_6472,N_8026);
and U11456 (N_11456,N_7496,N_8387);
or U11457 (N_11457,N_6006,N_6855);
nor U11458 (N_11458,N_7984,N_7767);
and U11459 (N_11459,N_7648,N_6094);
xor U11460 (N_11460,N_8542,N_6019);
nand U11461 (N_11461,N_7257,N_6774);
or U11462 (N_11462,N_6211,N_6288);
or U11463 (N_11463,N_7548,N_7572);
nor U11464 (N_11464,N_6372,N_7498);
and U11465 (N_11465,N_7049,N_7998);
nand U11466 (N_11466,N_6869,N_6603);
nand U11467 (N_11467,N_7144,N_7510);
nor U11468 (N_11468,N_8143,N_8514);
nand U11469 (N_11469,N_8215,N_6919);
nor U11470 (N_11470,N_6558,N_7908);
nor U11471 (N_11471,N_6418,N_8017);
nor U11472 (N_11472,N_7873,N_7009);
and U11473 (N_11473,N_8551,N_8702);
or U11474 (N_11474,N_6969,N_7917);
nor U11475 (N_11475,N_6038,N_7820);
and U11476 (N_11476,N_8440,N_6872);
nor U11477 (N_11477,N_6590,N_7525);
or U11478 (N_11478,N_8851,N_7643);
or U11479 (N_11479,N_6437,N_8882);
nor U11480 (N_11480,N_6989,N_8480);
nor U11481 (N_11481,N_6510,N_6048);
nand U11482 (N_11482,N_8257,N_8805);
or U11483 (N_11483,N_6004,N_7370);
and U11484 (N_11484,N_7834,N_6659);
and U11485 (N_11485,N_8848,N_8011);
or U11486 (N_11486,N_7383,N_7568);
nand U11487 (N_11487,N_8414,N_6233);
nor U11488 (N_11488,N_6683,N_8748);
nor U11489 (N_11489,N_8144,N_6856);
and U11490 (N_11490,N_7696,N_6980);
or U11491 (N_11491,N_7435,N_6777);
or U11492 (N_11492,N_8073,N_6279);
and U11493 (N_11493,N_8925,N_6968);
nand U11494 (N_11494,N_8548,N_6244);
nand U11495 (N_11495,N_8791,N_8383);
nand U11496 (N_11496,N_6022,N_6441);
and U11497 (N_11497,N_7602,N_6003);
nor U11498 (N_11498,N_8796,N_6079);
nand U11499 (N_11499,N_6000,N_8097);
nor U11500 (N_11500,N_8640,N_7105);
and U11501 (N_11501,N_6571,N_6231);
or U11502 (N_11502,N_6696,N_8572);
or U11503 (N_11503,N_8174,N_8090);
nand U11504 (N_11504,N_8749,N_8497);
nor U11505 (N_11505,N_6033,N_8633);
nor U11506 (N_11506,N_6616,N_7213);
or U11507 (N_11507,N_7423,N_6386);
or U11508 (N_11508,N_7145,N_7023);
nor U11509 (N_11509,N_6078,N_6955);
or U11510 (N_11510,N_6738,N_8719);
or U11511 (N_11511,N_6560,N_6815);
xor U11512 (N_11512,N_8480,N_6714);
and U11513 (N_11513,N_7442,N_8354);
and U11514 (N_11514,N_7287,N_7828);
nand U11515 (N_11515,N_7310,N_8006);
and U11516 (N_11516,N_7653,N_6987);
or U11517 (N_11517,N_8079,N_7384);
or U11518 (N_11518,N_6833,N_7889);
nor U11519 (N_11519,N_7255,N_7815);
and U11520 (N_11520,N_7708,N_7575);
or U11521 (N_11521,N_8577,N_7700);
and U11522 (N_11522,N_7730,N_6881);
xor U11523 (N_11523,N_7487,N_7352);
nor U11524 (N_11524,N_6017,N_8611);
nand U11525 (N_11525,N_7161,N_7024);
nor U11526 (N_11526,N_6809,N_7244);
nand U11527 (N_11527,N_6979,N_7526);
nor U11528 (N_11528,N_6571,N_8535);
or U11529 (N_11529,N_7691,N_6230);
and U11530 (N_11530,N_6265,N_7655);
nor U11531 (N_11531,N_6886,N_7241);
nand U11532 (N_11532,N_6510,N_8186);
nor U11533 (N_11533,N_7794,N_7765);
and U11534 (N_11534,N_7131,N_7281);
or U11535 (N_11535,N_8216,N_7522);
xor U11536 (N_11536,N_8382,N_6070);
nor U11537 (N_11537,N_7335,N_6818);
nand U11538 (N_11538,N_8064,N_8862);
nand U11539 (N_11539,N_6185,N_7364);
xor U11540 (N_11540,N_8230,N_7123);
and U11541 (N_11541,N_7113,N_7443);
xor U11542 (N_11542,N_6592,N_8378);
and U11543 (N_11543,N_7533,N_6458);
or U11544 (N_11544,N_7368,N_6855);
or U11545 (N_11545,N_6568,N_8628);
or U11546 (N_11546,N_7991,N_7684);
and U11547 (N_11547,N_7294,N_8337);
and U11548 (N_11548,N_8796,N_6378);
xor U11549 (N_11549,N_7085,N_6328);
nand U11550 (N_11550,N_7545,N_6726);
nor U11551 (N_11551,N_8839,N_8262);
and U11552 (N_11552,N_8312,N_6700);
or U11553 (N_11553,N_7644,N_8843);
nand U11554 (N_11554,N_8271,N_8262);
or U11555 (N_11555,N_8155,N_6150);
and U11556 (N_11556,N_7046,N_7239);
or U11557 (N_11557,N_7419,N_8094);
and U11558 (N_11558,N_8621,N_7586);
or U11559 (N_11559,N_6105,N_7965);
or U11560 (N_11560,N_6194,N_8315);
nand U11561 (N_11561,N_8429,N_7889);
nor U11562 (N_11562,N_7884,N_7542);
nor U11563 (N_11563,N_6016,N_8902);
and U11564 (N_11564,N_6737,N_6999);
and U11565 (N_11565,N_6062,N_6199);
nor U11566 (N_11566,N_7404,N_6898);
nor U11567 (N_11567,N_7902,N_7770);
and U11568 (N_11568,N_8251,N_8071);
nor U11569 (N_11569,N_8935,N_6645);
and U11570 (N_11570,N_7489,N_8092);
xor U11571 (N_11571,N_7051,N_8618);
nand U11572 (N_11572,N_7342,N_8105);
and U11573 (N_11573,N_8822,N_8541);
nand U11574 (N_11574,N_7818,N_7224);
nor U11575 (N_11575,N_7894,N_7241);
or U11576 (N_11576,N_8314,N_7403);
nand U11577 (N_11577,N_7446,N_6734);
or U11578 (N_11578,N_8718,N_6815);
nand U11579 (N_11579,N_8269,N_7328);
xor U11580 (N_11580,N_6494,N_7926);
or U11581 (N_11581,N_6003,N_6851);
nand U11582 (N_11582,N_7626,N_6481);
and U11583 (N_11583,N_7380,N_7363);
or U11584 (N_11584,N_7101,N_7296);
nand U11585 (N_11585,N_8912,N_6818);
nor U11586 (N_11586,N_7112,N_7098);
and U11587 (N_11587,N_7129,N_8314);
nand U11588 (N_11588,N_6383,N_8132);
or U11589 (N_11589,N_8328,N_6594);
or U11590 (N_11590,N_7245,N_8755);
nand U11591 (N_11591,N_6753,N_7187);
nand U11592 (N_11592,N_7327,N_6350);
or U11593 (N_11593,N_7204,N_7838);
and U11594 (N_11594,N_6694,N_6932);
xor U11595 (N_11595,N_7069,N_7686);
nor U11596 (N_11596,N_7591,N_8114);
and U11597 (N_11597,N_7774,N_8757);
nor U11598 (N_11598,N_7593,N_7495);
xnor U11599 (N_11599,N_6145,N_6250);
or U11600 (N_11600,N_7803,N_8991);
and U11601 (N_11601,N_6459,N_8198);
and U11602 (N_11602,N_8142,N_7058);
or U11603 (N_11603,N_7180,N_7593);
or U11604 (N_11604,N_8883,N_7110);
nor U11605 (N_11605,N_7315,N_7783);
xor U11606 (N_11606,N_6234,N_7172);
nand U11607 (N_11607,N_6357,N_6754);
or U11608 (N_11608,N_6533,N_7068);
nand U11609 (N_11609,N_6258,N_6254);
xor U11610 (N_11610,N_7520,N_6802);
nand U11611 (N_11611,N_6336,N_8772);
or U11612 (N_11612,N_8944,N_7738);
and U11613 (N_11613,N_6927,N_7304);
and U11614 (N_11614,N_8438,N_6817);
nand U11615 (N_11615,N_8046,N_8574);
nand U11616 (N_11616,N_6045,N_8018);
nor U11617 (N_11617,N_8372,N_7276);
or U11618 (N_11618,N_7768,N_7624);
or U11619 (N_11619,N_8870,N_6400);
nor U11620 (N_11620,N_7369,N_6045);
and U11621 (N_11621,N_8751,N_8486);
and U11622 (N_11622,N_6242,N_8283);
or U11623 (N_11623,N_6398,N_8305);
and U11624 (N_11624,N_7779,N_7486);
or U11625 (N_11625,N_6836,N_7828);
nor U11626 (N_11626,N_8978,N_7335);
or U11627 (N_11627,N_7046,N_6688);
or U11628 (N_11628,N_6744,N_7963);
or U11629 (N_11629,N_7094,N_8594);
or U11630 (N_11630,N_7171,N_8450);
or U11631 (N_11631,N_7611,N_8181);
nor U11632 (N_11632,N_8417,N_8586);
and U11633 (N_11633,N_7622,N_8332);
or U11634 (N_11634,N_8161,N_8971);
nor U11635 (N_11635,N_6129,N_8972);
nor U11636 (N_11636,N_7612,N_6869);
nor U11637 (N_11637,N_7667,N_7268);
or U11638 (N_11638,N_7251,N_7711);
nor U11639 (N_11639,N_6668,N_8298);
nand U11640 (N_11640,N_8562,N_8938);
nand U11641 (N_11641,N_6757,N_7163);
nand U11642 (N_11642,N_6541,N_7305);
nand U11643 (N_11643,N_7856,N_8871);
and U11644 (N_11644,N_7762,N_8847);
and U11645 (N_11645,N_6008,N_8301);
nor U11646 (N_11646,N_7206,N_7457);
nand U11647 (N_11647,N_7299,N_6500);
or U11648 (N_11648,N_6171,N_7370);
nand U11649 (N_11649,N_8150,N_8417);
nand U11650 (N_11650,N_6750,N_6089);
and U11651 (N_11651,N_8683,N_8423);
nand U11652 (N_11652,N_6755,N_8520);
nor U11653 (N_11653,N_7879,N_7786);
and U11654 (N_11654,N_6151,N_7692);
nand U11655 (N_11655,N_7431,N_8252);
nand U11656 (N_11656,N_6766,N_7414);
nand U11657 (N_11657,N_6153,N_7288);
nand U11658 (N_11658,N_7996,N_8556);
and U11659 (N_11659,N_8008,N_7278);
and U11660 (N_11660,N_7173,N_6621);
or U11661 (N_11661,N_6033,N_7327);
nor U11662 (N_11662,N_8363,N_6974);
nor U11663 (N_11663,N_8760,N_6225);
nand U11664 (N_11664,N_8929,N_7499);
and U11665 (N_11665,N_8453,N_6707);
xnor U11666 (N_11666,N_7835,N_7750);
or U11667 (N_11667,N_8000,N_7831);
or U11668 (N_11668,N_7267,N_7883);
or U11669 (N_11669,N_6118,N_7827);
xor U11670 (N_11670,N_7234,N_6098);
nand U11671 (N_11671,N_8363,N_6339);
or U11672 (N_11672,N_6080,N_7308);
nor U11673 (N_11673,N_6578,N_6314);
nor U11674 (N_11674,N_7901,N_8193);
xor U11675 (N_11675,N_6406,N_7451);
xnor U11676 (N_11676,N_7870,N_7546);
nand U11677 (N_11677,N_8311,N_7508);
nor U11678 (N_11678,N_6493,N_6809);
nor U11679 (N_11679,N_8135,N_8541);
and U11680 (N_11680,N_7599,N_7259);
nor U11681 (N_11681,N_6505,N_6043);
xnor U11682 (N_11682,N_6509,N_7406);
nand U11683 (N_11683,N_6650,N_6516);
and U11684 (N_11684,N_6046,N_7493);
xnor U11685 (N_11685,N_7881,N_7721);
nor U11686 (N_11686,N_6027,N_8080);
or U11687 (N_11687,N_7073,N_7638);
and U11688 (N_11688,N_6367,N_7461);
or U11689 (N_11689,N_7966,N_6168);
or U11690 (N_11690,N_6636,N_8229);
or U11691 (N_11691,N_6665,N_6074);
or U11692 (N_11692,N_7300,N_7746);
and U11693 (N_11693,N_8059,N_8738);
nand U11694 (N_11694,N_6654,N_7984);
and U11695 (N_11695,N_7081,N_8070);
xor U11696 (N_11696,N_7089,N_8089);
or U11697 (N_11697,N_7893,N_6868);
and U11698 (N_11698,N_7376,N_6269);
or U11699 (N_11699,N_6853,N_7318);
nand U11700 (N_11700,N_8878,N_6998);
xnor U11701 (N_11701,N_7167,N_6044);
and U11702 (N_11702,N_7723,N_8865);
nor U11703 (N_11703,N_6736,N_7321);
or U11704 (N_11704,N_6265,N_6289);
and U11705 (N_11705,N_6569,N_7503);
nor U11706 (N_11706,N_6561,N_6039);
nor U11707 (N_11707,N_8261,N_8768);
or U11708 (N_11708,N_7188,N_8006);
nor U11709 (N_11709,N_7206,N_6743);
and U11710 (N_11710,N_8662,N_6386);
nor U11711 (N_11711,N_6781,N_7712);
and U11712 (N_11712,N_7880,N_8523);
nor U11713 (N_11713,N_6109,N_8919);
nand U11714 (N_11714,N_6550,N_8164);
nand U11715 (N_11715,N_7536,N_8980);
nand U11716 (N_11716,N_7044,N_6800);
and U11717 (N_11717,N_7867,N_8248);
or U11718 (N_11718,N_6502,N_6591);
and U11719 (N_11719,N_6347,N_6596);
or U11720 (N_11720,N_6595,N_7013);
and U11721 (N_11721,N_7053,N_6060);
nor U11722 (N_11722,N_6765,N_6174);
nand U11723 (N_11723,N_7868,N_8127);
nor U11724 (N_11724,N_8661,N_6544);
or U11725 (N_11725,N_7174,N_8318);
nand U11726 (N_11726,N_8531,N_8888);
xnor U11727 (N_11727,N_6269,N_8757);
nand U11728 (N_11728,N_8107,N_6727);
or U11729 (N_11729,N_8481,N_8259);
or U11730 (N_11730,N_6982,N_6311);
nor U11731 (N_11731,N_6589,N_8490);
and U11732 (N_11732,N_7652,N_8912);
nand U11733 (N_11733,N_6539,N_7212);
or U11734 (N_11734,N_7385,N_8954);
nor U11735 (N_11735,N_6727,N_8185);
nor U11736 (N_11736,N_7925,N_6246);
xnor U11737 (N_11737,N_6530,N_6608);
or U11738 (N_11738,N_7395,N_8261);
nor U11739 (N_11739,N_7294,N_6210);
nor U11740 (N_11740,N_6415,N_8421);
and U11741 (N_11741,N_8226,N_6532);
and U11742 (N_11742,N_6615,N_7299);
xnor U11743 (N_11743,N_6103,N_8314);
nor U11744 (N_11744,N_8855,N_7454);
nand U11745 (N_11745,N_6267,N_8562);
or U11746 (N_11746,N_7449,N_8959);
nor U11747 (N_11747,N_8802,N_7747);
or U11748 (N_11748,N_6615,N_8576);
and U11749 (N_11749,N_7278,N_7858);
and U11750 (N_11750,N_7107,N_6254);
xor U11751 (N_11751,N_7315,N_8068);
or U11752 (N_11752,N_8732,N_6466);
xor U11753 (N_11753,N_7534,N_6541);
nor U11754 (N_11754,N_8810,N_8011);
nor U11755 (N_11755,N_8109,N_6988);
nand U11756 (N_11756,N_8680,N_6546);
or U11757 (N_11757,N_6650,N_7015);
or U11758 (N_11758,N_8778,N_7478);
nor U11759 (N_11759,N_8431,N_6682);
nand U11760 (N_11760,N_8810,N_6378);
xnor U11761 (N_11761,N_7106,N_6915);
and U11762 (N_11762,N_7758,N_7823);
nand U11763 (N_11763,N_7392,N_7634);
or U11764 (N_11764,N_6762,N_7559);
and U11765 (N_11765,N_6406,N_7650);
and U11766 (N_11766,N_6957,N_7836);
and U11767 (N_11767,N_6522,N_8482);
or U11768 (N_11768,N_7500,N_8551);
and U11769 (N_11769,N_6609,N_6920);
nor U11770 (N_11770,N_6900,N_6699);
xnor U11771 (N_11771,N_8772,N_7930);
xnor U11772 (N_11772,N_7015,N_6566);
or U11773 (N_11773,N_6590,N_6525);
nand U11774 (N_11774,N_8050,N_7041);
nor U11775 (N_11775,N_8806,N_6623);
nor U11776 (N_11776,N_7373,N_8464);
nor U11777 (N_11777,N_6833,N_8743);
and U11778 (N_11778,N_8398,N_7431);
or U11779 (N_11779,N_7227,N_6219);
and U11780 (N_11780,N_8182,N_6489);
and U11781 (N_11781,N_7038,N_7567);
nor U11782 (N_11782,N_8370,N_6449);
nor U11783 (N_11783,N_8377,N_6637);
nor U11784 (N_11784,N_6563,N_8461);
nor U11785 (N_11785,N_7007,N_7735);
nand U11786 (N_11786,N_8621,N_7119);
or U11787 (N_11787,N_7992,N_7145);
xnor U11788 (N_11788,N_8667,N_8849);
nor U11789 (N_11789,N_7158,N_6062);
or U11790 (N_11790,N_7408,N_7444);
nand U11791 (N_11791,N_8375,N_6438);
and U11792 (N_11792,N_6129,N_7435);
or U11793 (N_11793,N_8517,N_6270);
nand U11794 (N_11794,N_8549,N_7136);
nand U11795 (N_11795,N_6994,N_8864);
or U11796 (N_11796,N_6667,N_7830);
or U11797 (N_11797,N_8707,N_7493);
and U11798 (N_11798,N_7351,N_7852);
nand U11799 (N_11799,N_7140,N_7275);
nand U11800 (N_11800,N_6276,N_8927);
or U11801 (N_11801,N_7740,N_8945);
nand U11802 (N_11802,N_7425,N_6955);
or U11803 (N_11803,N_7611,N_6643);
or U11804 (N_11804,N_6264,N_6317);
nand U11805 (N_11805,N_8056,N_7868);
or U11806 (N_11806,N_7527,N_8893);
and U11807 (N_11807,N_7163,N_6992);
nor U11808 (N_11808,N_8735,N_8552);
nor U11809 (N_11809,N_6230,N_8217);
nor U11810 (N_11810,N_8936,N_8998);
and U11811 (N_11811,N_6356,N_6726);
nor U11812 (N_11812,N_8278,N_8668);
or U11813 (N_11813,N_7829,N_7549);
nor U11814 (N_11814,N_6491,N_7389);
and U11815 (N_11815,N_7894,N_6362);
nor U11816 (N_11816,N_8851,N_8990);
or U11817 (N_11817,N_6886,N_7134);
or U11818 (N_11818,N_6264,N_7465);
nand U11819 (N_11819,N_6453,N_8588);
or U11820 (N_11820,N_7804,N_6975);
nor U11821 (N_11821,N_6713,N_8805);
xnor U11822 (N_11822,N_8634,N_6868);
nor U11823 (N_11823,N_7561,N_8487);
nand U11824 (N_11824,N_6485,N_7869);
and U11825 (N_11825,N_6407,N_6095);
and U11826 (N_11826,N_7292,N_6412);
xor U11827 (N_11827,N_8976,N_8404);
and U11828 (N_11828,N_6069,N_6598);
nor U11829 (N_11829,N_8501,N_6477);
nor U11830 (N_11830,N_7688,N_7219);
and U11831 (N_11831,N_7812,N_6037);
nor U11832 (N_11832,N_6033,N_8163);
nand U11833 (N_11833,N_7249,N_6092);
or U11834 (N_11834,N_7239,N_7250);
nor U11835 (N_11835,N_8098,N_8273);
and U11836 (N_11836,N_6736,N_6129);
xor U11837 (N_11837,N_7937,N_6070);
nor U11838 (N_11838,N_7976,N_7970);
nor U11839 (N_11839,N_6870,N_7839);
nand U11840 (N_11840,N_7333,N_8930);
nand U11841 (N_11841,N_7248,N_8784);
or U11842 (N_11842,N_6857,N_6032);
or U11843 (N_11843,N_6649,N_7558);
nor U11844 (N_11844,N_6217,N_7941);
and U11845 (N_11845,N_7250,N_7578);
or U11846 (N_11846,N_7216,N_7221);
or U11847 (N_11847,N_6326,N_7542);
nor U11848 (N_11848,N_7374,N_6292);
or U11849 (N_11849,N_6145,N_6769);
and U11850 (N_11850,N_6074,N_6802);
nor U11851 (N_11851,N_8131,N_7248);
nor U11852 (N_11852,N_8515,N_8900);
and U11853 (N_11853,N_7903,N_7128);
or U11854 (N_11854,N_8424,N_8977);
and U11855 (N_11855,N_7438,N_6392);
or U11856 (N_11856,N_6006,N_6564);
or U11857 (N_11857,N_8530,N_7223);
and U11858 (N_11858,N_8250,N_8324);
and U11859 (N_11859,N_8193,N_8087);
nand U11860 (N_11860,N_6500,N_7820);
nor U11861 (N_11861,N_8387,N_8606);
nor U11862 (N_11862,N_6024,N_7152);
and U11863 (N_11863,N_6595,N_6997);
nor U11864 (N_11864,N_7144,N_6500);
xnor U11865 (N_11865,N_8189,N_7652);
nor U11866 (N_11866,N_8240,N_6926);
nor U11867 (N_11867,N_6747,N_8761);
nor U11868 (N_11868,N_6285,N_7203);
nor U11869 (N_11869,N_8717,N_6997);
nor U11870 (N_11870,N_7330,N_8668);
nor U11871 (N_11871,N_7886,N_6794);
or U11872 (N_11872,N_8103,N_6973);
xnor U11873 (N_11873,N_8671,N_6657);
and U11874 (N_11874,N_8930,N_8676);
or U11875 (N_11875,N_7555,N_8656);
or U11876 (N_11876,N_8190,N_8407);
or U11877 (N_11877,N_8339,N_7485);
nand U11878 (N_11878,N_7859,N_8838);
xor U11879 (N_11879,N_7079,N_8522);
nand U11880 (N_11880,N_6340,N_8983);
nor U11881 (N_11881,N_6368,N_7980);
or U11882 (N_11882,N_6214,N_6414);
nand U11883 (N_11883,N_6780,N_8348);
nor U11884 (N_11884,N_7238,N_7241);
and U11885 (N_11885,N_8315,N_6995);
and U11886 (N_11886,N_8907,N_8245);
nor U11887 (N_11887,N_7010,N_7097);
or U11888 (N_11888,N_7919,N_8044);
nor U11889 (N_11889,N_7224,N_6968);
xnor U11890 (N_11890,N_8714,N_6426);
and U11891 (N_11891,N_7131,N_8724);
and U11892 (N_11892,N_8353,N_6914);
or U11893 (N_11893,N_8114,N_8150);
xor U11894 (N_11894,N_7088,N_7504);
and U11895 (N_11895,N_6100,N_7312);
or U11896 (N_11896,N_7082,N_6547);
and U11897 (N_11897,N_8890,N_8999);
or U11898 (N_11898,N_7472,N_7235);
nor U11899 (N_11899,N_8939,N_7928);
and U11900 (N_11900,N_7222,N_6723);
nand U11901 (N_11901,N_8709,N_8145);
or U11902 (N_11902,N_8751,N_8092);
nand U11903 (N_11903,N_6961,N_8636);
xnor U11904 (N_11904,N_7440,N_6049);
or U11905 (N_11905,N_7274,N_6296);
xor U11906 (N_11906,N_6664,N_8113);
or U11907 (N_11907,N_8353,N_8314);
or U11908 (N_11908,N_7993,N_8581);
and U11909 (N_11909,N_7983,N_7932);
or U11910 (N_11910,N_8405,N_8927);
nor U11911 (N_11911,N_8220,N_6743);
nand U11912 (N_11912,N_8066,N_6855);
nand U11913 (N_11913,N_7954,N_8902);
xor U11914 (N_11914,N_7957,N_7703);
and U11915 (N_11915,N_8741,N_7098);
nand U11916 (N_11916,N_6132,N_7640);
nand U11917 (N_11917,N_7188,N_6499);
xnor U11918 (N_11918,N_7254,N_6057);
and U11919 (N_11919,N_8353,N_7942);
nor U11920 (N_11920,N_7869,N_7476);
or U11921 (N_11921,N_7476,N_6665);
nor U11922 (N_11922,N_6709,N_6145);
and U11923 (N_11923,N_7339,N_6715);
nor U11924 (N_11924,N_6850,N_8594);
and U11925 (N_11925,N_8653,N_7285);
or U11926 (N_11926,N_8489,N_6252);
and U11927 (N_11927,N_7462,N_6367);
nand U11928 (N_11928,N_7841,N_6967);
nor U11929 (N_11929,N_6536,N_8375);
and U11930 (N_11930,N_7657,N_6987);
xor U11931 (N_11931,N_8060,N_8646);
nand U11932 (N_11932,N_7352,N_6912);
nand U11933 (N_11933,N_6148,N_6247);
nand U11934 (N_11934,N_8214,N_7790);
and U11935 (N_11935,N_7321,N_6190);
or U11936 (N_11936,N_7719,N_8633);
and U11937 (N_11937,N_6746,N_7685);
nand U11938 (N_11938,N_7399,N_6325);
or U11939 (N_11939,N_7105,N_8031);
nand U11940 (N_11940,N_8893,N_8723);
xnor U11941 (N_11941,N_8206,N_7137);
xnor U11942 (N_11942,N_8412,N_6098);
nand U11943 (N_11943,N_6940,N_7578);
or U11944 (N_11944,N_8846,N_7952);
nand U11945 (N_11945,N_8197,N_6573);
nand U11946 (N_11946,N_8320,N_8704);
nor U11947 (N_11947,N_7103,N_8130);
nor U11948 (N_11948,N_7479,N_8527);
or U11949 (N_11949,N_6691,N_7814);
nand U11950 (N_11950,N_6516,N_8383);
or U11951 (N_11951,N_7653,N_7689);
nor U11952 (N_11952,N_7774,N_8181);
nand U11953 (N_11953,N_8665,N_7931);
or U11954 (N_11954,N_7632,N_7739);
and U11955 (N_11955,N_7698,N_7729);
xor U11956 (N_11956,N_6893,N_6066);
xnor U11957 (N_11957,N_7547,N_6045);
nor U11958 (N_11958,N_7434,N_8143);
and U11959 (N_11959,N_8756,N_6795);
nand U11960 (N_11960,N_8495,N_7271);
nand U11961 (N_11961,N_7896,N_8267);
and U11962 (N_11962,N_6220,N_8418);
or U11963 (N_11963,N_8805,N_8480);
and U11964 (N_11964,N_8122,N_6866);
nor U11965 (N_11965,N_7671,N_8318);
and U11966 (N_11966,N_8403,N_6450);
xor U11967 (N_11967,N_8648,N_8952);
nand U11968 (N_11968,N_8503,N_8924);
nand U11969 (N_11969,N_6947,N_8157);
nand U11970 (N_11970,N_7958,N_6234);
and U11971 (N_11971,N_6661,N_8492);
nor U11972 (N_11972,N_8473,N_8743);
and U11973 (N_11973,N_8374,N_6031);
nand U11974 (N_11974,N_6430,N_7741);
and U11975 (N_11975,N_6820,N_6683);
or U11976 (N_11976,N_6922,N_8597);
nand U11977 (N_11977,N_6887,N_7072);
or U11978 (N_11978,N_6905,N_7895);
nor U11979 (N_11979,N_8047,N_8748);
nor U11980 (N_11980,N_6919,N_7956);
or U11981 (N_11981,N_7144,N_7984);
nand U11982 (N_11982,N_7886,N_7404);
nor U11983 (N_11983,N_6321,N_6540);
xor U11984 (N_11984,N_6329,N_8547);
and U11985 (N_11985,N_7338,N_8527);
or U11986 (N_11986,N_6358,N_7375);
nand U11987 (N_11987,N_7932,N_6503);
nor U11988 (N_11988,N_7235,N_7488);
or U11989 (N_11989,N_6825,N_8026);
and U11990 (N_11990,N_7511,N_7353);
or U11991 (N_11991,N_7384,N_7275);
and U11992 (N_11992,N_8020,N_7508);
nor U11993 (N_11993,N_6082,N_8812);
nor U11994 (N_11994,N_6017,N_7484);
xor U11995 (N_11995,N_7189,N_7686);
or U11996 (N_11996,N_7660,N_6746);
and U11997 (N_11997,N_7725,N_7700);
or U11998 (N_11998,N_7513,N_7873);
nor U11999 (N_11999,N_7842,N_6088);
nor U12000 (N_12000,N_11448,N_10307);
nor U12001 (N_12001,N_11482,N_9212);
or U12002 (N_12002,N_11905,N_10077);
or U12003 (N_12003,N_9761,N_9178);
nor U12004 (N_12004,N_10853,N_9953);
nand U12005 (N_12005,N_11276,N_11500);
or U12006 (N_12006,N_9543,N_11970);
and U12007 (N_12007,N_11785,N_9088);
nand U12008 (N_12008,N_11220,N_11731);
and U12009 (N_12009,N_11441,N_11579);
nor U12010 (N_12010,N_11615,N_11527);
or U12011 (N_12011,N_11042,N_10009);
nor U12012 (N_12012,N_10066,N_11906);
nand U12013 (N_12013,N_10492,N_11384);
and U12014 (N_12014,N_11090,N_10396);
nor U12015 (N_12015,N_10131,N_11987);
nand U12016 (N_12016,N_10632,N_9840);
nor U12017 (N_12017,N_9157,N_9272);
nor U12018 (N_12018,N_10942,N_9738);
and U12019 (N_12019,N_9964,N_11577);
or U12020 (N_12020,N_10812,N_10173);
nor U12021 (N_12021,N_11281,N_10777);
or U12022 (N_12022,N_9805,N_11036);
and U12023 (N_12023,N_10969,N_11822);
and U12024 (N_12024,N_9483,N_11857);
nand U12025 (N_12025,N_9059,N_11889);
nand U12026 (N_12026,N_10222,N_10638);
and U12027 (N_12027,N_11188,N_11844);
nand U12028 (N_12028,N_10020,N_9806);
nor U12029 (N_12029,N_10138,N_11138);
and U12030 (N_12030,N_11287,N_10398);
or U12031 (N_12031,N_9347,N_10167);
or U12032 (N_12032,N_11122,N_10677);
xnor U12033 (N_12033,N_11403,N_9714);
or U12034 (N_12034,N_10185,N_11823);
nand U12035 (N_12035,N_9165,N_10986);
nand U12036 (N_12036,N_10019,N_9139);
nor U12037 (N_12037,N_11072,N_9441);
or U12038 (N_12038,N_10027,N_10482);
or U12039 (N_12039,N_10051,N_9175);
nor U12040 (N_12040,N_9872,N_11911);
nand U12041 (N_12041,N_10663,N_10116);
or U12042 (N_12042,N_10792,N_11428);
or U12043 (N_12043,N_9900,N_9439);
xor U12044 (N_12044,N_10617,N_11427);
nor U12045 (N_12045,N_11267,N_11759);
nor U12046 (N_12046,N_10878,N_9916);
nor U12047 (N_12047,N_9952,N_11768);
or U12048 (N_12048,N_10060,N_10514);
or U12049 (N_12049,N_9885,N_9002);
nand U12050 (N_12050,N_11440,N_11841);
or U12051 (N_12051,N_11039,N_10428);
and U12052 (N_12052,N_11582,N_10523);
nor U12053 (N_12053,N_11076,N_9834);
or U12054 (N_12054,N_9592,N_9531);
and U12055 (N_12055,N_10321,N_9263);
nand U12056 (N_12056,N_10725,N_10723);
nor U12057 (N_12057,N_10856,N_11132);
or U12058 (N_12058,N_11912,N_11873);
or U12059 (N_12059,N_10050,N_10274);
and U12060 (N_12060,N_9809,N_10443);
nand U12061 (N_12061,N_9475,N_10956);
nor U12062 (N_12062,N_11474,N_10933);
and U12063 (N_12063,N_10798,N_10434);
and U12064 (N_12064,N_11801,N_11203);
or U12065 (N_12065,N_10404,N_11169);
or U12066 (N_12066,N_9598,N_9903);
nand U12067 (N_12067,N_10742,N_10685);
nand U12068 (N_12068,N_10953,N_11364);
nand U12069 (N_12069,N_10362,N_9436);
xor U12070 (N_12070,N_11610,N_9889);
and U12071 (N_12071,N_9216,N_10955);
and U12072 (N_12072,N_9315,N_9676);
nand U12073 (N_12073,N_9381,N_9637);
nand U12074 (N_12074,N_11189,N_10268);
and U12075 (N_12075,N_9351,N_10254);
or U12076 (N_12076,N_9253,N_10401);
and U12077 (N_12077,N_9061,N_10213);
nand U12078 (N_12078,N_11985,N_11758);
nand U12079 (N_12079,N_9433,N_9181);
nor U12080 (N_12080,N_11517,N_9003);
nor U12081 (N_12081,N_9939,N_10640);
nor U12082 (N_12082,N_9249,N_10745);
nor U12083 (N_12083,N_10872,N_9070);
and U12084 (N_12084,N_11134,N_9756);
or U12085 (N_12085,N_10505,N_10360);
and U12086 (N_12086,N_9682,N_10882);
and U12087 (N_12087,N_10111,N_11174);
nand U12088 (N_12088,N_10822,N_11376);
and U12089 (N_12089,N_11549,N_9521);
or U12090 (N_12090,N_11454,N_9584);
nand U12091 (N_12091,N_11321,N_9461);
xnor U12092 (N_12092,N_10573,N_11054);
or U12093 (N_12093,N_9015,N_10394);
nand U12094 (N_12094,N_9678,N_10898);
nand U12095 (N_12095,N_11583,N_9367);
nand U12096 (N_12096,N_9813,N_10200);
nor U12097 (N_12097,N_10603,N_11730);
and U12098 (N_12098,N_11111,N_11994);
or U12099 (N_12099,N_11261,N_9286);
and U12100 (N_12100,N_9213,N_11125);
or U12101 (N_12101,N_9202,N_11308);
nor U12102 (N_12102,N_10769,N_10072);
and U12103 (N_12103,N_10546,N_10276);
nand U12104 (N_12104,N_10824,N_11946);
and U12105 (N_12105,N_11317,N_11824);
nand U12106 (N_12106,N_9874,N_9364);
nor U12107 (N_12107,N_9402,N_10080);
nand U12108 (N_12108,N_11605,N_10214);
nand U12109 (N_12109,N_11791,N_9743);
nand U12110 (N_12110,N_10493,N_9228);
and U12111 (N_12111,N_9773,N_9236);
nand U12112 (N_12112,N_11638,N_10304);
and U12113 (N_12113,N_9265,N_9371);
or U12114 (N_12114,N_11502,N_9824);
and U12115 (N_12115,N_9753,N_10188);
xor U12116 (N_12116,N_9944,N_10481);
nor U12117 (N_12117,N_9186,N_10251);
or U12118 (N_12118,N_9593,N_9241);
or U12119 (N_12119,N_9512,N_11473);
nor U12120 (N_12120,N_9276,N_10599);
or U12121 (N_12121,N_11266,N_9231);
nand U12122 (N_12122,N_10292,N_9163);
or U12123 (N_12123,N_11709,N_9452);
nand U12124 (N_12124,N_11435,N_11986);
nand U12125 (N_12125,N_10311,N_9618);
nor U12126 (N_12126,N_10296,N_10497);
or U12127 (N_12127,N_9414,N_10002);
nor U12128 (N_12128,N_11116,N_9579);
nor U12129 (N_12129,N_9481,N_10896);
or U12130 (N_12130,N_9324,N_11762);
nand U12131 (N_12131,N_9852,N_10923);
nand U12132 (N_12132,N_11957,N_11350);
nand U12133 (N_12133,N_10449,N_10595);
and U12134 (N_12134,N_11271,N_9026);
nor U12135 (N_12135,N_10682,N_11277);
or U12136 (N_12136,N_11247,N_9039);
or U12137 (N_12137,N_9879,N_10684);
or U12138 (N_12138,N_11333,N_10548);
and U12139 (N_12139,N_10840,N_11932);
or U12140 (N_12140,N_11504,N_9387);
nand U12141 (N_12141,N_11108,N_11655);
nand U12142 (N_12142,N_11621,N_9655);
and U12143 (N_12143,N_11982,N_11816);
nand U12144 (N_12144,N_9901,N_11499);
and U12145 (N_12145,N_11078,N_11388);
nor U12146 (N_12146,N_11493,N_11687);
and U12147 (N_12147,N_9049,N_11828);
and U12148 (N_12148,N_10089,N_11636);
and U12149 (N_12149,N_10110,N_10978);
or U12150 (N_12150,N_11130,N_9455);
and U12151 (N_12151,N_10155,N_11180);
xor U12152 (N_12152,N_11217,N_11066);
or U12153 (N_12153,N_9140,N_10120);
nor U12154 (N_12154,N_9501,N_11850);
nand U12155 (N_12155,N_11306,N_10561);
xor U12156 (N_12156,N_10577,N_10176);
and U12157 (N_12157,N_11442,N_9426);
nor U12158 (N_12158,N_11962,N_11097);
nand U12159 (N_12159,N_10193,N_9014);
and U12160 (N_12160,N_10436,N_9240);
or U12161 (N_12161,N_10132,N_11774);
or U12162 (N_12162,N_9894,N_11914);
xnor U12163 (N_12163,N_10984,N_11784);
nand U12164 (N_12164,N_9559,N_10737);
nand U12165 (N_12165,N_10618,N_11264);
xnor U12166 (N_12166,N_11236,N_11398);
and U12167 (N_12167,N_9118,N_9029);
xnor U12168 (N_12168,N_10946,N_11954);
nand U12169 (N_12169,N_11127,N_11006);
and U12170 (N_12170,N_9326,N_10907);
or U12171 (N_12171,N_10863,N_11327);
and U12172 (N_12172,N_9938,N_10258);
or U12173 (N_12173,N_10588,N_11222);
nor U12174 (N_12174,N_9526,N_9179);
or U12175 (N_12175,N_11164,N_9660);
nor U12176 (N_12176,N_9319,N_10536);
or U12177 (N_12177,N_11597,N_11748);
xor U12178 (N_12178,N_10761,N_11926);
nor U12179 (N_12179,N_11811,N_11349);
xor U12180 (N_12180,N_10044,N_10951);
nand U12181 (N_12181,N_10526,N_9079);
and U12182 (N_12182,N_11852,N_10478);
and U12183 (N_12183,N_9052,N_11898);
nand U12184 (N_12184,N_11311,N_10147);
or U12185 (N_12185,N_11034,N_11556);
nor U12186 (N_12186,N_10438,N_11543);
xor U12187 (N_12187,N_9233,N_9060);
xnor U12188 (N_12188,N_10294,N_9605);
xor U12189 (N_12189,N_11901,N_11681);
nor U12190 (N_12190,N_11386,N_11790);
or U12191 (N_12191,N_11980,N_9835);
and U12192 (N_12192,N_11046,N_11197);
nand U12193 (N_12193,N_11481,N_10234);
nand U12194 (N_12194,N_10062,N_11148);
nor U12195 (N_12195,N_11848,N_11967);
nor U12196 (N_12196,N_9292,N_10619);
nor U12197 (N_12197,N_9106,N_10064);
xnor U12198 (N_12198,N_9707,N_9159);
nand U12199 (N_12199,N_11369,N_10578);
nor U12200 (N_12200,N_9502,N_10842);
nor U12201 (N_12201,N_9604,N_10847);
and U12202 (N_12202,N_9812,N_10952);
nand U12203 (N_12203,N_11686,N_11747);
nor U12204 (N_12204,N_9293,N_11918);
nand U12205 (N_12205,N_10017,N_9195);
and U12206 (N_12206,N_11018,N_11477);
nor U12207 (N_12207,N_11870,N_11834);
or U12208 (N_12208,N_11456,N_9842);
and U12209 (N_12209,N_9398,N_9784);
or U12210 (N_12210,N_9899,N_9205);
or U12211 (N_12211,N_11729,N_9078);
nor U12212 (N_12212,N_10779,N_11113);
nor U12213 (N_12213,N_9831,N_9736);
xor U12214 (N_12214,N_9416,N_11230);
or U12215 (N_12215,N_11678,N_9620);
nand U12216 (N_12216,N_9645,N_11783);
or U12217 (N_12217,N_11601,N_9480);
nor U12218 (N_12218,N_10437,N_10506);
nand U12219 (N_12219,N_9574,N_9582);
or U12220 (N_12220,N_9551,N_11891);
or U12221 (N_12221,N_10270,N_10718);
nor U12222 (N_12222,N_10248,N_11890);
nor U12223 (N_12223,N_11953,N_10145);
and U12224 (N_12224,N_9599,N_11329);
or U12225 (N_12225,N_10457,N_11325);
and U12226 (N_12226,N_9130,N_11566);
nand U12227 (N_12227,N_9010,N_9558);
xor U12228 (N_12228,N_9575,N_10369);
or U12229 (N_12229,N_11862,N_10832);
and U12230 (N_12230,N_10650,N_9578);
or U12231 (N_12231,N_9105,N_10750);
nor U12232 (N_12232,N_9415,N_9121);
or U12233 (N_12233,N_10287,N_10560);
xor U12234 (N_12234,N_9065,N_10701);
nand U12235 (N_12235,N_9362,N_10332);
nor U12236 (N_12236,N_10297,N_10339);
and U12237 (N_12237,N_10759,N_10889);
nor U12238 (N_12238,N_10717,N_11272);
or U12239 (N_12239,N_9602,N_9820);
or U12240 (N_12240,N_9494,N_11830);
and U12241 (N_12241,N_9383,N_10722);
nor U12242 (N_12242,N_10883,N_9765);
nor U12243 (N_12243,N_11209,N_11307);
or U12244 (N_12244,N_10117,N_10743);
and U12245 (N_12245,N_9344,N_11089);
nand U12246 (N_12246,N_9643,N_11143);
or U12247 (N_12247,N_11245,N_9606);
nand U12248 (N_12248,N_9142,N_9495);
nand U12249 (N_12249,N_11592,N_10865);
nor U12250 (N_12250,N_11546,N_10411);
and U12251 (N_12251,N_11486,N_9571);
xnor U12252 (N_12252,N_9177,N_9173);
and U12253 (N_12253,N_10586,N_9244);
nor U12254 (N_12254,N_11951,N_9400);
or U12255 (N_12255,N_9112,N_11219);
or U12256 (N_12256,N_11623,N_11728);
nand U12257 (N_12257,N_10754,N_10881);
nor U12258 (N_12258,N_11205,N_9093);
xor U12259 (N_12259,N_9023,N_9595);
nand U12260 (N_12260,N_10309,N_11609);
xnor U12261 (N_12261,N_10753,N_9208);
nand U12262 (N_12262,N_9927,N_10053);
nor U12263 (N_12263,N_11255,N_10991);
nor U12264 (N_12264,N_10756,N_11381);
nand U12265 (N_12265,N_10197,N_10610);
nor U12266 (N_12266,N_10460,N_11160);
nor U12267 (N_12267,N_10129,N_11304);
and U12268 (N_12268,N_9149,N_10585);
nand U12269 (N_12269,N_11375,N_10263);
nor U12270 (N_12270,N_9500,N_9227);
nand U12271 (N_12271,N_9154,N_10508);
nor U12272 (N_12272,N_11224,N_10075);
and U12273 (N_12273,N_11140,N_10144);
nand U12274 (N_12274,N_10710,N_11706);
or U12275 (N_12275,N_10305,N_9697);
nand U12276 (N_12276,N_10078,N_10741);
nor U12277 (N_12277,N_11101,N_11518);
or U12278 (N_12278,N_11256,N_11528);
nor U12279 (N_12279,N_9392,N_11952);
and U12280 (N_12280,N_9300,N_9905);
and U12281 (N_12281,N_9096,N_9138);
and U12282 (N_12282,N_9745,N_10999);
nor U12283 (N_12283,N_10563,N_9336);
nor U12284 (N_12284,N_9919,N_10327);
nor U12285 (N_12285,N_10272,N_10574);
nor U12286 (N_12286,N_10797,N_11789);
nor U12287 (N_12287,N_9379,N_10049);
nand U12288 (N_12288,N_10819,N_9285);
and U12289 (N_12289,N_9020,N_11231);
and U12290 (N_12290,N_11600,N_9148);
or U12291 (N_12291,N_11563,N_10232);
nor U12292 (N_12292,N_9691,N_11001);
nand U12293 (N_12293,N_10996,N_9548);
or U12294 (N_12294,N_10974,N_11507);
and U12295 (N_12295,N_9825,N_9295);
and U12296 (N_12296,N_9162,N_9127);
and U12297 (N_12297,N_10781,N_10802);
or U12298 (N_12298,N_10105,N_11447);
xnor U12299 (N_12299,N_11562,N_10476);
nor U12300 (N_12300,N_11254,N_9073);
nor U12301 (N_12301,N_9283,N_10054);
xnor U12302 (N_12302,N_11930,N_9926);
xor U12303 (N_12303,N_9522,N_9378);
nor U12304 (N_12304,N_10553,N_11040);
nor U12305 (N_12305,N_11379,N_10712);
or U12306 (N_12306,N_9679,N_10024);
nand U12307 (N_12307,N_9920,N_9430);
nand U12308 (N_12308,N_11648,N_9935);
or U12309 (N_12309,N_10337,N_9038);
nor U12310 (N_12310,N_9853,N_9696);
or U12311 (N_12311,N_10336,N_11494);
or U12312 (N_12312,N_11360,N_11988);
and U12313 (N_12313,N_10765,N_10874);
nor U12314 (N_12314,N_11478,N_11679);
nor U12315 (N_12315,N_9477,N_9719);
and U12316 (N_12316,N_9349,N_9051);
xnor U12317 (N_12317,N_11925,N_11192);
and U12318 (N_12318,N_10930,N_11511);
and U12319 (N_12319,N_10830,N_10491);
and U12320 (N_12320,N_11243,N_10661);
or U12321 (N_12321,N_11720,N_10273);
nand U12322 (N_12322,N_9811,N_11893);
and U12323 (N_12323,N_10215,N_9866);
nand U12324 (N_12324,N_10036,N_9573);
nor U12325 (N_12325,N_9766,N_9983);
or U12326 (N_12326,N_9591,N_11022);
or U12327 (N_12327,N_10099,N_11956);
nand U12328 (N_12328,N_9911,N_11115);
and U12329 (N_12329,N_11885,N_9530);
nor U12330 (N_12330,N_11743,N_10844);
nor U12331 (N_12331,N_10003,N_9126);
nand U12332 (N_12332,N_10525,N_10180);
xnor U12333 (N_12333,N_11644,N_10736);
nand U12334 (N_12334,N_9200,N_10624);
nand U12335 (N_12335,N_9675,N_10043);
and U12336 (N_12336,N_10121,N_9373);
nand U12337 (N_12337,N_11475,N_10347);
or U12338 (N_12338,N_9160,N_9056);
and U12339 (N_12339,N_11087,N_9497);
nor U12340 (N_12340,N_11662,N_10995);
nor U12341 (N_12341,N_9391,N_11766);
or U12342 (N_12342,N_9504,N_10607);
nand U12343 (N_12343,N_9459,N_11061);
or U12344 (N_12344,N_10890,N_10390);
nor U12345 (N_12345,N_10079,N_11241);
or U12346 (N_12346,N_11080,N_10137);
and U12347 (N_12347,N_10417,N_10266);
or U12348 (N_12348,N_9837,N_9053);
and U12349 (N_12349,N_9103,N_9796);
nand U12350 (N_12350,N_9062,N_9961);
xor U12351 (N_12351,N_11351,N_9668);
nand U12352 (N_12352,N_9978,N_10450);
nand U12353 (N_12353,N_10261,N_11515);
and U12354 (N_12354,N_11630,N_10562);
nand U12355 (N_12355,N_9528,N_11634);
nand U12356 (N_12356,N_11365,N_11249);
and U12357 (N_12357,N_10922,N_10947);
and U12358 (N_12358,N_11257,N_9438);
nand U12359 (N_12359,N_11826,N_11539);
nor U12360 (N_12360,N_11691,N_9485);
nor U12361 (N_12361,N_9529,N_11663);
or U12362 (N_12362,N_9050,N_11059);
and U12363 (N_12363,N_10739,N_10480);
nor U12364 (N_12364,N_11095,N_9445);
nor U12365 (N_12365,N_10864,N_9778);
nand U12366 (N_12366,N_10299,N_9124);
nor U12367 (N_12367,N_9956,N_9854);
and U12368 (N_12368,N_10157,N_10979);
nor U12369 (N_12369,N_11452,N_11645);
and U12370 (N_12370,N_9058,N_11124);
or U12371 (N_12371,N_10389,N_10683);
or U12372 (N_12372,N_11689,N_11451);
or U12373 (N_12373,N_10782,N_11651);
and U12374 (N_12374,N_10503,N_9995);
nor U12375 (N_12375,N_10047,N_11856);
and U12376 (N_12376,N_9246,N_9337);
nor U12377 (N_12377,N_11204,N_11781);
or U12378 (N_12378,N_11410,N_10662);
or U12379 (N_12379,N_9449,N_10366);
nor U12380 (N_12380,N_10937,N_10286);
nor U12381 (N_12381,N_10186,N_10870);
nand U12382 (N_12382,N_9016,N_11736);
and U12383 (N_12383,N_10228,N_9792);
and U12384 (N_12384,N_9284,N_11541);
and U12385 (N_12385,N_11752,N_11433);
or U12386 (N_12386,N_10895,N_9589);
nor U12387 (N_12387,N_10811,N_9942);
nand U12388 (N_12388,N_10988,N_9429);
and U12389 (N_12389,N_10735,N_10423);
and U12390 (N_12390,N_10410,N_10418);
nor U12391 (N_12391,N_10342,N_9612);
nand U12392 (N_12392,N_11996,N_9258);
and U12393 (N_12393,N_11860,N_10647);
or U12394 (N_12394,N_11868,N_10634);
nand U12395 (N_12395,N_9590,N_10928);
or U12396 (N_12396,N_11426,N_11966);
nor U12397 (N_12397,N_10859,N_9537);
and U12398 (N_12398,N_11286,N_9462);
and U12399 (N_12399,N_10380,N_10317);
and U12400 (N_12400,N_11575,N_9252);
nor U12401 (N_12401,N_9305,N_10744);
or U12402 (N_12402,N_9182,N_11593);
xnor U12403 (N_12403,N_11314,N_11104);
nor U12404 (N_12404,N_11538,N_10190);
nor U12405 (N_12405,N_11401,N_10789);
or U12406 (N_12406,N_10444,N_10925);
nand U12407 (N_12407,N_11552,N_11782);
and U12408 (N_12408,N_11027,N_9151);
xnor U12409 (N_12409,N_9856,N_9539);
or U12410 (N_12410,N_11278,N_10720);
nor U12411 (N_12411,N_9777,N_9486);
or U12412 (N_12412,N_10852,N_10912);
nand U12413 (N_12413,N_11847,N_10554);
nor U12414 (N_12414,N_10333,N_9012);
nor U12415 (N_12415,N_11806,N_11118);
nor U12416 (N_12416,N_9467,N_11855);
nand U12417 (N_12417,N_10775,N_11015);
nor U12418 (N_12418,N_11414,N_11128);
and U12419 (N_12419,N_9851,N_11156);
nor U12420 (N_12420,N_9787,N_11722);
and U12421 (N_12421,N_10076,N_9962);
and U12422 (N_12422,N_9623,N_11081);
and U12423 (N_12423,N_11010,N_11126);
and U12424 (N_12424,N_10689,N_11050);
nand U12425 (N_12425,N_9304,N_9794);
nand U12426 (N_12426,N_9490,N_9380);
and U12427 (N_12427,N_10537,N_11310);
and U12428 (N_12428,N_11313,N_11359);
nor U12429 (N_12429,N_9167,N_10026);
nor U12430 (N_12430,N_11484,N_10081);
or U12431 (N_12431,N_11107,N_9239);
xnor U12432 (N_12432,N_9546,N_11771);
nand U12433 (N_12433,N_11353,N_10746);
xor U12434 (N_12434,N_9072,N_10748);
and U12435 (N_12435,N_10166,N_9210);
nand U12436 (N_12436,N_10971,N_10245);
and U12437 (N_12437,N_9683,N_9915);
nand U12438 (N_12438,N_9224,N_10733);
and U12439 (N_12439,N_11469,N_9703);
and U12440 (N_12440,N_10393,N_9384);
xnor U12441 (N_12441,N_10122,N_11740);
and U12442 (N_12442,N_9921,N_9338);
nor U12443 (N_12443,N_10729,N_11657);
xor U12444 (N_12444,N_10218,N_10343);
or U12445 (N_12445,N_10106,N_10581);
nand U12446 (N_12446,N_10221,N_9715);
nand U12447 (N_12447,N_11028,N_11936);
and U12448 (N_12448,N_11288,N_9608);
nand U12449 (N_12449,N_11643,N_10379);
nand U12450 (N_12450,N_11355,N_9909);
nand U12451 (N_12451,N_10539,N_9999);
or U12452 (N_12452,N_9568,N_10855);
nand U12453 (N_12453,N_9453,N_9071);
or U12454 (N_12454,N_11041,N_11235);
or U12455 (N_12455,N_9564,N_11817);
or U12456 (N_12456,N_10447,N_9583);
nor U12457 (N_12457,N_11029,N_9829);
or U12458 (N_12458,N_10242,N_11279);
or U12459 (N_12459,N_10641,N_11165);
or U12460 (N_12460,N_9622,N_10945);
nor U12461 (N_12461,N_10916,N_9170);
nand U12462 (N_12462,N_10814,N_10244);
nor U12463 (N_12463,N_9363,N_9994);
nand U12464 (N_12464,N_10635,N_11646);
or U12465 (N_12465,N_10948,N_10894);
nor U12466 (N_12466,N_9299,N_10397);
xor U12467 (N_12467,N_10648,N_11417);
xnor U12468 (N_12468,N_10101,N_10156);
or U12469 (N_12469,N_9279,N_9783);
xnor U12470 (N_12470,N_11305,N_9199);
or U12471 (N_12471,N_9960,N_11032);
nand U12472 (N_12472,N_9638,N_11733);
and U12473 (N_12473,N_10601,N_9185);
and U12474 (N_12474,N_9041,N_9720);
nor U12475 (N_12475,N_10582,N_10614);
nor U12476 (N_12476,N_11596,N_10202);
nand U12477 (N_12477,N_11769,N_10283);
nand U12478 (N_12478,N_9247,N_9774);
nand U12479 (N_12479,N_9022,N_11900);
and U12480 (N_12480,N_10096,N_9097);
nand U12481 (N_12481,N_11700,N_9189);
or U12482 (N_12482,N_11263,N_9048);
nand U12483 (N_12483,N_11086,N_9764);
or U12484 (N_12484,N_9844,N_10289);
and U12485 (N_12485,N_10055,N_11488);
and U12486 (N_12486,N_11434,N_11883);
nor U12487 (N_12487,N_9870,N_9552);
or U12488 (N_12488,N_11569,N_10758);
xor U12489 (N_12489,N_10615,N_10686);
nor U12490 (N_12490,N_11688,N_11135);
and U12491 (N_12491,N_10331,N_9063);
nand U12492 (N_12492,N_11470,N_9465);
and U12493 (N_12493,N_10467,N_11234);
nand U12494 (N_12494,N_11377,N_11370);
or U12495 (N_12495,N_10322,N_9094);
nor U12496 (N_12496,N_11069,N_11529);
nor U12497 (N_12497,N_9759,N_11888);
nor U12498 (N_12498,N_10584,N_10238);
nand U12499 (N_12499,N_10994,N_9751);
nand U12500 (N_12500,N_11757,N_11411);
nor U12501 (N_12501,N_10230,N_9800);
nor U12502 (N_12502,N_10773,N_10616);
xnor U12503 (N_12503,N_9187,N_9587);
nor U12504 (N_12504,N_9068,N_9913);
and U12505 (N_12505,N_10407,N_11338);
nand U12506 (N_12506,N_10869,N_11929);
and U12507 (N_12507,N_9116,N_10306);
nand U12508 (N_12508,N_11829,N_11959);
nor U12509 (N_12509,N_11382,N_10082);
nor U12510 (N_12510,N_10767,N_11777);
or U12511 (N_12511,N_10123,N_9632);
xnor U12512 (N_12512,N_10669,N_9451);
nor U12513 (N_12513,N_9630,N_11404);
xor U12514 (N_12514,N_10471,N_10198);
or U12515 (N_12515,N_11843,N_9356);
nor U12516 (N_12516,N_9168,N_9488);
or U12517 (N_12517,N_10083,N_11301);
nand U12518 (N_12518,N_10402,N_11437);
and U12519 (N_12519,N_9701,N_10152);
xor U12520 (N_12520,N_11735,N_10113);
or U12521 (N_12521,N_10866,N_10124);
or U12522 (N_12522,N_11978,N_11323);
and U12523 (N_12523,N_9193,N_11550);
and U12524 (N_12524,N_9621,N_11030);
nor U12525 (N_12525,N_10657,N_10579);
and U12526 (N_12526,N_11400,N_10087);
or U12527 (N_12527,N_11136,N_9456);
nand U12528 (N_12528,N_10602,N_11618);
and U12529 (N_12529,N_10237,N_11865);
nand U12530 (N_12530,N_11331,N_10357);
xnor U12531 (N_12531,N_10241,N_11664);
xor U12532 (N_12532,N_11702,N_9875);
and U12533 (N_12533,N_11472,N_9498);
nand U12534 (N_12534,N_9998,N_11340);
xor U12535 (N_12535,N_9183,N_9515);
nand U12536 (N_12536,N_10039,N_10495);
xor U12537 (N_12537,N_10732,N_10243);
nor U12538 (N_12538,N_10353,N_11803);
nand U12539 (N_12539,N_9664,N_11580);
or U12540 (N_12540,N_9607,N_10382);
and U12541 (N_12541,N_9700,N_9728);
or U12542 (N_12542,N_11439,N_10637);
nand U12543 (N_12543,N_9479,N_10281);
and U12544 (N_12544,N_11613,N_10494);
and U12545 (N_12545,N_10665,N_10259);
or U12546 (N_12546,N_10567,N_11269);
nor U12547 (N_12547,N_11058,N_10126);
and U12548 (N_12548,N_9633,N_10821);
nor U12549 (N_12549,N_9358,N_11821);
xor U12550 (N_12550,N_10544,N_11068);
and U12551 (N_12551,N_9350,N_10045);
and U12552 (N_12552,N_10141,N_9095);
and U12553 (N_12553,N_10968,N_11225);
and U12554 (N_12554,N_10207,N_9506);
nor U12555 (N_12555,N_10088,N_11751);
nor U12556 (N_12556,N_9718,N_11878);
nor U12557 (N_12557,N_11732,N_11356);
or U12558 (N_12558,N_11449,N_10597);
nor U12559 (N_12559,N_11055,N_9000);
and U12560 (N_12560,N_9006,N_9217);
nor U12561 (N_12561,N_10693,N_10386);
or U12562 (N_12562,N_9656,N_11693);
nand U12563 (N_12563,N_9146,N_10919);
and U12564 (N_12564,N_9113,N_11248);
nor U12565 (N_12565,N_10372,N_11955);
xor U12566 (N_12566,N_11144,N_11285);
nand U12567 (N_12567,N_11316,N_9925);
or U12568 (N_12568,N_9847,N_9685);
nor U12569 (N_12569,N_11933,N_9102);
xnor U12570 (N_12570,N_9080,N_11492);
and U12571 (N_12571,N_10810,N_10031);
or U12572 (N_12572,N_9802,N_9731);
nor U12573 (N_12573,N_10879,N_9503);
and U12574 (N_12574,N_11468,N_9520);
or U12575 (N_12575,N_10489,N_11024);
xnor U12576 (N_12576,N_9828,N_10345);
nor U12577 (N_12577,N_11207,N_9366);
nor U12578 (N_12578,N_9448,N_9544);
nand U12579 (N_12579,N_11780,N_11520);
or U12580 (N_12580,N_11182,N_10593);
nor U12581 (N_12581,N_10959,N_10531);
nand U12582 (N_12582,N_11616,N_10596);
or U12583 (N_12583,N_9666,N_9799);
nand U12584 (N_12584,N_10470,N_11176);
xnor U12585 (N_12585,N_10097,N_9108);
or U12586 (N_12586,N_10931,N_11282);
or U12587 (N_12587,N_11837,N_11070);
xor U12588 (N_12588,N_11226,N_9721);
and U12589 (N_12589,N_11578,N_10171);
nor U12590 (N_12590,N_11354,N_11166);
xor U12591 (N_12591,N_10358,N_11739);
or U12592 (N_12592,N_11631,N_11315);
nor U12593 (N_12593,N_9740,N_11778);
and U12594 (N_12594,N_10818,N_9694);
nand U12595 (N_12595,N_11869,N_11797);
or U12596 (N_12596,N_11827,N_9788);
xor U12597 (N_12597,N_11344,N_9369);
and U12598 (N_12598,N_10006,N_9585);
nand U12599 (N_12599,N_10313,N_11984);
xnor U12600 (N_12600,N_11048,N_11756);
nand U12601 (N_12601,N_11589,N_9968);
nor U12602 (N_12602,N_9422,N_10691);
nand U12603 (N_12603,N_10162,N_11971);
or U12604 (N_12604,N_9150,N_9242);
nand U12605 (N_12605,N_9982,N_10041);
nor U12606 (N_12606,N_11362,N_9087);
nor U12607 (N_12607,N_10085,N_9511);
or U12608 (N_12608,N_10642,N_11859);
nor U12609 (N_12609,N_10042,N_11014);
nor U12610 (N_12610,N_11009,N_9290);
or U12611 (N_12611,N_11438,N_9036);
nand U12612 (N_12612,N_11721,N_11742);
or U12613 (N_12613,N_9849,N_11296);
nand U12614 (N_12614,N_10007,N_10592);
or U12615 (N_12615,N_9411,N_10678);
xnor U12616 (N_12616,N_10178,N_11117);
nand U12617 (N_12617,N_9626,N_9918);
nor U12618 (N_12618,N_9119,N_11794);
nand U12619 (N_12619,N_10359,N_10671);
nand U12620 (N_12620,N_10412,N_11895);
nor U12621 (N_12621,N_11496,N_9807);
nand U12622 (N_12622,N_9267,N_11917);
and U12623 (N_12623,N_10277,N_11526);
or U12624 (N_12624,N_10021,N_9662);
nor U12625 (N_12625,N_10316,N_11309);
or U12626 (N_12626,N_10826,N_9460);
or U12627 (N_12627,N_10250,N_9752);
nor U12628 (N_12628,N_9013,N_10149);
nor U12629 (N_12629,N_10210,N_9225);
nand U12630 (N_12630,N_11491,N_11611);
nor U12631 (N_12631,N_9262,N_10688);
nor U12632 (N_12632,N_10790,N_9355);
or U12633 (N_12633,N_9839,N_9354);
and U12634 (N_12634,N_9101,N_10334);
or U12635 (N_12635,N_11835,N_11016);
nor U12636 (N_12636,N_10545,N_9545);
nand U12637 (N_12637,N_11788,N_10212);
and U12638 (N_12638,N_9042,N_9321);
nand U12639 (N_12639,N_9945,N_11997);
nand U12640 (N_12640,N_10308,N_10355);
and U12641 (N_12641,N_9427,N_11990);
and U12642 (N_12642,N_10154,N_10246);
and U12643 (N_12643,N_10236,N_9680);
nor U12644 (N_12644,N_10057,N_9444);
and U12645 (N_12645,N_10547,N_11102);
and U12646 (N_12646,N_11669,N_10828);
nor U12647 (N_12647,N_10627,N_10365);
or U12648 (N_12648,N_11710,N_11692);
and U12649 (N_12649,N_11519,N_10487);
nor U12650 (N_12650,N_9716,N_11775);
and U12651 (N_12651,N_9527,N_11208);
or U12652 (N_12652,N_10008,N_11715);
or U12653 (N_12653,N_11897,N_11142);
xor U12654 (N_12654,N_11430,N_10034);
or U12655 (N_12655,N_9412,N_10473);
nand U12656 (N_12656,N_11239,N_11573);
and U12657 (N_12657,N_10674,N_11832);
nor U12658 (N_12658,N_9143,N_9642);
xor U12659 (N_12659,N_11367,N_10760);
and U12660 (N_12660,N_9176,N_10174);
xnor U12661 (N_12661,N_11088,N_11011);
nand U12662 (N_12662,N_9803,N_9891);
nor U12663 (N_12663,N_10836,N_9074);
nor U12664 (N_12664,N_10269,N_9781);
nor U12665 (N_12665,N_10766,N_10472);
nand U12666 (N_12666,N_11060,N_9505);
xnor U12667 (N_12667,N_11322,N_9437);
xor U12668 (N_12668,N_11250,N_10451);
or U12669 (N_12669,N_11738,N_9397);
or U12670 (N_12670,N_9147,N_11553);
or U12671 (N_12671,N_10981,N_9755);
nor U12672 (N_12672,N_10967,N_9328);
nand U12673 (N_12673,N_9360,N_10892);
nor U12674 (N_12674,N_11585,N_11564);
or U12675 (N_12675,N_10675,N_11274);
and U12676 (N_12676,N_10862,N_9732);
nand U12677 (N_12677,N_11455,N_9421);
nor U12678 (N_12678,N_11465,N_9207);
xnor U12679 (N_12679,N_11260,N_9464);
or U12680 (N_12680,N_9550,N_9382);
xnor U12681 (N_12681,N_11043,N_10328);
and U12682 (N_12682,N_11942,N_9555);
nand U12683 (N_12683,N_10605,N_11445);
and U12684 (N_12684,N_10764,N_10061);
and U12685 (N_12685,N_9695,N_10194);
nor U12686 (N_12686,N_11602,N_9836);
or U12687 (N_12687,N_10056,N_11071);
nor U12688 (N_12688,N_11606,N_11571);
or U12689 (N_12689,N_10474,N_9237);
and U12690 (N_12690,N_11607,N_10441);
nand U12691 (N_12691,N_11290,N_9737);
or U12692 (N_12692,N_10954,N_11884);
nor U12693 (N_12693,N_10667,N_11194);
and U12694 (N_12694,N_9873,N_9388);
nand U12695 (N_12695,N_9793,N_10373);
and U12696 (N_12696,N_9128,N_11227);
nand U12697 (N_12697,N_11961,N_11694);
nand U12698 (N_12698,N_9772,N_10927);
or U12699 (N_12699,N_10783,N_11851);
or U12700 (N_12700,N_9814,N_10608);
xor U12701 (N_12701,N_11591,N_11512);
nand U12702 (N_12702,N_11421,N_11557);
xor U12703 (N_12703,N_10629,N_11002);
or U12704 (N_12704,N_9507,N_9357);
and U12705 (N_12705,N_10206,N_9432);
or U12706 (N_12706,N_9724,N_9572);
nand U12707 (N_12707,N_10534,N_10583);
and U12708 (N_12708,N_10517,N_9446);
nand U12709 (N_12709,N_9989,N_10885);
or U12710 (N_12710,N_11853,N_11627);
or U12711 (N_12711,N_11941,N_11708);
or U12712 (N_12712,N_9109,N_11005);
and U12713 (N_12713,N_11074,N_11608);
and U12714 (N_12714,N_11718,N_10168);
or U12715 (N_12715,N_9287,N_11975);
or U12716 (N_12716,N_11291,N_9846);
nand U12717 (N_12717,N_10091,N_10681);
and U12718 (N_12718,N_9209,N_9312);
nand U12719 (N_12719,N_10977,N_10416);
nand U12720 (N_12720,N_11444,N_11073);
nor U12721 (N_12721,N_9818,N_9385);
and U12722 (N_12722,N_11150,N_11622);
nand U12723 (N_12723,N_10664,N_11863);
nor U12724 (N_12724,N_10267,N_11000);
nor U12725 (N_12725,N_11283,N_10512);
and U12726 (N_12726,N_11096,N_9841);
nor U12727 (N_12727,N_10463,N_11624);
and U12728 (N_12728,N_11408,N_10184);
nand U12729 (N_12729,N_9523,N_10216);
xnor U12730 (N_12730,N_10529,N_9393);
or U12731 (N_12731,N_9986,N_11017);
nand U12732 (N_12732,N_11836,N_10676);
nand U12733 (N_12733,N_11628,N_9979);
or U12734 (N_12734,N_10854,N_10385);
nor U12735 (N_12735,N_9567,N_11133);
nand U12736 (N_12736,N_11424,N_9723);
and U12737 (N_12737,N_10659,N_10247);
nand U12738 (N_12738,N_11214,N_10800);
xor U12739 (N_12739,N_10070,N_9708);
nor U12740 (N_12740,N_10442,N_10172);
xnor U12741 (N_12741,N_9767,N_9322);
and U12742 (N_12742,N_9370,N_9257);
or U12743 (N_12743,N_10791,N_11170);
and U12744 (N_12744,N_10374,N_11516);
nor U12745 (N_12745,N_11332,N_9992);
nand U12746 (N_12746,N_11763,N_10960);
xnor U12747 (N_12747,N_10338,N_9586);
and U12748 (N_12748,N_9191,N_10483);
and U12749 (N_12749,N_11003,N_9469);
nand U12750 (N_12750,N_10040,N_9862);
nor U12751 (N_12751,N_10698,N_11812);
or U12752 (N_12752,N_10558,N_11268);
nor U12753 (N_12753,N_9822,N_9884);
and U12754 (N_12754,N_9565,N_10552);
nor U12755 (N_12755,N_11007,N_9308);
or U12756 (N_12756,N_9457,N_11749);
or U12757 (N_12757,N_10350,N_11157);
nor U12758 (N_12758,N_9137,N_10301);
nor U12759 (N_12759,N_9924,N_9760);
xor U12760 (N_12760,N_11303,N_10058);
xor U12761 (N_12761,N_11818,N_9327);
or U12762 (N_12762,N_11162,N_10426);
xnor U12763 (N_12763,N_10290,N_10884);
and U12764 (N_12764,N_10012,N_10911);
and U12765 (N_12765,N_10805,N_10074);
or U12766 (N_12766,N_11764,N_9034);
xor U12767 (N_12767,N_10465,N_9219);
nand U12768 (N_12768,N_9898,N_11904);
nor U12769 (N_12769,N_10413,N_11787);
and U12770 (N_12770,N_9341,N_11800);
or U12771 (N_12771,N_10303,N_11431);
nand U12772 (N_12772,N_10653,N_9008);
and U12773 (N_12773,N_10420,N_11259);
nor U12774 (N_12774,N_9860,N_11184);
or U12775 (N_12775,N_11924,N_11503);
nor U12776 (N_12776,N_9273,N_9763);
nand U12777 (N_12777,N_9307,N_10909);
nand U12778 (N_12778,N_10565,N_9172);
nand U12779 (N_12779,N_9817,N_10330);
and U12780 (N_12780,N_10899,N_11960);
and U12781 (N_12781,N_10867,N_11594);
or U12782 (N_12782,N_10405,N_11021);
nor U12783 (N_12783,N_10115,N_9110);
xor U12784 (N_12784,N_9115,N_9203);
or U12785 (N_12785,N_11530,N_10351);
or U12786 (N_12786,N_11792,N_10507);
and U12787 (N_12787,N_9932,N_9152);
nor U12788 (N_12788,N_10073,N_11674);
nand U12789 (N_12789,N_11161,N_10738);
xor U12790 (N_12790,N_9922,N_9248);
or U12791 (N_12791,N_10265,N_11212);
and U12792 (N_12792,N_11213,N_9291);
nand U12793 (N_12793,N_11347,N_10048);
nand U12794 (N_12794,N_9288,N_11083);
nor U12795 (N_12795,N_11809,N_11395);
nor U12796 (N_12796,N_11831,N_11446);
or U12797 (N_12797,N_10564,N_11654);
nand U12798 (N_12798,N_9597,N_9786);
xnor U12799 (N_12799,N_11668,N_10356);
or U12800 (N_12800,N_11717,N_9955);
and U12801 (N_12801,N_11119,N_9727);
nand U12802 (N_12802,N_11324,N_11659);
or U12803 (N_12803,N_11233,N_11544);
nand U12804 (N_12804,N_10432,N_10183);
nor U12805 (N_12805,N_9076,N_9484);
nand U12806 (N_12806,N_11581,N_11295);
or U12807 (N_12807,N_10570,N_11649);
and U12808 (N_12808,N_10917,N_9904);
nor U12809 (N_12809,N_10985,N_9334);
and U12810 (N_12810,N_11913,N_10611);
or U12811 (N_12811,N_9428,N_10841);
or U12812 (N_12812,N_10949,N_10164);
or U12813 (N_12813,N_9211,N_11141);
or U12814 (N_12814,N_10538,N_11206);
and U12815 (N_12815,N_9089,N_11525);
or U12816 (N_12816,N_9677,N_10224);
and U12817 (N_12817,N_10958,N_9663);
nand U12818 (N_12818,N_10231,N_10086);
nand U12819 (N_12819,N_9040,N_9625);
nor U12820 (N_12820,N_11838,N_10182);
and U12821 (N_12821,N_9735,N_11498);
or U12822 (N_12822,N_11420,N_10658);
nor U12823 (N_12823,N_11232,N_9024);
or U12824 (N_12824,N_10376,N_10177);
xor U12825 (N_12825,N_11840,N_10103);
nor U12826 (N_12826,N_10858,N_9596);
or U12827 (N_12827,N_9746,N_9365);
nor U12828 (N_12828,N_9085,N_10191);
and U12829 (N_12829,N_9425,N_11436);
nand U12830 (N_12830,N_11719,N_9730);
or U12831 (N_12831,N_10459,N_9055);
nand U12832 (N_12832,N_9867,N_9282);
nand U12833 (N_12833,N_9156,N_9882);
or U12834 (N_12834,N_11665,N_9243);
and U12835 (N_12835,N_9007,N_11336);
and U12836 (N_12836,N_11218,N_10458);
or U12837 (N_12837,N_9009,N_11944);
or U12838 (N_12838,N_10279,N_9340);
nand U12839 (N_12839,N_10780,N_9232);
nand U12840 (N_12840,N_9458,N_10114);
and U12841 (N_12841,N_9496,N_11385);
nor U12842 (N_12842,N_10600,N_9821);
and U12843 (N_12843,N_10260,N_10408);
or U12844 (N_12844,N_11196,N_10486);
nor U12845 (N_12845,N_9580,N_11008);
and U12846 (N_12846,N_10857,N_11641);
and U12847 (N_12847,N_11983,N_10118);
and U12848 (N_12848,N_10695,N_10477);
or U12849 (N_12849,N_10130,N_9726);
xor U12850 (N_12850,N_10488,N_10400);
or U12851 (N_12851,N_11509,N_10098);
and U12852 (N_12852,N_9946,N_10707);
and U12853 (N_12853,N_9454,N_10572);
xor U12854 (N_12854,N_9779,N_9967);
and U12855 (N_12855,N_10868,N_11670);
nor U12856 (N_12856,N_10032,N_9681);
nand U12857 (N_12857,N_11755,N_10532);
nor U12858 (N_12858,N_10521,N_10871);
xor U12859 (N_12859,N_11545,N_10571);
nand U12860 (N_12860,N_11337,N_10112);
or U12861 (N_12861,N_11228,N_11346);
xnor U12862 (N_12862,N_10796,N_11820);
nor U12863 (N_12863,N_11551,N_11877);
and U12864 (N_12864,N_9722,N_10621);
nor U12865 (N_12865,N_11025,N_10921);
nand U12866 (N_12866,N_11675,N_10594);
or U12867 (N_12867,N_10704,N_10018);
xor U12868 (N_12868,N_11063,N_10346);
nand U12869 (N_12869,N_9712,N_9789);
or U12870 (N_12870,N_11123,N_10719);
and U12871 (N_12871,N_9489,N_11513);
nand U12872 (N_12872,N_9396,N_10628);
nor U12873 (N_12873,N_11297,N_11348);
nor U12874 (N_12874,N_10731,N_10740);
nand U12875 (N_12875,N_9896,N_10774);
and U12876 (N_12876,N_10004,N_10566);
and U12877 (N_12877,N_11147,N_9035);
nand U12878 (N_12878,N_11020,N_9320);
and U12879 (N_12879,N_10630,N_9850);
or U12880 (N_12880,N_11396,N_9468);
nand U12881 (N_12881,N_9832,N_10575);
xor U12882 (N_12882,N_9084,N_11252);
nand U12883 (N_12883,N_9883,N_9969);
xnor U12884 (N_12884,N_9611,N_11407);
xor U12885 (N_12885,N_10464,N_10014);
nor U12886 (N_12886,N_9091,N_10786);
or U12887 (N_12887,N_9890,N_9562);
xor U12888 (N_12888,N_10502,N_11560);
and U12889 (N_12889,N_9037,N_9153);
xnor U12890 (N_12890,N_11019,N_10672);
xnor U12891 (N_12891,N_10419,N_11576);
nor U12892 (N_12892,N_9180,N_9954);
and U12893 (N_12893,N_9541,N_10848);
or U12894 (N_12894,N_10709,N_11796);
nand U12895 (N_12895,N_11968,N_10381);
nor U12896 (N_12896,N_10905,N_10367);
or U12897 (N_12897,N_9368,N_11620);
or U12898 (N_12898,N_11726,N_11195);
and U12899 (N_12899,N_10749,N_10589);
and U12900 (N_12900,N_10140,N_10104);
or U12901 (N_12901,N_10587,N_10046);
xnor U12902 (N_12902,N_10944,N_11139);
or U12903 (N_12903,N_9266,N_11588);
or U12904 (N_12904,N_11599,N_10414);
and U12905 (N_12905,N_9985,N_9930);
nand U12906 (N_12906,N_9902,N_10335);
or U12907 (N_12907,N_9540,N_11555);
nand U12908 (N_12908,N_10843,N_9734);
nand U12909 (N_12909,N_9206,N_9892);
or U12910 (N_12910,N_11023,N_10315);
and U12911 (N_12911,N_11619,N_11079);
or U12912 (N_12912,N_10724,N_10941);
nand U12913 (N_12913,N_9419,N_10875);
or U12914 (N_12914,N_9361,N_11745);
nand U12915 (N_12915,N_11052,N_11650);
and U12916 (N_12916,N_9670,N_11339);
nor U12917 (N_12917,N_9823,N_9201);
nor U12918 (N_12918,N_11053,N_11056);
or U12919 (N_12919,N_9343,N_9158);
nor U12920 (N_12920,N_10037,N_9819);
xnor U12921 (N_12921,N_9044,N_11871);
xnor U12922 (N_12922,N_11510,N_9260);
or U12923 (N_12923,N_10181,N_10623);
and U12924 (N_12924,N_9709,N_11242);
xnor U12925 (N_12925,N_10820,N_9086);
xor U12926 (N_12926,N_11793,N_11887);
or U12927 (N_12927,N_9294,N_11258);
nor U12928 (N_12928,N_11476,N_11899);
nand U12929 (N_12929,N_10770,N_9482);
nor U12930 (N_12930,N_11772,N_10490);
and U12931 (N_12931,N_10341,N_11713);
nand U12932 (N_12932,N_10613,N_9988);
and U12933 (N_12933,N_9519,N_10891);
nand U12934 (N_12934,N_10440,N_9155);
or U12935 (N_12935,N_10233,N_9310);
xnor U12936 (N_12936,N_10849,N_10835);
nand U12937 (N_12937,N_11565,N_9406);
and U12938 (N_12938,N_9372,N_11705);
nand U12939 (N_12939,N_9859,N_11808);
or U12940 (N_12940,N_11558,N_10806);
xnor U12941 (N_12941,N_11112,N_9509);
nand U12942 (N_12942,N_9629,N_11062);
nor U12943 (N_12943,N_10326,N_10785);
nand U12944 (N_12944,N_9404,N_10804);
and U12945 (N_12945,N_10013,N_11992);
xnor U12946 (N_12946,N_11949,N_9566);
nand U12947 (N_12947,N_10801,N_10391);
and U12948 (N_12948,N_10591,N_11149);
nor U12949 (N_12949,N_11167,N_11383);
and U12950 (N_12950,N_11244,N_9235);
and U12951 (N_12951,N_10511,N_10520);
nand U12952 (N_12952,N_10293,N_11031);
or U12953 (N_12953,N_11460,N_10651);
nand U12954 (N_12954,N_9303,N_11737);
and U12955 (N_12955,N_11652,N_9331);
or U12956 (N_12956,N_10975,N_10455);
nor U12957 (N_12957,N_10150,N_10649);
or U12958 (N_12958,N_10943,N_9518);
nor U12959 (N_12959,N_9476,N_11858);
xor U12960 (N_12960,N_11845,N_11814);
nand U12961 (N_12961,N_9762,N_9401);
nor U12962 (N_12962,N_9650,N_10913);
or U12963 (N_12963,N_9220,N_10399);
nor U12964 (N_12964,N_10323,N_9298);
or U12965 (N_12965,N_10620,N_9868);
and U12966 (N_12966,N_9741,N_11698);
nand U12967 (N_12967,N_9653,N_10030);
and U12968 (N_12968,N_11672,N_10622);
nand U12969 (N_12969,N_9991,N_11934);
nand U12970 (N_12970,N_9277,N_11938);
nand U12971 (N_12971,N_11795,N_9346);
nand U12972 (N_12972,N_10102,N_10901);
and U12973 (N_12973,N_11487,N_10011);
nor U12974 (N_12974,N_11201,N_11584);
xnor U12975 (N_12975,N_9325,N_11839);
nand U12976 (N_12976,N_10625,N_9594);
or U12977 (N_12977,N_9032,N_9111);
and U12978 (N_12978,N_10509,N_10431);
nor U12979 (N_12979,N_10329,N_9390);
nand U12980 (N_12980,N_10485,N_9815);
and U12981 (N_12981,N_9066,N_10361);
or U12982 (N_12982,N_10364,N_9880);
or U12983 (N_12983,N_10496,N_9135);
nor U12984 (N_12984,N_10711,N_10325);
and U12985 (N_12985,N_10639,N_10501);
and U12986 (N_12986,N_9627,N_10370);
and U12987 (N_12987,N_11372,N_10435);
or U12988 (N_12988,N_11330,N_11366);
and U12989 (N_12989,N_11229,N_10271);
xor U12990 (N_12990,N_10429,N_10500);
and U12991 (N_12991,N_11026,N_11635);
and U12992 (N_12992,N_10752,N_10543);
or U12993 (N_12993,N_11919,N_9542);
nand U12994 (N_12994,N_11485,N_9547);
and U12995 (N_12995,N_10108,N_10092);
nor U12996 (N_12996,N_10446,N_11461);
and U12997 (N_12997,N_9997,N_9443);
or U12998 (N_12998,N_10371,N_11483);
and U12999 (N_12999,N_10877,N_10023);
or U13000 (N_13000,N_10706,N_9554);
nand U13001 (N_13001,N_11100,N_11617);
or U13002 (N_13002,N_10015,N_9616);
nor U13003 (N_13003,N_9897,N_10929);
nand U13004 (N_13004,N_9030,N_9409);
xor U13005 (N_13005,N_11854,N_9957);
nand U13006 (N_13006,N_11701,N_11159);
and U13007 (N_13007,N_10987,N_10915);
and U13008 (N_13008,N_9693,N_9229);
nor U13009 (N_13009,N_10421,N_10606);
nand U13010 (N_13010,N_10965,N_10755);
and U13011 (N_13011,N_10957,N_10747);
xor U13012 (N_13012,N_11965,N_11471);
and U13013 (N_13013,N_11881,N_10384);
nor U13014 (N_13014,N_11479,N_11202);
or U13015 (N_13015,N_9264,N_11037);
and U13016 (N_13016,N_11075,N_9987);
xnor U13017 (N_13017,N_11923,N_10716);
and U13018 (N_13018,N_11524,N_10886);
nand U13019 (N_13019,N_10000,N_9043);
nand U13020 (N_13020,N_11432,N_9895);
nand U13021 (N_13021,N_10001,N_10993);
or U13022 (N_13022,N_9192,N_11462);
or U13023 (N_13023,N_9514,N_9776);
or U13024 (N_13024,N_9474,N_11685);
xor U13025 (N_13025,N_9827,N_11091);
nand U13026 (N_13026,N_10713,N_10199);
or U13027 (N_13027,N_10763,N_11390);
and U13028 (N_13028,N_9936,N_11921);
xnor U13029 (N_13029,N_11328,N_10498);
and U13030 (N_13030,N_10298,N_10694);
nand U13031 (N_13031,N_9563,N_11931);
nor U13032 (N_13032,N_9281,N_9858);
and U13033 (N_13033,N_10255,N_9188);
and U13034 (N_13034,N_11537,N_11909);
nand U13035 (N_13035,N_9804,N_11013);
and U13036 (N_13036,N_11872,N_10084);
and U13037 (N_13037,N_10972,N_11825);
nor U13038 (N_13038,N_11875,N_9424);
nand U13039 (N_13039,N_10795,N_9510);
nor U13040 (N_13040,N_10227,N_10976);
nand U13041 (N_13041,N_9600,N_10910);
and U13042 (N_13042,N_10090,N_11561);
or U13043 (N_13043,N_11813,N_11989);
nand U13044 (N_13044,N_10656,N_10604);
xor U13045 (N_13045,N_11038,N_9641);
xor U13046 (N_13046,N_11958,N_9259);
xor U13047 (N_13047,N_9940,N_11753);
and U13048 (N_13048,N_10163,N_9375);
nor U13049 (N_13049,N_11805,N_11193);
and U13050 (N_13050,N_9933,N_10643);
nor U13051 (N_13051,N_9654,N_10908);
or U13052 (N_13052,N_9943,N_9881);
xor U13053 (N_13053,N_10787,N_11199);
nor U13054 (N_13054,N_11677,N_9865);
xor U13055 (N_13055,N_10468,N_10148);
and U13056 (N_13056,N_11976,N_9423);
nand U13057 (N_13057,N_10757,N_11405);
or U13058 (N_13058,N_11554,N_10285);
nor U13059 (N_13059,N_11416,N_11633);
nand U13060 (N_13060,N_10751,N_9791);
nand U13061 (N_13061,N_11033,N_9493);
or U13062 (N_13062,N_11341,N_10555);
or U13063 (N_13063,N_9353,N_9125);
nor U13064 (N_13064,N_9215,N_9297);
nand U13065 (N_13065,N_9610,N_11704);
nand U13066 (N_13066,N_10966,N_11647);
and U13067 (N_13067,N_9635,N_9619);
nor U13068 (N_13068,N_9976,N_10702);
nor U13069 (N_13069,N_9704,N_10170);
or U13070 (N_13070,N_9648,N_9318);
and U13071 (N_13071,N_9780,N_11216);
nand U13072 (N_13072,N_9413,N_11570);
nor U13073 (N_13073,N_10980,N_9302);
nand U13074 (N_13074,N_11497,N_11892);
nand U13075 (N_13075,N_11394,N_11210);
or U13076 (N_13076,N_11464,N_11371);
nor U13077 (N_13077,N_9348,N_9004);
nand U13078 (N_13078,N_9775,N_11453);
nor U13079 (N_13079,N_10179,N_11343);
nor U13080 (N_13080,N_9742,N_9122);
nor U13081 (N_13081,N_11799,N_10375);
nor U13082 (N_13082,N_9064,N_10406);
nor U13083 (N_13083,N_9535,N_10768);
or U13084 (N_13084,N_11907,N_10484);
and U13085 (N_13085,N_11937,N_9974);
xnor U13086 (N_13086,N_11667,N_9405);
and U13087 (N_13087,N_9339,N_9790);
nor U13088 (N_13088,N_10016,N_11879);
and U13089 (N_13089,N_9377,N_9931);
nor U13090 (N_13090,N_9197,N_9887);
and U13091 (N_13091,N_9614,N_9099);
or U13092 (N_13092,N_11508,N_9782);
nand U13093 (N_13093,N_9171,N_9317);
and U13094 (N_13094,N_11640,N_10135);
nor U13095 (N_13095,N_10282,N_11972);
xor U13096 (N_13096,N_9958,N_11387);
nand U13097 (N_13097,N_9739,N_9878);
nor U13098 (N_13098,N_10302,N_10809);
nor U13099 (N_13099,N_10504,N_10454);
or U13100 (N_13100,N_10159,N_9472);
or U13101 (N_13101,N_10668,N_9603);
and U13102 (N_13102,N_11137,N_11939);
xor U13103 (N_13103,N_11595,N_11450);
nand U13104 (N_13104,N_10673,N_10652);
or U13105 (N_13105,N_9553,N_11625);
nand U13106 (N_13106,N_11773,N_11637);
and U13107 (N_13107,N_9164,N_9403);
and U13108 (N_13108,N_9083,N_11489);
or U13109 (N_13109,N_9657,N_9971);
nor U13110 (N_13110,N_10817,N_11146);
or U13111 (N_13111,N_11711,N_11154);
or U13112 (N_13112,N_9081,N_11298);
or U13113 (N_13113,N_9394,N_9769);
nand U13114 (N_13114,N_10970,N_9561);
and U13115 (N_13115,N_9250,N_9082);
or U13116 (N_13116,N_11335,N_10816);
nand U13117 (N_13117,N_9254,N_11612);
or U13118 (N_13118,N_11402,N_11696);
nor U13119 (N_13119,N_9990,N_11413);
or U13120 (N_13120,N_11238,N_11065);
nand U13121 (N_13121,N_9758,N_9688);
nor U13122 (N_13122,N_9661,N_10580);
and U13123 (N_13123,N_9963,N_10938);
nand U13124 (N_13124,N_11680,N_11363);
or U13125 (N_13125,N_10264,N_10201);
nand U13126 (N_13126,N_10939,N_9532);
or U13127 (N_13127,N_11767,N_9669);
nor U13128 (N_13128,N_9311,N_9549);
nor U13129 (N_13129,N_11786,N_10196);
or U13130 (N_13130,N_11275,N_9624);
xor U13131 (N_13131,N_10721,N_11172);
or U13132 (N_13132,N_11653,N_10961);
nand U13133 (N_13133,N_9937,N_9744);
or U13134 (N_13134,N_9748,N_11963);
nor U13135 (N_13135,N_10240,N_11695);
or U13136 (N_13136,N_11393,N_10387);
nand U13137 (N_13137,N_10107,N_10893);
nand U13138 (N_13138,N_10010,N_11666);
or U13139 (N_13139,N_10291,N_10324);
and U13140 (N_13140,N_9141,N_10708);
nand U13141 (N_13141,N_11969,N_9410);
or U13142 (N_13142,N_10990,N_11598);
nor U13143 (N_13143,N_10973,N_11723);
xor U13144 (N_13144,N_11947,N_11406);
nand U13145 (N_13145,N_9359,N_11882);
or U13146 (N_13146,N_10530,N_11798);
or U13147 (N_13147,N_10533,N_11109);
or U13148 (N_13148,N_10692,N_9830);
nor U13149 (N_13149,N_9534,N_10368);
nand U13150 (N_13150,N_11380,N_11682);
and U13151 (N_13151,N_10466,N_9959);
or U13152 (N_13152,N_10793,N_11153);
and U13153 (N_13153,N_11200,N_11155);
xnor U13154 (N_13154,N_11419,N_11163);
nand U13155 (N_13155,N_11099,N_9117);
nor U13156 (N_13156,N_9785,N_11185);
or U13157 (N_13157,N_9628,N_11035);
and U13158 (N_13158,N_10300,N_10519);
nor U13159 (N_13159,N_11760,N_10136);
xnor U13160 (N_13160,N_9533,N_10195);
and U13161 (N_13161,N_10612,N_10550);
or U13162 (N_13162,N_10771,N_11948);
nand U13163 (N_13163,N_9190,N_10646);
and U13164 (N_13164,N_11103,N_11121);
and U13165 (N_13165,N_9408,N_9492);
or U13166 (N_13166,N_11833,N_9214);
and U13167 (N_13167,N_11734,N_9692);
and U13168 (N_13168,N_11867,N_10906);
or U13169 (N_13169,N_9435,N_10697);
and U13170 (N_13170,N_10318,N_10655);
or U13171 (N_13171,N_9386,N_11051);
or U13172 (N_13172,N_9031,N_11590);
nand U13173 (N_13173,N_9977,N_11361);
nor U13174 (N_13174,N_9649,N_11874);
nor U13175 (N_13175,N_11908,N_9395);
or U13176 (N_13176,N_9517,N_11684);
and U13177 (N_13177,N_10815,N_10189);
nand U13178 (N_13178,N_10095,N_9768);
and U13179 (N_13179,N_9161,N_9487);
xnor U13180 (N_13180,N_11098,N_9687);
and U13181 (N_13181,N_11105,N_11389);
nor U13182 (N_13182,N_9928,N_10139);
nor U13183 (N_13183,N_11505,N_10203);
nand U13184 (N_13184,N_11044,N_10065);
or U13185 (N_13185,N_11974,N_11810);
or U13186 (N_13186,N_10143,N_11547);
or U13187 (N_13187,N_11495,N_10823);
nand U13188 (N_13188,N_9673,N_9057);
nand U13189 (N_13189,N_11521,N_10424);
or U13190 (N_13190,N_9194,N_11293);
and U13191 (N_13191,N_11466,N_10528);
nor U13192 (N_13192,N_11876,N_11866);
nor U13193 (N_13193,N_9473,N_11639);
nor U13194 (N_13194,N_11262,N_10344);
xor U13195 (N_13195,N_11673,N_10220);
nand U13196 (N_13196,N_9713,N_10452);
nor U13197 (N_13197,N_9729,N_11973);
nand U13198 (N_13198,N_10699,N_9104);
nor U13199 (N_13199,N_9981,N_10433);
nand U13200 (N_13200,N_9471,N_11724);
or U13201 (N_13201,N_9975,N_9417);
or U13202 (N_13202,N_10513,N_9757);
and U13203 (N_13203,N_10825,N_9389);
nand U13204 (N_13204,N_10275,N_10772);
nor U13205 (N_13205,N_9011,N_9184);
and U13206 (N_13206,N_11480,N_11981);
xor U13207 (N_13207,N_11690,N_9996);
nand U13208 (N_13208,N_11864,N_11045);
xor U13209 (N_13209,N_9450,N_11712);
nor U13210 (N_13210,N_11746,N_10644);
xor U13211 (N_13211,N_9631,N_10146);
nand U13212 (N_13212,N_11815,N_10515);
nand U13213 (N_13213,N_11714,N_9352);
or U13214 (N_13214,N_10631,N_9871);
nor U13215 (N_13215,N_11092,N_9984);
or U13216 (N_13216,N_9888,N_9771);
xor U13217 (N_13217,N_9864,N_9749);
and U13218 (N_13218,N_10069,N_11057);
xnor U13219 (N_13219,N_9028,N_9886);
or U13220 (N_13220,N_9581,N_10861);
or U13221 (N_13221,N_9647,N_9434);
and U13222 (N_13222,N_10252,N_9556);
or U13223 (N_13223,N_11418,N_10109);
nor U13224 (N_13224,N_11656,N_11120);
and U13225 (N_13225,N_11312,N_11084);
or U13226 (N_13226,N_11501,N_10799);
nor U13227 (N_13227,N_10187,N_10160);
xnor U13228 (N_13228,N_11977,N_11979);
and U13229 (N_13229,N_11744,N_9524);
nand U13230 (N_13230,N_11085,N_10415);
nor U13231 (N_13231,N_10209,N_10924);
and U13232 (N_13232,N_9136,N_11660);
xor U13233 (N_13233,N_9166,N_10409);
nor U13234 (N_13234,N_10425,N_9144);
and U13235 (N_13235,N_9274,N_9634);
nor U13236 (N_13236,N_10837,N_10295);
and U13237 (N_13237,N_9330,N_11896);
xnor U13238 (N_13238,N_9686,N_11548);
nand U13239 (N_13239,N_10262,N_11443);
nand U13240 (N_13240,N_9280,N_11765);
nand U13241 (N_13241,N_10278,N_11943);
nand U13242 (N_13242,N_10256,N_11289);
or U13243 (N_13243,N_11425,N_10063);
nand U13244 (N_13244,N_9075,N_9950);
or U13245 (N_13245,N_9538,N_10989);
or U13246 (N_13246,N_9478,N_10093);
and U13247 (N_13247,N_11357,N_11409);
nor U13248 (N_13248,N_9754,N_9335);
nand U13249 (N_13249,N_9536,N_11614);
xor U13250 (N_13250,N_9333,N_11177);
nand U13251 (N_13251,N_11251,N_11175);
nor U13252 (N_13252,N_10225,N_10728);
or U13253 (N_13253,N_11993,N_11064);
nand U13254 (N_13254,N_11849,N_9218);
and U13255 (N_13255,N_11067,N_9569);
nor U13256 (N_13256,N_10950,N_10834);
nand U13257 (N_13257,N_9238,N_10762);
nor U13258 (N_13258,N_10936,N_10654);
nand U13259 (N_13259,N_9934,N_11215);
xor U13260 (N_13260,N_11299,N_11273);
nand U13261 (N_13261,N_11940,N_10833);
nand U13262 (N_13262,N_10461,N_11151);
or U13263 (N_13263,N_9877,N_9949);
and U13264 (N_13264,N_9017,N_9710);
xor U13265 (N_13265,N_9770,N_9808);
nor U13266 (N_13266,N_10551,N_10052);
nor U13267 (N_13267,N_9491,N_11999);
and U13268 (N_13268,N_11415,N_11514);
nor U13269 (N_13269,N_11114,N_11842);
and U13270 (N_13270,N_10319,N_11211);
or U13271 (N_13271,N_9848,N_9923);
nand U13272 (N_13272,N_10469,N_10151);
and U13273 (N_13273,N_11292,N_9499);
or U13274 (N_13274,N_11094,N_10059);
nand U13275 (N_13275,N_11093,N_10235);
and U13276 (N_13276,N_11110,N_10208);
or U13277 (N_13277,N_11457,N_9316);
or U13278 (N_13278,N_9090,N_9861);
nand U13279 (N_13279,N_11523,N_10935);
and U13280 (N_13280,N_11707,N_10257);
and U13281 (N_13281,N_11334,N_9965);
nand U13282 (N_13282,N_9588,N_11604);
and U13283 (N_13283,N_10734,N_10636);
or U13284 (N_13284,N_11459,N_9045);
nand U13285 (N_13285,N_10094,N_9033);
or U13286 (N_13286,N_10900,N_10831);
nor U13287 (N_13287,N_10169,N_11725);
nand U13288 (N_13288,N_10071,N_9711);
nand U13289 (N_13289,N_11145,N_10516);
and U13290 (N_13290,N_10829,N_10778);
nand U13291 (N_13291,N_10029,N_9021);
or U13292 (N_13292,N_10838,N_9018);
nor U13293 (N_13293,N_11572,N_11178);
and U13294 (N_13294,N_9966,N_10535);
and U13295 (N_13295,N_9420,N_11342);
and U13296 (N_13296,N_11326,N_10609);
and U13297 (N_13297,N_11804,N_9332);
nand U13298 (N_13298,N_11779,N_9833);
and U13299 (N_13299,N_11568,N_9196);
nand U13300 (N_13300,N_10100,N_9615);
xor U13301 (N_13301,N_10590,N_9234);
and U13302 (N_13302,N_9798,N_11240);
and U13303 (N_13303,N_10158,N_11542);
and U13304 (N_13304,N_11998,N_10902);
nor U13305 (N_13305,N_9100,N_11392);
or U13306 (N_13306,N_9646,N_11522);
or U13307 (N_13307,N_10038,N_11770);
or U13308 (N_13308,N_11173,N_9747);
nand U13309 (N_13309,N_10690,N_10448);
or U13310 (N_13310,N_9659,N_11991);
xor U13311 (N_13311,N_10992,N_11536);
and U13312 (N_13312,N_11302,N_10703);
or U13313 (N_13313,N_10217,N_9296);
and U13314 (N_13314,N_9609,N_9725);
or U13315 (N_13315,N_10312,N_11703);
and U13316 (N_13316,N_9001,N_11004);
nand U13317 (N_13317,N_11319,N_10192);
nand U13318 (N_13318,N_11886,N_9869);
or U13319 (N_13319,N_10223,N_10310);
nor U13320 (N_13320,N_10846,N_10204);
nand U13321 (N_13321,N_11532,N_9067);
nand U13322 (N_13322,N_9951,N_11819);
xnor U13323 (N_13323,N_9684,N_9702);
xor U13324 (N_13324,N_11198,N_10794);
or U13325 (N_13325,N_9223,N_10557);
or U13326 (N_13326,N_9314,N_9107);
nand U13327 (N_13327,N_9672,N_9698);
nor U13328 (N_13328,N_11280,N_11190);
and U13329 (N_13329,N_10352,N_10803);
nor U13330 (N_13330,N_9047,N_11429);
nor U13331 (N_13331,N_11423,N_10175);
or U13332 (N_13332,N_9174,N_11995);
nand U13333 (N_13333,N_9345,N_11586);
xor U13334 (N_13334,N_10022,N_10880);
or U13335 (N_13335,N_9133,N_10827);
nand U13336 (N_13336,N_10784,N_9652);
nor U13337 (N_13337,N_10559,N_9617);
and U13338 (N_13338,N_11129,N_11171);
nand U13339 (N_13339,N_10963,N_10576);
xor U13340 (N_13340,N_11535,N_11903);
nand U13341 (N_13341,N_10888,N_10904);
nor U13342 (N_13342,N_11506,N_11358);
nand U13343 (N_13343,N_11927,N_11158);
nand U13344 (N_13344,N_10542,N_11658);
nand U13345 (N_13345,N_10430,N_10518);
and U13346 (N_13346,N_9313,N_9374);
xor U13347 (N_13347,N_10133,N_11077);
and U13348 (N_13348,N_10445,N_9750);
nand U13349 (N_13349,N_9306,N_10851);
or U13350 (N_13350,N_10918,N_9271);
nand U13351 (N_13351,N_9440,N_10161);
nor U13352 (N_13352,N_10377,N_10932);
and U13353 (N_13353,N_11422,N_11463);
and U13354 (N_13354,N_10730,N_9092);
xor U13355 (N_13355,N_10349,N_10549);
or U13356 (N_13356,N_10320,N_9342);
and U13357 (N_13357,N_9129,N_9447);
and U13358 (N_13358,N_10598,N_9706);
and U13359 (N_13359,N_11397,N_9644);
and U13360 (N_13360,N_10633,N_11300);
nand U13361 (N_13361,N_9120,N_9256);
nor U13362 (N_13362,N_10249,N_9908);
nand U13363 (N_13363,N_9601,N_10153);
nor U13364 (N_13364,N_10696,N_10462);
and U13365 (N_13365,N_9907,N_11352);
or U13366 (N_13366,N_10914,N_11270);
or U13367 (N_13367,N_10527,N_10280);
nand U13368 (N_13368,N_9665,N_11391);
nor U13369 (N_13369,N_10028,N_9893);
and U13370 (N_13370,N_11378,N_9516);
and U13371 (N_13371,N_9972,N_10726);
or U13372 (N_13372,N_11490,N_11928);
and U13373 (N_13373,N_9689,N_10211);
or U13374 (N_13374,N_10392,N_11776);
or U13375 (N_13375,N_11727,N_11626);
nand U13376 (N_13376,N_9651,N_10934);
xor U13377 (N_13377,N_10903,N_10005);
or U13378 (N_13378,N_10998,N_9255);
xnor U13379 (N_13379,N_9019,N_9268);
or U13380 (N_13380,N_9301,N_10860);
nor U13381 (N_13381,N_10067,N_10284);
nand U13382 (N_13382,N_11861,N_11894);
or U13383 (N_13383,N_10219,N_11223);
nand U13384 (N_13384,N_10033,N_11131);
or U13385 (N_13385,N_9513,N_11699);
nand U13386 (N_13386,N_11574,N_9376);
nor U13387 (N_13387,N_10926,N_10383);
xnor U13388 (N_13388,N_10388,N_10670);
xnor U13389 (N_13389,N_9671,N_9463);
and U13390 (N_13390,N_10714,N_10229);
or U13391 (N_13391,N_9123,N_10119);
or U13392 (N_13392,N_9699,N_10679);
nand U13393 (N_13393,N_10687,N_10314);
xor U13394 (N_13394,N_11629,N_11587);
or U13395 (N_13395,N_9077,N_10422);
nor U13396 (N_13396,N_9278,N_11284);
nand U13397 (N_13397,N_9797,N_10165);
xnor U13398 (N_13398,N_10439,N_10239);
and U13399 (N_13399,N_10568,N_10524);
nand U13400 (N_13400,N_10839,N_10727);
nand U13401 (N_13401,N_9941,N_10569);
nand U13402 (N_13402,N_10128,N_11187);
nand U13403 (N_13403,N_10873,N_11179);
nor U13404 (N_13404,N_9131,N_9838);
nor U13405 (N_13405,N_10025,N_11676);
or U13406 (N_13406,N_9134,N_11603);
xor U13407 (N_13407,N_9230,N_10660);
nor U13408 (N_13408,N_11916,N_9251);
or U13409 (N_13409,N_9169,N_9863);
or U13410 (N_13410,N_9309,N_11318);
nor U13411 (N_13411,N_9980,N_10982);
nor U13412 (N_13412,N_9525,N_11374);
or U13413 (N_13413,N_10808,N_11106);
or U13414 (N_13414,N_10456,N_9560);
and U13415 (N_13415,N_10125,N_10363);
nand U13416 (N_13416,N_10940,N_11761);
or U13417 (N_13417,N_9025,N_11399);
or U13418 (N_13418,N_11642,N_9929);
and U13419 (N_13419,N_11559,N_11935);
or U13420 (N_13420,N_9069,N_10897);
or U13421 (N_13421,N_10354,N_11534);
nor U13422 (N_13422,N_11467,N_11412);
or U13423 (N_13423,N_9204,N_9221);
and U13424 (N_13424,N_10453,N_11950);
nor U13425 (N_13425,N_9289,N_11807);
or U13426 (N_13426,N_11922,N_10378);
and U13427 (N_13427,N_11683,N_10645);
xnor U13428 (N_13428,N_10813,N_11368);
nor U13429 (N_13429,N_10997,N_11294);
or U13430 (N_13430,N_9947,N_9054);
nand U13431 (N_13431,N_10962,N_9914);
xnor U13432 (N_13432,N_9399,N_9114);
and U13433 (N_13433,N_11754,N_10127);
nand U13434 (N_13434,N_9577,N_10845);
nand U13435 (N_13435,N_9855,N_9508);
nor U13436 (N_13436,N_10403,N_11253);
nor U13437 (N_13437,N_9910,N_11964);
or U13438 (N_13438,N_9323,N_10348);
or U13439 (N_13439,N_11880,N_9407);
nand U13440 (N_13440,N_9993,N_10475);
nor U13441 (N_13441,N_11902,N_10626);
or U13442 (N_13442,N_11915,N_10705);
or U13443 (N_13443,N_10134,N_9442);
xnor U13444 (N_13444,N_9132,N_11697);
nand U13445 (N_13445,N_11246,N_11910);
and U13446 (N_13446,N_10253,N_11540);
nor U13447 (N_13447,N_9795,N_9329);
and U13448 (N_13448,N_11567,N_10700);
nor U13449 (N_13449,N_9717,N_11945);
nand U13450 (N_13450,N_11320,N_9973);
nand U13451 (N_13451,N_9261,N_11741);
or U13452 (N_13452,N_10522,N_9198);
nor U13453 (N_13453,N_9816,N_10887);
or U13454 (N_13454,N_10666,N_9733);
or U13455 (N_13455,N_11049,N_10556);
nand U13456 (N_13456,N_10479,N_9466);
nor U13457 (N_13457,N_9005,N_9690);
nand U13458 (N_13458,N_10427,N_11168);
nor U13459 (N_13459,N_9636,N_9826);
or U13460 (N_13460,N_10205,N_9270);
and U13461 (N_13461,N_11531,N_9027);
or U13462 (N_13462,N_11152,N_11716);
or U13463 (N_13463,N_9667,N_10340);
and U13464 (N_13464,N_11265,N_10540);
nand U13465 (N_13465,N_11345,N_9912);
nand U13466 (N_13466,N_9843,N_10499);
and U13467 (N_13467,N_9876,N_11671);
and U13468 (N_13468,N_9245,N_9674);
or U13469 (N_13469,N_10541,N_11802);
xor U13470 (N_13470,N_10035,N_9613);
nand U13471 (N_13471,N_11458,N_9275);
nor U13472 (N_13472,N_9098,N_10715);
or U13473 (N_13473,N_11082,N_10288);
nor U13474 (N_13474,N_9906,N_10510);
xor U13475 (N_13475,N_11750,N_10395);
nor U13476 (N_13476,N_10680,N_11012);
nor U13477 (N_13477,N_10807,N_9470);
and U13478 (N_13478,N_11237,N_11661);
or U13479 (N_13479,N_10876,N_10920);
and U13480 (N_13480,N_11920,N_9418);
and U13481 (N_13481,N_11186,N_9226);
xor U13482 (N_13482,N_10983,N_9658);
nand U13483 (N_13483,N_9145,N_10850);
and U13484 (N_13484,N_11181,N_9801);
xnor U13485 (N_13485,N_10776,N_10964);
nor U13486 (N_13486,N_9705,N_9857);
and U13487 (N_13487,N_9431,N_9576);
nor U13488 (N_13488,N_9222,N_9810);
and U13489 (N_13489,N_9917,N_11191);
nor U13490 (N_13490,N_11183,N_9970);
and U13491 (N_13491,N_11221,N_9269);
nor U13492 (N_13492,N_9845,N_11533);
nor U13493 (N_13493,N_11047,N_9046);
nor U13494 (N_13494,N_9640,N_9557);
or U13495 (N_13495,N_9639,N_11632);
xnor U13496 (N_13496,N_11373,N_9948);
nor U13497 (N_13497,N_11846,N_10226);
nor U13498 (N_13498,N_10788,N_10142);
and U13499 (N_13499,N_9570,N_10068);
and U13500 (N_13500,N_9844,N_10655);
or U13501 (N_13501,N_10995,N_11520);
nand U13502 (N_13502,N_9878,N_11794);
xor U13503 (N_13503,N_11800,N_10177);
nand U13504 (N_13504,N_9591,N_10838);
xor U13505 (N_13505,N_10924,N_11007);
nand U13506 (N_13506,N_9693,N_9890);
nor U13507 (N_13507,N_11457,N_10643);
nand U13508 (N_13508,N_11553,N_10752);
nand U13509 (N_13509,N_9455,N_9806);
nor U13510 (N_13510,N_9141,N_9522);
nand U13511 (N_13511,N_10064,N_10382);
and U13512 (N_13512,N_11858,N_11073);
xor U13513 (N_13513,N_10157,N_11536);
xor U13514 (N_13514,N_10845,N_9300);
nand U13515 (N_13515,N_9146,N_9853);
and U13516 (N_13516,N_10514,N_11257);
nor U13517 (N_13517,N_10110,N_11083);
or U13518 (N_13518,N_11367,N_11108);
or U13519 (N_13519,N_11360,N_10717);
xnor U13520 (N_13520,N_11726,N_9520);
nor U13521 (N_13521,N_9108,N_9563);
xor U13522 (N_13522,N_10203,N_11773);
and U13523 (N_13523,N_11644,N_11857);
nor U13524 (N_13524,N_11483,N_10027);
or U13525 (N_13525,N_9158,N_9705);
nand U13526 (N_13526,N_11445,N_10905);
nand U13527 (N_13527,N_9853,N_11357);
and U13528 (N_13528,N_11553,N_10053);
and U13529 (N_13529,N_9093,N_11827);
or U13530 (N_13530,N_11598,N_11058);
nand U13531 (N_13531,N_10831,N_10582);
xnor U13532 (N_13532,N_9401,N_9763);
or U13533 (N_13533,N_9084,N_9578);
and U13534 (N_13534,N_10064,N_9601);
or U13535 (N_13535,N_11323,N_9872);
nor U13536 (N_13536,N_9417,N_10028);
or U13537 (N_13537,N_9417,N_11062);
xor U13538 (N_13538,N_9952,N_11566);
nor U13539 (N_13539,N_11414,N_9954);
and U13540 (N_13540,N_9108,N_9415);
and U13541 (N_13541,N_10847,N_10513);
and U13542 (N_13542,N_11434,N_10101);
nor U13543 (N_13543,N_10801,N_9351);
or U13544 (N_13544,N_9879,N_11704);
nand U13545 (N_13545,N_11035,N_10153);
and U13546 (N_13546,N_10757,N_11882);
nor U13547 (N_13547,N_10308,N_10356);
or U13548 (N_13548,N_11294,N_11537);
and U13549 (N_13549,N_9858,N_11128);
and U13550 (N_13550,N_9401,N_11741);
nand U13551 (N_13551,N_9898,N_9891);
and U13552 (N_13552,N_9652,N_11719);
nor U13553 (N_13553,N_10009,N_10500);
or U13554 (N_13554,N_11025,N_9922);
and U13555 (N_13555,N_11932,N_9738);
or U13556 (N_13556,N_10514,N_11846);
and U13557 (N_13557,N_11952,N_9946);
or U13558 (N_13558,N_11840,N_9025);
or U13559 (N_13559,N_10635,N_9162);
nand U13560 (N_13560,N_10209,N_9640);
and U13561 (N_13561,N_11802,N_11487);
nor U13562 (N_13562,N_9029,N_10468);
xnor U13563 (N_13563,N_10787,N_11467);
nor U13564 (N_13564,N_9980,N_9093);
or U13565 (N_13565,N_11876,N_9837);
or U13566 (N_13566,N_11418,N_9761);
nand U13567 (N_13567,N_11066,N_9593);
and U13568 (N_13568,N_9618,N_9936);
and U13569 (N_13569,N_10740,N_10537);
nand U13570 (N_13570,N_9056,N_11782);
xor U13571 (N_13571,N_10345,N_11543);
nand U13572 (N_13572,N_11558,N_10420);
nor U13573 (N_13573,N_9697,N_9832);
and U13574 (N_13574,N_10457,N_10751);
nand U13575 (N_13575,N_11166,N_11297);
and U13576 (N_13576,N_11860,N_11142);
nand U13577 (N_13577,N_11459,N_11000);
and U13578 (N_13578,N_11792,N_10198);
xnor U13579 (N_13579,N_10636,N_11283);
or U13580 (N_13580,N_10922,N_9563);
xor U13581 (N_13581,N_10672,N_10553);
and U13582 (N_13582,N_9364,N_9572);
xnor U13583 (N_13583,N_9315,N_9497);
nor U13584 (N_13584,N_10752,N_9641);
nor U13585 (N_13585,N_10918,N_10670);
nor U13586 (N_13586,N_9195,N_10577);
and U13587 (N_13587,N_9552,N_11232);
nor U13588 (N_13588,N_11307,N_9312);
xor U13589 (N_13589,N_10913,N_10472);
and U13590 (N_13590,N_9743,N_10528);
or U13591 (N_13591,N_10097,N_9529);
nor U13592 (N_13592,N_11020,N_9048);
nor U13593 (N_13593,N_9878,N_9143);
nor U13594 (N_13594,N_10717,N_10217);
xor U13595 (N_13595,N_11844,N_10721);
and U13596 (N_13596,N_9657,N_11571);
xor U13597 (N_13597,N_10205,N_9153);
or U13598 (N_13598,N_9423,N_9024);
or U13599 (N_13599,N_9765,N_11127);
and U13600 (N_13600,N_10606,N_11861);
or U13601 (N_13601,N_9484,N_11506);
or U13602 (N_13602,N_11690,N_10326);
and U13603 (N_13603,N_11596,N_10279);
or U13604 (N_13604,N_11032,N_11244);
and U13605 (N_13605,N_9035,N_9790);
nor U13606 (N_13606,N_11439,N_10076);
xnor U13607 (N_13607,N_11818,N_9177);
xnor U13608 (N_13608,N_9936,N_10741);
or U13609 (N_13609,N_11005,N_9402);
nand U13610 (N_13610,N_9547,N_11042);
or U13611 (N_13611,N_11843,N_10157);
or U13612 (N_13612,N_11731,N_10323);
or U13613 (N_13613,N_10370,N_11936);
nand U13614 (N_13614,N_10993,N_10963);
or U13615 (N_13615,N_10756,N_10529);
or U13616 (N_13616,N_9549,N_9587);
nor U13617 (N_13617,N_11253,N_11762);
nor U13618 (N_13618,N_9729,N_10299);
nor U13619 (N_13619,N_9196,N_10405);
or U13620 (N_13620,N_9384,N_9381);
nand U13621 (N_13621,N_9616,N_10038);
nor U13622 (N_13622,N_10337,N_11856);
and U13623 (N_13623,N_9274,N_9841);
and U13624 (N_13624,N_10773,N_11399);
and U13625 (N_13625,N_11573,N_10479);
and U13626 (N_13626,N_9806,N_11999);
nor U13627 (N_13627,N_9338,N_9799);
nand U13628 (N_13628,N_11021,N_9590);
and U13629 (N_13629,N_9996,N_10446);
nand U13630 (N_13630,N_9800,N_11603);
nand U13631 (N_13631,N_11297,N_11897);
nand U13632 (N_13632,N_10509,N_11242);
nand U13633 (N_13633,N_11709,N_11495);
or U13634 (N_13634,N_9311,N_10429);
nor U13635 (N_13635,N_10119,N_10889);
nand U13636 (N_13636,N_9125,N_11250);
nand U13637 (N_13637,N_9593,N_9068);
nand U13638 (N_13638,N_9926,N_10719);
nand U13639 (N_13639,N_9893,N_11229);
or U13640 (N_13640,N_10217,N_10007);
xor U13641 (N_13641,N_10908,N_10139);
and U13642 (N_13642,N_9302,N_11931);
and U13643 (N_13643,N_11434,N_11926);
or U13644 (N_13644,N_9824,N_9333);
or U13645 (N_13645,N_10790,N_10331);
or U13646 (N_13646,N_9525,N_11913);
or U13647 (N_13647,N_11138,N_9462);
nand U13648 (N_13648,N_9821,N_9006);
and U13649 (N_13649,N_10364,N_10365);
nor U13650 (N_13650,N_10683,N_10321);
or U13651 (N_13651,N_11619,N_10364);
or U13652 (N_13652,N_9301,N_9471);
xnor U13653 (N_13653,N_11979,N_11450);
and U13654 (N_13654,N_10968,N_11854);
and U13655 (N_13655,N_11452,N_11417);
xnor U13656 (N_13656,N_10803,N_11499);
nand U13657 (N_13657,N_11491,N_9471);
or U13658 (N_13658,N_10687,N_10664);
nand U13659 (N_13659,N_11696,N_11494);
and U13660 (N_13660,N_10389,N_10175);
nor U13661 (N_13661,N_10547,N_9847);
or U13662 (N_13662,N_10738,N_9742);
nand U13663 (N_13663,N_10967,N_10083);
nor U13664 (N_13664,N_9721,N_11167);
nor U13665 (N_13665,N_11332,N_11761);
nor U13666 (N_13666,N_11156,N_11014);
and U13667 (N_13667,N_10715,N_11286);
nor U13668 (N_13668,N_9331,N_10814);
or U13669 (N_13669,N_10683,N_10979);
nor U13670 (N_13670,N_11791,N_11904);
and U13671 (N_13671,N_11920,N_10931);
nand U13672 (N_13672,N_10032,N_10354);
nor U13673 (N_13673,N_11470,N_9177);
nand U13674 (N_13674,N_11178,N_11724);
and U13675 (N_13675,N_10262,N_9960);
nor U13676 (N_13676,N_9324,N_11454);
and U13677 (N_13677,N_10370,N_9365);
and U13678 (N_13678,N_10202,N_11603);
nand U13679 (N_13679,N_9796,N_11208);
or U13680 (N_13680,N_9590,N_11252);
or U13681 (N_13681,N_10443,N_9972);
and U13682 (N_13682,N_9339,N_9189);
or U13683 (N_13683,N_11732,N_10691);
or U13684 (N_13684,N_11234,N_10364);
and U13685 (N_13685,N_9079,N_10894);
or U13686 (N_13686,N_10021,N_10509);
nand U13687 (N_13687,N_9561,N_11441);
nand U13688 (N_13688,N_10425,N_10154);
xnor U13689 (N_13689,N_9748,N_11210);
nand U13690 (N_13690,N_11599,N_11898);
xor U13691 (N_13691,N_10908,N_10954);
nor U13692 (N_13692,N_10285,N_11753);
nor U13693 (N_13693,N_9810,N_9874);
nand U13694 (N_13694,N_10162,N_10015);
nor U13695 (N_13695,N_10764,N_10883);
nand U13696 (N_13696,N_11765,N_11282);
and U13697 (N_13697,N_11138,N_11961);
nand U13698 (N_13698,N_9106,N_11244);
nand U13699 (N_13699,N_9275,N_10085);
and U13700 (N_13700,N_10761,N_11512);
xnor U13701 (N_13701,N_11462,N_10659);
or U13702 (N_13702,N_9042,N_9190);
xnor U13703 (N_13703,N_11053,N_11251);
and U13704 (N_13704,N_9652,N_9025);
and U13705 (N_13705,N_11462,N_10351);
xnor U13706 (N_13706,N_9524,N_11609);
and U13707 (N_13707,N_9652,N_11101);
nand U13708 (N_13708,N_10221,N_11518);
xnor U13709 (N_13709,N_10744,N_9694);
and U13710 (N_13710,N_10159,N_9099);
nand U13711 (N_13711,N_11901,N_10108);
nor U13712 (N_13712,N_11829,N_9228);
nand U13713 (N_13713,N_10646,N_9536);
or U13714 (N_13714,N_10513,N_10596);
nand U13715 (N_13715,N_11387,N_10601);
and U13716 (N_13716,N_11709,N_10094);
nand U13717 (N_13717,N_9077,N_10723);
nor U13718 (N_13718,N_10624,N_10565);
nand U13719 (N_13719,N_11628,N_11715);
xnor U13720 (N_13720,N_9534,N_10500);
nand U13721 (N_13721,N_11122,N_9604);
nand U13722 (N_13722,N_10882,N_11773);
nand U13723 (N_13723,N_9021,N_11693);
and U13724 (N_13724,N_10878,N_9389);
or U13725 (N_13725,N_10340,N_9414);
and U13726 (N_13726,N_11309,N_10613);
nor U13727 (N_13727,N_10081,N_10250);
or U13728 (N_13728,N_9878,N_9380);
or U13729 (N_13729,N_11144,N_11798);
nor U13730 (N_13730,N_9821,N_9815);
nor U13731 (N_13731,N_10335,N_11480);
nand U13732 (N_13732,N_11859,N_9380);
and U13733 (N_13733,N_9000,N_9862);
and U13734 (N_13734,N_9192,N_11200);
xnor U13735 (N_13735,N_11849,N_10370);
nor U13736 (N_13736,N_10948,N_10858);
nand U13737 (N_13737,N_11632,N_11793);
nor U13738 (N_13738,N_11062,N_10211);
nor U13739 (N_13739,N_9180,N_11632);
nand U13740 (N_13740,N_10803,N_10789);
and U13741 (N_13741,N_10929,N_10781);
and U13742 (N_13742,N_10306,N_10785);
nor U13743 (N_13743,N_11527,N_11923);
or U13744 (N_13744,N_11048,N_10064);
or U13745 (N_13745,N_11303,N_11143);
nor U13746 (N_13746,N_11475,N_10263);
and U13747 (N_13747,N_10881,N_10817);
nand U13748 (N_13748,N_9216,N_10433);
and U13749 (N_13749,N_10134,N_9676);
nor U13750 (N_13750,N_9473,N_11990);
nor U13751 (N_13751,N_9334,N_9348);
or U13752 (N_13752,N_9584,N_10554);
and U13753 (N_13753,N_10981,N_10119);
xor U13754 (N_13754,N_9305,N_11781);
and U13755 (N_13755,N_11937,N_11735);
nand U13756 (N_13756,N_11909,N_11926);
or U13757 (N_13757,N_10599,N_11388);
or U13758 (N_13758,N_10086,N_9222);
and U13759 (N_13759,N_9024,N_11784);
nor U13760 (N_13760,N_10532,N_10261);
nor U13761 (N_13761,N_9621,N_11626);
nand U13762 (N_13762,N_11893,N_10595);
and U13763 (N_13763,N_9271,N_11279);
nor U13764 (N_13764,N_10972,N_9745);
nand U13765 (N_13765,N_11141,N_9280);
or U13766 (N_13766,N_11879,N_11408);
or U13767 (N_13767,N_10732,N_11795);
or U13768 (N_13768,N_11167,N_10027);
nor U13769 (N_13769,N_9325,N_10195);
nand U13770 (N_13770,N_10513,N_10742);
xnor U13771 (N_13771,N_9253,N_10409);
or U13772 (N_13772,N_10032,N_9170);
nor U13773 (N_13773,N_9719,N_9066);
nand U13774 (N_13774,N_11628,N_9521);
nor U13775 (N_13775,N_10543,N_10491);
nand U13776 (N_13776,N_9825,N_10243);
nand U13777 (N_13777,N_9493,N_10230);
or U13778 (N_13778,N_11950,N_10648);
nor U13779 (N_13779,N_11214,N_9547);
nand U13780 (N_13780,N_10552,N_11701);
and U13781 (N_13781,N_9437,N_11149);
or U13782 (N_13782,N_10351,N_10235);
nand U13783 (N_13783,N_11604,N_10680);
or U13784 (N_13784,N_10523,N_10353);
and U13785 (N_13785,N_10543,N_9855);
or U13786 (N_13786,N_9951,N_9521);
and U13787 (N_13787,N_9448,N_9997);
and U13788 (N_13788,N_11085,N_9373);
and U13789 (N_13789,N_9533,N_11242);
and U13790 (N_13790,N_11962,N_9207);
and U13791 (N_13791,N_10064,N_11037);
xor U13792 (N_13792,N_10510,N_9249);
nand U13793 (N_13793,N_10070,N_10425);
nand U13794 (N_13794,N_9012,N_9988);
or U13795 (N_13795,N_11484,N_10863);
nand U13796 (N_13796,N_10469,N_10860);
and U13797 (N_13797,N_10388,N_9607);
and U13798 (N_13798,N_9609,N_10372);
and U13799 (N_13799,N_9748,N_10791);
nor U13800 (N_13800,N_10500,N_10879);
or U13801 (N_13801,N_11016,N_10127);
nor U13802 (N_13802,N_11398,N_10519);
nor U13803 (N_13803,N_11269,N_10626);
nor U13804 (N_13804,N_9915,N_10646);
nand U13805 (N_13805,N_11479,N_10400);
or U13806 (N_13806,N_11333,N_10900);
nand U13807 (N_13807,N_10850,N_11751);
nor U13808 (N_13808,N_10343,N_11440);
nand U13809 (N_13809,N_9962,N_11942);
or U13810 (N_13810,N_9603,N_11565);
and U13811 (N_13811,N_10442,N_10223);
and U13812 (N_13812,N_9101,N_11673);
or U13813 (N_13813,N_11730,N_9107);
or U13814 (N_13814,N_9623,N_11476);
xnor U13815 (N_13815,N_9272,N_10876);
xnor U13816 (N_13816,N_9229,N_10646);
or U13817 (N_13817,N_10130,N_11425);
xor U13818 (N_13818,N_9080,N_11586);
xor U13819 (N_13819,N_10559,N_9804);
or U13820 (N_13820,N_11488,N_9109);
or U13821 (N_13821,N_10377,N_11999);
and U13822 (N_13822,N_11165,N_11205);
and U13823 (N_13823,N_11357,N_10133);
xor U13824 (N_13824,N_9390,N_10851);
nor U13825 (N_13825,N_11020,N_10574);
or U13826 (N_13826,N_10378,N_11502);
nand U13827 (N_13827,N_10021,N_9201);
or U13828 (N_13828,N_11454,N_9602);
nor U13829 (N_13829,N_11020,N_11493);
xnor U13830 (N_13830,N_9791,N_10601);
nand U13831 (N_13831,N_9658,N_11280);
xor U13832 (N_13832,N_9325,N_11153);
or U13833 (N_13833,N_10972,N_11489);
nand U13834 (N_13834,N_10243,N_11924);
or U13835 (N_13835,N_10718,N_11136);
and U13836 (N_13836,N_10081,N_9148);
xor U13837 (N_13837,N_10574,N_11632);
nand U13838 (N_13838,N_9541,N_9221);
nor U13839 (N_13839,N_10375,N_11421);
nand U13840 (N_13840,N_9627,N_11450);
nor U13841 (N_13841,N_10585,N_10951);
and U13842 (N_13842,N_10852,N_11456);
nor U13843 (N_13843,N_9536,N_9978);
nor U13844 (N_13844,N_10182,N_10055);
and U13845 (N_13845,N_10610,N_11384);
nor U13846 (N_13846,N_10567,N_11074);
or U13847 (N_13847,N_9941,N_11676);
or U13848 (N_13848,N_10502,N_9033);
or U13849 (N_13849,N_11604,N_9944);
and U13850 (N_13850,N_11331,N_10738);
xnor U13851 (N_13851,N_9342,N_10974);
or U13852 (N_13852,N_11165,N_10263);
or U13853 (N_13853,N_9398,N_11026);
xor U13854 (N_13854,N_9447,N_11582);
and U13855 (N_13855,N_11003,N_10196);
or U13856 (N_13856,N_10869,N_10086);
xnor U13857 (N_13857,N_9784,N_11558);
and U13858 (N_13858,N_9276,N_11804);
and U13859 (N_13859,N_11785,N_10619);
and U13860 (N_13860,N_11536,N_11460);
or U13861 (N_13861,N_10530,N_9271);
xor U13862 (N_13862,N_11182,N_11278);
nor U13863 (N_13863,N_10261,N_9526);
or U13864 (N_13864,N_11156,N_10300);
nor U13865 (N_13865,N_9485,N_11977);
and U13866 (N_13866,N_9580,N_10257);
nor U13867 (N_13867,N_9538,N_11008);
nor U13868 (N_13868,N_9892,N_9032);
or U13869 (N_13869,N_11278,N_9489);
nand U13870 (N_13870,N_9828,N_11634);
xor U13871 (N_13871,N_10519,N_9875);
and U13872 (N_13872,N_10104,N_9774);
and U13873 (N_13873,N_11756,N_10188);
nor U13874 (N_13874,N_9957,N_11685);
and U13875 (N_13875,N_9604,N_9943);
nor U13876 (N_13876,N_10459,N_9760);
or U13877 (N_13877,N_10465,N_10908);
nand U13878 (N_13878,N_10572,N_9797);
and U13879 (N_13879,N_10948,N_10774);
or U13880 (N_13880,N_11937,N_9283);
and U13881 (N_13881,N_11373,N_9607);
and U13882 (N_13882,N_10928,N_10531);
nand U13883 (N_13883,N_9248,N_11669);
nor U13884 (N_13884,N_9662,N_10662);
or U13885 (N_13885,N_11104,N_10683);
or U13886 (N_13886,N_10762,N_10172);
nor U13887 (N_13887,N_9268,N_11508);
xnor U13888 (N_13888,N_10042,N_11558);
nand U13889 (N_13889,N_9433,N_11565);
or U13890 (N_13890,N_10049,N_9595);
or U13891 (N_13891,N_11387,N_11481);
nor U13892 (N_13892,N_10904,N_10321);
or U13893 (N_13893,N_10240,N_9841);
xor U13894 (N_13894,N_11197,N_10206);
and U13895 (N_13895,N_10023,N_9505);
and U13896 (N_13896,N_11515,N_9028);
and U13897 (N_13897,N_11744,N_9607);
nand U13898 (N_13898,N_11019,N_11984);
nor U13899 (N_13899,N_11658,N_11387);
and U13900 (N_13900,N_10201,N_9343);
nor U13901 (N_13901,N_11030,N_11985);
nand U13902 (N_13902,N_9423,N_11704);
or U13903 (N_13903,N_11133,N_11129);
nor U13904 (N_13904,N_10781,N_11571);
and U13905 (N_13905,N_11523,N_9948);
nand U13906 (N_13906,N_11417,N_9794);
nand U13907 (N_13907,N_11163,N_10770);
xnor U13908 (N_13908,N_10113,N_10041);
xnor U13909 (N_13909,N_10297,N_10895);
and U13910 (N_13910,N_11559,N_10166);
nor U13911 (N_13911,N_9057,N_9734);
nor U13912 (N_13912,N_9361,N_9133);
or U13913 (N_13913,N_9837,N_9389);
nand U13914 (N_13914,N_9694,N_11618);
or U13915 (N_13915,N_10916,N_9109);
and U13916 (N_13916,N_9567,N_9076);
nand U13917 (N_13917,N_9560,N_9522);
and U13918 (N_13918,N_11919,N_11097);
xor U13919 (N_13919,N_11609,N_10664);
nand U13920 (N_13920,N_10410,N_11940);
nor U13921 (N_13921,N_10175,N_11727);
xnor U13922 (N_13922,N_10234,N_11595);
and U13923 (N_13923,N_9096,N_10476);
nor U13924 (N_13924,N_9568,N_11907);
or U13925 (N_13925,N_9988,N_9499);
nor U13926 (N_13926,N_9198,N_10381);
xnor U13927 (N_13927,N_10752,N_11294);
nor U13928 (N_13928,N_10698,N_11319);
nand U13929 (N_13929,N_10504,N_11679);
and U13930 (N_13930,N_11606,N_11347);
and U13931 (N_13931,N_10532,N_11449);
and U13932 (N_13932,N_11020,N_9842);
and U13933 (N_13933,N_10859,N_9821);
or U13934 (N_13934,N_11543,N_11158);
nand U13935 (N_13935,N_10936,N_9026);
xnor U13936 (N_13936,N_9193,N_11517);
nand U13937 (N_13937,N_9426,N_10830);
xnor U13938 (N_13938,N_10389,N_11204);
and U13939 (N_13939,N_9201,N_10022);
nand U13940 (N_13940,N_9422,N_10378);
and U13941 (N_13941,N_11775,N_9708);
and U13942 (N_13942,N_11623,N_10885);
nor U13943 (N_13943,N_11541,N_10069);
nor U13944 (N_13944,N_10297,N_10721);
nor U13945 (N_13945,N_9310,N_11088);
xor U13946 (N_13946,N_10846,N_10959);
xor U13947 (N_13947,N_9022,N_11631);
and U13948 (N_13948,N_11135,N_11541);
xnor U13949 (N_13949,N_11461,N_9399);
or U13950 (N_13950,N_10590,N_11594);
nand U13951 (N_13951,N_11094,N_10781);
xor U13952 (N_13952,N_11631,N_9646);
nand U13953 (N_13953,N_10546,N_11998);
or U13954 (N_13954,N_11422,N_11714);
nand U13955 (N_13955,N_9719,N_11302);
or U13956 (N_13956,N_9344,N_9275);
and U13957 (N_13957,N_10863,N_11734);
nand U13958 (N_13958,N_9817,N_10929);
nor U13959 (N_13959,N_9254,N_11024);
nand U13960 (N_13960,N_10015,N_11308);
nand U13961 (N_13961,N_11672,N_9058);
nand U13962 (N_13962,N_9754,N_9359);
and U13963 (N_13963,N_10869,N_9877);
xor U13964 (N_13964,N_10910,N_11660);
and U13965 (N_13965,N_10520,N_10111);
or U13966 (N_13966,N_11599,N_9938);
and U13967 (N_13967,N_10868,N_9708);
or U13968 (N_13968,N_10537,N_10601);
nor U13969 (N_13969,N_9020,N_11085);
nor U13970 (N_13970,N_11896,N_9338);
nand U13971 (N_13971,N_11456,N_11266);
xnor U13972 (N_13972,N_10761,N_10245);
or U13973 (N_13973,N_11118,N_9481);
nand U13974 (N_13974,N_9756,N_11533);
nor U13975 (N_13975,N_11170,N_11106);
or U13976 (N_13976,N_9469,N_10570);
nand U13977 (N_13977,N_9315,N_11257);
and U13978 (N_13978,N_10173,N_11945);
nand U13979 (N_13979,N_10723,N_9597);
or U13980 (N_13980,N_9498,N_11618);
nand U13981 (N_13981,N_11299,N_10458);
and U13982 (N_13982,N_10010,N_11293);
nand U13983 (N_13983,N_9717,N_11387);
or U13984 (N_13984,N_10975,N_9029);
or U13985 (N_13985,N_10672,N_9266);
nand U13986 (N_13986,N_11057,N_11779);
or U13987 (N_13987,N_10392,N_10287);
and U13988 (N_13988,N_10624,N_10211);
xor U13989 (N_13989,N_10372,N_9430);
and U13990 (N_13990,N_10029,N_9626);
xnor U13991 (N_13991,N_10831,N_9791);
or U13992 (N_13992,N_10912,N_9771);
and U13993 (N_13993,N_11065,N_9365);
nand U13994 (N_13994,N_11945,N_9933);
nand U13995 (N_13995,N_11931,N_10762);
nor U13996 (N_13996,N_11790,N_9271);
or U13997 (N_13997,N_9241,N_10121);
xnor U13998 (N_13998,N_9925,N_11443);
nand U13999 (N_13999,N_10572,N_9650);
and U14000 (N_14000,N_9075,N_9363);
nor U14001 (N_14001,N_9650,N_9096);
nand U14002 (N_14002,N_11488,N_9776);
nor U14003 (N_14003,N_9961,N_9526);
or U14004 (N_14004,N_11699,N_9322);
nor U14005 (N_14005,N_10904,N_10521);
nor U14006 (N_14006,N_9597,N_9949);
nor U14007 (N_14007,N_10012,N_10676);
nand U14008 (N_14008,N_9054,N_11887);
nand U14009 (N_14009,N_9029,N_11339);
xor U14010 (N_14010,N_9510,N_10698);
nand U14011 (N_14011,N_9949,N_11932);
nor U14012 (N_14012,N_9727,N_11369);
nand U14013 (N_14013,N_9363,N_10015);
or U14014 (N_14014,N_9195,N_11383);
and U14015 (N_14015,N_9440,N_9558);
xnor U14016 (N_14016,N_10547,N_9120);
and U14017 (N_14017,N_11141,N_9692);
and U14018 (N_14018,N_10838,N_11532);
nor U14019 (N_14019,N_9993,N_9367);
nor U14020 (N_14020,N_11774,N_9022);
and U14021 (N_14021,N_10480,N_11816);
or U14022 (N_14022,N_9095,N_11976);
or U14023 (N_14023,N_9720,N_10706);
nand U14024 (N_14024,N_11408,N_11947);
and U14025 (N_14025,N_10539,N_10559);
and U14026 (N_14026,N_10361,N_9955);
and U14027 (N_14027,N_10868,N_11471);
nor U14028 (N_14028,N_10180,N_10537);
and U14029 (N_14029,N_9756,N_9033);
and U14030 (N_14030,N_9144,N_11707);
xor U14031 (N_14031,N_9243,N_11368);
xor U14032 (N_14032,N_10847,N_11002);
xor U14033 (N_14033,N_10959,N_11315);
nor U14034 (N_14034,N_9207,N_10978);
and U14035 (N_14035,N_10611,N_11230);
nor U14036 (N_14036,N_11768,N_10386);
or U14037 (N_14037,N_9869,N_10481);
or U14038 (N_14038,N_10636,N_10573);
nor U14039 (N_14039,N_9038,N_9307);
nor U14040 (N_14040,N_10287,N_11665);
nand U14041 (N_14041,N_9892,N_10251);
nand U14042 (N_14042,N_10157,N_10630);
nor U14043 (N_14043,N_10397,N_11945);
nor U14044 (N_14044,N_9279,N_11578);
xor U14045 (N_14045,N_9486,N_11881);
or U14046 (N_14046,N_11226,N_11294);
and U14047 (N_14047,N_9764,N_9701);
nand U14048 (N_14048,N_9968,N_10594);
and U14049 (N_14049,N_10261,N_11413);
xnor U14050 (N_14050,N_11799,N_10139);
or U14051 (N_14051,N_9325,N_11503);
or U14052 (N_14052,N_11041,N_9176);
nor U14053 (N_14053,N_10468,N_11799);
or U14054 (N_14054,N_9700,N_11623);
or U14055 (N_14055,N_11144,N_10082);
and U14056 (N_14056,N_9914,N_10969);
nand U14057 (N_14057,N_11829,N_11744);
or U14058 (N_14058,N_11991,N_11771);
or U14059 (N_14059,N_10386,N_9652);
or U14060 (N_14060,N_10760,N_9679);
and U14061 (N_14061,N_9013,N_11303);
nor U14062 (N_14062,N_9380,N_11924);
nand U14063 (N_14063,N_9455,N_11804);
nor U14064 (N_14064,N_11669,N_10676);
xnor U14065 (N_14065,N_9745,N_9202);
and U14066 (N_14066,N_9937,N_11099);
nand U14067 (N_14067,N_10481,N_10872);
nor U14068 (N_14068,N_10667,N_9117);
and U14069 (N_14069,N_10812,N_11328);
xnor U14070 (N_14070,N_10072,N_11730);
or U14071 (N_14071,N_10355,N_9326);
or U14072 (N_14072,N_9396,N_11665);
and U14073 (N_14073,N_9360,N_10627);
or U14074 (N_14074,N_10016,N_11438);
or U14075 (N_14075,N_10965,N_11235);
or U14076 (N_14076,N_9267,N_10593);
nand U14077 (N_14077,N_10411,N_10194);
or U14078 (N_14078,N_11684,N_10645);
nand U14079 (N_14079,N_10262,N_11960);
and U14080 (N_14080,N_11315,N_10053);
nand U14081 (N_14081,N_11206,N_9750);
nand U14082 (N_14082,N_10280,N_10857);
nor U14083 (N_14083,N_11137,N_10413);
or U14084 (N_14084,N_11851,N_9865);
or U14085 (N_14085,N_10853,N_10324);
and U14086 (N_14086,N_11965,N_10247);
or U14087 (N_14087,N_10684,N_11885);
nand U14088 (N_14088,N_9288,N_9025);
nor U14089 (N_14089,N_9797,N_9327);
and U14090 (N_14090,N_11543,N_10021);
nor U14091 (N_14091,N_11569,N_9514);
nor U14092 (N_14092,N_11971,N_9492);
nor U14093 (N_14093,N_9535,N_11146);
or U14094 (N_14094,N_9029,N_10846);
or U14095 (N_14095,N_10529,N_10309);
nand U14096 (N_14096,N_11061,N_10982);
or U14097 (N_14097,N_9841,N_10235);
nor U14098 (N_14098,N_10772,N_10999);
nor U14099 (N_14099,N_11979,N_10257);
and U14100 (N_14100,N_9351,N_11646);
nand U14101 (N_14101,N_11265,N_9053);
or U14102 (N_14102,N_10279,N_9660);
or U14103 (N_14103,N_10325,N_11652);
or U14104 (N_14104,N_11689,N_10074);
xor U14105 (N_14105,N_11203,N_11213);
nand U14106 (N_14106,N_9450,N_11042);
or U14107 (N_14107,N_9778,N_9935);
nand U14108 (N_14108,N_9604,N_9428);
nor U14109 (N_14109,N_11089,N_10577);
or U14110 (N_14110,N_9478,N_11596);
nor U14111 (N_14111,N_10139,N_11471);
or U14112 (N_14112,N_11035,N_10834);
nand U14113 (N_14113,N_10595,N_11376);
and U14114 (N_14114,N_10631,N_10127);
or U14115 (N_14115,N_9630,N_10441);
or U14116 (N_14116,N_9365,N_11361);
nor U14117 (N_14117,N_10902,N_9975);
or U14118 (N_14118,N_9531,N_11239);
xnor U14119 (N_14119,N_9014,N_11666);
nand U14120 (N_14120,N_9233,N_11845);
nand U14121 (N_14121,N_11570,N_10629);
or U14122 (N_14122,N_11165,N_11325);
nor U14123 (N_14123,N_10932,N_11660);
or U14124 (N_14124,N_11664,N_11126);
nor U14125 (N_14125,N_9478,N_10431);
and U14126 (N_14126,N_10109,N_10266);
and U14127 (N_14127,N_11821,N_11442);
and U14128 (N_14128,N_10737,N_10645);
nand U14129 (N_14129,N_10044,N_11323);
nand U14130 (N_14130,N_9041,N_9215);
nor U14131 (N_14131,N_11172,N_11176);
nor U14132 (N_14132,N_11670,N_11723);
and U14133 (N_14133,N_10817,N_9149);
or U14134 (N_14134,N_11902,N_11037);
nand U14135 (N_14135,N_9479,N_9734);
xnor U14136 (N_14136,N_9373,N_10421);
xor U14137 (N_14137,N_10333,N_9165);
or U14138 (N_14138,N_9677,N_11957);
nand U14139 (N_14139,N_9952,N_9714);
nand U14140 (N_14140,N_11413,N_9957);
and U14141 (N_14141,N_9925,N_9502);
or U14142 (N_14142,N_11747,N_11313);
nand U14143 (N_14143,N_9589,N_11317);
nand U14144 (N_14144,N_9019,N_10745);
nand U14145 (N_14145,N_11829,N_11224);
nor U14146 (N_14146,N_11585,N_10391);
and U14147 (N_14147,N_10413,N_11155);
and U14148 (N_14148,N_10630,N_11803);
nand U14149 (N_14149,N_9145,N_11971);
or U14150 (N_14150,N_10145,N_10104);
nor U14151 (N_14151,N_11553,N_9226);
and U14152 (N_14152,N_10854,N_10201);
or U14153 (N_14153,N_10126,N_9548);
and U14154 (N_14154,N_11612,N_11402);
nor U14155 (N_14155,N_9130,N_9016);
and U14156 (N_14156,N_11376,N_11040);
nor U14157 (N_14157,N_10062,N_9991);
or U14158 (N_14158,N_9544,N_11822);
nand U14159 (N_14159,N_9465,N_9610);
and U14160 (N_14160,N_10297,N_9781);
and U14161 (N_14161,N_9038,N_10160);
nand U14162 (N_14162,N_10878,N_10928);
nor U14163 (N_14163,N_11324,N_9313);
and U14164 (N_14164,N_10172,N_9316);
xor U14165 (N_14165,N_11201,N_9602);
nor U14166 (N_14166,N_9088,N_9647);
and U14167 (N_14167,N_9477,N_9481);
and U14168 (N_14168,N_11167,N_11320);
nor U14169 (N_14169,N_9333,N_10837);
or U14170 (N_14170,N_9563,N_10428);
nor U14171 (N_14171,N_9363,N_11401);
nor U14172 (N_14172,N_9395,N_11969);
nor U14173 (N_14173,N_11024,N_10609);
and U14174 (N_14174,N_10998,N_9847);
nor U14175 (N_14175,N_9284,N_9031);
and U14176 (N_14176,N_11172,N_10069);
nand U14177 (N_14177,N_10793,N_11846);
and U14178 (N_14178,N_9810,N_10900);
nor U14179 (N_14179,N_10390,N_9324);
or U14180 (N_14180,N_9804,N_11019);
nor U14181 (N_14181,N_9619,N_11797);
and U14182 (N_14182,N_11674,N_10733);
nor U14183 (N_14183,N_11113,N_11449);
nand U14184 (N_14184,N_10681,N_11009);
nor U14185 (N_14185,N_9291,N_11047);
nand U14186 (N_14186,N_10899,N_10973);
and U14187 (N_14187,N_10522,N_9484);
or U14188 (N_14188,N_10628,N_9518);
or U14189 (N_14189,N_11197,N_10089);
nand U14190 (N_14190,N_9719,N_10859);
and U14191 (N_14191,N_9794,N_9624);
nor U14192 (N_14192,N_10592,N_11744);
nand U14193 (N_14193,N_11234,N_9537);
nand U14194 (N_14194,N_9082,N_11812);
nand U14195 (N_14195,N_11940,N_11058);
and U14196 (N_14196,N_11692,N_10543);
nand U14197 (N_14197,N_9377,N_9374);
nor U14198 (N_14198,N_9790,N_9991);
or U14199 (N_14199,N_9786,N_10417);
and U14200 (N_14200,N_10821,N_10419);
or U14201 (N_14201,N_9102,N_10178);
and U14202 (N_14202,N_11309,N_10739);
nand U14203 (N_14203,N_10373,N_10543);
nor U14204 (N_14204,N_11440,N_9750);
nor U14205 (N_14205,N_11805,N_9198);
and U14206 (N_14206,N_9416,N_9030);
xor U14207 (N_14207,N_10893,N_10043);
or U14208 (N_14208,N_11217,N_11570);
and U14209 (N_14209,N_10149,N_11426);
or U14210 (N_14210,N_9831,N_9630);
nor U14211 (N_14211,N_10347,N_11098);
or U14212 (N_14212,N_9022,N_11498);
nor U14213 (N_14213,N_11363,N_10402);
or U14214 (N_14214,N_10534,N_11202);
xor U14215 (N_14215,N_11587,N_10757);
nand U14216 (N_14216,N_9606,N_9999);
and U14217 (N_14217,N_11877,N_9121);
nand U14218 (N_14218,N_10386,N_9284);
nand U14219 (N_14219,N_11934,N_9643);
and U14220 (N_14220,N_11500,N_10433);
nor U14221 (N_14221,N_9988,N_10676);
nand U14222 (N_14222,N_10895,N_11199);
xor U14223 (N_14223,N_11873,N_11946);
and U14224 (N_14224,N_11169,N_10442);
nor U14225 (N_14225,N_11917,N_11890);
and U14226 (N_14226,N_11630,N_10980);
or U14227 (N_14227,N_11606,N_9084);
or U14228 (N_14228,N_10100,N_10645);
and U14229 (N_14229,N_10320,N_11376);
and U14230 (N_14230,N_11697,N_9531);
nand U14231 (N_14231,N_11956,N_11021);
xnor U14232 (N_14232,N_11865,N_9671);
and U14233 (N_14233,N_11887,N_9104);
nand U14234 (N_14234,N_10334,N_11767);
xor U14235 (N_14235,N_9037,N_11866);
or U14236 (N_14236,N_9789,N_11607);
xnor U14237 (N_14237,N_10303,N_11303);
and U14238 (N_14238,N_10208,N_10065);
nor U14239 (N_14239,N_10691,N_9006);
xnor U14240 (N_14240,N_9567,N_9033);
and U14241 (N_14241,N_9225,N_11989);
nand U14242 (N_14242,N_9928,N_11150);
xor U14243 (N_14243,N_10110,N_11927);
xor U14244 (N_14244,N_11038,N_10207);
nand U14245 (N_14245,N_10807,N_11602);
xnor U14246 (N_14246,N_11000,N_9594);
and U14247 (N_14247,N_11685,N_11311);
xnor U14248 (N_14248,N_11793,N_9308);
or U14249 (N_14249,N_9629,N_9490);
nor U14250 (N_14250,N_10354,N_9152);
or U14251 (N_14251,N_11355,N_10897);
and U14252 (N_14252,N_9127,N_11194);
nand U14253 (N_14253,N_9849,N_9532);
nand U14254 (N_14254,N_9488,N_9861);
or U14255 (N_14255,N_10680,N_11590);
nand U14256 (N_14256,N_9029,N_9641);
or U14257 (N_14257,N_9086,N_11615);
xor U14258 (N_14258,N_9560,N_9312);
xor U14259 (N_14259,N_10220,N_9372);
or U14260 (N_14260,N_9286,N_11337);
or U14261 (N_14261,N_11295,N_10484);
nor U14262 (N_14262,N_11732,N_10932);
and U14263 (N_14263,N_11317,N_9949);
or U14264 (N_14264,N_9571,N_9277);
nand U14265 (N_14265,N_10731,N_10871);
and U14266 (N_14266,N_9884,N_10174);
or U14267 (N_14267,N_11102,N_10961);
and U14268 (N_14268,N_10896,N_10305);
nand U14269 (N_14269,N_11694,N_10796);
nor U14270 (N_14270,N_10056,N_10895);
nand U14271 (N_14271,N_11438,N_9505);
nor U14272 (N_14272,N_9043,N_11020);
nand U14273 (N_14273,N_10211,N_9457);
nand U14274 (N_14274,N_11421,N_11222);
xnor U14275 (N_14275,N_9969,N_9238);
or U14276 (N_14276,N_11706,N_10468);
nor U14277 (N_14277,N_9730,N_10978);
nor U14278 (N_14278,N_11948,N_9878);
xor U14279 (N_14279,N_11147,N_9015);
nor U14280 (N_14280,N_9329,N_9630);
nor U14281 (N_14281,N_11640,N_9985);
nand U14282 (N_14282,N_9218,N_11440);
and U14283 (N_14283,N_10302,N_10170);
or U14284 (N_14284,N_10012,N_10252);
nor U14285 (N_14285,N_10364,N_9698);
nand U14286 (N_14286,N_10933,N_10974);
nor U14287 (N_14287,N_11623,N_9492);
nor U14288 (N_14288,N_10536,N_11097);
xnor U14289 (N_14289,N_11593,N_10175);
nand U14290 (N_14290,N_9736,N_11269);
xor U14291 (N_14291,N_11524,N_9855);
or U14292 (N_14292,N_11592,N_10653);
nand U14293 (N_14293,N_9215,N_10324);
or U14294 (N_14294,N_9204,N_9814);
nor U14295 (N_14295,N_10852,N_11373);
and U14296 (N_14296,N_9653,N_9968);
or U14297 (N_14297,N_11049,N_11292);
xnor U14298 (N_14298,N_9785,N_9879);
nor U14299 (N_14299,N_10573,N_10377);
and U14300 (N_14300,N_11446,N_9049);
nor U14301 (N_14301,N_10790,N_10884);
nor U14302 (N_14302,N_10422,N_11653);
nor U14303 (N_14303,N_9871,N_11965);
or U14304 (N_14304,N_11974,N_9133);
xnor U14305 (N_14305,N_9585,N_9892);
nand U14306 (N_14306,N_10766,N_9012);
xor U14307 (N_14307,N_9329,N_9477);
nand U14308 (N_14308,N_10513,N_9002);
xnor U14309 (N_14309,N_11384,N_10972);
xnor U14310 (N_14310,N_9448,N_10097);
or U14311 (N_14311,N_10555,N_9167);
nand U14312 (N_14312,N_10245,N_11162);
nand U14313 (N_14313,N_10798,N_10578);
or U14314 (N_14314,N_9444,N_10791);
and U14315 (N_14315,N_10773,N_10287);
and U14316 (N_14316,N_9754,N_10461);
nor U14317 (N_14317,N_9832,N_11427);
or U14318 (N_14318,N_11175,N_10789);
nand U14319 (N_14319,N_11016,N_11709);
and U14320 (N_14320,N_10187,N_10252);
or U14321 (N_14321,N_11584,N_9670);
or U14322 (N_14322,N_10845,N_10027);
xnor U14323 (N_14323,N_11964,N_9482);
nand U14324 (N_14324,N_11179,N_10286);
nor U14325 (N_14325,N_11744,N_9661);
xnor U14326 (N_14326,N_10889,N_9260);
nor U14327 (N_14327,N_11128,N_10000);
xnor U14328 (N_14328,N_9043,N_10024);
nand U14329 (N_14329,N_11862,N_9323);
and U14330 (N_14330,N_9663,N_9519);
nor U14331 (N_14331,N_10268,N_10277);
and U14332 (N_14332,N_11745,N_11552);
and U14333 (N_14333,N_9366,N_10052);
or U14334 (N_14334,N_10346,N_10967);
xnor U14335 (N_14335,N_11607,N_10769);
or U14336 (N_14336,N_11055,N_10105);
and U14337 (N_14337,N_10403,N_11081);
nor U14338 (N_14338,N_9239,N_10168);
nor U14339 (N_14339,N_10652,N_10261);
nor U14340 (N_14340,N_9069,N_9065);
nand U14341 (N_14341,N_11663,N_11236);
or U14342 (N_14342,N_11193,N_10140);
and U14343 (N_14343,N_11794,N_9050);
nor U14344 (N_14344,N_10448,N_9947);
nand U14345 (N_14345,N_9804,N_11433);
nor U14346 (N_14346,N_10826,N_11567);
or U14347 (N_14347,N_11439,N_10259);
or U14348 (N_14348,N_10319,N_11439);
or U14349 (N_14349,N_11080,N_9489);
or U14350 (N_14350,N_9516,N_9075);
or U14351 (N_14351,N_11227,N_10064);
nor U14352 (N_14352,N_11636,N_10685);
or U14353 (N_14353,N_11678,N_11556);
nand U14354 (N_14354,N_11614,N_9411);
or U14355 (N_14355,N_9938,N_9882);
nor U14356 (N_14356,N_9184,N_11244);
nor U14357 (N_14357,N_10401,N_9483);
nor U14358 (N_14358,N_11533,N_11310);
and U14359 (N_14359,N_9383,N_10478);
nand U14360 (N_14360,N_10443,N_10472);
nand U14361 (N_14361,N_9978,N_10905);
and U14362 (N_14362,N_9016,N_10825);
or U14363 (N_14363,N_9436,N_9997);
nand U14364 (N_14364,N_9862,N_10209);
and U14365 (N_14365,N_10344,N_9780);
nand U14366 (N_14366,N_9536,N_9471);
nor U14367 (N_14367,N_10906,N_9969);
nor U14368 (N_14368,N_11189,N_11960);
nor U14369 (N_14369,N_11821,N_10883);
nor U14370 (N_14370,N_11037,N_11310);
and U14371 (N_14371,N_10110,N_10462);
nand U14372 (N_14372,N_10256,N_10243);
nand U14373 (N_14373,N_11143,N_11761);
nand U14374 (N_14374,N_9636,N_11256);
nand U14375 (N_14375,N_11213,N_9042);
xnor U14376 (N_14376,N_10869,N_11107);
nand U14377 (N_14377,N_11566,N_9354);
or U14378 (N_14378,N_9348,N_11680);
or U14379 (N_14379,N_9435,N_9881);
and U14380 (N_14380,N_11991,N_10000);
nor U14381 (N_14381,N_9533,N_10227);
xnor U14382 (N_14382,N_10802,N_11391);
nor U14383 (N_14383,N_11783,N_9233);
and U14384 (N_14384,N_11962,N_10818);
and U14385 (N_14385,N_10539,N_11918);
nand U14386 (N_14386,N_10067,N_9513);
nor U14387 (N_14387,N_9347,N_10296);
or U14388 (N_14388,N_11109,N_10271);
and U14389 (N_14389,N_11168,N_9493);
xnor U14390 (N_14390,N_9945,N_9200);
and U14391 (N_14391,N_9392,N_10928);
nor U14392 (N_14392,N_9310,N_10979);
and U14393 (N_14393,N_9129,N_9908);
nand U14394 (N_14394,N_10382,N_10182);
or U14395 (N_14395,N_11660,N_10287);
nor U14396 (N_14396,N_11586,N_11391);
xnor U14397 (N_14397,N_9043,N_11455);
xnor U14398 (N_14398,N_9354,N_9998);
nand U14399 (N_14399,N_10822,N_10270);
or U14400 (N_14400,N_10617,N_11864);
xnor U14401 (N_14401,N_9608,N_9280);
and U14402 (N_14402,N_11782,N_11209);
nor U14403 (N_14403,N_10571,N_9888);
and U14404 (N_14404,N_10475,N_10973);
xnor U14405 (N_14405,N_11893,N_9407);
or U14406 (N_14406,N_11143,N_11489);
nand U14407 (N_14407,N_11280,N_9185);
xor U14408 (N_14408,N_9189,N_11591);
nor U14409 (N_14409,N_10240,N_9861);
or U14410 (N_14410,N_11277,N_10179);
or U14411 (N_14411,N_10721,N_11651);
and U14412 (N_14412,N_9095,N_11273);
or U14413 (N_14413,N_9327,N_9718);
or U14414 (N_14414,N_9595,N_9224);
and U14415 (N_14415,N_11239,N_11067);
and U14416 (N_14416,N_9804,N_9297);
or U14417 (N_14417,N_11261,N_11282);
and U14418 (N_14418,N_9244,N_9843);
or U14419 (N_14419,N_9434,N_10898);
nor U14420 (N_14420,N_11330,N_9862);
nor U14421 (N_14421,N_11980,N_9873);
nand U14422 (N_14422,N_9222,N_11980);
or U14423 (N_14423,N_9099,N_9363);
or U14424 (N_14424,N_11470,N_9823);
or U14425 (N_14425,N_10536,N_9328);
nand U14426 (N_14426,N_9121,N_9510);
and U14427 (N_14427,N_9332,N_11421);
nor U14428 (N_14428,N_9161,N_11535);
nor U14429 (N_14429,N_9532,N_11727);
or U14430 (N_14430,N_9542,N_9533);
and U14431 (N_14431,N_11486,N_11176);
nor U14432 (N_14432,N_11252,N_9058);
or U14433 (N_14433,N_9889,N_10637);
nand U14434 (N_14434,N_9594,N_9791);
nor U14435 (N_14435,N_9900,N_9176);
and U14436 (N_14436,N_11637,N_9189);
xnor U14437 (N_14437,N_9943,N_10011);
nand U14438 (N_14438,N_10457,N_10042);
and U14439 (N_14439,N_9975,N_10162);
xnor U14440 (N_14440,N_9575,N_11725);
nand U14441 (N_14441,N_10630,N_11988);
or U14442 (N_14442,N_11144,N_9618);
and U14443 (N_14443,N_10282,N_11282);
nand U14444 (N_14444,N_9052,N_9560);
or U14445 (N_14445,N_10872,N_9142);
or U14446 (N_14446,N_11497,N_10426);
nand U14447 (N_14447,N_10147,N_11583);
nor U14448 (N_14448,N_9734,N_9175);
and U14449 (N_14449,N_11890,N_10416);
xor U14450 (N_14450,N_9858,N_11976);
nor U14451 (N_14451,N_10568,N_11213);
nor U14452 (N_14452,N_10212,N_9622);
or U14453 (N_14453,N_10816,N_9451);
nor U14454 (N_14454,N_9249,N_11761);
nor U14455 (N_14455,N_10446,N_9875);
and U14456 (N_14456,N_10721,N_11528);
nand U14457 (N_14457,N_11573,N_11092);
xor U14458 (N_14458,N_10191,N_9792);
and U14459 (N_14459,N_9874,N_9578);
and U14460 (N_14460,N_9203,N_11246);
xnor U14461 (N_14461,N_11543,N_9525);
and U14462 (N_14462,N_10660,N_9502);
xnor U14463 (N_14463,N_11443,N_11435);
and U14464 (N_14464,N_10220,N_9189);
or U14465 (N_14465,N_9979,N_11055);
and U14466 (N_14466,N_10008,N_10441);
nor U14467 (N_14467,N_10508,N_11174);
nor U14468 (N_14468,N_10891,N_11723);
or U14469 (N_14469,N_10768,N_11430);
and U14470 (N_14470,N_11457,N_10503);
nand U14471 (N_14471,N_11447,N_9312);
and U14472 (N_14472,N_11041,N_11481);
nor U14473 (N_14473,N_11441,N_9992);
nand U14474 (N_14474,N_10493,N_9124);
and U14475 (N_14475,N_11107,N_9702);
nand U14476 (N_14476,N_10779,N_10365);
nand U14477 (N_14477,N_11821,N_11065);
nor U14478 (N_14478,N_10673,N_10912);
and U14479 (N_14479,N_9178,N_9078);
and U14480 (N_14480,N_9719,N_9772);
nand U14481 (N_14481,N_9946,N_10377);
xor U14482 (N_14482,N_9812,N_9070);
and U14483 (N_14483,N_9852,N_9350);
or U14484 (N_14484,N_11383,N_10730);
or U14485 (N_14485,N_10656,N_9004);
nand U14486 (N_14486,N_11583,N_11197);
or U14487 (N_14487,N_11779,N_9763);
and U14488 (N_14488,N_9517,N_9238);
nand U14489 (N_14489,N_9620,N_11956);
nand U14490 (N_14490,N_10269,N_11718);
nor U14491 (N_14491,N_9605,N_10841);
nor U14492 (N_14492,N_10803,N_10830);
or U14493 (N_14493,N_9387,N_11774);
nor U14494 (N_14494,N_11201,N_11786);
nand U14495 (N_14495,N_9179,N_9129);
nor U14496 (N_14496,N_10953,N_11819);
nor U14497 (N_14497,N_11513,N_10509);
nor U14498 (N_14498,N_9685,N_10043);
and U14499 (N_14499,N_9577,N_9748);
or U14500 (N_14500,N_10000,N_9326);
and U14501 (N_14501,N_10429,N_11476);
nor U14502 (N_14502,N_11243,N_11053);
or U14503 (N_14503,N_11167,N_9604);
nor U14504 (N_14504,N_11358,N_9404);
nor U14505 (N_14505,N_9947,N_10644);
nor U14506 (N_14506,N_11477,N_10683);
nand U14507 (N_14507,N_11147,N_9896);
nor U14508 (N_14508,N_9057,N_11876);
nand U14509 (N_14509,N_9195,N_9242);
and U14510 (N_14510,N_9134,N_10858);
nand U14511 (N_14511,N_11403,N_10528);
nand U14512 (N_14512,N_10259,N_10924);
xnor U14513 (N_14513,N_10304,N_9993);
or U14514 (N_14514,N_11443,N_10225);
xnor U14515 (N_14515,N_11955,N_10386);
and U14516 (N_14516,N_11931,N_10180);
nand U14517 (N_14517,N_10700,N_9148);
xnor U14518 (N_14518,N_11172,N_11447);
nand U14519 (N_14519,N_11125,N_10259);
or U14520 (N_14520,N_11068,N_11849);
and U14521 (N_14521,N_9503,N_9236);
or U14522 (N_14522,N_10818,N_10072);
nor U14523 (N_14523,N_9228,N_11535);
nor U14524 (N_14524,N_10950,N_9702);
nor U14525 (N_14525,N_11280,N_10906);
nor U14526 (N_14526,N_9458,N_11657);
nand U14527 (N_14527,N_11727,N_10421);
and U14528 (N_14528,N_10919,N_9968);
nand U14529 (N_14529,N_9693,N_9213);
xnor U14530 (N_14530,N_10608,N_11219);
and U14531 (N_14531,N_10726,N_10669);
nand U14532 (N_14532,N_11970,N_10116);
nand U14533 (N_14533,N_10569,N_9109);
nor U14534 (N_14534,N_10706,N_9508);
and U14535 (N_14535,N_11544,N_9965);
or U14536 (N_14536,N_10422,N_10287);
and U14537 (N_14537,N_11387,N_10588);
nand U14538 (N_14538,N_10987,N_10415);
nand U14539 (N_14539,N_11478,N_9748);
nor U14540 (N_14540,N_10075,N_11281);
nand U14541 (N_14541,N_9079,N_9397);
and U14542 (N_14542,N_11878,N_9906);
and U14543 (N_14543,N_11596,N_11965);
nor U14544 (N_14544,N_9297,N_11658);
or U14545 (N_14545,N_11451,N_10928);
and U14546 (N_14546,N_11587,N_9309);
nor U14547 (N_14547,N_9771,N_10726);
nand U14548 (N_14548,N_10403,N_9637);
nand U14549 (N_14549,N_10446,N_10340);
and U14550 (N_14550,N_9539,N_9242);
and U14551 (N_14551,N_11362,N_9488);
nand U14552 (N_14552,N_11732,N_10037);
or U14553 (N_14553,N_9613,N_9340);
and U14554 (N_14554,N_10492,N_11748);
nand U14555 (N_14555,N_11266,N_11509);
or U14556 (N_14556,N_11104,N_9636);
nand U14557 (N_14557,N_10167,N_10434);
and U14558 (N_14558,N_11148,N_10096);
and U14559 (N_14559,N_11912,N_9450);
or U14560 (N_14560,N_9261,N_11965);
nand U14561 (N_14561,N_9808,N_9693);
nand U14562 (N_14562,N_11965,N_10903);
nor U14563 (N_14563,N_9006,N_10650);
nor U14564 (N_14564,N_9677,N_9129);
or U14565 (N_14565,N_10527,N_11525);
nor U14566 (N_14566,N_11110,N_9328);
nand U14567 (N_14567,N_9351,N_10671);
nand U14568 (N_14568,N_10088,N_9793);
nand U14569 (N_14569,N_11014,N_10966);
nor U14570 (N_14570,N_10968,N_10032);
and U14571 (N_14571,N_9746,N_9293);
or U14572 (N_14572,N_11519,N_11054);
nand U14573 (N_14573,N_11631,N_10786);
nand U14574 (N_14574,N_11767,N_11093);
nor U14575 (N_14575,N_9335,N_11786);
or U14576 (N_14576,N_10208,N_11706);
nand U14577 (N_14577,N_9855,N_9334);
nor U14578 (N_14578,N_11143,N_10055);
or U14579 (N_14579,N_10004,N_10149);
and U14580 (N_14580,N_11145,N_11515);
and U14581 (N_14581,N_10340,N_11785);
nor U14582 (N_14582,N_11463,N_11008);
or U14583 (N_14583,N_9605,N_11438);
and U14584 (N_14584,N_11067,N_11814);
or U14585 (N_14585,N_10384,N_9765);
nor U14586 (N_14586,N_10180,N_10869);
nor U14587 (N_14587,N_11877,N_9198);
or U14588 (N_14588,N_9181,N_9645);
nor U14589 (N_14589,N_10111,N_10390);
and U14590 (N_14590,N_10778,N_11989);
xnor U14591 (N_14591,N_11240,N_9486);
or U14592 (N_14592,N_10656,N_11056);
or U14593 (N_14593,N_9442,N_11350);
or U14594 (N_14594,N_11890,N_9871);
and U14595 (N_14595,N_11741,N_9313);
and U14596 (N_14596,N_10864,N_10967);
nor U14597 (N_14597,N_10997,N_11646);
and U14598 (N_14598,N_10511,N_10945);
nand U14599 (N_14599,N_11488,N_9338);
or U14600 (N_14600,N_9994,N_10735);
nor U14601 (N_14601,N_9875,N_11368);
or U14602 (N_14602,N_10162,N_9654);
xnor U14603 (N_14603,N_9606,N_10149);
and U14604 (N_14604,N_9742,N_11082);
nor U14605 (N_14605,N_10056,N_10886);
and U14606 (N_14606,N_9235,N_10090);
nor U14607 (N_14607,N_11131,N_10667);
nand U14608 (N_14608,N_9921,N_9524);
or U14609 (N_14609,N_10099,N_9582);
and U14610 (N_14610,N_11576,N_10880);
or U14611 (N_14611,N_10134,N_9738);
nand U14612 (N_14612,N_11348,N_9841);
or U14613 (N_14613,N_10301,N_11159);
nand U14614 (N_14614,N_10578,N_11051);
nor U14615 (N_14615,N_11094,N_11993);
nor U14616 (N_14616,N_9500,N_9382);
nand U14617 (N_14617,N_10638,N_9649);
and U14618 (N_14618,N_11129,N_9173);
or U14619 (N_14619,N_10818,N_9699);
or U14620 (N_14620,N_10991,N_9057);
nor U14621 (N_14621,N_11355,N_9596);
xnor U14622 (N_14622,N_11547,N_9851);
nor U14623 (N_14623,N_9320,N_10874);
or U14624 (N_14624,N_11199,N_10374);
nor U14625 (N_14625,N_10723,N_11613);
and U14626 (N_14626,N_9271,N_11976);
nand U14627 (N_14627,N_10591,N_11668);
nand U14628 (N_14628,N_9947,N_11819);
and U14629 (N_14629,N_9708,N_11894);
xnor U14630 (N_14630,N_10992,N_11821);
nor U14631 (N_14631,N_11107,N_11620);
and U14632 (N_14632,N_11325,N_10414);
nor U14633 (N_14633,N_10964,N_10983);
nand U14634 (N_14634,N_10185,N_11148);
nor U14635 (N_14635,N_10598,N_9196);
nor U14636 (N_14636,N_11728,N_11329);
nand U14637 (N_14637,N_10824,N_9848);
nand U14638 (N_14638,N_10244,N_10188);
nand U14639 (N_14639,N_9342,N_11846);
nor U14640 (N_14640,N_9463,N_9817);
xnor U14641 (N_14641,N_11467,N_9656);
or U14642 (N_14642,N_10918,N_10053);
nor U14643 (N_14643,N_9713,N_10435);
or U14644 (N_14644,N_11205,N_10367);
nand U14645 (N_14645,N_9064,N_11273);
nor U14646 (N_14646,N_9433,N_10310);
nor U14647 (N_14647,N_9972,N_10803);
nor U14648 (N_14648,N_11495,N_10177);
nor U14649 (N_14649,N_9196,N_11805);
or U14650 (N_14650,N_10910,N_11914);
or U14651 (N_14651,N_9927,N_11111);
nor U14652 (N_14652,N_11808,N_10999);
and U14653 (N_14653,N_11127,N_10696);
nor U14654 (N_14654,N_10142,N_10184);
and U14655 (N_14655,N_10957,N_11583);
xnor U14656 (N_14656,N_11105,N_11749);
and U14657 (N_14657,N_10262,N_11258);
nand U14658 (N_14658,N_11956,N_11043);
nor U14659 (N_14659,N_10508,N_10138);
nand U14660 (N_14660,N_11197,N_11196);
nor U14661 (N_14661,N_10215,N_10803);
nand U14662 (N_14662,N_9245,N_9794);
nor U14663 (N_14663,N_11641,N_10577);
and U14664 (N_14664,N_9836,N_9372);
or U14665 (N_14665,N_9468,N_9406);
nor U14666 (N_14666,N_9016,N_11094);
nand U14667 (N_14667,N_11588,N_11976);
or U14668 (N_14668,N_11359,N_9300);
xor U14669 (N_14669,N_10781,N_9914);
xnor U14670 (N_14670,N_10870,N_9936);
nand U14671 (N_14671,N_9413,N_11787);
nor U14672 (N_14672,N_11175,N_11863);
and U14673 (N_14673,N_10457,N_10016);
or U14674 (N_14674,N_10839,N_9560);
and U14675 (N_14675,N_9308,N_10193);
and U14676 (N_14676,N_9091,N_10086);
and U14677 (N_14677,N_9536,N_10320);
and U14678 (N_14678,N_9817,N_10051);
nand U14679 (N_14679,N_10275,N_9205);
or U14680 (N_14680,N_9201,N_11242);
and U14681 (N_14681,N_10735,N_10544);
or U14682 (N_14682,N_10861,N_11896);
and U14683 (N_14683,N_11076,N_10499);
or U14684 (N_14684,N_11398,N_9694);
nand U14685 (N_14685,N_9583,N_9271);
nor U14686 (N_14686,N_9271,N_9083);
or U14687 (N_14687,N_10965,N_10208);
and U14688 (N_14688,N_9635,N_9367);
nand U14689 (N_14689,N_11684,N_9438);
nor U14690 (N_14690,N_10758,N_10777);
nor U14691 (N_14691,N_10235,N_10933);
xor U14692 (N_14692,N_10460,N_9716);
nor U14693 (N_14693,N_9871,N_9339);
nor U14694 (N_14694,N_11714,N_11739);
and U14695 (N_14695,N_10468,N_11945);
nor U14696 (N_14696,N_11607,N_11332);
or U14697 (N_14697,N_10541,N_11433);
nor U14698 (N_14698,N_10157,N_9813);
nand U14699 (N_14699,N_11841,N_10505);
nor U14700 (N_14700,N_9581,N_10946);
or U14701 (N_14701,N_11425,N_11878);
or U14702 (N_14702,N_9740,N_11406);
and U14703 (N_14703,N_10040,N_10191);
or U14704 (N_14704,N_9448,N_9802);
or U14705 (N_14705,N_10637,N_10609);
xor U14706 (N_14706,N_11488,N_10631);
nor U14707 (N_14707,N_9986,N_11290);
nand U14708 (N_14708,N_9288,N_10486);
xor U14709 (N_14709,N_10260,N_9274);
and U14710 (N_14710,N_9902,N_11539);
and U14711 (N_14711,N_11120,N_11167);
nand U14712 (N_14712,N_9194,N_9182);
nand U14713 (N_14713,N_10335,N_11453);
nand U14714 (N_14714,N_11307,N_9831);
and U14715 (N_14715,N_11057,N_10062);
or U14716 (N_14716,N_9502,N_9522);
or U14717 (N_14717,N_10608,N_10234);
and U14718 (N_14718,N_10588,N_9461);
nor U14719 (N_14719,N_11119,N_9656);
nand U14720 (N_14720,N_10593,N_11278);
or U14721 (N_14721,N_9887,N_10449);
nor U14722 (N_14722,N_10900,N_10048);
or U14723 (N_14723,N_10526,N_10741);
nand U14724 (N_14724,N_9603,N_9414);
or U14725 (N_14725,N_10943,N_11352);
nor U14726 (N_14726,N_11114,N_10262);
or U14727 (N_14727,N_10092,N_11144);
and U14728 (N_14728,N_10933,N_10059);
and U14729 (N_14729,N_11630,N_9367);
and U14730 (N_14730,N_11878,N_9775);
xor U14731 (N_14731,N_11634,N_10553);
or U14732 (N_14732,N_11002,N_11457);
xnor U14733 (N_14733,N_9832,N_10457);
or U14734 (N_14734,N_9532,N_10516);
xnor U14735 (N_14735,N_9001,N_10969);
nand U14736 (N_14736,N_10657,N_9122);
nand U14737 (N_14737,N_10315,N_11191);
xor U14738 (N_14738,N_10360,N_10784);
and U14739 (N_14739,N_9469,N_10405);
nand U14740 (N_14740,N_9838,N_10336);
or U14741 (N_14741,N_11726,N_9632);
nor U14742 (N_14742,N_9168,N_11335);
nand U14743 (N_14743,N_9259,N_11649);
xor U14744 (N_14744,N_10189,N_9925);
nor U14745 (N_14745,N_11810,N_10152);
nor U14746 (N_14746,N_10766,N_10287);
nand U14747 (N_14747,N_10179,N_11147);
and U14748 (N_14748,N_9644,N_10248);
and U14749 (N_14749,N_10311,N_10784);
or U14750 (N_14750,N_11169,N_9755);
xor U14751 (N_14751,N_11868,N_11209);
nand U14752 (N_14752,N_10798,N_11630);
nor U14753 (N_14753,N_9942,N_10576);
and U14754 (N_14754,N_9537,N_9726);
nor U14755 (N_14755,N_9369,N_11401);
or U14756 (N_14756,N_9608,N_9109);
xnor U14757 (N_14757,N_10078,N_9267);
nand U14758 (N_14758,N_11661,N_11561);
nor U14759 (N_14759,N_11122,N_10680);
and U14760 (N_14760,N_10878,N_10459);
nand U14761 (N_14761,N_11089,N_9674);
and U14762 (N_14762,N_10352,N_9597);
nand U14763 (N_14763,N_11817,N_9927);
or U14764 (N_14764,N_10341,N_9483);
nor U14765 (N_14765,N_10790,N_11467);
nor U14766 (N_14766,N_10216,N_10565);
nand U14767 (N_14767,N_11814,N_9246);
and U14768 (N_14768,N_11367,N_11585);
nand U14769 (N_14769,N_11189,N_10292);
or U14770 (N_14770,N_10129,N_9717);
and U14771 (N_14771,N_11279,N_9604);
and U14772 (N_14772,N_11043,N_10681);
nand U14773 (N_14773,N_11547,N_9985);
and U14774 (N_14774,N_9245,N_10876);
or U14775 (N_14775,N_11581,N_10648);
or U14776 (N_14776,N_11000,N_11814);
and U14777 (N_14777,N_9222,N_11298);
nand U14778 (N_14778,N_11515,N_9556);
nor U14779 (N_14779,N_10407,N_9860);
and U14780 (N_14780,N_11412,N_10717);
nor U14781 (N_14781,N_11837,N_10669);
and U14782 (N_14782,N_11103,N_11793);
and U14783 (N_14783,N_9231,N_11574);
nand U14784 (N_14784,N_10971,N_10485);
nor U14785 (N_14785,N_11371,N_10477);
nand U14786 (N_14786,N_11343,N_9008);
and U14787 (N_14787,N_11077,N_11416);
or U14788 (N_14788,N_11495,N_11458);
and U14789 (N_14789,N_9255,N_11764);
nand U14790 (N_14790,N_9464,N_11289);
and U14791 (N_14791,N_9522,N_9047);
nand U14792 (N_14792,N_10188,N_11016);
and U14793 (N_14793,N_11083,N_9976);
or U14794 (N_14794,N_11913,N_11192);
nor U14795 (N_14795,N_11495,N_11932);
nand U14796 (N_14796,N_9952,N_9973);
nand U14797 (N_14797,N_10606,N_10267);
nand U14798 (N_14798,N_11329,N_11996);
nand U14799 (N_14799,N_11707,N_11844);
and U14800 (N_14800,N_10011,N_11884);
or U14801 (N_14801,N_9227,N_11135);
nand U14802 (N_14802,N_10688,N_11131);
nand U14803 (N_14803,N_10121,N_9475);
nand U14804 (N_14804,N_9536,N_11952);
or U14805 (N_14805,N_10869,N_10675);
or U14806 (N_14806,N_10347,N_10228);
nand U14807 (N_14807,N_9790,N_10364);
xnor U14808 (N_14808,N_11223,N_11056);
nor U14809 (N_14809,N_9466,N_10697);
nand U14810 (N_14810,N_10718,N_9777);
or U14811 (N_14811,N_9339,N_11366);
xor U14812 (N_14812,N_11991,N_11151);
nor U14813 (N_14813,N_9673,N_11251);
nand U14814 (N_14814,N_9166,N_10028);
nand U14815 (N_14815,N_9585,N_11795);
or U14816 (N_14816,N_11832,N_9114);
xnor U14817 (N_14817,N_10922,N_9397);
nor U14818 (N_14818,N_9998,N_10393);
nand U14819 (N_14819,N_10477,N_9065);
and U14820 (N_14820,N_10852,N_9746);
and U14821 (N_14821,N_11612,N_11890);
nor U14822 (N_14822,N_10629,N_9944);
nand U14823 (N_14823,N_10281,N_11523);
nor U14824 (N_14824,N_9358,N_11036);
nand U14825 (N_14825,N_11491,N_10023);
and U14826 (N_14826,N_11885,N_10463);
and U14827 (N_14827,N_10686,N_9228);
nand U14828 (N_14828,N_9620,N_9464);
nand U14829 (N_14829,N_11644,N_11404);
or U14830 (N_14830,N_11541,N_10281);
nor U14831 (N_14831,N_10230,N_11522);
or U14832 (N_14832,N_10329,N_11274);
xnor U14833 (N_14833,N_9489,N_9681);
xnor U14834 (N_14834,N_9557,N_10924);
nand U14835 (N_14835,N_10089,N_9504);
xnor U14836 (N_14836,N_10523,N_11193);
or U14837 (N_14837,N_10369,N_11496);
nor U14838 (N_14838,N_11238,N_9348);
or U14839 (N_14839,N_9823,N_10115);
xor U14840 (N_14840,N_10738,N_11621);
and U14841 (N_14841,N_11741,N_10494);
or U14842 (N_14842,N_9532,N_11894);
nand U14843 (N_14843,N_11373,N_11219);
nor U14844 (N_14844,N_9343,N_9950);
nand U14845 (N_14845,N_9038,N_9520);
or U14846 (N_14846,N_10398,N_10747);
or U14847 (N_14847,N_10872,N_9525);
and U14848 (N_14848,N_11385,N_9991);
nand U14849 (N_14849,N_10850,N_9025);
and U14850 (N_14850,N_10838,N_10916);
or U14851 (N_14851,N_11580,N_10050);
xnor U14852 (N_14852,N_9671,N_10412);
nand U14853 (N_14853,N_10331,N_9514);
and U14854 (N_14854,N_11913,N_10377);
nand U14855 (N_14855,N_11541,N_10064);
nand U14856 (N_14856,N_9525,N_11489);
nor U14857 (N_14857,N_9087,N_9316);
nor U14858 (N_14858,N_10025,N_11629);
or U14859 (N_14859,N_9837,N_11401);
or U14860 (N_14860,N_10248,N_11566);
nor U14861 (N_14861,N_10992,N_11440);
nand U14862 (N_14862,N_11088,N_10378);
and U14863 (N_14863,N_11842,N_9218);
or U14864 (N_14864,N_10299,N_9127);
nor U14865 (N_14865,N_9058,N_9675);
and U14866 (N_14866,N_10031,N_11242);
xnor U14867 (N_14867,N_10124,N_10816);
and U14868 (N_14868,N_11435,N_9824);
nor U14869 (N_14869,N_11861,N_9394);
nor U14870 (N_14870,N_10434,N_10355);
nor U14871 (N_14871,N_11684,N_10996);
and U14872 (N_14872,N_11562,N_9257);
and U14873 (N_14873,N_11076,N_11314);
or U14874 (N_14874,N_10785,N_11179);
or U14875 (N_14875,N_11722,N_9610);
nand U14876 (N_14876,N_9556,N_9918);
and U14877 (N_14877,N_10988,N_9664);
and U14878 (N_14878,N_10629,N_9596);
and U14879 (N_14879,N_11771,N_10384);
xnor U14880 (N_14880,N_10467,N_11306);
or U14881 (N_14881,N_9815,N_10171);
xor U14882 (N_14882,N_10124,N_11158);
and U14883 (N_14883,N_9600,N_9851);
nand U14884 (N_14884,N_10138,N_11498);
or U14885 (N_14885,N_11987,N_10307);
and U14886 (N_14886,N_10761,N_11078);
or U14887 (N_14887,N_11471,N_9148);
xnor U14888 (N_14888,N_11901,N_10477);
or U14889 (N_14889,N_9341,N_11339);
nor U14890 (N_14890,N_10974,N_9598);
or U14891 (N_14891,N_10505,N_10390);
nand U14892 (N_14892,N_11196,N_11354);
nor U14893 (N_14893,N_9574,N_10932);
nand U14894 (N_14894,N_9480,N_10012);
nand U14895 (N_14895,N_11814,N_9382);
nor U14896 (N_14896,N_11737,N_10539);
nand U14897 (N_14897,N_9834,N_10363);
nor U14898 (N_14898,N_10127,N_11059);
nand U14899 (N_14899,N_10232,N_9024);
or U14900 (N_14900,N_9465,N_11771);
nand U14901 (N_14901,N_10268,N_9886);
nand U14902 (N_14902,N_9905,N_9206);
xnor U14903 (N_14903,N_9113,N_10507);
and U14904 (N_14904,N_9689,N_10389);
and U14905 (N_14905,N_9720,N_10915);
nor U14906 (N_14906,N_10576,N_10340);
xor U14907 (N_14907,N_11826,N_11311);
nor U14908 (N_14908,N_10807,N_9206);
nand U14909 (N_14909,N_11886,N_11312);
nand U14910 (N_14910,N_9176,N_10189);
and U14911 (N_14911,N_9305,N_10523);
nor U14912 (N_14912,N_10177,N_9531);
and U14913 (N_14913,N_9313,N_10284);
and U14914 (N_14914,N_10631,N_9623);
nor U14915 (N_14915,N_9100,N_10806);
and U14916 (N_14916,N_11644,N_11055);
or U14917 (N_14917,N_10074,N_10568);
nand U14918 (N_14918,N_11181,N_11589);
nand U14919 (N_14919,N_9250,N_10683);
or U14920 (N_14920,N_11486,N_9761);
nor U14921 (N_14921,N_11342,N_9460);
or U14922 (N_14922,N_10352,N_10347);
xnor U14923 (N_14923,N_9998,N_10769);
nor U14924 (N_14924,N_10238,N_9921);
and U14925 (N_14925,N_10878,N_11508);
or U14926 (N_14926,N_11878,N_9418);
nand U14927 (N_14927,N_10768,N_11634);
and U14928 (N_14928,N_9109,N_9658);
nand U14929 (N_14929,N_10247,N_10538);
nand U14930 (N_14930,N_10733,N_11351);
nor U14931 (N_14931,N_10194,N_9228);
and U14932 (N_14932,N_9869,N_11387);
or U14933 (N_14933,N_11924,N_9903);
or U14934 (N_14934,N_11235,N_9050);
nor U14935 (N_14935,N_11778,N_11020);
nand U14936 (N_14936,N_11275,N_11727);
or U14937 (N_14937,N_11103,N_10523);
and U14938 (N_14938,N_11185,N_9487);
nand U14939 (N_14939,N_9430,N_10850);
and U14940 (N_14940,N_9715,N_11971);
or U14941 (N_14941,N_10804,N_10758);
nor U14942 (N_14942,N_11024,N_10716);
and U14943 (N_14943,N_9803,N_10520);
or U14944 (N_14944,N_11743,N_10885);
nand U14945 (N_14945,N_11846,N_9410);
xnor U14946 (N_14946,N_10150,N_9465);
or U14947 (N_14947,N_10760,N_11566);
or U14948 (N_14948,N_10598,N_11509);
nand U14949 (N_14949,N_10966,N_11183);
xor U14950 (N_14950,N_10823,N_10695);
nor U14951 (N_14951,N_9669,N_11449);
or U14952 (N_14952,N_9147,N_10630);
and U14953 (N_14953,N_10427,N_11162);
nand U14954 (N_14954,N_10837,N_10124);
or U14955 (N_14955,N_11965,N_10380);
nor U14956 (N_14956,N_11896,N_10426);
nand U14957 (N_14957,N_11749,N_11030);
nand U14958 (N_14958,N_11397,N_10193);
nor U14959 (N_14959,N_10189,N_10577);
and U14960 (N_14960,N_11176,N_11801);
and U14961 (N_14961,N_9354,N_9795);
or U14962 (N_14962,N_11353,N_11315);
nor U14963 (N_14963,N_11270,N_11063);
or U14964 (N_14964,N_10988,N_11107);
and U14965 (N_14965,N_11231,N_11977);
or U14966 (N_14966,N_11691,N_10644);
nand U14967 (N_14967,N_10866,N_9684);
nor U14968 (N_14968,N_10932,N_11897);
nand U14969 (N_14969,N_11530,N_9344);
nand U14970 (N_14970,N_11248,N_10566);
and U14971 (N_14971,N_11091,N_9939);
and U14972 (N_14972,N_9359,N_10735);
or U14973 (N_14973,N_9159,N_11351);
nor U14974 (N_14974,N_11210,N_11764);
nor U14975 (N_14975,N_10616,N_10388);
nand U14976 (N_14976,N_10585,N_9630);
xnor U14977 (N_14977,N_10452,N_10609);
nor U14978 (N_14978,N_11224,N_11139);
nand U14979 (N_14979,N_10377,N_10732);
or U14980 (N_14980,N_11023,N_10618);
and U14981 (N_14981,N_9590,N_11173);
nand U14982 (N_14982,N_10198,N_10956);
nor U14983 (N_14983,N_10864,N_9743);
nand U14984 (N_14984,N_9959,N_10868);
nor U14985 (N_14985,N_9163,N_10877);
nor U14986 (N_14986,N_9416,N_9075);
nand U14987 (N_14987,N_9375,N_10132);
nor U14988 (N_14988,N_9319,N_11740);
nand U14989 (N_14989,N_10423,N_9957);
xor U14990 (N_14990,N_10823,N_11503);
and U14991 (N_14991,N_10836,N_11692);
and U14992 (N_14992,N_11665,N_11129);
or U14993 (N_14993,N_9094,N_11196);
xor U14994 (N_14994,N_10201,N_11882);
xor U14995 (N_14995,N_10397,N_10904);
or U14996 (N_14996,N_9421,N_10281);
nor U14997 (N_14997,N_11057,N_11906);
nand U14998 (N_14998,N_11218,N_9860);
and U14999 (N_14999,N_10953,N_9447);
nor UO_0 (O_0,N_13908,N_12896);
nand UO_1 (O_1,N_13238,N_12447);
or UO_2 (O_2,N_14079,N_14250);
nand UO_3 (O_3,N_14662,N_14465);
or UO_4 (O_4,N_12308,N_12962);
nor UO_5 (O_5,N_13287,N_14221);
nor UO_6 (O_6,N_14558,N_13781);
nor UO_7 (O_7,N_13638,N_13269);
nand UO_8 (O_8,N_13526,N_12608);
nand UO_9 (O_9,N_12458,N_13285);
nand UO_10 (O_10,N_12049,N_13227);
or UO_11 (O_11,N_13691,N_14811);
and UO_12 (O_12,N_13099,N_13124);
and UO_13 (O_13,N_13839,N_13532);
nand UO_14 (O_14,N_14833,N_12392);
and UO_15 (O_15,N_12290,N_12052);
nand UO_16 (O_16,N_12620,N_13832);
or UO_17 (O_17,N_12588,N_13658);
nor UO_18 (O_18,N_13898,N_14908);
or UO_19 (O_19,N_12941,N_12938);
and UO_20 (O_20,N_13553,N_13828);
nand UO_21 (O_21,N_14059,N_13655);
xnor UO_22 (O_22,N_14522,N_13092);
and UO_23 (O_23,N_12110,N_12966);
or UO_24 (O_24,N_14876,N_14557);
or UO_25 (O_25,N_13510,N_14860);
xnor UO_26 (O_26,N_14169,N_12274);
or UO_27 (O_27,N_14652,N_14252);
xnor UO_28 (O_28,N_13405,N_12200);
or UO_29 (O_29,N_12516,N_14341);
and UO_30 (O_30,N_13882,N_14783);
nor UO_31 (O_31,N_13799,N_14339);
nand UO_32 (O_32,N_14236,N_14987);
or UO_33 (O_33,N_13231,N_13897);
xor UO_34 (O_34,N_13556,N_14620);
and UO_35 (O_35,N_12641,N_13086);
nor UO_36 (O_36,N_14589,N_13535);
or UO_37 (O_37,N_12639,N_14807);
and UO_38 (O_38,N_13743,N_12340);
or UO_39 (O_39,N_12659,N_14259);
and UO_40 (O_40,N_14568,N_14004);
nor UO_41 (O_41,N_13793,N_14520);
nor UO_42 (O_42,N_12387,N_14832);
or UO_43 (O_43,N_14028,N_12633);
nand UO_44 (O_44,N_13083,N_12336);
and UO_45 (O_45,N_14460,N_13049);
nor UO_46 (O_46,N_13712,N_12397);
and UO_47 (O_47,N_13926,N_12517);
and UO_48 (O_48,N_13198,N_14921);
nor UO_49 (O_49,N_14668,N_12804);
nand UO_50 (O_50,N_12578,N_13782);
nand UO_51 (O_51,N_13278,N_13318);
xor UO_52 (O_52,N_13126,N_14730);
nand UO_53 (O_53,N_14477,N_13867);
or UO_54 (O_54,N_12495,N_14065);
xnor UO_55 (O_55,N_14181,N_12982);
xor UO_56 (O_56,N_14809,N_14296);
xor UO_57 (O_57,N_14591,N_14162);
and UO_58 (O_58,N_13180,N_14886);
nor UO_59 (O_59,N_13737,N_12506);
nor UO_60 (O_60,N_13215,N_13572);
or UO_61 (O_61,N_12202,N_14732);
nor UO_62 (O_62,N_12269,N_13508);
nor UO_63 (O_63,N_12595,N_13626);
nand UO_64 (O_64,N_12898,N_13449);
and UO_65 (O_65,N_14316,N_14818);
nand UO_66 (O_66,N_14952,N_12788);
nand UO_67 (O_67,N_14442,N_12039);
or UO_68 (O_68,N_14450,N_13790);
or UO_69 (O_69,N_13068,N_12078);
and UO_70 (O_70,N_13438,N_14814);
nor UO_71 (O_71,N_13938,N_13317);
nand UO_72 (O_72,N_14869,N_13052);
and UO_73 (O_73,N_13309,N_13389);
xnor UO_74 (O_74,N_12371,N_12131);
or UO_75 (O_75,N_13656,N_13365);
nand UO_76 (O_76,N_14214,N_12405);
nand UO_77 (O_77,N_12163,N_14417);
or UO_78 (O_78,N_13053,N_14610);
or UO_79 (O_79,N_13232,N_14267);
or UO_80 (O_80,N_13750,N_14973);
nor UO_81 (O_81,N_12558,N_14717);
or UO_82 (O_82,N_12768,N_14381);
or UO_83 (O_83,N_14999,N_12561);
xor UO_84 (O_84,N_14953,N_12278);
nor UO_85 (O_85,N_13156,N_13073);
nor UO_86 (O_86,N_13878,N_13697);
nor UO_87 (O_87,N_12007,N_12453);
and UO_88 (O_88,N_13142,N_14331);
and UO_89 (O_89,N_12210,N_14085);
xor UO_90 (O_90,N_13200,N_12499);
xnor UO_91 (O_91,N_13015,N_12243);
nor UO_92 (O_92,N_13613,N_12207);
and UO_93 (O_93,N_14487,N_14362);
and UO_94 (O_94,N_14293,N_14102);
nand UO_95 (O_95,N_14824,N_12760);
nor UO_96 (O_96,N_14258,N_14910);
or UO_97 (O_97,N_14675,N_12010);
xor UO_98 (O_98,N_14974,N_14769);
nand UO_99 (O_99,N_13182,N_13672);
nand UO_100 (O_100,N_13186,N_13384);
or UO_101 (O_101,N_14976,N_14173);
or UO_102 (O_102,N_12801,N_13536);
xnor UO_103 (O_103,N_12309,N_14640);
or UO_104 (O_104,N_12892,N_12944);
nand UO_105 (O_105,N_14344,N_14333);
nor UO_106 (O_106,N_14555,N_13950);
nor UO_107 (O_107,N_13701,N_14384);
xor UO_108 (O_108,N_13006,N_13847);
xnor UO_109 (O_109,N_14737,N_13944);
or UO_110 (O_110,N_12741,N_14899);
and UO_111 (O_111,N_12067,N_14884);
nand UO_112 (O_112,N_13353,N_13197);
and UO_113 (O_113,N_14398,N_13632);
and UO_114 (O_114,N_12234,N_12347);
nand UO_115 (O_115,N_12632,N_14639);
xnor UO_116 (O_116,N_13034,N_13393);
and UO_117 (O_117,N_14549,N_14038);
or UO_118 (O_118,N_12777,N_14285);
nor UO_119 (O_119,N_12754,N_14171);
and UO_120 (O_120,N_13968,N_12687);
nand UO_121 (O_121,N_14220,N_12033);
nand UO_122 (O_122,N_12329,N_14887);
xor UO_123 (O_123,N_12541,N_12077);
nor UO_124 (O_124,N_12122,N_14629);
nand UO_125 (O_125,N_14033,N_13071);
and UO_126 (O_126,N_12912,N_13481);
nor UO_127 (O_127,N_13139,N_14667);
nor UO_128 (O_128,N_13520,N_14034);
nand UO_129 (O_129,N_13096,N_14932);
xnor UO_130 (O_130,N_12988,N_13599);
nor UO_131 (O_131,N_13751,N_14305);
nor UO_132 (O_132,N_12865,N_14847);
and UO_133 (O_133,N_13112,N_12648);
and UO_134 (O_134,N_14215,N_12034);
nand UO_135 (O_135,N_13966,N_12601);
xor UO_136 (O_136,N_12083,N_14705);
nand UO_137 (O_137,N_13177,N_13304);
and UO_138 (O_138,N_12220,N_14361);
nor UO_139 (O_139,N_14068,N_14801);
or UO_140 (O_140,N_12197,N_14888);
nor UO_141 (O_141,N_12255,N_13945);
nor UO_142 (O_142,N_13334,N_13690);
xor UO_143 (O_143,N_13943,N_12625);
and UO_144 (O_144,N_12799,N_13522);
nor UO_145 (O_145,N_14495,N_12539);
nor UO_146 (O_146,N_12719,N_14321);
xnor UO_147 (O_147,N_12520,N_13284);
nand UO_148 (O_148,N_12203,N_13918);
and UO_149 (O_149,N_12266,N_13964);
and UO_150 (O_150,N_13970,N_13814);
or UO_151 (O_151,N_13994,N_13028);
nand UO_152 (O_152,N_13218,N_12820);
nor UO_153 (O_153,N_12054,N_13903);
nand UO_154 (O_154,N_14133,N_14759);
and UO_155 (O_155,N_12664,N_12045);
nor UO_156 (O_156,N_13797,N_12808);
nand UO_157 (O_157,N_14441,N_14157);
and UO_158 (O_158,N_13732,N_14731);
nor UO_159 (O_159,N_12649,N_13044);
nand UO_160 (O_160,N_14790,N_13446);
or UO_161 (O_161,N_12745,N_12024);
and UO_162 (O_162,N_13603,N_13758);
nand UO_163 (O_163,N_14686,N_12380);
and UO_164 (O_164,N_12008,N_14660);
and UO_165 (O_165,N_12891,N_14587);
or UO_166 (O_166,N_13120,N_14604);
nand UO_167 (O_167,N_13233,N_13490);
and UO_168 (O_168,N_13720,N_12750);
nor UO_169 (O_169,N_14193,N_13519);
nand UO_170 (O_170,N_14197,N_13072);
or UO_171 (O_171,N_13229,N_12361);
or UO_172 (O_172,N_13596,N_12463);
and UO_173 (O_173,N_14020,N_14622);
nand UO_174 (O_174,N_14284,N_13128);
or UO_175 (O_175,N_12908,N_14377);
nor UO_176 (O_176,N_12021,N_14946);
and UO_177 (O_177,N_14454,N_13116);
nand UO_178 (O_178,N_13211,N_14388);
and UO_179 (O_179,N_13713,N_14778);
nand UO_180 (O_180,N_12116,N_14349);
and UO_181 (O_181,N_13900,N_13779);
nor UO_182 (O_182,N_12417,N_14708);
nand UO_183 (O_183,N_12334,N_12927);
nor UO_184 (O_184,N_13352,N_14984);
and UO_185 (O_185,N_12888,N_13528);
nor UO_186 (O_186,N_14436,N_13696);
nand UO_187 (O_187,N_14325,N_13913);
nor UO_188 (O_188,N_14338,N_12529);
nand UO_189 (O_189,N_12698,N_12064);
nand UO_190 (O_190,N_12814,N_14222);
or UO_191 (O_191,N_13456,N_13412);
nor UO_192 (O_192,N_12422,N_12752);
and UO_193 (O_193,N_14613,N_12838);
or UO_194 (O_194,N_12259,N_12365);
xor UO_195 (O_195,N_13999,N_13702);
nand UO_196 (O_196,N_13400,N_13552);
nand UO_197 (O_197,N_13948,N_13498);
nand UO_198 (O_198,N_12088,N_12240);
nor UO_199 (O_199,N_14843,N_14593);
and UO_200 (O_200,N_13753,N_14617);
or UO_201 (O_201,N_13949,N_13833);
nor UO_202 (O_202,N_14095,N_13491);
nor UO_203 (O_203,N_14890,N_12963);
xor UO_204 (O_204,N_14294,N_12974);
and UO_205 (O_205,N_13167,N_13382);
xnor UO_206 (O_206,N_12564,N_12803);
and UO_207 (O_207,N_12983,N_14143);
or UO_208 (O_208,N_12947,N_14393);
xnor UO_209 (O_209,N_13383,N_12035);
nor UO_210 (O_210,N_12886,N_14019);
nor UO_211 (O_211,N_13496,N_13499);
nor UO_212 (O_212,N_12261,N_13140);
or UO_213 (O_213,N_12840,N_12626);
nand UO_214 (O_214,N_14641,N_12844);
or UO_215 (O_215,N_12644,N_13005);
nor UO_216 (O_216,N_12480,N_14043);
and UO_217 (O_217,N_13051,N_12001);
nor UO_218 (O_218,N_13248,N_12829);
and UO_219 (O_219,N_12043,N_13335);
or UO_220 (O_220,N_12487,N_13623);
nand UO_221 (O_221,N_12575,N_12776);
or UO_222 (O_222,N_12473,N_13978);
and UO_223 (O_223,N_12426,N_14096);
or UO_224 (O_224,N_13069,N_14712);
and UO_225 (O_225,N_12695,N_13663);
or UO_226 (O_226,N_14141,N_12350);
nand UO_227 (O_227,N_13735,N_12222);
and UO_228 (O_228,N_14868,N_12618);
nor UO_229 (O_229,N_13346,N_13617);
xnor UO_230 (O_230,N_14468,N_13630);
or UO_231 (O_231,N_14158,N_13547);
and UO_232 (O_232,N_13721,N_13056);
xnor UO_233 (O_233,N_13609,N_13018);
nand UO_234 (O_234,N_14088,N_14430);
and UO_235 (O_235,N_13150,N_14392);
or UO_236 (O_236,N_12469,N_13776);
and UO_237 (O_237,N_13555,N_14047);
and UO_238 (O_238,N_14894,N_14146);
nor UO_239 (O_239,N_12374,N_14155);
nor UO_240 (O_240,N_13286,N_14201);
nor UO_241 (O_241,N_14838,N_13095);
and UO_242 (O_242,N_12859,N_12174);
and UO_243 (O_243,N_14202,N_13157);
or UO_244 (O_244,N_14409,N_12009);
or UO_245 (O_245,N_12032,N_14751);
or UO_246 (O_246,N_14334,N_13322);
and UO_247 (O_247,N_13694,N_13893);
and UO_248 (O_248,N_13674,N_14231);
nor UO_249 (O_249,N_14094,N_12419);
nand UO_250 (O_250,N_14251,N_12522);
nor UO_251 (O_251,N_14056,N_12738);
and UO_252 (O_252,N_14014,N_13969);
and UO_253 (O_253,N_13250,N_12399);
or UO_254 (O_254,N_12688,N_13298);
and UO_255 (O_255,N_12931,N_14839);
nor UO_256 (O_256,N_13469,N_14722);
or UO_257 (O_257,N_13419,N_12500);
nand UO_258 (O_258,N_13635,N_12398);
nand UO_259 (O_259,N_12589,N_13660);
nor UO_260 (O_260,N_13507,N_13710);
nand UO_261 (O_261,N_14343,N_12985);
xnor UO_262 (O_262,N_12494,N_14186);
or UO_263 (O_263,N_12680,N_14656);
nand UO_264 (O_264,N_14916,N_12766);
xnor UO_265 (O_265,N_12530,N_14788);
nand UO_266 (O_266,N_12742,N_13870);
nor UO_267 (O_267,N_13641,N_12345);
and UO_268 (O_268,N_13879,N_14434);
or UO_269 (O_269,N_13187,N_14996);
or UO_270 (O_270,N_13729,N_12646);
nor UO_271 (O_271,N_13026,N_14831);
nand UO_272 (O_272,N_14103,N_12383);
nand UO_273 (O_273,N_14299,N_13646);
and UO_274 (O_274,N_14954,N_13173);
and UO_275 (O_275,N_13319,N_13762);
nor UO_276 (O_276,N_13835,N_14947);
and UO_277 (O_277,N_12519,N_12903);
or UO_278 (O_278,N_13461,N_12662);
and UO_279 (O_279,N_12882,N_14590);
and UO_280 (O_280,N_14718,N_12136);
and UO_281 (O_281,N_14484,N_12976);
or UO_282 (O_282,N_12895,N_14951);
nor UO_283 (O_283,N_12604,N_12735);
xnor UO_284 (O_284,N_14342,N_13889);
or UO_285 (O_285,N_14904,N_14612);
and UO_286 (O_286,N_12421,N_12102);
nand UO_287 (O_287,N_14725,N_14402);
nor UO_288 (O_288,N_14758,N_12536);
or UO_289 (O_289,N_13416,N_14998);
or UO_290 (O_290,N_13002,N_13350);
nand UO_291 (O_291,N_12123,N_12733);
or UO_292 (O_292,N_13460,N_12094);
nand UO_293 (O_293,N_12030,N_13965);
nand UO_294 (O_294,N_13385,N_13470);
and UO_295 (O_295,N_13927,N_12438);
or UO_296 (O_296,N_13208,N_14961);
nor UO_297 (O_297,N_13117,N_14723);
nor UO_298 (O_298,N_14665,N_12609);
nor UO_299 (O_299,N_13752,N_12250);
or UO_300 (O_300,N_13806,N_13653);
or UO_301 (O_301,N_14885,N_14923);
or UO_302 (O_302,N_14217,N_14407);
nand UO_303 (O_303,N_13136,N_12691);
or UO_304 (O_304,N_12711,N_13910);
nand UO_305 (O_305,N_14914,N_12171);
xnor UO_306 (O_306,N_14000,N_12022);
nand UO_307 (O_307,N_13807,N_13819);
nor UO_308 (O_308,N_14435,N_12429);
xor UO_309 (O_309,N_12180,N_13363);
nor UO_310 (O_310,N_14235,N_13820);
and UO_311 (O_311,N_13447,N_14965);
nand UO_312 (O_312,N_14073,N_13853);
nand UO_313 (O_313,N_13291,N_14556);
nand UO_314 (O_314,N_12304,N_14672);
nor UO_315 (O_315,N_12277,N_14286);
and UO_316 (O_316,N_12228,N_12343);
nand UO_317 (O_317,N_13024,N_14208);
or UO_318 (O_318,N_12323,N_13967);
nand UO_319 (O_319,N_13714,N_12349);
and UO_320 (O_320,N_12806,N_13974);
nor UO_321 (O_321,N_12224,N_12322);
nor UO_322 (O_322,N_12932,N_13736);
or UO_323 (O_323,N_14658,N_13722);
nor UO_324 (O_324,N_14364,N_12928);
nand UO_325 (O_325,N_12362,N_13669);
and UO_326 (O_326,N_14109,N_13122);
nand UO_327 (O_327,N_12360,N_13105);
nand UO_328 (O_328,N_14849,N_12000);
nor UO_329 (O_329,N_12684,N_13109);
or UO_330 (O_330,N_12969,N_12562);
nor UO_331 (O_331,N_12843,N_14741);
or UO_332 (O_332,N_12679,N_13562);
nand UO_333 (O_333,N_14880,N_12379);
or UO_334 (O_334,N_13257,N_12979);
xnor UO_335 (O_335,N_13864,N_14142);
and UO_336 (O_336,N_13682,N_12491);
and UO_337 (O_337,N_14359,N_12297);
and UO_338 (O_338,N_12005,N_14927);
and UO_339 (O_339,N_14076,N_14470);
nand UO_340 (O_340,N_13225,N_12787);
nor UO_341 (O_341,N_14992,N_14949);
and UO_342 (O_342,N_13260,N_13076);
or UO_343 (O_343,N_12701,N_12521);
nand UO_344 (O_344,N_13295,N_12574);
nor UO_345 (O_345,N_14988,N_14871);
nand UO_346 (O_346,N_14785,N_14154);
nor UO_347 (O_347,N_13444,N_14663);
xnor UO_348 (O_348,N_13516,N_14913);
xor UO_349 (O_349,N_12337,N_14503);
nand UO_350 (O_350,N_12702,N_14905);
or UO_351 (O_351,N_14982,N_14950);
nor UO_352 (O_352,N_14330,N_14453);
or UO_353 (O_353,N_14968,N_13571);
nand UO_354 (O_354,N_12954,N_13206);
nand UO_355 (O_355,N_13530,N_12040);
nor UO_356 (O_356,N_14791,N_13217);
nor UO_357 (O_357,N_13786,N_12864);
or UO_358 (O_358,N_12845,N_14599);
or UO_359 (O_359,N_13642,N_14755);
and UO_360 (O_360,N_12977,N_12211);
nand UO_361 (O_361,N_13524,N_13754);
nand UO_362 (O_362,N_12214,N_12716);
and UO_363 (O_363,N_13021,N_14491);
xor UO_364 (O_364,N_14606,N_14067);
or UO_365 (O_365,N_14767,N_14086);
nand UO_366 (O_366,N_13203,N_14579);
and UO_367 (O_367,N_12998,N_13022);
and UO_368 (O_368,N_13125,N_12879);
or UO_369 (O_369,N_14699,N_14114);
and UO_370 (O_370,N_14931,N_12472);
or UO_371 (O_371,N_12786,N_12128);
and UO_372 (O_372,N_14496,N_13244);
or UO_373 (O_373,N_12660,N_12580);
nand UO_374 (O_374,N_14623,N_12948);
nand UO_375 (O_375,N_14489,N_12016);
nand UO_376 (O_376,N_14499,N_13281);
nor UO_377 (O_377,N_13147,N_13940);
nor UO_378 (O_378,N_14308,N_12743);
or UO_379 (O_379,N_14850,N_13375);
xnor UO_380 (O_380,N_12586,N_13860);
xnor UO_381 (O_381,N_14415,N_12942);
xor UO_382 (O_382,N_14255,N_13100);
and UO_383 (O_383,N_14238,N_12540);
nor UO_384 (O_384,N_12263,N_13598);
and UO_385 (O_385,N_12771,N_14304);
or UO_386 (O_386,N_13282,N_13445);
nand UO_387 (O_387,N_14892,N_12183);
nand UO_388 (O_388,N_13240,N_14837);
xnor UO_389 (O_389,N_12086,N_12490);
nand UO_390 (O_390,N_13894,N_12201);
or UO_391 (O_391,N_13012,N_14097);
or UO_392 (O_392,N_14355,N_13747);
or UO_393 (O_393,N_14408,N_13418);
and UO_394 (O_394,N_13262,N_14414);
xnor UO_395 (O_395,N_12582,N_13627);
xnor UO_396 (O_396,N_13379,N_12185);
nor UO_397 (O_397,N_14633,N_14775);
or UO_398 (O_398,N_14479,N_14041);
nand UO_399 (O_399,N_12746,N_14352);
or UO_400 (O_400,N_13473,N_14175);
nand UO_401 (O_401,N_13141,N_14071);
or UO_402 (O_402,N_12599,N_13110);
and UO_403 (O_403,N_12025,N_13388);
or UO_404 (O_404,N_12736,N_12456);
and UO_405 (O_405,N_14649,N_12717);
nor UO_406 (O_406,N_13356,N_14264);
xnor UO_407 (O_407,N_13132,N_12946);
nand UO_408 (O_408,N_13414,N_13146);
and UO_409 (O_409,N_12241,N_14875);
nor UO_410 (O_410,N_14830,N_12055);
nor UO_411 (O_411,N_12189,N_14118);
nand UO_412 (O_412,N_14955,N_13153);
nor UO_413 (O_413,N_14419,N_14403);
nand UO_414 (O_414,N_13858,N_12342);
and UO_415 (O_415,N_12177,N_12591);
or UO_416 (O_416,N_13851,N_12437);
or UO_417 (O_417,N_13265,N_12957);
and UO_418 (O_418,N_14077,N_13990);
and UO_419 (O_419,N_14821,N_14091);
or UO_420 (O_420,N_13176,N_14529);
nor UO_421 (O_421,N_12098,N_13805);
and UO_422 (O_422,N_14099,N_13671);
nor UO_423 (O_423,N_13035,N_12284);
nor UO_424 (O_424,N_12643,N_13339);
xor UO_425 (O_425,N_13154,N_14716);
nand UO_426 (O_426,N_12440,N_12556);
and UO_427 (O_427,N_13594,N_12002);
or UO_428 (O_428,N_12156,N_12666);
and UO_429 (O_429,N_13583,N_13725);
or UO_430 (O_430,N_12554,N_12272);
and UO_431 (O_431,N_14650,N_13149);
nor UO_432 (O_432,N_14780,N_13667);
nand UO_433 (O_433,N_12195,N_13822);
xnor UO_434 (O_434,N_12471,N_13395);
nand UO_435 (O_435,N_14152,N_13560);
nand UO_436 (O_436,N_12512,N_13324);
nor UO_437 (O_437,N_14366,N_12720);
and UO_438 (O_438,N_13728,N_14291);
nand UO_439 (O_439,N_12312,N_13953);
xnor UO_440 (O_440,N_12479,N_14163);
xnor UO_441 (O_441,N_13791,N_14159);
or UO_442 (O_442,N_12690,N_13774);
and UO_443 (O_443,N_12503,N_12921);
xnor UO_444 (O_444,N_14789,N_12467);
or UO_445 (O_445,N_13249,N_12668);
xor UO_446 (O_446,N_12231,N_14054);
nand UO_447 (O_447,N_12148,N_12138);
nor UO_448 (O_448,N_13031,N_13130);
or UO_449 (O_449,N_13801,N_14371);
xor UO_450 (O_450,N_14140,N_13152);
and UO_451 (O_451,N_13045,N_12769);
nand UO_452 (O_452,N_14834,N_12774);
or UO_453 (O_453,N_14792,N_13606);
nor UO_454 (O_454,N_13123,N_12542);
nor UO_455 (O_455,N_13330,N_12810);
xor UO_456 (O_456,N_13253,N_14995);
or UO_457 (O_457,N_13995,N_14439);
and UO_458 (O_458,N_13545,N_12739);
nor UO_459 (O_459,N_14756,N_12455);
and UO_460 (O_460,N_13947,N_12454);
nand UO_461 (O_461,N_14265,N_12109);
nor UO_462 (O_462,N_13133,N_12074);
nand UO_463 (O_463,N_12511,N_13289);
nor UO_464 (O_464,N_12204,N_13796);
or UO_465 (O_465,N_13463,N_14160);
and UO_466 (O_466,N_12598,N_12728);
nand UO_467 (O_467,N_13573,N_14196);
and UO_468 (O_468,N_12925,N_12433);
nand UO_469 (O_469,N_13258,N_14538);
and UO_470 (O_470,N_13033,N_12264);
or UO_471 (O_471,N_12610,N_14474);
xnor UO_472 (O_472,N_13237,N_13201);
and UO_473 (O_473,N_14287,N_13001);
nand UO_474 (O_474,N_13849,N_14124);
or UO_475 (O_475,N_14768,N_14332);
nor UO_476 (O_476,N_14478,N_12172);
nor UO_477 (O_477,N_12442,N_13550);
and UO_478 (O_478,N_13517,N_14926);
and UO_479 (O_479,N_12873,N_13242);
nand UO_480 (O_480,N_13081,N_13778);
nor UO_481 (O_481,N_14989,N_14446);
nand UO_482 (O_482,N_13195,N_12747);
nor UO_483 (O_483,N_13955,N_14156);
and UO_484 (O_484,N_12121,N_14482);
and UO_485 (O_485,N_13880,N_13676);
nand UO_486 (O_486,N_12410,N_12909);
or UO_487 (O_487,N_12108,N_13474);
nand UO_488 (O_488,N_13094,N_13928);
or UO_489 (O_489,N_14323,N_13301);
xor UO_490 (O_490,N_14037,N_13810);
nand UO_491 (O_491,N_12945,N_13794);
or UO_492 (O_492,N_14681,N_12492);
and UO_493 (O_493,N_13693,N_13825);
or UO_494 (O_494,N_13220,N_12670);
or UO_495 (O_495,N_13325,N_12685);
nand UO_496 (O_496,N_14506,N_14177);
or UO_497 (O_497,N_13429,N_14375);
and UO_498 (O_498,N_13888,N_14544);
nor UO_499 (O_499,N_14570,N_12727);
nor UO_500 (O_500,N_14205,N_12451);
and UO_501 (O_501,N_12028,N_13299);
and UO_502 (O_502,N_13360,N_14721);
nand UO_503 (O_503,N_13397,N_13380);
nor UO_504 (O_504,N_14011,N_13462);
nand UO_505 (O_505,N_12647,N_14327);
or UO_506 (O_506,N_13436,N_14507);
nand UO_507 (O_507,N_13221,N_12862);
or UO_508 (O_508,N_12911,N_14353);
nor UO_509 (O_509,N_12987,N_12640);
nand UO_510 (O_510,N_13840,N_14523);
nand UO_511 (O_511,N_13929,N_13951);
xor UO_512 (O_512,N_13707,N_13019);
nor UO_513 (O_513,N_14456,N_13738);
and UO_514 (O_514,N_14936,N_14219);
or UO_515 (O_515,N_12481,N_12097);
xor UO_516 (O_516,N_12151,N_13270);
nor UO_517 (O_517,N_14621,N_13312);
xnor UO_518 (O_518,N_12295,N_14720);
and UO_519 (O_519,N_14190,N_14695);
nor UO_520 (O_520,N_12420,N_14314);
nor UO_521 (O_521,N_12310,N_13486);
nand UO_522 (O_522,N_12816,N_12006);
nand UO_523 (O_523,N_13621,N_14087);
nand UO_524 (O_524,N_14112,N_12393);
or UO_525 (O_525,N_12584,N_12069);
nor UO_526 (O_526,N_12215,N_13523);
nor UO_527 (O_527,N_12622,N_14464);
nor UO_528 (O_528,N_13158,N_12444);
or UO_529 (O_529,N_13209,N_13297);
and UO_530 (O_530,N_12676,N_13219);
nand UO_531 (O_531,N_13804,N_13064);
or UO_532 (O_532,N_13196,N_12568);
nand UO_533 (O_533,N_14859,N_13692);
nor UO_534 (O_534,N_14081,N_13578);
or UO_535 (O_535,N_14107,N_12856);
and UO_536 (O_536,N_12412,N_12877);
nand UO_537 (O_537,N_14203,N_13687);
or UO_538 (O_538,N_14745,N_12567);
nor UO_539 (O_539,N_14248,N_12683);
xor UO_540 (O_540,N_12939,N_12518);
and UO_541 (O_541,N_13563,N_14851);
and UO_542 (O_542,N_14929,N_12286);
nand UO_543 (O_543,N_14661,N_13962);
nor UO_544 (O_544,N_13543,N_14324);
or UO_545 (O_545,N_13040,N_14137);
or UO_546 (O_546,N_12524,N_13235);
and UO_547 (O_547,N_14609,N_13254);
or UO_548 (O_548,N_12436,N_14760);
nand UO_549 (O_549,N_13351,N_14298);
nor UO_550 (O_550,N_14684,N_14089);
xor UO_551 (O_551,N_14796,N_12497);
and UO_552 (O_552,N_14270,N_14282);
and UO_553 (O_553,N_13424,N_13595);
and UO_554 (O_554,N_14879,N_14057);
xor UO_555 (O_555,N_14611,N_12150);
nor UO_556 (O_556,N_12370,N_14654);
nand UO_557 (O_557,N_13746,N_14711);
nor UO_558 (O_558,N_12046,N_13885);
nand UO_559 (O_559,N_13294,N_13426);
or UO_560 (O_560,N_14689,N_14659);
nor UO_561 (O_561,N_12675,N_12906);
nand UO_562 (O_562,N_13090,N_12548);
nor UO_563 (O_563,N_14426,N_14404);
and UO_564 (O_564,N_13997,N_13430);
nand UO_565 (O_565,N_12872,N_14933);
nor UO_566 (O_566,N_12459,N_13433);
nor UO_567 (O_567,N_12192,N_14438);
nor UO_568 (O_568,N_14883,N_13194);
or UO_569 (O_569,N_12894,N_12441);
and UO_570 (O_570,N_12606,N_14704);
or UO_571 (O_571,N_13611,N_13493);
and UO_572 (O_572,N_13011,N_12176);
and UO_573 (O_573,N_12861,N_14505);
nor UO_574 (O_574,N_12645,N_12461);
xnor UO_575 (O_575,N_13812,N_13391);
nand UO_576 (O_576,N_13003,N_14182);
nor UO_577 (O_577,N_14480,N_13061);
nand UO_578 (O_578,N_12607,N_13204);
nand UO_579 (O_579,N_13214,N_12770);
or UO_580 (O_580,N_14084,N_12173);
nand UO_581 (O_581,N_13210,N_13717);
xor UO_582 (O_582,N_13163,N_13347);
nand UO_583 (O_583,N_12179,N_12279);
and UO_584 (O_584,N_14249,N_13368);
nand UO_585 (O_585,N_12325,N_13645);
nand UO_586 (O_586,N_13946,N_13467);
xor UO_587 (O_587,N_14782,N_12373);
and UO_588 (O_588,N_14064,N_14254);
nor UO_589 (O_589,N_14906,N_14511);
or UO_590 (O_590,N_12085,N_12686);
or UO_591 (O_591,N_13981,N_13681);
or UO_592 (O_592,N_14626,N_13772);
or UO_593 (O_593,N_12205,N_12273);
nor UO_594 (O_594,N_12191,N_14645);
or UO_595 (O_595,N_13700,N_14433);
or UO_596 (O_596,N_14230,N_14977);
or UO_597 (O_597,N_13868,N_12658);
or UO_598 (O_598,N_12830,N_13979);
xor UO_599 (O_599,N_13009,N_13841);
nand UO_600 (O_600,N_12155,N_14376);
and UO_601 (O_601,N_13537,N_14753);
or UO_602 (O_602,N_14498,N_12445);
nand UO_603 (O_603,N_12407,N_12302);
and UO_604 (O_604,N_13371,N_14893);
xnor UO_605 (O_605,N_13057,N_12612);
and UO_606 (O_606,N_13581,N_13976);
or UO_607 (O_607,N_12020,N_12199);
or UO_608 (O_608,N_13933,N_13652);
nor UO_609 (O_609,N_14136,N_13151);
nand UO_610 (O_610,N_12216,N_12068);
and UO_611 (O_611,N_14147,N_14896);
and UO_612 (O_612,N_13307,N_14389);
and UO_613 (O_613,N_14794,N_12635);
xnor UO_614 (O_614,N_12364,N_14452);
xor UO_615 (O_615,N_14198,N_14713);
nand UO_616 (O_616,N_14601,N_14986);
xor UO_617 (O_617,N_14062,N_14260);
and UO_618 (O_618,N_13305,N_13895);
nand UO_619 (O_619,N_14049,N_14799);
nand UO_620 (O_620,N_14696,N_12624);
and UO_621 (O_621,N_12315,N_12029);
or UO_622 (O_622,N_13887,N_13127);
nand UO_623 (O_623,N_14483,N_14853);
or UO_624 (O_624,N_13328,N_14535);
and UO_625 (O_625,N_14052,N_14981);
or UO_626 (O_626,N_13355,N_12117);
or UO_627 (O_627,N_12823,N_12485);
xnor UO_628 (O_628,N_14237,N_14437);
or UO_629 (O_629,N_12917,N_12807);
and UO_630 (O_630,N_12508,N_12933);
nand UO_631 (O_631,N_14310,N_13431);
or UO_632 (O_632,N_14669,N_12395);
nor UO_633 (O_633,N_12565,N_14774);
or UO_634 (O_634,N_12999,N_13811);
or UO_635 (O_635,N_12375,N_12827);
nor UO_636 (O_636,N_14582,N_12496);
nand UO_637 (O_637,N_14597,N_13783);
or UO_638 (O_638,N_12423,N_12338);
nand UO_639 (O_639,N_13016,N_13205);
nor UO_640 (O_640,N_12353,N_14174);
or UO_641 (O_641,N_14090,N_14687);
nor UO_642 (O_642,N_12368,N_13857);
nor UO_643 (O_643,N_14706,N_13925);
nor UO_644 (O_644,N_13677,N_13077);
and UO_645 (O_645,N_13310,N_13472);
nor UO_646 (O_646,N_14228,N_13020);
nor UO_647 (O_647,N_13715,N_14979);
and UO_648 (O_648,N_13089,N_13337);
nor UO_649 (O_649,N_13919,N_14030);
or UO_650 (O_650,N_12835,N_14312);
and UO_651 (O_651,N_12206,N_14069);
or UO_652 (O_652,N_14566,N_12825);
or UO_653 (O_653,N_13525,N_14471);
nand UO_654 (O_654,N_13952,N_13364);
or UO_655 (O_655,N_12093,N_12306);
nor UO_656 (O_656,N_12318,N_12615);
or UO_657 (O_657,N_14559,N_12846);
and UO_658 (O_658,N_13896,N_13457);
nand UO_659 (O_659,N_12837,N_14701);
nand UO_660 (O_660,N_14815,N_12722);
or UO_661 (O_661,N_14542,N_12793);
or UO_662 (O_662,N_14564,N_14239);
or UO_663 (O_663,N_13129,N_12141);
nor UO_664 (O_664,N_12531,N_12693);
and UO_665 (O_665,N_14545,N_12430);
and UO_666 (O_666,N_12959,N_13106);
or UO_667 (O_667,N_14592,N_13039);
nand UO_668 (O_668,N_13354,N_13155);
nand UO_669 (O_669,N_14715,N_13567);
nor UO_670 (O_670,N_12332,N_13080);
nor UO_671 (O_671,N_13876,N_12681);
nor UO_672 (O_672,N_12884,N_13531);
nor UO_673 (O_673,N_13922,N_14881);
and UO_674 (O_674,N_13427,N_14856);
xnor UO_675 (O_675,N_12061,N_12474);
and UO_676 (O_676,N_13394,N_14448);
nor UO_677 (O_677,N_14967,N_13800);
and UO_678 (O_678,N_12378,N_14710);
nand UO_679 (O_679,N_12981,N_12817);
or UO_680 (O_680,N_14416,N_14993);
xnor UO_681 (O_681,N_13251,N_12973);
or UO_682 (O_682,N_12505,N_14677);
and UO_683 (O_683,N_14541,N_14340);
or UO_684 (O_684,N_14144,N_14042);
nor UO_685 (O_685,N_14120,N_13538);
xnor UO_686 (O_686,N_14280,N_13873);
and UO_687 (O_687,N_14105,N_13111);
and UO_688 (O_688,N_12486,N_12106);
and UO_689 (O_689,N_14382,N_12293);
or UO_690 (O_690,N_12725,N_12775);
nand UO_691 (O_691,N_13245,N_13138);
or UO_692 (O_692,N_12080,N_13376);
nand UO_693 (O_693,N_13875,N_13622);
or UO_694 (O_694,N_13326,N_13074);
or UO_695 (O_695,N_12922,N_14111);
and UO_696 (O_696,N_14490,N_14131);
xnor UO_697 (O_697,N_13514,N_12587);
or UO_698 (O_698,N_12143,N_13234);
nor UO_699 (O_699,N_14707,N_14106);
nor UO_700 (O_700,N_12357,N_13802);
or UO_701 (O_701,N_12756,N_12634);
nand UO_702 (O_702,N_14827,N_13554);
nand UO_703 (O_703,N_14588,N_13678);
or UO_704 (O_704,N_14719,N_13280);
nor UO_705 (O_705,N_13010,N_13861);
xor UO_706 (O_706,N_13527,N_12653);
nand UO_707 (O_707,N_13175,N_14431);
or UO_708 (O_708,N_13345,N_14029);
nor UO_709 (O_709,N_14051,N_14846);
and UO_710 (O_710,N_13332,N_14966);
nand UO_711 (O_711,N_13370,N_13785);
and UO_712 (O_712,N_13293,N_13769);
or UO_713 (O_713,N_14600,N_12652);
or UO_714 (O_714,N_13963,N_13592);
nand UO_715 (O_715,N_14007,N_13359);
or UO_716 (O_716,N_12044,N_12048);
and UO_717 (O_717,N_12858,N_12144);
or UO_718 (O_718,N_14941,N_12961);
nand UO_719 (O_719,N_14060,N_12314);
nand UO_720 (O_720,N_13357,N_12972);
nand UO_721 (O_721,N_12344,N_14734);
nor UO_722 (O_722,N_12782,N_12401);
nand UO_723 (O_723,N_14918,N_13458);
or UO_724 (O_724,N_13975,N_14922);
nand UO_725 (O_725,N_12706,N_12415);
xnor UO_726 (O_726,N_14671,N_13649);
nor UO_727 (O_727,N_13726,N_12994);
nand UO_728 (O_728,N_14309,N_12388);
or UO_729 (O_729,N_14003,N_13871);
or UO_730 (O_730,N_13048,N_14781);
xnor UO_731 (O_731,N_14036,N_12710);
nand UO_732 (O_732,N_12301,N_13343);
or UO_733 (O_733,N_14816,N_13763);
and UO_734 (O_734,N_12547,N_13041);
nor UO_735 (O_735,N_12789,N_12071);
or UO_736 (O_736,N_12753,N_14802);
or UO_737 (O_737,N_13954,N_14519);
and UO_738 (O_738,N_13892,N_13450);
xnor UO_739 (O_739,N_14528,N_13580);
and UO_740 (O_740,N_12970,N_13620);
or UO_741 (O_741,N_14165,N_12260);
and UO_742 (O_742,N_13865,N_13629);
or UO_743 (O_743,N_14319,N_14421);
or UO_744 (O_744,N_12363,N_14379);
or UO_745 (O_745,N_13546,N_13143);
xnor UO_746 (O_746,N_13213,N_12715);
nor UO_747 (O_747,N_12047,N_14346);
nor UO_748 (O_748,N_14550,N_14018);
or UO_749 (O_749,N_13273,N_13296);
nand UO_750 (O_750,N_13777,N_13809);
or UO_751 (O_751,N_14191,N_13760);
and UO_752 (O_752,N_13991,N_12167);
or UO_753 (O_753,N_13703,N_13684);
xnor UO_754 (O_754,N_13259,N_12305);
nand UO_755 (O_755,N_14930,N_14812);
or UO_756 (O_756,N_12217,N_12213);
nor UO_757 (O_757,N_13386,N_14845);
or UO_758 (O_758,N_14634,N_14469);
nand UO_759 (O_759,N_14180,N_12339);
or UO_760 (O_760,N_14045,N_14023);
or UO_761 (O_761,N_12427,N_13848);
nand UO_762 (O_762,N_14098,N_13484);
and UO_763 (O_763,N_12208,N_12790);
nand UO_764 (O_764,N_13521,N_12854);
xor UO_765 (O_765,N_12245,N_13568);
and UO_766 (O_766,N_14678,N_14288);
nor UO_767 (O_767,N_12682,N_13387);
nor UO_768 (O_768,N_12256,N_14027);
or UO_769 (O_769,N_13957,N_12832);
nor UO_770 (O_770,N_13171,N_14560);
xnor UO_771 (O_771,N_12826,N_12307);
nor UO_772 (O_772,N_14631,N_13495);
nand UO_773 (O_773,N_14497,N_13960);
nor UO_774 (O_774,N_14583,N_12936);
nor UO_775 (O_775,N_13756,N_14153);
nand UO_776 (O_776,N_14614,N_14501);
nand UO_777 (O_777,N_14602,N_14822);
nand UO_778 (O_778,N_13668,N_14554);
xnor UO_779 (O_779,N_13813,N_14595);
or UO_780 (O_780,N_12113,N_12737);
or UO_781 (O_781,N_12878,N_14357);
nand UO_782 (O_782,N_14857,N_12317);
and UO_783 (O_783,N_14900,N_12755);
or UO_784 (O_784,N_13134,N_12051);
nand UO_785 (O_785,N_12800,N_13659);
nand UO_786 (O_786,N_13539,N_14543);
and UO_787 (O_787,N_12821,N_13185);
or UO_788 (O_788,N_13585,N_12311);
nor UO_789 (O_789,N_13855,N_12283);
xor UO_790 (O_790,N_14673,N_12718);
or UO_791 (O_791,N_13640,N_12538);
nand UO_792 (O_792,N_12124,N_14113);
and UO_793 (O_793,N_12603,N_13850);
xor UO_794 (O_794,N_13004,N_13428);
or UO_795 (O_795,N_12251,N_12139);
or UO_796 (O_796,N_12740,N_14272);
and UO_797 (O_797,N_14729,N_13723);
nand UO_798 (O_798,N_12457,N_13959);
nor UO_799 (O_799,N_13787,N_14139);
and UO_800 (O_800,N_12285,N_12993);
nand UO_801 (O_801,N_12893,N_13891);
nand UO_802 (O_802,N_12450,N_14971);
nor UO_803 (O_803,N_13277,N_12327);
and UO_804 (O_804,N_12324,N_12075);
nor UO_805 (O_805,N_13561,N_13193);
and UO_806 (O_806,N_13492,N_12899);
or UO_807 (O_807,N_12478,N_14647);
or UO_808 (O_808,N_13261,N_12763);
or UO_809 (O_809,N_14690,N_12133);
nor UO_810 (O_810,N_13559,N_13733);
xor UO_811 (O_811,N_14326,N_12470);
xnor UO_812 (O_812,N_13471,N_14363);
or UO_813 (O_813,N_12619,N_12239);
nor UO_814 (O_814,N_14078,N_14763);
nor UO_815 (O_815,N_14048,N_13181);
or UO_816 (O_816,N_14540,N_13615);
nor UO_817 (O_817,N_12372,N_14939);
nor UO_818 (O_818,N_12855,N_14682);
xnor UO_819 (O_819,N_12237,N_14347);
nand UO_820 (O_820,N_13078,N_12851);
xor UO_821 (O_821,N_12298,N_12227);
or UO_822 (O_822,N_12798,N_12950);
or UO_823 (O_823,N_13619,N_13390);
or UO_824 (O_824,N_13378,N_13610);
and UO_825 (O_825,N_12581,N_12654);
nor UO_826 (O_826,N_12056,N_14279);
nor UO_827 (O_827,N_12705,N_13453);
or UO_828 (O_828,N_14277,N_14997);
xor UO_829 (O_829,N_14844,N_13212);
xor UO_830 (O_830,N_14798,N_13362);
nand UO_831 (O_831,N_14066,N_14247);
and UO_832 (O_832,N_12918,N_14691);
nand UO_833 (O_833,N_12280,N_14206);
nor UO_834 (O_834,N_12592,N_12852);
nand UO_835 (O_835,N_13466,N_13789);
xnor UO_836 (O_836,N_12870,N_14213);
xor UO_837 (O_837,N_12848,N_13937);
nor UO_838 (O_838,N_12700,N_12159);
nand UO_839 (O_839,N_14727,N_14624);
and UO_840 (O_840,N_14373,N_12560);
and UO_841 (O_841,N_14127,N_13906);
and UO_842 (O_842,N_14183,N_12291);
and UO_843 (O_843,N_12980,N_13098);
and UO_844 (O_844,N_14990,N_13403);
and UO_845 (O_845,N_14164,N_14991);
nand UO_846 (O_846,N_13494,N_14370);
xor UO_847 (O_847,N_14122,N_13744);
nand UO_848 (O_848,N_13941,N_14608);
and UO_849 (O_849,N_12073,N_12623);
and UO_850 (O_850,N_12761,N_12570);
nand UO_851 (O_851,N_12638,N_14110);
and UO_852 (O_852,N_13631,N_13113);
nor UO_853 (O_853,N_14736,N_14225);
and UO_854 (O_854,N_13600,N_13836);
nand UO_855 (O_855,N_12477,N_12650);
or UO_856 (O_856,N_14742,N_14017);
or UO_857 (O_857,N_14411,N_12188);
nor UO_858 (O_858,N_14700,N_14396);
nor UO_859 (O_859,N_12004,N_12394);
nor UO_860 (O_860,N_12079,N_14810);
nor UO_861 (O_861,N_14149,N_13683);
nand UO_862 (O_862,N_14960,N_13636);
nand UO_863 (O_863,N_14009,N_12513);
nor UO_864 (O_864,N_13795,N_12778);
or UO_865 (O_865,N_12535,N_13934);
nor UO_866 (O_866,N_12232,N_13070);
nor UO_867 (O_867,N_12875,N_13834);
nor UO_868 (O_868,N_12537,N_12792);
or UO_869 (O_869,N_13059,N_13501);
nor UO_870 (O_870,N_12866,N_12355);
nand UO_871 (O_871,N_12813,N_12089);
or UO_872 (O_872,N_13874,N_14093);
and UO_873 (O_873,N_12667,N_13731);
or UO_874 (O_874,N_14618,N_14771);
or UO_875 (O_875,N_12871,N_13119);
and UO_876 (O_876,N_14638,N_12611);
and UO_877 (O_877,N_13101,N_13165);
nand UO_878 (O_878,N_12571,N_13478);
nand UO_879 (O_879,N_12990,N_14516);
nor UO_880 (O_880,N_12084,N_12627);
nor UO_881 (O_881,N_12390,N_14605);
or UO_882 (O_882,N_12221,N_14728);
nor UO_883 (O_883,N_12149,N_13169);
and UO_884 (O_884,N_13905,N_13909);
or UO_885 (O_885,N_12744,N_12510);
or UO_886 (O_886,N_12498,N_13992);
nand UO_887 (O_887,N_13358,N_14864);
and UO_888 (O_888,N_13942,N_14646);
nand UO_889 (O_889,N_14348,N_12907);
or UO_890 (O_890,N_13452,N_14233);
nand UO_891 (O_891,N_14536,N_14234);
and UO_892 (O_892,N_13422,N_13775);
xnor UO_893 (O_893,N_14702,N_12406);
or UO_894 (O_894,N_12689,N_13988);
or UO_895 (O_895,N_14268,N_14472);
or UO_896 (O_896,N_12527,N_13439);
nor UO_897 (O_897,N_13884,N_14481);
nor UO_898 (O_898,N_13917,N_13179);
nor UO_899 (O_899,N_12012,N_12515);
and UO_900 (O_900,N_13716,N_12063);
or UO_901 (O_901,N_14356,N_12414);
and UO_902 (O_902,N_13529,N_12439);
and UO_903 (O_903,N_12316,N_14978);
or UO_904 (O_904,N_12377,N_13843);
or UO_905 (O_905,N_14777,N_12996);
or UO_906 (O_906,N_12557,N_13637);
nor UO_907 (O_907,N_12111,N_14246);
and UO_908 (O_908,N_12992,N_14256);
nand UO_909 (O_909,N_12673,N_13097);
and UO_910 (O_910,N_14301,N_14548);
nand UO_911 (O_911,N_13103,N_12613);
nor UO_912 (O_912,N_13973,N_14517);
nor UO_913 (O_913,N_13647,N_12193);
and UO_914 (O_914,N_14651,N_14709);
or UO_915 (O_915,N_12066,N_14387);
or UO_916 (O_916,N_13614,N_14970);
or UO_917 (O_917,N_12585,N_13192);
and UO_918 (O_918,N_13482,N_13664);
and UO_919 (O_919,N_13916,N_12014);
and UO_920 (O_920,N_13755,N_13174);
nand UO_921 (O_921,N_14872,N_14466);
nand UO_922 (O_922,N_14297,N_13477);
nor UO_923 (O_923,N_13255,N_13829);
nand UO_924 (O_924,N_12924,N_14873);
nand UO_925 (O_925,N_14311,N_13256);
and UO_926 (O_926,N_14485,N_13292);
and UO_927 (O_927,N_13252,N_12348);
and UO_928 (O_928,N_14130,N_13425);
nor UO_929 (O_929,N_12657,N_14500);
xor UO_930 (O_930,N_13079,N_14274);
or UO_931 (O_931,N_12424,N_13989);
or UO_932 (O_932,N_13476,N_14895);
nor UO_933 (O_933,N_12287,N_14026);
nor UO_934 (O_934,N_14467,N_14518);
and UO_935 (O_935,N_13327,N_12130);
nor UO_936 (O_936,N_12590,N_13348);
nand UO_937 (O_937,N_14117,N_13007);
nand UO_938 (O_938,N_14150,N_14757);
or UO_939 (O_939,N_13373,N_14300);
and UO_940 (O_940,N_14766,N_12132);
nor UO_941 (O_941,N_12874,N_14380);
nand UO_942 (O_942,N_13228,N_14283);
nor UO_943 (O_943,N_14750,N_13306);
nor UO_944 (O_944,N_13199,N_13091);
nor UO_945 (O_945,N_13549,N_13844);
nand UO_946 (O_946,N_12271,N_13036);
nor UO_947 (O_947,N_13587,N_13688);
nor UO_948 (O_948,N_14972,N_14773);
nor UO_949 (O_949,N_13706,N_14172);
nor UO_950 (O_950,N_13689,N_14882);
xnor UO_951 (O_951,N_13216,N_12493);
or UO_952 (O_952,N_13730,N_12460);
or UO_953 (O_953,N_12734,N_12225);
and UO_954 (O_954,N_12352,N_12418);
and UO_955 (O_955,N_13593,N_13971);
nand UO_956 (O_956,N_13066,N_13686);
and UO_957 (O_957,N_14962,N_14943);
nor UO_958 (O_958,N_14637,N_13872);
nor UO_959 (O_959,N_12834,N_14532);
and UO_960 (O_960,N_12965,N_14058);
nor UO_961 (O_961,N_13582,N_12767);
and UO_962 (O_962,N_12762,N_12549);
nor UO_963 (O_963,N_14787,N_12796);
and UO_964 (O_964,N_13168,N_12857);
and UO_965 (O_965,N_14121,N_14935);
nand UO_966 (O_966,N_14625,N_13341);
nor UO_967 (O_967,N_12818,N_14533);
and UO_968 (O_968,N_12881,N_12276);
xnor UO_969 (O_969,N_14565,N_14132);
and UO_970 (O_970,N_12464,N_14176);
and UO_971 (O_971,N_12569,N_14793);
nor UO_972 (O_972,N_12937,N_12087);
nand UO_973 (O_973,N_12065,N_13602);
or UO_974 (O_974,N_13734,N_13283);
and UO_975 (O_975,N_14227,N_13060);
nand UO_976 (O_976,N_12435,N_13821);
xor UO_977 (O_977,N_12351,N_13344);
and UO_978 (O_978,N_12194,N_14693);
nand UO_979 (O_979,N_14369,N_12443);
nand UO_980 (O_980,N_14082,N_14050);
and UO_981 (O_981,N_14770,N_14510);
nand UO_982 (O_982,N_13564,N_13374);
nand UO_983 (O_983,N_14956,N_12253);
or UO_984 (O_984,N_12704,N_12696);
or UO_985 (O_985,N_12773,N_13590);
or UO_986 (O_986,N_12218,N_12070);
nand UO_987 (O_987,N_12452,N_13724);
or UO_988 (O_988,N_12616,N_14575);
nand UO_989 (O_989,N_13046,N_12841);
xor UO_990 (O_990,N_13742,N_12989);
and UO_991 (O_991,N_13014,N_14515);
or UO_992 (O_992,N_14586,N_12897);
or UO_993 (O_993,N_12573,N_13666);
or UO_994 (O_994,N_14261,N_14166);
xnor UO_995 (O_995,N_12238,N_14360);
or UO_996 (O_996,N_12819,N_12246);
nor UO_997 (O_997,N_12057,N_14494);
or UO_998 (O_998,N_12003,N_14318);
nand UO_999 (O_999,N_14428,N_12449);
nand UO_1000 (O_1000,N_14108,N_12572);
nor UO_1001 (O_1001,N_12916,N_13993);
or UO_1002 (O_1002,N_13118,N_12432);
nor UO_1003 (O_1003,N_14642,N_12783);
or UO_1004 (O_1004,N_14619,N_14394);
nor UO_1005 (O_1005,N_14271,N_12904);
and UO_1006 (O_1006,N_13842,N_14493);
and UO_1007 (O_1007,N_13483,N_12081);
and UO_1008 (O_1008,N_12815,N_13616);
or UO_1009 (O_1009,N_13063,N_14273);
xnor UO_1010 (O_1010,N_12960,N_14063);
or UO_1011 (O_1011,N_12198,N_14210);
nor UO_1012 (O_1012,N_12027,N_14607);
nand UO_1013 (O_1013,N_12389,N_12956);
nand UO_1014 (O_1014,N_14276,N_14290);
nand UO_1015 (O_1015,N_13575,N_14975);
and UO_1016 (O_1016,N_14919,N_14917);
and UO_1017 (O_1017,N_14275,N_13302);
or UO_1018 (O_1018,N_13935,N_14825);
nand UO_1019 (O_1019,N_14655,N_12181);
nor UO_1020 (O_1020,N_13679,N_14378);
nor UO_1021 (O_1021,N_12784,N_12661);
nand UO_1022 (O_1022,N_12577,N_14400);
nand UO_1023 (O_1023,N_14295,N_13831);
nand UO_1024 (O_1024,N_14138,N_12226);
xor UO_1025 (O_1025,N_14938,N_12828);
or UO_1026 (O_1026,N_13166,N_13223);
or UO_1027 (O_1027,N_14934,N_14584);
and UO_1028 (O_1028,N_14924,N_12062);
xnor UO_1029 (O_1029,N_14385,N_13639);
and UO_1030 (O_1030,N_14746,N_12853);
nand UO_1031 (O_1031,N_13628,N_14101);
or UO_1032 (O_1032,N_12731,N_13489);
nor UO_1033 (O_1033,N_12651,N_13961);
or UO_1034 (O_1034,N_13115,N_13932);
or UO_1035 (O_1035,N_13846,N_14572);
and UO_1036 (O_1036,N_12160,N_13511);
and UO_1037 (O_1037,N_14915,N_12757);
and UO_1038 (O_1038,N_12617,N_12488);
or UO_1039 (O_1039,N_13415,N_12563);
or UO_1040 (O_1040,N_13408,N_12190);
xor UO_1041 (O_1041,N_14666,N_13054);
or UO_1042 (O_1042,N_13670,N_12839);
nand UO_1043 (O_1043,N_13290,N_12883);
or UO_1044 (O_1044,N_12594,N_14547);
or UO_1045 (O_1045,N_12703,N_14901);
nand UO_1046 (O_1046,N_13601,N_12885);
nor UO_1047 (O_1047,N_13243,N_12166);
nand UO_1048 (O_1048,N_13673,N_13191);
nand UO_1049 (O_1049,N_14643,N_12209);
nor UO_1050 (O_1050,N_14459,N_13859);
nor UO_1051 (O_1051,N_14209,N_13654);
and UO_1052 (O_1052,N_13454,N_13224);
nor UO_1053 (O_1053,N_13170,N_13323);
xor UO_1054 (O_1054,N_12262,N_13705);
nand UO_1055 (O_1055,N_12105,N_12596);
or UO_1056 (O_1056,N_13381,N_14476);
and UO_1057 (O_1057,N_13161,N_13958);
nor UO_1058 (O_1058,N_13333,N_13534);
and UO_1059 (O_1059,N_14218,N_12384);
nor UO_1060 (O_1060,N_12212,N_12403);
nor UO_1061 (O_1061,N_14425,N_14534);
nor UO_1062 (O_1062,N_14269,N_13230);
or UO_1063 (O_1063,N_12267,N_13067);
or UO_1064 (O_1064,N_14676,N_13506);
nand UO_1065 (O_1065,N_12157,N_13316);
nand UO_1066 (O_1066,N_14350,N_13648);
and UO_1067 (O_1067,N_13085,N_14135);
and UO_1068 (O_1068,N_13008,N_12031);
xor UO_1069 (O_1069,N_14463,N_13798);
and UO_1070 (O_1070,N_12713,N_14567);
nand UO_1071 (O_1071,N_14195,N_12483);
and UO_1072 (O_1072,N_12013,N_12553);
and UO_1073 (O_1073,N_12178,N_14509);
nand UO_1074 (O_1074,N_13856,N_13441);
and UO_1075 (O_1075,N_13464,N_14898);
or UO_1076 (O_1076,N_12952,N_13901);
and UO_1077 (O_1077,N_13037,N_13263);
or UO_1078 (O_1078,N_13459,N_13956);
and UO_1079 (O_1079,N_13930,N_14432);
nand UO_1080 (O_1080,N_14855,N_14891);
and UO_1081 (O_1081,N_14189,N_13643);
nand UO_1082 (O_1082,N_12242,N_14983);
and UO_1083 (O_1083,N_12165,N_12101);
nand UO_1084 (O_1084,N_14401,N_13366);
or UO_1085 (O_1085,N_12772,N_12356);
nand UO_1086 (O_1086,N_13788,N_14576);
xor UO_1087 (O_1087,N_14253,N_14188);
and UO_1088 (O_1088,N_14281,N_14074);
nor UO_1089 (O_1089,N_12811,N_13410);
nand UO_1090 (O_1090,N_13480,N_14817);
nand UO_1091 (O_1091,N_12555,N_14670);
nand UO_1092 (O_1092,N_14546,N_14241);
nand UO_1093 (O_1093,N_13808,N_14125);
nor UO_1094 (O_1094,N_14075,N_12822);
or UO_1095 (O_1095,N_13644,N_14942);
and UO_1096 (O_1096,N_13336,N_12672);
or UO_1097 (O_1097,N_13881,N_12764);
nand UO_1098 (O_1098,N_12431,N_13331);
and UO_1099 (O_1099,N_13027,N_14289);
nand UO_1100 (O_1100,N_14909,N_12748);
or UO_1101 (O_1101,N_12934,N_13745);
and UO_1102 (O_1102,N_13497,N_13503);
nand UO_1103 (O_1103,N_13665,N_13984);
nor UO_1104 (O_1104,N_14870,N_14070);
nor UO_1105 (O_1105,N_13164,N_12484);
nand UO_1106 (O_1106,N_12534,N_13340);
nand UO_1107 (O_1107,N_14021,N_12724);
and UO_1108 (O_1108,N_12502,N_14354);
nand UO_1109 (O_1109,N_14266,N_13500);
and UO_1110 (O_1110,N_13420,N_14329);
nand UO_1111 (O_1111,N_12164,N_13597);
nand UO_1112 (O_1112,N_12507,N_12158);
or UO_1113 (O_1113,N_12949,N_14786);
and UO_1114 (O_1114,N_14738,N_13093);
or UO_1115 (O_1115,N_12869,N_12971);
xor UO_1116 (O_1116,N_14399,N_13055);
or UO_1117 (O_1117,N_14148,N_13924);
and UO_1118 (O_1118,N_13661,N_12809);
nand UO_1119 (O_1119,N_12137,N_12268);
nor UO_1120 (O_1120,N_12824,N_12694);
nor UO_1121 (O_1121,N_12354,N_13137);
nor UO_1122 (O_1122,N_14391,N_13566);
nor UO_1123 (O_1123,N_14553,N_12780);
and UO_1124 (O_1124,N_12465,N_12341);
and UO_1125 (O_1125,N_13768,N_12275);
nand UO_1126 (O_1126,N_14032,N_12292);
nand UO_1127 (O_1127,N_13058,N_13396);
nand UO_1128 (O_1128,N_13612,N_12135);
nand UO_1129 (O_1129,N_14445,N_12299);
or UO_1130 (O_1130,N_12408,N_13401);
nor UO_1131 (O_1131,N_14744,N_13038);
and UO_1132 (O_1132,N_14514,N_12289);
or UO_1133 (O_1133,N_12118,N_14386);
nand UO_1134 (O_1134,N_13488,N_14524);
nand UO_1135 (O_1135,N_13025,N_12059);
nor UO_1136 (O_1136,N_14854,N_12546);
nor UO_1137 (O_1137,N_12600,N_12448);
nor UO_1138 (O_1138,N_13518,N_14948);
nor UO_1139 (O_1139,N_13207,N_12233);
and UO_1140 (O_1140,N_12759,N_12678);
or UO_1141 (O_1141,N_12697,N_14561);
and UO_1142 (O_1142,N_13434,N_12147);
or UO_1143 (O_1143,N_14216,N_13711);
nor UO_1144 (O_1144,N_14072,N_14508);
and UO_1145 (O_1145,N_13082,N_12489);
nand UO_1146 (O_1146,N_13367,N_12642);
nor UO_1147 (O_1147,N_13784,N_14012);
and UO_1148 (O_1148,N_12597,N_13308);
nor UO_1149 (O_1149,N_12257,N_14703);
or UO_1150 (O_1150,N_13108,N_14245);
nor UO_1151 (O_1151,N_14161,N_14963);
nor UO_1152 (O_1152,N_13982,N_13589);
or UO_1153 (O_1153,N_14940,N_14877);
or UO_1154 (O_1154,N_13544,N_12663);
or UO_1155 (O_1155,N_14199,N_14836);
and UO_1156 (O_1156,N_13321,N_12425);
or UO_1157 (O_1157,N_12751,N_14653);
nor UO_1158 (O_1158,N_14005,N_14129);
nor UO_1159 (O_1159,N_12416,N_13588);
nor UO_1160 (O_1160,N_13657,N_13709);
nor UO_1161 (O_1161,N_14779,N_12015);
nor UO_1162 (O_1162,N_13435,N_13650);
and UO_1163 (O_1163,N_13675,N_13275);
and UO_1164 (O_1164,N_13417,N_14874);
nor UO_1165 (O_1165,N_14367,N_13792);
or UO_1166 (O_1166,N_14920,N_13369);
nor UO_1167 (O_1167,N_12605,N_13862);
or UO_1168 (O_1168,N_14351,N_13817);
or UO_1169 (O_1169,N_14539,N_14585);
nand UO_1170 (O_1170,N_14632,N_14861);
or UO_1171 (O_1171,N_13131,N_13264);
and UO_1172 (O_1172,N_14776,N_13226);
nor UO_1173 (O_1173,N_12975,N_12475);
nand UO_1174 (O_1174,N_12099,N_13586);
nor UO_1175 (O_1175,N_13000,N_14015);
or UO_1176 (O_1176,N_12184,N_13455);
or UO_1177 (O_1177,N_13320,N_13983);
nand UO_1178 (O_1178,N_13504,N_14134);
or UO_1179 (O_1179,N_12709,N_14080);
nor UO_1180 (O_1180,N_13314,N_13088);
or UO_1181 (O_1181,N_14492,N_13998);
nor UO_1182 (O_1182,N_12802,N_12229);
or UO_1183 (O_1183,N_13803,N_12628);
xnor UO_1184 (O_1184,N_12019,N_14244);
nor UO_1185 (O_1185,N_14903,N_12732);
nor UO_1186 (O_1186,N_12726,N_12997);
and UO_1187 (O_1187,N_14862,N_12254);
nor UO_1188 (O_1188,N_14800,N_12244);
or UO_1189 (O_1189,N_14170,N_12629);
nand UO_1190 (O_1190,N_12168,N_12107);
or UO_1191 (O_1191,N_14504,N_12929);
or UO_1192 (O_1192,N_13985,N_14828);
or UO_1193 (O_1193,N_14303,N_12011);
nor UO_1194 (O_1194,N_14486,N_12712);
nor UO_1195 (O_1195,N_13574,N_14461);
and UO_1196 (O_1196,N_14337,N_12196);
nand UO_1197 (O_1197,N_14168,N_13107);
nand UO_1198 (O_1198,N_14628,N_12902);
nand UO_1199 (O_1199,N_14184,N_12905);
nor UO_1200 (O_1200,N_14320,N_13902);
or UO_1201 (O_1201,N_13342,N_14679);
or UO_1202 (O_1202,N_14462,N_12915);
and UO_1203 (O_1203,N_14928,N_12076);
nand UO_1204 (O_1204,N_14100,N_14024);
nand UO_1205 (O_1205,N_13402,N_14803);
nand UO_1206 (O_1206,N_12114,N_13451);
and UO_1207 (O_1207,N_14858,N_13533);
nand UO_1208 (O_1208,N_13300,N_14212);
nand UO_1209 (O_1209,N_14714,N_13188);
xnor UO_1210 (O_1210,N_14035,N_14739);
nand UO_1211 (O_1211,N_13815,N_12785);
and UO_1212 (O_1212,N_13440,N_12402);
nor UO_1213 (O_1213,N_12860,N_13759);
nand UO_1214 (O_1214,N_12863,N_12920);
and UO_1215 (O_1215,N_14055,N_12466);
or UO_1216 (O_1216,N_13830,N_12037);
nor UO_1217 (O_1217,N_12621,N_12129);
nor UO_1218 (O_1218,N_12385,N_12282);
or UO_1219 (O_1219,N_13837,N_12409);
or UO_1220 (O_1220,N_14512,N_14317);
nor UO_1221 (O_1221,N_14390,N_12186);
or UO_1222 (O_1222,N_14937,N_14603);
nor UO_1223 (O_1223,N_12758,N_12926);
or UO_1224 (O_1224,N_12175,N_14412);
nor UO_1225 (O_1225,N_14747,N_12182);
or UO_1226 (O_1226,N_12545,N_12091);
or UO_1227 (O_1227,N_13740,N_12552);
nand UO_1228 (O_1228,N_13695,N_12836);
nand UO_1229 (O_1229,N_13023,N_13565);
nor UO_1230 (O_1230,N_14031,N_14226);
nand UO_1231 (O_1231,N_13980,N_13315);
nand UO_1232 (O_1232,N_12146,N_12955);
and UO_1233 (O_1233,N_14865,N_12593);
and UO_1234 (O_1234,N_13542,N_13409);
and UO_1235 (O_1235,N_14473,N_13749);
or UO_1236 (O_1236,N_14569,N_12145);
nor UO_1237 (O_1237,N_12434,N_14053);
nor UO_1238 (O_1238,N_14345,N_13551);
xnor UO_1239 (O_1239,N_14179,N_12923);
nand UO_1240 (O_1240,N_12428,N_12321);
nor UO_1241 (O_1241,N_13121,N_14959);
nand UO_1242 (O_1242,N_13239,N_13160);
xnor UO_1243 (O_1243,N_12161,N_14527);
and UO_1244 (O_1244,N_12602,N_12636);
or UO_1245 (O_1245,N_13765,N_13921);
nor UO_1246 (O_1246,N_12140,N_13303);
nor UO_1247 (O_1247,N_12533,N_12951);
nand UO_1248 (O_1248,N_13279,N_14578);
or UO_1249 (O_1249,N_13114,N_13162);
and UO_1250 (O_1250,N_14907,N_14200);
and UO_1251 (O_1251,N_14680,N_12369);
or UO_1252 (O_1252,N_14262,N_14410);
nor UO_1253 (O_1253,N_12296,N_12319);
nor UO_1254 (O_1254,N_13685,N_14944);
and UO_1255 (O_1255,N_12104,N_13866);
and UO_1256 (O_1256,N_14405,N_13406);
nor UO_1257 (O_1257,N_13349,N_13392);
nand UO_1258 (O_1258,N_14128,N_13042);
nor UO_1259 (O_1259,N_14115,N_14257);
or UO_1260 (O_1260,N_12103,N_12404);
nand UO_1261 (O_1261,N_13569,N_14040);
or UO_1262 (O_1262,N_14574,N_14513);
or UO_1263 (O_1263,N_12154,N_14243);
and UO_1264 (O_1264,N_12162,N_13883);
nand UO_1265 (O_1265,N_12249,N_12092);
xor UO_1266 (O_1266,N_14531,N_13558);
and UO_1267 (O_1267,N_12991,N_14224);
nand UO_1268 (O_1268,N_14664,N_14636);
or UO_1269 (O_1269,N_12995,N_14232);
nor UO_1270 (O_1270,N_13920,N_14229);
or UO_1271 (O_1271,N_13845,N_12677);
nor UO_1272 (O_1272,N_12366,N_12142);
nand UO_1273 (O_1273,N_13579,N_13399);
and UO_1274 (O_1274,N_13145,N_13767);
nand UO_1275 (O_1275,N_13869,N_12714);
and UO_1276 (O_1276,N_14594,N_14863);
or UO_1277 (O_1277,N_12671,N_14223);
nor UO_1278 (O_1278,N_14322,N_14001);
and UO_1279 (O_1279,N_12914,N_12391);
or UO_1280 (O_1280,N_13246,N_14406);
nor UO_1281 (O_1281,N_12913,N_14475);
xnor UO_1282 (O_1282,N_13680,N_14083);
or UO_1283 (O_1283,N_12637,N_14902);
and UO_1284 (O_1284,N_12359,N_12730);
nor UO_1285 (O_1285,N_14525,N_13886);
nand UO_1286 (O_1286,N_12576,N_12476);
and UO_1287 (O_1287,N_12326,N_12930);
nand UO_1288 (O_1288,N_13827,N_14735);
and UO_1289 (O_1289,N_12381,N_13605);
and UO_1290 (O_1290,N_14985,N_12125);
or UO_1291 (O_1291,N_12523,N_13996);
nand UO_1292 (O_1292,N_14784,N_14674);
xor UO_1293 (O_1293,N_14187,N_13576);
and UO_1294 (O_1294,N_14630,N_14424);
or UO_1295 (O_1295,N_14749,N_13202);
and UO_1296 (O_1296,N_14764,N_14733);
nor UO_1297 (O_1297,N_12501,N_14167);
nand UO_1298 (O_1298,N_12023,N_14911);
or UO_1299 (O_1299,N_13271,N_13421);
and UO_1300 (O_1300,N_12812,N_14372);
and UO_1301 (O_1301,N_14455,N_12984);
xor UO_1302 (O_1302,N_13502,N_14598);
and UO_1303 (O_1303,N_12779,N_14573);
or UO_1304 (O_1304,N_12935,N_14313);
nor UO_1305 (O_1305,N_14795,N_12842);
or UO_1306 (O_1306,N_14840,N_14823);
and UO_1307 (O_1307,N_12669,N_12462);
xnor UO_1308 (O_1308,N_14013,N_14683);
or UO_1309 (O_1309,N_13515,N_14819);
or UO_1310 (O_1310,N_14627,N_13222);
nand UO_1311 (O_1311,N_13184,N_13479);
nor UO_1312 (O_1312,N_14418,N_12223);
and UO_1313 (O_1313,N_12958,N_14092);
and UO_1314 (O_1314,N_14648,N_12631);
or UO_1315 (O_1315,N_14443,N_13423);
xor UO_1316 (O_1316,N_13189,N_13577);
nand UO_1317 (O_1317,N_13548,N_13377);
nor UO_1318 (O_1318,N_13708,N_14743);
nand UO_1319 (O_1319,N_12528,N_12090);
or UO_1320 (O_1320,N_14335,N_14842);
and UO_1321 (O_1321,N_14644,N_12252);
and UO_1322 (O_1322,N_12544,N_12112);
and UO_1323 (O_1323,N_14964,N_14292);
nor UO_1324 (O_1324,N_14867,N_14685);
nor UO_1325 (O_1325,N_12797,N_13633);
xor UO_1326 (O_1326,N_12230,N_14365);
nand UO_1327 (O_1327,N_13247,N_13739);
nand UO_1328 (O_1328,N_14263,N_13183);
nand UO_1329 (O_1329,N_12036,N_13986);
nand UO_1330 (O_1330,N_14829,N_13013);
nor UO_1331 (O_1331,N_12303,N_12270);
nor UO_1332 (O_1332,N_14119,N_12526);
nand UO_1333 (O_1333,N_14835,N_13904);
and UO_1334 (O_1334,N_12446,N_14383);
and UO_1335 (O_1335,N_12665,N_14635);
nor UO_1336 (O_1336,N_12265,N_14820);
nor UO_1337 (O_1337,N_13923,N_13651);
nand UO_1338 (O_1338,N_12018,N_14761);
and UO_1339 (O_1339,N_13911,N_13719);
nor UO_1340 (O_1340,N_14307,N_13372);
nand UO_1341 (O_1341,N_14427,N_13407);
and UO_1342 (O_1342,N_14697,N_13475);
or UO_1343 (O_1343,N_14451,N_13266);
or UO_1344 (O_1344,N_12096,N_12880);
or UO_1345 (O_1345,N_12833,N_14440);
and UO_1346 (O_1346,N_12868,N_13313);
nor UO_1347 (O_1347,N_13432,N_14980);
or UO_1348 (O_1348,N_13413,N_12805);
nand UO_1349 (O_1349,N_13770,N_14457);
nand UO_1350 (O_1350,N_13443,N_13513);
nor UO_1351 (O_1351,N_12919,N_12910);
and UO_1352 (O_1352,N_12358,N_12889);
nand UO_1353 (O_1353,N_13826,N_13771);
and UO_1354 (O_1354,N_12674,N_14563);
or UO_1355 (O_1355,N_13540,N_13764);
nor UO_1356 (O_1356,N_13268,N_14551);
nor UO_1357 (O_1357,N_12367,N_13584);
or UO_1358 (O_1358,N_14526,N_12017);
or UO_1359 (O_1359,N_12115,N_13102);
xor UO_1360 (O_1360,N_12781,N_12849);
nand UO_1361 (O_1361,N_14848,N_13936);
and UO_1362 (O_1362,N_12058,N_12551);
or UO_1363 (O_1363,N_13288,N_13178);
nor UO_1364 (O_1364,N_13135,N_12082);
nand UO_1365 (O_1365,N_13863,N_14994);
nor UO_1366 (O_1366,N_13718,N_13075);
and UO_1367 (O_1367,N_14336,N_12281);
or UO_1368 (O_1368,N_14008,N_14969);
and UO_1369 (O_1369,N_13914,N_14765);
nand UO_1370 (O_1370,N_12134,N_14615);
or UO_1371 (O_1371,N_14278,N_14302);
xnor UO_1372 (O_1372,N_13043,N_12038);
or UO_1373 (O_1373,N_12041,N_12550);
nand UO_1374 (O_1374,N_14740,N_13487);
nand UO_1375 (O_1375,N_13442,N_14726);
nand UO_1376 (O_1376,N_12978,N_12236);
or UO_1377 (O_1377,N_13625,N_13773);
nand UO_1378 (O_1378,N_13816,N_14315);
nor UO_1379 (O_1379,N_13404,N_14724);
nand UO_1380 (O_1380,N_14151,N_13766);
or UO_1381 (O_1381,N_14211,N_14192);
nor UO_1382 (O_1382,N_14925,N_12382);
nand UO_1383 (O_1383,N_13852,N_14502);
nor UO_1384 (O_1384,N_12794,N_12100);
or UO_1385 (O_1385,N_13468,N_13505);
or UO_1386 (O_1386,N_14804,N_13065);
or UO_1387 (O_1387,N_12831,N_13854);
nor UO_1388 (O_1388,N_14866,N_14145);
nor UO_1389 (O_1389,N_12729,N_12514);
nor UO_1390 (O_1390,N_13032,N_14688);
xnor UO_1391 (O_1391,N_12791,N_13877);
nor UO_1392 (O_1392,N_12127,N_12411);
nand UO_1393 (O_1393,N_12721,N_12900);
nand UO_1394 (O_1394,N_13890,N_13838);
and UO_1395 (O_1395,N_12346,N_13047);
nand UO_1396 (O_1396,N_12614,N_13748);
and UO_1397 (O_1397,N_14061,N_12876);
nand UO_1398 (O_1398,N_14368,N_13329);
or UO_1399 (O_1399,N_13338,N_13311);
nor UO_1400 (O_1400,N_12723,N_12765);
nor UO_1401 (O_1401,N_12543,N_14374);
nor UO_1402 (O_1402,N_12509,N_14447);
xor UO_1403 (O_1403,N_14444,N_12692);
or UO_1404 (O_1404,N_14957,N_13987);
nand UO_1405 (O_1405,N_13780,N_14657);
nand UO_1406 (O_1406,N_13029,N_13624);
nor UO_1407 (O_1407,N_13604,N_13741);
nor UO_1408 (O_1408,N_14006,N_13144);
and UO_1409 (O_1409,N_12847,N_13448);
nor UO_1410 (O_1410,N_12566,N_12288);
nand UO_1411 (O_1411,N_12901,N_14692);
nand UO_1412 (O_1412,N_14116,N_14458);
nand UO_1413 (O_1413,N_12320,N_14194);
or UO_1414 (O_1414,N_13465,N_13274);
and UO_1415 (O_1415,N_13050,N_14123);
nor UO_1416 (O_1416,N_13267,N_13699);
and UO_1417 (O_1417,N_12749,N_14748);
xnor UO_1418 (O_1418,N_13437,N_14826);
and UO_1419 (O_1419,N_14185,N_14806);
nand UO_1420 (O_1420,N_12330,N_14104);
nor UO_1421 (O_1421,N_12525,N_12708);
nand UO_1422 (O_1422,N_14488,N_13276);
or UO_1423 (O_1423,N_13104,N_14420);
or UO_1424 (O_1424,N_14616,N_14562);
nor UO_1425 (O_1425,N_12468,N_13361);
or UO_1426 (O_1426,N_14596,N_14878);
nor UO_1427 (O_1427,N_14422,N_13570);
nand UO_1428 (O_1428,N_14581,N_14207);
and UO_1429 (O_1429,N_13704,N_14552);
nor UO_1430 (O_1430,N_12119,N_12699);
xor UO_1431 (O_1431,N_14694,N_12247);
and UO_1432 (O_1432,N_12967,N_14046);
or UO_1433 (O_1433,N_12333,N_12026);
or UO_1434 (O_1434,N_14762,N_12579);
xor UO_1435 (O_1435,N_12504,N_14022);
xor UO_1436 (O_1436,N_12795,N_12053);
and UO_1437 (O_1437,N_13148,N_13618);
nor UO_1438 (O_1438,N_12050,N_14306);
nand UO_1439 (O_1439,N_14912,N_12300);
or UO_1440 (O_1440,N_14449,N_13272);
or UO_1441 (O_1441,N_13541,N_13017);
xnor UO_1442 (O_1442,N_12656,N_13608);
or UO_1443 (O_1443,N_14039,N_14808);
nand UO_1444 (O_1444,N_14577,N_14413);
nor UO_1445 (O_1445,N_14889,N_14044);
nand UO_1446 (O_1446,N_14897,N_12482);
nor UO_1447 (O_1447,N_14204,N_14429);
nor UO_1448 (O_1448,N_14010,N_14025);
or UO_1449 (O_1449,N_14852,N_14328);
and UO_1450 (O_1450,N_13915,N_13190);
nor UO_1451 (O_1451,N_14537,N_12120);
or UO_1452 (O_1452,N_13172,N_13939);
xnor UO_1453 (O_1453,N_12258,N_12386);
nor UO_1454 (O_1454,N_12095,N_12890);
and UO_1455 (O_1455,N_12986,N_13398);
or UO_1456 (O_1456,N_12953,N_12583);
nor UO_1457 (O_1457,N_14698,N_14126);
or UO_1458 (O_1458,N_12170,N_14242);
and UO_1459 (O_1459,N_12413,N_13607);
or UO_1460 (O_1460,N_13236,N_12532);
and UO_1461 (O_1461,N_12376,N_12887);
nor UO_1462 (O_1462,N_13062,N_13907);
nor UO_1463 (O_1463,N_12655,N_14530);
nor UO_1464 (O_1464,N_14423,N_12169);
nor UO_1465 (O_1465,N_13698,N_13557);
nor UO_1466 (O_1466,N_12940,N_12850);
and UO_1467 (O_1467,N_12072,N_13030);
nor UO_1468 (O_1468,N_12331,N_12248);
and UO_1469 (O_1469,N_12187,N_12152);
nand UO_1470 (O_1470,N_14002,N_13485);
and UO_1471 (O_1471,N_14016,N_13912);
xnor UO_1472 (O_1472,N_13509,N_13159);
nor UO_1473 (O_1473,N_14571,N_12235);
nand UO_1474 (O_1474,N_12559,N_12400);
nor UO_1475 (O_1475,N_13931,N_14580);
nor UO_1476 (O_1476,N_14521,N_14813);
and UO_1477 (O_1477,N_12294,N_13411);
nor UO_1478 (O_1478,N_13824,N_12328);
nand UO_1479 (O_1479,N_14841,N_14797);
nand UO_1480 (O_1480,N_13087,N_12396);
or UO_1481 (O_1481,N_13757,N_12060);
and UO_1482 (O_1482,N_14772,N_12153);
nand UO_1483 (O_1483,N_13662,N_12219);
and UO_1484 (O_1484,N_13634,N_14945);
nand UO_1485 (O_1485,N_13084,N_13823);
nand UO_1486 (O_1486,N_12964,N_12630);
or UO_1487 (O_1487,N_13727,N_12707);
nand UO_1488 (O_1488,N_14397,N_14805);
nand UO_1489 (O_1489,N_12335,N_14178);
nor UO_1490 (O_1490,N_14358,N_13512);
and UO_1491 (O_1491,N_14754,N_14240);
nand UO_1492 (O_1492,N_13241,N_12867);
and UO_1493 (O_1493,N_13977,N_13972);
or UO_1494 (O_1494,N_13591,N_13761);
nor UO_1495 (O_1495,N_14752,N_12968);
and UO_1496 (O_1496,N_13899,N_12943);
nor UO_1497 (O_1497,N_12313,N_14958);
nand UO_1498 (O_1498,N_12126,N_12042);
xnor UO_1499 (O_1499,N_13818,N_14395);
nand UO_1500 (O_1500,N_13631,N_12497);
or UO_1501 (O_1501,N_14057,N_14069);
nand UO_1502 (O_1502,N_12210,N_14462);
nor UO_1503 (O_1503,N_14549,N_12918);
nand UO_1504 (O_1504,N_13838,N_13174);
or UO_1505 (O_1505,N_14156,N_14961);
nand UO_1506 (O_1506,N_14379,N_14746);
or UO_1507 (O_1507,N_14131,N_13169);
nand UO_1508 (O_1508,N_13764,N_13687);
nor UO_1509 (O_1509,N_14010,N_14540);
or UO_1510 (O_1510,N_14884,N_12350);
nand UO_1511 (O_1511,N_14207,N_14255);
nor UO_1512 (O_1512,N_14257,N_14870);
nor UO_1513 (O_1513,N_12095,N_13002);
nand UO_1514 (O_1514,N_14057,N_12492);
nor UO_1515 (O_1515,N_14869,N_14722);
and UO_1516 (O_1516,N_12846,N_14936);
nor UO_1517 (O_1517,N_13024,N_14683);
xnor UO_1518 (O_1518,N_13572,N_13317);
xnor UO_1519 (O_1519,N_12784,N_12576);
or UO_1520 (O_1520,N_12405,N_13426);
or UO_1521 (O_1521,N_14724,N_13067);
and UO_1522 (O_1522,N_13953,N_12960);
nand UO_1523 (O_1523,N_13860,N_14557);
nand UO_1524 (O_1524,N_12407,N_14935);
xor UO_1525 (O_1525,N_13846,N_14436);
and UO_1526 (O_1526,N_14502,N_13434);
or UO_1527 (O_1527,N_12899,N_14761);
and UO_1528 (O_1528,N_13202,N_14502);
nor UO_1529 (O_1529,N_13765,N_13125);
or UO_1530 (O_1530,N_13781,N_12057);
nand UO_1531 (O_1531,N_14781,N_12935);
xor UO_1532 (O_1532,N_14335,N_14243);
nor UO_1533 (O_1533,N_14830,N_14207);
nor UO_1534 (O_1534,N_12216,N_13605);
and UO_1535 (O_1535,N_13868,N_12417);
or UO_1536 (O_1536,N_13136,N_14692);
nor UO_1537 (O_1537,N_13545,N_12775);
nand UO_1538 (O_1538,N_14650,N_12167);
or UO_1539 (O_1539,N_13803,N_13150);
nor UO_1540 (O_1540,N_12615,N_12226);
or UO_1541 (O_1541,N_14197,N_12891);
and UO_1542 (O_1542,N_14680,N_12491);
nand UO_1543 (O_1543,N_12291,N_14999);
nand UO_1544 (O_1544,N_12313,N_14375);
nor UO_1545 (O_1545,N_13273,N_12428);
nand UO_1546 (O_1546,N_14690,N_12270);
nor UO_1547 (O_1547,N_14402,N_13653);
xnor UO_1548 (O_1548,N_14907,N_14148);
nor UO_1549 (O_1549,N_14293,N_14659);
or UO_1550 (O_1550,N_14650,N_12013);
nand UO_1551 (O_1551,N_13820,N_12128);
xnor UO_1552 (O_1552,N_13837,N_12024);
and UO_1553 (O_1553,N_14854,N_12701);
nor UO_1554 (O_1554,N_12308,N_12164);
nand UO_1555 (O_1555,N_14313,N_14843);
nor UO_1556 (O_1556,N_12722,N_12355);
and UO_1557 (O_1557,N_14553,N_13606);
xnor UO_1558 (O_1558,N_14453,N_13806);
nor UO_1559 (O_1559,N_12505,N_12836);
nor UO_1560 (O_1560,N_13009,N_14174);
or UO_1561 (O_1561,N_14063,N_12830);
nand UO_1562 (O_1562,N_13188,N_12456);
nor UO_1563 (O_1563,N_12450,N_14495);
xnor UO_1564 (O_1564,N_13393,N_12604);
nand UO_1565 (O_1565,N_13838,N_12211);
and UO_1566 (O_1566,N_13022,N_12113);
or UO_1567 (O_1567,N_13943,N_13849);
nor UO_1568 (O_1568,N_13094,N_13848);
or UO_1569 (O_1569,N_12269,N_13193);
and UO_1570 (O_1570,N_13365,N_14837);
xnor UO_1571 (O_1571,N_13142,N_14005);
nor UO_1572 (O_1572,N_13521,N_12222);
or UO_1573 (O_1573,N_12604,N_14264);
or UO_1574 (O_1574,N_14614,N_13155);
xnor UO_1575 (O_1575,N_14974,N_13363);
xnor UO_1576 (O_1576,N_13880,N_14842);
and UO_1577 (O_1577,N_14359,N_12250);
or UO_1578 (O_1578,N_13413,N_14626);
nand UO_1579 (O_1579,N_14055,N_12314);
and UO_1580 (O_1580,N_13103,N_13100);
nand UO_1581 (O_1581,N_12938,N_12054);
and UO_1582 (O_1582,N_13700,N_12462);
and UO_1583 (O_1583,N_14568,N_14067);
or UO_1584 (O_1584,N_12425,N_12013);
nor UO_1585 (O_1585,N_13890,N_14994);
and UO_1586 (O_1586,N_12939,N_13222);
or UO_1587 (O_1587,N_13835,N_12997);
nand UO_1588 (O_1588,N_13835,N_13068);
nor UO_1589 (O_1589,N_14600,N_14193);
xnor UO_1590 (O_1590,N_14390,N_12197);
or UO_1591 (O_1591,N_13923,N_13536);
nand UO_1592 (O_1592,N_14168,N_14985);
and UO_1593 (O_1593,N_13845,N_12640);
or UO_1594 (O_1594,N_14787,N_13202);
nand UO_1595 (O_1595,N_14450,N_12909);
and UO_1596 (O_1596,N_12648,N_14055);
or UO_1597 (O_1597,N_14781,N_13736);
nand UO_1598 (O_1598,N_13225,N_13343);
nor UO_1599 (O_1599,N_13662,N_12604);
and UO_1600 (O_1600,N_14080,N_14874);
and UO_1601 (O_1601,N_13670,N_14409);
nor UO_1602 (O_1602,N_14183,N_14625);
xor UO_1603 (O_1603,N_12033,N_14137);
nor UO_1604 (O_1604,N_14291,N_13107);
nand UO_1605 (O_1605,N_13194,N_13258);
nor UO_1606 (O_1606,N_13120,N_12335);
nor UO_1607 (O_1607,N_13811,N_14254);
and UO_1608 (O_1608,N_14351,N_13597);
and UO_1609 (O_1609,N_13364,N_13917);
nand UO_1610 (O_1610,N_12967,N_12517);
and UO_1611 (O_1611,N_13267,N_12388);
and UO_1612 (O_1612,N_12466,N_12229);
nand UO_1613 (O_1613,N_12817,N_12201);
or UO_1614 (O_1614,N_13784,N_13838);
or UO_1615 (O_1615,N_12328,N_14191);
nand UO_1616 (O_1616,N_12715,N_12912);
nand UO_1617 (O_1617,N_13587,N_13755);
or UO_1618 (O_1618,N_12139,N_12988);
nand UO_1619 (O_1619,N_14571,N_12529);
nor UO_1620 (O_1620,N_14476,N_12466);
nor UO_1621 (O_1621,N_14673,N_12987);
or UO_1622 (O_1622,N_14028,N_13488);
and UO_1623 (O_1623,N_14717,N_12755);
xnor UO_1624 (O_1624,N_13727,N_14901);
and UO_1625 (O_1625,N_12889,N_12891);
nor UO_1626 (O_1626,N_12619,N_14794);
or UO_1627 (O_1627,N_14290,N_13787);
nor UO_1628 (O_1628,N_14323,N_12464);
and UO_1629 (O_1629,N_12693,N_12784);
nor UO_1630 (O_1630,N_12325,N_12258);
and UO_1631 (O_1631,N_13255,N_12772);
and UO_1632 (O_1632,N_14238,N_12817);
and UO_1633 (O_1633,N_12563,N_12302);
or UO_1634 (O_1634,N_12585,N_13151);
or UO_1635 (O_1635,N_12518,N_13475);
xnor UO_1636 (O_1636,N_12731,N_12169);
nand UO_1637 (O_1637,N_12530,N_14361);
or UO_1638 (O_1638,N_13533,N_13403);
xor UO_1639 (O_1639,N_13176,N_12929);
nand UO_1640 (O_1640,N_13379,N_12602);
xor UO_1641 (O_1641,N_14359,N_13787);
or UO_1642 (O_1642,N_14616,N_12873);
and UO_1643 (O_1643,N_14101,N_14290);
nor UO_1644 (O_1644,N_13560,N_13320);
and UO_1645 (O_1645,N_13370,N_14908);
and UO_1646 (O_1646,N_14920,N_13939);
nand UO_1647 (O_1647,N_12417,N_14540);
nor UO_1648 (O_1648,N_13505,N_12284);
and UO_1649 (O_1649,N_13507,N_13799);
nand UO_1650 (O_1650,N_13969,N_14514);
or UO_1651 (O_1651,N_12538,N_13217);
and UO_1652 (O_1652,N_14153,N_14775);
and UO_1653 (O_1653,N_12058,N_13914);
nor UO_1654 (O_1654,N_12302,N_13153);
nor UO_1655 (O_1655,N_12564,N_12839);
and UO_1656 (O_1656,N_12777,N_14004);
nor UO_1657 (O_1657,N_12311,N_14418);
or UO_1658 (O_1658,N_14119,N_13232);
or UO_1659 (O_1659,N_12934,N_13973);
nor UO_1660 (O_1660,N_13094,N_14067);
and UO_1661 (O_1661,N_14335,N_13580);
nor UO_1662 (O_1662,N_13450,N_12466);
and UO_1663 (O_1663,N_12537,N_13133);
or UO_1664 (O_1664,N_14824,N_13074);
nand UO_1665 (O_1665,N_13048,N_14544);
or UO_1666 (O_1666,N_14246,N_13915);
nor UO_1667 (O_1667,N_12105,N_14878);
or UO_1668 (O_1668,N_13827,N_12535);
nand UO_1669 (O_1669,N_12804,N_12750);
or UO_1670 (O_1670,N_13636,N_13872);
nand UO_1671 (O_1671,N_13462,N_14600);
or UO_1672 (O_1672,N_13783,N_12404);
nor UO_1673 (O_1673,N_14016,N_14554);
xor UO_1674 (O_1674,N_13108,N_12016);
or UO_1675 (O_1675,N_13195,N_12528);
or UO_1676 (O_1676,N_13150,N_14206);
nor UO_1677 (O_1677,N_12341,N_13560);
or UO_1678 (O_1678,N_14135,N_12763);
and UO_1679 (O_1679,N_12421,N_14717);
or UO_1680 (O_1680,N_12185,N_14379);
and UO_1681 (O_1681,N_12446,N_12194);
or UO_1682 (O_1682,N_12336,N_14816);
and UO_1683 (O_1683,N_13639,N_13057);
nor UO_1684 (O_1684,N_12721,N_14822);
nor UO_1685 (O_1685,N_14070,N_13897);
or UO_1686 (O_1686,N_12748,N_12568);
nor UO_1687 (O_1687,N_14973,N_12402);
nor UO_1688 (O_1688,N_12212,N_14122);
nor UO_1689 (O_1689,N_13112,N_12947);
and UO_1690 (O_1690,N_14102,N_13221);
and UO_1691 (O_1691,N_12462,N_12370);
nand UO_1692 (O_1692,N_13229,N_12489);
nor UO_1693 (O_1693,N_14753,N_14061);
nor UO_1694 (O_1694,N_14882,N_14497);
and UO_1695 (O_1695,N_13736,N_14222);
nand UO_1696 (O_1696,N_12939,N_13508);
and UO_1697 (O_1697,N_12647,N_13369);
nand UO_1698 (O_1698,N_13881,N_13556);
and UO_1699 (O_1699,N_14788,N_12578);
or UO_1700 (O_1700,N_12231,N_14778);
nor UO_1701 (O_1701,N_14947,N_14491);
and UO_1702 (O_1702,N_14589,N_13586);
nor UO_1703 (O_1703,N_13214,N_13414);
or UO_1704 (O_1704,N_14952,N_12606);
nand UO_1705 (O_1705,N_12501,N_13420);
nor UO_1706 (O_1706,N_12918,N_13571);
or UO_1707 (O_1707,N_13032,N_14169);
nand UO_1708 (O_1708,N_13029,N_12178);
nor UO_1709 (O_1709,N_14443,N_14029);
xnor UO_1710 (O_1710,N_13161,N_12565);
nand UO_1711 (O_1711,N_13707,N_13896);
or UO_1712 (O_1712,N_14878,N_14104);
nand UO_1713 (O_1713,N_12966,N_12868);
or UO_1714 (O_1714,N_12678,N_13180);
nor UO_1715 (O_1715,N_13973,N_14522);
xnor UO_1716 (O_1716,N_14568,N_13998);
nor UO_1717 (O_1717,N_13312,N_12988);
xor UO_1718 (O_1718,N_12991,N_14783);
nand UO_1719 (O_1719,N_13462,N_14923);
xor UO_1720 (O_1720,N_14354,N_13631);
and UO_1721 (O_1721,N_13039,N_14736);
nand UO_1722 (O_1722,N_13588,N_12507);
or UO_1723 (O_1723,N_14355,N_13401);
nand UO_1724 (O_1724,N_14734,N_12902);
nor UO_1725 (O_1725,N_12430,N_14824);
xnor UO_1726 (O_1726,N_14896,N_13489);
or UO_1727 (O_1727,N_13580,N_14174);
nand UO_1728 (O_1728,N_13637,N_12746);
nand UO_1729 (O_1729,N_14660,N_12265);
xor UO_1730 (O_1730,N_12973,N_14725);
or UO_1731 (O_1731,N_13895,N_13333);
and UO_1732 (O_1732,N_13493,N_13873);
nand UO_1733 (O_1733,N_14494,N_13815);
or UO_1734 (O_1734,N_13249,N_13658);
nor UO_1735 (O_1735,N_14367,N_14593);
or UO_1736 (O_1736,N_12235,N_12208);
nor UO_1737 (O_1737,N_14719,N_13826);
xor UO_1738 (O_1738,N_13757,N_13946);
nor UO_1739 (O_1739,N_13709,N_14211);
or UO_1740 (O_1740,N_14007,N_14937);
nor UO_1741 (O_1741,N_12264,N_14229);
and UO_1742 (O_1742,N_12236,N_12520);
nor UO_1743 (O_1743,N_14161,N_12241);
and UO_1744 (O_1744,N_14163,N_12917);
and UO_1745 (O_1745,N_14815,N_13969);
nand UO_1746 (O_1746,N_13407,N_13760);
or UO_1747 (O_1747,N_14894,N_12032);
or UO_1748 (O_1748,N_14767,N_14827);
xnor UO_1749 (O_1749,N_12649,N_14628);
nand UO_1750 (O_1750,N_14768,N_12547);
nand UO_1751 (O_1751,N_12567,N_14877);
and UO_1752 (O_1752,N_12277,N_13161);
or UO_1753 (O_1753,N_12473,N_14223);
nor UO_1754 (O_1754,N_13815,N_14778);
nand UO_1755 (O_1755,N_13542,N_14247);
or UO_1756 (O_1756,N_13580,N_13245);
xor UO_1757 (O_1757,N_14769,N_14886);
nand UO_1758 (O_1758,N_13679,N_12578);
xor UO_1759 (O_1759,N_14183,N_13073);
nor UO_1760 (O_1760,N_12670,N_14830);
and UO_1761 (O_1761,N_13559,N_13683);
and UO_1762 (O_1762,N_13248,N_12121);
nor UO_1763 (O_1763,N_12978,N_14931);
nor UO_1764 (O_1764,N_12756,N_13324);
xor UO_1765 (O_1765,N_13534,N_12323);
nor UO_1766 (O_1766,N_13789,N_13885);
nand UO_1767 (O_1767,N_14163,N_13174);
and UO_1768 (O_1768,N_13529,N_13337);
or UO_1769 (O_1769,N_13083,N_12622);
or UO_1770 (O_1770,N_14498,N_14321);
nor UO_1771 (O_1771,N_14338,N_14196);
nor UO_1772 (O_1772,N_14783,N_14747);
and UO_1773 (O_1773,N_13462,N_13837);
nand UO_1774 (O_1774,N_13627,N_12900);
or UO_1775 (O_1775,N_13753,N_12697);
nor UO_1776 (O_1776,N_12446,N_12047);
nand UO_1777 (O_1777,N_12620,N_13586);
xnor UO_1778 (O_1778,N_14375,N_12526);
and UO_1779 (O_1779,N_13751,N_12167);
or UO_1780 (O_1780,N_12908,N_12876);
xnor UO_1781 (O_1781,N_14720,N_14579);
or UO_1782 (O_1782,N_14861,N_12471);
xor UO_1783 (O_1783,N_14850,N_14811);
xor UO_1784 (O_1784,N_14278,N_14515);
or UO_1785 (O_1785,N_12139,N_12770);
nor UO_1786 (O_1786,N_12197,N_13174);
or UO_1787 (O_1787,N_12854,N_13617);
nand UO_1788 (O_1788,N_12176,N_14912);
or UO_1789 (O_1789,N_13707,N_12969);
or UO_1790 (O_1790,N_14306,N_12340);
and UO_1791 (O_1791,N_13362,N_13902);
nor UO_1792 (O_1792,N_12250,N_12912);
xor UO_1793 (O_1793,N_13417,N_14007);
and UO_1794 (O_1794,N_12900,N_14198);
nand UO_1795 (O_1795,N_13074,N_13214);
and UO_1796 (O_1796,N_13449,N_14440);
xnor UO_1797 (O_1797,N_13627,N_13623);
nand UO_1798 (O_1798,N_12824,N_14957);
nor UO_1799 (O_1799,N_12899,N_12388);
xnor UO_1800 (O_1800,N_14325,N_13859);
or UO_1801 (O_1801,N_14155,N_12505);
or UO_1802 (O_1802,N_13068,N_12049);
nand UO_1803 (O_1803,N_14191,N_13840);
nor UO_1804 (O_1804,N_14327,N_12207);
nand UO_1805 (O_1805,N_14980,N_14742);
nand UO_1806 (O_1806,N_12221,N_13669);
nand UO_1807 (O_1807,N_12007,N_14201);
and UO_1808 (O_1808,N_13391,N_12990);
or UO_1809 (O_1809,N_14878,N_14901);
nand UO_1810 (O_1810,N_13460,N_12169);
nor UO_1811 (O_1811,N_14828,N_13281);
nand UO_1812 (O_1812,N_12011,N_14092);
and UO_1813 (O_1813,N_14996,N_13451);
nor UO_1814 (O_1814,N_14489,N_13706);
nor UO_1815 (O_1815,N_14097,N_14927);
nor UO_1816 (O_1816,N_14001,N_12108);
xor UO_1817 (O_1817,N_13271,N_14258);
nor UO_1818 (O_1818,N_12596,N_13314);
xnor UO_1819 (O_1819,N_14043,N_13967);
nor UO_1820 (O_1820,N_14741,N_12212);
nand UO_1821 (O_1821,N_14387,N_14382);
or UO_1822 (O_1822,N_12722,N_13925);
nor UO_1823 (O_1823,N_14645,N_12210);
and UO_1824 (O_1824,N_13579,N_13228);
or UO_1825 (O_1825,N_13960,N_14562);
nand UO_1826 (O_1826,N_12050,N_12244);
or UO_1827 (O_1827,N_13341,N_12756);
or UO_1828 (O_1828,N_12445,N_12258);
or UO_1829 (O_1829,N_13566,N_14807);
and UO_1830 (O_1830,N_13381,N_12305);
and UO_1831 (O_1831,N_13622,N_14657);
and UO_1832 (O_1832,N_12281,N_14898);
nand UO_1833 (O_1833,N_14773,N_14993);
nor UO_1834 (O_1834,N_12351,N_12550);
and UO_1835 (O_1835,N_12993,N_14746);
nor UO_1836 (O_1836,N_14351,N_12723);
nor UO_1837 (O_1837,N_13841,N_13271);
nor UO_1838 (O_1838,N_13916,N_14692);
or UO_1839 (O_1839,N_12622,N_13936);
nor UO_1840 (O_1840,N_12898,N_12540);
nand UO_1841 (O_1841,N_12688,N_14763);
nor UO_1842 (O_1842,N_14327,N_14370);
or UO_1843 (O_1843,N_14356,N_14431);
or UO_1844 (O_1844,N_12015,N_14642);
nand UO_1845 (O_1845,N_13136,N_12019);
nand UO_1846 (O_1846,N_13856,N_12656);
nand UO_1847 (O_1847,N_14697,N_13377);
xnor UO_1848 (O_1848,N_14129,N_14461);
or UO_1849 (O_1849,N_12527,N_12514);
and UO_1850 (O_1850,N_13824,N_12940);
and UO_1851 (O_1851,N_13513,N_12587);
nand UO_1852 (O_1852,N_13516,N_12715);
and UO_1853 (O_1853,N_13540,N_13072);
xnor UO_1854 (O_1854,N_14690,N_14013);
nand UO_1855 (O_1855,N_14642,N_12918);
or UO_1856 (O_1856,N_14405,N_12593);
nand UO_1857 (O_1857,N_12794,N_14791);
nand UO_1858 (O_1858,N_13229,N_12981);
nor UO_1859 (O_1859,N_12151,N_13564);
nor UO_1860 (O_1860,N_12041,N_13672);
nand UO_1861 (O_1861,N_13808,N_13880);
nor UO_1862 (O_1862,N_13066,N_12242);
nor UO_1863 (O_1863,N_12121,N_13743);
nor UO_1864 (O_1864,N_13391,N_14568);
and UO_1865 (O_1865,N_14889,N_12280);
nand UO_1866 (O_1866,N_14820,N_12350);
nand UO_1867 (O_1867,N_13610,N_13549);
or UO_1868 (O_1868,N_14737,N_13810);
nor UO_1869 (O_1869,N_13299,N_14284);
nand UO_1870 (O_1870,N_12629,N_12705);
nand UO_1871 (O_1871,N_13452,N_13381);
and UO_1872 (O_1872,N_12084,N_13945);
and UO_1873 (O_1873,N_13825,N_12892);
and UO_1874 (O_1874,N_12045,N_14015);
and UO_1875 (O_1875,N_13243,N_12188);
and UO_1876 (O_1876,N_13324,N_14536);
and UO_1877 (O_1877,N_12304,N_14177);
nand UO_1878 (O_1878,N_13126,N_12790);
nor UO_1879 (O_1879,N_14183,N_13652);
and UO_1880 (O_1880,N_12117,N_12533);
and UO_1881 (O_1881,N_12187,N_13499);
nand UO_1882 (O_1882,N_12848,N_13504);
or UO_1883 (O_1883,N_12726,N_14879);
or UO_1884 (O_1884,N_12363,N_14902);
and UO_1885 (O_1885,N_13458,N_14250);
nand UO_1886 (O_1886,N_13332,N_12344);
xor UO_1887 (O_1887,N_12772,N_14847);
nor UO_1888 (O_1888,N_14908,N_14726);
nand UO_1889 (O_1889,N_14945,N_14102);
and UO_1890 (O_1890,N_12751,N_12586);
and UO_1891 (O_1891,N_13644,N_12961);
nand UO_1892 (O_1892,N_12792,N_12695);
or UO_1893 (O_1893,N_14240,N_13826);
and UO_1894 (O_1894,N_12518,N_13921);
nor UO_1895 (O_1895,N_13714,N_12571);
or UO_1896 (O_1896,N_14593,N_13974);
nand UO_1897 (O_1897,N_12281,N_12725);
nor UO_1898 (O_1898,N_13524,N_13234);
or UO_1899 (O_1899,N_12437,N_12159);
xor UO_1900 (O_1900,N_12199,N_12555);
nor UO_1901 (O_1901,N_12715,N_13349);
xor UO_1902 (O_1902,N_14212,N_13987);
or UO_1903 (O_1903,N_14574,N_12018);
nand UO_1904 (O_1904,N_13682,N_13569);
nor UO_1905 (O_1905,N_14605,N_14915);
nand UO_1906 (O_1906,N_13648,N_12803);
xor UO_1907 (O_1907,N_13532,N_14757);
nor UO_1908 (O_1908,N_14262,N_12730);
nand UO_1909 (O_1909,N_14313,N_13273);
and UO_1910 (O_1910,N_12679,N_12457);
or UO_1911 (O_1911,N_12212,N_12746);
nand UO_1912 (O_1912,N_14941,N_13451);
nor UO_1913 (O_1913,N_14413,N_14765);
or UO_1914 (O_1914,N_12485,N_13360);
nor UO_1915 (O_1915,N_13681,N_13566);
nand UO_1916 (O_1916,N_14934,N_13703);
nand UO_1917 (O_1917,N_12940,N_12535);
nand UO_1918 (O_1918,N_13615,N_14976);
nor UO_1919 (O_1919,N_12771,N_13242);
or UO_1920 (O_1920,N_14370,N_12096);
or UO_1921 (O_1921,N_14020,N_14548);
and UO_1922 (O_1922,N_13234,N_14642);
and UO_1923 (O_1923,N_14744,N_14807);
or UO_1924 (O_1924,N_13446,N_14672);
and UO_1925 (O_1925,N_12140,N_12054);
xnor UO_1926 (O_1926,N_14737,N_13876);
or UO_1927 (O_1927,N_13073,N_13129);
nand UO_1928 (O_1928,N_14908,N_14011);
xnor UO_1929 (O_1929,N_14938,N_12361);
nor UO_1930 (O_1930,N_14642,N_12930);
and UO_1931 (O_1931,N_14166,N_13886);
or UO_1932 (O_1932,N_12018,N_12117);
or UO_1933 (O_1933,N_14429,N_14835);
and UO_1934 (O_1934,N_13527,N_14660);
nand UO_1935 (O_1935,N_14280,N_13133);
xor UO_1936 (O_1936,N_14398,N_13391);
nand UO_1937 (O_1937,N_14285,N_12696);
or UO_1938 (O_1938,N_14940,N_13196);
xor UO_1939 (O_1939,N_14694,N_12610);
or UO_1940 (O_1940,N_13645,N_12688);
nor UO_1941 (O_1941,N_13654,N_14901);
nand UO_1942 (O_1942,N_12203,N_14480);
or UO_1943 (O_1943,N_12279,N_13484);
and UO_1944 (O_1944,N_14414,N_14952);
and UO_1945 (O_1945,N_12482,N_14674);
and UO_1946 (O_1946,N_13705,N_12063);
and UO_1947 (O_1947,N_12820,N_14347);
or UO_1948 (O_1948,N_14013,N_14614);
nor UO_1949 (O_1949,N_14324,N_13746);
xor UO_1950 (O_1950,N_14993,N_14105);
nor UO_1951 (O_1951,N_12538,N_12224);
and UO_1952 (O_1952,N_14699,N_13219);
nand UO_1953 (O_1953,N_12930,N_12205);
nor UO_1954 (O_1954,N_12875,N_14944);
nor UO_1955 (O_1955,N_12756,N_13625);
xnor UO_1956 (O_1956,N_14773,N_14999);
and UO_1957 (O_1957,N_13534,N_13437);
xor UO_1958 (O_1958,N_14303,N_13590);
nor UO_1959 (O_1959,N_12138,N_13890);
and UO_1960 (O_1960,N_12670,N_13809);
and UO_1961 (O_1961,N_12983,N_14243);
nand UO_1962 (O_1962,N_13108,N_13814);
nor UO_1963 (O_1963,N_14221,N_14800);
nor UO_1964 (O_1964,N_13512,N_13103);
xor UO_1965 (O_1965,N_12201,N_13410);
nor UO_1966 (O_1966,N_13889,N_14472);
or UO_1967 (O_1967,N_12384,N_12393);
and UO_1968 (O_1968,N_13792,N_12053);
nor UO_1969 (O_1969,N_12680,N_13679);
nor UO_1970 (O_1970,N_14227,N_14997);
nand UO_1971 (O_1971,N_13869,N_13589);
or UO_1972 (O_1972,N_14899,N_14359);
nor UO_1973 (O_1973,N_13336,N_13421);
and UO_1974 (O_1974,N_14562,N_13722);
nor UO_1975 (O_1975,N_12246,N_14142);
nor UO_1976 (O_1976,N_13314,N_13589);
nand UO_1977 (O_1977,N_13777,N_14672);
and UO_1978 (O_1978,N_12472,N_12191);
or UO_1979 (O_1979,N_14022,N_12498);
and UO_1980 (O_1980,N_12476,N_14699);
nand UO_1981 (O_1981,N_12732,N_13086);
and UO_1982 (O_1982,N_12743,N_13385);
nand UO_1983 (O_1983,N_12962,N_14250);
and UO_1984 (O_1984,N_14676,N_12200);
and UO_1985 (O_1985,N_12255,N_13484);
and UO_1986 (O_1986,N_13187,N_12100);
or UO_1987 (O_1987,N_13754,N_14165);
nor UO_1988 (O_1988,N_12498,N_14285);
nor UO_1989 (O_1989,N_13217,N_12239);
nor UO_1990 (O_1990,N_14793,N_13626);
or UO_1991 (O_1991,N_13194,N_13468);
nand UO_1992 (O_1992,N_13867,N_12235);
xnor UO_1993 (O_1993,N_12538,N_12111);
xnor UO_1994 (O_1994,N_13122,N_12099);
and UO_1995 (O_1995,N_14766,N_13321);
and UO_1996 (O_1996,N_14336,N_12005);
xnor UO_1997 (O_1997,N_12088,N_13129);
nor UO_1998 (O_1998,N_13964,N_14081);
and UO_1999 (O_1999,N_14184,N_12206);
endmodule