module basic_2500_25000_3000_40_levels_10xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
xor U0 (N_0,In_2230,In_1077);
nor U1 (N_1,In_2346,In_400);
xor U2 (N_2,In_602,In_1284);
xnor U3 (N_3,In_1453,In_2395);
nand U4 (N_4,In_1395,In_1369);
or U5 (N_5,In_1278,In_841);
or U6 (N_6,In_192,In_1089);
nor U7 (N_7,In_851,In_1196);
nor U8 (N_8,In_405,In_853);
nand U9 (N_9,In_1000,In_1379);
nand U10 (N_10,In_1399,In_1195);
nor U11 (N_11,In_807,In_1597);
and U12 (N_12,In_1824,In_689);
nand U13 (N_13,In_1047,In_366);
and U14 (N_14,In_1811,In_2349);
xnor U15 (N_15,In_765,In_1964);
xnor U16 (N_16,In_825,In_1793);
and U17 (N_17,In_791,In_395);
xor U18 (N_18,In_1560,In_532);
nand U19 (N_19,In_2152,In_2248);
xnor U20 (N_20,In_1303,In_615);
xnor U21 (N_21,In_2436,In_1896);
nand U22 (N_22,In_241,In_844);
xor U23 (N_23,In_2244,In_69);
or U24 (N_24,In_418,In_1889);
nand U25 (N_25,In_885,In_1677);
or U26 (N_26,In_565,In_1416);
nor U27 (N_27,In_1070,In_2344);
and U28 (N_28,In_1311,In_1853);
and U29 (N_29,In_2474,In_2100);
nor U30 (N_30,In_2410,In_2191);
xnor U31 (N_31,In_1402,In_1866);
or U32 (N_32,In_421,In_16);
nor U33 (N_33,In_1767,In_652);
nor U34 (N_34,In_2083,In_68);
and U35 (N_35,In_2110,In_500);
or U36 (N_36,In_1271,In_848);
or U37 (N_37,In_518,In_1299);
nor U38 (N_38,In_352,In_353);
nor U39 (N_39,In_137,In_2310);
nand U40 (N_40,In_951,In_2352);
nor U41 (N_41,In_525,In_1334);
nand U42 (N_42,In_1740,In_2124);
and U43 (N_43,In_1405,In_1795);
and U44 (N_44,In_285,In_1673);
or U45 (N_45,In_2207,In_1428);
nand U46 (N_46,In_19,In_1729);
xor U47 (N_47,In_437,In_2296);
xnor U48 (N_48,In_691,In_1883);
nand U49 (N_49,In_1342,In_1653);
nor U50 (N_50,In_2287,In_2336);
nand U51 (N_51,In_222,In_1873);
nand U52 (N_52,In_2351,In_750);
and U53 (N_53,In_876,In_1612);
nand U54 (N_54,In_1063,In_1247);
nor U55 (N_55,In_2113,In_202);
xnor U56 (N_56,In_155,In_2449);
nor U57 (N_57,In_1878,In_2357);
xor U58 (N_58,In_2123,In_1174);
and U59 (N_59,In_1587,In_2243);
xor U60 (N_60,In_917,In_1952);
nand U61 (N_61,In_977,In_799);
or U62 (N_62,In_2046,In_2013);
nand U63 (N_63,In_2014,In_1482);
and U64 (N_64,In_2127,In_2224);
or U65 (N_65,In_1323,In_1121);
or U66 (N_66,In_1851,In_296);
nor U67 (N_67,In_1013,In_1185);
xor U68 (N_68,In_2183,In_601);
and U69 (N_69,In_244,In_1854);
and U70 (N_70,In_10,In_2094);
xor U71 (N_71,In_1689,In_37);
and U72 (N_72,In_840,In_1909);
or U73 (N_73,In_2266,In_987);
xnor U74 (N_74,In_1202,In_2313);
nand U75 (N_75,In_1512,In_217);
and U76 (N_76,In_1627,In_2140);
or U77 (N_77,In_469,In_3);
xor U78 (N_78,In_533,In_588);
and U79 (N_79,In_1559,In_1037);
nor U80 (N_80,In_1274,In_213);
and U81 (N_81,In_862,In_764);
nor U82 (N_82,In_2086,In_179);
and U83 (N_83,In_997,In_1745);
and U84 (N_84,In_2034,In_1118);
xor U85 (N_85,In_173,In_2220);
nor U86 (N_86,In_684,In_1444);
nand U87 (N_87,In_2467,In_436);
xnor U88 (N_88,In_242,In_749);
nor U89 (N_89,In_214,In_77);
xor U90 (N_90,In_2148,In_786);
or U91 (N_91,In_1298,In_2223);
and U92 (N_92,In_664,In_540);
nand U93 (N_93,In_1921,In_967);
and U94 (N_94,In_1862,In_892);
nand U95 (N_95,In_1357,In_252);
nand U96 (N_96,In_1204,In_585);
nor U97 (N_97,In_1438,In_729);
nand U98 (N_98,In_524,In_118);
nor U99 (N_99,In_1147,In_1979);
nor U100 (N_100,In_830,In_649);
nor U101 (N_101,In_1136,In_669);
and U102 (N_102,In_1844,In_555);
nor U103 (N_103,In_1434,In_446);
and U104 (N_104,In_1131,In_2389);
or U105 (N_105,In_1385,In_1557);
xor U106 (N_106,In_546,In_2259);
xor U107 (N_107,In_1447,In_1309);
or U108 (N_108,In_2033,In_1965);
nand U109 (N_109,In_2036,In_866);
or U110 (N_110,In_1578,In_1211);
nor U111 (N_111,In_32,In_1315);
and U112 (N_112,In_483,In_550);
nand U113 (N_113,In_1924,In_2356);
nor U114 (N_114,In_1771,In_371);
nand U115 (N_115,In_466,In_695);
and U116 (N_116,In_2279,In_1799);
nor U117 (N_117,In_171,In_2067);
xnor U118 (N_118,In_2380,In_281);
or U119 (N_119,In_1625,In_337);
nor U120 (N_120,In_598,In_508);
nor U121 (N_121,In_1652,In_519);
and U122 (N_122,In_2403,In_2325);
nor U123 (N_123,In_1456,In_1800);
nor U124 (N_124,In_597,In_578);
xor U125 (N_125,In_341,In_275);
nand U126 (N_126,In_460,In_1540);
nand U127 (N_127,In_1642,In_2070);
nand U128 (N_128,In_2294,In_1571);
nand U129 (N_129,In_2002,In_2493);
nor U130 (N_130,In_1207,In_1582);
xnor U131 (N_131,In_2396,In_526);
nand U132 (N_132,In_170,In_710);
or U133 (N_133,In_1472,In_407);
and U134 (N_134,In_2234,In_1111);
and U135 (N_135,In_109,In_732);
xnor U136 (N_136,In_59,In_186);
nand U137 (N_137,In_1259,In_2055);
nand U138 (N_138,In_2470,In_425);
nor U139 (N_139,In_302,In_1057);
or U140 (N_140,In_333,In_2334);
or U141 (N_141,In_1029,In_2114);
xor U142 (N_142,In_1125,In_2017);
nor U143 (N_143,In_1806,In_1364);
or U144 (N_144,In_2052,In_1366);
nor U145 (N_145,In_1233,In_1160);
or U146 (N_146,In_1452,In_1940);
or U147 (N_147,In_2097,In_2328);
nand U148 (N_148,In_1473,In_1935);
and U149 (N_149,In_1213,In_864);
xor U150 (N_150,In_1167,In_968);
nand U151 (N_151,In_1317,In_2487);
nand U152 (N_152,In_2242,In_1182);
nor U153 (N_153,In_1017,In_75);
nor U154 (N_154,In_295,In_2044);
nand U155 (N_155,In_2262,In_2477);
xor U156 (N_156,In_826,In_1508);
nor U157 (N_157,In_2193,In_1801);
or U158 (N_158,In_625,In_2289);
and U159 (N_159,In_415,In_307);
xor U160 (N_160,In_1216,In_1318);
nand U161 (N_161,In_632,In_1151);
nand U162 (N_162,In_2054,In_326);
and U163 (N_163,In_2031,In_1388);
and U164 (N_164,In_419,In_1992);
and U165 (N_165,In_1887,In_1258);
xor U166 (N_166,In_922,In_283);
nor U167 (N_167,In_551,In_1114);
or U168 (N_168,In_838,In_1078);
and U169 (N_169,In_2197,In_2393);
or U170 (N_170,In_1923,In_1474);
nand U171 (N_171,In_384,In_2150);
nor U172 (N_172,In_2051,In_1297);
nor U173 (N_173,In_2378,In_880);
nand U174 (N_174,In_2306,In_1825);
and U175 (N_175,In_1632,In_809);
or U176 (N_176,In_584,In_231);
xor U177 (N_177,In_2457,In_1647);
nand U178 (N_178,In_660,In_1218);
xnor U179 (N_179,In_2324,In_1228);
xor U180 (N_180,In_2414,In_1351);
nor U181 (N_181,In_45,In_362);
xor U182 (N_182,In_752,In_1948);
and U183 (N_183,In_347,In_1927);
nand U184 (N_184,In_449,In_1367);
xor U185 (N_185,In_1529,In_2442);
and U186 (N_186,In_1613,In_1648);
or U187 (N_187,In_630,In_736);
nor U188 (N_188,In_1208,In_1930);
or U189 (N_189,In_2348,In_1765);
nor U190 (N_190,In_2450,In_638);
nand U191 (N_191,In_639,In_1698);
xor U192 (N_192,In_1541,In_1725);
nand U193 (N_193,In_2060,In_388);
or U194 (N_194,In_380,In_401);
nor U195 (N_195,In_1591,In_1294);
or U196 (N_196,In_2232,In_276);
or U197 (N_197,In_636,In_855);
nor U198 (N_198,In_1250,In_1143);
and U199 (N_199,In_611,In_1814);
xor U200 (N_200,In_210,In_1050);
nand U201 (N_201,In_1676,In_1550);
and U202 (N_202,In_1127,In_132);
and U203 (N_203,In_2292,In_1764);
xor U204 (N_204,In_2432,In_1490);
and U205 (N_205,In_368,In_948);
or U206 (N_206,In_1594,In_795);
nor U207 (N_207,In_2181,In_81);
and U208 (N_208,In_988,In_1024);
nand U209 (N_209,In_2337,In_1021);
nand U210 (N_210,In_1120,In_1713);
nand U211 (N_211,In_129,In_412);
or U212 (N_212,In_1062,In_683);
nor U213 (N_213,In_1105,In_2156);
nand U214 (N_214,In_34,In_1598);
nor U215 (N_215,In_1968,In_2120);
nand U216 (N_216,In_2409,In_1535);
nor U217 (N_217,In_1688,In_1290);
nor U218 (N_218,In_272,In_190);
or U219 (N_219,In_846,In_1789);
nor U220 (N_220,In_1865,In_1666);
or U221 (N_221,In_1545,In_1007);
xor U222 (N_222,In_2275,In_2362);
or U223 (N_223,In_725,In_2219);
nand U224 (N_224,In_268,In_1224);
and U225 (N_225,In_2195,In_43);
and U226 (N_226,In_663,In_2479);
or U227 (N_227,In_2173,In_2321);
or U228 (N_228,In_97,In_1590);
or U229 (N_229,In_2129,In_1156);
and U230 (N_230,In_1069,In_293);
nor U231 (N_231,In_2043,In_1630);
nand U232 (N_232,In_2343,In_1847);
or U233 (N_233,In_2130,In_769);
nand U234 (N_234,In_1735,In_1994);
nand U235 (N_235,In_87,In_46);
nor U236 (N_236,In_1092,In_1929);
nand U237 (N_237,In_22,In_1701);
and U238 (N_238,In_49,In_1392);
nor U239 (N_239,In_2471,In_2061);
nor U240 (N_240,In_2006,In_1991);
or U241 (N_241,In_650,In_1197);
nand U242 (N_242,In_1237,In_1702);
nand U243 (N_243,In_1857,In_2466);
nand U244 (N_244,In_2452,In_2270);
nand U245 (N_245,In_2415,In_334);
and U246 (N_246,In_901,In_2285);
xnor U247 (N_247,In_811,In_775);
nand U248 (N_248,In_290,In_989);
or U249 (N_249,In_2441,In_394);
nand U250 (N_250,In_378,In_816);
and U251 (N_251,In_1645,In_544);
and U252 (N_252,In_1506,In_298);
and U253 (N_253,In_2048,In_1374);
xor U254 (N_254,In_1633,In_1051);
nand U255 (N_255,In_1983,In_1068);
nand U256 (N_256,In_1813,In_1011);
xor U257 (N_257,In_345,In_1236);
xor U258 (N_258,In_1717,In_1526);
xnor U259 (N_259,In_1919,In_376);
nor U260 (N_260,In_392,In_1389);
nand U261 (N_261,In_974,In_7);
and U262 (N_262,In_1030,In_1358);
nand U263 (N_263,In_2162,In_2330);
xnor U264 (N_264,In_1019,In_2288);
or U265 (N_265,In_1465,In_628);
or U266 (N_266,In_1699,In_1839);
or U267 (N_267,In_939,In_125);
nand U268 (N_268,In_1723,In_1706);
and U269 (N_269,In_82,In_616);
and U270 (N_270,In_2167,In_1908);
nand U271 (N_271,In_975,In_724);
or U272 (N_272,In_1959,In_1544);
nand U273 (N_273,In_2421,In_703);
nor U274 (N_274,In_682,In_648);
nand U275 (N_275,In_372,In_1241);
nand U276 (N_276,In_596,In_1296);
xnor U277 (N_277,In_488,In_50);
nor U278 (N_278,In_1422,In_1523);
nand U279 (N_279,In_1410,In_2253);
nand U280 (N_280,In_1166,In_1432);
xor U281 (N_281,In_1175,In_1468);
or U282 (N_282,In_1396,In_2280);
xnor U283 (N_283,In_719,In_2072);
and U284 (N_284,In_2354,In_879);
nor U285 (N_285,In_2082,In_317);
nor U286 (N_286,In_1882,In_1184);
nor U287 (N_287,In_516,In_1020);
xnor U288 (N_288,In_1818,In_1724);
and U289 (N_289,In_557,In_2136);
nand U290 (N_290,In_340,In_2009);
and U291 (N_291,In_463,In_1957);
nand U292 (N_292,In_1662,In_956);
nand U293 (N_293,In_1090,In_356);
and U294 (N_294,In_1322,In_847);
or U295 (N_295,In_2360,In_2087);
nand U296 (N_296,In_733,In_2342);
xnor U297 (N_297,In_2430,In_1257);
nand U298 (N_298,In_1275,In_1163);
or U299 (N_299,In_2426,In_1477);
nor U300 (N_300,In_1770,In_1904);
xor U301 (N_301,In_1816,In_995);
or U302 (N_302,In_146,In_1435);
xnor U303 (N_303,In_163,In_1718);
nand U304 (N_304,In_1665,In_1073);
and U305 (N_305,In_93,In_135);
xor U306 (N_306,In_382,In_1171);
or U307 (N_307,In_172,In_274);
or U308 (N_308,In_1762,In_2160);
xnor U309 (N_309,In_409,In_91);
and U310 (N_310,In_64,In_969);
or U311 (N_311,In_531,In_72);
nor U312 (N_312,In_1335,In_911);
and U313 (N_313,In_324,In_2369);
and U314 (N_314,In_1346,In_600);
nand U315 (N_315,In_2093,In_496);
nand U316 (N_316,In_1514,In_837);
nor U317 (N_317,In_286,In_1549);
nand U318 (N_318,In_1552,In_2390);
nor U319 (N_319,In_1668,In_127);
and U320 (N_320,In_1010,In_2199);
nor U321 (N_321,In_666,In_1144);
xnor U322 (N_322,In_796,In_1530);
nor U323 (N_323,In_918,In_1531);
or U324 (N_324,In_1015,In_1727);
nand U325 (N_325,In_1329,In_2433);
or U326 (N_326,In_965,In_1933);
or U327 (N_327,In_2298,In_1892);
and U328 (N_328,In_2042,In_359);
and U329 (N_329,In_130,In_330);
xnor U330 (N_330,In_692,In_623);
and U331 (N_331,In_1087,In_2134);
and U332 (N_332,In_406,In_888);
xnor U333 (N_333,In_2299,In_604);
xor U334 (N_334,In_2235,In_2018);
and U335 (N_335,In_103,In_1758);
nand U336 (N_336,In_349,In_929);
or U337 (N_337,In_983,In_89);
nand U338 (N_338,In_2165,In_1664);
or U339 (N_339,In_553,In_723);
xnor U340 (N_340,In_1394,In_1577);
xor U341 (N_341,In_2458,In_581);
xor U342 (N_342,In_1067,In_1373);
or U343 (N_343,In_2122,In_2028);
and U344 (N_344,In_1522,In_537);
nor U345 (N_345,In_1270,In_2260);
xnor U346 (N_346,In_2020,In_2071);
nor U347 (N_347,In_2454,In_1451);
nor U348 (N_348,In_1895,In_646);
or U349 (N_349,In_1609,In_755);
nor U350 (N_350,In_574,In_506);
or U351 (N_351,In_819,In_1333);
nand U352 (N_352,In_1621,In_514);
and U353 (N_353,In_731,In_2374);
nor U354 (N_354,In_1169,In_2464);
xnor U355 (N_355,In_1501,In_963);
xor U356 (N_356,In_2213,In_481);
and U357 (N_357,In_2121,In_1567);
or U358 (N_358,In_2168,In_1926);
nor U359 (N_359,In_1542,In_709);
and U360 (N_360,In_1788,In_2332);
or U361 (N_361,In_1489,In_2040);
and U362 (N_362,In_389,In_1097);
and U363 (N_363,In_1235,In_2112);
nor U364 (N_364,In_2143,In_1843);
or U365 (N_365,In_1263,In_836);
nor U366 (N_366,In_2025,In_1859);
xor U367 (N_367,In_925,In_2364);
xnor U368 (N_368,In_679,In_402);
or U369 (N_369,In_735,In_1215);
nor U370 (N_370,In_1797,In_1977);
and U371 (N_371,In_2226,In_2420);
nor U372 (N_372,In_883,In_1879);
xnor U373 (N_373,In_453,In_358);
nor U374 (N_374,In_2145,In_424);
nand U375 (N_375,In_538,In_586);
nand U376 (N_376,In_1960,In_1565);
nor U377 (N_377,In_2473,In_1503);
or U378 (N_378,In_614,In_1918);
nor U379 (N_379,In_1424,In_250);
nand U380 (N_380,In_1832,In_354);
xor U381 (N_381,In_1365,In_2021);
and U382 (N_382,In_687,In_1446);
nand U383 (N_383,In_872,In_1190);
and U384 (N_384,In_2338,In_1354);
or U385 (N_385,In_2315,In_808);
and U386 (N_386,In_502,In_2367);
xnor U387 (N_387,In_696,In_2175);
or U388 (N_388,In_1352,In_727);
and U389 (N_389,In_845,In_1411);
nand U390 (N_390,In_1200,In_908);
nor U391 (N_391,In_1186,In_1679);
and U392 (N_392,In_1807,In_1491);
nand U393 (N_393,In_465,In_1230);
xnor U394 (N_394,In_2178,In_668);
nor U395 (N_395,In_2440,In_954);
nand U396 (N_396,In_292,In_2406);
nand U397 (N_397,In_78,In_914);
nor U398 (N_398,In_79,In_1148);
and U399 (N_399,In_715,In_2462);
or U400 (N_400,In_2335,In_2428);
nand U401 (N_401,In_2290,In_1109);
xor U402 (N_402,In_928,In_20);
xor U403 (N_403,In_2350,In_953);
or U404 (N_404,In_924,In_2203);
or U405 (N_405,In_504,In_1976);
or U406 (N_406,In_2490,In_1611);
nand U407 (N_407,In_306,In_693);
nand U408 (N_408,In_1476,In_1761);
nor U409 (N_409,In_993,In_365);
and U410 (N_410,In_261,In_2375);
xnor U411 (N_411,In_1440,In_1459);
nor U412 (N_412,In_2491,In_145);
and U413 (N_413,In_1561,In_1916);
nor U414 (N_414,In_1016,In_2483);
or U415 (N_415,In_694,In_13);
nor U416 (N_416,In_667,In_1589);
or U417 (N_417,In_2221,In_489);
xor U418 (N_418,In_2188,In_592);
xor U419 (N_419,In_1573,In_1742);
or U420 (N_420,In_780,In_282);
nor U421 (N_421,In_657,In_624);
xor U422 (N_422,In_2465,In_2251);
or U423 (N_423,In_673,In_910);
and U424 (N_424,In_70,In_442);
xnor U425 (N_425,In_2455,In_631);
xor U426 (N_426,In_1980,In_99);
or U427 (N_427,In_2267,In_742);
xnor U428 (N_428,In_1743,In_2016);
xnor U429 (N_429,In_1802,In_2023);
nor U430 (N_430,In_184,In_1641);
and U431 (N_431,In_2258,In_2166);
or U432 (N_432,In_512,In_2102);
and U433 (N_433,In_2116,In_1769);
and U434 (N_434,In_1722,In_120);
nor U435 (N_435,In_219,In_1116);
or U436 (N_436,In_321,In_748);
xor U437 (N_437,In_1488,In_1599);
and U438 (N_438,In_279,In_1112);
and U439 (N_439,In_613,In_1480);
or U440 (N_440,In_932,In_1584);
or U441 (N_441,In_1942,In_232);
and U442 (N_442,In_1040,In_2322);
nor U443 (N_443,In_945,In_2247);
nand U444 (N_444,In_92,In_573);
and U445 (N_445,In_2045,In_2125);
xnor U446 (N_446,In_2495,In_1359);
or U447 (N_447,In_1176,In_964);
or U448 (N_448,In_111,In_1546);
nand U449 (N_449,In_868,In_2416);
xnor U450 (N_450,In_804,In_1507);
and U451 (N_451,In_1220,In_2012);
xnor U452 (N_452,In_534,In_48);
or U453 (N_453,In_1400,In_610);
nand U454 (N_454,In_289,In_1433);
xor U455 (N_455,In_1307,In_416);
xnor U456 (N_456,In_27,In_1135);
nand U457 (N_457,In_161,In_2485);
and U458 (N_458,In_311,In_528);
nand U459 (N_459,In_1782,In_1046);
nand U460 (N_460,In_590,In_738);
xor U461 (N_461,In_1987,In_2497);
nor U462 (N_462,In_671,In_299);
nor U463 (N_463,In_873,In_1055);
or U464 (N_464,In_1846,In_745);
and U465 (N_465,In_1312,In_789);
nand U466 (N_466,In_2076,In_1128);
nor U467 (N_467,In_1036,In_1194);
nor U468 (N_468,In_379,In_547);
nor U469 (N_469,In_823,In_1310);
nand U470 (N_470,In_344,In_1654);
or U471 (N_471,In_1243,In_2439);
or U472 (N_472,In_2399,In_1527);
nand U473 (N_473,In_1255,In_1331);
nor U474 (N_474,In_1860,In_2066);
nand U475 (N_475,In_1988,In_595);
nor U476 (N_476,In_484,In_1970);
nor U477 (N_477,In_480,In_1915);
xor U478 (N_478,In_477,In_1353);
or U479 (N_479,In_834,In_2373);
xor U480 (N_480,In_1781,In_327);
xnor U481 (N_481,In_1371,In_653);
or U482 (N_482,In_1886,In_567);
and U483 (N_483,In_0,In_2307);
nor U484 (N_484,In_2202,In_478);
nand U485 (N_485,In_788,In_1912);
and U486 (N_486,In_1414,In_1426);
and U487 (N_487,In_1272,In_981);
nor U488 (N_488,In_2229,In_1624);
xor U489 (N_489,In_2499,In_95);
or U490 (N_490,In_558,In_1657);
and U491 (N_491,In_1033,In_1044);
xnor U492 (N_492,In_2208,In_1146);
nor U493 (N_493,In_1326,In_1083);
xnor U494 (N_494,In_1242,In_1917);
and U495 (N_495,In_96,In_1252);
xor U496 (N_496,In_2405,In_434);
and U497 (N_497,In_2276,In_447);
or U498 (N_498,In_1821,In_1052);
and U499 (N_499,In_143,In_134);
or U500 (N_500,In_1034,In_433);
nor U501 (N_501,In_1517,In_674);
nor U502 (N_502,In_426,In_1906);
xnor U503 (N_503,In_2463,In_1786);
xor U504 (N_504,In_1875,In_1803);
xor U505 (N_505,In_1709,In_1292);
and U506 (N_506,In_1268,In_2238);
and U507 (N_507,In_973,In_1295);
xnor U508 (N_508,In_350,In_1437);
nor U509 (N_509,In_117,In_2318);
xor U510 (N_510,In_1449,In_776);
nor U511 (N_511,In_2359,In_1752);
and U512 (N_512,In_2039,In_454);
nand U513 (N_513,In_1479,In_2469);
nor U514 (N_514,In_2101,In_589);
nand U515 (N_515,In_935,In_1515);
xor U516 (N_516,In_2233,In_1617);
nand U517 (N_517,In_1925,In_1386);
or U518 (N_518,In_2264,In_462);
nor U519 (N_519,In_2089,In_1219);
nand U520 (N_520,In_1784,In_1443);
nand U521 (N_521,In_2099,In_1967);
and U522 (N_522,In_1817,In_827);
nor U523 (N_523,In_2119,In_2481);
or U524 (N_524,In_877,In_874);
or U525 (N_525,In_1458,In_309);
nand U526 (N_526,In_2079,In_2278);
and U527 (N_527,In_238,In_88);
or U528 (N_528,In_331,In_1093);
nor U529 (N_529,In_1695,In_2381);
or U530 (N_530,In_737,In_1640);
nor U531 (N_531,In_606,In_762);
nor U532 (N_532,In_479,In_2468);
xnor U533 (N_533,In_21,In_385);
and U534 (N_534,In_642,In_2118);
nor U535 (N_535,In_2400,In_1694);
or U536 (N_536,In_2333,In_681);
and U537 (N_537,In_970,In_1377);
xnor U538 (N_538,In_2331,In_1989);
and U539 (N_539,In_881,In_870);
xnor U540 (N_540,In_2053,In_2157);
nor U541 (N_541,In_2447,In_2304);
xor U542 (N_542,In_2418,In_774);
nand U543 (N_543,In_1783,In_404);
xnor U544 (N_544,In_2177,In_1993);
nand U545 (N_545,In_1570,In_1);
nor U546 (N_546,In_1248,In_2303);
or U547 (N_547,In_711,In_47);
xor U548 (N_548,In_1731,In_2010);
xnor U549 (N_549,In_1893,In_1026);
nand U550 (N_550,In_60,In_255);
nand U551 (N_551,In_1280,In_1525);
nor U552 (N_552,In_618,In_18);
xor U553 (N_553,In_1622,In_599);
and U554 (N_554,In_2486,In_226);
and U555 (N_555,In_280,In_1119);
or U556 (N_556,In_1301,In_2392);
and U557 (N_557,In_2158,In_562);
xnor U558 (N_558,In_367,In_1355);
xor U559 (N_559,In_2170,In_1191);
xnor U560 (N_560,In_2309,In_1283);
xnor U561 (N_561,In_1586,In_144);
nor U562 (N_562,In_2323,In_139);
and U563 (N_563,In_63,In_726);
nor U564 (N_564,In_2035,In_545);
nand U565 (N_565,In_235,In_1461);
xnor U566 (N_566,In_1539,In_1672);
nand U567 (N_567,In_1716,In_1823);
or U568 (N_568,In_1249,In_246);
xnor U569 (N_569,In_1707,In_33);
nor U570 (N_570,In_722,In_2004);
and U571 (N_571,In_1958,In_149);
or U572 (N_572,In_1868,In_110);
and U573 (N_573,In_1509,In_443);
nand U574 (N_574,In_157,In_1172);
or U575 (N_575,In_1401,In_2312);
or U576 (N_576,In_1221,In_1644);
or U577 (N_577,In_563,In_1043);
nand U578 (N_578,In_2137,In_1798);
or U579 (N_579,In_943,In_1282);
xor U580 (N_580,In_626,In_106);
nand U581 (N_581,In_100,In_1635);
and U582 (N_582,In_112,In_438);
nand U583 (N_583,In_1705,In_952);
xnor U584 (N_584,In_201,In_781);
or U585 (N_585,In_1867,In_1683);
nor U586 (N_586,In_1619,In_1075);
nor U587 (N_587,In_1870,In_148);
nor U588 (N_588,In_760,In_1132);
nor U589 (N_589,In_1922,In_253);
and U590 (N_590,In_1790,In_121);
and U591 (N_591,In_361,In_2489);
nand U592 (N_592,In_1441,In_1804);
nand U593 (N_593,In_1950,In_915);
or U594 (N_594,In_1203,In_1500);
nand U595 (N_595,In_2057,In_1408);
nor U596 (N_596,In_1238,In_1475);
or U597 (N_597,In_42,In_1686);
nor U598 (N_598,In_1025,In_1888);
or U599 (N_599,In_821,In_1287);
or U600 (N_600,In_1041,In_1792);
nand U601 (N_601,In_1431,In_549);
nor U602 (N_602,In_985,In_230);
xnor U603 (N_603,In_224,In_15);
xor U604 (N_604,In_1406,In_383);
or U605 (N_605,In_5,In_1080);
xnor U606 (N_606,In_1493,In_1142);
xor U607 (N_607,In_2417,In_2271);
and U608 (N_608,In_757,In_1754);
nand U609 (N_609,In_2142,In_784);
nor U610 (N_610,In_2363,In_1834);
nand U611 (N_611,In_1656,In_820);
nor U612 (N_612,In_116,In_1902);
nor U613 (N_613,In_194,In_1520);
and U614 (N_614,In_1183,In_1244);
nand U615 (N_615,In_2425,In_535);
or U616 (N_616,In_39,In_1685);
xor U617 (N_617,In_609,In_278);
nor U618 (N_618,In_1123,In_1462);
xor U619 (N_619,In_1498,In_721);
nor U620 (N_620,In_265,In_1678);
nand U621 (N_621,In_284,In_342);
or U622 (N_622,In_1349,In_491);
xor U623 (N_623,In_759,In_2088);
and U624 (N_624,In_131,In_1830);
nor U625 (N_625,N_463,N_458);
and U626 (N_626,N_171,In_860);
or U627 (N_627,In_2210,In_575);
and U628 (N_628,In_569,In_1251);
or U629 (N_629,In_2090,In_2383);
xor U630 (N_630,N_67,In_1747);
nand U631 (N_631,N_394,In_249);
or U632 (N_632,In_2106,In_867);
nand U633 (N_633,N_494,N_123);
or U634 (N_634,In_54,In_2327);
nor U635 (N_635,N_82,In_1978);
nand U636 (N_636,N_206,In_1494);
nand U637 (N_637,In_2347,In_1324);
nor U638 (N_638,In_572,In_1061);
nand U639 (N_639,In_1894,In_62);
or U640 (N_640,In_818,N_75);
nand U641 (N_641,In_1181,In_2236);
or U642 (N_642,In_474,N_480);
nor U643 (N_643,N_146,In_955);
nor U644 (N_644,In_976,N_231);
xor U645 (N_645,N_105,N_449);
nand U646 (N_646,In_1460,In_1537);
nand U647 (N_647,In_472,In_2078);
nand U648 (N_648,In_1084,In_1605);
nand U649 (N_649,In_1650,In_1534);
nand U650 (N_650,In_36,N_308);
nand U651 (N_651,In_2339,In_960);
and U652 (N_652,In_1532,In_1890);
and U653 (N_653,In_1913,In_2480);
or U654 (N_654,In_1210,In_2214);
xnor U655 (N_655,In_1115,N_447);
or U656 (N_656,In_166,In_758);
xnor U657 (N_657,In_1658,N_608);
nand U658 (N_658,In_822,In_90);
or U659 (N_659,In_2008,N_439);
nand U660 (N_660,N_535,In_271);
xor U661 (N_661,In_893,In_783);
nand U662 (N_662,N_47,In_28);
and U663 (N_663,In_1623,N_419);
nand U664 (N_664,N_484,In_916);
nand U665 (N_665,N_441,In_29);
and U666 (N_666,In_1999,In_2172);
nand U667 (N_667,N_385,In_770);
nor U668 (N_668,In_2075,In_1995);
or U669 (N_669,In_1634,In_1720);
nand U670 (N_670,In_2341,N_8);
or U671 (N_671,N_233,N_468);
or U672 (N_672,In_308,N_173);
and U673 (N_673,In_2402,In_2407);
nor U674 (N_674,N_425,N_96);
or U675 (N_675,In_497,N_309);
nand U676 (N_676,In_1975,In_662);
nand U677 (N_677,N_428,In_1614);
nor U678 (N_678,N_257,N_489);
nor U679 (N_679,In_1356,In_2423);
and U680 (N_680,In_1547,N_345);
or U681 (N_681,In_2404,In_1603);
xor U682 (N_682,In_971,N_359);
nand U683 (N_683,In_114,N_129);
nand U684 (N_684,N_70,In_1738);
or U685 (N_685,N_336,In_661);
or U686 (N_686,In_513,In_1177);
or U687 (N_687,In_998,In_1066);
xor U688 (N_688,N_284,N_88);
nor U689 (N_689,In_771,N_142);
nand U690 (N_690,In_810,In_714);
nor U691 (N_691,N_470,In_451);
or U692 (N_692,In_1231,In_2095);
nand U693 (N_693,In_1751,In_1225);
nor U694 (N_694,In_946,In_2050);
xor U695 (N_695,N_137,In_2190);
xor U696 (N_696,N_438,In_961);
nor U697 (N_697,In_1777,In_133);
xor U698 (N_698,N_311,N_620);
and U699 (N_699,In_793,In_1234);
nand U700 (N_700,N_337,In_17);
and U701 (N_701,N_65,In_1516);
and U702 (N_702,In_2412,In_262);
and U703 (N_703,N_327,In_697);
nand U704 (N_704,N_567,N_261);
and U705 (N_705,In_1376,N_85);
and U706 (N_706,In_267,In_1393);
and U707 (N_707,In_665,N_52);
or U708 (N_708,In_152,In_1332);
nand U709 (N_709,In_593,In_2317);
xnor U710 (N_710,In_1566,In_854);
xnor U711 (N_711,In_369,In_1336);
and U712 (N_712,N_530,N_350);
and U713 (N_713,In_999,In_2117);
nand U714 (N_714,N_303,In_1809);
and U715 (N_715,In_236,N_175);
xor U716 (N_716,In_343,In_832);
and U717 (N_717,N_555,In_1154);
nand U718 (N_718,In_2387,In_445);
nor U719 (N_719,In_958,In_761);
nor U720 (N_720,In_857,In_53);
nor U721 (N_721,In_794,In_884);
nor U722 (N_722,N_424,In_2163);
nand U723 (N_723,In_1058,In_2261);
or U724 (N_724,In_552,In_1165);
nand U725 (N_725,N_242,In_420);
xor U726 (N_726,In_1361,In_2429);
or U727 (N_727,N_48,N_411);
nand U728 (N_728,N_454,In_2272);
nor U729 (N_729,In_1291,In_1099);
or U730 (N_730,In_1188,In_1969);
nand U731 (N_731,In_1226,In_2345);
and U732 (N_732,N_56,In_1126);
nand U733 (N_733,N_2,In_1961);
nand U734 (N_734,In_800,In_1256);
nand U735 (N_735,N_491,N_550);
xnor U736 (N_736,In_1596,N_191);
nand U737 (N_737,In_1056,In_875);
nand U738 (N_738,N_471,In_529);
and U739 (N_739,In_1279,In_741);
and U740 (N_740,N_141,In_523);
xor U741 (N_741,In_408,N_443);
and U742 (N_742,In_889,In_566);
xnor U743 (N_743,In_1576,In_1157);
and U744 (N_744,In_1065,N_585);
nand U745 (N_745,N_456,N_176);
nand U746 (N_746,In_169,N_273);
nor U747 (N_747,In_1528,N_130);
nor U748 (N_748,In_1338,In_338);
nor U749 (N_749,In_1427,In_1002);
nor U750 (N_750,In_2422,In_490);
nor U751 (N_751,In_1982,In_429);
and U752 (N_752,N_103,In_1732);
nor U753 (N_753,In_1316,In_790);
xnor U754 (N_754,In_1604,N_317);
xor U755 (N_755,In_843,N_510);
xor U756 (N_756,In_1054,In_1152);
nand U757 (N_757,N_217,N_253);
or U758 (N_758,In_1240,In_1744);
nor U759 (N_759,In_777,N_114);
nor U760 (N_760,In_1497,N_219);
nand U761 (N_761,In_1649,In_2314);
and U762 (N_762,In_2431,In_1937);
nor U763 (N_763,N_571,N_237);
or U764 (N_764,In_1956,In_1031);
nor U765 (N_765,N_334,In_237);
and U766 (N_766,N_54,In_645);
nand U767 (N_767,In_912,N_312);
and U768 (N_768,In_1341,N_109);
nor U769 (N_769,In_1553,In_1984);
and U770 (N_770,In_174,N_466);
and U771 (N_771,In_448,In_1693);
nor U772 (N_772,N_315,In_1660);
xnor U773 (N_773,In_1363,In_399);
xnor U774 (N_774,In_2268,In_1502);
or U775 (N_775,In_499,In_233);
and U776 (N_776,N_12,In_142);
or U777 (N_777,N_351,In_1189);
nand U778 (N_778,In_1554,N_483);
nand U779 (N_779,In_1733,N_182);
nand U780 (N_780,In_2492,In_2159);
nor U781 (N_781,In_2273,In_905);
or U782 (N_782,N_364,N_73);
xnor U783 (N_783,N_507,In_704);
or U784 (N_784,In_1840,N_262);
xor U785 (N_785,In_2164,In_1778);
or U786 (N_786,N_254,N_586);
or U787 (N_787,In_1254,N_331);
or U788 (N_788,In_2496,In_2059);
xnor U789 (N_789,In_1712,In_699);
xnor U790 (N_790,N_479,N_583);
or U791 (N_791,In_1419,N_560);
nand U792 (N_792,In_211,N_393);
nand U793 (N_793,In_1384,In_2030);
xnor U794 (N_794,In_2019,N_133);
nor U795 (N_795,N_172,In_2187);
nand U796 (N_796,In_2361,N_538);
nor U797 (N_797,In_740,N_348);
or U798 (N_798,In_896,N_529);
nor U799 (N_799,N_258,N_66);
nor U800 (N_800,In_304,In_2027);
or U801 (N_801,N_297,In_1639);
and U802 (N_802,In_1748,N_360);
nor U803 (N_803,In_30,In_897);
or U804 (N_804,N_316,In_1403);
and U805 (N_805,In_1006,In_35);
or U806 (N_806,In_1885,In_2286);
xor U807 (N_807,N_581,In_227);
nand U808 (N_808,In_1305,N_396);
xor U809 (N_809,In_2022,In_351);
nand U810 (N_810,In_942,In_457);
or U811 (N_811,In_1556,In_138);
nand U812 (N_812,In_986,N_383);
nand U813 (N_813,In_539,In_743);
and U814 (N_814,In_1418,In_1700);
nor U815 (N_815,N_473,In_2269);
or U816 (N_816,In_1463,In_782);
nand U817 (N_817,N_545,In_577);
nand U818 (N_818,N_392,In_373);
or U819 (N_819,In_1321,N_220);
or U820 (N_820,N_595,In_2198);
xnor U821 (N_821,N_49,In_2358);
or U822 (N_822,N_404,In_1442);
or U823 (N_823,In_1035,In_387);
and U824 (N_824,In_339,In_1102);
xnor U825 (N_825,In_1643,N_255);
nand U826 (N_826,In_672,In_1193);
and U827 (N_827,In_2494,In_1757);
and U828 (N_828,In_1574,N_24);
nor U829 (N_829,In_2126,In_1362);
xor U830 (N_830,In_1504,In_620);
nor U831 (N_831,In_1420,N_347);
xnor U832 (N_832,N_509,In_2161);
nand U833 (N_833,N_95,In_1928);
and U834 (N_834,N_579,N_128);
xor U835 (N_835,In_57,In_787);
nor U836 (N_836,In_920,In_124);
xor U837 (N_837,N_247,N_611);
nand U838 (N_838,In_1827,In_579);
xor U839 (N_839,In_754,In_205);
xor U840 (N_840,In_1130,In_303);
xnor U841 (N_841,N_162,In_1139);
nand U842 (N_842,In_1785,In_659);
xor U843 (N_843,N_278,N_578);
nor U844 (N_844,In_1253,In_2011);
xor U845 (N_845,N_305,In_108);
and U846 (N_846,N_248,In_2206);
nor U847 (N_847,In_319,In_619);
xnor U848 (N_848,In_414,In_2180);
or U849 (N_849,N_136,In_1773);
nand U850 (N_850,N_416,In_1874);
nand U851 (N_851,In_83,N_120);
nor U852 (N_852,In_323,In_842);
xor U853 (N_853,In_1651,In_1293);
or U854 (N_854,In_1325,In_1768);
nor U855 (N_855,In_1606,N_329);
or U856 (N_856,In_1098,In_2038);
or U857 (N_857,In_1739,In_71);
nor U858 (N_858,N_614,In_31);
and U859 (N_859,N_314,N_263);
xnor U860 (N_860,N_22,In_2250);
or U861 (N_861,In_1631,In_785);
xnor U862 (N_862,In_348,In_390);
nor U863 (N_863,In_2305,In_2302);
nand U864 (N_864,N_157,In_470);
nor U865 (N_865,In_1113,In_2277);
and U866 (N_866,In_1837,In_940);
or U867 (N_867,In_1521,N_161);
or U868 (N_868,In_318,N_169);
and U869 (N_869,N_207,In_1511);
or U870 (N_870,In_766,In_346);
nor U871 (N_871,N_572,N_553);
or U872 (N_872,N_577,N_600);
or U873 (N_873,In_1246,In_1518);
xnor U874 (N_874,In_159,In_1690);
xnor U875 (N_875,N_166,In_1760);
nand U876 (N_876,In_1495,In_1505);
nand U877 (N_877,In_1947,In_1519);
or U878 (N_878,In_655,N_38);
nand U879 (N_879,N_406,In_1187);
or U880 (N_880,N_310,In_435);
nand U881 (N_881,In_907,In_1936);
and U882 (N_882,N_72,In_126);
xnor U883 (N_883,In_1663,N_221);
or U884 (N_884,In_1049,In_927);
or U885 (N_885,N_493,N_541);
xnor U886 (N_886,In_1881,In_957);
or U887 (N_887,N_9,N_324);
xor U888 (N_888,In_6,In_641);
nor U889 (N_889,N_117,In_2241);
nor U890 (N_890,N_402,In_763);
xor U891 (N_891,N_546,N_565);
and U892 (N_892,N_432,N_405);
or U893 (N_893,N_525,In_2385);
or U894 (N_894,N_506,N_164);
or U895 (N_895,In_467,In_128);
nor U896 (N_896,In_1684,In_1996);
nand U897 (N_897,In_1898,In_2209);
xor U898 (N_898,In_162,N_343);
and U899 (N_899,N_64,In_495);
nor U900 (N_900,In_2169,N_260);
or U901 (N_901,N_356,In_605);
nor U902 (N_902,In_1655,In_150);
nor U903 (N_903,N_226,In_1608);
nor U904 (N_904,In_938,N_33);
nor U905 (N_905,In_1387,N_395);
nand U906 (N_906,In_2424,In_328);
nor U907 (N_907,In_1812,In_1610);
or U908 (N_908,N_462,In_2041);
nor U909 (N_909,In_1079,In_2049);
and U910 (N_910,In_1038,In_1593);
or U911 (N_911,N_478,In_439);
nor U912 (N_912,N_218,In_2077);
nor U913 (N_913,In_702,N_26);
nor U914 (N_914,In_895,N_605);
nor U915 (N_915,In_1564,In_1319);
or U916 (N_916,In_188,In_891);
or U917 (N_917,In_1710,In_444);
xnor U918 (N_918,In_1192,In_2189);
xnor U919 (N_919,N_301,In_294);
xor U920 (N_920,In_815,In_1749);
nand U921 (N_921,In_1538,In_966);
nand U922 (N_922,In_1869,N_618);
or U923 (N_923,In_559,In_744);
nor U924 (N_924,In_2092,In_1327);
nor U925 (N_925,In_1133,In_1140);
xnor U926 (N_926,N_288,In_651);
nor U927 (N_927,In_254,N_251);
and U928 (N_928,In_2384,In_1615);
nand U929 (N_929,N_104,In_991);
and U930 (N_930,N_43,N_372);
nor U931 (N_931,In_1421,In_2154);
nand U932 (N_932,N_298,In_1572);
or U933 (N_933,In_1409,N_554);
or U934 (N_934,In_1838,N_234);
xnor U935 (N_935,In_1217,In_2311);
nor U936 (N_936,In_658,In_1345);
and U937 (N_937,In_1510,In_2217);
and U938 (N_938,N_346,In_944);
nor U939 (N_939,In_305,In_1302);
nor U940 (N_940,In_2291,N_126);
or U941 (N_941,In_1581,In_2459);
xor U942 (N_942,In_2015,In_225);
xor U943 (N_943,In_1064,In_1129);
or U944 (N_944,In_1383,N_259);
or U945 (N_945,N_410,N_16);
or U946 (N_946,In_2111,N_341);
or U947 (N_947,In_849,In_1763);
xor U948 (N_948,N_515,N_568);
or U949 (N_949,N_589,In_1304);
xor U950 (N_950,In_530,N_241);
xnor U951 (N_951,In_2293,In_2029);
nand U952 (N_952,N_467,In_1555);
nand U953 (N_953,N_413,In_1951);
and U954 (N_954,N_124,In_1766);
nand U955 (N_955,In_1696,N_59);
nand U956 (N_956,N_597,N_100);
nand U957 (N_957,N_542,N_436);
nand U958 (N_958,N_412,In_1232);
nor U959 (N_959,In_1448,In_1728);
nor U960 (N_960,N_353,In_1772);
nand U961 (N_961,In_921,In_1018);
nand U962 (N_962,In_2081,In_806);
nand U963 (N_963,In_751,In_1831);
nor U964 (N_964,In_982,In_1845);
nor U965 (N_965,In_617,In_2265);
and U966 (N_966,In_1168,In_1138);
nand U967 (N_967,N_17,In_979);
nand U968 (N_968,In_1153,In_153);
nand U969 (N_969,In_260,In_2062);
nor U970 (N_970,In_637,In_1466);
xor U971 (N_971,In_1966,In_492);
or U972 (N_972,In_2453,In_1884);
and U973 (N_973,N_211,In_2460);
or U974 (N_974,In_747,In_1990);
and U975 (N_975,N_584,N_87);
nor U976 (N_976,In_332,In_950);
or U977 (N_977,In_200,In_1714);
and U978 (N_978,N_80,In_322);
or U979 (N_979,In_423,In_1450);
nor U980 (N_980,In_906,In_1158);
nor U981 (N_981,In_768,In_507);
or U982 (N_982,In_670,N_528);
nand U983 (N_983,In_2171,N_99);
and U984 (N_984,In_2445,In_1481);
or U985 (N_985,In_288,N_318);
nand U986 (N_986,In_1946,In_1891);
xor U987 (N_987,In_959,In_417);
or U988 (N_988,N_374,In_1398);
and U989 (N_989,N_184,In_992);
or U990 (N_990,In_165,N_152);
xor U991 (N_991,N_603,In_2068);
xor U992 (N_992,In_561,In_141);
nand U993 (N_993,In_493,N_28);
and U994 (N_994,In_115,In_1855);
xor U995 (N_995,In_2001,In_1900);
nor U996 (N_996,In_1580,In_65);
or U997 (N_997,N_401,In_1145);
and U998 (N_998,In_2228,In_158);
and U999 (N_999,In_1585,N_62);
and U1000 (N_1000,In_1134,In_1071);
or U1001 (N_1001,In_1730,In_640);
or U1002 (N_1002,N_596,N_592);
and U1003 (N_1003,N_369,In_2215);
nand U1004 (N_1004,In_2446,N_623);
nand U1005 (N_1005,In_2133,N_83);
or U1006 (N_1006,In_2326,N_526);
nand U1007 (N_1007,N_204,In_2115);
xnor U1008 (N_1008,In_1288,In_259);
xor U1009 (N_1009,In_1464,In_403);
or U1010 (N_1010,N_299,In_1638);
or U1011 (N_1011,In_256,N_434);
nor U1012 (N_1012,In_1430,In_2456);
or U1013 (N_1013,N_476,In_542);
xnor U1014 (N_1014,In_1796,In_26);
and U1015 (N_1015,In_792,In_413);
nand U1016 (N_1016,In_1005,In_2249);
and U1017 (N_1017,N_14,In_1938);
nor U1018 (N_1018,N_181,In_2204);
nor U1019 (N_1019,In_919,N_504);
or U1020 (N_1020,In_1637,N_264);
or U1021 (N_1021,N_373,In_325);
xnor U1022 (N_1022,N_1,N_144);
and U1023 (N_1023,In_175,N_461);
xnor U1024 (N_1024,N_222,N_193);
and U1025 (N_1025,In_2135,N_472);
xnor U1026 (N_1026,In_878,N_403);
or U1027 (N_1027,In_2107,In_1949);
nand U1028 (N_1028,In_1903,N_534);
nor U1029 (N_1029,In_1277,In_852);
nor U1030 (N_1030,N_10,N_268);
or U1031 (N_1031,In_1558,In_101);
and U1032 (N_1032,In_1822,In_167);
nand U1033 (N_1033,In_1391,In_2320);
or U1034 (N_1034,In_1022,In_1810);
xor U1035 (N_1035,In_1469,In_548);
or U1036 (N_1036,N_452,N_76);
nand U1037 (N_1037,N_203,In_270);
nand U1038 (N_1038,N_238,N_132);
nor U1039 (N_1039,In_1934,N_167);
and U1040 (N_1040,In_1239,N_368);
nand U1041 (N_1041,In_773,In_858);
nand U1042 (N_1042,N_492,In_41);
or U1043 (N_1043,In_707,In_1897);
nor U1044 (N_1044,N_236,In_1931);
nor U1045 (N_1045,In_2394,N_576);
nand U1046 (N_1046,In_104,In_2074);
nor U1047 (N_1047,In_1042,In_398);
or U1048 (N_1048,In_273,N_230);
or U1049 (N_1049,In_8,N_588);
nor U1050 (N_1050,In_2488,In_2355);
nand U1051 (N_1051,N_41,In_66);
xnor U1052 (N_1052,N_205,In_377);
xnor U1053 (N_1053,In_198,In_107);
nand U1054 (N_1054,N_290,In_428);
or U1055 (N_1055,N_287,In_2476);
nand U1056 (N_1056,In_24,In_1850);
nor U1057 (N_1057,In_2316,N_519);
or U1058 (N_1058,In_264,In_1380);
nor U1059 (N_1059,In_772,N_397);
xnor U1060 (N_1060,In_1081,N_422);
or U1061 (N_1061,In_1626,In_1543);
or U1062 (N_1062,In_1741,In_2146);
and U1063 (N_1063,N_147,In_2382);
nand U1064 (N_1064,In_2401,In_316);
or U1065 (N_1065,In_509,N_332);
and U1066 (N_1066,In_1164,N_79);
nand U1067 (N_1067,N_197,In_886);
nor U1068 (N_1068,N_450,N_279);
nand U1069 (N_1069,N_178,In_1091);
and U1070 (N_1070,In_498,N_399);
xnor U1071 (N_1071,In_690,In_56);
nand U1072 (N_1072,In_485,N_415);
xnor U1073 (N_1073,In_1155,In_228);
xnor U1074 (N_1074,In_2005,In_1575);
or U1075 (N_1075,In_2155,In_1836);
nand U1076 (N_1076,In_269,N_617);
or U1077 (N_1077,N_20,In_1286);
and U1078 (N_1078,N_556,In_1170);
nand U1079 (N_1079,N_296,In_1941);
nand U1080 (N_1080,In_1682,In_287);
nor U1081 (N_1081,N_201,In_1791);
xnor U1082 (N_1082,In_140,In_1704);
or U1083 (N_1083,In_949,In_1141);
nand U1084 (N_1084,In_84,In_813);
nand U1085 (N_1085,N_469,In_1390);
or U1086 (N_1086,In_2185,In_300);
or U1087 (N_1087,In_386,In_1397);
or U1088 (N_1088,In_521,In_183);
xnor U1089 (N_1089,N_3,In_2056);
nand U1090 (N_1090,N_186,In_1161);
nor U1091 (N_1091,In_803,In_2073);
nor U1092 (N_1092,In_582,In_2368);
or U1093 (N_1093,N_97,N_482);
nand U1094 (N_1094,In_1340,N_602);
xnor U1095 (N_1095,In_2239,N_282);
or U1096 (N_1096,In_734,N_51);
and U1097 (N_1097,In_996,N_185);
nor U1098 (N_1098,N_420,In_2085);
nor U1099 (N_1099,N_503,In_248);
and U1100 (N_1100,In_458,In_1425);
nor U1101 (N_1101,N_570,In_1588);
nor U1102 (N_1102,In_1378,In_933);
nand U1103 (N_1103,In_2427,In_1162);
xor U1104 (N_1104,N_266,N_517);
or U1105 (N_1105,In_486,In_1944);
or U1106 (N_1106,In_2065,In_310);
nand U1107 (N_1107,In_1262,In_1150);
and U1108 (N_1108,In_247,N_612);
nor U1109 (N_1109,In_1628,In_1375);
xor U1110 (N_1110,In_74,N_125);
nand U1111 (N_1111,N_621,In_1173);
xor U1112 (N_1112,In_1669,In_1229);
or U1113 (N_1113,In_1308,In_635);
and U1114 (N_1114,N_485,In_1985);
and U1115 (N_1115,In_2222,N_112);
or U1116 (N_1116,In_1939,In_2372);
nand U1117 (N_1117,In_2069,In_1780);
nand U1118 (N_1118,In_947,N_557);
xnor U1119 (N_1119,In_1027,In_297);
and U1120 (N_1120,In_1276,In_1680);
or U1121 (N_1121,N_379,N_295);
nor U1122 (N_1122,In_720,In_554);
nor U1123 (N_1123,N_382,In_1963);
xnor U1124 (N_1124,In_1600,In_1212);
xor U1125 (N_1125,In_580,N_209);
nor U1126 (N_1126,In_1439,In_468);
and U1127 (N_1127,N_165,In_335);
or U1128 (N_1128,In_2200,In_1899);
or U1129 (N_1129,In_1085,In_320);
and U1130 (N_1130,N_501,N_291);
and U1131 (N_1131,N_239,In_1997);
nand U1132 (N_1132,In_1674,In_1214);
or U1133 (N_1133,N_335,In_177);
and U1134 (N_1134,N_232,In_923);
or U1135 (N_1135,N_155,In_430);
and U1136 (N_1136,In_2196,In_1776);
nand U1137 (N_1137,In_431,N_378);
nand U1138 (N_1138,In_700,N_322);
and U1139 (N_1139,N_442,In_1986);
and U1140 (N_1140,In_51,N_69);
nand U1141 (N_1141,N_281,N_371);
and U1142 (N_1142,In_594,In_1445);
nand U1143 (N_1143,In_1267,In_937);
and U1144 (N_1144,In_1028,N_340);
xnor U1145 (N_1145,In_1101,N_294);
or U1146 (N_1146,N_569,In_2461);
nand U1147 (N_1147,N_27,In_2192);
nor U1148 (N_1148,In_1199,In_1486);
or U1149 (N_1149,In_902,In_656);
and U1150 (N_1150,N_326,In_1719);
xnor U1151 (N_1151,In_778,In_156);
xnor U1152 (N_1152,In_1370,In_1088);
xor U1153 (N_1153,In_1330,In_2174);
xor U1154 (N_1154,In_903,N_223);
and U1155 (N_1155,N_194,N_225);
xor U1156 (N_1156,In_2300,In_930);
nor U1157 (N_1157,N_150,In_2435);
nand U1158 (N_1158,In_1998,N_516);
xnor U1159 (N_1159,In_1266,N_562);
or U1160 (N_1160,In_452,N_559);
and U1161 (N_1161,In_154,N_609);
and U1162 (N_1162,In_2419,In_1708);
xnor U1163 (N_1163,In_972,In_1955);
or U1164 (N_1164,In_1945,N_487);
nor U1165 (N_1165,In_1629,N_44);
nor U1166 (N_1166,In_455,N_0);
or U1167 (N_1167,In_1858,N_35);
and U1168 (N_1168,In_1618,In_515);
nor U1169 (N_1169,In_2283,In_1269);
nor U1170 (N_1170,In_1607,N_19);
and U1171 (N_1171,In_2377,N_544);
and U1172 (N_1172,N_92,In_2184);
xnor U1173 (N_1173,In_536,In_1412);
nor U1174 (N_1174,In_2246,N_440);
xor U1175 (N_1175,N_537,In_2281);
nor U1176 (N_1176,N_102,In_718);
or U1177 (N_1177,N_499,N_307);
nor U1178 (N_1178,N_159,In_52);
xor U1179 (N_1179,N_50,In_798);
xnor U1180 (N_1180,In_370,In_2064);
or U1181 (N_1181,In_871,In_583);
or U1182 (N_1182,In_1094,N_116);
and U1183 (N_1183,In_1048,N_246);
nor U1184 (N_1184,In_801,In_1137);
or U1185 (N_1185,In_1750,In_381);
nand U1186 (N_1186,In_1382,In_612);
or U1187 (N_1187,In_314,N_199);
nor U1188 (N_1188,N_77,In_1009);
and U1189 (N_1189,In_4,In_2329);
xnor U1190 (N_1190,In_1159,N_86);
and U1191 (N_1191,In_301,N_333);
or U1192 (N_1192,In_1914,In_629);
nor U1193 (N_1193,N_156,N_6);
xor U1194 (N_1194,In_746,N_512);
and U1195 (N_1195,N_418,In_1863);
nand U1196 (N_1196,N_275,In_1852);
nand U1197 (N_1197,In_1039,N_240);
nand U1198 (N_1198,N_437,N_551);
or U1199 (N_1199,In_2000,In_189);
or U1200 (N_1200,N_270,In_1053);
nor U1201 (N_1201,In_587,N_423);
xor U1202 (N_1202,In_1004,N_342);
or U1203 (N_1203,In_203,In_621);
nand U1204 (N_1204,In_2301,N_582);
or U1205 (N_1205,N_409,In_12);
and U1206 (N_1206,In_2282,In_2478);
or U1207 (N_1207,In_2003,N_195);
nor U1208 (N_1208,In_2443,In_1060);
nand U1209 (N_1209,N_384,N_457);
and U1210 (N_1210,In_2194,In_2103);
nor U1211 (N_1211,In_1273,In_355);
and U1212 (N_1212,In_1045,N_58);
and U1213 (N_1213,N_229,In_1646);
nand U1214 (N_1214,In_2411,N_63);
xnor U1215 (N_1215,In_329,N_154);
and U1216 (N_1216,In_2295,In_9);
and U1217 (N_1217,N_448,In_994);
or U1218 (N_1218,N_25,In_1681);
xor U1219 (N_1219,In_1471,In_1616);
and U1220 (N_1220,In_1108,In_654);
or U1221 (N_1221,N_451,In_427);
xnor U1222 (N_1222,In_560,N_619);
xnor U1223 (N_1223,N_622,In_1602);
nor U1224 (N_1224,In_1954,N_601);
nand U1225 (N_1225,N_274,N_108);
nand U1226 (N_1226,N_358,In_1943);
and U1227 (N_1227,In_2245,In_2);
nor U1228 (N_1228,In_2252,In_229);
nand U1229 (N_1229,In_1003,In_622);
nand U1230 (N_1230,In_2105,N_57);
and U1231 (N_1231,In_1794,N_163);
or U1232 (N_1232,N_119,N_289);
and U1233 (N_1233,In_2201,In_634);
nand U1234 (N_1234,N_558,N_344);
nand U1235 (N_1235,In_220,N_446);
xnor U1236 (N_1236,In_216,In_1849);
or U1237 (N_1237,N_514,In_1692);
xor U1238 (N_1238,N_139,In_1313);
and U1239 (N_1239,In_1348,N_30);
xnor U1240 (N_1240,N_252,N_313);
xor U1241 (N_1241,In_151,In_2231);
and U1242 (N_1242,N_536,N_180);
and U1243 (N_1243,In_14,In_1551);
xnor U1244 (N_1244,N_573,In_122);
nor U1245 (N_1245,N_74,In_644);
nand U1246 (N_1246,In_1910,In_2131);
nor U1247 (N_1247,In_1223,In_119);
xor U1248 (N_1248,N_216,In_2371);
nor U1249 (N_1249,In_1289,N_101);
and U1250 (N_1250,In_2472,In_94);
xor U1251 (N_1251,N_196,N_1242);
nand U1252 (N_1252,N_692,N_1049);
nor U1253 (N_1253,N_98,N_189);
and U1254 (N_1254,In_2237,N_115);
or U1255 (N_1255,N_751,In_2128);
or U1256 (N_1256,In_1703,N_709);
nor U1257 (N_1257,N_352,N_829);
nand U1258 (N_1258,N_840,N_776);
or U1259 (N_1259,N_690,N_794);
nor U1260 (N_1260,N_435,N_675);
xor U1261 (N_1261,In_204,N_215);
and U1262 (N_1262,N_767,In_839);
xnor U1263 (N_1263,In_767,In_779);
or U1264 (N_1264,N_989,N_304);
nand U1265 (N_1265,N_68,N_1058);
nor U1266 (N_1266,N_791,N_798);
or U1267 (N_1267,N_391,N_818);
and U1268 (N_1268,N_177,In_1864);
xnor U1269 (N_1269,N_60,N_1249);
and U1270 (N_1270,In_730,N_1031);
nor U1271 (N_1271,N_477,In_206);
nor U1272 (N_1272,N_1081,In_2058);
xnor U1273 (N_1273,N_963,In_2144);
and U1274 (N_1274,N_1084,In_1306);
nand U1275 (N_1275,N_964,N_1141);
nand U1276 (N_1276,N_755,In_556);
nor U1277 (N_1277,N_639,N_668);
or U1278 (N_1278,N_256,N_782);
or U1279 (N_1279,N_1202,N_407);
nand U1280 (N_1280,N_1183,N_630);
nand U1281 (N_1281,N_148,N_812);
nand U1282 (N_1282,N_1135,N_743);
nand U1283 (N_1283,N_1123,In_1261);
and U1284 (N_1284,N_160,N_946);
nand U1285 (N_1285,N_886,N_736);
and U1286 (N_1286,N_1113,N_210);
xor U1287 (N_1287,N_681,N_1157);
nor U1288 (N_1288,In_712,In_2388);
nand U1289 (N_1289,In_2437,N_953);
nand U1290 (N_1290,N_1194,In_1721);
xor U1291 (N_1291,N_190,In_11);
and U1292 (N_1292,N_1119,N_1064);
nor U1293 (N_1293,In_510,N_660);
nor U1294 (N_1294,N_903,In_441);
nor U1295 (N_1295,N_375,N_1230);
or U1296 (N_1296,N_1037,N_1021);
xnor U1297 (N_1297,In_86,In_1023);
xor U1298 (N_1298,In_1300,In_1110);
nor U1299 (N_1299,N_1088,In_257);
and U1300 (N_1300,N_21,N_361);
and U1301 (N_1301,In_2216,In_1726);
xor U1302 (N_1302,In_73,N_465);
nor U1303 (N_1303,N_1114,N_912);
nor U1304 (N_1304,In_1524,N_227);
nor U1305 (N_1305,In_647,N_1196);
and U1306 (N_1306,In_1972,In_2370);
xor U1307 (N_1307,N_844,In_209);
or U1308 (N_1308,In_708,N_122);
xor U1309 (N_1309,N_780,N_656);
xor U1310 (N_1310,In_1492,N_1002);
xnor U1311 (N_1311,N_267,In_375);
and U1312 (N_1312,In_1971,In_2080);
nor U1313 (N_1313,N_1190,N_521);
or U1314 (N_1314,N_749,In_1149);
xnor U1315 (N_1315,In_2218,N_1011);
and U1316 (N_1316,N_78,In_833);
and U1317 (N_1317,In_1436,N_1187);
nor U1318 (N_1318,N_1105,N_46);
xnor U1319 (N_1319,N_627,N_1087);
xnor U1320 (N_1320,N_1147,N_905);
and U1321 (N_1321,N_1034,In_828);
nor U1322 (N_1322,N_1211,N_408);
nor U1323 (N_1323,N_1038,N_249);
xnor U1324 (N_1324,N_1056,N_914);
nor U1325 (N_1325,In_931,N_1017);
nor U1326 (N_1326,In_80,N_13);
or U1327 (N_1327,N_982,N_1215);
or U1328 (N_1328,N_320,N_1166);
and U1329 (N_1329,N_978,N_824);
xor U1330 (N_1330,N_670,N_1239);
and U1331 (N_1331,N_1096,N_1152);
nand U1332 (N_1332,N_934,N_673);
nand U1333 (N_1333,N_213,N_575);
or U1334 (N_1334,In_1826,N_956);
and U1335 (N_1335,N_661,N_928);
and U1336 (N_1336,N_1047,In_2141);
nand U1337 (N_1337,N_677,N_710);
nor U1338 (N_1338,In_199,N_417);
nand U1339 (N_1339,N_1244,In_2151);
nor U1340 (N_1340,In_698,In_1711);
nor U1341 (N_1341,N_430,N_1167);
or U1342 (N_1342,N_629,N_722);
xnor U1343 (N_1343,N_111,N_663);
xnor U1344 (N_1344,In_182,N_981);
nor U1345 (N_1345,N_752,N_857);
or U1346 (N_1346,N_868,In_1423);
xnor U1347 (N_1347,N_907,In_856);
nor U1348 (N_1348,N_390,N_887);
xor U1349 (N_1349,N_93,In_898);
xor U1350 (N_1350,In_1671,N_276);
and U1351 (N_1351,In_1072,N_822);
nand U1352 (N_1352,In_58,N_387);
or U1353 (N_1353,N_727,In_23);
xnor U1354 (N_1354,N_856,N_804);
nand U1355 (N_1355,N_1205,N_1132);
nand U1356 (N_1356,N_1228,N_626);
nor U1357 (N_1357,N_662,In_814);
nor U1358 (N_1358,In_1568,N_84);
and U1359 (N_1359,In_517,N_55);
or U1360 (N_1360,In_185,N_153);
nand U1361 (N_1361,N_979,In_1670);
or U1362 (N_1362,N_682,In_1533);
nand U1363 (N_1363,N_563,N_1158);
or U1364 (N_1364,N_871,In_1106);
nor U1365 (N_1365,In_1636,N_1007);
nor U1366 (N_1366,N_796,In_1872);
xor U1367 (N_1367,N_958,In_1407);
nor U1368 (N_1368,In_756,N_962);
nand U1369 (N_1369,N_587,N_1090);
xor U1370 (N_1370,N_1137,In_1227);
and U1371 (N_1371,In_1457,In_440);
xor U1372 (N_1372,N_1010,N_1125);
and U1373 (N_1373,In_869,N_878);
nor U1374 (N_1374,In_397,N_431);
nor U1375 (N_1375,N_547,In_2026);
nor U1376 (N_1376,In_863,N_781);
and U1377 (N_1377,N_854,In_1201);
or U1378 (N_1378,In_1245,N_1101);
or U1379 (N_1379,N_730,In_2366);
and U1380 (N_1380,N_1035,N_695);
and U1381 (N_1381,In_1687,N_877);
xnor U1382 (N_1382,N_398,N_616);
nor U1383 (N_1383,In_450,N_355);
or U1384 (N_1384,N_968,N_269);
xnor U1385 (N_1385,N_1062,N_811);
nor U1386 (N_1386,N_145,N_362);
and U1387 (N_1387,In_1180,In_2379);
or U1388 (N_1388,N_18,N_726);
nor U1389 (N_1389,N_659,N_635);
or U1390 (N_1390,In_2498,N_739);
xor U1391 (N_1391,N_183,N_518);
nor U1392 (N_1392,In_1835,N_23);
nor U1393 (N_1393,N_740,In_1715);
nand U1394 (N_1394,In_432,N_890);
nor U1395 (N_1395,In_1082,In_1842);
nand U1396 (N_1396,N_976,N_813);
xnor U1397 (N_1397,N_140,N_513);
nor U1398 (N_1398,N_935,N_292);
nand U1399 (N_1399,N_1041,In_1981);
nand U1400 (N_1400,N_858,N_870);
xnor U1401 (N_1401,In_1008,N_961);
nand U1402 (N_1402,In_494,N_604);
xnor U1403 (N_1403,N_841,N_994);
nand U1404 (N_1404,N_1120,N_1209);
nor U1405 (N_1405,N_993,In_941);
and U1406 (N_1406,N_872,N_703);
or U1407 (N_1407,N_36,In_487);
nor U1408 (N_1408,N_1069,N_1188);
nor U1409 (N_1409,In_2308,N_945);
or U1410 (N_1410,In_208,N_1046);
and U1411 (N_1411,N_899,N_1036);
or U1412 (N_1412,In_266,N_941);
and U1413 (N_1413,In_1347,N_107);
and U1414 (N_1414,N_1076,N_1203);
nor U1415 (N_1415,N_884,N_1159);
nor U1416 (N_1416,In_1737,N_771);
and U1417 (N_1417,N_977,N_599);
or U1418 (N_1418,N_669,N_1027);
or U1419 (N_1419,In_180,In_1381);
nor U1420 (N_1420,In_464,N_1082);
xor U1421 (N_1421,In_102,N_202);
or U1422 (N_1422,N_971,N_495);
nand U1423 (N_1423,N_293,N_121);
or U1424 (N_1424,N_650,N_1186);
nand U1425 (N_1425,In_1974,N_915);
xnor U1426 (N_1426,N_932,In_701);
nand U1427 (N_1427,In_422,N_665);
and U1428 (N_1428,N_834,N_806);
nand U1429 (N_1429,N_893,N_634);
xor U1430 (N_1430,N_732,In_887);
or U1431 (N_1431,N_944,N_1029);
and U1432 (N_1432,In_393,N_1138);
or U1433 (N_1433,In_187,N_498);
and U1434 (N_1434,N_481,N_947);
and U1435 (N_1435,In_2254,N_1172);
nand U1436 (N_1436,In_1281,In_239);
xor U1437 (N_1437,In_2227,N_1164);
or U1438 (N_1438,N_1216,N_1191);
nor U1439 (N_1439,N_386,In_1096);
nor U1440 (N_1440,N_879,N_1104);
xnor U1441 (N_1441,In_1759,N_833);
nor U1442 (N_1442,In_728,In_797);
xnor U1443 (N_1443,N_734,In_2147);
or U1444 (N_1444,N_725,N_496);
nor U1445 (N_1445,N_110,In_1911);
xnor U1446 (N_1446,N_1079,In_1962);
or U1447 (N_1447,In_900,N_738);
and U1448 (N_1448,In_1734,N_502);
and U1449 (N_1449,N_859,N_357);
and U1450 (N_1450,N_939,N_678);
or U1451 (N_1451,N_1127,N_633);
nand U1452 (N_1452,N_867,In_1339);
xnor U1453 (N_1453,N_885,N_745);
xor U1454 (N_1454,N_32,In_1973);
nand U1455 (N_1455,In_1736,N_852);
nor U1456 (N_1456,N_214,N_951);
or U1457 (N_1457,In_1746,N_552);
nor U1458 (N_1458,In_859,N_625);
nand U1459 (N_1459,N_339,N_645);
nor U1460 (N_1460,In_1001,N_224);
nor U1461 (N_1461,N_149,In_277);
xor U1462 (N_1462,N_674,N_540);
and U1463 (N_1463,N_1221,N_790);
xnor U1464 (N_1464,N_1004,In_223);
and U1465 (N_1465,N_904,In_2098);
nand U1466 (N_1466,In_1871,In_1828);
and U1467 (N_1467,N_1165,N_1055);
or U1468 (N_1468,In_2091,In_1372);
nand U1469 (N_1469,In_1417,In_1496);
xor U1470 (N_1470,In_1198,In_1014);
xnor U1471 (N_1471,In_984,In_136);
xnor U1472 (N_1472,In_105,N_762);
nand U1473 (N_1473,N_991,In_1815);
xor U1474 (N_1474,N_655,N_706);
xnor U1475 (N_1475,In_2149,In_243);
or U1476 (N_1476,N_913,In_482);
nor U1477 (N_1477,N_1161,In_1513);
or U1478 (N_1478,N_644,In_1178);
or U1479 (N_1479,N_574,In_608);
and U1480 (N_1480,N_1059,N_1028);
xnor U1481 (N_1481,In_1264,N_511);
xor U1482 (N_1482,In_234,In_147);
or U1483 (N_1483,N_208,N_920);
nand U1484 (N_1484,N_658,N_720);
and U1485 (N_1485,In_1876,In_181);
or U1486 (N_1486,N_363,N_1030);
or U1487 (N_1487,In_527,In_476);
or U1488 (N_1488,In_2386,N_948);
nand U1489 (N_1489,N_1219,In_909);
and U1490 (N_1490,N_733,N_775);
or U1491 (N_1491,In_2138,N_694);
nand U1492 (N_1492,In_503,In_2032);
nor U1493 (N_1493,N_1179,N_37);
xor U1494 (N_1494,In_1100,N_966);
and U1495 (N_1495,In_25,N_786);
and U1496 (N_1496,N_960,In_1841);
or U1497 (N_1497,In_1320,N_1052);
nand U1498 (N_1498,N_1111,N_975);
and U1499 (N_1499,N_91,In_1455);
nand U1500 (N_1500,N_170,N_711);
xor U1501 (N_1501,N_1097,N_651);
nor U1502 (N_1502,N_328,In_2434);
or U1503 (N_1503,N_768,In_520);
nand U1504 (N_1504,In_1483,N_680);
xor U1505 (N_1505,N_500,N_135);
nor U1506 (N_1506,N_937,N_286);
or U1507 (N_1507,N_919,In_1536);
and U1508 (N_1508,N_922,N_803);
xor U1509 (N_1509,N_647,In_713);
and U1510 (N_1510,In_85,N_81);
nor U1511 (N_1511,In_2484,N_188);
nand U1512 (N_1512,N_632,N_365);
nand U1513 (N_1513,In_1756,In_501);
nor U1514 (N_1514,In_336,N_637);
nor U1515 (N_1515,N_134,N_1229);
xnor U1516 (N_1516,N_1177,N_783);
or U1517 (N_1517,N_967,In_1487);
nor U1518 (N_1518,N_127,N_272);
xor U1519 (N_1519,In_1753,N_696);
nand U1520 (N_1520,N_929,N_1181);
nand U1521 (N_1521,N_624,N_1122);
or U1522 (N_1522,N_1083,In_802);
nand U1523 (N_1523,N_90,N_1023);
xnor U1524 (N_1524,N_992,N_1234);
nor U1525 (N_1525,N_192,In_1819);
and U1526 (N_1526,N_931,N_1149);
xnor U1527 (N_1527,N_787,N_549);
xor U1528 (N_1528,In_471,N_837);
and U1529 (N_1529,N_497,In_1901);
xnor U1530 (N_1530,N_983,In_1059);
xor U1531 (N_1531,N_715,N_527);
nor U1532 (N_1532,In_1675,N_89);
xnor U1533 (N_1533,N_760,N_869);
xnor U1534 (N_1534,N_1128,In_360);
xnor U1535 (N_1535,In_570,N_1223);
nand U1536 (N_1536,N_721,N_1192);
or U1537 (N_1537,N_1130,N_366);
or U1538 (N_1538,N_1222,N_708);
nand U1539 (N_1539,N_388,N_831);
or U1540 (N_1540,In_2475,N_816);
or U1541 (N_1541,N_1174,N_784);
or U1542 (N_1542,N_764,N_367);
nor U1543 (N_1543,N_613,In_61);
nand U1544 (N_1544,N_11,N_1126);
nor U1545 (N_1545,In_2319,N_370);
nor U1546 (N_1546,N_785,N_1225);
nand U1547 (N_1547,In_2438,N_843);
nor U1548 (N_1548,In_2104,N_761);
and U1549 (N_1549,N_737,In_1076);
and U1550 (N_1550,N_1162,N_896);
xor U1551 (N_1551,N_704,In_1209);
or U1552 (N_1552,N_860,N_1012);
xor U1553 (N_1553,In_291,N_1247);
nor U1554 (N_1554,In_76,N_349);
nor U1555 (N_1555,N_377,In_1222);
xnor U1556 (N_1556,N_1155,In_2212);
and U1557 (N_1557,N_380,N_543);
xnor U1558 (N_1558,N_1060,N_325);
or U1559 (N_1559,In_40,N_750);
xnor U1560 (N_1560,In_38,N_828);
xnor U1561 (N_1561,N_488,N_713);
xnor U1562 (N_1562,N_1014,N_1144);
xor U1563 (N_1563,In_374,N_777);
nand U1564 (N_1564,In_739,N_1018);
and U1565 (N_1565,N_1232,N_849);
and U1566 (N_1566,In_221,In_1667);
xor U1567 (N_1567,N_113,In_1601);
nand U1568 (N_1568,N_900,N_846);
or U1569 (N_1569,In_603,In_473);
and U1570 (N_1570,N_652,N_862);
nand U1571 (N_1571,N_642,N_1180);
nand U1572 (N_1572,N_910,N_707);
nand U1573 (N_1573,In_571,N_797);
nor U1574 (N_1574,In_2376,N_1110);
nor U1575 (N_1575,In_882,N_1108);
nor U1576 (N_1576,N_598,N_1019);
xor U1577 (N_1577,N_1042,In_1103);
nand U1578 (N_1578,N_486,In_686);
and U1579 (N_1579,In_2448,In_1467);
and U1580 (N_1580,N_593,N_889);
nor U1581 (N_1581,N_808,In_835);
nand U1582 (N_1582,N_39,N_1070);
nand U1583 (N_1583,In_2482,N_1067);
nor U1584 (N_1584,In_364,N_998);
and U1585 (N_1585,N_925,In_2186);
nor U1586 (N_1586,In_2007,In_817);
nor U1587 (N_1587,In_1470,N_1201);
nand U1588 (N_1588,N_980,In_2397);
and U1589 (N_1589,N_873,N_1100);
nand U1590 (N_1590,N_143,N_1106);
or U1591 (N_1591,N_71,In_2274);
or U1592 (N_1592,N_942,N_453);
and U1593 (N_1593,In_1861,In_627);
xnor U1594 (N_1594,N_744,In_962);
or U1595 (N_1595,In_705,N_747);
xor U1596 (N_1596,In_980,N_815);
xnor U1597 (N_1597,N_933,N_381);
xnor U1598 (N_1598,N_895,N_689);
nor U1599 (N_1599,N_901,In_168);
nand U1600 (N_1600,N_1153,N_4);
and U1601 (N_1601,N_817,N_748);
nand U1602 (N_1602,N_591,In_607);
nand U1603 (N_1603,N_693,N_1214);
and U1604 (N_1604,N_271,N_823);
nand U1605 (N_1605,N_1043,In_1413);
and U1606 (N_1606,N_523,In_753);
xnor U1607 (N_1607,In_1562,N_810);
xor U1608 (N_1608,In_1856,N_1226);
xnor U1609 (N_1609,In_2139,N_1243);
nand U1610 (N_1610,In_1548,N_283);
nand U1611 (N_1611,In_2037,N_1025);
xnor U1612 (N_1612,N_29,N_997);
xor U1613 (N_1613,N_522,N_1173);
and U1614 (N_1614,N_909,In_1583);
nand U1615 (N_1615,In_899,N_1148);
nand U1616 (N_1616,N_974,In_1485);
xnor U1617 (N_1617,N_724,N_94);
or U1618 (N_1618,In_2255,In_1563);
or U1619 (N_1619,In_1579,N_1065);
xnor U1620 (N_1620,N_1080,In_2211);
nor U1621 (N_1621,In_936,In_67);
and U1622 (N_1622,N_847,N_524);
nand U1623 (N_1623,N_758,In_1905);
nand U1624 (N_1624,In_1124,In_904);
nand U1625 (N_1625,In_1877,N_1217);
or U1626 (N_1626,In_824,N_917);
nand U1627 (N_1627,N_1142,N_174);
and U1628 (N_1628,N_1116,N_1176);
nor U1629 (N_1629,In_2084,N_1238);
and U1630 (N_1630,N_950,N_985);
and U1631 (N_1631,N_1197,N_1039);
nor U1632 (N_1632,N_539,In_1343);
or U1633 (N_1633,N_805,N_1109);
xnor U1634 (N_1634,In_2047,In_2109);
and U1635 (N_1635,In_195,N_421);
or U1636 (N_1636,N_228,In_716);
nand U1637 (N_1637,N_1051,In_2340);
and U1638 (N_1638,N_848,N_243);
xnor U1639 (N_1639,In_1415,N_475);
and U1640 (N_1640,In_2108,N_444);
xnor U1641 (N_1641,N_1213,N_338);
xnor U1642 (N_1642,N_921,In_1360);
nor U1643 (N_1643,In_191,N_926);
xor U1644 (N_1644,N_1139,N_938);
xor U1645 (N_1645,N_778,N_323);
xor U1646 (N_1646,N_548,N_1066);
nor U1647 (N_1647,N_1077,In_812);
nand U1648 (N_1648,N_936,N_984);
xnor U1649 (N_1649,N_779,N_1134);
and U1650 (N_1650,In_2365,N_200);
or U1651 (N_1651,In_831,In_1344);
and U1652 (N_1652,N_106,In_2024);
nor U1653 (N_1653,In_688,N_45);
or U1654 (N_1654,N_1118,N_1103);
xor U1655 (N_1655,In_1953,In_2263);
xor U1656 (N_1656,N_1003,In_564);
xnor U1657 (N_1657,N_198,N_1044);
or U1658 (N_1658,N_684,N_1145);
and U1659 (N_1659,N_773,In_676);
and U1660 (N_1660,N_15,N_118);
or U1661 (N_1661,In_1117,In_913);
nor U1662 (N_1662,N_235,N_999);
or U1663 (N_1663,N_679,N_1020);
nor U1664 (N_1664,In_212,N_1008);
nand U1665 (N_1665,In_680,In_1260);
nand U1666 (N_1666,N_1024,In_850);
xor U1667 (N_1667,N_1089,N_168);
nor U1668 (N_1668,In_633,N_965);
nand U1669 (N_1669,N_34,In_2096);
and U1670 (N_1670,In_706,N_1212);
xnor U1671 (N_1671,In_461,In_363);
nor U1672 (N_1672,N_1195,In_1032);
and U1673 (N_1673,N_31,N_1054);
xor U1674 (N_1674,In_1337,N_1227);
nor U1675 (N_1675,N_687,N_1143);
xor U1676 (N_1676,N_699,In_207);
nand U1677 (N_1677,N_990,In_215);
or U1678 (N_1678,N_531,N_590);
nor U1679 (N_1679,N_741,N_300);
or U1680 (N_1680,N_433,In_315);
and U1681 (N_1681,In_1661,N_959);
or U1682 (N_1682,In_934,In_1907);
xnor U1683 (N_1683,N_770,N_863);
nand U1684 (N_1684,N_881,In_717);
nor U1685 (N_1685,In_1484,N_880);
xor U1686 (N_1686,In_2391,In_411);
nor U1687 (N_1687,N_763,N_654);
nor U1688 (N_1688,N_1093,N_1032);
nor U1689 (N_1689,In_391,In_1691);
and U1690 (N_1690,N_1146,N_1236);
and U1691 (N_1691,N_158,N_1075);
xor U1692 (N_1692,N_1199,N_717);
and U1693 (N_1693,N_1006,N_801);
and U1694 (N_1694,N_1175,In_1368);
or U1695 (N_1695,N_244,In_677);
xor U1696 (N_1696,N_714,N_864);
nand U1697 (N_1697,In_2408,In_1659);
xnor U1698 (N_1698,N_842,N_561);
nand U1699 (N_1699,N_533,In_2284);
xor U1700 (N_1700,N_875,N_1163);
nand U1701 (N_1701,N_1200,In_829);
or U1702 (N_1702,In_678,N_735);
xor U1703 (N_1703,N_955,N_1210);
and U1704 (N_1704,N_649,In_1569);
nand U1705 (N_1705,N_911,N_839);
or U1706 (N_1706,N_389,N_376);
xor U1707 (N_1707,N_902,N_1178);
nor U1708 (N_1708,N_330,N_1207);
xnor U1709 (N_1709,N_972,N_1218);
nand U1710 (N_1710,In_263,In_123);
or U1711 (N_1711,N_1091,N_1102);
nor U1712 (N_1712,N_643,In_55);
or U1713 (N_1713,N_400,N_866);
or U1714 (N_1714,N_807,N_1098);
nor U1715 (N_1715,N_594,In_197);
and U1716 (N_1716,In_1805,N_564);
xnor U1717 (N_1717,N_698,N_1050);
nand U1718 (N_1718,In_1478,N_1129);
nor U1719 (N_1719,N_508,N_943);
and U1720 (N_1720,N_1184,N_792);
nand U1721 (N_1721,N_1000,N_1198);
nand U1722 (N_1722,N_319,N_212);
xor U1723 (N_1723,N_474,N_61);
and U1724 (N_1724,N_1168,N_1094);
xnor U1725 (N_1725,In_1104,N_1246);
or U1726 (N_1726,N_5,In_1787);
nand U1727 (N_1727,In_2444,In_2413);
nor U1728 (N_1728,N_131,N_795);
nand U1729 (N_1729,In_312,In_511);
nor U1730 (N_1730,In_459,In_2179);
xnor U1731 (N_1731,In_1265,In_313);
or U1732 (N_1732,N_1131,N_426);
xnor U1733 (N_1733,In_2398,In_1808);
or U1734 (N_1734,N_742,N_1016);
or U1735 (N_1735,N_187,N_1154);
or U1736 (N_1736,N_1224,In_576);
nor U1737 (N_1737,N_628,N_1231);
nor U1738 (N_1738,N_916,N_638);
nor U1739 (N_1739,N_850,In_543);
nand U1740 (N_1740,N_701,In_113);
and U1741 (N_1741,N_728,N_1233);
and U1742 (N_1742,N_799,N_719);
or U1743 (N_1743,In_1205,N_427);
xnor U1744 (N_1744,N_179,N_908);
nor U1745 (N_1745,In_1328,N_1124);
and U1746 (N_1746,In_1779,N_1182);
nor U1747 (N_1747,N_1193,In_1880);
xor U1748 (N_1748,In_2240,N_1073);
nor U1749 (N_1749,In_410,In_98);
and U1750 (N_1750,In_1107,N_995);
xor U1751 (N_1751,N_1206,In_505);
or U1752 (N_1752,N_769,N_671);
or U1753 (N_1753,In_1755,N_888);
xor U1754 (N_1754,N_1022,N_321);
nand U1755 (N_1755,N_631,In_178);
nor U1756 (N_1756,N_1040,N_1099);
or U1757 (N_1757,N_1248,N_969);
or U1758 (N_1758,In_1620,N_265);
and U1759 (N_1759,In_218,N_672);
and U1760 (N_1760,N_766,In_865);
and U1761 (N_1761,N_1005,N_1133);
xnor U1762 (N_1762,N_505,N_865);
xnor U1763 (N_1763,N_1220,In_2153);
xor U1764 (N_1764,N_809,N_606);
and U1765 (N_1765,N_836,N_1189);
xnor U1766 (N_1766,In_1829,In_1350);
nor U1767 (N_1767,N_1208,N_354);
nor U1768 (N_1768,N_927,N_53);
nand U1769 (N_1769,N_1237,N_1013);
or U1770 (N_1770,In_2176,N_1045);
or U1771 (N_1771,N_756,N_702);
nand U1772 (N_1772,N_1033,N_753);
and U1773 (N_1773,N_1140,N_646);
and U1774 (N_1774,N_683,N_906);
xnor U1775 (N_1775,N_876,N_607);
and U1776 (N_1776,N_970,N_688);
and U1777 (N_1777,N_610,N_774);
and U1778 (N_1778,N_459,N_723);
nand U1779 (N_1779,N_918,N_835);
nor U1780 (N_1780,N_250,N_657);
and U1781 (N_1781,N_464,In_805);
xor U1782 (N_1782,N_685,N_285);
xor U1783 (N_1783,N_986,N_1240);
nand U1784 (N_1784,N_138,N_1061);
and U1785 (N_1785,N_455,In_164);
xor U1786 (N_1786,In_568,N_718);
and U1787 (N_1787,In_675,In_522);
and U1788 (N_1788,N_800,In_1920);
xor U1789 (N_1789,In_890,N_302);
or U1790 (N_1790,N_820,N_460);
xor U1791 (N_1791,N_1117,N_636);
and U1792 (N_1792,N_1072,N_532);
nor U1793 (N_1793,In_1012,In_978);
nor U1794 (N_1794,N_1241,N_1170);
nor U1795 (N_1795,N_40,N_280);
xnor U1796 (N_1796,N_930,N_793);
xor U1797 (N_1797,N_1171,In_1454);
or U1798 (N_1798,In_193,In_894);
nor U1799 (N_1799,N_729,In_1592);
nor U1800 (N_1800,N_802,N_754);
xnor U1801 (N_1801,In_591,N_883);
nor U1802 (N_1802,In_1285,In_685);
and U1803 (N_1803,In_196,N_891);
nor U1804 (N_1804,In_541,N_1150);
or U1805 (N_1805,N_1063,In_2225);
nand U1806 (N_1806,N_1074,N_957);
xnor U1807 (N_1807,N_1169,In_2256);
and U1808 (N_1808,In_475,N_855);
xor U1809 (N_1809,In_1074,N_691);
and U1810 (N_1810,N_765,N_861);
or U1811 (N_1811,N_580,N_1068);
nand U1812 (N_1812,N_1009,In_926);
nand U1813 (N_1813,In_1833,N_705);
xor U1814 (N_1814,N_1204,N_277);
and U1815 (N_1815,N_615,N_788);
and U1816 (N_1816,In_396,N_151);
nand U1817 (N_1817,In_1086,N_826);
nand U1818 (N_1818,In_1206,In_1595);
xor U1819 (N_1819,N_897,N_1071);
or U1820 (N_1820,N_1001,N_789);
nor U1821 (N_1821,In_176,N_306);
and U1822 (N_1822,N_827,In_2132);
nor U1823 (N_1823,N_949,N_666);
xnor U1824 (N_1824,N_566,N_1136);
and U1825 (N_1825,N_1107,In_1697);
xnor U1826 (N_1826,In_240,In_245);
and U1827 (N_1827,N_648,N_851);
and U1828 (N_1828,In_2257,N_1015);
nand U1829 (N_1829,In_258,N_892);
xor U1830 (N_1830,In_1179,N_1115);
nor U1831 (N_1831,N_759,N_814);
xnor U1832 (N_1832,N_712,N_825);
and U1833 (N_1833,N_1156,N_924);
or U1834 (N_1834,N_874,N_882);
xor U1835 (N_1835,N_731,In_456);
nor U1836 (N_1836,In_1404,N_1151);
nand U1837 (N_1837,N_641,N_1092);
and U1838 (N_1838,N_697,N_490);
nor U1839 (N_1839,N_716,N_1048);
nor U1840 (N_1840,N_1245,N_832);
or U1841 (N_1841,N_952,In_44);
xnor U1842 (N_1842,In_1314,N_1026);
and U1843 (N_1843,In_2353,N_1112);
xnor U1844 (N_1844,In_1499,N_1235);
xnor U1845 (N_1845,N_746,In_1095);
and U1846 (N_1846,N_700,In_2063);
and U1847 (N_1847,In_1122,In_1774);
nor U1848 (N_1848,N_640,In_990);
and U1849 (N_1849,N_830,In_861);
xor U1850 (N_1850,In_2182,N_445);
xor U1851 (N_1851,N_821,N_7);
nor U1852 (N_1852,In_1848,N_1121);
nor U1853 (N_1853,In_2297,N_988);
nand U1854 (N_1854,N_1095,N_853);
nor U1855 (N_1855,N_42,N_1160);
and U1856 (N_1856,N_245,N_996);
xor U1857 (N_1857,N_429,N_894);
xnor U1858 (N_1858,N_1085,N_819);
nor U1859 (N_1859,N_940,In_357);
nor U1860 (N_1860,N_757,N_1185);
or U1861 (N_1861,N_954,In_1429);
nor U1862 (N_1862,N_520,N_1057);
nor U1863 (N_1863,N_772,N_987);
nor U1864 (N_1864,N_664,N_667);
nand U1865 (N_1865,In_2451,N_845);
or U1866 (N_1866,N_676,N_1086);
nor U1867 (N_1867,In_1820,In_1932);
nor U1868 (N_1868,N_1053,In_2205);
and U1869 (N_1869,N_686,In_251);
xnor U1870 (N_1870,N_1078,N_653);
nand U1871 (N_1871,N_414,N_898);
nand U1872 (N_1872,In_643,In_160);
and U1873 (N_1873,N_973,N_838);
and U1874 (N_1874,In_1775,N_923);
nor U1875 (N_1875,N_1473,N_1599);
and U1876 (N_1876,N_1554,N_1639);
xnor U1877 (N_1877,N_1729,N_1764);
nand U1878 (N_1878,N_1714,N_1534);
and U1879 (N_1879,N_1442,N_1389);
nand U1880 (N_1880,N_1564,N_1835);
nor U1881 (N_1881,N_1438,N_1316);
nor U1882 (N_1882,N_1850,N_1419);
xor U1883 (N_1883,N_1526,N_1431);
and U1884 (N_1884,N_1254,N_1313);
or U1885 (N_1885,N_1331,N_1754);
or U1886 (N_1886,N_1642,N_1339);
or U1887 (N_1887,N_1761,N_1620);
or U1888 (N_1888,N_1377,N_1359);
nor U1889 (N_1889,N_1463,N_1700);
and U1890 (N_1890,N_1420,N_1383);
or U1891 (N_1891,N_1696,N_1371);
nand U1892 (N_1892,N_1296,N_1660);
or U1893 (N_1893,N_1776,N_1657);
xor U1894 (N_1894,N_1386,N_1605);
and U1895 (N_1895,N_1816,N_1509);
nor U1896 (N_1896,N_1868,N_1464);
nor U1897 (N_1897,N_1460,N_1810);
xnor U1898 (N_1898,N_1662,N_1822);
xnor U1899 (N_1899,N_1370,N_1833);
xnor U1900 (N_1900,N_1784,N_1646);
or U1901 (N_1901,N_1837,N_1306);
xnor U1902 (N_1902,N_1797,N_1286);
or U1903 (N_1903,N_1786,N_1732);
or U1904 (N_1904,N_1256,N_1703);
nand U1905 (N_1905,N_1427,N_1796);
nor U1906 (N_1906,N_1399,N_1602);
nor U1907 (N_1907,N_1329,N_1505);
xnor U1908 (N_1908,N_1302,N_1622);
nand U1909 (N_1909,N_1255,N_1684);
nand U1910 (N_1910,N_1475,N_1310);
or U1911 (N_1911,N_1624,N_1576);
nor U1912 (N_1912,N_1317,N_1635);
xor U1913 (N_1913,N_1452,N_1756);
xor U1914 (N_1914,N_1731,N_1297);
nand U1915 (N_1915,N_1841,N_1767);
or U1916 (N_1916,N_1529,N_1572);
or U1917 (N_1917,N_1577,N_1437);
nand U1918 (N_1918,N_1787,N_1445);
nand U1919 (N_1919,N_1493,N_1395);
nor U1920 (N_1920,N_1540,N_1533);
and U1921 (N_1921,N_1504,N_1798);
nand U1922 (N_1922,N_1697,N_1677);
nor U1923 (N_1923,N_1503,N_1280);
nor U1924 (N_1924,N_1544,N_1751);
nand U1925 (N_1925,N_1406,N_1332);
nand U1926 (N_1926,N_1461,N_1632);
xor U1927 (N_1927,N_1330,N_1869);
xnor U1928 (N_1928,N_1573,N_1644);
or U1929 (N_1929,N_1307,N_1670);
nor U1930 (N_1930,N_1708,N_1396);
or U1931 (N_1931,N_1552,N_1318);
and U1932 (N_1932,N_1537,N_1855);
nor U1933 (N_1933,N_1748,N_1785);
and U1934 (N_1934,N_1768,N_1511);
and U1935 (N_1935,N_1827,N_1518);
nand U1936 (N_1936,N_1823,N_1749);
xor U1937 (N_1937,N_1268,N_1309);
nor U1938 (N_1938,N_1421,N_1365);
nor U1939 (N_1939,N_1337,N_1600);
xor U1940 (N_1940,N_1272,N_1556);
nor U1941 (N_1941,N_1707,N_1536);
nor U1942 (N_1942,N_1448,N_1400);
xnor U1943 (N_1943,N_1303,N_1342);
nor U1944 (N_1944,N_1580,N_1857);
xor U1945 (N_1945,N_1683,N_1375);
nor U1946 (N_1946,N_1560,N_1496);
nand U1947 (N_1947,N_1704,N_1671);
nor U1948 (N_1948,N_1575,N_1736);
and U1949 (N_1949,N_1746,N_1269);
and U1950 (N_1950,N_1369,N_1451);
xnor U1951 (N_1951,N_1291,N_1539);
nor U1952 (N_1952,N_1282,N_1743);
and U1953 (N_1953,N_1251,N_1739);
nor U1954 (N_1954,N_1488,N_1323);
xnor U1955 (N_1955,N_1804,N_1727);
or U1956 (N_1956,N_1257,N_1393);
xor U1957 (N_1957,N_1565,N_1742);
xor U1958 (N_1958,N_1434,N_1324);
nand U1959 (N_1959,N_1410,N_1344);
nand U1960 (N_1960,N_1631,N_1470);
xor U1961 (N_1961,N_1363,N_1347);
nor U1962 (N_1962,N_1333,N_1455);
nor U1963 (N_1963,N_1312,N_1740);
nand U1964 (N_1964,N_1718,N_1640);
and U1965 (N_1965,N_1374,N_1450);
nand U1966 (N_1966,N_1555,N_1681);
nor U1967 (N_1967,N_1766,N_1354);
xor U1968 (N_1968,N_1724,N_1801);
nor U1969 (N_1969,N_1382,N_1691);
xor U1970 (N_1970,N_1710,N_1528);
and U1971 (N_1971,N_1426,N_1259);
nand U1972 (N_1972,N_1569,N_1356);
and U1973 (N_1973,N_1826,N_1474);
xor U1974 (N_1974,N_1527,N_1870);
or U1975 (N_1975,N_1638,N_1851);
nor U1976 (N_1976,N_1430,N_1659);
xor U1977 (N_1977,N_1424,N_1672);
nor U1978 (N_1978,N_1562,N_1558);
and U1979 (N_1979,N_1828,N_1489);
and U1980 (N_1980,N_1583,N_1561);
xnor U1981 (N_1981,N_1838,N_1779);
and U1982 (N_1982,N_1874,N_1679);
nand U1983 (N_1983,N_1295,N_1721);
nor U1984 (N_1984,N_1627,N_1531);
or U1985 (N_1985,N_1597,N_1458);
xor U1986 (N_1986,N_1601,N_1871);
or U1987 (N_1987,N_1336,N_1477);
xor U1988 (N_1988,N_1520,N_1654);
or U1989 (N_1989,N_1772,N_1262);
xnor U1990 (N_1990,N_1692,N_1701);
nand U1991 (N_1991,N_1522,N_1472);
and U1992 (N_1992,N_1791,N_1273);
and U1993 (N_1993,N_1405,N_1865);
or U1994 (N_1994,N_1446,N_1608);
xor U1995 (N_1995,N_1340,N_1765);
xnor U1996 (N_1996,N_1319,N_1849);
nand U1997 (N_1997,N_1719,N_1480);
and U1998 (N_1998,N_1250,N_1546);
or U1999 (N_1999,N_1471,N_1422);
or U2000 (N_2000,N_1266,N_1780);
or U2001 (N_2001,N_1686,N_1858);
or U2002 (N_2002,N_1532,N_1832);
xnor U2003 (N_2003,N_1275,N_1397);
xnor U2004 (N_2004,N_1469,N_1416);
or U2005 (N_2005,N_1497,N_1360);
nor U2006 (N_2006,N_1549,N_1637);
xnor U2007 (N_2007,N_1320,N_1521);
and U2008 (N_2008,N_1690,N_1843);
nand U2009 (N_2009,N_1428,N_1315);
and U2010 (N_2010,N_1283,N_1813);
nand U2011 (N_2011,N_1769,N_1584);
and U2012 (N_2012,N_1479,N_1423);
or U2013 (N_2013,N_1321,N_1260);
nor U2014 (N_2014,N_1633,N_1346);
xor U2015 (N_2015,N_1550,N_1680);
nand U2016 (N_2016,N_1433,N_1304);
nand U2017 (N_2017,N_1694,N_1789);
nand U2018 (N_2018,N_1376,N_1563);
and U2019 (N_2019,N_1278,N_1634);
nand U2020 (N_2020,N_1414,N_1417);
nand U2021 (N_2021,N_1621,N_1587);
nand U2022 (N_2022,N_1723,N_1459);
xor U2023 (N_2023,N_1398,N_1567);
nor U2024 (N_2024,N_1799,N_1844);
or U2025 (N_2025,N_1808,N_1378);
or U2026 (N_2026,N_1263,N_1656);
nand U2027 (N_2027,N_1817,N_1334);
xnor U2028 (N_2028,N_1792,N_1643);
nand U2029 (N_2029,N_1741,N_1343);
and U2030 (N_2030,N_1593,N_1326);
and U2031 (N_2031,N_1525,N_1862);
nand U2032 (N_2032,N_1391,N_1647);
nand U2033 (N_2033,N_1863,N_1778);
nor U2034 (N_2034,N_1650,N_1722);
xor U2035 (N_2035,N_1839,N_1847);
nor U2036 (N_2036,N_1325,N_1341);
and U2037 (N_2037,N_1372,N_1502);
nor U2038 (N_2038,N_1454,N_1384);
xnor U2039 (N_2039,N_1604,N_1803);
xnor U2040 (N_2040,N_1538,N_1289);
and U2041 (N_2041,N_1628,N_1611);
or U2042 (N_2042,N_1411,N_1689);
xnor U2043 (N_2043,N_1665,N_1308);
and U2044 (N_2044,N_1355,N_1500);
and U2045 (N_2045,N_1253,N_1759);
nor U2046 (N_2046,N_1335,N_1413);
xnor U2047 (N_2047,N_1818,N_1501);
nand U2048 (N_2048,N_1294,N_1693);
and U2049 (N_2049,N_1629,N_1802);
or U2050 (N_2050,N_1793,N_1814);
or U2051 (N_2051,N_1606,N_1588);
nor U2052 (N_2052,N_1351,N_1733);
xor U2053 (N_2053,N_1812,N_1566);
nand U2054 (N_2054,N_1506,N_1831);
nand U2055 (N_2055,N_1626,N_1436);
and U2056 (N_2056,N_1492,N_1735);
nand U2057 (N_2057,N_1571,N_1425);
nand U2058 (N_2058,N_1578,N_1774);
xnor U2059 (N_2059,N_1311,N_1512);
and U2060 (N_2060,N_1846,N_1598);
xor U2061 (N_2061,N_1364,N_1491);
xor U2062 (N_2062,N_1595,N_1866);
nor U2063 (N_2063,N_1401,N_1668);
nand U2064 (N_2064,N_1547,N_1495);
or U2065 (N_2065,N_1819,N_1806);
and U2066 (N_2066,N_1292,N_1702);
nor U2067 (N_2067,N_1805,N_1353);
nand U2068 (N_2068,N_1664,N_1387);
nand U2069 (N_2069,N_1392,N_1581);
xnor U2070 (N_2070,N_1607,N_1777);
nand U2071 (N_2071,N_1585,N_1623);
xor U2072 (N_2072,N_1568,N_1687);
xor U2073 (N_2073,N_1698,N_1782);
or U2074 (N_2074,N_1695,N_1730);
and U2075 (N_2075,N_1612,N_1551);
nor U2076 (N_2076,N_1379,N_1390);
xor U2077 (N_2077,N_1755,N_1557);
or U2078 (N_2078,N_1468,N_1781);
and U2079 (N_2079,N_1328,N_1630);
xor U2080 (N_2080,N_1720,N_1747);
nand U2081 (N_2081,N_1264,N_1845);
nand U2082 (N_2082,N_1441,N_1852);
xor U2083 (N_2083,N_1271,N_1494);
nand U2084 (N_2084,N_1825,N_1610);
xor U2085 (N_2085,N_1834,N_1590);
and U2086 (N_2086,N_1699,N_1728);
and U2087 (N_2087,N_1788,N_1745);
and U2088 (N_2088,N_1443,N_1367);
or U2089 (N_2089,N_1478,N_1658);
or U2090 (N_2090,N_1675,N_1465);
and U2091 (N_2091,N_1820,N_1449);
or U2092 (N_2092,N_1842,N_1873);
nor U2093 (N_2093,N_1456,N_1362);
xnor U2094 (N_2094,N_1617,N_1807);
or U2095 (N_2095,N_1542,N_1481);
and U2096 (N_2096,N_1361,N_1553);
nand U2097 (N_2097,N_1327,N_1574);
nor U2098 (N_2098,N_1403,N_1366);
xor U2099 (N_2099,N_1457,N_1757);
xnor U2100 (N_2100,N_1795,N_1678);
nand U2101 (N_2101,N_1655,N_1661);
xor U2102 (N_2102,N_1439,N_1758);
nand U2103 (N_2103,N_1482,N_1763);
nand U2104 (N_2104,N_1523,N_1407);
nor U2105 (N_2105,N_1815,N_1811);
nand U2106 (N_2106,N_1753,N_1636);
and U2107 (N_2107,N_1252,N_1760);
xor U2108 (N_2108,N_1408,N_1618);
xor U2109 (N_2109,N_1284,N_1653);
nor U2110 (N_2110,N_1669,N_1609);
nand U2111 (N_2111,N_1840,N_1388);
nand U2112 (N_2112,N_1486,N_1548);
xnor U2113 (N_2113,N_1867,N_1864);
or U2114 (N_2114,N_1288,N_1510);
nand U2115 (N_2115,N_1582,N_1715);
nand U2116 (N_2116,N_1649,N_1591);
nor U2117 (N_2117,N_1594,N_1619);
nor U2118 (N_2118,N_1373,N_1444);
or U2119 (N_2119,N_1716,N_1645);
nand U2120 (N_2120,N_1872,N_1349);
nor U2121 (N_2121,N_1380,N_1734);
nor U2122 (N_2122,N_1385,N_1290);
or U2123 (N_2123,N_1462,N_1499);
nor U2124 (N_2124,N_1648,N_1281);
xor U2125 (N_2125,N_1752,N_1824);
nor U2126 (N_2126,N_1614,N_1484);
and U2127 (N_2127,N_1712,N_1530);
xnor U2128 (N_2128,N_1412,N_1579);
and U2129 (N_2129,N_1652,N_1314);
and U2130 (N_2130,N_1616,N_1485);
nor U2131 (N_2131,N_1770,N_1545);
xor U2132 (N_2132,N_1592,N_1663);
or U2133 (N_2133,N_1498,N_1709);
xnor U2134 (N_2134,N_1322,N_1513);
or U2135 (N_2135,N_1570,N_1711);
nor U2136 (N_2136,N_1404,N_1809);
or U2137 (N_2137,N_1771,N_1535);
nand U2138 (N_2138,N_1685,N_1358);
nor U2139 (N_2139,N_1524,N_1666);
xor U2140 (N_2140,N_1762,N_1853);
nor U2141 (N_2141,N_1453,N_1298);
and U2142 (N_2142,N_1267,N_1368);
xnor U2143 (N_2143,N_1829,N_1277);
and U2144 (N_2144,N_1507,N_1300);
nor U2145 (N_2145,N_1673,N_1466);
and U2146 (N_2146,N_1790,N_1514);
xnor U2147 (N_2147,N_1848,N_1402);
or U2148 (N_2148,N_1287,N_1651);
or U2149 (N_2149,N_1490,N_1350);
or U2150 (N_2150,N_1483,N_1276);
nor U2151 (N_2151,N_1856,N_1299);
or U2152 (N_2152,N_1476,N_1674);
or U2153 (N_2153,N_1861,N_1625);
or U2154 (N_2154,N_1738,N_1800);
nor U2155 (N_2155,N_1821,N_1338);
and U2156 (N_2156,N_1345,N_1261);
or U2157 (N_2157,N_1744,N_1301);
or U2158 (N_2158,N_1429,N_1750);
xnor U2159 (N_2159,N_1596,N_1258);
nand U2160 (N_2160,N_1541,N_1706);
nor U2161 (N_2161,N_1682,N_1418);
or U2162 (N_2162,N_1836,N_1381);
nand U2163 (N_2163,N_1517,N_1860);
and U2164 (N_2164,N_1265,N_1676);
nor U2165 (N_2165,N_1794,N_1516);
nand U2166 (N_2166,N_1352,N_1519);
or U2167 (N_2167,N_1603,N_1667);
xnor U2168 (N_2168,N_1357,N_1717);
or U2169 (N_2169,N_1274,N_1285);
or U2170 (N_2170,N_1775,N_1559);
or U2171 (N_2171,N_1543,N_1725);
xnor U2172 (N_2172,N_1487,N_1415);
nand U2173 (N_2173,N_1589,N_1508);
or U2174 (N_2174,N_1713,N_1394);
nor U2175 (N_2175,N_1705,N_1783);
and U2176 (N_2176,N_1447,N_1773);
nor U2177 (N_2177,N_1726,N_1467);
or U2178 (N_2178,N_1854,N_1293);
and U2179 (N_2179,N_1515,N_1688);
xnor U2180 (N_2180,N_1279,N_1432);
nor U2181 (N_2181,N_1830,N_1613);
nor U2182 (N_2182,N_1409,N_1615);
xor U2183 (N_2183,N_1440,N_1641);
xor U2184 (N_2184,N_1737,N_1859);
nor U2185 (N_2185,N_1270,N_1348);
and U2186 (N_2186,N_1435,N_1305);
and U2187 (N_2187,N_1586,N_1319);
or U2188 (N_2188,N_1694,N_1559);
or U2189 (N_2189,N_1275,N_1846);
xor U2190 (N_2190,N_1466,N_1359);
xor U2191 (N_2191,N_1614,N_1686);
and U2192 (N_2192,N_1501,N_1342);
or U2193 (N_2193,N_1684,N_1507);
xnor U2194 (N_2194,N_1589,N_1832);
and U2195 (N_2195,N_1290,N_1493);
or U2196 (N_2196,N_1712,N_1544);
and U2197 (N_2197,N_1469,N_1549);
xnor U2198 (N_2198,N_1726,N_1694);
nand U2199 (N_2199,N_1869,N_1848);
xor U2200 (N_2200,N_1583,N_1445);
nor U2201 (N_2201,N_1603,N_1734);
and U2202 (N_2202,N_1628,N_1576);
nor U2203 (N_2203,N_1358,N_1594);
nor U2204 (N_2204,N_1451,N_1518);
or U2205 (N_2205,N_1440,N_1432);
nand U2206 (N_2206,N_1366,N_1549);
nand U2207 (N_2207,N_1395,N_1631);
nor U2208 (N_2208,N_1524,N_1328);
or U2209 (N_2209,N_1360,N_1329);
or U2210 (N_2210,N_1315,N_1774);
or U2211 (N_2211,N_1684,N_1775);
nand U2212 (N_2212,N_1505,N_1465);
and U2213 (N_2213,N_1331,N_1500);
xnor U2214 (N_2214,N_1850,N_1436);
nand U2215 (N_2215,N_1304,N_1806);
xnor U2216 (N_2216,N_1587,N_1686);
and U2217 (N_2217,N_1679,N_1464);
and U2218 (N_2218,N_1840,N_1592);
xor U2219 (N_2219,N_1731,N_1446);
and U2220 (N_2220,N_1867,N_1556);
and U2221 (N_2221,N_1345,N_1386);
nor U2222 (N_2222,N_1570,N_1553);
nor U2223 (N_2223,N_1512,N_1408);
or U2224 (N_2224,N_1782,N_1523);
xnor U2225 (N_2225,N_1431,N_1695);
or U2226 (N_2226,N_1860,N_1808);
or U2227 (N_2227,N_1649,N_1613);
or U2228 (N_2228,N_1864,N_1379);
nor U2229 (N_2229,N_1798,N_1484);
nand U2230 (N_2230,N_1741,N_1408);
xor U2231 (N_2231,N_1823,N_1710);
xnor U2232 (N_2232,N_1291,N_1498);
and U2233 (N_2233,N_1773,N_1571);
xor U2234 (N_2234,N_1308,N_1519);
and U2235 (N_2235,N_1733,N_1366);
or U2236 (N_2236,N_1673,N_1484);
nor U2237 (N_2237,N_1337,N_1424);
nor U2238 (N_2238,N_1812,N_1392);
xor U2239 (N_2239,N_1505,N_1753);
and U2240 (N_2240,N_1695,N_1775);
and U2241 (N_2241,N_1340,N_1402);
xor U2242 (N_2242,N_1687,N_1681);
and U2243 (N_2243,N_1528,N_1347);
xnor U2244 (N_2244,N_1505,N_1773);
nand U2245 (N_2245,N_1335,N_1574);
or U2246 (N_2246,N_1714,N_1513);
nand U2247 (N_2247,N_1410,N_1862);
xor U2248 (N_2248,N_1793,N_1447);
xnor U2249 (N_2249,N_1849,N_1431);
and U2250 (N_2250,N_1318,N_1467);
or U2251 (N_2251,N_1304,N_1268);
nor U2252 (N_2252,N_1703,N_1848);
and U2253 (N_2253,N_1753,N_1569);
nand U2254 (N_2254,N_1523,N_1465);
xor U2255 (N_2255,N_1374,N_1460);
nor U2256 (N_2256,N_1696,N_1619);
and U2257 (N_2257,N_1761,N_1683);
or U2258 (N_2258,N_1820,N_1341);
nand U2259 (N_2259,N_1307,N_1388);
nand U2260 (N_2260,N_1605,N_1575);
or U2261 (N_2261,N_1680,N_1427);
xor U2262 (N_2262,N_1638,N_1495);
nand U2263 (N_2263,N_1436,N_1762);
xor U2264 (N_2264,N_1313,N_1748);
and U2265 (N_2265,N_1503,N_1787);
or U2266 (N_2266,N_1794,N_1677);
nand U2267 (N_2267,N_1839,N_1627);
nor U2268 (N_2268,N_1585,N_1622);
nand U2269 (N_2269,N_1744,N_1861);
and U2270 (N_2270,N_1253,N_1413);
xor U2271 (N_2271,N_1733,N_1462);
nand U2272 (N_2272,N_1789,N_1870);
nand U2273 (N_2273,N_1802,N_1764);
nand U2274 (N_2274,N_1486,N_1516);
or U2275 (N_2275,N_1574,N_1606);
or U2276 (N_2276,N_1848,N_1374);
or U2277 (N_2277,N_1679,N_1809);
xor U2278 (N_2278,N_1384,N_1795);
xnor U2279 (N_2279,N_1766,N_1283);
and U2280 (N_2280,N_1491,N_1584);
nor U2281 (N_2281,N_1534,N_1872);
xnor U2282 (N_2282,N_1318,N_1263);
or U2283 (N_2283,N_1536,N_1534);
and U2284 (N_2284,N_1722,N_1648);
or U2285 (N_2285,N_1849,N_1546);
xor U2286 (N_2286,N_1455,N_1281);
xnor U2287 (N_2287,N_1544,N_1349);
nand U2288 (N_2288,N_1722,N_1749);
or U2289 (N_2289,N_1411,N_1849);
xnor U2290 (N_2290,N_1751,N_1287);
and U2291 (N_2291,N_1437,N_1806);
xnor U2292 (N_2292,N_1438,N_1470);
and U2293 (N_2293,N_1831,N_1874);
nor U2294 (N_2294,N_1454,N_1467);
xor U2295 (N_2295,N_1350,N_1633);
nor U2296 (N_2296,N_1376,N_1743);
or U2297 (N_2297,N_1872,N_1251);
nor U2298 (N_2298,N_1730,N_1281);
or U2299 (N_2299,N_1359,N_1382);
or U2300 (N_2300,N_1691,N_1815);
nand U2301 (N_2301,N_1618,N_1251);
nand U2302 (N_2302,N_1256,N_1472);
or U2303 (N_2303,N_1870,N_1681);
or U2304 (N_2304,N_1416,N_1594);
nand U2305 (N_2305,N_1305,N_1475);
xnor U2306 (N_2306,N_1332,N_1816);
xor U2307 (N_2307,N_1729,N_1753);
and U2308 (N_2308,N_1692,N_1645);
or U2309 (N_2309,N_1505,N_1831);
xnor U2310 (N_2310,N_1605,N_1496);
nor U2311 (N_2311,N_1569,N_1408);
and U2312 (N_2312,N_1575,N_1413);
xnor U2313 (N_2313,N_1869,N_1716);
nand U2314 (N_2314,N_1504,N_1430);
nor U2315 (N_2315,N_1688,N_1571);
and U2316 (N_2316,N_1552,N_1765);
or U2317 (N_2317,N_1559,N_1493);
xor U2318 (N_2318,N_1433,N_1737);
or U2319 (N_2319,N_1637,N_1797);
xor U2320 (N_2320,N_1582,N_1834);
and U2321 (N_2321,N_1386,N_1696);
and U2322 (N_2322,N_1454,N_1599);
and U2323 (N_2323,N_1390,N_1315);
nor U2324 (N_2324,N_1772,N_1731);
or U2325 (N_2325,N_1867,N_1825);
or U2326 (N_2326,N_1667,N_1262);
and U2327 (N_2327,N_1269,N_1329);
nor U2328 (N_2328,N_1320,N_1801);
and U2329 (N_2329,N_1825,N_1419);
and U2330 (N_2330,N_1659,N_1745);
xnor U2331 (N_2331,N_1624,N_1782);
nor U2332 (N_2332,N_1480,N_1636);
or U2333 (N_2333,N_1578,N_1509);
nand U2334 (N_2334,N_1291,N_1255);
and U2335 (N_2335,N_1570,N_1741);
nand U2336 (N_2336,N_1784,N_1418);
nand U2337 (N_2337,N_1781,N_1251);
or U2338 (N_2338,N_1747,N_1412);
nand U2339 (N_2339,N_1266,N_1770);
nor U2340 (N_2340,N_1421,N_1534);
or U2341 (N_2341,N_1610,N_1577);
nor U2342 (N_2342,N_1512,N_1308);
and U2343 (N_2343,N_1410,N_1760);
and U2344 (N_2344,N_1439,N_1738);
and U2345 (N_2345,N_1716,N_1695);
or U2346 (N_2346,N_1476,N_1732);
xnor U2347 (N_2347,N_1627,N_1485);
nand U2348 (N_2348,N_1674,N_1838);
or U2349 (N_2349,N_1661,N_1657);
xor U2350 (N_2350,N_1340,N_1824);
nand U2351 (N_2351,N_1279,N_1387);
xor U2352 (N_2352,N_1711,N_1709);
xnor U2353 (N_2353,N_1425,N_1814);
and U2354 (N_2354,N_1276,N_1461);
xnor U2355 (N_2355,N_1610,N_1482);
and U2356 (N_2356,N_1815,N_1648);
xor U2357 (N_2357,N_1293,N_1793);
nor U2358 (N_2358,N_1691,N_1608);
or U2359 (N_2359,N_1647,N_1407);
xor U2360 (N_2360,N_1849,N_1743);
or U2361 (N_2361,N_1586,N_1818);
or U2362 (N_2362,N_1825,N_1361);
nand U2363 (N_2363,N_1448,N_1671);
nand U2364 (N_2364,N_1295,N_1848);
or U2365 (N_2365,N_1782,N_1391);
nand U2366 (N_2366,N_1576,N_1524);
xnor U2367 (N_2367,N_1591,N_1433);
and U2368 (N_2368,N_1288,N_1577);
or U2369 (N_2369,N_1447,N_1304);
nand U2370 (N_2370,N_1746,N_1328);
and U2371 (N_2371,N_1859,N_1264);
xor U2372 (N_2372,N_1376,N_1801);
xor U2373 (N_2373,N_1832,N_1370);
nand U2374 (N_2374,N_1372,N_1850);
xor U2375 (N_2375,N_1581,N_1252);
or U2376 (N_2376,N_1527,N_1290);
nor U2377 (N_2377,N_1677,N_1630);
or U2378 (N_2378,N_1550,N_1786);
nor U2379 (N_2379,N_1285,N_1627);
and U2380 (N_2380,N_1519,N_1707);
xor U2381 (N_2381,N_1553,N_1577);
and U2382 (N_2382,N_1754,N_1633);
nor U2383 (N_2383,N_1567,N_1451);
or U2384 (N_2384,N_1645,N_1482);
and U2385 (N_2385,N_1362,N_1508);
xor U2386 (N_2386,N_1499,N_1287);
and U2387 (N_2387,N_1857,N_1385);
and U2388 (N_2388,N_1595,N_1300);
or U2389 (N_2389,N_1563,N_1626);
and U2390 (N_2390,N_1859,N_1295);
nand U2391 (N_2391,N_1688,N_1549);
or U2392 (N_2392,N_1504,N_1776);
nand U2393 (N_2393,N_1568,N_1376);
xnor U2394 (N_2394,N_1450,N_1511);
xor U2395 (N_2395,N_1531,N_1524);
xor U2396 (N_2396,N_1764,N_1809);
nor U2397 (N_2397,N_1301,N_1446);
nand U2398 (N_2398,N_1652,N_1486);
nor U2399 (N_2399,N_1341,N_1723);
or U2400 (N_2400,N_1407,N_1358);
nand U2401 (N_2401,N_1575,N_1825);
xnor U2402 (N_2402,N_1652,N_1668);
nand U2403 (N_2403,N_1358,N_1715);
nand U2404 (N_2404,N_1655,N_1795);
xor U2405 (N_2405,N_1352,N_1763);
or U2406 (N_2406,N_1724,N_1469);
and U2407 (N_2407,N_1809,N_1811);
nand U2408 (N_2408,N_1647,N_1665);
nor U2409 (N_2409,N_1332,N_1850);
nor U2410 (N_2410,N_1505,N_1619);
or U2411 (N_2411,N_1396,N_1250);
nor U2412 (N_2412,N_1841,N_1700);
nand U2413 (N_2413,N_1444,N_1461);
or U2414 (N_2414,N_1505,N_1536);
and U2415 (N_2415,N_1802,N_1394);
nand U2416 (N_2416,N_1329,N_1795);
or U2417 (N_2417,N_1722,N_1573);
nand U2418 (N_2418,N_1380,N_1643);
or U2419 (N_2419,N_1500,N_1715);
xnor U2420 (N_2420,N_1622,N_1274);
nand U2421 (N_2421,N_1711,N_1484);
xor U2422 (N_2422,N_1544,N_1691);
xnor U2423 (N_2423,N_1376,N_1496);
nand U2424 (N_2424,N_1777,N_1365);
or U2425 (N_2425,N_1769,N_1317);
nor U2426 (N_2426,N_1751,N_1435);
nor U2427 (N_2427,N_1774,N_1841);
or U2428 (N_2428,N_1384,N_1405);
nor U2429 (N_2429,N_1337,N_1287);
xnor U2430 (N_2430,N_1604,N_1743);
or U2431 (N_2431,N_1656,N_1549);
and U2432 (N_2432,N_1313,N_1784);
nor U2433 (N_2433,N_1282,N_1591);
nand U2434 (N_2434,N_1610,N_1341);
and U2435 (N_2435,N_1712,N_1414);
and U2436 (N_2436,N_1516,N_1472);
and U2437 (N_2437,N_1757,N_1665);
nor U2438 (N_2438,N_1721,N_1633);
nand U2439 (N_2439,N_1874,N_1382);
or U2440 (N_2440,N_1519,N_1324);
nand U2441 (N_2441,N_1684,N_1561);
xor U2442 (N_2442,N_1602,N_1469);
and U2443 (N_2443,N_1270,N_1278);
and U2444 (N_2444,N_1474,N_1677);
nand U2445 (N_2445,N_1309,N_1654);
nor U2446 (N_2446,N_1763,N_1631);
or U2447 (N_2447,N_1834,N_1726);
and U2448 (N_2448,N_1354,N_1483);
or U2449 (N_2449,N_1395,N_1715);
and U2450 (N_2450,N_1556,N_1395);
nand U2451 (N_2451,N_1836,N_1308);
nor U2452 (N_2452,N_1768,N_1654);
xnor U2453 (N_2453,N_1354,N_1567);
xnor U2454 (N_2454,N_1308,N_1762);
and U2455 (N_2455,N_1530,N_1475);
nor U2456 (N_2456,N_1604,N_1478);
nor U2457 (N_2457,N_1680,N_1717);
nor U2458 (N_2458,N_1383,N_1456);
xnor U2459 (N_2459,N_1714,N_1609);
or U2460 (N_2460,N_1854,N_1305);
xor U2461 (N_2461,N_1390,N_1545);
and U2462 (N_2462,N_1471,N_1689);
and U2463 (N_2463,N_1492,N_1289);
or U2464 (N_2464,N_1292,N_1566);
nand U2465 (N_2465,N_1607,N_1408);
and U2466 (N_2466,N_1397,N_1465);
nand U2467 (N_2467,N_1826,N_1674);
or U2468 (N_2468,N_1305,N_1530);
xnor U2469 (N_2469,N_1387,N_1265);
and U2470 (N_2470,N_1361,N_1782);
nor U2471 (N_2471,N_1590,N_1511);
xor U2472 (N_2472,N_1869,N_1658);
xnor U2473 (N_2473,N_1804,N_1754);
and U2474 (N_2474,N_1395,N_1508);
or U2475 (N_2475,N_1397,N_1416);
nor U2476 (N_2476,N_1721,N_1273);
or U2477 (N_2477,N_1732,N_1838);
or U2478 (N_2478,N_1517,N_1568);
or U2479 (N_2479,N_1273,N_1456);
xnor U2480 (N_2480,N_1581,N_1345);
nor U2481 (N_2481,N_1405,N_1847);
xnor U2482 (N_2482,N_1459,N_1493);
xnor U2483 (N_2483,N_1815,N_1433);
and U2484 (N_2484,N_1478,N_1417);
xnor U2485 (N_2485,N_1439,N_1743);
xnor U2486 (N_2486,N_1291,N_1563);
or U2487 (N_2487,N_1726,N_1800);
and U2488 (N_2488,N_1710,N_1315);
nand U2489 (N_2489,N_1459,N_1685);
nor U2490 (N_2490,N_1328,N_1275);
nor U2491 (N_2491,N_1811,N_1728);
nor U2492 (N_2492,N_1502,N_1374);
nand U2493 (N_2493,N_1292,N_1644);
or U2494 (N_2494,N_1561,N_1393);
nand U2495 (N_2495,N_1683,N_1281);
or U2496 (N_2496,N_1507,N_1327);
and U2497 (N_2497,N_1813,N_1386);
or U2498 (N_2498,N_1366,N_1464);
xor U2499 (N_2499,N_1432,N_1624);
nor U2500 (N_2500,N_1999,N_1930);
or U2501 (N_2501,N_2319,N_2036);
and U2502 (N_2502,N_2366,N_2171);
or U2503 (N_2503,N_2302,N_2151);
or U2504 (N_2504,N_2138,N_2196);
or U2505 (N_2505,N_1876,N_2423);
nand U2506 (N_2506,N_2383,N_2445);
nor U2507 (N_2507,N_2463,N_1907);
nand U2508 (N_2508,N_2386,N_2051);
and U2509 (N_2509,N_1929,N_2128);
nand U2510 (N_2510,N_2472,N_2117);
xor U2511 (N_2511,N_2040,N_2481);
nand U2512 (N_2512,N_2052,N_2275);
nor U2513 (N_2513,N_2178,N_2216);
or U2514 (N_2514,N_2371,N_1931);
or U2515 (N_2515,N_2426,N_2210);
nor U2516 (N_2516,N_2400,N_2301);
nor U2517 (N_2517,N_1901,N_2172);
and U2518 (N_2518,N_2049,N_2390);
xor U2519 (N_2519,N_2235,N_2233);
and U2520 (N_2520,N_2430,N_2041);
nand U2521 (N_2521,N_2376,N_2341);
or U2522 (N_2522,N_2057,N_2267);
xnor U2523 (N_2523,N_2250,N_1989);
nand U2524 (N_2524,N_2114,N_2339);
or U2525 (N_2525,N_2355,N_2300);
or U2526 (N_2526,N_2308,N_2285);
xnor U2527 (N_2527,N_2115,N_2175);
xnor U2528 (N_2528,N_2498,N_2450);
nor U2529 (N_2529,N_2225,N_1944);
nand U2530 (N_2530,N_2101,N_2050);
and U2531 (N_2531,N_2044,N_1909);
and U2532 (N_2532,N_2195,N_2042);
nand U2533 (N_2533,N_2217,N_2095);
and U2534 (N_2534,N_2224,N_2353);
and U2535 (N_2535,N_2268,N_1972);
nor U2536 (N_2536,N_2137,N_2311);
nand U2537 (N_2537,N_2009,N_2454);
nor U2538 (N_2538,N_2278,N_2062);
nand U2539 (N_2539,N_2082,N_2168);
xor U2540 (N_2540,N_2358,N_2088);
and U2541 (N_2541,N_2098,N_1880);
xor U2542 (N_2542,N_1978,N_2008);
nor U2543 (N_2543,N_2466,N_2262);
nand U2544 (N_2544,N_1890,N_2428);
or U2545 (N_2545,N_2438,N_1977);
nor U2546 (N_2546,N_2477,N_2211);
nand U2547 (N_2547,N_2401,N_1886);
xnor U2548 (N_2548,N_1953,N_2149);
and U2549 (N_2549,N_2134,N_2435);
xor U2550 (N_2550,N_2294,N_2414);
nor U2551 (N_2551,N_1904,N_2242);
nor U2552 (N_2552,N_2393,N_2464);
or U2553 (N_2553,N_2075,N_2251);
nand U2554 (N_2554,N_2465,N_2013);
nand U2555 (N_2555,N_2019,N_2150);
and U2556 (N_2556,N_2391,N_2360);
nand U2557 (N_2557,N_2127,N_1969);
or U2558 (N_2558,N_2432,N_2327);
nand U2559 (N_2559,N_1920,N_1885);
nand U2560 (N_2560,N_1985,N_2367);
xnor U2561 (N_2561,N_2192,N_2399);
nor U2562 (N_2562,N_2133,N_1893);
nor U2563 (N_2563,N_2298,N_1877);
nor U2564 (N_2564,N_2347,N_2475);
and U2565 (N_2565,N_1970,N_2204);
nand U2566 (N_2566,N_2462,N_2107);
nor U2567 (N_2567,N_2229,N_2072);
xor U2568 (N_2568,N_2370,N_1905);
nor U2569 (N_2569,N_2187,N_2316);
nor U2570 (N_2570,N_2304,N_2410);
xor U2571 (N_2571,N_2048,N_2324);
nand U2572 (N_2572,N_2344,N_2015);
and U2573 (N_2573,N_2154,N_2110);
or U2574 (N_2574,N_1964,N_2299);
nand U2575 (N_2575,N_2310,N_2482);
xnor U2576 (N_2576,N_1908,N_2499);
or U2577 (N_2577,N_2484,N_2193);
xnor U2578 (N_2578,N_1959,N_2120);
xnor U2579 (N_2579,N_2334,N_2007);
or U2580 (N_2580,N_2018,N_2495);
and U2581 (N_2581,N_2378,N_2024);
xor U2582 (N_2582,N_2361,N_2349);
or U2583 (N_2583,N_2159,N_2429);
or U2584 (N_2584,N_2081,N_1888);
nand U2585 (N_2585,N_2102,N_2086);
or U2586 (N_2586,N_2436,N_2116);
and U2587 (N_2587,N_2295,N_2248);
and U2588 (N_2588,N_2470,N_1912);
nand U2589 (N_2589,N_2173,N_2286);
nand U2590 (N_2590,N_2345,N_2274);
nor U2591 (N_2591,N_2080,N_1965);
and U2592 (N_2592,N_2119,N_2130);
nor U2593 (N_2593,N_1975,N_2025);
and U2594 (N_2594,N_2074,N_2092);
and U2595 (N_2595,N_2326,N_1891);
and U2596 (N_2596,N_2314,N_2212);
nand U2597 (N_2597,N_2201,N_2460);
xnor U2598 (N_2598,N_2241,N_2238);
and U2599 (N_2599,N_2028,N_2160);
nor U2600 (N_2600,N_2179,N_2090);
and U2601 (N_2601,N_2185,N_2017);
and U2602 (N_2602,N_2169,N_1988);
xnor U2603 (N_2603,N_2280,N_1884);
or U2604 (N_2604,N_2255,N_1949);
xor U2605 (N_2605,N_2317,N_2152);
or U2606 (N_2606,N_2143,N_2408);
nor U2607 (N_2607,N_2321,N_1941);
xnor U2608 (N_2608,N_2232,N_2068);
nor U2609 (N_2609,N_2109,N_2406);
xor U2610 (N_2610,N_1936,N_2003);
xor U2611 (N_2611,N_2365,N_2077);
xor U2612 (N_2612,N_2162,N_2253);
xor U2613 (N_2613,N_1987,N_2097);
xor U2614 (N_2614,N_2340,N_2087);
or U2615 (N_2615,N_1992,N_1932);
or U2616 (N_2616,N_2263,N_2440);
or U2617 (N_2617,N_1956,N_2407);
xor U2618 (N_2618,N_2281,N_2014);
and U2619 (N_2619,N_2444,N_2461);
xor U2620 (N_2620,N_2244,N_2228);
xnor U2621 (N_2621,N_2483,N_2157);
nor U2622 (N_2622,N_2431,N_2213);
or U2623 (N_2623,N_2166,N_1923);
xnor U2624 (N_2624,N_2234,N_2348);
or U2625 (N_2625,N_1973,N_2288);
nor U2626 (N_2626,N_1982,N_1960);
and U2627 (N_2627,N_1979,N_2227);
xor U2628 (N_2628,N_1957,N_1948);
or U2629 (N_2629,N_2079,N_2387);
and U2630 (N_2630,N_2479,N_2485);
xnor U2631 (N_2631,N_1955,N_2441);
and U2632 (N_2632,N_2389,N_2337);
and U2633 (N_2633,N_2118,N_1947);
and U2634 (N_2634,N_2146,N_2384);
xor U2635 (N_2635,N_2059,N_1950);
and U2636 (N_2636,N_2382,N_2420);
xnor U2637 (N_2637,N_1937,N_2437);
and U2638 (N_2638,N_2289,N_2106);
or U2639 (N_2639,N_1916,N_1952);
nor U2640 (N_2640,N_2427,N_2357);
or U2641 (N_2641,N_1983,N_2270);
and U2642 (N_2642,N_2397,N_2247);
and U2643 (N_2643,N_2329,N_2273);
or U2644 (N_2644,N_2473,N_2089);
xor U2645 (N_2645,N_1951,N_2027);
and U2646 (N_2646,N_2336,N_2125);
xor U2647 (N_2647,N_2103,N_2207);
nand U2648 (N_2648,N_2452,N_2409);
xnor U2649 (N_2649,N_2418,N_2331);
and U2650 (N_2650,N_1993,N_2372);
or U2651 (N_2651,N_1926,N_2226);
or U2652 (N_2652,N_1990,N_2279);
nor U2653 (N_2653,N_2395,N_2377);
or U2654 (N_2654,N_2184,N_2352);
xor U2655 (N_2655,N_2307,N_1906);
nor U2656 (N_2656,N_1879,N_2064);
and U2657 (N_2657,N_2342,N_2455);
and U2658 (N_2658,N_2148,N_2290);
or U2659 (N_2659,N_2139,N_2188);
xnor U2660 (N_2660,N_2328,N_2209);
xnor U2661 (N_2661,N_2412,N_2039);
or U2662 (N_2662,N_1971,N_2140);
nor U2663 (N_2663,N_1986,N_2487);
xor U2664 (N_2664,N_2197,N_1974);
nand U2665 (N_2665,N_2396,N_1934);
and U2666 (N_2666,N_1910,N_2385);
nand U2667 (N_2667,N_2005,N_2419);
nor U2668 (N_2668,N_2156,N_2182);
nor U2669 (N_2669,N_1958,N_1961);
or U2670 (N_2670,N_2416,N_2434);
and U2671 (N_2671,N_2394,N_2056);
and U2672 (N_2672,N_2373,N_2076);
nand U2673 (N_2673,N_2121,N_2252);
and U2674 (N_2674,N_2046,N_1967);
nand U2675 (N_2675,N_2266,N_1946);
or U2676 (N_2676,N_2451,N_2313);
xor U2677 (N_2677,N_2002,N_2231);
nor U2678 (N_2678,N_1902,N_1976);
or U2679 (N_2679,N_1917,N_2392);
or U2680 (N_2680,N_2021,N_2291);
nand U2681 (N_2681,N_2239,N_2272);
xnor U2682 (N_2682,N_2065,N_2260);
nor U2683 (N_2683,N_2142,N_2332);
nor U2684 (N_2684,N_2144,N_2369);
nor U2685 (N_2685,N_2218,N_2066);
or U2686 (N_2686,N_2493,N_2404);
and U2687 (N_2687,N_2402,N_2323);
and U2688 (N_2688,N_2011,N_2257);
xnor U2689 (N_2689,N_2053,N_1991);
xnor U2690 (N_2690,N_1984,N_2132);
nor U2691 (N_2691,N_2006,N_2265);
or U2692 (N_2692,N_1878,N_1922);
xnor U2693 (N_2693,N_1962,N_1994);
nand U2694 (N_2694,N_1966,N_2354);
nand U2695 (N_2695,N_2422,N_2359);
and U2696 (N_2696,N_2029,N_2067);
or U2697 (N_2697,N_2292,N_1881);
nand U2698 (N_2698,N_1924,N_2403);
nor U2699 (N_2699,N_2026,N_2236);
and U2700 (N_2700,N_2163,N_2073);
or U2701 (N_2701,N_2282,N_2381);
xor U2702 (N_2702,N_2186,N_2442);
nor U2703 (N_2703,N_2047,N_2237);
and U2704 (N_2704,N_2456,N_2276);
nand U2705 (N_2705,N_1938,N_2190);
nand U2706 (N_2706,N_2259,N_1892);
nand U2707 (N_2707,N_1913,N_2258);
nor U2708 (N_2708,N_2122,N_1896);
nand U2709 (N_2709,N_1940,N_2467);
or U2710 (N_2710,N_2045,N_2012);
nand U2711 (N_2711,N_2283,N_2063);
nor U2712 (N_2712,N_1997,N_2459);
xor U2713 (N_2713,N_2091,N_2447);
or U2714 (N_2714,N_1980,N_2468);
or U2715 (N_2715,N_2368,N_2058);
and U2716 (N_2716,N_2164,N_2170);
nor U2717 (N_2717,N_1927,N_2060);
and U2718 (N_2718,N_1882,N_2034);
nand U2719 (N_2719,N_2246,N_2411);
and U2720 (N_2720,N_2489,N_2112);
nor U2721 (N_2721,N_2322,N_2476);
or U2722 (N_2722,N_2004,N_1943);
nand U2723 (N_2723,N_2126,N_2105);
and U2724 (N_2724,N_2099,N_2240);
or U2725 (N_2725,N_2458,N_2351);
and U2726 (N_2726,N_2271,N_1998);
nand U2727 (N_2727,N_2448,N_2296);
nor U2728 (N_2728,N_2131,N_2415);
or U2729 (N_2729,N_2312,N_2123);
xor U2730 (N_2730,N_2153,N_2083);
or U2731 (N_2731,N_2261,N_2165);
or U2732 (N_2732,N_2453,N_2205);
nand U2733 (N_2733,N_2030,N_2035);
nand U2734 (N_2734,N_2471,N_1996);
nand U2735 (N_2735,N_2199,N_2449);
nand U2736 (N_2736,N_1942,N_2486);
or U2737 (N_2737,N_2001,N_2023);
or U2738 (N_2738,N_2335,N_2364);
xnor U2739 (N_2739,N_2135,N_2497);
or U2740 (N_2740,N_2136,N_2303);
nand U2741 (N_2741,N_2043,N_2494);
nor U2742 (N_2742,N_2287,N_2439);
or U2743 (N_2743,N_2256,N_2297);
xor U2744 (N_2744,N_2085,N_1919);
and U2745 (N_2745,N_2309,N_2177);
nand U2746 (N_2746,N_2433,N_2306);
nor U2747 (N_2747,N_2264,N_2147);
and U2748 (N_2748,N_2398,N_2037);
xor U2749 (N_2749,N_2033,N_2254);
nor U2750 (N_2750,N_2061,N_2069);
nand U2751 (N_2751,N_2469,N_2492);
xnor U2752 (N_2752,N_2093,N_2388);
or U2753 (N_2753,N_1915,N_2183);
xnor U2754 (N_2754,N_2100,N_2284);
nand U2755 (N_2755,N_2198,N_2315);
or U2756 (N_2756,N_2474,N_2054);
nor U2757 (N_2757,N_2016,N_1875);
xnor U2758 (N_2758,N_2363,N_2496);
nand U2759 (N_2759,N_2078,N_1898);
nor U2760 (N_2760,N_2031,N_2070);
xnor U2761 (N_2761,N_2343,N_2022);
and U2762 (N_2762,N_2222,N_2333);
nand U2763 (N_2763,N_2374,N_2141);
or U2764 (N_2764,N_1911,N_2379);
and U2765 (N_2765,N_2491,N_2446);
nor U2766 (N_2766,N_1900,N_2490);
and U2767 (N_2767,N_1968,N_2320);
nand U2768 (N_2768,N_2330,N_1933);
and U2769 (N_2769,N_2375,N_2181);
nor U2770 (N_2770,N_2155,N_2424);
xnor U2771 (N_2771,N_2071,N_2425);
or U2772 (N_2772,N_2269,N_2305);
or U2773 (N_2773,N_1945,N_2338);
and U2774 (N_2774,N_1899,N_1995);
xnor U2775 (N_2775,N_2220,N_2219);
and U2776 (N_2776,N_2208,N_1895);
xnor U2777 (N_2777,N_1887,N_2215);
and U2778 (N_2778,N_2245,N_2405);
nor U2779 (N_2779,N_2161,N_2200);
nand U2780 (N_2780,N_2223,N_2380);
nand U2781 (N_2781,N_1883,N_1954);
nand U2782 (N_2782,N_2111,N_2096);
and U2783 (N_2783,N_2202,N_2167);
xor U2784 (N_2784,N_1939,N_1918);
or U2785 (N_2785,N_2206,N_2000);
nor U2786 (N_2786,N_2176,N_2488);
and U2787 (N_2787,N_2191,N_1925);
nor U2788 (N_2788,N_2350,N_2180);
or U2789 (N_2789,N_2318,N_2194);
or U2790 (N_2790,N_1935,N_2032);
xor U2791 (N_2791,N_2108,N_2038);
xnor U2792 (N_2792,N_2480,N_1928);
and U2793 (N_2793,N_2084,N_2249);
xnor U2794 (N_2794,N_2413,N_1921);
xnor U2795 (N_2795,N_1894,N_2129);
or U2796 (N_2796,N_2145,N_2293);
or U2797 (N_2797,N_2158,N_1914);
and U2798 (N_2798,N_1903,N_2221);
or U2799 (N_2799,N_2362,N_2113);
xor U2800 (N_2800,N_2421,N_2243);
and U2801 (N_2801,N_2325,N_1981);
or U2802 (N_2802,N_1889,N_2457);
and U2803 (N_2803,N_1897,N_1963);
nand U2804 (N_2804,N_2010,N_2094);
nand U2805 (N_2805,N_2124,N_2203);
nand U2806 (N_2806,N_2230,N_2055);
and U2807 (N_2807,N_2356,N_2478);
or U2808 (N_2808,N_2104,N_2417);
xor U2809 (N_2809,N_2189,N_2214);
or U2810 (N_2810,N_2020,N_2443);
nand U2811 (N_2811,N_2277,N_2346);
nand U2812 (N_2812,N_2174,N_2142);
xnor U2813 (N_2813,N_2357,N_2246);
nand U2814 (N_2814,N_1974,N_2416);
nand U2815 (N_2815,N_2385,N_2413);
nor U2816 (N_2816,N_2388,N_2318);
or U2817 (N_2817,N_2094,N_2005);
nand U2818 (N_2818,N_1895,N_2085);
nand U2819 (N_2819,N_2034,N_1900);
nand U2820 (N_2820,N_2272,N_1959);
xor U2821 (N_2821,N_2201,N_1987);
or U2822 (N_2822,N_2484,N_2065);
or U2823 (N_2823,N_2086,N_1986);
and U2824 (N_2824,N_1930,N_1972);
nor U2825 (N_2825,N_2069,N_2019);
nand U2826 (N_2826,N_2309,N_2297);
nand U2827 (N_2827,N_2435,N_2208);
nand U2828 (N_2828,N_2087,N_2465);
or U2829 (N_2829,N_2463,N_2012);
nor U2830 (N_2830,N_2432,N_2137);
nor U2831 (N_2831,N_2210,N_2253);
xor U2832 (N_2832,N_2361,N_2455);
nor U2833 (N_2833,N_2323,N_2046);
xnor U2834 (N_2834,N_2386,N_1996);
nor U2835 (N_2835,N_2018,N_2005);
nor U2836 (N_2836,N_2405,N_2099);
xor U2837 (N_2837,N_1915,N_2041);
nor U2838 (N_2838,N_1977,N_1934);
nor U2839 (N_2839,N_1917,N_1938);
and U2840 (N_2840,N_2293,N_1876);
or U2841 (N_2841,N_2096,N_2240);
xor U2842 (N_2842,N_2097,N_1955);
or U2843 (N_2843,N_1957,N_2160);
nor U2844 (N_2844,N_2182,N_2152);
nand U2845 (N_2845,N_2153,N_2252);
or U2846 (N_2846,N_2052,N_2261);
xor U2847 (N_2847,N_2195,N_2103);
or U2848 (N_2848,N_2450,N_2197);
or U2849 (N_2849,N_1987,N_2170);
nand U2850 (N_2850,N_2347,N_2064);
nor U2851 (N_2851,N_2470,N_2038);
xnor U2852 (N_2852,N_2434,N_2170);
xnor U2853 (N_2853,N_1966,N_1953);
nand U2854 (N_2854,N_1992,N_2380);
xnor U2855 (N_2855,N_1963,N_1948);
or U2856 (N_2856,N_2303,N_2341);
or U2857 (N_2857,N_2206,N_2373);
nand U2858 (N_2858,N_2132,N_2110);
nor U2859 (N_2859,N_1994,N_2108);
nand U2860 (N_2860,N_2142,N_1949);
and U2861 (N_2861,N_2099,N_2043);
or U2862 (N_2862,N_2176,N_2162);
or U2863 (N_2863,N_2228,N_2494);
xor U2864 (N_2864,N_1997,N_2261);
xor U2865 (N_2865,N_1923,N_2418);
nor U2866 (N_2866,N_1957,N_2263);
nand U2867 (N_2867,N_2330,N_2257);
nor U2868 (N_2868,N_2004,N_2146);
nor U2869 (N_2869,N_2176,N_2197);
nor U2870 (N_2870,N_1883,N_2429);
nor U2871 (N_2871,N_1969,N_2449);
nand U2872 (N_2872,N_2050,N_2296);
nand U2873 (N_2873,N_1927,N_2288);
or U2874 (N_2874,N_2059,N_2442);
or U2875 (N_2875,N_2260,N_2099);
nor U2876 (N_2876,N_2022,N_2261);
xnor U2877 (N_2877,N_2176,N_2484);
xor U2878 (N_2878,N_2421,N_2064);
xnor U2879 (N_2879,N_2045,N_1900);
xnor U2880 (N_2880,N_1943,N_2182);
nand U2881 (N_2881,N_2215,N_2302);
or U2882 (N_2882,N_2109,N_1915);
nor U2883 (N_2883,N_1916,N_2154);
or U2884 (N_2884,N_2225,N_2474);
nand U2885 (N_2885,N_2092,N_2486);
nand U2886 (N_2886,N_1996,N_2109);
xor U2887 (N_2887,N_2446,N_2119);
nand U2888 (N_2888,N_1960,N_2372);
nand U2889 (N_2889,N_2453,N_2301);
or U2890 (N_2890,N_2462,N_2082);
xor U2891 (N_2891,N_2184,N_2249);
nor U2892 (N_2892,N_2127,N_2083);
and U2893 (N_2893,N_2148,N_1895);
or U2894 (N_2894,N_2157,N_2097);
or U2895 (N_2895,N_2302,N_1927);
nand U2896 (N_2896,N_2491,N_2495);
nand U2897 (N_2897,N_1993,N_2315);
or U2898 (N_2898,N_1910,N_2205);
or U2899 (N_2899,N_2129,N_1912);
nor U2900 (N_2900,N_2459,N_2343);
and U2901 (N_2901,N_2373,N_2469);
or U2902 (N_2902,N_2224,N_2492);
and U2903 (N_2903,N_2373,N_2248);
nand U2904 (N_2904,N_2414,N_1996);
or U2905 (N_2905,N_1904,N_1888);
nand U2906 (N_2906,N_1999,N_2110);
nand U2907 (N_2907,N_2099,N_2160);
and U2908 (N_2908,N_1961,N_2245);
or U2909 (N_2909,N_2175,N_2179);
and U2910 (N_2910,N_2426,N_2340);
nor U2911 (N_2911,N_2441,N_2315);
xnor U2912 (N_2912,N_2299,N_2382);
or U2913 (N_2913,N_2100,N_2371);
or U2914 (N_2914,N_2220,N_2189);
nand U2915 (N_2915,N_2290,N_2046);
nor U2916 (N_2916,N_2348,N_2198);
nor U2917 (N_2917,N_2036,N_2092);
and U2918 (N_2918,N_2379,N_2348);
xor U2919 (N_2919,N_1926,N_2359);
or U2920 (N_2920,N_1977,N_2482);
nand U2921 (N_2921,N_2341,N_2368);
nor U2922 (N_2922,N_2142,N_2073);
or U2923 (N_2923,N_2333,N_2476);
nor U2924 (N_2924,N_2309,N_2399);
and U2925 (N_2925,N_2028,N_2470);
or U2926 (N_2926,N_1919,N_2121);
nand U2927 (N_2927,N_1955,N_2315);
nor U2928 (N_2928,N_2322,N_2368);
nor U2929 (N_2929,N_2261,N_1951);
and U2930 (N_2930,N_2212,N_2147);
or U2931 (N_2931,N_2274,N_1978);
xnor U2932 (N_2932,N_2470,N_2229);
nand U2933 (N_2933,N_1917,N_2314);
or U2934 (N_2934,N_2223,N_2209);
xnor U2935 (N_2935,N_2410,N_2088);
nand U2936 (N_2936,N_2066,N_2261);
nor U2937 (N_2937,N_1965,N_2172);
or U2938 (N_2938,N_2209,N_2334);
and U2939 (N_2939,N_2180,N_2064);
xnor U2940 (N_2940,N_2105,N_2379);
xor U2941 (N_2941,N_2101,N_1946);
nor U2942 (N_2942,N_2062,N_2374);
or U2943 (N_2943,N_2496,N_2331);
xor U2944 (N_2944,N_2064,N_1932);
xor U2945 (N_2945,N_2457,N_2261);
nand U2946 (N_2946,N_2091,N_1964);
and U2947 (N_2947,N_1988,N_1948);
and U2948 (N_2948,N_2067,N_2451);
nor U2949 (N_2949,N_1982,N_1919);
or U2950 (N_2950,N_2305,N_2349);
nand U2951 (N_2951,N_2139,N_2346);
and U2952 (N_2952,N_2334,N_2078);
xnor U2953 (N_2953,N_1917,N_2422);
xor U2954 (N_2954,N_2023,N_2051);
and U2955 (N_2955,N_2018,N_1953);
and U2956 (N_2956,N_2315,N_2126);
nor U2957 (N_2957,N_2100,N_2396);
nand U2958 (N_2958,N_2198,N_2069);
nand U2959 (N_2959,N_2299,N_2267);
or U2960 (N_2960,N_1941,N_2436);
nor U2961 (N_2961,N_2270,N_1969);
xnor U2962 (N_2962,N_1931,N_2327);
or U2963 (N_2963,N_2126,N_2229);
nand U2964 (N_2964,N_1946,N_2405);
xnor U2965 (N_2965,N_2326,N_2460);
or U2966 (N_2966,N_2442,N_2079);
xnor U2967 (N_2967,N_2018,N_1930);
or U2968 (N_2968,N_2253,N_2206);
nor U2969 (N_2969,N_2034,N_1916);
xor U2970 (N_2970,N_2324,N_2241);
or U2971 (N_2971,N_2480,N_2151);
xnor U2972 (N_2972,N_2336,N_2354);
and U2973 (N_2973,N_2465,N_2464);
nand U2974 (N_2974,N_1905,N_2162);
nand U2975 (N_2975,N_1937,N_2495);
and U2976 (N_2976,N_1933,N_1998);
xor U2977 (N_2977,N_1930,N_2463);
and U2978 (N_2978,N_2349,N_2078);
and U2979 (N_2979,N_2158,N_2304);
xor U2980 (N_2980,N_2026,N_1968);
nor U2981 (N_2981,N_2048,N_2425);
xor U2982 (N_2982,N_2408,N_1922);
xnor U2983 (N_2983,N_2199,N_2454);
or U2984 (N_2984,N_1947,N_2279);
xnor U2985 (N_2985,N_2198,N_2378);
xor U2986 (N_2986,N_2419,N_2202);
nand U2987 (N_2987,N_2165,N_2463);
or U2988 (N_2988,N_2013,N_1902);
or U2989 (N_2989,N_2497,N_2066);
or U2990 (N_2990,N_1912,N_2050);
nand U2991 (N_2991,N_2454,N_2048);
xor U2992 (N_2992,N_1949,N_2477);
xnor U2993 (N_2993,N_2370,N_1940);
nor U2994 (N_2994,N_1971,N_2460);
or U2995 (N_2995,N_1977,N_1933);
nor U2996 (N_2996,N_2170,N_2475);
xor U2997 (N_2997,N_2125,N_2218);
or U2998 (N_2998,N_2073,N_2070);
xnor U2999 (N_2999,N_2031,N_1983);
and U3000 (N_3000,N_2472,N_2151);
nand U3001 (N_3001,N_2084,N_2492);
xor U3002 (N_3002,N_1875,N_2416);
nor U3003 (N_3003,N_1935,N_2303);
or U3004 (N_3004,N_2046,N_1889);
and U3005 (N_3005,N_1949,N_2330);
nand U3006 (N_3006,N_2271,N_2252);
nor U3007 (N_3007,N_1939,N_2040);
nor U3008 (N_3008,N_2375,N_2091);
or U3009 (N_3009,N_2403,N_1912);
xor U3010 (N_3010,N_2174,N_2273);
or U3011 (N_3011,N_1995,N_2140);
xnor U3012 (N_3012,N_2140,N_2472);
xnor U3013 (N_3013,N_2456,N_2203);
or U3014 (N_3014,N_2477,N_1981);
nand U3015 (N_3015,N_2338,N_1986);
and U3016 (N_3016,N_2284,N_2418);
and U3017 (N_3017,N_2383,N_2389);
xor U3018 (N_3018,N_1883,N_2330);
xnor U3019 (N_3019,N_2446,N_1938);
nor U3020 (N_3020,N_2191,N_1882);
xnor U3021 (N_3021,N_2425,N_1913);
nor U3022 (N_3022,N_2252,N_2409);
nor U3023 (N_3023,N_2129,N_2116);
or U3024 (N_3024,N_2026,N_2404);
xnor U3025 (N_3025,N_2305,N_2047);
nor U3026 (N_3026,N_2393,N_2123);
or U3027 (N_3027,N_2093,N_2006);
and U3028 (N_3028,N_2421,N_2454);
xor U3029 (N_3029,N_2288,N_2056);
and U3030 (N_3030,N_2433,N_2031);
and U3031 (N_3031,N_2437,N_2338);
xor U3032 (N_3032,N_2376,N_2299);
nor U3033 (N_3033,N_2497,N_1993);
nor U3034 (N_3034,N_2314,N_2302);
or U3035 (N_3035,N_2165,N_2109);
or U3036 (N_3036,N_2199,N_2065);
nor U3037 (N_3037,N_1985,N_2423);
xor U3038 (N_3038,N_2029,N_2426);
nand U3039 (N_3039,N_2047,N_2430);
and U3040 (N_3040,N_2460,N_2398);
nor U3041 (N_3041,N_2139,N_2286);
and U3042 (N_3042,N_2244,N_2460);
and U3043 (N_3043,N_2074,N_2485);
nand U3044 (N_3044,N_2149,N_2487);
xor U3045 (N_3045,N_2349,N_2056);
nand U3046 (N_3046,N_2483,N_2071);
or U3047 (N_3047,N_2263,N_2182);
and U3048 (N_3048,N_1975,N_2329);
nor U3049 (N_3049,N_2068,N_2110);
and U3050 (N_3050,N_2248,N_2397);
xor U3051 (N_3051,N_2440,N_2136);
nand U3052 (N_3052,N_2026,N_2040);
nor U3053 (N_3053,N_2483,N_2326);
xnor U3054 (N_3054,N_2454,N_2114);
nand U3055 (N_3055,N_2258,N_2102);
and U3056 (N_3056,N_2269,N_2462);
nor U3057 (N_3057,N_2180,N_2173);
nor U3058 (N_3058,N_2295,N_2171);
xnor U3059 (N_3059,N_1987,N_2195);
nand U3060 (N_3060,N_2383,N_2300);
nand U3061 (N_3061,N_2453,N_2350);
nor U3062 (N_3062,N_2172,N_2389);
nand U3063 (N_3063,N_2012,N_2493);
nor U3064 (N_3064,N_2163,N_2045);
xor U3065 (N_3065,N_2059,N_2258);
or U3066 (N_3066,N_1877,N_2113);
and U3067 (N_3067,N_2033,N_2200);
nand U3068 (N_3068,N_2355,N_1955);
or U3069 (N_3069,N_2085,N_2340);
or U3070 (N_3070,N_2191,N_2021);
and U3071 (N_3071,N_2000,N_2388);
nor U3072 (N_3072,N_2262,N_1892);
and U3073 (N_3073,N_2229,N_1879);
nand U3074 (N_3074,N_2433,N_1972);
nand U3075 (N_3075,N_2050,N_2214);
xnor U3076 (N_3076,N_2069,N_1911);
and U3077 (N_3077,N_2020,N_2149);
xnor U3078 (N_3078,N_2140,N_2414);
and U3079 (N_3079,N_2458,N_2318);
nand U3080 (N_3080,N_2103,N_2153);
nor U3081 (N_3081,N_2379,N_2321);
xor U3082 (N_3082,N_1995,N_2105);
or U3083 (N_3083,N_2407,N_2399);
or U3084 (N_3084,N_2398,N_2410);
xor U3085 (N_3085,N_2171,N_2488);
xnor U3086 (N_3086,N_2436,N_2289);
nor U3087 (N_3087,N_2389,N_2283);
nor U3088 (N_3088,N_2385,N_2335);
nor U3089 (N_3089,N_2173,N_2456);
nor U3090 (N_3090,N_2187,N_2064);
and U3091 (N_3091,N_2477,N_2204);
and U3092 (N_3092,N_2204,N_2116);
or U3093 (N_3093,N_2266,N_2015);
nand U3094 (N_3094,N_2069,N_2264);
and U3095 (N_3095,N_2065,N_2284);
nand U3096 (N_3096,N_2472,N_2323);
xnor U3097 (N_3097,N_2087,N_2385);
nor U3098 (N_3098,N_2102,N_2414);
xor U3099 (N_3099,N_2176,N_1897);
nand U3100 (N_3100,N_2271,N_2015);
or U3101 (N_3101,N_2365,N_2395);
xnor U3102 (N_3102,N_2197,N_1963);
or U3103 (N_3103,N_1878,N_2499);
nand U3104 (N_3104,N_2338,N_2025);
or U3105 (N_3105,N_1905,N_2014);
nand U3106 (N_3106,N_1899,N_1955);
and U3107 (N_3107,N_2109,N_2198);
nor U3108 (N_3108,N_2003,N_2389);
nor U3109 (N_3109,N_2284,N_2244);
xor U3110 (N_3110,N_1880,N_2259);
or U3111 (N_3111,N_2282,N_2193);
and U3112 (N_3112,N_1960,N_2064);
xor U3113 (N_3113,N_2412,N_2074);
nor U3114 (N_3114,N_2096,N_1917);
or U3115 (N_3115,N_2059,N_2229);
xor U3116 (N_3116,N_2126,N_2415);
xnor U3117 (N_3117,N_2094,N_2244);
nand U3118 (N_3118,N_2269,N_2140);
xnor U3119 (N_3119,N_2162,N_2032);
or U3120 (N_3120,N_1933,N_2491);
nand U3121 (N_3121,N_2220,N_2150);
nand U3122 (N_3122,N_2172,N_1970);
nor U3123 (N_3123,N_2066,N_2442);
xor U3124 (N_3124,N_2330,N_2469);
nor U3125 (N_3125,N_3016,N_2662);
nor U3126 (N_3126,N_2565,N_2622);
and U3127 (N_3127,N_3116,N_2883);
xor U3128 (N_3128,N_3035,N_2770);
or U3129 (N_3129,N_2516,N_2660);
nor U3130 (N_3130,N_2913,N_2994);
nor U3131 (N_3131,N_2553,N_2764);
and U3132 (N_3132,N_2875,N_3013);
and U3133 (N_3133,N_2851,N_2942);
xor U3134 (N_3134,N_2608,N_2776);
or U3135 (N_3135,N_2984,N_3081);
and U3136 (N_3136,N_2576,N_2784);
or U3137 (N_3137,N_2733,N_2872);
or U3138 (N_3138,N_2932,N_2647);
and U3139 (N_3139,N_2893,N_2876);
and U3140 (N_3140,N_2822,N_2807);
or U3141 (N_3141,N_3056,N_3122);
nor U3142 (N_3142,N_2869,N_2732);
nor U3143 (N_3143,N_2987,N_3042);
or U3144 (N_3144,N_2537,N_2930);
or U3145 (N_3145,N_3043,N_2960);
and U3146 (N_3146,N_3039,N_2914);
nand U3147 (N_3147,N_3015,N_2670);
and U3148 (N_3148,N_3024,N_2898);
xnor U3149 (N_3149,N_2561,N_2642);
nor U3150 (N_3150,N_2825,N_3031);
xor U3151 (N_3151,N_2800,N_2551);
nor U3152 (N_3152,N_2916,N_2743);
and U3153 (N_3153,N_2862,N_3046);
xor U3154 (N_3154,N_3113,N_2767);
or U3155 (N_3155,N_2538,N_2755);
or U3156 (N_3156,N_2992,N_3096);
nor U3157 (N_3157,N_2939,N_2635);
xor U3158 (N_3158,N_2886,N_2737);
and U3159 (N_3159,N_3073,N_2688);
or U3160 (N_3160,N_2997,N_2915);
xnor U3161 (N_3161,N_2759,N_3062);
nor U3162 (N_3162,N_2588,N_3004);
or U3163 (N_3163,N_2777,N_2967);
nand U3164 (N_3164,N_3050,N_2760);
xnor U3165 (N_3165,N_2510,N_2547);
nand U3166 (N_3166,N_2958,N_2607);
nand U3167 (N_3167,N_2781,N_3103);
nand U3168 (N_3168,N_2559,N_2936);
xnor U3169 (N_3169,N_2909,N_2650);
xor U3170 (N_3170,N_3040,N_2697);
xnor U3171 (N_3171,N_2836,N_2792);
or U3172 (N_3172,N_2736,N_2723);
xnor U3173 (N_3173,N_2679,N_2587);
nor U3174 (N_3174,N_3099,N_2560);
and U3175 (N_3175,N_3089,N_2704);
and U3176 (N_3176,N_3036,N_3071);
nand U3177 (N_3177,N_3064,N_2933);
nand U3178 (N_3178,N_2797,N_2630);
or U3179 (N_3179,N_2756,N_2597);
or U3180 (N_3180,N_2899,N_2721);
and U3181 (N_3181,N_2625,N_2941);
nor U3182 (N_3182,N_2712,N_3101);
nor U3183 (N_3183,N_2602,N_2885);
nor U3184 (N_3184,N_2680,N_2705);
or U3185 (N_3185,N_3027,N_3001);
or U3186 (N_3186,N_2605,N_3077);
nand U3187 (N_3187,N_2891,N_2586);
and U3188 (N_3188,N_2549,N_3105);
or U3189 (N_3189,N_2956,N_2754);
or U3190 (N_3190,N_2703,N_2813);
nand U3191 (N_3191,N_2888,N_3048);
nand U3192 (N_3192,N_2791,N_3028);
and U3193 (N_3193,N_2534,N_2848);
or U3194 (N_3194,N_2830,N_3005);
and U3195 (N_3195,N_2502,N_2711);
nor U3196 (N_3196,N_2707,N_2852);
nor U3197 (N_3197,N_2540,N_3025);
or U3198 (N_3198,N_2867,N_3102);
nand U3199 (N_3199,N_2975,N_2773);
xor U3200 (N_3200,N_2603,N_2990);
and U3201 (N_3201,N_2908,N_2833);
or U3202 (N_3202,N_2782,N_2877);
nand U3203 (N_3203,N_2779,N_2722);
nor U3204 (N_3204,N_2817,N_2550);
nor U3205 (N_3205,N_2708,N_3061);
and U3206 (N_3206,N_2738,N_3037);
and U3207 (N_3207,N_2887,N_2674);
and U3208 (N_3208,N_2988,N_2512);
xnor U3209 (N_3209,N_2793,N_3010);
nor U3210 (N_3210,N_2959,N_2881);
nor U3211 (N_3211,N_2815,N_2904);
nor U3212 (N_3212,N_3114,N_3087);
and U3213 (N_3213,N_2644,N_2826);
nor U3214 (N_3214,N_2824,N_2879);
nand U3215 (N_3215,N_2573,N_2971);
nor U3216 (N_3216,N_3038,N_2526);
nor U3217 (N_3217,N_2974,N_2818);
xnor U3218 (N_3218,N_2774,N_2805);
xor U3219 (N_3219,N_2977,N_2799);
nor U3220 (N_3220,N_2530,N_2541);
or U3221 (N_3221,N_2900,N_2798);
or U3222 (N_3222,N_2716,N_2574);
nor U3223 (N_3223,N_2517,N_3119);
or U3224 (N_3224,N_2922,N_2804);
xor U3225 (N_3225,N_3044,N_2570);
nand U3226 (N_3226,N_2567,N_3084);
nand U3227 (N_3227,N_2558,N_2533);
and U3228 (N_3228,N_2522,N_2785);
and U3229 (N_3229,N_2726,N_2884);
or U3230 (N_3230,N_2715,N_3095);
nand U3231 (N_3231,N_2969,N_3076);
nor U3232 (N_3232,N_2860,N_2931);
and U3233 (N_3233,N_2861,N_2944);
and U3234 (N_3234,N_2903,N_2693);
xnor U3235 (N_3235,N_2532,N_2649);
nand U3236 (N_3236,N_2866,N_2746);
nand U3237 (N_3237,N_2664,N_2921);
nand U3238 (N_3238,N_2518,N_2882);
and U3239 (N_3239,N_2810,N_2957);
nand U3240 (N_3240,N_2762,N_3063);
xnor U3241 (N_3241,N_2575,N_3093);
nand U3242 (N_3242,N_2802,N_2927);
nand U3243 (N_3243,N_2741,N_2878);
or U3244 (N_3244,N_2686,N_2968);
nor U3245 (N_3245,N_2896,N_2717);
or U3246 (N_3246,N_2528,N_2970);
xor U3247 (N_3247,N_2695,N_2819);
nor U3248 (N_3248,N_3022,N_3051);
nand U3249 (N_3249,N_2778,N_2965);
or U3250 (N_3250,N_2521,N_3019);
nor U3251 (N_3251,N_2613,N_3108);
nand U3252 (N_3252,N_3023,N_2581);
xnor U3253 (N_3253,N_2681,N_2769);
nand U3254 (N_3254,N_3026,N_2657);
nand U3255 (N_3255,N_2911,N_2897);
nor U3256 (N_3256,N_2656,N_2728);
nand U3257 (N_3257,N_2617,N_2783);
xnor U3258 (N_3258,N_3069,N_3110);
or U3259 (N_3259,N_2973,N_3032);
nand U3260 (N_3260,N_2545,N_2689);
nor U3261 (N_3261,N_2951,N_2513);
and U3262 (N_3262,N_2803,N_2548);
and U3263 (N_3263,N_3017,N_2604);
and U3264 (N_3264,N_2980,N_2870);
xnor U3265 (N_3265,N_2788,N_2752);
nor U3266 (N_3266,N_2906,N_2683);
or U3267 (N_3267,N_3065,N_2691);
or U3268 (N_3268,N_2854,N_3052);
nor U3269 (N_3269,N_2655,N_2591);
nor U3270 (N_3270,N_2566,N_2672);
or U3271 (N_3271,N_3124,N_3118);
nand U3272 (N_3272,N_2511,N_2859);
and U3273 (N_3273,N_2606,N_2639);
nand U3274 (N_3274,N_2850,N_2814);
xor U3275 (N_3275,N_2827,N_2938);
nand U3276 (N_3276,N_2734,N_2535);
and U3277 (N_3277,N_2641,N_3053);
nand U3278 (N_3278,N_3080,N_2757);
xnor U3279 (N_3279,N_2843,N_2562);
nand U3280 (N_3280,N_3111,N_2621);
nor U3281 (N_3281,N_2963,N_2620);
xor U3282 (N_3282,N_2787,N_3029);
nand U3283 (N_3283,N_2976,N_2811);
nor U3284 (N_3284,N_2555,N_2895);
nand U3285 (N_3285,N_2694,N_2614);
and U3286 (N_3286,N_3088,N_3068);
and U3287 (N_3287,N_2648,N_2790);
or U3288 (N_3288,N_3109,N_2678);
or U3289 (N_3289,N_2636,N_2593);
or U3290 (N_3290,N_2753,N_2982);
nand U3291 (N_3291,N_2600,N_2514);
nor U3292 (N_3292,N_2789,N_2643);
nand U3293 (N_3293,N_2934,N_2569);
nor U3294 (N_3294,N_2889,N_2706);
and U3295 (N_3295,N_2701,N_3120);
nor U3296 (N_3296,N_2945,N_2991);
or U3297 (N_3297,N_3054,N_2582);
xor U3298 (N_3298,N_3034,N_2966);
nand U3299 (N_3299,N_2552,N_2610);
or U3300 (N_3300,N_2742,N_2508);
nor U3301 (N_3301,N_3021,N_2720);
nand U3302 (N_3302,N_2501,N_2844);
xor U3303 (N_3303,N_2673,N_3107);
xnor U3304 (N_3304,N_2954,N_2868);
or U3305 (N_3305,N_2544,N_2685);
nand U3306 (N_3306,N_2920,N_2698);
xnor U3307 (N_3307,N_2923,N_2961);
xor U3308 (N_3308,N_3020,N_2831);
xor U3309 (N_3309,N_2853,N_3094);
xnor U3310 (N_3310,N_2629,N_3100);
and U3311 (N_3311,N_2633,N_2506);
or U3312 (N_3312,N_2972,N_2529);
or U3313 (N_3313,N_2775,N_2740);
xor U3314 (N_3314,N_2985,N_2557);
and U3315 (N_3315,N_2536,N_2627);
nor U3316 (N_3316,N_2739,N_2735);
xor U3317 (N_3317,N_2585,N_2834);
or U3318 (N_3318,N_2806,N_2816);
or U3319 (N_3319,N_2952,N_2761);
or U3320 (N_3320,N_2667,N_2858);
or U3321 (N_3321,N_2626,N_2794);
xor U3322 (N_3322,N_2531,N_2955);
and U3323 (N_3323,N_2999,N_2863);
nand U3324 (N_3324,N_2590,N_3060);
and U3325 (N_3325,N_2786,N_3047);
and U3326 (N_3326,N_2820,N_2675);
nor U3327 (N_3327,N_2725,N_2856);
and U3328 (N_3328,N_3007,N_2796);
and U3329 (N_3329,N_2577,N_3002);
xnor U3330 (N_3330,N_2616,N_2946);
nand U3331 (N_3331,N_2948,N_2926);
nor U3332 (N_3332,N_2835,N_3098);
or U3333 (N_3333,N_2519,N_3033);
xor U3334 (N_3334,N_3003,N_2828);
and U3335 (N_3335,N_2509,N_2727);
or U3336 (N_3336,N_2663,N_3074);
nor U3337 (N_3337,N_2771,N_2995);
xnor U3338 (N_3338,N_3086,N_2696);
nor U3339 (N_3339,N_2857,N_2890);
and U3340 (N_3340,N_2809,N_3006);
nand U3341 (N_3341,N_2747,N_2964);
or U3342 (N_3342,N_2543,N_3079);
nor U3343 (N_3343,N_2571,N_2669);
and U3344 (N_3344,N_2594,N_2619);
xnor U3345 (N_3345,N_2823,N_2631);
nor U3346 (N_3346,N_2702,N_2837);
and U3347 (N_3347,N_2865,N_2515);
and U3348 (N_3348,N_3014,N_3070);
and U3349 (N_3349,N_2873,N_2808);
or U3350 (N_3350,N_2661,N_3121);
nand U3351 (N_3351,N_2950,N_2986);
or U3352 (N_3352,N_2847,N_2578);
xor U3353 (N_3353,N_2855,N_2652);
and U3354 (N_3354,N_2615,N_2611);
nand U3355 (N_3355,N_3058,N_2996);
xnor U3356 (N_3356,N_2910,N_2919);
or U3357 (N_3357,N_3104,N_2947);
or U3358 (N_3358,N_2692,N_2840);
nor U3359 (N_3359,N_2979,N_2632);
nand U3360 (N_3360,N_3055,N_2949);
nand U3361 (N_3361,N_2713,N_2596);
xnor U3362 (N_3362,N_3012,N_2524);
nand U3363 (N_3363,N_2612,N_2758);
xnor U3364 (N_3364,N_3066,N_2654);
or U3365 (N_3365,N_2699,N_2943);
nand U3366 (N_3366,N_2993,N_2719);
xnor U3367 (N_3367,N_3083,N_3092);
or U3368 (N_3368,N_2902,N_2682);
or U3369 (N_3369,N_2821,N_2894);
xnor U3370 (N_3370,N_3123,N_3117);
nand U3371 (N_3371,N_2507,N_2580);
nand U3372 (N_3372,N_2520,N_2842);
or U3373 (N_3373,N_2918,N_2568);
or U3374 (N_3374,N_2928,N_2583);
and U3375 (N_3375,N_2556,N_2504);
nor U3376 (N_3376,N_2589,N_2832);
and U3377 (N_3377,N_2772,N_2666);
and U3378 (N_3378,N_2634,N_2653);
nand U3379 (N_3379,N_2687,N_2849);
nor U3380 (N_3380,N_2925,N_2645);
and U3381 (N_3381,N_2812,N_3041);
nor U3382 (N_3382,N_2729,N_2609);
nor U3383 (N_3383,N_2845,N_2592);
and U3384 (N_3384,N_2623,N_2525);
and U3385 (N_3385,N_2795,N_3059);
nor U3386 (N_3386,N_2953,N_2584);
xor U3387 (N_3387,N_2523,N_3078);
and U3388 (N_3388,N_2595,N_3115);
nand U3389 (N_3389,N_2554,N_3049);
and U3390 (N_3390,N_3082,N_3112);
nor U3391 (N_3391,N_3057,N_2709);
nand U3392 (N_3392,N_2780,N_2766);
nand U3393 (N_3393,N_2765,N_2981);
nand U3394 (N_3394,N_3097,N_3008);
nor U3395 (N_3395,N_3085,N_2838);
or U3396 (N_3396,N_2880,N_2730);
nor U3397 (N_3397,N_2637,N_2677);
nor U3398 (N_3398,N_2745,N_2658);
and U3399 (N_3399,N_3030,N_2724);
nor U3400 (N_3400,N_3072,N_2751);
and U3401 (N_3401,N_2718,N_2700);
and U3402 (N_3402,N_2998,N_3106);
and U3403 (N_3403,N_2564,N_2500);
xor U3404 (N_3404,N_2989,N_2714);
nand U3405 (N_3405,N_2676,N_3045);
or U3406 (N_3406,N_2542,N_2572);
xor U3407 (N_3407,N_3018,N_2763);
nor U3408 (N_3408,N_2628,N_2905);
nand U3409 (N_3409,N_3075,N_2801);
nor U3410 (N_3410,N_2505,N_2937);
nor U3411 (N_3411,N_2640,N_2907);
or U3412 (N_3412,N_2829,N_2579);
nand U3413 (N_3413,N_2768,N_2598);
nand U3414 (N_3414,N_2962,N_2917);
nor U3415 (N_3415,N_2841,N_2874);
and U3416 (N_3416,N_2599,N_2527);
or U3417 (N_3417,N_2651,N_2924);
or U3418 (N_3418,N_2749,N_2839);
nand U3419 (N_3419,N_2935,N_2563);
nand U3420 (N_3420,N_2601,N_2912);
xor U3421 (N_3421,N_2638,N_2539);
nand U3422 (N_3422,N_2983,N_2503);
xor U3423 (N_3423,N_2646,N_3009);
and U3424 (N_3424,N_2748,N_2871);
or U3425 (N_3425,N_3000,N_2744);
nor U3426 (N_3426,N_2665,N_2864);
nor U3427 (N_3427,N_3011,N_3067);
or U3428 (N_3428,N_2671,N_2901);
nor U3429 (N_3429,N_3090,N_2659);
or U3430 (N_3430,N_2618,N_2668);
or U3431 (N_3431,N_3091,N_2978);
xor U3432 (N_3432,N_2929,N_2892);
and U3433 (N_3433,N_2546,N_2684);
and U3434 (N_3434,N_2690,N_2710);
or U3435 (N_3435,N_2846,N_2750);
nand U3436 (N_3436,N_2624,N_2731);
xnor U3437 (N_3437,N_2940,N_2747);
nor U3438 (N_3438,N_2875,N_2818);
or U3439 (N_3439,N_2884,N_2546);
and U3440 (N_3440,N_3050,N_2591);
and U3441 (N_3441,N_2977,N_2785);
or U3442 (N_3442,N_2627,N_2500);
or U3443 (N_3443,N_2843,N_2756);
nor U3444 (N_3444,N_3034,N_2581);
or U3445 (N_3445,N_3059,N_2744);
and U3446 (N_3446,N_2552,N_2876);
nor U3447 (N_3447,N_2725,N_3086);
nor U3448 (N_3448,N_3050,N_2830);
or U3449 (N_3449,N_2710,N_2587);
xor U3450 (N_3450,N_2529,N_2830);
nand U3451 (N_3451,N_2814,N_3073);
xnor U3452 (N_3452,N_2714,N_3093);
nor U3453 (N_3453,N_2885,N_2674);
or U3454 (N_3454,N_2628,N_2738);
and U3455 (N_3455,N_2828,N_2899);
nor U3456 (N_3456,N_2689,N_2643);
and U3457 (N_3457,N_2690,N_2806);
xnor U3458 (N_3458,N_2590,N_2670);
nor U3459 (N_3459,N_2633,N_2647);
and U3460 (N_3460,N_2710,N_2657);
nor U3461 (N_3461,N_2985,N_3035);
xnor U3462 (N_3462,N_3083,N_3003);
and U3463 (N_3463,N_3008,N_2660);
xnor U3464 (N_3464,N_2956,N_2531);
or U3465 (N_3465,N_2551,N_2721);
nor U3466 (N_3466,N_2722,N_2591);
and U3467 (N_3467,N_2538,N_2765);
nand U3468 (N_3468,N_2726,N_2655);
nor U3469 (N_3469,N_2672,N_2976);
and U3470 (N_3470,N_2559,N_3072);
xnor U3471 (N_3471,N_2536,N_2920);
xnor U3472 (N_3472,N_2737,N_2539);
nand U3473 (N_3473,N_3000,N_2881);
nor U3474 (N_3474,N_3009,N_2984);
nor U3475 (N_3475,N_2862,N_2866);
or U3476 (N_3476,N_2880,N_2574);
and U3477 (N_3477,N_2520,N_2975);
nor U3478 (N_3478,N_2585,N_2830);
and U3479 (N_3479,N_2659,N_2733);
or U3480 (N_3480,N_3043,N_3077);
xnor U3481 (N_3481,N_2787,N_2889);
or U3482 (N_3482,N_2732,N_3119);
or U3483 (N_3483,N_2619,N_2810);
and U3484 (N_3484,N_2699,N_2760);
xnor U3485 (N_3485,N_2853,N_2859);
nor U3486 (N_3486,N_2657,N_2594);
or U3487 (N_3487,N_2764,N_2982);
xnor U3488 (N_3488,N_3088,N_2599);
or U3489 (N_3489,N_2608,N_2945);
nor U3490 (N_3490,N_3083,N_2778);
or U3491 (N_3491,N_2834,N_2681);
nor U3492 (N_3492,N_2801,N_2874);
nor U3493 (N_3493,N_2643,N_3011);
nor U3494 (N_3494,N_2652,N_2509);
and U3495 (N_3495,N_2713,N_2568);
nand U3496 (N_3496,N_2979,N_2620);
nand U3497 (N_3497,N_2941,N_2505);
nand U3498 (N_3498,N_2844,N_2996);
or U3499 (N_3499,N_2762,N_2849);
or U3500 (N_3500,N_3111,N_2953);
nor U3501 (N_3501,N_3009,N_2889);
or U3502 (N_3502,N_2689,N_2650);
and U3503 (N_3503,N_2952,N_2798);
xor U3504 (N_3504,N_2740,N_2879);
nand U3505 (N_3505,N_2585,N_3035);
xor U3506 (N_3506,N_2706,N_2850);
nand U3507 (N_3507,N_2978,N_2817);
nand U3508 (N_3508,N_2706,N_2903);
nand U3509 (N_3509,N_2539,N_2863);
and U3510 (N_3510,N_2916,N_2862);
xor U3511 (N_3511,N_2684,N_3032);
or U3512 (N_3512,N_2579,N_3117);
or U3513 (N_3513,N_3044,N_2678);
or U3514 (N_3514,N_2589,N_2980);
nand U3515 (N_3515,N_2820,N_2870);
and U3516 (N_3516,N_2625,N_3108);
or U3517 (N_3517,N_2519,N_3110);
nand U3518 (N_3518,N_2544,N_2553);
nor U3519 (N_3519,N_3121,N_2541);
and U3520 (N_3520,N_2974,N_2887);
nand U3521 (N_3521,N_2789,N_2781);
or U3522 (N_3522,N_3033,N_2802);
xnor U3523 (N_3523,N_2993,N_2904);
or U3524 (N_3524,N_2595,N_2724);
xnor U3525 (N_3525,N_2900,N_2786);
xor U3526 (N_3526,N_2808,N_3041);
and U3527 (N_3527,N_2761,N_3051);
nand U3528 (N_3528,N_2777,N_2848);
xnor U3529 (N_3529,N_3047,N_2862);
and U3530 (N_3530,N_3043,N_2522);
nand U3531 (N_3531,N_2678,N_3025);
and U3532 (N_3532,N_2714,N_2748);
or U3533 (N_3533,N_2843,N_2537);
nand U3534 (N_3534,N_2693,N_2765);
or U3535 (N_3535,N_2568,N_2612);
nor U3536 (N_3536,N_2672,N_2935);
nand U3537 (N_3537,N_2946,N_2970);
and U3538 (N_3538,N_2557,N_2944);
xor U3539 (N_3539,N_2579,N_2924);
xor U3540 (N_3540,N_2978,N_2905);
or U3541 (N_3541,N_2927,N_2872);
and U3542 (N_3542,N_2616,N_2909);
nor U3543 (N_3543,N_2902,N_2697);
and U3544 (N_3544,N_2563,N_2726);
or U3545 (N_3545,N_2978,N_2942);
nand U3546 (N_3546,N_2679,N_2870);
nor U3547 (N_3547,N_2766,N_2679);
nor U3548 (N_3548,N_2514,N_2812);
nor U3549 (N_3549,N_3097,N_2683);
nor U3550 (N_3550,N_2900,N_3062);
and U3551 (N_3551,N_3082,N_2745);
xor U3552 (N_3552,N_2696,N_2584);
or U3553 (N_3553,N_3070,N_2803);
or U3554 (N_3554,N_3034,N_2706);
nand U3555 (N_3555,N_2616,N_3041);
nor U3556 (N_3556,N_3038,N_2932);
or U3557 (N_3557,N_3014,N_3013);
or U3558 (N_3558,N_2544,N_3081);
nor U3559 (N_3559,N_2847,N_2955);
xnor U3560 (N_3560,N_2624,N_3091);
xnor U3561 (N_3561,N_3033,N_2943);
or U3562 (N_3562,N_2932,N_2880);
and U3563 (N_3563,N_2909,N_2725);
nor U3564 (N_3564,N_2850,N_3059);
and U3565 (N_3565,N_2942,N_2705);
xor U3566 (N_3566,N_2756,N_2508);
or U3567 (N_3567,N_2660,N_2919);
nor U3568 (N_3568,N_2954,N_2525);
xnor U3569 (N_3569,N_2870,N_2647);
and U3570 (N_3570,N_2971,N_2963);
xnor U3571 (N_3571,N_3119,N_2758);
nor U3572 (N_3572,N_3047,N_3032);
or U3573 (N_3573,N_2890,N_2776);
xnor U3574 (N_3574,N_2868,N_3075);
nand U3575 (N_3575,N_2973,N_2733);
or U3576 (N_3576,N_2859,N_2785);
nor U3577 (N_3577,N_3114,N_3033);
or U3578 (N_3578,N_2870,N_3072);
and U3579 (N_3579,N_2532,N_2814);
nand U3580 (N_3580,N_2514,N_2914);
nand U3581 (N_3581,N_3003,N_2671);
nor U3582 (N_3582,N_2597,N_2870);
or U3583 (N_3583,N_2888,N_2809);
and U3584 (N_3584,N_2623,N_2761);
nand U3585 (N_3585,N_2536,N_2711);
or U3586 (N_3586,N_3058,N_2617);
nor U3587 (N_3587,N_2826,N_2623);
nand U3588 (N_3588,N_2869,N_2873);
xnor U3589 (N_3589,N_2875,N_2530);
nor U3590 (N_3590,N_2830,N_2894);
nor U3591 (N_3591,N_2784,N_2797);
and U3592 (N_3592,N_2892,N_2529);
and U3593 (N_3593,N_3109,N_2636);
nand U3594 (N_3594,N_2647,N_2501);
xnor U3595 (N_3595,N_2610,N_3068);
xnor U3596 (N_3596,N_2918,N_2927);
or U3597 (N_3597,N_2730,N_2656);
nor U3598 (N_3598,N_2896,N_3118);
or U3599 (N_3599,N_2842,N_2956);
nand U3600 (N_3600,N_2537,N_3074);
nor U3601 (N_3601,N_2770,N_2667);
or U3602 (N_3602,N_2634,N_2547);
xnor U3603 (N_3603,N_2904,N_2939);
and U3604 (N_3604,N_2966,N_3065);
nor U3605 (N_3605,N_2785,N_2735);
xnor U3606 (N_3606,N_2718,N_2851);
nor U3607 (N_3607,N_2701,N_3096);
and U3608 (N_3608,N_2671,N_2970);
or U3609 (N_3609,N_2750,N_2814);
or U3610 (N_3610,N_2593,N_2561);
nor U3611 (N_3611,N_2827,N_2933);
and U3612 (N_3612,N_2718,N_2520);
and U3613 (N_3613,N_3056,N_2602);
or U3614 (N_3614,N_2744,N_2575);
xnor U3615 (N_3615,N_2702,N_2886);
xor U3616 (N_3616,N_2664,N_3105);
nor U3617 (N_3617,N_2839,N_2523);
nor U3618 (N_3618,N_2825,N_2620);
nor U3619 (N_3619,N_2987,N_2902);
nor U3620 (N_3620,N_2598,N_2549);
and U3621 (N_3621,N_2932,N_2530);
and U3622 (N_3622,N_2598,N_2984);
nor U3623 (N_3623,N_2982,N_2991);
nand U3624 (N_3624,N_3026,N_3009);
or U3625 (N_3625,N_2739,N_3001);
xnor U3626 (N_3626,N_2645,N_2791);
xor U3627 (N_3627,N_2981,N_2903);
xor U3628 (N_3628,N_2773,N_2898);
xnor U3629 (N_3629,N_2774,N_2889);
and U3630 (N_3630,N_2650,N_2852);
xnor U3631 (N_3631,N_3001,N_2679);
nand U3632 (N_3632,N_2831,N_2511);
nand U3633 (N_3633,N_3049,N_2705);
and U3634 (N_3634,N_3113,N_2525);
or U3635 (N_3635,N_3093,N_2698);
nor U3636 (N_3636,N_2819,N_2685);
nor U3637 (N_3637,N_2901,N_2708);
xnor U3638 (N_3638,N_2633,N_2508);
nor U3639 (N_3639,N_2852,N_2989);
xnor U3640 (N_3640,N_2536,N_2756);
nand U3641 (N_3641,N_2806,N_3008);
or U3642 (N_3642,N_2635,N_2694);
nor U3643 (N_3643,N_3102,N_2699);
xnor U3644 (N_3644,N_2533,N_3103);
or U3645 (N_3645,N_2695,N_3083);
xnor U3646 (N_3646,N_2891,N_2905);
or U3647 (N_3647,N_2574,N_2805);
nor U3648 (N_3648,N_2613,N_2597);
and U3649 (N_3649,N_2827,N_2794);
nand U3650 (N_3650,N_3008,N_2618);
xnor U3651 (N_3651,N_2687,N_2925);
or U3652 (N_3652,N_2655,N_2880);
xnor U3653 (N_3653,N_2588,N_3028);
nand U3654 (N_3654,N_2647,N_2755);
nor U3655 (N_3655,N_2777,N_2675);
and U3656 (N_3656,N_2686,N_2760);
or U3657 (N_3657,N_2776,N_2686);
xnor U3658 (N_3658,N_3091,N_2505);
xor U3659 (N_3659,N_2857,N_3042);
and U3660 (N_3660,N_2563,N_2626);
nand U3661 (N_3661,N_3074,N_3102);
or U3662 (N_3662,N_2930,N_2943);
xnor U3663 (N_3663,N_2943,N_2755);
and U3664 (N_3664,N_3080,N_2731);
or U3665 (N_3665,N_2732,N_3099);
nor U3666 (N_3666,N_2764,N_2890);
nor U3667 (N_3667,N_2805,N_2821);
or U3668 (N_3668,N_2535,N_3034);
or U3669 (N_3669,N_2634,N_2641);
nor U3670 (N_3670,N_2906,N_3094);
nor U3671 (N_3671,N_2989,N_3100);
nor U3672 (N_3672,N_2760,N_2731);
and U3673 (N_3673,N_2729,N_2924);
or U3674 (N_3674,N_2828,N_2750);
or U3675 (N_3675,N_2859,N_2618);
xnor U3676 (N_3676,N_2660,N_2817);
and U3677 (N_3677,N_2898,N_2928);
or U3678 (N_3678,N_2606,N_2660);
or U3679 (N_3679,N_3069,N_2588);
nor U3680 (N_3680,N_3025,N_2864);
nand U3681 (N_3681,N_2869,N_2648);
xor U3682 (N_3682,N_3052,N_3079);
xnor U3683 (N_3683,N_2662,N_2531);
or U3684 (N_3684,N_3081,N_3068);
and U3685 (N_3685,N_2865,N_2878);
or U3686 (N_3686,N_2684,N_3052);
xor U3687 (N_3687,N_3098,N_2814);
nor U3688 (N_3688,N_2935,N_3110);
nand U3689 (N_3689,N_2895,N_3072);
or U3690 (N_3690,N_2665,N_2572);
or U3691 (N_3691,N_2772,N_2671);
and U3692 (N_3692,N_2683,N_2647);
xnor U3693 (N_3693,N_2745,N_2515);
xnor U3694 (N_3694,N_2834,N_2919);
xnor U3695 (N_3695,N_2544,N_2994);
nor U3696 (N_3696,N_2886,N_2951);
or U3697 (N_3697,N_2887,N_2670);
or U3698 (N_3698,N_2532,N_2621);
or U3699 (N_3699,N_2740,N_2560);
nand U3700 (N_3700,N_2597,N_2788);
and U3701 (N_3701,N_2884,N_2684);
xnor U3702 (N_3702,N_2537,N_2543);
nand U3703 (N_3703,N_2933,N_3022);
or U3704 (N_3704,N_3115,N_2744);
nor U3705 (N_3705,N_2561,N_2607);
and U3706 (N_3706,N_2956,N_2642);
and U3707 (N_3707,N_2778,N_2945);
or U3708 (N_3708,N_2750,N_2516);
nand U3709 (N_3709,N_2603,N_3020);
nand U3710 (N_3710,N_2688,N_3065);
xnor U3711 (N_3711,N_2581,N_3040);
nand U3712 (N_3712,N_2688,N_2972);
xnor U3713 (N_3713,N_2963,N_2713);
nor U3714 (N_3714,N_2756,N_3112);
and U3715 (N_3715,N_2959,N_2995);
and U3716 (N_3716,N_3070,N_2962);
nand U3717 (N_3717,N_2500,N_2702);
xor U3718 (N_3718,N_2862,N_2531);
xnor U3719 (N_3719,N_2586,N_2711);
xnor U3720 (N_3720,N_2547,N_3120);
and U3721 (N_3721,N_3029,N_3069);
and U3722 (N_3722,N_2897,N_2600);
xnor U3723 (N_3723,N_3076,N_3049);
or U3724 (N_3724,N_2850,N_2736);
and U3725 (N_3725,N_2974,N_2684);
nand U3726 (N_3726,N_3093,N_3042);
and U3727 (N_3727,N_3051,N_2762);
nor U3728 (N_3728,N_3003,N_2701);
or U3729 (N_3729,N_2836,N_2974);
and U3730 (N_3730,N_3103,N_2590);
nand U3731 (N_3731,N_2716,N_2886);
and U3732 (N_3732,N_2982,N_2769);
xor U3733 (N_3733,N_3078,N_2682);
or U3734 (N_3734,N_2959,N_2640);
and U3735 (N_3735,N_2589,N_2907);
and U3736 (N_3736,N_2795,N_2943);
nor U3737 (N_3737,N_2626,N_2506);
or U3738 (N_3738,N_2538,N_2852);
and U3739 (N_3739,N_2959,N_2509);
and U3740 (N_3740,N_2831,N_2537);
nand U3741 (N_3741,N_2890,N_2667);
nand U3742 (N_3742,N_3116,N_2873);
or U3743 (N_3743,N_2533,N_2971);
nand U3744 (N_3744,N_2857,N_2952);
xnor U3745 (N_3745,N_2771,N_2606);
xnor U3746 (N_3746,N_3123,N_3115);
nand U3747 (N_3747,N_3034,N_2925);
nor U3748 (N_3748,N_2913,N_2919);
nor U3749 (N_3749,N_3057,N_2787);
nand U3750 (N_3750,N_3455,N_3462);
nand U3751 (N_3751,N_3629,N_3696);
and U3752 (N_3752,N_3568,N_3396);
nand U3753 (N_3753,N_3137,N_3173);
nor U3754 (N_3754,N_3418,N_3521);
nor U3755 (N_3755,N_3704,N_3168);
and U3756 (N_3756,N_3698,N_3519);
nor U3757 (N_3757,N_3339,N_3201);
nand U3758 (N_3758,N_3391,N_3524);
and U3759 (N_3759,N_3588,N_3139);
and U3760 (N_3760,N_3196,N_3281);
or U3761 (N_3761,N_3374,N_3152);
and U3762 (N_3762,N_3371,N_3631);
nand U3763 (N_3763,N_3620,N_3270);
or U3764 (N_3764,N_3708,N_3537);
nand U3765 (N_3765,N_3590,N_3660);
nand U3766 (N_3766,N_3197,N_3285);
nand U3767 (N_3767,N_3184,N_3609);
and U3768 (N_3768,N_3233,N_3558);
nor U3769 (N_3769,N_3202,N_3130);
and U3770 (N_3770,N_3439,N_3287);
nand U3771 (N_3771,N_3164,N_3358);
or U3772 (N_3772,N_3487,N_3292);
xnor U3773 (N_3773,N_3236,N_3464);
and U3774 (N_3774,N_3740,N_3195);
and U3775 (N_3775,N_3344,N_3650);
or U3776 (N_3776,N_3315,N_3158);
xor U3777 (N_3777,N_3536,N_3389);
xor U3778 (N_3778,N_3433,N_3509);
xnor U3779 (N_3779,N_3141,N_3526);
nor U3780 (N_3780,N_3730,N_3375);
nand U3781 (N_3781,N_3720,N_3587);
nand U3782 (N_3782,N_3366,N_3557);
nor U3783 (N_3783,N_3484,N_3503);
and U3784 (N_3784,N_3316,N_3299);
xor U3785 (N_3785,N_3486,N_3240);
and U3786 (N_3786,N_3692,N_3129);
and U3787 (N_3787,N_3157,N_3624);
and U3788 (N_3788,N_3435,N_3382);
or U3789 (N_3789,N_3589,N_3518);
nand U3790 (N_3790,N_3289,N_3501);
and U3791 (N_3791,N_3482,N_3125);
and U3792 (N_3792,N_3363,N_3739);
nand U3793 (N_3793,N_3434,N_3512);
or U3794 (N_3794,N_3467,N_3269);
or U3795 (N_3795,N_3662,N_3387);
xor U3796 (N_3796,N_3694,N_3255);
xor U3797 (N_3797,N_3454,N_3697);
nor U3798 (N_3798,N_3528,N_3460);
nor U3799 (N_3799,N_3290,N_3563);
nand U3800 (N_3800,N_3329,N_3659);
nand U3801 (N_3801,N_3428,N_3722);
nor U3802 (N_3802,N_3317,N_3397);
nor U3803 (N_3803,N_3161,N_3733);
nor U3804 (N_3804,N_3407,N_3209);
or U3805 (N_3805,N_3180,N_3525);
xnor U3806 (N_3806,N_3639,N_3472);
nor U3807 (N_3807,N_3737,N_3594);
and U3808 (N_3808,N_3672,N_3386);
nor U3809 (N_3809,N_3146,N_3261);
nand U3810 (N_3810,N_3179,N_3400);
nand U3811 (N_3811,N_3301,N_3716);
xnor U3812 (N_3812,N_3551,N_3309);
xnor U3813 (N_3813,N_3303,N_3187);
or U3814 (N_3814,N_3291,N_3426);
xnor U3815 (N_3815,N_3284,N_3674);
nor U3816 (N_3816,N_3262,N_3468);
or U3817 (N_3817,N_3461,N_3183);
or U3818 (N_3818,N_3547,N_3367);
nor U3819 (N_3819,N_3142,N_3127);
and U3820 (N_3820,N_3627,N_3520);
nor U3821 (N_3821,N_3369,N_3225);
or U3822 (N_3822,N_3295,N_3586);
and U3823 (N_3823,N_3390,N_3268);
nand U3824 (N_3824,N_3610,N_3686);
nand U3825 (N_3825,N_3444,N_3388);
or U3826 (N_3826,N_3505,N_3148);
nor U3827 (N_3827,N_3442,N_3746);
nor U3828 (N_3828,N_3438,N_3178);
xor U3829 (N_3829,N_3326,N_3492);
xnor U3830 (N_3830,N_3741,N_3699);
or U3831 (N_3831,N_3649,N_3241);
or U3832 (N_3832,N_3279,N_3684);
nor U3833 (N_3833,N_3293,N_3381);
nor U3834 (N_3834,N_3258,N_3300);
and U3835 (N_3835,N_3453,N_3565);
and U3836 (N_3836,N_3630,N_3669);
and U3837 (N_3837,N_3147,N_3191);
nand U3838 (N_3838,N_3656,N_3638);
nand U3839 (N_3839,N_3224,N_3530);
nor U3840 (N_3840,N_3711,N_3721);
and U3841 (N_3841,N_3266,N_3393);
xor U3842 (N_3842,N_3600,N_3687);
or U3843 (N_3843,N_3223,N_3471);
nor U3844 (N_3844,N_3320,N_3625);
xnor U3845 (N_3845,N_3443,N_3194);
nor U3846 (N_3846,N_3712,N_3459);
or U3847 (N_3847,N_3569,N_3166);
nor U3848 (N_3848,N_3411,N_3437);
or U3849 (N_3849,N_3465,N_3652);
and U3850 (N_3850,N_3286,N_3377);
xnor U3851 (N_3851,N_3218,N_3481);
and U3852 (N_3852,N_3275,N_3305);
or U3853 (N_3853,N_3477,N_3655);
nor U3854 (N_3854,N_3145,N_3614);
xor U3855 (N_3855,N_3334,N_3661);
nand U3856 (N_3856,N_3582,N_3506);
and U3857 (N_3857,N_3496,N_3342);
xor U3858 (N_3858,N_3634,N_3345);
and U3859 (N_3859,N_3420,N_3507);
nor U3860 (N_3860,N_3497,N_3333);
and U3861 (N_3861,N_3228,N_3608);
nor U3862 (N_3862,N_3237,N_3713);
or U3863 (N_3863,N_3304,N_3748);
or U3864 (N_3864,N_3579,N_3214);
or U3865 (N_3865,N_3250,N_3338);
nand U3866 (N_3866,N_3440,N_3622);
and U3867 (N_3867,N_3384,N_3606);
nor U3868 (N_3868,N_3667,N_3278);
nand U3869 (N_3869,N_3330,N_3226);
xnor U3870 (N_3870,N_3576,N_3372);
xor U3871 (N_3871,N_3283,N_3504);
or U3872 (N_3872,N_3126,N_3522);
nand U3873 (N_3873,N_3364,N_3714);
nand U3874 (N_3874,N_3319,N_3540);
nand U3875 (N_3875,N_3131,N_3539);
or U3876 (N_3876,N_3210,N_3273);
xor U3877 (N_3877,N_3176,N_3402);
nor U3878 (N_3878,N_3355,N_3688);
nand U3879 (N_3879,N_3153,N_3401);
and U3880 (N_3880,N_3679,N_3222);
and U3881 (N_3881,N_3474,N_3331);
and U3882 (N_3882,N_3172,N_3128);
or U3883 (N_3883,N_3668,N_3691);
and U3884 (N_3884,N_3695,N_3412);
and U3885 (N_3885,N_3626,N_3596);
nor U3886 (N_3886,N_3735,N_3405);
nand U3887 (N_3887,N_3533,N_3644);
and U3888 (N_3888,N_3546,N_3419);
nand U3889 (N_3889,N_3404,N_3312);
xor U3890 (N_3890,N_3206,N_3149);
and U3891 (N_3891,N_3370,N_3188);
or U3892 (N_3892,N_3406,N_3570);
nand U3893 (N_3893,N_3246,N_3318);
or U3894 (N_3894,N_3361,N_3595);
nor U3895 (N_3895,N_3532,N_3616);
or U3896 (N_3896,N_3227,N_3591);
or U3897 (N_3897,N_3621,N_3491);
and U3898 (N_3898,N_3365,N_3445);
nand U3899 (N_3899,N_3463,N_3478);
or U3900 (N_3900,N_3257,N_3346);
and U3901 (N_3901,N_3550,N_3671);
and U3902 (N_3902,N_3336,N_3651);
nor U3903 (N_3903,N_3607,N_3494);
nand U3904 (N_3904,N_3562,N_3154);
and U3905 (N_3905,N_3357,N_3171);
nand U3906 (N_3906,N_3552,N_3205);
nor U3907 (N_3907,N_3378,N_3220);
xor U3908 (N_3908,N_3360,N_3738);
nor U3909 (N_3909,N_3272,N_3677);
and U3910 (N_3910,N_3527,N_3643);
nor U3911 (N_3911,N_3162,N_3208);
and U3912 (N_3912,N_3362,N_3637);
or U3913 (N_3913,N_3247,N_3203);
nor U3914 (N_3914,N_3423,N_3383);
nor U3915 (N_3915,N_3466,N_3151);
or U3916 (N_3916,N_3654,N_3658);
or U3917 (N_3917,N_3430,N_3717);
xor U3918 (N_3918,N_3745,N_3580);
and U3919 (N_3919,N_3617,N_3376);
nor U3920 (N_3920,N_3488,N_3581);
and U3921 (N_3921,N_3310,N_3545);
xnor U3922 (N_3922,N_3215,N_3700);
nand U3923 (N_3923,N_3690,N_3709);
or U3924 (N_3924,N_3186,N_3200);
xnor U3925 (N_3925,N_3743,N_3447);
or U3926 (N_3926,N_3256,N_3458);
nor U3927 (N_3927,N_3707,N_3603);
or U3928 (N_3928,N_3598,N_3744);
or U3929 (N_3929,N_3409,N_3410);
and U3930 (N_3930,N_3475,N_3456);
nand U3931 (N_3931,N_3457,N_3192);
nor U3932 (N_3932,N_3726,N_3559);
xor U3933 (N_3933,N_3238,N_3216);
or U3934 (N_3934,N_3615,N_3483);
or U3935 (N_3935,N_3259,N_3427);
nand U3936 (N_3936,N_3647,N_3431);
nor U3937 (N_3937,N_3633,N_3623);
nand U3938 (N_3938,N_3715,N_3432);
nand U3939 (N_3939,N_3544,N_3140);
or U3940 (N_3940,N_3719,N_3543);
and U3941 (N_3941,N_3710,N_3156);
nor U3942 (N_3942,N_3498,N_3325);
or U3943 (N_3943,N_3231,N_3341);
and U3944 (N_3944,N_3676,N_3198);
nor U3945 (N_3945,N_3485,N_3324);
or U3946 (N_3946,N_3235,N_3599);
and U3947 (N_3947,N_3703,N_3619);
xor U3948 (N_3948,N_3251,N_3514);
xor U3949 (N_3949,N_3648,N_3601);
nand U3950 (N_3950,N_3340,N_3204);
nand U3951 (N_3951,N_3480,N_3332);
nand U3952 (N_3952,N_3189,N_3605);
and U3953 (N_3953,N_3451,N_3239);
xnor U3954 (N_3954,N_3260,N_3354);
or U3955 (N_3955,N_3274,N_3664);
nand U3956 (N_3956,N_3727,N_3271);
nand U3957 (N_3957,N_3470,N_3243);
nor U3958 (N_3958,N_3327,N_3379);
and U3959 (N_3959,N_3348,N_3288);
nand U3960 (N_3960,N_3573,N_3489);
nor U3961 (N_3961,N_3693,N_3701);
nor U3962 (N_3962,N_3294,N_3181);
xor U3963 (N_3963,N_3385,N_3725);
xor U3964 (N_3964,N_3408,N_3160);
xor U3965 (N_3965,N_3252,N_3495);
nand U3966 (N_3966,N_3473,N_3207);
and U3967 (N_3967,N_3297,N_3417);
nand U3968 (N_3968,N_3185,N_3135);
xnor U3969 (N_3969,N_3567,N_3490);
nand U3970 (N_3970,N_3542,N_3734);
nand U3971 (N_3971,N_3469,N_3585);
nand U3972 (N_3972,N_3531,N_3229);
nor U3973 (N_3973,N_3612,N_3347);
and U3974 (N_3974,N_3296,N_3429);
xor U3975 (N_3975,N_3403,N_3584);
or U3976 (N_3976,N_3602,N_3618);
xor U3977 (N_3977,N_3450,N_3555);
xnor U3978 (N_3978,N_3307,N_3636);
nor U3979 (N_3979,N_3380,N_3425);
and U3980 (N_3980,N_3446,N_3513);
nor U3981 (N_3981,N_3583,N_3508);
nand U3982 (N_3982,N_3144,N_3199);
nor U3983 (N_3983,N_3165,N_3424);
xnor U3984 (N_3984,N_3337,N_3723);
nor U3985 (N_3985,N_3449,N_3311);
nand U3986 (N_3986,N_3645,N_3133);
or U3987 (N_3987,N_3553,N_3675);
nor U3988 (N_3988,N_3175,N_3232);
nand U3989 (N_3989,N_3242,N_3592);
or U3990 (N_3990,N_3663,N_3352);
xnor U3991 (N_3991,N_3155,N_3476);
and U3992 (N_3992,N_3276,N_3234);
nand U3993 (N_3993,N_3193,N_3323);
xor U3994 (N_3994,N_3136,N_3577);
xor U3995 (N_3995,N_3705,N_3499);
or U3996 (N_3996,N_3143,N_3516);
or U3997 (N_3997,N_3416,N_3441);
nor U3998 (N_3998,N_3217,N_3732);
and U3999 (N_3999,N_3670,N_3306);
or U4000 (N_4000,N_3150,N_3353);
xor U4001 (N_4001,N_3502,N_3138);
nand U4002 (N_4002,N_3302,N_3373);
and U4003 (N_4003,N_3398,N_3736);
nand U4004 (N_4004,N_3190,N_3574);
nor U4005 (N_4005,N_3263,N_3448);
nand U4006 (N_4006,N_3628,N_3182);
or U4007 (N_4007,N_3249,N_3349);
nand U4008 (N_4008,N_3724,N_3666);
nand U4009 (N_4009,N_3604,N_3685);
xor U4010 (N_4010,N_3523,N_3493);
and U4011 (N_4011,N_3350,N_3510);
or U4012 (N_4012,N_3665,N_3728);
or U4013 (N_4013,N_3174,N_3575);
or U4014 (N_4014,N_3566,N_3702);
or U4015 (N_4015,N_3248,N_3298);
or U4016 (N_4016,N_3556,N_3395);
nand U4017 (N_4017,N_3632,N_3351);
nand U4018 (N_4018,N_3548,N_3535);
or U4019 (N_4019,N_3515,N_3541);
nand U4020 (N_4020,N_3511,N_3163);
nor U4021 (N_4021,N_3265,N_3635);
nor U4022 (N_4022,N_3413,N_3322);
nor U4023 (N_4023,N_3641,N_3731);
xnor U4024 (N_4024,N_3132,N_3421);
xor U4025 (N_4025,N_3177,N_3593);
nor U4026 (N_4026,N_3282,N_3706);
xnor U4027 (N_4027,N_3529,N_3747);
nor U4028 (N_4028,N_3392,N_3356);
nor U4029 (N_4029,N_3673,N_3749);
or U4030 (N_4030,N_3313,N_3729);
and U4031 (N_4031,N_3742,N_3245);
xnor U4032 (N_4032,N_3682,N_3399);
or U4033 (N_4033,N_3335,N_3640);
or U4034 (N_4034,N_3653,N_3267);
nand U4035 (N_4035,N_3212,N_3718);
nand U4036 (N_4036,N_3328,N_3230);
and U4037 (N_4037,N_3415,N_3169);
nand U4038 (N_4038,N_3689,N_3452);
xnor U4039 (N_4039,N_3611,N_3549);
xor U4040 (N_4040,N_3646,N_3642);
and U4041 (N_4041,N_3134,N_3564);
xor U4042 (N_4042,N_3479,N_3534);
or U4043 (N_4043,N_3683,N_3254);
nor U4044 (N_4044,N_3554,N_3500);
nor U4045 (N_4045,N_3170,N_3680);
and U4046 (N_4046,N_3221,N_3422);
xor U4047 (N_4047,N_3277,N_3213);
nor U4048 (N_4048,N_3681,N_3167);
nand U4049 (N_4049,N_3264,N_3572);
nand U4050 (N_4050,N_3560,N_3538);
nand U4051 (N_4051,N_3517,N_3561);
xor U4052 (N_4052,N_3368,N_3343);
nor U4053 (N_4053,N_3211,N_3578);
nor U4054 (N_4054,N_3359,N_3613);
nor U4055 (N_4055,N_3678,N_3597);
nor U4056 (N_4056,N_3321,N_3414);
nand U4057 (N_4057,N_3159,N_3394);
nand U4058 (N_4058,N_3280,N_3657);
and U4059 (N_4059,N_3308,N_3436);
nor U4060 (N_4060,N_3219,N_3244);
nand U4061 (N_4061,N_3253,N_3571);
or U4062 (N_4062,N_3314,N_3741);
or U4063 (N_4063,N_3489,N_3324);
xor U4064 (N_4064,N_3659,N_3427);
nand U4065 (N_4065,N_3296,N_3180);
nor U4066 (N_4066,N_3749,N_3637);
and U4067 (N_4067,N_3378,N_3686);
and U4068 (N_4068,N_3373,N_3520);
xnor U4069 (N_4069,N_3439,N_3715);
xor U4070 (N_4070,N_3245,N_3662);
nand U4071 (N_4071,N_3207,N_3183);
and U4072 (N_4072,N_3172,N_3639);
or U4073 (N_4073,N_3534,N_3251);
xor U4074 (N_4074,N_3431,N_3421);
xnor U4075 (N_4075,N_3186,N_3318);
nand U4076 (N_4076,N_3449,N_3547);
nor U4077 (N_4077,N_3155,N_3667);
nand U4078 (N_4078,N_3632,N_3335);
nor U4079 (N_4079,N_3569,N_3139);
and U4080 (N_4080,N_3214,N_3304);
or U4081 (N_4081,N_3532,N_3607);
nand U4082 (N_4082,N_3573,N_3319);
xor U4083 (N_4083,N_3288,N_3318);
xnor U4084 (N_4084,N_3532,N_3149);
and U4085 (N_4085,N_3552,N_3684);
xor U4086 (N_4086,N_3449,N_3206);
nor U4087 (N_4087,N_3449,N_3281);
or U4088 (N_4088,N_3165,N_3555);
and U4089 (N_4089,N_3268,N_3369);
xnor U4090 (N_4090,N_3378,N_3126);
xnor U4091 (N_4091,N_3602,N_3748);
or U4092 (N_4092,N_3580,N_3699);
or U4093 (N_4093,N_3429,N_3316);
nor U4094 (N_4094,N_3476,N_3580);
and U4095 (N_4095,N_3512,N_3242);
and U4096 (N_4096,N_3511,N_3694);
nand U4097 (N_4097,N_3374,N_3550);
nand U4098 (N_4098,N_3746,N_3657);
nand U4099 (N_4099,N_3640,N_3611);
nor U4100 (N_4100,N_3449,N_3443);
xnor U4101 (N_4101,N_3170,N_3145);
or U4102 (N_4102,N_3642,N_3127);
nand U4103 (N_4103,N_3664,N_3475);
nor U4104 (N_4104,N_3280,N_3468);
or U4105 (N_4105,N_3404,N_3233);
and U4106 (N_4106,N_3560,N_3541);
or U4107 (N_4107,N_3563,N_3645);
nand U4108 (N_4108,N_3559,N_3596);
nand U4109 (N_4109,N_3244,N_3675);
and U4110 (N_4110,N_3450,N_3149);
or U4111 (N_4111,N_3483,N_3135);
nor U4112 (N_4112,N_3624,N_3407);
and U4113 (N_4113,N_3131,N_3404);
nor U4114 (N_4114,N_3143,N_3609);
xor U4115 (N_4115,N_3256,N_3631);
or U4116 (N_4116,N_3539,N_3274);
xnor U4117 (N_4117,N_3136,N_3508);
nand U4118 (N_4118,N_3685,N_3543);
nor U4119 (N_4119,N_3348,N_3628);
or U4120 (N_4120,N_3235,N_3660);
nor U4121 (N_4121,N_3600,N_3712);
xnor U4122 (N_4122,N_3725,N_3568);
nand U4123 (N_4123,N_3271,N_3374);
or U4124 (N_4124,N_3441,N_3403);
or U4125 (N_4125,N_3270,N_3567);
nand U4126 (N_4126,N_3669,N_3459);
or U4127 (N_4127,N_3397,N_3649);
nand U4128 (N_4128,N_3532,N_3623);
nand U4129 (N_4129,N_3597,N_3705);
nand U4130 (N_4130,N_3171,N_3251);
nor U4131 (N_4131,N_3395,N_3130);
or U4132 (N_4132,N_3577,N_3368);
xor U4133 (N_4133,N_3541,N_3322);
xnor U4134 (N_4134,N_3671,N_3312);
and U4135 (N_4135,N_3395,N_3513);
or U4136 (N_4136,N_3603,N_3415);
nand U4137 (N_4137,N_3228,N_3501);
or U4138 (N_4138,N_3391,N_3747);
xor U4139 (N_4139,N_3236,N_3738);
and U4140 (N_4140,N_3312,N_3287);
and U4141 (N_4141,N_3165,N_3327);
xor U4142 (N_4142,N_3449,N_3286);
xnor U4143 (N_4143,N_3435,N_3369);
nand U4144 (N_4144,N_3640,N_3695);
xnor U4145 (N_4145,N_3561,N_3615);
nor U4146 (N_4146,N_3476,N_3355);
nand U4147 (N_4147,N_3560,N_3440);
and U4148 (N_4148,N_3639,N_3327);
xor U4149 (N_4149,N_3474,N_3400);
xnor U4150 (N_4150,N_3655,N_3202);
nor U4151 (N_4151,N_3276,N_3310);
xnor U4152 (N_4152,N_3477,N_3414);
nor U4153 (N_4153,N_3247,N_3518);
or U4154 (N_4154,N_3359,N_3409);
and U4155 (N_4155,N_3434,N_3217);
and U4156 (N_4156,N_3468,N_3718);
and U4157 (N_4157,N_3678,N_3142);
nor U4158 (N_4158,N_3152,N_3687);
and U4159 (N_4159,N_3180,N_3288);
nand U4160 (N_4160,N_3684,N_3602);
nand U4161 (N_4161,N_3601,N_3395);
xnor U4162 (N_4162,N_3210,N_3208);
and U4163 (N_4163,N_3490,N_3616);
or U4164 (N_4164,N_3176,N_3158);
nand U4165 (N_4165,N_3378,N_3218);
nand U4166 (N_4166,N_3367,N_3360);
xor U4167 (N_4167,N_3464,N_3332);
nand U4168 (N_4168,N_3337,N_3298);
and U4169 (N_4169,N_3681,N_3261);
nand U4170 (N_4170,N_3715,N_3504);
or U4171 (N_4171,N_3278,N_3367);
or U4172 (N_4172,N_3736,N_3583);
or U4173 (N_4173,N_3367,N_3613);
xnor U4174 (N_4174,N_3326,N_3598);
xor U4175 (N_4175,N_3250,N_3470);
xor U4176 (N_4176,N_3152,N_3471);
nor U4177 (N_4177,N_3150,N_3365);
xnor U4178 (N_4178,N_3136,N_3233);
nand U4179 (N_4179,N_3315,N_3466);
or U4180 (N_4180,N_3526,N_3209);
nor U4181 (N_4181,N_3464,N_3705);
nand U4182 (N_4182,N_3422,N_3457);
and U4183 (N_4183,N_3363,N_3503);
xnor U4184 (N_4184,N_3361,N_3270);
xor U4185 (N_4185,N_3666,N_3195);
nand U4186 (N_4186,N_3689,N_3385);
xor U4187 (N_4187,N_3182,N_3584);
or U4188 (N_4188,N_3379,N_3255);
nor U4189 (N_4189,N_3357,N_3165);
or U4190 (N_4190,N_3170,N_3361);
or U4191 (N_4191,N_3305,N_3220);
nor U4192 (N_4192,N_3238,N_3600);
xnor U4193 (N_4193,N_3653,N_3255);
and U4194 (N_4194,N_3160,N_3395);
or U4195 (N_4195,N_3155,N_3279);
nand U4196 (N_4196,N_3202,N_3303);
nor U4197 (N_4197,N_3610,N_3334);
nor U4198 (N_4198,N_3382,N_3246);
xor U4199 (N_4199,N_3171,N_3157);
and U4200 (N_4200,N_3502,N_3220);
xor U4201 (N_4201,N_3523,N_3628);
nor U4202 (N_4202,N_3311,N_3541);
or U4203 (N_4203,N_3369,N_3552);
and U4204 (N_4204,N_3551,N_3279);
nor U4205 (N_4205,N_3651,N_3551);
nor U4206 (N_4206,N_3280,N_3146);
and U4207 (N_4207,N_3208,N_3373);
nand U4208 (N_4208,N_3692,N_3414);
nor U4209 (N_4209,N_3506,N_3693);
xor U4210 (N_4210,N_3316,N_3536);
and U4211 (N_4211,N_3516,N_3336);
nand U4212 (N_4212,N_3501,N_3343);
or U4213 (N_4213,N_3659,N_3414);
and U4214 (N_4214,N_3325,N_3698);
or U4215 (N_4215,N_3655,N_3399);
nor U4216 (N_4216,N_3182,N_3427);
or U4217 (N_4217,N_3343,N_3741);
or U4218 (N_4218,N_3255,N_3649);
and U4219 (N_4219,N_3448,N_3386);
nor U4220 (N_4220,N_3250,N_3330);
or U4221 (N_4221,N_3740,N_3267);
nor U4222 (N_4222,N_3702,N_3472);
nand U4223 (N_4223,N_3328,N_3172);
nor U4224 (N_4224,N_3452,N_3158);
and U4225 (N_4225,N_3470,N_3531);
or U4226 (N_4226,N_3386,N_3283);
nor U4227 (N_4227,N_3615,N_3286);
nand U4228 (N_4228,N_3198,N_3265);
or U4229 (N_4229,N_3287,N_3269);
xnor U4230 (N_4230,N_3507,N_3672);
and U4231 (N_4231,N_3217,N_3610);
xnor U4232 (N_4232,N_3300,N_3205);
and U4233 (N_4233,N_3387,N_3238);
nor U4234 (N_4234,N_3575,N_3252);
nand U4235 (N_4235,N_3342,N_3472);
or U4236 (N_4236,N_3162,N_3145);
and U4237 (N_4237,N_3628,N_3698);
nor U4238 (N_4238,N_3276,N_3237);
nand U4239 (N_4239,N_3695,N_3217);
nor U4240 (N_4240,N_3687,N_3150);
nor U4241 (N_4241,N_3578,N_3382);
nor U4242 (N_4242,N_3703,N_3234);
and U4243 (N_4243,N_3275,N_3453);
or U4244 (N_4244,N_3327,N_3247);
nor U4245 (N_4245,N_3280,N_3593);
and U4246 (N_4246,N_3198,N_3662);
nand U4247 (N_4247,N_3400,N_3500);
nand U4248 (N_4248,N_3481,N_3213);
xor U4249 (N_4249,N_3582,N_3504);
xnor U4250 (N_4250,N_3446,N_3288);
and U4251 (N_4251,N_3214,N_3660);
nand U4252 (N_4252,N_3511,N_3543);
nor U4253 (N_4253,N_3256,N_3586);
xnor U4254 (N_4254,N_3736,N_3408);
or U4255 (N_4255,N_3405,N_3745);
or U4256 (N_4256,N_3260,N_3715);
xnor U4257 (N_4257,N_3570,N_3639);
nor U4258 (N_4258,N_3279,N_3458);
nand U4259 (N_4259,N_3399,N_3358);
nand U4260 (N_4260,N_3380,N_3573);
or U4261 (N_4261,N_3528,N_3477);
xnor U4262 (N_4262,N_3593,N_3539);
nor U4263 (N_4263,N_3700,N_3746);
nand U4264 (N_4264,N_3509,N_3731);
nor U4265 (N_4265,N_3597,N_3646);
nand U4266 (N_4266,N_3336,N_3550);
xnor U4267 (N_4267,N_3662,N_3205);
nor U4268 (N_4268,N_3473,N_3489);
or U4269 (N_4269,N_3692,N_3554);
xnor U4270 (N_4270,N_3555,N_3158);
or U4271 (N_4271,N_3448,N_3435);
and U4272 (N_4272,N_3229,N_3700);
xnor U4273 (N_4273,N_3628,N_3595);
and U4274 (N_4274,N_3542,N_3701);
or U4275 (N_4275,N_3263,N_3647);
or U4276 (N_4276,N_3327,N_3311);
nor U4277 (N_4277,N_3320,N_3246);
nand U4278 (N_4278,N_3378,N_3190);
nand U4279 (N_4279,N_3425,N_3731);
or U4280 (N_4280,N_3622,N_3138);
nor U4281 (N_4281,N_3388,N_3458);
nand U4282 (N_4282,N_3254,N_3375);
and U4283 (N_4283,N_3326,N_3553);
nor U4284 (N_4284,N_3705,N_3396);
nor U4285 (N_4285,N_3666,N_3630);
nor U4286 (N_4286,N_3517,N_3418);
xnor U4287 (N_4287,N_3515,N_3442);
nand U4288 (N_4288,N_3640,N_3577);
nor U4289 (N_4289,N_3597,N_3287);
nor U4290 (N_4290,N_3393,N_3259);
nor U4291 (N_4291,N_3188,N_3738);
nor U4292 (N_4292,N_3585,N_3583);
nor U4293 (N_4293,N_3632,N_3294);
nor U4294 (N_4294,N_3279,N_3443);
xnor U4295 (N_4295,N_3729,N_3292);
xor U4296 (N_4296,N_3239,N_3220);
and U4297 (N_4297,N_3513,N_3492);
or U4298 (N_4298,N_3557,N_3523);
nor U4299 (N_4299,N_3326,N_3139);
or U4300 (N_4300,N_3131,N_3585);
nor U4301 (N_4301,N_3422,N_3335);
nor U4302 (N_4302,N_3188,N_3677);
nor U4303 (N_4303,N_3475,N_3662);
xor U4304 (N_4304,N_3206,N_3225);
nor U4305 (N_4305,N_3413,N_3441);
nor U4306 (N_4306,N_3589,N_3404);
nor U4307 (N_4307,N_3401,N_3125);
nor U4308 (N_4308,N_3316,N_3359);
or U4309 (N_4309,N_3273,N_3252);
nor U4310 (N_4310,N_3494,N_3724);
or U4311 (N_4311,N_3313,N_3507);
nand U4312 (N_4312,N_3234,N_3298);
and U4313 (N_4313,N_3675,N_3704);
and U4314 (N_4314,N_3192,N_3364);
xor U4315 (N_4315,N_3566,N_3206);
and U4316 (N_4316,N_3536,N_3153);
xnor U4317 (N_4317,N_3680,N_3498);
or U4318 (N_4318,N_3374,N_3594);
xor U4319 (N_4319,N_3290,N_3317);
or U4320 (N_4320,N_3535,N_3680);
nor U4321 (N_4321,N_3333,N_3336);
nand U4322 (N_4322,N_3530,N_3185);
xnor U4323 (N_4323,N_3144,N_3607);
nor U4324 (N_4324,N_3425,N_3745);
or U4325 (N_4325,N_3379,N_3653);
xor U4326 (N_4326,N_3213,N_3647);
and U4327 (N_4327,N_3700,N_3475);
nand U4328 (N_4328,N_3140,N_3610);
or U4329 (N_4329,N_3187,N_3134);
nor U4330 (N_4330,N_3239,N_3739);
xor U4331 (N_4331,N_3201,N_3522);
and U4332 (N_4332,N_3591,N_3176);
or U4333 (N_4333,N_3229,N_3316);
xor U4334 (N_4334,N_3597,N_3602);
nand U4335 (N_4335,N_3484,N_3464);
nor U4336 (N_4336,N_3534,N_3375);
and U4337 (N_4337,N_3173,N_3536);
and U4338 (N_4338,N_3488,N_3301);
xor U4339 (N_4339,N_3576,N_3231);
or U4340 (N_4340,N_3291,N_3545);
or U4341 (N_4341,N_3445,N_3131);
xnor U4342 (N_4342,N_3381,N_3249);
nor U4343 (N_4343,N_3364,N_3602);
nand U4344 (N_4344,N_3300,N_3479);
nor U4345 (N_4345,N_3395,N_3608);
xor U4346 (N_4346,N_3653,N_3679);
and U4347 (N_4347,N_3482,N_3377);
nand U4348 (N_4348,N_3397,N_3580);
nand U4349 (N_4349,N_3619,N_3668);
and U4350 (N_4350,N_3527,N_3362);
or U4351 (N_4351,N_3238,N_3591);
xnor U4352 (N_4352,N_3170,N_3605);
nor U4353 (N_4353,N_3614,N_3400);
xnor U4354 (N_4354,N_3126,N_3306);
xnor U4355 (N_4355,N_3396,N_3615);
xnor U4356 (N_4356,N_3704,N_3219);
nor U4357 (N_4357,N_3688,N_3385);
xnor U4358 (N_4358,N_3363,N_3179);
and U4359 (N_4359,N_3366,N_3376);
nand U4360 (N_4360,N_3720,N_3260);
nand U4361 (N_4361,N_3318,N_3344);
and U4362 (N_4362,N_3709,N_3190);
and U4363 (N_4363,N_3688,N_3449);
and U4364 (N_4364,N_3272,N_3434);
nand U4365 (N_4365,N_3663,N_3570);
xor U4366 (N_4366,N_3693,N_3427);
nor U4367 (N_4367,N_3128,N_3213);
nor U4368 (N_4368,N_3190,N_3686);
and U4369 (N_4369,N_3534,N_3364);
and U4370 (N_4370,N_3481,N_3445);
or U4371 (N_4371,N_3528,N_3284);
nor U4372 (N_4372,N_3182,N_3326);
and U4373 (N_4373,N_3283,N_3333);
xor U4374 (N_4374,N_3409,N_3207);
or U4375 (N_4375,N_3991,N_4249);
xor U4376 (N_4376,N_4011,N_4087);
or U4377 (N_4377,N_3796,N_4278);
and U4378 (N_4378,N_4136,N_4041);
or U4379 (N_4379,N_3975,N_4072);
xnor U4380 (N_4380,N_3876,N_4150);
nor U4381 (N_4381,N_4173,N_4361);
nor U4382 (N_4382,N_4130,N_3812);
nor U4383 (N_4383,N_3985,N_4276);
nor U4384 (N_4384,N_4143,N_3780);
and U4385 (N_4385,N_4074,N_3768);
nand U4386 (N_4386,N_3895,N_4079);
nor U4387 (N_4387,N_4201,N_3924);
and U4388 (N_4388,N_3830,N_3855);
or U4389 (N_4389,N_3996,N_4092);
and U4390 (N_4390,N_4005,N_3837);
or U4391 (N_4391,N_3937,N_4312);
nor U4392 (N_4392,N_4071,N_3992);
and U4393 (N_4393,N_4208,N_3874);
xor U4394 (N_4394,N_4162,N_4367);
or U4395 (N_4395,N_4153,N_4324);
nor U4396 (N_4396,N_3809,N_4023);
and U4397 (N_4397,N_3834,N_3930);
or U4398 (N_4398,N_4206,N_4047);
and U4399 (N_4399,N_4100,N_4154);
xnor U4400 (N_4400,N_3972,N_3964);
or U4401 (N_4401,N_3989,N_3841);
nor U4402 (N_4402,N_3944,N_4089);
nand U4403 (N_4403,N_4172,N_4081);
and U4404 (N_4404,N_3848,N_4053);
nor U4405 (N_4405,N_4068,N_3922);
and U4406 (N_4406,N_3808,N_4262);
xor U4407 (N_4407,N_4067,N_3942);
or U4408 (N_4408,N_3773,N_4106);
or U4409 (N_4409,N_3798,N_4204);
nor U4410 (N_4410,N_4099,N_3788);
nor U4411 (N_4411,N_4113,N_4165);
and U4412 (N_4412,N_3949,N_3760);
nor U4413 (N_4413,N_4066,N_4303);
nand U4414 (N_4414,N_4061,N_4024);
and U4415 (N_4415,N_3779,N_3983);
or U4416 (N_4416,N_4123,N_4213);
nand U4417 (N_4417,N_4097,N_4356);
and U4418 (N_4418,N_4290,N_4228);
xor U4419 (N_4419,N_4001,N_4245);
nor U4420 (N_4420,N_4317,N_3915);
or U4421 (N_4421,N_4372,N_4117);
nand U4422 (N_4422,N_4216,N_4291);
nand U4423 (N_4423,N_4225,N_4252);
xnor U4424 (N_4424,N_3884,N_3755);
nor U4425 (N_4425,N_4313,N_3952);
nor U4426 (N_4426,N_4366,N_4272);
nand U4427 (N_4427,N_4155,N_4301);
xor U4428 (N_4428,N_4064,N_4345);
nand U4429 (N_4429,N_4112,N_4084);
nand U4430 (N_4430,N_4088,N_3901);
xor U4431 (N_4431,N_4141,N_3849);
xor U4432 (N_4432,N_3894,N_4114);
nand U4433 (N_4433,N_4007,N_3969);
nor U4434 (N_4434,N_4027,N_4057);
nor U4435 (N_4435,N_4080,N_4120);
nand U4436 (N_4436,N_4355,N_4350);
or U4437 (N_4437,N_4091,N_3804);
nand U4438 (N_4438,N_4012,N_3977);
or U4439 (N_4439,N_4077,N_4287);
xor U4440 (N_4440,N_4098,N_4168);
and U4441 (N_4441,N_4016,N_4314);
and U4442 (N_4442,N_3858,N_3869);
nor U4443 (N_4443,N_3903,N_4368);
and U4444 (N_4444,N_3769,N_4343);
nor U4445 (N_4445,N_4248,N_4111);
nand U4446 (N_4446,N_4264,N_4184);
and U4447 (N_4447,N_3854,N_4363);
xor U4448 (N_4448,N_4360,N_3821);
xnor U4449 (N_4449,N_4102,N_4019);
nor U4450 (N_4450,N_3898,N_3963);
and U4451 (N_4451,N_4170,N_4175);
nand U4452 (N_4452,N_3899,N_3840);
xnor U4453 (N_4453,N_3851,N_3960);
or U4454 (N_4454,N_3881,N_3806);
xnor U4455 (N_4455,N_4302,N_4339);
nand U4456 (N_4456,N_4127,N_3973);
xor U4457 (N_4457,N_3825,N_4186);
or U4458 (N_4458,N_4199,N_4219);
nor U4459 (N_4459,N_4193,N_3792);
xor U4460 (N_4460,N_4212,N_4103);
and U4461 (N_4461,N_4348,N_4298);
or U4462 (N_4462,N_4310,N_3934);
xnor U4463 (N_4463,N_4347,N_4255);
nor U4464 (N_4464,N_3988,N_3998);
xnor U4465 (N_4465,N_4261,N_4257);
nor U4466 (N_4466,N_3883,N_3896);
nand U4467 (N_4467,N_3865,N_4236);
and U4468 (N_4468,N_3823,N_3947);
xnor U4469 (N_4469,N_3824,N_3868);
and U4470 (N_4470,N_3761,N_4226);
xnor U4471 (N_4471,N_3890,N_4002);
or U4472 (N_4472,N_3810,N_3800);
or U4473 (N_4473,N_4271,N_3897);
xnor U4474 (N_4474,N_4200,N_4029);
nand U4475 (N_4475,N_4144,N_3891);
and U4476 (N_4476,N_3911,N_4279);
nor U4477 (N_4477,N_4306,N_4233);
xnor U4478 (N_4478,N_4283,N_4058);
nor U4479 (N_4479,N_4056,N_3958);
xnor U4480 (N_4480,N_4232,N_4326);
and U4481 (N_4481,N_4185,N_4293);
xor U4482 (N_4482,N_4222,N_4282);
and U4483 (N_4483,N_4335,N_4353);
nor U4484 (N_4484,N_4296,N_3757);
or U4485 (N_4485,N_4336,N_3965);
xor U4486 (N_4486,N_4266,N_4297);
or U4487 (N_4487,N_4189,N_4094);
and U4488 (N_4488,N_4115,N_4256);
and U4489 (N_4489,N_4049,N_4242);
and U4490 (N_4490,N_3927,N_3926);
or U4491 (N_4491,N_4124,N_4331);
nand U4492 (N_4492,N_4018,N_4000);
xor U4493 (N_4493,N_3906,N_3940);
or U4494 (N_4494,N_4258,N_3815);
and U4495 (N_4495,N_4251,N_4122);
or U4496 (N_4496,N_4036,N_4260);
xor U4497 (N_4497,N_4359,N_4082);
or U4498 (N_4498,N_4017,N_3818);
xor U4499 (N_4499,N_4322,N_4161);
nor U4500 (N_4500,N_4022,N_3879);
xor U4501 (N_4501,N_4215,N_4070);
nand U4502 (N_4502,N_4054,N_3776);
nor U4503 (N_4503,N_4181,N_3982);
nand U4504 (N_4504,N_3900,N_4138);
nor U4505 (N_4505,N_4093,N_3756);
xnor U4506 (N_4506,N_3939,N_3893);
nand U4507 (N_4507,N_3902,N_4316);
xnor U4508 (N_4508,N_3850,N_4183);
nor U4509 (N_4509,N_3953,N_4267);
nor U4510 (N_4510,N_4220,N_4129);
nand U4511 (N_4511,N_4243,N_4163);
nand U4512 (N_4512,N_4030,N_3995);
xnor U4513 (N_4513,N_3888,N_4357);
nor U4514 (N_4514,N_3859,N_4171);
or U4515 (N_4515,N_4038,N_4116);
xnor U4516 (N_4516,N_4371,N_3785);
or U4517 (N_4517,N_4318,N_4148);
xor U4518 (N_4518,N_4031,N_4365);
and U4519 (N_4519,N_3856,N_4191);
xnor U4520 (N_4520,N_4275,N_3957);
nor U4521 (N_4521,N_3966,N_4274);
nor U4522 (N_4522,N_3753,N_3775);
nor U4523 (N_4523,N_4187,N_3971);
nor U4524 (N_4524,N_4341,N_4028);
xnor U4525 (N_4525,N_4358,N_4006);
or U4526 (N_4526,N_3778,N_4315);
nand U4527 (N_4527,N_4086,N_3774);
or U4528 (N_4528,N_4075,N_3961);
nor U4529 (N_4529,N_3931,N_3832);
and U4530 (N_4530,N_4224,N_3764);
xnor U4531 (N_4531,N_4132,N_4198);
and U4532 (N_4532,N_4166,N_4062);
nor U4533 (N_4533,N_3759,N_3771);
or U4534 (N_4534,N_3882,N_4128);
and U4535 (N_4535,N_4076,N_4037);
xnor U4536 (N_4536,N_3807,N_3801);
or U4537 (N_4537,N_4133,N_4020);
nor U4538 (N_4538,N_4137,N_3813);
nor U4539 (N_4539,N_3962,N_3852);
and U4540 (N_4540,N_4373,N_4003);
nand U4541 (N_4541,N_4065,N_3873);
nor U4542 (N_4542,N_4244,N_3872);
nand U4543 (N_4543,N_4334,N_3838);
nor U4544 (N_4544,N_3847,N_3880);
nand U4545 (N_4545,N_4051,N_3878);
nor U4546 (N_4546,N_4125,N_4195);
nand U4547 (N_4547,N_4351,N_4010);
or U4548 (N_4548,N_4192,N_4238);
or U4549 (N_4549,N_4330,N_4295);
xor U4550 (N_4550,N_3990,N_4259);
nor U4551 (N_4551,N_3870,N_4223);
and U4552 (N_4552,N_3875,N_3997);
and U4553 (N_4553,N_3943,N_4167);
xor U4554 (N_4554,N_4309,N_4033);
and U4555 (N_4555,N_4273,N_3904);
nor U4556 (N_4556,N_3861,N_4227);
and U4557 (N_4557,N_4327,N_4178);
nand U4558 (N_4558,N_3794,N_3803);
or U4559 (N_4559,N_4319,N_4042);
nand U4560 (N_4560,N_3795,N_3932);
nor U4561 (N_4561,N_3941,N_4308);
xnor U4562 (N_4562,N_4294,N_3802);
xor U4563 (N_4563,N_4032,N_4369);
and U4564 (N_4564,N_4340,N_4107);
nor U4565 (N_4565,N_4211,N_3829);
xnor U4566 (N_4566,N_3831,N_3820);
nor U4567 (N_4567,N_4048,N_3970);
and U4568 (N_4568,N_4134,N_3909);
nor U4569 (N_4569,N_3863,N_4337);
nand U4570 (N_4570,N_3968,N_3946);
nand U4571 (N_4571,N_4177,N_3763);
nand U4572 (N_4572,N_3784,N_3786);
nor U4573 (N_4573,N_4026,N_4299);
xnor U4574 (N_4574,N_4021,N_4139);
nor U4575 (N_4575,N_4069,N_4281);
or U4576 (N_4576,N_3836,N_4152);
xnor U4577 (N_4577,N_3754,N_3826);
nor U4578 (N_4578,N_4044,N_3912);
and U4579 (N_4579,N_3917,N_4253);
nor U4580 (N_4580,N_4202,N_4246);
and U4581 (N_4581,N_3828,N_4135);
or U4582 (N_4582,N_3822,N_4362);
nand U4583 (N_4583,N_3799,N_4118);
xor U4584 (N_4584,N_4025,N_4126);
nor U4585 (N_4585,N_3925,N_4333);
xor U4586 (N_4586,N_3956,N_4374);
xor U4587 (N_4587,N_4284,N_3762);
nand U4588 (N_4588,N_4108,N_3994);
xnor U4589 (N_4589,N_4209,N_4142);
xnor U4590 (N_4590,N_3777,N_4156);
xor U4591 (N_4591,N_4014,N_4231);
nor U4592 (N_4592,N_3827,N_3933);
xor U4593 (N_4593,N_3905,N_4105);
or U4594 (N_4594,N_4040,N_3770);
or U4595 (N_4595,N_4090,N_4332);
and U4596 (N_4596,N_3842,N_4197);
and U4597 (N_4597,N_4190,N_4164);
nor U4598 (N_4598,N_4352,N_4119);
nor U4599 (N_4599,N_3862,N_3833);
or U4600 (N_4600,N_3867,N_4342);
and U4601 (N_4601,N_4234,N_3919);
nand U4602 (N_4602,N_3853,N_4323);
xor U4603 (N_4603,N_4214,N_3864);
nor U4604 (N_4604,N_4078,N_4229);
or U4605 (N_4605,N_3819,N_4235);
nor U4606 (N_4606,N_4140,N_4083);
xnor U4607 (N_4607,N_4250,N_4147);
nor U4608 (N_4608,N_3923,N_3987);
nor U4609 (N_4609,N_3918,N_3766);
nor U4610 (N_4610,N_4059,N_4263);
or U4611 (N_4611,N_3866,N_4194);
and U4612 (N_4612,N_3954,N_4364);
or U4613 (N_4613,N_4045,N_4009);
or U4614 (N_4614,N_4159,N_3959);
or U4615 (N_4615,N_4354,N_4146);
nand U4616 (N_4616,N_4292,N_4060);
xnor U4617 (N_4617,N_4329,N_3984);
nand U4618 (N_4618,N_4004,N_4149);
nand U4619 (N_4619,N_3752,N_4269);
nand U4620 (N_4620,N_3999,N_3814);
nor U4621 (N_4621,N_4180,N_4240);
nor U4622 (N_4622,N_4109,N_3845);
nand U4623 (N_4623,N_4121,N_3791);
nand U4624 (N_4624,N_3758,N_4207);
nand U4625 (N_4625,N_3921,N_4338);
xor U4626 (N_4626,N_4370,N_3929);
xor U4627 (N_4627,N_3772,N_3765);
nor U4628 (N_4628,N_3913,N_3835);
or U4629 (N_4629,N_3935,N_3974);
xor U4630 (N_4630,N_3979,N_3967);
nand U4631 (N_4631,N_4046,N_4157);
xnor U4632 (N_4632,N_3751,N_3767);
and U4633 (N_4633,N_4268,N_4039);
xnor U4634 (N_4634,N_3797,N_3885);
and U4635 (N_4635,N_4203,N_3976);
nor U4636 (N_4636,N_4179,N_3916);
nor U4637 (N_4637,N_4328,N_3892);
and U4638 (N_4638,N_4218,N_4013);
nand U4639 (N_4639,N_4285,N_3889);
nand U4640 (N_4640,N_4239,N_3844);
and U4641 (N_4641,N_4096,N_3843);
or U4642 (N_4642,N_3907,N_4286);
xnor U4643 (N_4643,N_4055,N_3783);
nor U4644 (N_4644,N_3886,N_3781);
xnor U4645 (N_4645,N_4270,N_4160);
or U4646 (N_4646,N_4289,N_4131);
nor U4647 (N_4647,N_4085,N_3871);
xor U4648 (N_4648,N_4320,N_3993);
nand U4649 (N_4649,N_4280,N_4145);
and U4650 (N_4650,N_3980,N_4307);
nor U4651 (N_4651,N_4188,N_4104);
or U4652 (N_4652,N_4169,N_3920);
xnor U4653 (N_4653,N_4158,N_3936);
nand U4654 (N_4654,N_3914,N_3857);
nand U4655 (N_4655,N_4151,N_4015);
nand U4656 (N_4656,N_4304,N_4265);
nand U4657 (N_4657,N_3908,N_3787);
nand U4658 (N_4658,N_4325,N_4277);
or U4659 (N_4659,N_3811,N_4043);
nor U4660 (N_4660,N_3816,N_3846);
xor U4661 (N_4661,N_4050,N_3793);
xor U4662 (N_4662,N_4176,N_4237);
and U4663 (N_4663,N_3789,N_4095);
nor U4664 (N_4664,N_3950,N_3750);
xnor U4665 (N_4665,N_4344,N_3839);
nand U4666 (N_4666,N_4196,N_4101);
xnor U4667 (N_4667,N_3817,N_4008);
and U4668 (N_4668,N_4205,N_4241);
nand U4669 (N_4669,N_4210,N_3887);
and U4670 (N_4670,N_3948,N_4034);
xor U4671 (N_4671,N_4035,N_4230);
xnor U4672 (N_4672,N_4254,N_3938);
and U4673 (N_4673,N_3910,N_4321);
xor U4674 (N_4674,N_4349,N_4311);
or U4675 (N_4675,N_3986,N_4346);
nor U4676 (N_4676,N_3877,N_3951);
nor U4677 (N_4677,N_3782,N_4182);
nand U4678 (N_4678,N_4305,N_3860);
nor U4679 (N_4679,N_4110,N_3981);
and U4680 (N_4680,N_3928,N_3945);
xnor U4681 (N_4681,N_4288,N_4217);
nand U4682 (N_4682,N_3955,N_4300);
and U4683 (N_4683,N_4247,N_4052);
xnor U4684 (N_4684,N_3805,N_3790);
or U4685 (N_4685,N_4174,N_4073);
or U4686 (N_4686,N_3978,N_4063);
nor U4687 (N_4687,N_4221,N_4336);
nor U4688 (N_4688,N_4345,N_3975);
nor U4689 (N_4689,N_4058,N_3938);
and U4690 (N_4690,N_4072,N_4151);
nand U4691 (N_4691,N_3802,N_3876);
or U4692 (N_4692,N_3897,N_4238);
or U4693 (N_4693,N_4088,N_4119);
or U4694 (N_4694,N_4335,N_4332);
nor U4695 (N_4695,N_4305,N_4163);
or U4696 (N_4696,N_4352,N_3967);
and U4697 (N_4697,N_4050,N_4131);
xnor U4698 (N_4698,N_3789,N_3981);
nor U4699 (N_4699,N_3933,N_4154);
and U4700 (N_4700,N_3818,N_3900);
xor U4701 (N_4701,N_4042,N_4203);
or U4702 (N_4702,N_3756,N_4067);
or U4703 (N_4703,N_4239,N_4115);
xnor U4704 (N_4704,N_4320,N_3977);
and U4705 (N_4705,N_4269,N_4097);
nor U4706 (N_4706,N_3773,N_3935);
and U4707 (N_4707,N_4111,N_4075);
nor U4708 (N_4708,N_4313,N_3802);
nand U4709 (N_4709,N_4017,N_4137);
nand U4710 (N_4710,N_3978,N_4000);
or U4711 (N_4711,N_4011,N_4182);
and U4712 (N_4712,N_4197,N_4061);
or U4713 (N_4713,N_4362,N_4076);
nand U4714 (N_4714,N_3975,N_4368);
xnor U4715 (N_4715,N_3754,N_3847);
nor U4716 (N_4716,N_3897,N_3854);
nand U4717 (N_4717,N_4286,N_4356);
and U4718 (N_4718,N_3975,N_4128);
nor U4719 (N_4719,N_4175,N_3794);
and U4720 (N_4720,N_4061,N_3864);
nand U4721 (N_4721,N_4027,N_3970);
nor U4722 (N_4722,N_4122,N_3880);
xnor U4723 (N_4723,N_4173,N_3768);
xnor U4724 (N_4724,N_4351,N_4266);
xnor U4725 (N_4725,N_3942,N_4153);
nor U4726 (N_4726,N_4139,N_3819);
xnor U4727 (N_4727,N_4307,N_3773);
or U4728 (N_4728,N_3943,N_4359);
xnor U4729 (N_4729,N_4125,N_4005);
xor U4730 (N_4730,N_4029,N_3838);
nand U4731 (N_4731,N_3984,N_4339);
xnor U4732 (N_4732,N_4169,N_4298);
nor U4733 (N_4733,N_3880,N_4099);
or U4734 (N_4734,N_4044,N_4206);
or U4735 (N_4735,N_4215,N_3833);
or U4736 (N_4736,N_4302,N_4314);
nand U4737 (N_4737,N_4101,N_4064);
nor U4738 (N_4738,N_4239,N_4026);
or U4739 (N_4739,N_4108,N_4045);
xnor U4740 (N_4740,N_3927,N_3946);
or U4741 (N_4741,N_4240,N_4148);
or U4742 (N_4742,N_3942,N_3810);
or U4743 (N_4743,N_3970,N_3767);
and U4744 (N_4744,N_3792,N_3916);
and U4745 (N_4745,N_3837,N_3921);
and U4746 (N_4746,N_4166,N_3932);
or U4747 (N_4747,N_4141,N_4079);
and U4748 (N_4748,N_3847,N_4018);
and U4749 (N_4749,N_4078,N_4162);
nor U4750 (N_4750,N_4323,N_4218);
or U4751 (N_4751,N_4210,N_4272);
or U4752 (N_4752,N_4203,N_4246);
xnor U4753 (N_4753,N_4217,N_4207);
and U4754 (N_4754,N_4321,N_3843);
and U4755 (N_4755,N_3897,N_4356);
or U4756 (N_4756,N_4235,N_3900);
xor U4757 (N_4757,N_4013,N_4066);
or U4758 (N_4758,N_3869,N_3848);
nor U4759 (N_4759,N_3894,N_4010);
nand U4760 (N_4760,N_4205,N_4272);
nand U4761 (N_4761,N_4044,N_3884);
and U4762 (N_4762,N_4017,N_4262);
or U4763 (N_4763,N_4247,N_3939);
nand U4764 (N_4764,N_4154,N_4165);
nand U4765 (N_4765,N_4340,N_4309);
nor U4766 (N_4766,N_4053,N_4369);
nor U4767 (N_4767,N_4205,N_4260);
and U4768 (N_4768,N_4314,N_4022);
nand U4769 (N_4769,N_4126,N_4159);
xor U4770 (N_4770,N_4214,N_3920);
and U4771 (N_4771,N_4228,N_4102);
nand U4772 (N_4772,N_4060,N_4177);
or U4773 (N_4773,N_3897,N_4302);
nor U4774 (N_4774,N_3919,N_3974);
nor U4775 (N_4775,N_4071,N_3793);
xnor U4776 (N_4776,N_4290,N_3893);
xor U4777 (N_4777,N_3828,N_4120);
or U4778 (N_4778,N_4213,N_4324);
xnor U4779 (N_4779,N_3781,N_4273);
and U4780 (N_4780,N_3801,N_4232);
nand U4781 (N_4781,N_3833,N_4144);
nand U4782 (N_4782,N_4098,N_4292);
or U4783 (N_4783,N_4310,N_3966);
nand U4784 (N_4784,N_3919,N_4067);
nor U4785 (N_4785,N_3804,N_4334);
xor U4786 (N_4786,N_4163,N_4344);
nand U4787 (N_4787,N_4322,N_3868);
or U4788 (N_4788,N_3995,N_3992);
xor U4789 (N_4789,N_4140,N_4323);
or U4790 (N_4790,N_3755,N_3775);
or U4791 (N_4791,N_4134,N_4281);
or U4792 (N_4792,N_4336,N_3982);
nor U4793 (N_4793,N_4224,N_4213);
nand U4794 (N_4794,N_4282,N_3987);
xor U4795 (N_4795,N_3807,N_4366);
nor U4796 (N_4796,N_4327,N_4088);
nand U4797 (N_4797,N_4211,N_3969);
or U4798 (N_4798,N_4303,N_3875);
nor U4799 (N_4799,N_3875,N_3941);
or U4800 (N_4800,N_4311,N_3808);
nand U4801 (N_4801,N_4092,N_3974);
or U4802 (N_4802,N_4044,N_4166);
nor U4803 (N_4803,N_4091,N_4323);
nand U4804 (N_4804,N_3871,N_4064);
nand U4805 (N_4805,N_3925,N_4165);
and U4806 (N_4806,N_4346,N_4137);
or U4807 (N_4807,N_4034,N_3774);
and U4808 (N_4808,N_3996,N_3784);
nand U4809 (N_4809,N_4282,N_3970);
or U4810 (N_4810,N_4173,N_4248);
nand U4811 (N_4811,N_4026,N_4106);
nor U4812 (N_4812,N_4037,N_4372);
nor U4813 (N_4813,N_3994,N_3823);
and U4814 (N_4814,N_3970,N_4155);
xnor U4815 (N_4815,N_3843,N_3924);
xnor U4816 (N_4816,N_4019,N_4329);
and U4817 (N_4817,N_3803,N_4046);
nor U4818 (N_4818,N_3949,N_3768);
nand U4819 (N_4819,N_3966,N_4280);
xnor U4820 (N_4820,N_3970,N_3995);
nand U4821 (N_4821,N_3860,N_4057);
or U4822 (N_4822,N_4358,N_3794);
and U4823 (N_4823,N_4217,N_3906);
nor U4824 (N_4824,N_4336,N_4356);
and U4825 (N_4825,N_4094,N_3948);
or U4826 (N_4826,N_3750,N_4149);
or U4827 (N_4827,N_4201,N_3993);
nor U4828 (N_4828,N_4028,N_4296);
or U4829 (N_4829,N_3899,N_4007);
nand U4830 (N_4830,N_3789,N_3813);
nand U4831 (N_4831,N_3776,N_4304);
nor U4832 (N_4832,N_4330,N_3872);
nand U4833 (N_4833,N_4360,N_4101);
nor U4834 (N_4834,N_4295,N_4138);
or U4835 (N_4835,N_4188,N_4338);
or U4836 (N_4836,N_4032,N_3947);
xor U4837 (N_4837,N_4172,N_3798);
and U4838 (N_4838,N_4046,N_4146);
nand U4839 (N_4839,N_3996,N_4160);
xor U4840 (N_4840,N_4121,N_4163);
or U4841 (N_4841,N_4314,N_4144);
nand U4842 (N_4842,N_4120,N_4109);
nor U4843 (N_4843,N_3899,N_3902);
xnor U4844 (N_4844,N_4344,N_4034);
and U4845 (N_4845,N_4063,N_3764);
nand U4846 (N_4846,N_4042,N_4369);
xor U4847 (N_4847,N_3925,N_4115);
nand U4848 (N_4848,N_4189,N_4171);
or U4849 (N_4849,N_3871,N_4048);
nand U4850 (N_4850,N_4111,N_4249);
and U4851 (N_4851,N_3849,N_4039);
nor U4852 (N_4852,N_3885,N_4050);
nand U4853 (N_4853,N_4086,N_4068);
xnor U4854 (N_4854,N_4081,N_3769);
xor U4855 (N_4855,N_4000,N_4060);
and U4856 (N_4856,N_4340,N_3766);
xnor U4857 (N_4857,N_3939,N_3823);
and U4858 (N_4858,N_4140,N_3873);
nor U4859 (N_4859,N_3942,N_4126);
nand U4860 (N_4860,N_4146,N_4074);
nand U4861 (N_4861,N_4162,N_4100);
and U4862 (N_4862,N_3845,N_4283);
and U4863 (N_4863,N_4010,N_4199);
nand U4864 (N_4864,N_4270,N_4208);
or U4865 (N_4865,N_4095,N_4170);
nor U4866 (N_4866,N_4004,N_3793);
nand U4867 (N_4867,N_3918,N_4370);
or U4868 (N_4868,N_3956,N_4043);
nor U4869 (N_4869,N_4350,N_4002);
nand U4870 (N_4870,N_3804,N_4000);
nor U4871 (N_4871,N_4112,N_4005);
nor U4872 (N_4872,N_4083,N_4038);
or U4873 (N_4873,N_3886,N_3995);
nor U4874 (N_4874,N_4247,N_3783);
and U4875 (N_4875,N_3803,N_4304);
nor U4876 (N_4876,N_4032,N_4135);
or U4877 (N_4877,N_4207,N_3818);
nor U4878 (N_4878,N_4001,N_4113);
xnor U4879 (N_4879,N_3824,N_4178);
or U4880 (N_4880,N_3815,N_4372);
nor U4881 (N_4881,N_3877,N_4310);
or U4882 (N_4882,N_4016,N_4118);
and U4883 (N_4883,N_4196,N_3888);
and U4884 (N_4884,N_4191,N_3816);
xnor U4885 (N_4885,N_4116,N_4267);
or U4886 (N_4886,N_4359,N_4052);
nand U4887 (N_4887,N_4237,N_3993);
and U4888 (N_4888,N_4308,N_4014);
nor U4889 (N_4889,N_3961,N_4301);
and U4890 (N_4890,N_3759,N_4088);
nor U4891 (N_4891,N_4018,N_4322);
or U4892 (N_4892,N_3815,N_3985);
nand U4893 (N_4893,N_3834,N_4321);
nor U4894 (N_4894,N_4235,N_3800);
and U4895 (N_4895,N_4348,N_3843);
and U4896 (N_4896,N_4065,N_4322);
xnor U4897 (N_4897,N_4152,N_4021);
or U4898 (N_4898,N_3890,N_3902);
nor U4899 (N_4899,N_4284,N_4371);
and U4900 (N_4900,N_3751,N_3761);
or U4901 (N_4901,N_4214,N_4271);
xnor U4902 (N_4902,N_4254,N_3899);
and U4903 (N_4903,N_4368,N_4215);
and U4904 (N_4904,N_4120,N_3861);
and U4905 (N_4905,N_4153,N_3770);
xnor U4906 (N_4906,N_4061,N_3922);
nor U4907 (N_4907,N_4047,N_4342);
xnor U4908 (N_4908,N_3975,N_4064);
nand U4909 (N_4909,N_4295,N_4228);
nor U4910 (N_4910,N_3981,N_4041);
and U4911 (N_4911,N_4230,N_3889);
or U4912 (N_4912,N_4196,N_3883);
nor U4913 (N_4913,N_3760,N_4224);
nand U4914 (N_4914,N_3958,N_3961);
xnor U4915 (N_4915,N_4052,N_4257);
nand U4916 (N_4916,N_4002,N_4153);
or U4917 (N_4917,N_4174,N_3909);
and U4918 (N_4918,N_4124,N_3804);
or U4919 (N_4919,N_3915,N_3769);
nor U4920 (N_4920,N_3960,N_4030);
or U4921 (N_4921,N_3844,N_4161);
and U4922 (N_4922,N_4326,N_3864);
xor U4923 (N_4923,N_4193,N_4273);
and U4924 (N_4924,N_4082,N_3930);
xor U4925 (N_4925,N_4314,N_4015);
nor U4926 (N_4926,N_4148,N_4041);
or U4927 (N_4927,N_4165,N_4195);
or U4928 (N_4928,N_4090,N_4306);
nor U4929 (N_4929,N_3917,N_4327);
nor U4930 (N_4930,N_4309,N_3909);
xor U4931 (N_4931,N_4054,N_4005);
and U4932 (N_4932,N_4334,N_4275);
xor U4933 (N_4933,N_4061,N_4350);
nor U4934 (N_4934,N_4089,N_4031);
nor U4935 (N_4935,N_4198,N_3763);
and U4936 (N_4936,N_4233,N_4364);
xnor U4937 (N_4937,N_4253,N_4304);
nand U4938 (N_4938,N_4021,N_4251);
nor U4939 (N_4939,N_3915,N_4206);
or U4940 (N_4940,N_3881,N_4361);
and U4941 (N_4941,N_3896,N_3992);
and U4942 (N_4942,N_4043,N_3806);
nor U4943 (N_4943,N_4106,N_3801);
nand U4944 (N_4944,N_4309,N_4161);
and U4945 (N_4945,N_4372,N_3789);
or U4946 (N_4946,N_3818,N_3851);
nor U4947 (N_4947,N_4356,N_4148);
nor U4948 (N_4948,N_4171,N_3778);
or U4949 (N_4949,N_4303,N_4027);
nor U4950 (N_4950,N_3973,N_3804);
or U4951 (N_4951,N_4111,N_3865);
nand U4952 (N_4952,N_4312,N_3925);
nand U4953 (N_4953,N_4165,N_3852);
nand U4954 (N_4954,N_4161,N_4349);
nand U4955 (N_4955,N_4029,N_3879);
nand U4956 (N_4956,N_4109,N_4267);
and U4957 (N_4957,N_4078,N_4011);
nor U4958 (N_4958,N_4348,N_4337);
and U4959 (N_4959,N_3797,N_4356);
or U4960 (N_4960,N_4328,N_3837);
nand U4961 (N_4961,N_3864,N_4037);
xor U4962 (N_4962,N_4368,N_4352);
nand U4963 (N_4963,N_4035,N_3767);
and U4964 (N_4964,N_4001,N_4099);
nor U4965 (N_4965,N_3839,N_3924);
or U4966 (N_4966,N_4218,N_4110);
xnor U4967 (N_4967,N_4053,N_3776);
nand U4968 (N_4968,N_4370,N_3836);
or U4969 (N_4969,N_4348,N_3794);
or U4970 (N_4970,N_4040,N_4133);
nor U4971 (N_4971,N_3792,N_4298);
or U4972 (N_4972,N_3919,N_3863);
xor U4973 (N_4973,N_3903,N_3993);
or U4974 (N_4974,N_3856,N_4297);
nor U4975 (N_4975,N_3760,N_3770);
or U4976 (N_4976,N_4370,N_4165);
xnor U4977 (N_4977,N_4018,N_4012);
nand U4978 (N_4978,N_4161,N_3762);
and U4979 (N_4979,N_4110,N_4152);
nor U4980 (N_4980,N_4128,N_4215);
nand U4981 (N_4981,N_4361,N_4186);
or U4982 (N_4982,N_4241,N_4347);
xor U4983 (N_4983,N_4315,N_3791);
nor U4984 (N_4984,N_3909,N_4290);
nand U4985 (N_4985,N_4296,N_4128);
nor U4986 (N_4986,N_3759,N_3855);
nor U4987 (N_4987,N_3985,N_3876);
or U4988 (N_4988,N_3928,N_3871);
or U4989 (N_4989,N_3859,N_3956);
and U4990 (N_4990,N_4221,N_4363);
or U4991 (N_4991,N_4318,N_4032);
xor U4992 (N_4992,N_4285,N_4366);
nand U4993 (N_4993,N_3943,N_4173);
and U4994 (N_4994,N_4226,N_4028);
xnor U4995 (N_4995,N_4286,N_3824);
nor U4996 (N_4996,N_4086,N_3788);
nand U4997 (N_4997,N_4118,N_4292);
xor U4998 (N_4998,N_4075,N_3804);
nor U4999 (N_4999,N_4072,N_3756);
and U5000 (N_5000,N_4528,N_4861);
and U5001 (N_5001,N_4904,N_4740);
or U5002 (N_5002,N_4847,N_4809);
xnor U5003 (N_5003,N_4788,N_4666);
xnor U5004 (N_5004,N_4718,N_4520);
nand U5005 (N_5005,N_4697,N_4783);
xor U5006 (N_5006,N_4540,N_4558);
or U5007 (N_5007,N_4844,N_4796);
and U5008 (N_5008,N_4525,N_4482);
and U5009 (N_5009,N_4590,N_4874);
nand U5010 (N_5010,N_4687,N_4506);
xnor U5011 (N_5011,N_4815,N_4647);
nand U5012 (N_5012,N_4918,N_4742);
nand U5013 (N_5013,N_4767,N_4645);
xor U5014 (N_5014,N_4870,N_4532);
nor U5015 (N_5015,N_4680,N_4786);
or U5016 (N_5016,N_4485,N_4571);
nand U5017 (N_5017,N_4871,N_4704);
and U5018 (N_5018,N_4942,N_4863);
and U5019 (N_5019,N_4509,N_4657);
and U5020 (N_5020,N_4737,N_4500);
xor U5021 (N_5021,N_4919,N_4624);
nand U5022 (N_5022,N_4480,N_4574);
nor U5023 (N_5023,N_4854,N_4884);
nor U5024 (N_5024,N_4614,N_4518);
or U5025 (N_5025,N_4759,N_4576);
xor U5026 (N_5026,N_4495,N_4486);
nand U5027 (N_5027,N_4419,N_4489);
nand U5028 (N_5028,N_4632,N_4862);
and U5029 (N_5029,N_4834,N_4734);
nand U5030 (N_5030,N_4689,N_4722);
or U5031 (N_5031,N_4956,N_4967);
nor U5032 (N_5032,N_4693,N_4582);
nor U5033 (N_5033,N_4968,N_4387);
xnor U5034 (N_5034,N_4925,N_4597);
xnor U5035 (N_5035,N_4784,N_4463);
and U5036 (N_5036,N_4947,N_4619);
xnor U5037 (N_5037,N_4917,N_4801);
nand U5038 (N_5038,N_4700,N_4515);
and U5039 (N_5039,N_4642,N_4991);
nor U5040 (N_5040,N_4941,N_4720);
nor U5041 (N_5041,N_4466,N_4455);
xor U5042 (N_5042,N_4604,N_4444);
nor U5043 (N_5043,N_4996,N_4936);
or U5044 (N_5044,N_4866,N_4762);
nor U5045 (N_5045,N_4944,N_4885);
xor U5046 (N_5046,N_4504,N_4908);
and U5047 (N_5047,N_4430,N_4860);
xor U5048 (N_5048,N_4474,N_4600);
or U5049 (N_5049,N_4556,N_4608);
and U5050 (N_5050,N_4686,N_4530);
xor U5051 (N_5051,N_4450,N_4843);
xor U5052 (N_5052,N_4462,N_4554);
nor U5053 (N_5053,N_4502,N_4826);
nand U5054 (N_5054,N_4476,N_4977);
nor U5055 (N_5055,N_4706,N_4806);
nor U5056 (N_5056,N_4779,N_4541);
nand U5057 (N_5057,N_4688,N_4379);
nand U5058 (N_5058,N_4713,N_4460);
or U5059 (N_5059,N_4494,N_4751);
or U5060 (N_5060,N_4730,N_4529);
or U5061 (N_5061,N_4453,N_4551);
and U5062 (N_5062,N_4868,N_4431);
or U5063 (N_5063,N_4427,N_4385);
xnor U5064 (N_5064,N_4432,N_4452);
xor U5065 (N_5065,N_4878,N_4789);
xor U5066 (N_5066,N_4629,N_4490);
nor U5067 (N_5067,N_4933,N_4837);
xnor U5068 (N_5068,N_4418,N_4675);
nor U5069 (N_5069,N_4621,N_4875);
nand U5070 (N_5070,N_4993,N_4669);
xor U5071 (N_5071,N_4560,N_4577);
or U5072 (N_5072,N_4548,N_4840);
nand U5073 (N_5073,N_4916,N_4988);
nand U5074 (N_5074,N_4969,N_4910);
nand U5075 (N_5075,N_4683,N_4581);
nor U5076 (N_5076,N_4955,N_4957);
nor U5077 (N_5077,N_4733,N_4421);
nand U5078 (N_5078,N_4798,N_4924);
xnor U5079 (N_5079,N_4754,N_4596);
or U5080 (N_5080,N_4772,N_4999);
xor U5081 (N_5081,N_4838,N_4636);
and U5082 (N_5082,N_4867,N_4563);
nor U5083 (N_5083,N_4649,N_4685);
and U5084 (N_5084,N_4951,N_4975);
or U5085 (N_5085,N_4670,N_4488);
and U5086 (N_5086,N_4865,N_4543);
and U5087 (N_5087,N_4828,N_4731);
nand U5088 (N_5088,N_4561,N_4943);
or U5089 (N_5089,N_4952,N_4795);
and U5090 (N_5090,N_4710,N_4678);
nor U5091 (N_5091,N_4792,N_4816);
nand U5092 (N_5092,N_4507,N_4451);
nand U5093 (N_5093,N_4721,N_4709);
and U5094 (N_5094,N_4546,N_4959);
nor U5095 (N_5095,N_4876,N_4872);
xnor U5096 (N_5096,N_4493,N_4881);
or U5097 (N_5097,N_4818,N_4598);
and U5098 (N_5098,N_4660,N_4521);
nand U5099 (N_5099,N_4569,N_4705);
and U5100 (N_5100,N_4443,N_4814);
and U5101 (N_5101,N_4533,N_4800);
nand U5102 (N_5102,N_4416,N_4616);
and U5103 (N_5103,N_4426,N_4817);
nand U5104 (N_5104,N_4390,N_4777);
nor U5105 (N_5105,N_4813,N_4963);
xor U5106 (N_5106,N_4997,N_4778);
nand U5107 (N_5107,N_4932,N_4973);
xnor U5108 (N_5108,N_4668,N_4449);
or U5109 (N_5109,N_4447,N_4469);
nor U5110 (N_5110,N_4484,N_4573);
or U5111 (N_5111,N_4892,N_4694);
nand U5112 (N_5112,N_4656,N_4934);
nor U5113 (N_5113,N_4436,N_4827);
xor U5114 (N_5114,N_4637,N_4384);
and U5115 (N_5115,N_4939,N_4483);
nor U5116 (N_5116,N_4644,N_4728);
nor U5117 (N_5117,N_4425,N_4617);
and U5118 (N_5118,N_4412,N_4654);
xor U5119 (N_5119,N_4622,N_4897);
or U5120 (N_5120,N_4812,N_4930);
xnor U5121 (N_5121,N_4380,N_4699);
and U5122 (N_5122,N_4567,N_4458);
nand U5123 (N_5123,N_4921,N_4773);
nand U5124 (N_5124,N_4557,N_4756);
nor U5125 (N_5125,N_4625,N_4471);
nor U5126 (N_5126,N_4593,N_4682);
or U5127 (N_5127,N_4413,N_4791);
and U5128 (N_5128,N_4743,N_4607);
xnor U5129 (N_5129,N_4998,N_4691);
nand U5130 (N_5130,N_4994,N_4849);
and U5131 (N_5131,N_4513,N_4962);
and U5132 (N_5132,N_4664,N_4376);
and U5133 (N_5133,N_4510,N_4852);
and U5134 (N_5134,N_4765,N_4626);
nand U5135 (N_5135,N_4981,N_4831);
xor U5136 (N_5136,N_4652,N_4428);
nand U5137 (N_5137,N_4901,N_4785);
or U5138 (N_5138,N_4825,N_4768);
xnor U5139 (N_5139,N_4498,N_4946);
nand U5140 (N_5140,N_4445,N_4522);
or U5141 (N_5141,N_4880,N_4989);
nor U5142 (N_5142,N_4508,N_4900);
or U5143 (N_5143,N_4717,N_4491);
and U5144 (N_5144,N_4468,N_4725);
nor U5145 (N_5145,N_4404,N_4744);
nor U5146 (N_5146,N_4544,N_4984);
nand U5147 (N_5147,N_4399,N_4940);
or U5148 (N_5148,N_4650,N_4797);
and U5149 (N_5149,N_4553,N_4605);
and U5150 (N_5150,N_4928,N_4787);
and U5151 (N_5151,N_4757,N_4736);
and U5152 (N_5152,N_4873,N_4886);
xor U5153 (N_5153,N_4894,N_4763);
and U5154 (N_5154,N_4877,N_4732);
nand U5155 (N_5155,N_4512,N_4524);
nand U5156 (N_5156,N_4758,N_4905);
nor U5157 (N_5157,N_4475,N_4630);
and U5158 (N_5158,N_4702,N_4538);
nor U5159 (N_5159,N_4382,N_4594);
nor U5160 (N_5160,N_4437,N_4855);
nor U5161 (N_5161,N_4599,N_4401);
nand U5162 (N_5162,N_4411,N_4377);
and U5163 (N_5163,N_4954,N_4781);
xnor U5164 (N_5164,N_4770,N_4523);
or U5165 (N_5165,N_4679,N_4433);
and U5166 (N_5166,N_4403,N_4375);
xor U5167 (N_5167,N_4400,N_4889);
nor U5168 (N_5168,N_4627,N_4857);
and U5169 (N_5169,N_4931,N_4729);
nand U5170 (N_5170,N_4440,N_4646);
or U5171 (N_5171,N_4394,N_4464);
nand U5172 (N_5172,N_4961,N_4909);
or U5173 (N_5173,N_4842,N_4811);
nand U5174 (N_5174,N_4526,N_4535);
xnor U5175 (N_5175,N_4550,N_4850);
nand U5176 (N_5176,N_4673,N_4396);
xor U5177 (N_5177,N_4995,N_4695);
nor U5178 (N_5178,N_4985,N_4477);
nand U5179 (N_5179,N_4913,N_4676);
nand U5180 (N_5180,N_4496,N_4653);
xor U5181 (N_5181,N_4612,N_4803);
nand U5182 (N_5182,N_4566,N_4677);
nand U5183 (N_5183,N_4964,N_4423);
and U5184 (N_5184,N_4534,N_4711);
xor U5185 (N_5185,N_4979,N_4926);
or U5186 (N_5186,N_4807,N_4716);
and U5187 (N_5187,N_4591,N_4748);
or U5188 (N_5188,N_4992,N_4568);
nand U5189 (N_5189,N_4858,N_4820);
nand U5190 (N_5190,N_4393,N_4414);
and U5191 (N_5191,N_4948,N_4782);
or U5192 (N_5192,N_4639,N_4672);
or U5193 (N_5193,N_4378,N_4578);
xnor U5194 (N_5194,N_4580,N_4665);
nand U5195 (N_5195,N_4879,N_4461);
xor U5196 (N_5196,N_4392,N_4958);
nor U5197 (N_5197,N_4438,N_4835);
xor U5198 (N_5198,N_4606,N_4853);
xor U5199 (N_5199,N_4681,N_4775);
xnor U5200 (N_5200,N_4615,N_4986);
nand U5201 (N_5201,N_4896,N_4555);
or U5202 (N_5202,N_4603,N_4648);
xnor U5203 (N_5203,N_4741,N_4822);
or U5204 (N_5204,N_4406,N_4635);
or U5205 (N_5205,N_4552,N_4397);
or U5206 (N_5206,N_4755,N_4793);
or U5207 (N_5207,N_4658,N_4856);
xnor U5208 (N_5208,N_4620,N_4714);
and U5209 (N_5209,N_4457,N_4684);
nor U5210 (N_5210,N_4703,N_4902);
nand U5211 (N_5211,N_4836,N_4407);
nor U5212 (N_5212,N_4439,N_4769);
xor U5213 (N_5213,N_4888,N_4945);
nand U5214 (N_5214,N_4472,N_4634);
or U5215 (N_5215,N_4383,N_4389);
and U5216 (N_5216,N_4715,N_4895);
or U5217 (N_5217,N_4848,N_4887);
and U5218 (N_5218,N_4893,N_4570);
and U5219 (N_5219,N_4912,N_4422);
nor U5220 (N_5220,N_4559,N_4983);
or U5221 (N_5221,N_4592,N_4408);
nand U5222 (N_5222,N_4929,N_4511);
nor U5223 (N_5223,N_4752,N_4938);
nor U5224 (N_5224,N_4499,N_4572);
nor U5225 (N_5225,N_4771,N_4766);
nor U5226 (N_5226,N_4588,N_4503);
nand U5227 (N_5227,N_4388,N_4584);
nor U5228 (N_5228,N_4819,N_4846);
nor U5229 (N_5229,N_4671,N_4517);
xor U5230 (N_5230,N_4794,N_4545);
and U5231 (N_5231,N_4613,N_4920);
xor U5232 (N_5232,N_4833,N_4410);
and U5233 (N_5233,N_4381,N_4845);
or U5234 (N_5234,N_4586,N_4448);
and U5235 (N_5235,N_4898,N_4514);
nand U5236 (N_5236,N_4937,N_4505);
nor U5237 (N_5237,N_4478,N_4631);
xor U5238 (N_5238,N_4601,N_4602);
xnor U5239 (N_5239,N_4760,N_4883);
and U5240 (N_5240,N_4395,N_4640);
or U5241 (N_5241,N_4808,N_4698);
nand U5242 (N_5242,N_4802,N_4971);
xnor U5243 (N_5243,N_4927,N_4585);
nand U5244 (N_5244,N_4864,N_4970);
and U5245 (N_5245,N_4906,N_4537);
nor U5246 (N_5246,N_4978,N_4667);
nand U5247 (N_5247,N_4659,N_4527);
nor U5248 (N_5248,N_4859,N_4386);
xnor U5249 (N_5249,N_4456,N_4497);
and U5250 (N_5250,N_4911,N_4739);
nand U5251 (N_5251,N_4719,N_4974);
and U5252 (N_5252,N_4830,N_4804);
xor U5253 (N_5253,N_4549,N_4899);
xor U5254 (N_5254,N_4949,N_4610);
xor U5255 (N_5255,N_4547,N_4424);
and U5256 (N_5256,N_4405,N_4735);
xor U5257 (N_5257,N_4519,N_4536);
and U5258 (N_5258,N_4470,N_4750);
nor U5259 (N_5259,N_4935,N_4562);
nor U5260 (N_5260,N_4391,N_4575);
nand U5261 (N_5261,N_4583,N_4446);
and U5262 (N_5262,N_4662,N_4434);
and U5263 (N_5263,N_4539,N_4907);
or U5264 (N_5264,N_4780,N_4531);
or U5265 (N_5265,N_4790,N_4420);
nand U5266 (N_5266,N_4655,N_4821);
nand U5267 (N_5267,N_4841,N_4479);
or U5268 (N_5268,N_4589,N_4618);
nor U5269 (N_5269,N_4824,N_4441);
nand U5270 (N_5270,N_4542,N_4987);
nand U5271 (N_5271,N_4891,N_4473);
or U5272 (N_5272,N_4409,N_4922);
nor U5273 (N_5273,N_4501,N_4707);
nor U5274 (N_5274,N_4950,N_4839);
or U5275 (N_5275,N_4774,N_4823);
or U5276 (N_5276,N_4587,N_4454);
nor U5277 (N_5277,N_4829,N_4435);
and U5278 (N_5278,N_4799,N_4903);
and U5279 (N_5279,N_4579,N_4564);
xor U5280 (N_5280,N_4923,N_4980);
nor U5281 (N_5281,N_4805,N_4776);
nand U5282 (N_5282,N_4402,N_4661);
nor U5283 (N_5283,N_4745,N_4914);
nor U5284 (N_5284,N_4565,N_4976);
nor U5285 (N_5285,N_4727,N_4724);
or U5286 (N_5286,N_4915,N_4633);
nor U5287 (N_5287,N_4674,N_4415);
or U5288 (N_5288,N_4726,N_4663);
xnor U5289 (N_5289,N_4723,N_4609);
or U5290 (N_5290,N_4429,N_4465);
and U5291 (N_5291,N_4753,N_4712);
xnor U5292 (N_5292,N_4869,N_4708);
nand U5293 (N_5293,N_4761,N_4467);
xnor U5294 (N_5294,N_4417,N_4966);
xnor U5295 (N_5295,N_4442,N_4692);
xnor U5296 (N_5296,N_4481,N_4810);
or U5297 (N_5297,N_4651,N_4890);
and U5298 (N_5298,N_4965,N_4492);
nor U5299 (N_5299,N_4595,N_4960);
nor U5300 (N_5300,N_4487,N_4690);
nand U5301 (N_5301,N_4749,N_4643);
or U5302 (N_5302,N_4747,N_4516);
or U5303 (N_5303,N_4982,N_4611);
nor U5304 (N_5304,N_4851,N_4990);
and U5305 (N_5305,N_4696,N_4638);
or U5306 (N_5306,N_4972,N_4764);
xor U5307 (N_5307,N_4738,N_4628);
nor U5308 (N_5308,N_4398,N_4701);
and U5309 (N_5309,N_4953,N_4641);
nand U5310 (N_5310,N_4623,N_4882);
xnor U5311 (N_5311,N_4459,N_4832);
or U5312 (N_5312,N_4746,N_4876);
nand U5313 (N_5313,N_4645,N_4751);
nand U5314 (N_5314,N_4744,N_4868);
nor U5315 (N_5315,N_4936,N_4521);
or U5316 (N_5316,N_4681,N_4745);
nand U5317 (N_5317,N_4422,N_4729);
or U5318 (N_5318,N_4758,N_4836);
and U5319 (N_5319,N_4382,N_4757);
and U5320 (N_5320,N_4588,N_4863);
nor U5321 (N_5321,N_4628,N_4758);
nor U5322 (N_5322,N_4901,N_4508);
xnor U5323 (N_5323,N_4974,N_4546);
xor U5324 (N_5324,N_4614,N_4841);
or U5325 (N_5325,N_4510,N_4868);
nor U5326 (N_5326,N_4375,N_4720);
nor U5327 (N_5327,N_4791,N_4997);
or U5328 (N_5328,N_4495,N_4540);
and U5329 (N_5329,N_4715,N_4552);
xnor U5330 (N_5330,N_4631,N_4500);
nor U5331 (N_5331,N_4543,N_4399);
xnor U5332 (N_5332,N_4685,N_4489);
or U5333 (N_5333,N_4527,N_4417);
or U5334 (N_5334,N_4411,N_4712);
and U5335 (N_5335,N_4896,N_4741);
nand U5336 (N_5336,N_4426,N_4901);
nor U5337 (N_5337,N_4464,N_4750);
and U5338 (N_5338,N_4591,N_4883);
or U5339 (N_5339,N_4833,N_4620);
or U5340 (N_5340,N_4941,N_4441);
and U5341 (N_5341,N_4401,N_4667);
and U5342 (N_5342,N_4481,N_4799);
xor U5343 (N_5343,N_4873,N_4386);
nand U5344 (N_5344,N_4679,N_4576);
nand U5345 (N_5345,N_4834,N_4581);
and U5346 (N_5346,N_4759,N_4991);
nand U5347 (N_5347,N_4422,N_4828);
and U5348 (N_5348,N_4973,N_4945);
nor U5349 (N_5349,N_4898,N_4993);
nor U5350 (N_5350,N_4539,N_4684);
or U5351 (N_5351,N_4830,N_4821);
or U5352 (N_5352,N_4977,N_4414);
nand U5353 (N_5353,N_4678,N_4843);
or U5354 (N_5354,N_4484,N_4515);
nor U5355 (N_5355,N_4730,N_4457);
and U5356 (N_5356,N_4695,N_4395);
xnor U5357 (N_5357,N_4389,N_4808);
or U5358 (N_5358,N_4834,N_4511);
nand U5359 (N_5359,N_4981,N_4885);
xor U5360 (N_5360,N_4801,N_4799);
and U5361 (N_5361,N_4577,N_4864);
or U5362 (N_5362,N_4789,N_4936);
and U5363 (N_5363,N_4418,N_4683);
and U5364 (N_5364,N_4482,N_4743);
xor U5365 (N_5365,N_4925,N_4827);
xor U5366 (N_5366,N_4525,N_4953);
nand U5367 (N_5367,N_4601,N_4869);
xor U5368 (N_5368,N_4472,N_4618);
xor U5369 (N_5369,N_4907,N_4510);
nor U5370 (N_5370,N_4877,N_4397);
nand U5371 (N_5371,N_4894,N_4642);
nand U5372 (N_5372,N_4923,N_4822);
or U5373 (N_5373,N_4505,N_4949);
or U5374 (N_5374,N_4403,N_4558);
or U5375 (N_5375,N_4711,N_4802);
and U5376 (N_5376,N_4659,N_4605);
and U5377 (N_5377,N_4474,N_4640);
or U5378 (N_5378,N_4419,N_4469);
nand U5379 (N_5379,N_4816,N_4625);
nor U5380 (N_5380,N_4886,N_4755);
xnor U5381 (N_5381,N_4654,N_4682);
xnor U5382 (N_5382,N_4429,N_4809);
xor U5383 (N_5383,N_4425,N_4796);
or U5384 (N_5384,N_4446,N_4475);
xnor U5385 (N_5385,N_4939,N_4800);
nor U5386 (N_5386,N_4408,N_4787);
nor U5387 (N_5387,N_4617,N_4983);
or U5388 (N_5388,N_4604,N_4723);
nand U5389 (N_5389,N_4947,N_4437);
nor U5390 (N_5390,N_4586,N_4700);
nand U5391 (N_5391,N_4659,N_4884);
and U5392 (N_5392,N_4653,N_4838);
xnor U5393 (N_5393,N_4447,N_4970);
nand U5394 (N_5394,N_4943,N_4745);
nor U5395 (N_5395,N_4667,N_4472);
nand U5396 (N_5396,N_4719,N_4376);
xnor U5397 (N_5397,N_4861,N_4732);
and U5398 (N_5398,N_4743,N_4957);
or U5399 (N_5399,N_4480,N_4411);
nor U5400 (N_5400,N_4768,N_4766);
or U5401 (N_5401,N_4648,N_4889);
nand U5402 (N_5402,N_4679,N_4465);
xnor U5403 (N_5403,N_4585,N_4436);
and U5404 (N_5404,N_4686,N_4553);
xnor U5405 (N_5405,N_4582,N_4459);
nand U5406 (N_5406,N_4966,N_4920);
nor U5407 (N_5407,N_4829,N_4770);
and U5408 (N_5408,N_4821,N_4532);
and U5409 (N_5409,N_4727,N_4478);
or U5410 (N_5410,N_4451,N_4479);
or U5411 (N_5411,N_4750,N_4706);
xnor U5412 (N_5412,N_4403,N_4771);
or U5413 (N_5413,N_4808,N_4703);
nor U5414 (N_5414,N_4459,N_4518);
and U5415 (N_5415,N_4404,N_4768);
nand U5416 (N_5416,N_4728,N_4777);
nand U5417 (N_5417,N_4441,N_4485);
nor U5418 (N_5418,N_4640,N_4931);
and U5419 (N_5419,N_4581,N_4753);
nand U5420 (N_5420,N_4454,N_4964);
and U5421 (N_5421,N_4422,N_4676);
or U5422 (N_5422,N_4471,N_4944);
nor U5423 (N_5423,N_4554,N_4873);
and U5424 (N_5424,N_4678,N_4854);
nand U5425 (N_5425,N_4604,N_4424);
xnor U5426 (N_5426,N_4608,N_4776);
and U5427 (N_5427,N_4457,N_4541);
xor U5428 (N_5428,N_4597,N_4734);
nand U5429 (N_5429,N_4517,N_4872);
nor U5430 (N_5430,N_4593,N_4783);
nand U5431 (N_5431,N_4787,N_4756);
and U5432 (N_5432,N_4891,N_4408);
xor U5433 (N_5433,N_4418,N_4760);
and U5434 (N_5434,N_4733,N_4838);
or U5435 (N_5435,N_4440,N_4504);
nand U5436 (N_5436,N_4541,N_4787);
nor U5437 (N_5437,N_4933,N_4798);
nand U5438 (N_5438,N_4939,N_4725);
nand U5439 (N_5439,N_4530,N_4998);
nand U5440 (N_5440,N_4471,N_4483);
nand U5441 (N_5441,N_4429,N_4413);
nor U5442 (N_5442,N_4662,N_4964);
xnor U5443 (N_5443,N_4973,N_4991);
and U5444 (N_5444,N_4966,N_4661);
xnor U5445 (N_5445,N_4470,N_4422);
nor U5446 (N_5446,N_4714,N_4428);
xnor U5447 (N_5447,N_4886,N_4390);
nand U5448 (N_5448,N_4689,N_4618);
or U5449 (N_5449,N_4635,N_4971);
and U5450 (N_5450,N_4513,N_4709);
xnor U5451 (N_5451,N_4726,N_4910);
nand U5452 (N_5452,N_4841,N_4544);
xnor U5453 (N_5453,N_4669,N_4770);
xor U5454 (N_5454,N_4477,N_4855);
nand U5455 (N_5455,N_4777,N_4386);
or U5456 (N_5456,N_4920,N_4715);
or U5457 (N_5457,N_4414,N_4906);
and U5458 (N_5458,N_4885,N_4800);
or U5459 (N_5459,N_4478,N_4719);
or U5460 (N_5460,N_4391,N_4538);
and U5461 (N_5461,N_4794,N_4632);
xor U5462 (N_5462,N_4738,N_4841);
nor U5463 (N_5463,N_4941,N_4753);
xor U5464 (N_5464,N_4674,N_4823);
and U5465 (N_5465,N_4769,N_4683);
nor U5466 (N_5466,N_4981,N_4555);
and U5467 (N_5467,N_4446,N_4991);
and U5468 (N_5468,N_4931,N_4539);
xor U5469 (N_5469,N_4409,N_4564);
nor U5470 (N_5470,N_4685,N_4641);
or U5471 (N_5471,N_4473,N_4869);
and U5472 (N_5472,N_4503,N_4858);
and U5473 (N_5473,N_4553,N_4574);
and U5474 (N_5474,N_4964,N_4479);
xor U5475 (N_5475,N_4401,N_4425);
nor U5476 (N_5476,N_4811,N_4498);
xnor U5477 (N_5477,N_4610,N_4914);
or U5478 (N_5478,N_4684,N_4710);
xnor U5479 (N_5479,N_4460,N_4998);
or U5480 (N_5480,N_4640,N_4690);
xor U5481 (N_5481,N_4737,N_4556);
nor U5482 (N_5482,N_4610,N_4390);
xor U5483 (N_5483,N_4597,N_4423);
nand U5484 (N_5484,N_4585,N_4887);
nand U5485 (N_5485,N_4630,N_4896);
nand U5486 (N_5486,N_4940,N_4500);
or U5487 (N_5487,N_4418,N_4385);
or U5488 (N_5488,N_4925,N_4784);
or U5489 (N_5489,N_4773,N_4982);
nor U5490 (N_5490,N_4535,N_4627);
or U5491 (N_5491,N_4837,N_4677);
or U5492 (N_5492,N_4754,N_4881);
and U5493 (N_5493,N_4645,N_4817);
nand U5494 (N_5494,N_4834,N_4382);
and U5495 (N_5495,N_4821,N_4584);
nand U5496 (N_5496,N_4842,N_4570);
nor U5497 (N_5497,N_4391,N_4994);
nand U5498 (N_5498,N_4460,N_4789);
and U5499 (N_5499,N_4422,N_4464);
nand U5500 (N_5500,N_4873,N_4834);
nor U5501 (N_5501,N_4859,N_4824);
or U5502 (N_5502,N_4387,N_4636);
or U5503 (N_5503,N_4960,N_4716);
and U5504 (N_5504,N_4742,N_4659);
nand U5505 (N_5505,N_4574,N_4450);
and U5506 (N_5506,N_4660,N_4801);
xor U5507 (N_5507,N_4998,N_4442);
nor U5508 (N_5508,N_4578,N_4564);
xnor U5509 (N_5509,N_4504,N_4816);
nand U5510 (N_5510,N_4643,N_4658);
and U5511 (N_5511,N_4487,N_4443);
nand U5512 (N_5512,N_4586,N_4735);
xor U5513 (N_5513,N_4721,N_4609);
and U5514 (N_5514,N_4805,N_4511);
xor U5515 (N_5515,N_4557,N_4776);
or U5516 (N_5516,N_4388,N_4501);
nor U5517 (N_5517,N_4650,N_4997);
xnor U5518 (N_5518,N_4976,N_4715);
nand U5519 (N_5519,N_4906,N_4709);
and U5520 (N_5520,N_4633,N_4645);
xor U5521 (N_5521,N_4850,N_4591);
or U5522 (N_5522,N_4645,N_4574);
nor U5523 (N_5523,N_4853,N_4866);
xnor U5524 (N_5524,N_4677,N_4725);
or U5525 (N_5525,N_4465,N_4415);
nor U5526 (N_5526,N_4464,N_4822);
and U5527 (N_5527,N_4398,N_4784);
and U5528 (N_5528,N_4430,N_4450);
xor U5529 (N_5529,N_4655,N_4950);
xor U5530 (N_5530,N_4589,N_4911);
and U5531 (N_5531,N_4473,N_4457);
and U5532 (N_5532,N_4487,N_4376);
nand U5533 (N_5533,N_4798,N_4767);
and U5534 (N_5534,N_4759,N_4912);
or U5535 (N_5535,N_4656,N_4663);
nand U5536 (N_5536,N_4772,N_4878);
nand U5537 (N_5537,N_4941,N_4521);
nor U5538 (N_5538,N_4584,N_4983);
and U5539 (N_5539,N_4544,N_4643);
or U5540 (N_5540,N_4979,N_4981);
and U5541 (N_5541,N_4659,N_4610);
and U5542 (N_5542,N_4929,N_4489);
nand U5543 (N_5543,N_4495,N_4874);
xnor U5544 (N_5544,N_4820,N_4757);
and U5545 (N_5545,N_4936,N_4603);
or U5546 (N_5546,N_4541,N_4538);
nor U5547 (N_5547,N_4969,N_4634);
nor U5548 (N_5548,N_4635,N_4983);
and U5549 (N_5549,N_4403,N_4711);
xor U5550 (N_5550,N_4653,N_4843);
or U5551 (N_5551,N_4541,N_4652);
or U5552 (N_5552,N_4622,N_4882);
nand U5553 (N_5553,N_4457,N_4722);
or U5554 (N_5554,N_4910,N_4818);
or U5555 (N_5555,N_4926,N_4732);
and U5556 (N_5556,N_4595,N_4843);
or U5557 (N_5557,N_4818,N_4807);
nor U5558 (N_5558,N_4723,N_4656);
or U5559 (N_5559,N_4889,N_4595);
nor U5560 (N_5560,N_4714,N_4457);
or U5561 (N_5561,N_4956,N_4577);
xnor U5562 (N_5562,N_4817,N_4548);
or U5563 (N_5563,N_4375,N_4737);
nor U5564 (N_5564,N_4931,N_4890);
nand U5565 (N_5565,N_4497,N_4712);
nor U5566 (N_5566,N_4750,N_4473);
and U5567 (N_5567,N_4446,N_4690);
nor U5568 (N_5568,N_4928,N_4966);
nand U5569 (N_5569,N_4937,N_4603);
nand U5570 (N_5570,N_4451,N_4975);
or U5571 (N_5571,N_4981,N_4876);
nor U5572 (N_5572,N_4391,N_4694);
and U5573 (N_5573,N_4996,N_4414);
nor U5574 (N_5574,N_4666,N_4915);
xor U5575 (N_5575,N_4474,N_4665);
and U5576 (N_5576,N_4693,N_4821);
nand U5577 (N_5577,N_4833,N_4669);
nor U5578 (N_5578,N_4833,N_4602);
xor U5579 (N_5579,N_4720,N_4918);
xnor U5580 (N_5580,N_4517,N_4832);
nor U5581 (N_5581,N_4814,N_4536);
and U5582 (N_5582,N_4728,N_4599);
and U5583 (N_5583,N_4583,N_4826);
and U5584 (N_5584,N_4837,N_4581);
or U5585 (N_5585,N_4563,N_4560);
nand U5586 (N_5586,N_4747,N_4420);
or U5587 (N_5587,N_4407,N_4930);
or U5588 (N_5588,N_4486,N_4817);
or U5589 (N_5589,N_4916,N_4497);
and U5590 (N_5590,N_4868,N_4603);
xnor U5591 (N_5591,N_4892,N_4770);
and U5592 (N_5592,N_4493,N_4850);
and U5593 (N_5593,N_4997,N_4516);
or U5594 (N_5594,N_4922,N_4670);
and U5595 (N_5595,N_4563,N_4927);
or U5596 (N_5596,N_4436,N_4427);
nand U5597 (N_5597,N_4763,N_4670);
or U5598 (N_5598,N_4763,N_4868);
nand U5599 (N_5599,N_4443,N_4690);
nor U5600 (N_5600,N_4660,N_4462);
and U5601 (N_5601,N_4723,N_4580);
nand U5602 (N_5602,N_4934,N_4837);
nor U5603 (N_5603,N_4455,N_4861);
or U5604 (N_5604,N_4510,N_4843);
nand U5605 (N_5605,N_4751,N_4862);
xor U5606 (N_5606,N_4520,N_4878);
nor U5607 (N_5607,N_4418,N_4643);
or U5608 (N_5608,N_4652,N_4519);
nor U5609 (N_5609,N_4820,N_4880);
and U5610 (N_5610,N_4976,N_4646);
nand U5611 (N_5611,N_4928,N_4720);
nor U5612 (N_5612,N_4922,N_4382);
xor U5613 (N_5613,N_4872,N_4887);
and U5614 (N_5614,N_4375,N_4851);
or U5615 (N_5615,N_4857,N_4713);
nand U5616 (N_5616,N_4695,N_4690);
nand U5617 (N_5617,N_4813,N_4900);
or U5618 (N_5618,N_4483,N_4804);
xnor U5619 (N_5619,N_4448,N_4866);
nor U5620 (N_5620,N_4864,N_4941);
nand U5621 (N_5621,N_4742,N_4414);
nand U5622 (N_5622,N_4528,N_4914);
nand U5623 (N_5623,N_4999,N_4847);
nor U5624 (N_5624,N_4546,N_4533);
nand U5625 (N_5625,N_5152,N_5339);
and U5626 (N_5626,N_5555,N_5460);
nand U5627 (N_5627,N_5397,N_5146);
nor U5628 (N_5628,N_5316,N_5264);
nor U5629 (N_5629,N_5014,N_5482);
and U5630 (N_5630,N_5396,N_5539);
or U5631 (N_5631,N_5170,N_5150);
nor U5632 (N_5632,N_5068,N_5403);
xor U5633 (N_5633,N_5375,N_5439);
xnor U5634 (N_5634,N_5153,N_5090);
or U5635 (N_5635,N_5112,N_5273);
xnor U5636 (N_5636,N_5192,N_5006);
or U5637 (N_5637,N_5425,N_5334);
or U5638 (N_5638,N_5459,N_5290);
nor U5639 (N_5639,N_5147,N_5394);
xor U5640 (N_5640,N_5285,N_5590);
and U5641 (N_5641,N_5293,N_5114);
and U5642 (N_5642,N_5343,N_5051);
and U5643 (N_5643,N_5234,N_5021);
xor U5644 (N_5644,N_5072,N_5347);
nor U5645 (N_5645,N_5284,N_5614);
or U5646 (N_5646,N_5549,N_5158);
nor U5647 (N_5647,N_5538,N_5389);
nor U5648 (N_5648,N_5229,N_5294);
xor U5649 (N_5649,N_5364,N_5097);
or U5650 (N_5650,N_5160,N_5455);
nor U5651 (N_5651,N_5180,N_5600);
nand U5652 (N_5652,N_5233,N_5620);
or U5653 (N_5653,N_5226,N_5082);
nand U5654 (N_5654,N_5186,N_5207);
nor U5655 (N_5655,N_5346,N_5584);
or U5656 (N_5656,N_5028,N_5208);
xor U5657 (N_5657,N_5517,N_5122);
nand U5658 (N_5658,N_5324,N_5052);
xnor U5659 (N_5659,N_5322,N_5504);
or U5660 (N_5660,N_5002,N_5509);
xnor U5661 (N_5661,N_5329,N_5070);
or U5662 (N_5662,N_5193,N_5280);
xnor U5663 (N_5663,N_5369,N_5444);
or U5664 (N_5664,N_5326,N_5304);
nor U5665 (N_5665,N_5348,N_5438);
nand U5666 (N_5666,N_5536,N_5022);
xor U5667 (N_5667,N_5136,N_5544);
xnor U5668 (N_5668,N_5479,N_5011);
nand U5669 (N_5669,N_5278,N_5173);
nand U5670 (N_5670,N_5378,N_5104);
xor U5671 (N_5671,N_5059,N_5416);
and U5672 (N_5672,N_5044,N_5521);
nand U5673 (N_5673,N_5530,N_5048);
xor U5674 (N_5674,N_5622,N_5528);
or U5675 (N_5675,N_5360,N_5015);
and U5676 (N_5676,N_5001,N_5610);
and U5677 (N_5677,N_5457,N_5286);
or U5678 (N_5678,N_5105,N_5300);
nand U5679 (N_5679,N_5215,N_5308);
or U5680 (N_5680,N_5239,N_5107);
xnor U5681 (N_5681,N_5100,N_5182);
nor U5682 (N_5682,N_5592,N_5237);
or U5683 (N_5683,N_5451,N_5143);
or U5684 (N_5684,N_5499,N_5349);
and U5685 (N_5685,N_5217,N_5311);
or U5686 (N_5686,N_5032,N_5593);
and U5687 (N_5687,N_5363,N_5566);
or U5688 (N_5688,N_5024,N_5253);
nor U5689 (N_5689,N_5008,N_5075);
and U5690 (N_5690,N_5195,N_5135);
xor U5691 (N_5691,N_5058,N_5354);
and U5692 (N_5692,N_5098,N_5310);
nor U5693 (N_5693,N_5385,N_5250);
and U5694 (N_5694,N_5529,N_5081);
nor U5695 (N_5695,N_5312,N_5427);
nor U5696 (N_5696,N_5483,N_5548);
or U5697 (N_5697,N_5174,N_5093);
xnor U5698 (N_5698,N_5206,N_5611);
nor U5699 (N_5699,N_5288,N_5040);
or U5700 (N_5700,N_5084,N_5062);
nand U5701 (N_5701,N_5413,N_5115);
and U5702 (N_5702,N_5057,N_5505);
and U5703 (N_5703,N_5337,N_5606);
or U5704 (N_5704,N_5313,N_5594);
xor U5705 (N_5705,N_5398,N_5242);
xor U5706 (N_5706,N_5128,N_5252);
nand U5707 (N_5707,N_5492,N_5224);
or U5708 (N_5708,N_5241,N_5332);
nor U5709 (N_5709,N_5302,N_5359);
xnor U5710 (N_5710,N_5401,N_5315);
xor U5711 (N_5711,N_5066,N_5127);
and U5712 (N_5712,N_5410,N_5513);
or U5713 (N_5713,N_5069,N_5448);
or U5714 (N_5714,N_5004,N_5543);
nor U5715 (N_5715,N_5254,N_5520);
nor U5716 (N_5716,N_5382,N_5596);
xnor U5717 (N_5717,N_5301,N_5166);
xor U5718 (N_5718,N_5564,N_5036);
xor U5719 (N_5719,N_5540,N_5550);
nor U5720 (N_5720,N_5263,N_5144);
nand U5721 (N_5721,N_5018,N_5575);
and U5722 (N_5722,N_5465,N_5613);
and U5723 (N_5723,N_5362,N_5039);
xnor U5724 (N_5724,N_5094,N_5007);
xnor U5725 (N_5725,N_5145,N_5212);
xnor U5726 (N_5726,N_5442,N_5446);
nand U5727 (N_5727,N_5189,N_5623);
nor U5728 (N_5728,N_5279,N_5141);
nor U5729 (N_5729,N_5231,N_5541);
nand U5730 (N_5730,N_5088,N_5076);
or U5731 (N_5731,N_5325,N_5087);
xor U5732 (N_5732,N_5441,N_5338);
nor U5733 (N_5733,N_5571,N_5466);
xor U5734 (N_5734,N_5522,N_5214);
and U5735 (N_5735,N_5276,N_5467);
and U5736 (N_5736,N_5443,N_5198);
xnor U5737 (N_5737,N_5110,N_5358);
xor U5738 (N_5738,N_5533,N_5546);
xnor U5739 (N_5739,N_5169,N_5244);
or U5740 (N_5740,N_5336,N_5568);
xor U5741 (N_5741,N_5025,N_5489);
and U5742 (N_5742,N_5352,N_5383);
nor U5743 (N_5743,N_5461,N_5624);
nor U5744 (N_5744,N_5232,N_5559);
nand U5745 (N_5745,N_5140,N_5381);
and U5746 (N_5746,N_5271,N_5038);
nor U5747 (N_5747,N_5341,N_5464);
nor U5748 (N_5748,N_5010,N_5267);
xnor U5749 (N_5749,N_5142,N_5556);
and U5750 (N_5750,N_5605,N_5209);
and U5751 (N_5751,N_5295,N_5366);
nand U5752 (N_5752,N_5256,N_5553);
xnor U5753 (N_5753,N_5474,N_5420);
nand U5754 (N_5754,N_5298,N_5299);
and U5755 (N_5755,N_5203,N_5612);
and U5756 (N_5756,N_5527,N_5395);
or U5757 (N_5757,N_5379,N_5603);
xnor U5758 (N_5758,N_5317,N_5204);
nor U5759 (N_5759,N_5132,N_5523);
xor U5760 (N_5760,N_5109,N_5570);
nor U5761 (N_5761,N_5196,N_5003);
and U5762 (N_5762,N_5604,N_5175);
nand U5763 (N_5763,N_5376,N_5230);
or U5764 (N_5764,N_5181,N_5292);
nor U5765 (N_5765,N_5257,N_5200);
or U5766 (N_5766,N_5481,N_5532);
and U5767 (N_5767,N_5092,N_5370);
xor U5768 (N_5768,N_5275,N_5557);
or U5769 (N_5769,N_5131,N_5320);
or U5770 (N_5770,N_5415,N_5503);
xnor U5771 (N_5771,N_5309,N_5477);
nor U5772 (N_5772,N_5056,N_5030);
or U5773 (N_5773,N_5095,N_5249);
nand U5774 (N_5774,N_5155,N_5029);
and U5775 (N_5775,N_5582,N_5574);
xor U5776 (N_5776,N_5490,N_5113);
nand U5777 (N_5777,N_5586,N_5418);
or U5778 (N_5778,N_5524,N_5351);
nand U5779 (N_5779,N_5134,N_5017);
xor U5780 (N_5780,N_5116,N_5118);
nor U5781 (N_5781,N_5183,N_5515);
xor U5782 (N_5782,N_5246,N_5205);
or U5783 (N_5783,N_5130,N_5297);
and U5784 (N_5784,N_5031,N_5473);
or U5785 (N_5785,N_5367,N_5424);
and U5786 (N_5786,N_5488,N_5458);
and U5787 (N_5787,N_5621,N_5595);
xor U5788 (N_5788,N_5120,N_5373);
nand U5789 (N_5789,N_5519,N_5615);
and U5790 (N_5790,N_5163,N_5080);
xor U5791 (N_5791,N_5086,N_5171);
nor U5792 (N_5792,N_5512,N_5486);
and U5793 (N_5793,N_5067,N_5073);
xor U5794 (N_5794,N_5357,N_5417);
nand U5795 (N_5795,N_5476,N_5321);
nor U5796 (N_5796,N_5043,N_5047);
nor U5797 (N_5797,N_5162,N_5077);
xor U5798 (N_5798,N_5422,N_5510);
nor U5799 (N_5799,N_5560,N_5129);
nor U5800 (N_5800,N_5269,N_5138);
nand U5801 (N_5801,N_5272,N_5384);
and U5802 (N_5802,N_5314,N_5185);
nor U5803 (N_5803,N_5400,N_5139);
nand U5804 (N_5804,N_5259,N_5434);
nand U5805 (N_5805,N_5583,N_5000);
or U5806 (N_5806,N_5149,N_5580);
xnor U5807 (N_5807,N_5071,N_5050);
xnor U5808 (N_5808,N_5391,N_5041);
and U5809 (N_5809,N_5074,N_5046);
and U5810 (N_5810,N_5303,N_5390);
and U5811 (N_5811,N_5371,N_5511);
xor U5812 (N_5812,N_5531,N_5101);
nand U5813 (N_5813,N_5585,N_5344);
nor U5814 (N_5814,N_5251,N_5618);
or U5815 (N_5815,N_5156,N_5350);
or U5816 (N_5816,N_5061,N_5305);
or U5817 (N_5817,N_5091,N_5405);
nand U5818 (N_5818,N_5194,N_5589);
or U5819 (N_5819,N_5291,N_5345);
or U5820 (N_5820,N_5188,N_5306);
and U5821 (N_5821,N_5581,N_5261);
and U5822 (N_5822,N_5111,N_5197);
and U5823 (N_5823,N_5216,N_5437);
or U5824 (N_5824,N_5587,N_5484);
nor U5825 (N_5825,N_5108,N_5565);
nor U5826 (N_5826,N_5609,N_5498);
and U5827 (N_5827,N_5494,N_5023);
or U5828 (N_5828,N_5463,N_5578);
or U5829 (N_5829,N_5330,N_5616);
and U5830 (N_5830,N_5191,N_5323);
or U5831 (N_5831,N_5372,N_5165);
or U5832 (N_5832,N_5012,N_5423);
nor U5833 (N_5833,N_5579,N_5608);
nor U5834 (N_5834,N_5119,N_5368);
nand U5835 (N_5835,N_5535,N_5121);
nor U5836 (N_5836,N_5393,N_5013);
and U5837 (N_5837,N_5500,N_5355);
and U5838 (N_5838,N_5563,N_5471);
xnor U5839 (N_5839,N_5270,N_5340);
nor U5840 (N_5840,N_5296,N_5307);
and U5841 (N_5841,N_5356,N_5265);
or U5842 (N_5842,N_5445,N_5268);
or U5843 (N_5843,N_5331,N_5419);
nor U5844 (N_5844,N_5462,N_5495);
and U5845 (N_5845,N_5392,N_5247);
nand U5846 (N_5846,N_5468,N_5408);
xor U5847 (N_5847,N_5377,N_5485);
nor U5848 (N_5848,N_5172,N_5187);
xor U5849 (N_5849,N_5552,N_5055);
and U5850 (N_5850,N_5106,N_5019);
nand U5851 (N_5851,N_5409,N_5042);
nor U5852 (N_5852,N_5026,N_5222);
nand U5853 (N_5853,N_5167,N_5262);
or U5854 (N_5854,N_5404,N_5274);
or U5855 (N_5855,N_5085,N_5440);
xor U5856 (N_5856,N_5619,N_5033);
and U5857 (N_5857,N_5064,N_5281);
nand U5858 (N_5858,N_5353,N_5238);
and U5859 (N_5859,N_5456,N_5223);
or U5860 (N_5860,N_5065,N_5202);
xnor U5861 (N_5861,N_5374,N_5447);
nand U5862 (N_5862,N_5201,N_5475);
or U5863 (N_5863,N_5289,N_5049);
and U5864 (N_5864,N_5430,N_5508);
xnor U5865 (N_5865,N_5449,N_5327);
and U5866 (N_5866,N_5588,N_5157);
nand U5867 (N_5867,N_5573,N_5099);
and U5868 (N_5868,N_5426,N_5009);
or U5869 (N_5869,N_5542,N_5027);
and U5870 (N_5870,N_5501,N_5283);
nor U5871 (N_5871,N_5514,N_5572);
nand U5872 (N_5872,N_5245,N_5388);
or U5873 (N_5873,N_5277,N_5037);
nand U5874 (N_5874,N_5617,N_5534);
xor U5875 (N_5875,N_5429,N_5126);
xnor U5876 (N_5876,N_5599,N_5255);
or U5877 (N_5877,N_5569,N_5591);
xnor U5878 (N_5878,N_5103,N_5266);
xor U5879 (N_5879,N_5387,N_5518);
xor U5880 (N_5880,N_5179,N_5450);
and U5881 (N_5881,N_5221,N_5054);
xnor U5882 (N_5882,N_5335,N_5016);
and U5883 (N_5883,N_5491,N_5365);
and U5884 (N_5884,N_5598,N_5497);
nor U5885 (N_5885,N_5034,N_5380);
nand U5886 (N_5886,N_5328,N_5402);
and U5887 (N_5887,N_5562,N_5361);
nor U5888 (N_5888,N_5453,N_5063);
nor U5889 (N_5889,N_5005,N_5399);
xnor U5890 (N_5890,N_5545,N_5537);
nor U5891 (N_5891,N_5176,N_5220);
or U5892 (N_5892,N_5597,N_5507);
xor U5893 (N_5893,N_5516,N_5333);
nor U5894 (N_5894,N_5102,N_5161);
nor U5895 (N_5895,N_5228,N_5525);
or U5896 (N_5896,N_5454,N_5258);
xnor U5897 (N_5897,N_5502,N_5412);
and U5898 (N_5898,N_5260,N_5577);
nor U5899 (N_5899,N_5117,N_5506);
nand U5900 (N_5900,N_5218,N_5601);
and U5901 (N_5901,N_5225,N_5083);
xnor U5902 (N_5902,N_5159,N_5020);
nor U5903 (N_5903,N_5551,N_5414);
xor U5904 (N_5904,N_5602,N_5428);
nand U5905 (N_5905,N_5411,N_5436);
and U5906 (N_5906,N_5240,N_5211);
and U5907 (N_5907,N_5235,N_5168);
xnor U5908 (N_5908,N_5236,N_5227);
xnor U5909 (N_5909,N_5190,N_5607);
nor U5910 (N_5910,N_5470,N_5526);
nor U5911 (N_5911,N_5213,N_5124);
nor U5912 (N_5912,N_5406,N_5219);
and U5913 (N_5913,N_5096,N_5547);
nor U5914 (N_5914,N_5487,N_5342);
xnor U5915 (N_5915,N_5576,N_5386);
xnor U5916 (N_5916,N_5469,N_5089);
nand U5917 (N_5917,N_5567,N_5243);
or U5918 (N_5918,N_5199,N_5035);
nand U5919 (N_5919,N_5177,N_5561);
xnor U5920 (N_5920,N_5452,N_5496);
xor U5921 (N_5921,N_5154,N_5210);
and U5922 (N_5922,N_5435,N_5318);
and U5923 (N_5923,N_5558,N_5433);
nor U5924 (N_5924,N_5184,N_5319);
nor U5925 (N_5925,N_5431,N_5472);
and U5926 (N_5926,N_5079,N_5053);
xnor U5927 (N_5927,N_5133,N_5287);
and U5928 (N_5928,N_5554,N_5248);
or U5929 (N_5929,N_5493,N_5432);
nand U5930 (N_5930,N_5178,N_5478);
nand U5931 (N_5931,N_5137,N_5407);
or U5932 (N_5932,N_5282,N_5125);
xor U5933 (N_5933,N_5148,N_5421);
nand U5934 (N_5934,N_5045,N_5078);
and U5935 (N_5935,N_5164,N_5060);
nor U5936 (N_5936,N_5480,N_5123);
nor U5937 (N_5937,N_5151,N_5256);
nor U5938 (N_5938,N_5399,N_5203);
nor U5939 (N_5939,N_5014,N_5333);
or U5940 (N_5940,N_5396,N_5303);
nor U5941 (N_5941,N_5512,N_5044);
and U5942 (N_5942,N_5277,N_5141);
nand U5943 (N_5943,N_5580,N_5480);
xor U5944 (N_5944,N_5282,N_5611);
nand U5945 (N_5945,N_5217,N_5587);
nor U5946 (N_5946,N_5054,N_5196);
or U5947 (N_5947,N_5091,N_5546);
nand U5948 (N_5948,N_5026,N_5227);
and U5949 (N_5949,N_5217,N_5327);
nand U5950 (N_5950,N_5379,N_5008);
nor U5951 (N_5951,N_5432,N_5611);
xnor U5952 (N_5952,N_5431,N_5601);
and U5953 (N_5953,N_5561,N_5582);
nand U5954 (N_5954,N_5402,N_5340);
or U5955 (N_5955,N_5044,N_5361);
and U5956 (N_5956,N_5478,N_5483);
xnor U5957 (N_5957,N_5461,N_5332);
nor U5958 (N_5958,N_5488,N_5190);
nand U5959 (N_5959,N_5500,N_5115);
nor U5960 (N_5960,N_5563,N_5528);
nand U5961 (N_5961,N_5370,N_5534);
nand U5962 (N_5962,N_5492,N_5543);
nand U5963 (N_5963,N_5149,N_5366);
and U5964 (N_5964,N_5327,N_5072);
and U5965 (N_5965,N_5530,N_5540);
xnor U5966 (N_5966,N_5206,N_5608);
or U5967 (N_5967,N_5183,N_5460);
nor U5968 (N_5968,N_5545,N_5123);
xnor U5969 (N_5969,N_5370,N_5263);
and U5970 (N_5970,N_5098,N_5451);
and U5971 (N_5971,N_5387,N_5217);
xor U5972 (N_5972,N_5448,N_5490);
nand U5973 (N_5973,N_5393,N_5553);
or U5974 (N_5974,N_5044,N_5268);
nor U5975 (N_5975,N_5048,N_5015);
and U5976 (N_5976,N_5062,N_5186);
and U5977 (N_5977,N_5110,N_5474);
nand U5978 (N_5978,N_5507,N_5381);
or U5979 (N_5979,N_5544,N_5476);
xnor U5980 (N_5980,N_5274,N_5394);
or U5981 (N_5981,N_5339,N_5128);
or U5982 (N_5982,N_5376,N_5416);
nor U5983 (N_5983,N_5606,N_5477);
xnor U5984 (N_5984,N_5440,N_5484);
or U5985 (N_5985,N_5585,N_5516);
nor U5986 (N_5986,N_5133,N_5231);
nor U5987 (N_5987,N_5038,N_5474);
nand U5988 (N_5988,N_5439,N_5105);
xor U5989 (N_5989,N_5040,N_5539);
or U5990 (N_5990,N_5557,N_5428);
or U5991 (N_5991,N_5573,N_5302);
nor U5992 (N_5992,N_5523,N_5080);
nand U5993 (N_5993,N_5126,N_5183);
nand U5994 (N_5994,N_5101,N_5243);
and U5995 (N_5995,N_5080,N_5104);
or U5996 (N_5996,N_5592,N_5020);
xor U5997 (N_5997,N_5472,N_5246);
nor U5998 (N_5998,N_5527,N_5441);
and U5999 (N_5999,N_5068,N_5533);
nor U6000 (N_6000,N_5212,N_5250);
xor U6001 (N_6001,N_5386,N_5490);
or U6002 (N_6002,N_5078,N_5248);
nor U6003 (N_6003,N_5002,N_5160);
xnor U6004 (N_6004,N_5194,N_5340);
nand U6005 (N_6005,N_5461,N_5295);
and U6006 (N_6006,N_5347,N_5378);
or U6007 (N_6007,N_5027,N_5180);
xor U6008 (N_6008,N_5370,N_5220);
or U6009 (N_6009,N_5258,N_5569);
nor U6010 (N_6010,N_5409,N_5235);
and U6011 (N_6011,N_5101,N_5050);
xor U6012 (N_6012,N_5614,N_5501);
and U6013 (N_6013,N_5412,N_5445);
or U6014 (N_6014,N_5429,N_5226);
xor U6015 (N_6015,N_5190,N_5411);
nand U6016 (N_6016,N_5140,N_5218);
xor U6017 (N_6017,N_5556,N_5428);
xor U6018 (N_6018,N_5105,N_5474);
nand U6019 (N_6019,N_5170,N_5624);
and U6020 (N_6020,N_5020,N_5422);
nand U6021 (N_6021,N_5511,N_5375);
or U6022 (N_6022,N_5333,N_5403);
nor U6023 (N_6023,N_5503,N_5309);
or U6024 (N_6024,N_5486,N_5207);
xor U6025 (N_6025,N_5530,N_5086);
xnor U6026 (N_6026,N_5517,N_5335);
and U6027 (N_6027,N_5076,N_5574);
xor U6028 (N_6028,N_5563,N_5459);
nor U6029 (N_6029,N_5175,N_5569);
nor U6030 (N_6030,N_5453,N_5032);
or U6031 (N_6031,N_5220,N_5227);
and U6032 (N_6032,N_5252,N_5432);
xnor U6033 (N_6033,N_5480,N_5252);
or U6034 (N_6034,N_5003,N_5398);
nor U6035 (N_6035,N_5142,N_5131);
xor U6036 (N_6036,N_5296,N_5559);
xnor U6037 (N_6037,N_5182,N_5123);
or U6038 (N_6038,N_5152,N_5371);
and U6039 (N_6039,N_5612,N_5327);
nand U6040 (N_6040,N_5244,N_5172);
nand U6041 (N_6041,N_5594,N_5553);
and U6042 (N_6042,N_5340,N_5560);
nand U6043 (N_6043,N_5002,N_5213);
xor U6044 (N_6044,N_5338,N_5267);
or U6045 (N_6045,N_5450,N_5549);
nor U6046 (N_6046,N_5092,N_5347);
and U6047 (N_6047,N_5153,N_5165);
or U6048 (N_6048,N_5033,N_5385);
and U6049 (N_6049,N_5259,N_5538);
xor U6050 (N_6050,N_5119,N_5019);
xor U6051 (N_6051,N_5539,N_5505);
nand U6052 (N_6052,N_5284,N_5251);
xor U6053 (N_6053,N_5536,N_5414);
or U6054 (N_6054,N_5520,N_5478);
and U6055 (N_6055,N_5132,N_5426);
or U6056 (N_6056,N_5473,N_5552);
nand U6057 (N_6057,N_5613,N_5219);
xnor U6058 (N_6058,N_5132,N_5608);
xor U6059 (N_6059,N_5375,N_5549);
or U6060 (N_6060,N_5298,N_5393);
xor U6061 (N_6061,N_5174,N_5070);
and U6062 (N_6062,N_5152,N_5500);
nand U6063 (N_6063,N_5190,N_5150);
nand U6064 (N_6064,N_5472,N_5285);
and U6065 (N_6065,N_5152,N_5501);
xor U6066 (N_6066,N_5189,N_5162);
or U6067 (N_6067,N_5049,N_5447);
and U6068 (N_6068,N_5433,N_5165);
and U6069 (N_6069,N_5010,N_5096);
nand U6070 (N_6070,N_5271,N_5263);
nand U6071 (N_6071,N_5240,N_5163);
nor U6072 (N_6072,N_5526,N_5591);
nand U6073 (N_6073,N_5426,N_5036);
or U6074 (N_6074,N_5100,N_5204);
and U6075 (N_6075,N_5549,N_5462);
or U6076 (N_6076,N_5409,N_5624);
nand U6077 (N_6077,N_5372,N_5257);
nand U6078 (N_6078,N_5557,N_5445);
or U6079 (N_6079,N_5030,N_5115);
or U6080 (N_6080,N_5092,N_5477);
or U6081 (N_6081,N_5294,N_5373);
and U6082 (N_6082,N_5211,N_5067);
xor U6083 (N_6083,N_5353,N_5160);
and U6084 (N_6084,N_5600,N_5588);
or U6085 (N_6085,N_5199,N_5286);
nor U6086 (N_6086,N_5375,N_5579);
nand U6087 (N_6087,N_5381,N_5020);
xnor U6088 (N_6088,N_5379,N_5113);
nor U6089 (N_6089,N_5414,N_5510);
nand U6090 (N_6090,N_5552,N_5452);
or U6091 (N_6091,N_5007,N_5186);
nor U6092 (N_6092,N_5499,N_5541);
xor U6093 (N_6093,N_5232,N_5223);
nor U6094 (N_6094,N_5457,N_5236);
nand U6095 (N_6095,N_5020,N_5615);
nor U6096 (N_6096,N_5411,N_5502);
nor U6097 (N_6097,N_5318,N_5054);
or U6098 (N_6098,N_5591,N_5241);
or U6099 (N_6099,N_5152,N_5248);
or U6100 (N_6100,N_5532,N_5175);
and U6101 (N_6101,N_5281,N_5179);
xnor U6102 (N_6102,N_5021,N_5193);
xor U6103 (N_6103,N_5518,N_5123);
and U6104 (N_6104,N_5040,N_5433);
or U6105 (N_6105,N_5049,N_5199);
xnor U6106 (N_6106,N_5149,N_5370);
xnor U6107 (N_6107,N_5394,N_5306);
and U6108 (N_6108,N_5410,N_5531);
or U6109 (N_6109,N_5145,N_5455);
and U6110 (N_6110,N_5330,N_5082);
nor U6111 (N_6111,N_5511,N_5513);
and U6112 (N_6112,N_5489,N_5286);
nand U6113 (N_6113,N_5236,N_5434);
and U6114 (N_6114,N_5420,N_5023);
xor U6115 (N_6115,N_5348,N_5347);
xor U6116 (N_6116,N_5440,N_5454);
and U6117 (N_6117,N_5582,N_5293);
xor U6118 (N_6118,N_5018,N_5337);
or U6119 (N_6119,N_5579,N_5453);
nand U6120 (N_6120,N_5024,N_5002);
or U6121 (N_6121,N_5382,N_5614);
xor U6122 (N_6122,N_5170,N_5546);
xnor U6123 (N_6123,N_5413,N_5232);
and U6124 (N_6124,N_5017,N_5338);
or U6125 (N_6125,N_5457,N_5034);
or U6126 (N_6126,N_5601,N_5476);
xnor U6127 (N_6127,N_5218,N_5309);
or U6128 (N_6128,N_5606,N_5321);
and U6129 (N_6129,N_5148,N_5330);
nor U6130 (N_6130,N_5304,N_5139);
nor U6131 (N_6131,N_5466,N_5584);
and U6132 (N_6132,N_5483,N_5597);
xnor U6133 (N_6133,N_5371,N_5278);
and U6134 (N_6134,N_5546,N_5237);
or U6135 (N_6135,N_5401,N_5011);
and U6136 (N_6136,N_5296,N_5152);
or U6137 (N_6137,N_5286,N_5453);
nand U6138 (N_6138,N_5495,N_5457);
and U6139 (N_6139,N_5449,N_5016);
or U6140 (N_6140,N_5129,N_5156);
nor U6141 (N_6141,N_5226,N_5124);
nand U6142 (N_6142,N_5615,N_5326);
and U6143 (N_6143,N_5569,N_5271);
and U6144 (N_6144,N_5569,N_5466);
xor U6145 (N_6145,N_5344,N_5499);
nand U6146 (N_6146,N_5474,N_5537);
nand U6147 (N_6147,N_5612,N_5135);
nand U6148 (N_6148,N_5054,N_5275);
or U6149 (N_6149,N_5550,N_5158);
and U6150 (N_6150,N_5318,N_5475);
nor U6151 (N_6151,N_5500,N_5398);
or U6152 (N_6152,N_5192,N_5146);
nand U6153 (N_6153,N_5428,N_5528);
nand U6154 (N_6154,N_5318,N_5553);
and U6155 (N_6155,N_5451,N_5355);
nor U6156 (N_6156,N_5408,N_5143);
xor U6157 (N_6157,N_5386,N_5254);
and U6158 (N_6158,N_5369,N_5192);
or U6159 (N_6159,N_5316,N_5363);
and U6160 (N_6160,N_5001,N_5169);
and U6161 (N_6161,N_5589,N_5587);
nor U6162 (N_6162,N_5006,N_5185);
xor U6163 (N_6163,N_5112,N_5389);
or U6164 (N_6164,N_5386,N_5023);
xnor U6165 (N_6165,N_5601,N_5054);
or U6166 (N_6166,N_5421,N_5086);
nor U6167 (N_6167,N_5189,N_5494);
nor U6168 (N_6168,N_5137,N_5496);
or U6169 (N_6169,N_5484,N_5107);
nand U6170 (N_6170,N_5174,N_5175);
and U6171 (N_6171,N_5401,N_5232);
nor U6172 (N_6172,N_5541,N_5445);
and U6173 (N_6173,N_5321,N_5181);
nand U6174 (N_6174,N_5411,N_5459);
or U6175 (N_6175,N_5160,N_5320);
xnor U6176 (N_6176,N_5186,N_5173);
nor U6177 (N_6177,N_5455,N_5464);
nand U6178 (N_6178,N_5123,N_5120);
or U6179 (N_6179,N_5070,N_5235);
nand U6180 (N_6180,N_5337,N_5323);
nor U6181 (N_6181,N_5379,N_5314);
or U6182 (N_6182,N_5144,N_5030);
and U6183 (N_6183,N_5445,N_5094);
and U6184 (N_6184,N_5328,N_5473);
and U6185 (N_6185,N_5027,N_5456);
nand U6186 (N_6186,N_5481,N_5156);
nor U6187 (N_6187,N_5541,N_5085);
and U6188 (N_6188,N_5299,N_5203);
nor U6189 (N_6189,N_5432,N_5474);
or U6190 (N_6190,N_5192,N_5368);
or U6191 (N_6191,N_5100,N_5057);
xor U6192 (N_6192,N_5119,N_5412);
and U6193 (N_6193,N_5034,N_5439);
nor U6194 (N_6194,N_5097,N_5171);
nor U6195 (N_6195,N_5038,N_5118);
or U6196 (N_6196,N_5243,N_5544);
xnor U6197 (N_6197,N_5138,N_5364);
xor U6198 (N_6198,N_5424,N_5324);
or U6199 (N_6199,N_5070,N_5332);
xnor U6200 (N_6200,N_5031,N_5235);
nor U6201 (N_6201,N_5225,N_5002);
xnor U6202 (N_6202,N_5094,N_5438);
nand U6203 (N_6203,N_5192,N_5204);
nand U6204 (N_6204,N_5359,N_5570);
and U6205 (N_6205,N_5312,N_5065);
nand U6206 (N_6206,N_5259,N_5235);
xor U6207 (N_6207,N_5407,N_5516);
xnor U6208 (N_6208,N_5476,N_5324);
xnor U6209 (N_6209,N_5172,N_5414);
xor U6210 (N_6210,N_5265,N_5577);
xnor U6211 (N_6211,N_5030,N_5182);
or U6212 (N_6212,N_5347,N_5040);
nor U6213 (N_6213,N_5531,N_5253);
nand U6214 (N_6214,N_5320,N_5030);
xnor U6215 (N_6215,N_5208,N_5096);
and U6216 (N_6216,N_5209,N_5157);
and U6217 (N_6217,N_5276,N_5568);
nor U6218 (N_6218,N_5540,N_5185);
xor U6219 (N_6219,N_5364,N_5524);
and U6220 (N_6220,N_5268,N_5494);
xnor U6221 (N_6221,N_5474,N_5184);
or U6222 (N_6222,N_5014,N_5563);
nand U6223 (N_6223,N_5231,N_5107);
and U6224 (N_6224,N_5511,N_5451);
nand U6225 (N_6225,N_5169,N_5099);
nor U6226 (N_6226,N_5246,N_5206);
or U6227 (N_6227,N_5005,N_5100);
xor U6228 (N_6228,N_5106,N_5444);
or U6229 (N_6229,N_5619,N_5381);
and U6230 (N_6230,N_5035,N_5258);
or U6231 (N_6231,N_5423,N_5095);
xnor U6232 (N_6232,N_5121,N_5297);
xor U6233 (N_6233,N_5375,N_5542);
nor U6234 (N_6234,N_5303,N_5471);
nand U6235 (N_6235,N_5022,N_5208);
nand U6236 (N_6236,N_5136,N_5429);
or U6237 (N_6237,N_5616,N_5203);
xor U6238 (N_6238,N_5301,N_5053);
nor U6239 (N_6239,N_5195,N_5449);
xor U6240 (N_6240,N_5512,N_5212);
or U6241 (N_6241,N_5474,N_5004);
or U6242 (N_6242,N_5204,N_5457);
xnor U6243 (N_6243,N_5191,N_5070);
or U6244 (N_6244,N_5167,N_5476);
nor U6245 (N_6245,N_5024,N_5287);
nand U6246 (N_6246,N_5164,N_5530);
xnor U6247 (N_6247,N_5573,N_5309);
nand U6248 (N_6248,N_5424,N_5369);
and U6249 (N_6249,N_5051,N_5312);
or U6250 (N_6250,N_5921,N_6013);
and U6251 (N_6251,N_6209,N_6247);
or U6252 (N_6252,N_5962,N_5754);
and U6253 (N_6253,N_6212,N_6043);
xor U6254 (N_6254,N_6142,N_5839);
xnor U6255 (N_6255,N_5648,N_5865);
and U6256 (N_6256,N_5737,N_5944);
or U6257 (N_6257,N_5976,N_6031);
and U6258 (N_6258,N_5804,N_6235);
and U6259 (N_6259,N_6105,N_5999);
or U6260 (N_6260,N_6125,N_5798);
nor U6261 (N_6261,N_5776,N_5964);
nand U6262 (N_6262,N_5629,N_5914);
nor U6263 (N_6263,N_5645,N_6195);
and U6264 (N_6264,N_5949,N_5799);
nand U6265 (N_6265,N_6210,N_5739);
or U6266 (N_6266,N_5992,N_5929);
nand U6267 (N_6267,N_6158,N_6090);
nand U6268 (N_6268,N_5980,N_6204);
xor U6269 (N_6269,N_6166,N_5651);
nand U6270 (N_6270,N_6131,N_6191);
or U6271 (N_6271,N_6099,N_6050);
and U6272 (N_6272,N_5632,N_6044);
and U6273 (N_6273,N_6192,N_5708);
xnor U6274 (N_6274,N_5781,N_6104);
xor U6275 (N_6275,N_5698,N_6205);
nand U6276 (N_6276,N_6024,N_5675);
xnor U6277 (N_6277,N_6095,N_6202);
nor U6278 (N_6278,N_5926,N_6138);
xnor U6279 (N_6279,N_5749,N_6059);
nand U6280 (N_6280,N_6122,N_5889);
nor U6281 (N_6281,N_5762,N_6182);
xor U6282 (N_6282,N_6121,N_5990);
and U6283 (N_6283,N_6034,N_5679);
nor U6284 (N_6284,N_6221,N_5968);
xor U6285 (N_6285,N_5907,N_6147);
xor U6286 (N_6286,N_5979,N_5630);
xor U6287 (N_6287,N_5726,N_6120);
xnor U6288 (N_6288,N_6075,N_5959);
and U6289 (N_6289,N_6133,N_5786);
and U6290 (N_6290,N_6234,N_5869);
xor U6291 (N_6291,N_6239,N_5783);
or U6292 (N_6292,N_5901,N_5759);
nand U6293 (N_6293,N_6010,N_6162);
and U6294 (N_6294,N_6241,N_5843);
nor U6295 (N_6295,N_6160,N_5970);
nor U6296 (N_6296,N_5676,N_5880);
xor U6297 (N_6297,N_5899,N_5920);
and U6298 (N_6298,N_6096,N_5707);
or U6299 (N_6299,N_5891,N_5647);
and U6300 (N_6300,N_6098,N_6069);
nand U6301 (N_6301,N_5915,N_5761);
and U6302 (N_6302,N_5823,N_6225);
nand U6303 (N_6303,N_6020,N_6079);
xnor U6304 (N_6304,N_5795,N_6179);
xor U6305 (N_6305,N_6129,N_5702);
and U6306 (N_6306,N_5866,N_5625);
or U6307 (N_6307,N_5948,N_5879);
xnor U6308 (N_6308,N_5740,N_5838);
nand U6309 (N_6309,N_6119,N_5956);
nor U6310 (N_6310,N_5775,N_5745);
and U6311 (N_6311,N_6177,N_5688);
and U6312 (N_6312,N_5757,N_6085);
or U6313 (N_6313,N_5764,N_6027);
xnor U6314 (N_6314,N_6189,N_6100);
and U6315 (N_6315,N_6106,N_5912);
xnor U6316 (N_6316,N_6054,N_5670);
or U6317 (N_6317,N_6170,N_6021);
and U6318 (N_6318,N_6201,N_6011);
xnor U6319 (N_6319,N_6245,N_6089);
nand U6320 (N_6320,N_5834,N_5807);
xnor U6321 (N_6321,N_5793,N_5677);
xnor U6322 (N_6322,N_5649,N_5927);
xor U6323 (N_6323,N_5953,N_6042);
nand U6324 (N_6324,N_5911,N_6101);
and U6325 (N_6325,N_6035,N_6128);
or U6326 (N_6326,N_5996,N_5709);
xnor U6327 (N_6327,N_6146,N_5682);
and U6328 (N_6328,N_5893,N_5868);
nand U6329 (N_6329,N_6180,N_5773);
and U6330 (N_6330,N_6033,N_5994);
or U6331 (N_6331,N_5767,N_6224);
and U6332 (N_6332,N_5882,N_5644);
xnor U6333 (N_6333,N_6176,N_5642);
nand U6334 (N_6334,N_5963,N_5972);
or U6335 (N_6335,N_5842,N_5934);
nor U6336 (N_6336,N_6134,N_5824);
xnor U6337 (N_6337,N_6073,N_6248);
or U6338 (N_6338,N_5669,N_5732);
and U6339 (N_6339,N_5835,N_6091);
nor U6340 (N_6340,N_5957,N_6055);
xor U6341 (N_6341,N_5631,N_5888);
nand U6342 (N_6342,N_6148,N_6082);
and U6343 (N_6343,N_5690,N_5995);
nand U6344 (N_6344,N_5771,N_5801);
nand U6345 (N_6345,N_6064,N_5906);
nor U6346 (N_6346,N_5815,N_5951);
nor U6347 (N_6347,N_5816,N_5731);
xnor U6348 (N_6348,N_5984,N_5827);
nor U6349 (N_6349,N_5678,N_5989);
xor U6350 (N_6350,N_5736,N_5637);
nor U6351 (N_6351,N_5925,N_5860);
nand U6352 (N_6352,N_5993,N_5693);
and U6353 (N_6353,N_6203,N_5974);
nand U6354 (N_6354,N_6214,N_5986);
or U6355 (N_6355,N_6000,N_6113);
or U6356 (N_6356,N_6041,N_6156);
xor U6357 (N_6357,N_5727,N_5700);
or U6358 (N_6358,N_5943,N_5640);
nand U6359 (N_6359,N_5768,N_5978);
and U6360 (N_6360,N_6040,N_5704);
nand U6361 (N_6361,N_6143,N_5661);
and U6362 (N_6362,N_5738,N_6001);
xor U6363 (N_6363,N_5777,N_5735);
nor U6364 (N_6364,N_6109,N_6222);
nor U6365 (N_6365,N_5940,N_6008);
xor U6366 (N_6366,N_5744,N_5683);
or U6367 (N_6367,N_6172,N_5876);
nand U6368 (N_6368,N_5803,N_5750);
or U6369 (N_6369,N_5998,N_5917);
nand U6370 (N_6370,N_6127,N_5766);
nand U6371 (N_6371,N_5903,N_6110);
xor U6372 (N_6372,N_5955,N_6047);
and U6373 (N_6373,N_6130,N_5942);
nor U6374 (N_6374,N_5982,N_5784);
nor U6375 (N_6375,N_5855,N_5910);
nand U6376 (N_6376,N_5890,N_5791);
nor U6377 (N_6377,N_6052,N_5691);
or U6378 (N_6378,N_5713,N_5985);
nand U6379 (N_6379,N_5812,N_5908);
and U6380 (N_6380,N_5819,N_6074);
xnor U6381 (N_6381,N_6220,N_5946);
nor U6382 (N_6382,N_6032,N_6174);
nand U6383 (N_6383,N_5806,N_6002);
nand U6384 (N_6384,N_5861,N_5696);
nor U6385 (N_6385,N_5765,N_5825);
xor U6386 (N_6386,N_6218,N_5805);
nor U6387 (N_6387,N_6036,N_5660);
and U6388 (N_6388,N_6194,N_5681);
and U6389 (N_6389,N_6080,N_6028);
nand U6390 (N_6390,N_6161,N_6223);
nand U6391 (N_6391,N_5808,N_5634);
or U6392 (N_6392,N_5818,N_5780);
or U6393 (N_6393,N_6173,N_5883);
and U6394 (N_6394,N_5846,N_6145);
and U6395 (N_6395,N_5706,N_5840);
or U6396 (N_6396,N_5877,N_5932);
nor U6397 (N_6397,N_6111,N_5699);
xnor U6398 (N_6398,N_6048,N_6149);
nor U6399 (N_6399,N_5774,N_5686);
or U6400 (N_6400,N_6165,N_5663);
nor U6401 (N_6401,N_5997,N_6155);
and U6402 (N_6402,N_5725,N_5639);
nor U6403 (N_6403,N_5730,N_6232);
xor U6404 (N_6404,N_6231,N_5811);
nand U6405 (N_6405,N_5752,N_6057);
xnor U6406 (N_6406,N_5703,N_6115);
or U6407 (N_6407,N_5931,N_5900);
nor U6408 (N_6408,N_6066,N_6003);
and U6409 (N_6409,N_5933,N_5652);
nand U6410 (N_6410,N_5817,N_5965);
nor U6411 (N_6411,N_6084,N_5831);
nand U6412 (N_6412,N_6188,N_5822);
or U6413 (N_6413,N_5664,N_6168);
or U6414 (N_6414,N_6198,N_6193);
nor U6415 (N_6415,N_5919,N_5733);
nor U6416 (N_6416,N_6217,N_5837);
and U6417 (N_6417,N_5820,N_5705);
xnor U6418 (N_6418,N_5859,N_6190);
nand U6419 (N_6419,N_5857,N_6025);
and U6420 (N_6420,N_6123,N_5960);
nor U6421 (N_6421,N_5654,N_6086);
or U6422 (N_6422,N_6094,N_5896);
nor U6423 (N_6423,N_6062,N_5719);
nand U6424 (N_6424,N_6227,N_6230);
nor U6425 (N_6425,N_6244,N_5694);
or U6426 (N_6426,N_6068,N_5672);
or U6427 (N_6427,N_5887,N_5844);
nand U6428 (N_6428,N_6012,N_5924);
nand U6429 (N_6429,N_5656,N_5836);
nor U6430 (N_6430,N_6117,N_5692);
or U6431 (N_6431,N_5747,N_5809);
nor U6432 (N_6432,N_5828,N_6164);
xor U6433 (N_6433,N_5711,N_6151);
xnor U6434 (N_6434,N_5653,N_6200);
nand U6435 (N_6435,N_6005,N_5797);
or U6436 (N_6436,N_5902,N_5981);
and U6437 (N_6437,N_6083,N_6116);
xor U6438 (N_6438,N_5714,N_5941);
or U6439 (N_6439,N_6077,N_5895);
and U6440 (N_6440,N_6067,N_5668);
nand U6441 (N_6441,N_6242,N_5717);
and U6442 (N_6442,N_5778,N_6141);
and U6443 (N_6443,N_6019,N_6118);
nand U6444 (N_6444,N_5851,N_6018);
xor U6445 (N_6445,N_6207,N_6184);
and U6446 (N_6446,N_5734,N_5770);
nor U6447 (N_6447,N_5958,N_5988);
or U6448 (N_6448,N_5787,N_5751);
or U6449 (N_6449,N_6006,N_6014);
nand U6450 (N_6450,N_6015,N_6140);
or U6451 (N_6451,N_6215,N_6004);
nand U6452 (N_6452,N_5687,N_5885);
nor U6453 (N_6453,N_6022,N_5830);
and U6454 (N_6454,N_5638,N_5950);
nor U6455 (N_6455,N_6093,N_5872);
or U6456 (N_6456,N_6124,N_5850);
nand U6457 (N_6457,N_5758,N_6092);
and U6458 (N_6458,N_5636,N_5897);
and U6459 (N_6459,N_5969,N_6152);
nor U6460 (N_6460,N_6211,N_6175);
xor U6461 (N_6461,N_5674,N_5841);
nor U6462 (N_6462,N_6107,N_6087);
nand U6463 (N_6463,N_6061,N_5665);
and U6464 (N_6464,N_6039,N_6017);
and U6465 (N_6465,N_5863,N_5881);
and U6466 (N_6466,N_5646,N_5847);
xor U6467 (N_6467,N_5680,N_5659);
nor U6468 (N_6468,N_5643,N_5782);
nand U6469 (N_6469,N_6169,N_5633);
nor U6470 (N_6470,N_6114,N_6163);
nor U6471 (N_6471,N_5785,N_6126);
or U6472 (N_6472,N_5862,N_5728);
xor U6473 (N_6473,N_5821,N_6216);
nor U6474 (N_6474,N_6154,N_6030);
nor U6475 (N_6475,N_6243,N_6186);
or U6476 (N_6476,N_6132,N_5802);
nor U6477 (N_6477,N_6144,N_5667);
nor U6478 (N_6478,N_6136,N_6171);
xor U6479 (N_6479,N_6135,N_6060);
or U6480 (N_6480,N_5789,N_5769);
and U6481 (N_6481,N_6237,N_6226);
xor U6482 (N_6482,N_5810,N_5918);
nand U6483 (N_6483,N_6246,N_6007);
xnor U6484 (N_6484,N_5871,N_5878);
xor U6485 (N_6485,N_6240,N_5800);
xor U6486 (N_6486,N_5853,N_5790);
nor U6487 (N_6487,N_5715,N_5695);
and U6488 (N_6488,N_5813,N_5721);
nand U6489 (N_6489,N_5814,N_5779);
and U6490 (N_6490,N_5685,N_5845);
or U6491 (N_6491,N_5874,N_5892);
nor U6492 (N_6492,N_5858,N_5936);
xnor U6493 (N_6493,N_5720,N_6229);
and U6494 (N_6494,N_5898,N_6238);
and U6495 (N_6495,N_5975,N_5864);
nand U6496 (N_6496,N_5666,N_6088);
xor U6497 (N_6497,N_5722,N_5973);
and U6498 (N_6498,N_5987,N_5947);
nor U6499 (N_6499,N_5833,N_6236);
and U6500 (N_6500,N_6139,N_5966);
nor U6501 (N_6501,N_6072,N_6097);
or U6502 (N_6502,N_5954,N_5673);
nand U6503 (N_6503,N_6159,N_5635);
or U6504 (N_6504,N_5939,N_6009);
or U6505 (N_6505,N_5655,N_6197);
or U6506 (N_6506,N_5753,N_6029);
xor U6507 (N_6507,N_5961,N_6228);
nand U6508 (N_6508,N_5792,N_6023);
nor U6509 (N_6509,N_6070,N_5849);
or U6510 (N_6510,N_5716,N_5971);
xnor U6511 (N_6511,N_5697,N_6108);
nand U6512 (N_6512,N_5875,N_6026);
nand U6513 (N_6513,N_5712,N_5909);
nor U6514 (N_6514,N_6181,N_5904);
or U6515 (N_6515,N_6058,N_6016);
nor U6516 (N_6516,N_5742,N_6053);
or U6517 (N_6517,N_6056,N_5689);
and U6518 (N_6518,N_5627,N_5935);
xor U6519 (N_6519,N_5748,N_5626);
and U6520 (N_6520,N_5913,N_6233);
nand U6521 (N_6521,N_6076,N_6051);
or U6522 (N_6522,N_6178,N_6199);
xnor U6523 (N_6523,N_5894,N_5952);
nand U6524 (N_6524,N_5788,N_6150);
or U6525 (N_6525,N_6049,N_6208);
nand U6526 (N_6526,N_5867,N_5723);
nand U6527 (N_6527,N_5854,N_5873);
xor U6528 (N_6528,N_5641,N_5991);
nand U6529 (N_6529,N_5662,N_5657);
nor U6530 (N_6530,N_6157,N_5755);
xor U6531 (N_6531,N_5848,N_6046);
nor U6532 (N_6532,N_6078,N_5650);
nand U6533 (N_6533,N_6112,N_5763);
and U6534 (N_6534,N_6071,N_6187);
xor U6535 (N_6535,N_6249,N_5856);
or U6536 (N_6536,N_5826,N_5922);
or U6537 (N_6537,N_5756,N_6045);
xor U6538 (N_6538,N_5724,N_6213);
xor U6539 (N_6539,N_6038,N_6137);
and U6540 (N_6540,N_5760,N_5884);
nand U6541 (N_6541,N_5870,N_6102);
xor U6542 (N_6542,N_6081,N_5905);
or U6543 (N_6543,N_5983,N_6185);
nand U6544 (N_6544,N_5796,N_5938);
nand U6545 (N_6545,N_5746,N_6153);
xor U6546 (N_6546,N_6219,N_5794);
nand U6547 (N_6547,N_6063,N_5967);
nor U6548 (N_6548,N_5743,N_5671);
xor U6549 (N_6549,N_6103,N_6037);
nor U6550 (N_6550,N_5684,N_5937);
xnor U6551 (N_6551,N_5741,N_6196);
nand U6552 (N_6552,N_5923,N_5886);
nand U6553 (N_6553,N_5772,N_5628);
and U6554 (N_6554,N_5916,N_6065);
xor U6555 (N_6555,N_5945,N_5658);
or U6556 (N_6556,N_5729,N_5930);
nand U6557 (N_6557,N_6167,N_5829);
xnor U6558 (N_6558,N_5852,N_6183);
and U6559 (N_6559,N_5832,N_5718);
nand U6560 (N_6560,N_6206,N_5701);
nand U6561 (N_6561,N_5710,N_5977);
and U6562 (N_6562,N_5928,N_5705);
and U6563 (N_6563,N_5942,N_5812);
xor U6564 (N_6564,N_6168,N_6182);
nor U6565 (N_6565,N_6018,N_5662);
nand U6566 (N_6566,N_6101,N_5937);
or U6567 (N_6567,N_5753,N_6103);
nor U6568 (N_6568,N_6095,N_6135);
and U6569 (N_6569,N_6124,N_5942);
nor U6570 (N_6570,N_5855,N_5992);
nor U6571 (N_6571,N_6090,N_5747);
nand U6572 (N_6572,N_6068,N_5957);
nand U6573 (N_6573,N_5807,N_6152);
or U6574 (N_6574,N_6055,N_5842);
or U6575 (N_6575,N_6128,N_6040);
and U6576 (N_6576,N_5778,N_5904);
xnor U6577 (N_6577,N_6243,N_5889);
and U6578 (N_6578,N_5918,N_5966);
xor U6579 (N_6579,N_5832,N_5958);
xnor U6580 (N_6580,N_5803,N_6197);
xnor U6581 (N_6581,N_6005,N_5841);
and U6582 (N_6582,N_5829,N_6165);
nand U6583 (N_6583,N_5634,N_6000);
or U6584 (N_6584,N_5845,N_6057);
and U6585 (N_6585,N_6205,N_5874);
nand U6586 (N_6586,N_5731,N_6066);
xnor U6587 (N_6587,N_5812,N_6227);
and U6588 (N_6588,N_6153,N_5752);
xor U6589 (N_6589,N_5784,N_5734);
or U6590 (N_6590,N_6218,N_5913);
nor U6591 (N_6591,N_5824,N_5831);
xor U6592 (N_6592,N_5994,N_5785);
xor U6593 (N_6593,N_5819,N_5749);
nand U6594 (N_6594,N_6017,N_6214);
nor U6595 (N_6595,N_5845,N_5927);
nand U6596 (N_6596,N_6143,N_5816);
nand U6597 (N_6597,N_5738,N_5865);
and U6598 (N_6598,N_5861,N_6230);
xor U6599 (N_6599,N_5717,N_5845);
or U6600 (N_6600,N_5880,N_5804);
xor U6601 (N_6601,N_5900,N_6185);
nand U6602 (N_6602,N_6056,N_6104);
or U6603 (N_6603,N_5829,N_6152);
and U6604 (N_6604,N_5747,N_6016);
or U6605 (N_6605,N_5764,N_5783);
xnor U6606 (N_6606,N_5906,N_5880);
nor U6607 (N_6607,N_6071,N_5692);
or U6608 (N_6608,N_5845,N_6098);
nor U6609 (N_6609,N_5951,N_6131);
or U6610 (N_6610,N_5969,N_6140);
nor U6611 (N_6611,N_5716,N_5625);
and U6612 (N_6612,N_6150,N_6173);
and U6613 (N_6613,N_5907,N_5996);
and U6614 (N_6614,N_6004,N_5867);
xnor U6615 (N_6615,N_6242,N_5783);
and U6616 (N_6616,N_6060,N_6063);
or U6617 (N_6617,N_6134,N_5653);
and U6618 (N_6618,N_6113,N_5831);
nor U6619 (N_6619,N_5692,N_5759);
xnor U6620 (N_6620,N_5662,N_6148);
or U6621 (N_6621,N_5738,N_5786);
nand U6622 (N_6622,N_5816,N_6165);
xnor U6623 (N_6623,N_6222,N_6212);
nand U6624 (N_6624,N_5736,N_5979);
nor U6625 (N_6625,N_5732,N_6178);
or U6626 (N_6626,N_5797,N_6208);
nor U6627 (N_6627,N_6050,N_5764);
nor U6628 (N_6628,N_6152,N_5871);
and U6629 (N_6629,N_5848,N_5952);
nor U6630 (N_6630,N_5701,N_5854);
and U6631 (N_6631,N_5656,N_6043);
nor U6632 (N_6632,N_5640,N_5796);
or U6633 (N_6633,N_5659,N_5951);
nor U6634 (N_6634,N_5725,N_6030);
nor U6635 (N_6635,N_6079,N_6203);
and U6636 (N_6636,N_6167,N_6010);
and U6637 (N_6637,N_6019,N_5855);
and U6638 (N_6638,N_6190,N_5682);
and U6639 (N_6639,N_5829,N_6072);
nand U6640 (N_6640,N_6161,N_6024);
nor U6641 (N_6641,N_5654,N_5826);
xor U6642 (N_6642,N_6025,N_5851);
and U6643 (N_6643,N_5917,N_5945);
nor U6644 (N_6644,N_5855,N_5946);
nand U6645 (N_6645,N_6248,N_5843);
or U6646 (N_6646,N_5968,N_6042);
nand U6647 (N_6647,N_6099,N_6211);
xnor U6648 (N_6648,N_6249,N_5648);
nor U6649 (N_6649,N_5952,N_5739);
xnor U6650 (N_6650,N_6076,N_6131);
nor U6651 (N_6651,N_5796,N_6220);
xor U6652 (N_6652,N_6110,N_6003);
nand U6653 (N_6653,N_5792,N_5713);
or U6654 (N_6654,N_6145,N_5967);
nand U6655 (N_6655,N_5976,N_6188);
xor U6656 (N_6656,N_5987,N_5664);
xnor U6657 (N_6657,N_5900,N_5646);
or U6658 (N_6658,N_5844,N_6195);
or U6659 (N_6659,N_5926,N_5915);
nand U6660 (N_6660,N_5848,N_5781);
xnor U6661 (N_6661,N_6219,N_5679);
nor U6662 (N_6662,N_6228,N_6059);
and U6663 (N_6663,N_5877,N_5921);
or U6664 (N_6664,N_5979,N_6077);
nor U6665 (N_6665,N_5797,N_5762);
nor U6666 (N_6666,N_6107,N_6145);
nor U6667 (N_6667,N_5765,N_6190);
and U6668 (N_6668,N_5864,N_6024);
xnor U6669 (N_6669,N_5841,N_6213);
nand U6670 (N_6670,N_5912,N_6063);
nand U6671 (N_6671,N_6154,N_6071);
and U6672 (N_6672,N_5850,N_5656);
or U6673 (N_6673,N_5873,N_6248);
xor U6674 (N_6674,N_5852,N_5822);
nor U6675 (N_6675,N_6180,N_6199);
or U6676 (N_6676,N_5697,N_5662);
or U6677 (N_6677,N_6068,N_5656);
or U6678 (N_6678,N_6091,N_6002);
nand U6679 (N_6679,N_5709,N_6232);
nor U6680 (N_6680,N_5653,N_6167);
xnor U6681 (N_6681,N_5694,N_5735);
xnor U6682 (N_6682,N_5958,N_5653);
or U6683 (N_6683,N_5772,N_6091);
and U6684 (N_6684,N_5650,N_5686);
or U6685 (N_6685,N_5903,N_6098);
or U6686 (N_6686,N_5854,N_5716);
xor U6687 (N_6687,N_6151,N_6235);
nor U6688 (N_6688,N_5724,N_6056);
xor U6689 (N_6689,N_6205,N_6202);
nand U6690 (N_6690,N_6188,N_6184);
xnor U6691 (N_6691,N_5900,N_6227);
or U6692 (N_6692,N_6000,N_5704);
and U6693 (N_6693,N_5956,N_5957);
xnor U6694 (N_6694,N_5647,N_5878);
nor U6695 (N_6695,N_5996,N_6151);
xnor U6696 (N_6696,N_5795,N_6082);
nand U6697 (N_6697,N_6154,N_6051);
nor U6698 (N_6698,N_5686,N_5653);
and U6699 (N_6699,N_6059,N_5885);
or U6700 (N_6700,N_6015,N_5931);
nand U6701 (N_6701,N_6074,N_5931);
nor U6702 (N_6702,N_6043,N_6156);
or U6703 (N_6703,N_5851,N_6099);
nand U6704 (N_6704,N_5954,N_5939);
or U6705 (N_6705,N_5817,N_5632);
nand U6706 (N_6706,N_5757,N_5947);
or U6707 (N_6707,N_5977,N_5718);
xor U6708 (N_6708,N_5671,N_5865);
xnor U6709 (N_6709,N_5710,N_6221);
nor U6710 (N_6710,N_6049,N_6121);
nor U6711 (N_6711,N_5907,N_5978);
and U6712 (N_6712,N_5899,N_5701);
nor U6713 (N_6713,N_6222,N_6218);
nor U6714 (N_6714,N_5726,N_5844);
nor U6715 (N_6715,N_5790,N_6096);
nand U6716 (N_6716,N_5876,N_5905);
nor U6717 (N_6717,N_6066,N_5915);
and U6718 (N_6718,N_6220,N_6044);
or U6719 (N_6719,N_5698,N_6187);
nand U6720 (N_6720,N_6185,N_6131);
or U6721 (N_6721,N_5699,N_5737);
nor U6722 (N_6722,N_5662,N_5630);
nand U6723 (N_6723,N_5637,N_6150);
xor U6724 (N_6724,N_5994,N_6119);
and U6725 (N_6725,N_6090,N_5844);
nand U6726 (N_6726,N_6188,N_6149);
xor U6727 (N_6727,N_5852,N_5866);
nor U6728 (N_6728,N_6196,N_5748);
or U6729 (N_6729,N_5719,N_6183);
xor U6730 (N_6730,N_6032,N_5700);
and U6731 (N_6731,N_5720,N_6023);
or U6732 (N_6732,N_5641,N_5885);
and U6733 (N_6733,N_5646,N_5786);
and U6734 (N_6734,N_5882,N_6186);
nor U6735 (N_6735,N_5923,N_5977);
xnor U6736 (N_6736,N_5995,N_5729);
or U6737 (N_6737,N_6133,N_6057);
nor U6738 (N_6738,N_6077,N_5756);
and U6739 (N_6739,N_6098,N_5775);
nand U6740 (N_6740,N_5923,N_5710);
or U6741 (N_6741,N_6189,N_5863);
and U6742 (N_6742,N_5945,N_6191);
xor U6743 (N_6743,N_6217,N_5770);
nand U6744 (N_6744,N_6095,N_5743);
xor U6745 (N_6745,N_5672,N_6007);
and U6746 (N_6746,N_5738,N_5924);
xor U6747 (N_6747,N_6071,N_6004);
xor U6748 (N_6748,N_6152,N_6201);
nand U6749 (N_6749,N_6056,N_6125);
xnor U6750 (N_6750,N_5772,N_5826);
or U6751 (N_6751,N_6028,N_6130);
or U6752 (N_6752,N_6102,N_5843);
and U6753 (N_6753,N_5675,N_5850);
and U6754 (N_6754,N_6115,N_6246);
or U6755 (N_6755,N_5823,N_5873);
nand U6756 (N_6756,N_6052,N_6249);
and U6757 (N_6757,N_6072,N_5956);
or U6758 (N_6758,N_6069,N_5881);
xor U6759 (N_6759,N_6077,N_5944);
nor U6760 (N_6760,N_5888,N_6106);
xnor U6761 (N_6761,N_5755,N_5992);
nand U6762 (N_6762,N_5950,N_6222);
nand U6763 (N_6763,N_6023,N_5648);
nand U6764 (N_6764,N_5728,N_5781);
and U6765 (N_6765,N_6085,N_6171);
nand U6766 (N_6766,N_5815,N_6079);
or U6767 (N_6767,N_5885,N_5827);
nor U6768 (N_6768,N_5946,N_6121);
nand U6769 (N_6769,N_6063,N_5661);
and U6770 (N_6770,N_5721,N_5682);
xor U6771 (N_6771,N_5763,N_5837);
nand U6772 (N_6772,N_6004,N_5700);
nand U6773 (N_6773,N_6129,N_5936);
nor U6774 (N_6774,N_5729,N_6059);
or U6775 (N_6775,N_6195,N_6055);
xor U6776 (N_6776,N_6067,N_5848);
xor U6777 (N_6777,N_5648,N_5926);
nand U6778 (N_6778,N_5702,N_5699);
nor U6779 (N_6779,N_6209,N_6002);
nand U6780 (N_6780,N_5985,N_5895);
xor U6781 (N_6781,N_6030,N_5629);
nor U6782 (N_6782,N_5945,N_6078);
nand U6783 (N_6783,N_5941,N_5871);
and U6784 (N_6784,N_6181,N_5884);
nand U6785 (N_6785,N_5674,N_5635);
nor U6786 (N_6786,N_6141,N_5788);
or U6787 (N_6787,N_5762,N_5721);
nor U6788 (N_6788,N_6147,N_5668);
or U6789 (N_6789,N_5667,N_5990);
nand U6790 (N_6790,N_5706,N_6071);
and U6791 (N_6791,N_5676,N_6175);
xor U6792 (N_6792,N_5994,N_5888);
xor U6793 (N_6793,N_5854,N_5997);
xor U6794 (N_6794,N_5741,N_5932);
nand U6795 (N_6795,N_5818,N_6031);
nand U6796 (N_6796,N_5925,N_5678);
or U6797 (N_6797,N_5730,N_5896);
or U6798 (N_6798,N_5709,N_5920);
nor U6799 (N_6799,N_6064,N_6242);
xnor U6800 (N_6800,N_5628,N_5912);
and U6801 (N_6801,N_6012,N_5884);
nor U6802 (N_6802,N_5776,N_5761);
and U6803 (N_6803,N_5970,N_5766);
and U6804 (N_6804,N_5857,N_5808);
nor U6805 (N_6805,N_6247,N_5735);
nor U6806 (N_6806,N_5941,N_5660);
nand U6807 (N_6807,N_5689,N_6037);
xnor U6808 (N_6808,N_5995,N_5907);
xnor U6809 (N_6809,N_5831,N_5673);
and U6810 (N_6810,N_5644,N_5758);
xnor U6811 (N_6811,N_6060,N_6124);
nand U6812 (N_6812,N_5893,N_6066);
nand U6813 (N_6813,N_5639,N_6146);
xor U6814 (N_6814,N_5836,N_6144);
or U6815 (N_6815,N_6202,N_5817);
nand U6816 (N_6816,N_5945,N_6047);
and U6817 (N_6817,N_6030,N_5733);
and U6818 (N_6818,N_6046,N_6163);
or U6819 (N_6819,N_6193,N_5638);
xor U6820 (N_6820,N_6119,N_5684);
and U6821 (N_6821,N_6061,N_6032);
or U6822 (N_6822,N_6082,N_6223);
nor U6823 (N_6823,N_6156,N_6107);
nand U6824 (N_6824,N_5667,N_5870);
nor U6825 (N_6825,N_5808,N_6243);
nor U6826 (N_6826,N_5772,N_6108);
and U6827 (N_6827,N_6166,N_5723);
nand U6828 (N_6828,N_5687,N_5812);
xnor U6829 (N_6829,N_6125,N_5975);
and U6830 (N_6830,N_5787,N_6197);
xor U6831 (N_6831,N_5773,N_5882);
or U6832 (N_6832,N_5786,N_5833);
or U6833 (N_6833,N_5885,N_5905);
or U6834 (N_6834,N_6110,N_5986);
or U6835 (N_6835,N_5722,N_6188);
xor U6836 (N_6836,N_6213,N_6182);
nand U6837 (N_6837,N_6232,N_5847);
and U6838 (N_6838,N_6108,N_5850);
and U6839 (N_6839,N_5790,N_6040);
nand U6840 (N_6840,N_5985,N_5932);
and U6841 (N_6841,N_5679,N_6009);
xor U6842 (N_6842,N_5666,N_5742);
xor U6843 (N_6843,N_6035,N_6159);
or U6844 (N_6844,N_5755,N_5863);
or U6845 (N_6845,N_5705,N_6014);
xnor U6846 (N_6846,N_5677,N_6124);
nand U6847 (N_6847,N_6120,N_6215);
and U6848 (N_6848,N_5824,N_5702);
and U6849 (N_6849,N_5999,N_5789);
nor U6850 (N_6850,N_6060,N_5668);
nand U6851 (N_6851,N_5659,N_5688);
xnor U6852 (N_6852,N_5743,N_5995);
nand U6853 (N_6853,N_5837,N_5726);
nand U6854 (N_6854,N_6116,N_5631);
and U6855 (N_6855,N_5723,N_5698);
and U6856 (N_6856,N_5831,N_5915);
and U6857 (N_6857,N_5967,N_6012);
and U6858 (N_6858,N_6188,N_6198);
nand U6859 (N_6859,N_5921,N_5957);
or U6860 (N_6860,N_5657,N_5823);
nand U6861 (N_6861,N_5711,N_6239);
and U6862 (N_6862,N_5910,N_5746);
nor U6863 (N_6863,N_5667,N_6246);
nor U6864 (N_6864,N_6047,N_5668);
nor U6865 (N_6865,N_5849,N_6155);
or U6866 (N_6866,N_5721,N_5843);
xor U6867 (N_6867,N_5976,N_6043);
and U6868 (N_6868,N_6210,N_5659);
xnor U6869 (N_6869,N_6012,N_5642);
and U6870 (N_6870,N_6140,N_5950);
and U6871 (N_6871,N_5866,N_5999);
nand U6872 (N_6872,N_5753,N_5792);
nor U6873 (N_6873,N_5738,N_5757);
nor U6874 (N_6874,N_6085,N_5662);
nor U6875 (N_6875,N_6439,N_6529);
or U6876 (N_6876,N_6838,N_6555);
and U6877 (N_6877,N_6447,N_6738);
xor U6878 (N_6878,N_6771,N_6305);
xor U6879 (N_6879,N_6862,N_6369);
nor U6880 (N_6880,N_6778,N_6252);
xor U6881 (N_6881,N_6380,N_6490);
or U6882 (N_6882,N_6455,N_6541);
xor U6883 (N_6883,N_6390,N_6719);
or U6884 (N_6884,N_6621,N_6832);
nand U6885 (N_6885,N_6564,N_6487);
xor U6886 (N_6886,N_6589,N_6301);
or U6887 (N_6887,N_6826,N_6797);
or U6888 (N_6888,N_6553,N_6474);
or U6889 (N_6889,N_6491,N_6450);
nand U6890 (N_6890,N_6385,N_6693);
nand U6891 (N_6891,N_6342,N_6469);
nor U6892 (N_6892,N_6570,N_6731);
or U6893 (N_6893,N_6349,N_6427);
xnor U6894 (N_6894,N_6857,N_6560);
nor U6895 (N_6895,N_6300,N_6394);
nand U6896 (N_6896,N_6790,N_6714);
and U6897 (N_6897,N_6429,N_6355);
or U6898 (N_6898,N_6303,N_6255);
xnor U6899 (N_6899,N_6859,N_6651);
nand U6900 (N_6900,N_6416,N_6730);
or U6901 (N_6901,N_6554,N_6792);
nand U6902 (N_6902,N_6708,N_6434);
or U6903 (N_6903,N_6690,N_6291);
and U6904 (N_6904,N_6315,N_6330);
and U6905 (N_6905,N_6532,N_6260);
nor U6906 (N_6906,N_6298,N_6648);
or U6907 (N_6907,N_6584,N_6729);
and U6908 (N_6908,N_6578,N_6277);
or U6909 (N_6909,N_6765,N_6443);
nor U6910 (N_6910,N_6257,N_6863);
and U6911 (N_6911,N_6865,N_6759);
nand U6912 (N_6912,N_6327,N_6854);
and U6913 (N_6913,N_6425,N_6374);
nor U6914 (N_6914,N_6670,N_6281);
nor U6915 (N_6915,N_6351,N_6637);
nand U6916 (N_6916,N_6326,N_6420);
nor U6917 (N_6917,N_6353,N_6806);
and U6918 (N_6918,N_6754,N_6509);
xor U6919 (N_6919,N_6537,N_6461);
and U6920 (N_6920,N_6467,N_6337);
xor U6921 (N_6921,N_6830,N_6557);
nand U6922 (N_6922,N_6611,N_6649);
nand U6923 (N_6923,N_6415,N_6638);
nor U6924 (N_6924,N_6746,N_6744);
or U6925 (N_6925,N_6696,N_6251);
nor U6926 (N_6926,N_6462,N_6678);
or U6927 (N_6927,N_6680,N_6536);
xor U6928 (N_6928,N_6668,N_6727);
nor U6929 (N_6929,N_6659,N_6375);
and U6930 (N_6930,N_6336,N_6386);
and U6931 (N_6931,N_6606,N_6254);
and U6932 (N_6932,N_6413,N_6250);
or U6933 (N_6933,N_6702,N_6525);
nand U6934 (N_6934,N_6773,N_6829);
and U6935 (N_6935,N_6500,N_6675);
nor U6936 (N_6936,N_6745,N_6382);
nor U6937 (N_6937,N_6275,N_6314);
or U6938 (N_6938,N_6800,N_6840);
xnor U6939 (N_6939,N_6282,N_6712);
nand U6940 (N_6940,N_6607,N_6267);
and U6941 (N_6941,N_6852,N_6341);
xor U6942 (N_6942,N_6789,N_6313);
xnor U6943 (N_6943,N_6361,N_6444);
and U6944 (N_6944,N_6815,N_6694);
and U6945 (N_6945,N_6582,N_6835);
nand U6946 (N_6946,N_6470,N_6645);
xor U6947 (N_6947,N_6565,N_6686);
xnor U6948 (N_6948,N_6808,N_6288);
nand U6949 (N_6949,N_6665,N_6290);
xor U6950 (N_6950,N_6307,N_6874);
nor U6951 (N_6951,N_6843,N_6325);
nand U6952 (N_6952,N_6263,N_6398);
or U6953 (N_6953,N_6262,N_6407);
and U6954 (N_6954,N_6817,N_6869);
nand U6955 (N_6955,N_6734,N_6436);
nand U6956 (N_6956,N_6844,N_6741);
xnor U6957 (N_6957,N_6259,N_6373);
nand U6958 (N_6958,N_6867,N_6716);
and U6959 (N_6959,N_6454,N_6763);
nand U6960 (N_6960,N_6639,N_6682);
nand U6961 (N_6961,N_6404,N_6518);
or U6962 (N_6962,N_6842,N_6776);
and U6963 (N_6963,N_6476,N_6748);
nand U6964 (N_6964,N_6486,N_6624);
and U6965 (N_6965,N_6547,N_6562);
and U6966 (N_6966,N_6484,N_6475);
nand U6967 (N_6967,N_6673,N_6728);
or U6968 (N_6968,N_6586,N_6660);
xnor U6969 (N_6969,N_6677,N_6726);
nand U6970 (N_6970,N_6563,N_6317);
nand U6971 (N_6971,N_6402,N_6293);
or U6972 (N_6972,N_6850,N_6699);
or U6973 (N_6973,N_6704,N_6253);
nor U6974 (N_6974,N_6695,N_6672);
xor U6975 (N_6975,N_6451,N_6831);
nor U6976 (N_6976,N_6350,N_6456);
nor U6977 (N_6977,N_6412,N_6709);
nand U6978 (N_6978,N_6362,N_6600);
nand U6979 (N_6979,N_6596,N_6825);
and U6980 (N_6980,N_6737,N_6723);
nand U6981 (N_6981,N_6662,N_6417);
or U6982 (N_6982,N_6756,N_6583);
or U6983 (N_6983,N_6309,N_6345);
nand U6984 (N_6984,N_6616,N_6711);
xnor U6985 (N_6985,N_6318,N_6548);
and U6986 (N_6986,N_6837,N_6286);
nand U6987 (N_6987,N_6787,N_6441);
nand U6988 (N_6988,N_6569,N_6367);
xor U6989 (N_6989,N_6372,N_6633);
nor U6990 (N_6990,N_6595,N_6437);
nor U6991 (N_6991,N_6312,N_6834);
or U6992 (N_6992,N_6793,N_6483);
nand U6993 (N_6993,N_6848,N_6408);
nor U6994 (N_6994,N_6753,N_6632);
xnor U6995 (N_6995,N_6684,N_6409);
nor U6996 (N_6996,N_6268,N_6846);
xor U6997 (N_6997,N_6283,N_6365);
xor U6998 (N_6998,N_6505,N_6466);
xor U6999 (N_6999,N_6396,N_6747);
nand U7000 (N_7000,N_6331,N_6698);
and U7001 (N_7001,N_6647,N_6363);
xor U7002 (N_7002,N_6418,N_6428);
nand U7003 (N_7003,N_6501,N_6527);
nor U7004 (N_7004,N_6781,N_6605);
nor U7005 (N_7005,N_6706,N_6493);
xor U7006 (N_7006,N_6658,N_6406);
nand U7007 (N_7007,N_6533,N_6297);
nor U7008 (N_7008,N_6725,N_6489);
or U7009 (N_7009,N_6732,N_6598);
nor U7010 (N_7010,N_6807,N_6575);
and U7011 (N_7011,N_6513,N_6580);
xnor U7012 (N_7012,N_6335,N_6551);
xnor U7013 (N_7013,N_6609,N_6636);
nor U7014 (N_7014,N_6713,N_6435);
and U7015 (N_7015,N_6664,N_6669);
or U7016 (N_7016,N_6457,N_6344);
nand U7017 (N_7017,N_6332,N_6261);
and U7018 (N_7018,N_6587,N_6506);
xnor U7019 (N_7019,N_6674,N_6720);
xor U7020 (N_7020,N_6864,N_6641);
and U7021 (N_7021,N_6688,N_6517);
xnor U7022 (N_7022,N_6549,N_6357);
and U7023 (N_7023,N_6534,N_6608);
or U7024 (N_7024,N_6558,N_6308);
nor U7025 (N_7025,N_6739,N_6338);
xor U7026 (N_7026,N_6343,N_6640);
nor U7027 (N_7027,N_6858,N_6810);
or U7028 (N_7028,N_6284,N_6310);
nor U7029 (N_7029,N_6855,N_6453);
or U7030 (N_7030,N_6523,N_6324);
nand U7031 (N_7031,N_6368,N_6403);
nand U7032 (N_7032,N_6499,N_6784);
or U7033 (N_7033,N_6431,N_6497);
or U7034 (N_7034,N_6371,N_6594);
and U7035 (N_7035,N_6785,N_6340);
or U7036 (N_7036,N_6488,N_6507);
xnor U7037 (N_7037,N_6278,N_6836);
nor U7038 (N_7038,N_6572,N_6701);
and U7039 (N_7039,N_6603,N_6559);
and U7040 (N_7040,N_6410,N_6671);
and U7041 (N_7041,N_6322,N_6321);
nor U7042 (N_7042,N_6279,N_6516);
or U7043 (N_7043,N_6472,N_6574);
and U7044 (N_7044,N_6779,N_6514);
nand U7045 (N_7045,N_6473,N_6397);
nand U7046 (N_7046,N_6768,N_6576);
nand U7047 (N_7047,N_6285,N_6550);
xnor U7048 (N_7048,N_6526,N_6426);
nand U7049 (N_7049,N_6478,N_6568);
nor U7050 (N_7050,N_6306,N_6856);
nor U7051 (N_7051,N_6319,N_6623);
nor U7052 (N_7052,N_6370,N_6567);
or U7053 (N_7053,N_6522,N_6539);
or U7054 (N_7054,N_6430,N_6643);
or U7055 (N_7055,N_6347,N_6870);
and U7056 (N_7056,N_6873,N_6819);
xnor U7057 (N_7057,N_6543,N_6264);
or U7058 (N_7058,N_6528,N_6414);
xnor U7059 (N_7059,N_6795,N_6524);
nor U7060 (N_7060,N_6697,N_6346);
nand U7061 (N_7061,N_6510,N_6841);
and U7062 (N_7062,N_6400,N_6705);
or U7063 (N_7063,N_6788,N_6749);
xnor U7064 (N_7064,N_6588,N_6740);
nand U7065 (N_7065,N_6601,N_6614);
nor U7066 (N_7066,N_6724,N_6799);
nor U7067 (N_7067,N_6530,N_6610);
nand U7068 (N_7068,N_6666,N_6389);
nand U7069 (N_7069,N_6828,N_6777);
and U7070 (N_7070,N_6692,N_6783);
nand U7071 (N_7071,N_6449,N_6667);
and U7072 (N_7072,N_6392,N_6460);
or U7073 (N_7073,N_6395,N_6766);
or U7074 (N_7074,N_6780,N_6683);
xnor U7075 (N_7075,N_6366,N_6540);
xor U7076 (N_7076,N_6861,N_6635);
nor U7077 (N_7077,N_6715,N_6717);
xor U7078 (N_7078,N_6774,N_6794);
or U7079 (N_7079,N_6604,N_6851);
xnor U7080 (N_7080,N_6742,N_6269);
xor U7081 (N_7081,N_6360,N_6498);
nor U7082 (N_7082,N_6591,N_6770);
nor U7083 (N_7083,N_6833,N_6294);
nand U7084 (N_7084,N_6654,N_6512);
and U7085 (N_7085,N_6802,N_6258);
nor U7086 (N_7086,N_6761,N_6280);
or U7087 (N_7087,N_6579,N_6617);
nor U7088 (N_7088,N_6265,N_6359);
nand U7089 (N_7089,N_6270,N_6612);
and U7090 (N_7090,N_6676,N_6494);
xor U7091 (N_7091,N_6348,N_6289);
nor U7092 (N_7092,N_6276,N_6471);
and U7093 (N_7093,N_6791,N_6383);
xnor U7094 (N_7094,N_6440,N_6256);
and U7095 (N_7095,N_6764,N_6821);
nor U7096 (N_7096,N_6707,N_6381);
nor U7097 (N_7097,N_6722,N_6503);
xor U7098 (N_7098,N_6847,N_6772);
and U7099 (N_7099,N_6377,N_6468);
and U7100 (N_7100,N_6519,N_6590);
nor U7101 (N_7101,N_6657,N_6511);
nand U7102 (N_7102,N_6703,N_6845);
or U7103 (N_7103,N_6538,N_6274);
and U7104 (N_7104,N_6401,N_6482);
nor U7105 (N_7105,N_6464,N_6422);
or U7106 (N_7106,N_6546,N_6266);
nand U7107 (N_7107,N_6760,N_6718);
nor U7108 (N_7108,N_6743,N_6423);
or U7109 (N_7109,N_6767,N_6508);
or U7110 (N_7110,N_6320,N_6271);
nor U7111 (N_7111,N_6629,N_6689);
and U7112 (N_7112,N_6631,N_6515);
xor U7113 (N_7113,N_6818,N_6311);
xnor U7114 (N_7114,N_6376,N_6465);
nand U7115 (N_7115,N_6656,N_6812);
nor U7116 (N_7116,N_6811,N_6803);
or U7117 (N_7117,N_6459,N_6521);
xnor U7118 (N_7118,N_6552,N_6292);
nand U7119 (N_7119,N_6801,N_6295);
and U7120 (N_7120,N_6827,N_6504);
and U7121 (N_7121,N_6796,N_6782);
and U7122 (N_7122,N_6642,N_6872);
or U7123 (N_7123,N_6544,N_6329);
nor U7124 (N_7124,N_6650,N_6424);
nand U7125 (N_7125,N_6438,N_6691);
nand U7126 (N_7126,N_6751,N_6721);
and U7127 (N_7127,N_6333,N_6571);
or U7128 (N_7128,N_6387,N_6805);
nand U7129 (N_7129,N_6700,N_6334);
nor U7130 (N_7130,N_6628,N_6809);
and U7131 (N_7131,N_6736,N_6822);
nand U7132 (N_7132,N_6419,N_6581);
nand U7133 (N_7133,N_6687,N_6405);
nand U7134 (N_7134,N_6585,N_6433);
nand U7135 (N_7135,N_6492,N_6354);
nand U7136 (N_7136,N_6593,N_6393);
and U7137 (N_7137,N_6384,N_6813);
or U7138 (N_7138,N_6710,N_6411);
and U7139 (N_7139,N_6520,N_6531);
nor U7140 (N_7140,N_6620,N_6496);
or U7141 (N_7141,N_6823,N_6597);
and U7142 (N_7142,N_6733,N_6304);
nor U7143 (N_7143,N_6839,N_6445);
xnor U7144 (N_7144,N_6485,N_6273);
xnor U7145 (N_7145,N_6757,N_6762);
or U7146 (N_7146,N_6655,N_6618);
xor U7147 (N_7147,N_6871,N_6646);
nor U7148 (N_7148,N_6679,N_6356);
or U7149 (N_7149,N_6302,N_6615);
xor U7150 (N_7150,N_6630,N_6339);
and U7151 (N_7151,N_6458,N_6542);
and U7152 (N_7152,N_6625,N_6622);
or U7153 (N_7153,N_6364,N_6853);
or U7154 (N_7154,N_6352,N_6619);
or U7155 (N_7155,N_6446,N_6328);
xnor U7156 (N_7156,N_6442,N_6663);
nor U7157 (N_7157,N_6816,N_6849);
nand U7158 (N_7158,N_6860,N_6755);
or U7159 (N_7159,N_6432,N_6634);
xnor U7160 (N_7160,N_6681,N_6556);
and U7161 (N_7161,N_6358,N_6653);
xor U7162 (N_7162,N_6452,N_6866);
and U7163 (N_7163,N_6566,N_6626);
and U7164 (N_7164,N_6758,N_6479);
nand U7165 (N_7165,N_6480,N_6868);
nand U7166 (N_7166,N_6463,N_6379);
nand U7167 (N_7167,N_6824,N_6502);
xnor U7168 (N_7168,N_6391,N_6577);
nor U7169 (N_7169,N_6561,N_6272);
xor U7170 (N_7170,N_6644,N_6752);
nor U7171 (N_7171,N_6592,N_6775);
xnor U7172 (N_7172,N_6323,N_6599);
nor U7173 (N_7173,N_6573,N_6735);
nor U7174 (N_7174,N_6535,N_6448);
or U7175 (N_7175,N_6804,N_6798);
and U7176 (N_7176,N_6477,N_6296);
or U7177 (N_7177,N_6814,N_6299);
xnor U7178 (N_7178,N_6786,N_6613);
nor U7179 (N_7179,N_6685,N_6545);
and U7180 (N_7180,N_6652,N_6602);
and U7181 (N_7181,N_6481,N_6627);
xor U7182 (N_7182,N_6661,N_6399);
nand U7183 (N_7183,N_6750,N_6316);
nor U7184 (N_7184,N_6388,N_6820);
xor U7185 (N_7185,N_6287,N_6378);
xnor U7186 (N_7186,N_6421,N_6769);
nand U7187 (N_7187,N_6495,N_6472);
nor U7188 (N_7188,N_6841,N_6817);
and U7189 (N_7189,N_6859,N_6856);
and U7190 (N_7190,N_6257,N_6418);
nor U7191 (N_7191,N_6431,N_6572);
and U7192 (N_7192,N_6706,N_6345);
xor U7193 (N_7193,N_6806,N_6765);
and U7194 (N_7194,N_6445,N_6651);
nor U7195 (N_7195,N_6460,N_6828);
nor U7196 (N_7196,N_6513,N_6678);
or U7197 (N_7197,N_6681,N_6317);
nor U7198 (N_7198,N_6492,N_6819);
nor U7199 (N_7199,N_6563,N_6724);
xor U7200 (N_7200,N_6256,N_6710);
nand U7201 (N_7201,N_6529,N_6311);
and U7202 (N_7202,N_6643,N_6633);
xnor U7203 (N_7203,N_6573,N_6341);
and U7204 (N_7204,N_6824,N_6456);
or U7205 (N_7205,N_6364,N_6780);
and U7206 (N_7206,N_6694,N_6691);
nand U7207 (N_7207,N_6730,N_6812);
xor U7208 (N_7208,N_6439,N_6638);
nand U7209 (N_7209,N_6548,N_6494);
xnor U7210 (N_7210,N_6363,N_6850);
or U7211 (N_7211,N_6712,N_6292);
nand U7212 (N_7212,N_6592,N_6426);
or U7213 (N_7213,N_6346,N_6562);
xor U7214 (N_7214,N_6827,N_6351);
nor U7215 (N_7215,N_6846,N_6415);
nor U7216 (N_7216,N_6694,N_6700);
nand U7217 (N_7217,N_6681,N_6780);
xnor U7218 (N_7218,N_6587,N_6797);
or U7219 (N_7219,N_6384,N_6606);
and U7220 (N_7220,N_6586,N_6459);
xor U7221 (N_7221,N_6696,N_6727);
and U7222 (N_7222,N_6453,N_6397);
and U7223 (N_7223,N_6345,N_6864);
or U7224 (N_7224,N_6382,N_6522);
or U7225 (N_7225,N_6582,N_6770);
and U7226 (N_7226,N_6349,N_6367);
or U7227 (N_7227,N_6389,N_6430);
nand U7228 (N_7228,N_6786,N_6865);
nand U7229 (N_7229,N_6570,N_6385);
nor U7230 (N_7230,N_6416,N_6782);
xnor U7231 (N_7231,N_6462,N_6802);
or U7232 (N_7232,N_6384,N_6427);
or U7233 (N_7233,N_6863,N_6803);
nand U7234 (N_7234,N_6690,N_6383);
or U7235 (N_7235,N_6272,N_6749);
xor U7236 (N_7236,N_6418,N_6545);
and U7237 (N_7237,N_6843,N_6477);
or U7238 (N_7238,N_6800,N_6295);
or U7239 (N_7239,N_6642,N_6727);
xor U7240 (N_7240,N_6418,N_6836);
nand U7241 (N_7241,N_6650,N_6438);
or U7242 (N_7242,N_6709,N_6398);
nand U7243 (N_7243,N_6653,N_6784);
and U7244 (N_7244,N_6727,N_6466);
or U7245 (N_7245,N_6725,N_6637);
nand U7246 (N_7246,N_6523,N_6693);
nor U7247 (N_7247,N_6514,N_6664);
or U7248 (N_7248,N_6839,N_6256);
nand U7249 (N_7249,N_6257,N_6500);
or U7250 (N_7250,N_6614,N_6480);
and U7251 (N_7251,N_6276,N_6529);
or U7252 (N_7252,N_6256,N_6754);
nor U7253 (N_7253,N_6825,N_6527);
nor U7254 (N_7254,N_6722,N_6758);
xnor U7255 (N_7255,N_6781,N_6448);
nand U7256 (N_7256,N_6565,N_6674);
and U7257 (N_7257,N_6629,N_6301);
or U7258 (N_7258,N_6672,N_6304);
and U7259 (N_7259,N_6844,N_6765);
xnor U7260 (N_7260,N_6414,N_6372);
nand U7261 (N_7261,N_6725,N_6764);
xnor U7262 (N_7262,N_6722,N_6732);
xor U7263 (N_7263,N_6348,N_6442);
nand U7264 (N_7264,N_6596,N_6502);
nor U7265 (N_7265,N_6570,N_6336);
nand U7266 (N_7266,N_6588,N_6702);
or U7267 (N_7267,N_6778,N_6762);
and U7268 (N_7268,N_6395,N_6872);
or U7269 (N_7269,N_6437,N_6602);
nand U7270 (N_7270,N_6870,N_6793);
nor U7271 (N_7271,N_6517,N_6850);
xnor U7272 (N_7272,N_6274,N_6770);
xor U7273 (N_7273,N_6660,N_6646);
nor U7274 (N_7274,N_6258,N_6642);
xnor U7275 (N_7275,N_6268,N_6488);
xor U7276 (N_7276,N_6496,N_6462);
xor U7277 (N_7277,N_6800,N_6780);
xor U7278 (N_7278,N_6491,N_6709);
nand U7279 (N_7279,N_6660,N_6554);
nor U7280 (N_7280,N_6389,N_6669);
and U7281 (N_7281,N_6480,N_6401);
xnor U7282 (N_7282,N_6691,N_6399);
nor U7283 (N_7283,N_6777,N_6506);
or U7284 (N_7284,N_6863,N_6725);
or U7285 (N_7285,N_6757,N_6626);
xor U7286 (N_7286,N_6614,N_6694);
and U7287 (N_7287,N_6464,N_6543);
or U7288 (N_7288,N_6600,N_6792);
nor U7289 (N_7289,N_6813,N_6690);
nand U7290 (N_7290,N_6747,N_6675);
nor U7291 (N_7291,N_6494,N_6486);
or U7292 (N_7292,N_6473,N_6482);
nand U7293 (N_7293,N_6750,N_6848);
xnor U7294 (N_7294,N_6464,N_6663);
or U7295 (N_7295,N_6774,N_6702);
or U7296 (N_7296,N_6803,N_6693);
and U7297 (N_7297,N_6326,N_6468);
or U7298 (N_7298,N_6703,N_6594);
and U7299 (N_7299,N_6668,N_6654);
nand U7300 (N_7300,N_6621,N_6709);
and U7301 (N_7301,N_6552,N_6505);
or U7302 (N_7302,N_6854,N_6275);
and U7303 (N_7303,N_6738,N_6391);
and U7304 (N_7304,N_6760,N_6723);
xor U7305 (N_7305,N_6715,N_6839);
nand U7306 (N_7306,N_6788,N_6815);
nor U7307 (N_7307,N_6416,N_6251);
nand U7308 (N_7308,N_6418,N_6827);
nand U7309 (N_7309,N_6629,N_6270);
nand U7310 (N_7310,N_6639,N_6744);
nor U7311 (N_7311,N_6455,N_6808);
nor U7312 (N_7312,N_6679,N_6683);
xnor U7313 (N_7313,N_6271,N_6442);
nor U7314 (N_7314,N_6855,N_6739);
or U7315 (N_7315,N_6431,N_6765);
nor U7316 (N_7316,N_6577,N_6851);
nor U7317 (N_7317,N_6661,N_6826);
and U7318 (N_7318,N_6664,N_6334);
and U7319 (N_7319,N_6522,N_6793);
xor U7320 (N_7320,N_6362,N_6513);
and U7321 (N_7321,N_6631,N_6355);
and U7322 (N_7322,N_6483,N_6563);
nor U7323 (N_7323,N_6603,N_6726);
and U7324 (N_7324,N_6622,N_6260);
xnor U7325 (N_7325,N_6382,N_6443);
xor U7326 (N_7326,N_6866,N_6782);
nor U7327 (N_7327,N_6802,N_6627);
xnor U7328 (N_7328,N_6613,N_6508);
xor U7329 (N_7329,N_6392,N_6566);
xor U7330 (N_7330,N_6404,N_6309);
and U7331 (N_7331,N_6273,N_6537);
and U7332 (N_7332,N_6362,N_6308);
nor U7333 (N_7333,N_6559,N_6493);
or U7334 (N_7334,N_6576,N_6860);
xor U7335 (N_7335,N_6298,N_6431);
nand U7336 (N_7336,N_6862,N_6538);
nor U7337 (N_7337,N_6669,N_6386);
nor U7338 (N_7338,N_6494,N_6401);
nand U7339 (N_7339,N_6621,N_6484);
xor U7340 (N_7340,N_6822,N_6701);
and U7341 (N_7341,N_6828,N_6826);
or U7342 (N_7342,N_6738,N_6766);
xnor U7343 (N_7343,N_6669,N_6568);
or U7344 (N_7344,N_6256,N_6685);
nor U7345 (N_7345,N_6260,N_6447);
xnor U7346 (N_7346,N_6391,N_6815);
xnor U7347 (N_7347,N_6609,N_6312);
or U7348 (N_7348,N_6274,N_6699);
xnor U7349 (N_7349,N_6273,N_6867);
xor U7350 (N_7350,N_6469,N_6646);
or U7351 (N_7351,N_6561,N_6254);
and U7352 (N_7352,N_6784,N_6645);
xor U7353 (N_7353,N_6407,N_6563);
xnor U7354 (N_7354,N_6346,N_6731);
xnor U7355 (N_7355,N_6539,N_6717);
nand U7356 (N_7356,N_6790,N_6649);
nand U7357 (N_7357,N_6871,N_6723);
xor U7358 (N_7358,N_6795,N_6310);
xor U7359 (N_7359,N_6563,N_6496);
and U7360 (N_7360,N_6642,N_6719);
xnor U7361 (N_7361,N_6259,N_6554);
nor U7362 (N_7362,N_6849,N_6740);
xnor U7363 (N_7363,N_6672,N_6355);
or U7364 (N_7364,N_6418,N_6282);
xnor U7365 (N_7365,N_6314,N_6786);
nand U7366 (N_7366,N_6709,N_6644);
and U7367 (N_7367,N_6276,N_6472);
xor U7368 (N_7368,N_6507,N_6426);
xor U7369 (N_7369,N_6855,N_6460);
xnor U7370 (N_7370,N_6426,N_6614);
or U7371 (N_7371,N_6325,N_6403);
nand U7372 (N_7372,N_6576,N_6529);
nor U7373 (N_7373,N_6384,N_6790);
nor U7374 (N_7374,N_6409,N_6449);
nor U7375 (N_7375,N_6448,N_6872);
nand U7376 (N_7376,N_6311,N_6369);
nand U7377 (N_7377,N_6752,N_6510);
and U7378 (N_7378,N_6375,N_6855);
or U7379 (N_7379,N_6672,N_6767);
nand U7380 (N_7380,N_6372,N_6736);
and U7381 (N_7381,N_6307,N_6337);
nor U7382 (N_7382,N_6337,N_6440);
and U7383 (N_7383,N_6276,N_6360);
and U7384 (N_7384,N_6421,N_6277);
nand U7385 (N_7385,N_6572,N_6292);
or U7386 (N_7386,N_6442,N_6320);
nor U7387 (N_7387,N_6548,N_6314);
xor U7388 (N_7388,N_6346,N_6743);
xor U7389 (N_7389,N_6786,N_6611);
and U7390 (N_7390,N_6509,N_6786);
nor U7391 (N_7391,N_6789,N_6480);
or U7392 (N_7392,N_6626,N_6516);
and U7393 (N_7393,N_6847,N_6431);
nor U7394 (N_7394,N_6524,N_6638);
and U7395 (N_7395,N_6448,N_6444);
nor U7396 (N_7396,N_6652,N_6864);
nand U7397 (N_7397,N_6533,N_6818);
or U7398 (N_7398,N_6807,N_6775);
nand U7399 (N_7399,N_6437,N_6279);
or U7400 (N_7400,N_6344,N_6412);
nor U7401 (N_7401,N_6566,N_6364);
xor U7402 (N_7402,N_6816,N_6350);
and U7403 (N_7403,N_6763,N_6259);
xnor U7404 (N_7404,N_6555,N_6342);
nor U7405 (N_7405,N_6431,N_6265);
nor U7406 (N_7406,N_6626,N_6560);
nand U7407 (N_7407,N_6455,N_6768);
xor U7408 (N_7408,N_6494,N_6354);
nor U7409 (N_7409,N_6330,N_6299);
xnor U7410 (N_7410,N_6565,N_6722);
xor U7411 (N_7411,N_6492,N_6790);
nand U7412 (N_7412,N_6723,N_6646);
nand U7413 (N_7413,N_6590,N_6794);
nor U7414 (N_7414,N_6543,N_6654);
or U7415 (N_7415,N_6708,N_6711);
nor U7416 (N_7416,N_6732,N_6300);
or U7417 (N_7417,N_6734,N_6574);
xnor U7418 (N_7418,N_6736,N_6267);
xnor U7419 (N_7419,N_6251,N_6460);
nand U7420 (N_7420,N_6509,N_6363);
or U7421 (N_7421,N_6256,N_6520);
and U7422 (N_7422,N_6287,N_6435);
or U7423 (N_7423,N_6261,N_6768);
nor U7424 (N_7424,N_6498,N_6331);
xnor U7425 (N_7425,N_6261,N_6635);
or U7426 (N_7426,N_6585,N_6272);
nor U7427 (N_7427,N_6798,N_6688);
and U7428 (N_7428,N_6757,N_6383);
nor U7429 (N_7429,N_6458,N_6284);
and U7430 (N_7430,N_6675,N_6365);
nand U7431 (N_7431,N_6697,N_6632);
nor U7432 (N_7432,N_6446,N_6749);
nor U7433 (N_7433,N_6852,N_6563);
nor U7434 (N_7434,N_6730,N_6726);
and U7435 (N_7435,N_6539,N_6643);
or U7436 (N_7436,N_6454,N_6268);
xor U7437 (N_7437,N_6653,N_6379);
nand U7438 (N_7438,N_6362,N_6314);
or U7439 (N_7439,N_6460,N_6532);
or U7440 (N_7440,N_6272,N_6354);
nor U7441 (N_7441,N_6507,N_6803);
or U7442 (N_7442,N_6517,N_6819);
and U7443 (N_7443,N_6521,N_6604);
xnor U7444 (N_7444,N_6381,N_6709);
and U7445 (N_7445,N_6283,N_6705);
xor U7446 (N_7446,N_6598,N_6435);
or U7447 (N_7447,N_6774,N_6573);
and U7448 (N_7448,N_6370,N_6346);
and U7449 (N_7449,N_6747,N_6765);
xnor U7450 (N_7450,N_6840,N_6854);
or U7451 (N_7451,N_6403,N_6803);
and U7452 (N_7452,N_6839,N_6403);
xor U7453 (N_7453,N_6575,N_6322);
and U7454 (N_7454,N_6661,N_6816);
nand U7455 (N_7455,N_6652,N_6704);
or U7456 (N_7456,N_6381,N_6634);
and U7457 (N_7457,N_6403,N_6604);
nand U7458 (N_7458,N_6284,N_6684);
nand U7459 (N_7459,N_6434,N_6754);
or U7460 (N_7460,N_6376,N_6780);
nor U7461 (N_7461,N_6269,N_6514);
nand U7462 (N_7462,N_6502,N_6797);
xnor U7463 (N_7463,N_6706,N_6719);
nor U7464 (N_7464,N_6343,N_6805);
xnor U7465 (N_7465,N_6605,N_6525);
xnor U7466 (N_7466,N_6632,N_6628);
xnor U7467 (N_7467,N_6669,N_6384);
or U7468 (N_7468,N_6854,N_6314);
or U7469 (N_7469,N_6340,N_6478);
xor U7470 (N_7470,N_6278,N_6601);
nand U7471 (N_7471,N_6831,N_6606);
or U7472 (N_7472,N_6418,N_6566);
nor U7473 (N_7473,N_6597,N_6648);
nand U7474 (N_7474,N_6510,N_6284);
or U7475 (N_7475,N_6539,N_6793);
xor U7476 (N_7476,N_6621,N_6439);
xor U7477 (N_7477,N_6440,N_6524);
or U7478 (N_7478,N_6412,N_6313);
nand U7479 (N_7479,N_6661,N_6539);
nor U7480 (N_7480,N_6827,N_6789);
xnor U7481 (N_7481,N_6268,N_6736);
and U7482 (N_7482,N_6793,N_6318);
nand U7483 (N_7483,N_6462,N_6450);
nand U7484 (N_7484,N_6513,N_6568);
xor U7485 (N_7485,N_6448,N_6318);
nor U7486 (N_7486,N_6345,N_6511);
xor U7487 (N_7487,N_6468,N_6513);
or U7488 (N_7488,N_6601,N_6329);
or U7489 (N_7489,N_6508,N_6777);
nand U7490 (N_7490,N_6258,N_6333);
nor U7491 (N_7491,N_6441,N_6537);
and U7492 (N_7492,N_6502,N_6283);
nor U7493 (N_7493,N_6634,N_6594);
and U7494 (N_7494,N_6691,N_6797);
nand U7495 (N_7495,N_6467,N_6755);
nand U7496 (N_7496,N_6261,N_6352);
nor U7497 (N_7497,N_6298,N_6451);
nor U7498 (N_7498,N_6283,N_6690);
xnor U7499 (N_7499,N_6612,N_6545);
nand U7500 (N_7500,N_7390,N_6984);
and U7501 (N_7501,N_7454,N_7153);
and U7502 (N_7502,N_7415,N_7258);
nand U7503 (N_7503,N_7309,N_6941);
nand U7504 (N_7504,N_7354,N_7130);
nand U7505 (N_7505,N_7154,N_6998);
and U7506 (N_7506,N_6953,N_6895);
xor U7507 (N_7507,N_7393,N_6928);
or U7508 (N_7508,N_7324,N_7321);
xnor U7509 (N_7509,N_7001,N_7301);
or U7510 (N_7510,N_6948,N_7084);
nand U7511 (N_7511,N_7275,N_7072);
xnor U7512 (N_7512,N_7289,N_7155);
and U7513 (N_7513,N_7240,N_6892);
nor U7514 (N_7514,N_6996,N_7458);
xor U7515 (N_7515,N_7238,N_7210);
nor U7516 (N_7516,N_7299,N_7097);
or U7517 (N_7517,N_7171,N_7000);
and U7518 (N_7518,N_7316,N_7423);
nand U7519 (N_7519,N_7222,N_7022);
nand U7520 (N_7520,N_7284,N_7455);
and U7521 (N_7521,N_7392,N_7464);
nor U7522 (N_7522,N_7334,N_7091);
nor U7523 (N_7523,N_7055,N_7208);
or U7524 (N_7524,N_7217,N_7338);
nor U7525 (N_7525,N_7252,N_6964);
nor U7526 (N_7526,N_7361,N_7092);
nor U7527 (N_7527,N_6889,N_7119);
or U7528 (N_7528,N_7140,N_7305);
nor U7529 (N_7529,N_7215,N_7213);
nand U7530 (N_7530,N_7136,N_7133);
and U7531 (N_7531,N_7046,N_7068);
and U7532 (N_7532,N_6885,N_7282);
xor U7533 (N_7533,N_7152,N_6969);
nand U7534 (N_7534,N_7443,N_7486);
nand U7535 (N_7535,N_7247,N_7298);
nand U7536 (N_7536,N_7012,N_7164);
nor U7537 (N_7537,N_7228,N_6923);
and U7538 (N_7538,N_7048,N_7043);
and U7539 (N_7539,N_6902,N_6972);
or U7540 (N_7540,N_7452,N_6921);
xor U7541 (N_7541,N_6999,N_6992);
nand U7542 (N_7542,N_7403,N_7336);
and U7543 (N_7543,N_7015,N_7371);
or U7544 (N_7544,N_7113,N_7101);
or U7545 (N_7545,N_7404,N_6907);
xor U7546 (N_7546,N_7462,N_7008);
and U7547 (N_7547,N_7434,N_7420);
and U7548 (N_7548,N_7107,N_7399);
or U7549 (N_7549,N_7435,N_7329);
nor U7550 (N_7550,N_6922,N_7496);
nor U7551 (N_7551,N_6960,N_7003);
and U7552 (N_7552,N_6875,N_7168);
nor U7553 (N_7553,N_7019,N_7424);
nor U7554 (N_7554,N_7359,N_7187);
nand U7555 (N_7555,N_7366,N_7206);
xnor U7556 (N_7556,N_6990,N_6942);
and U7557 (N_7557,N_7492,N_7451);
or U7558 (N_7558,N_7069,N_7417);
nand U7559 (N_7559,N_7353,N_7388);
or U7560 (N_7560,N_7195,N_6956);
nand U7561 (N_7561,N_7202,N_6913);
or U7562 (N_7562,N_7378,N_6890);
nor U7563 (N_7563,N_7010,N_6888);
nor U7564 (N_7564,N_7478,N_7271);
nand U7565 (N_7565,N_6965,N_7088);
nor U7566 (N_7566,N_7445,N_7192);
nand U7567 (N_7567,N_7444,N_7216);
nand U7568 (N_7568,N_7108,N_7146);
nor U7569 (N_7569,N_7115,N_7065);
nor U7570 (N_7570,N_7332,N_7036);
nand U7571 (N_7571,N_7441,N_7469);
or U7572 (N_7572,N_7197,N_7315);
and U7573 (N_7573,N_6976,N_7158);
nand U7574 (N_7574,N_7314,N_7104);
nor U7575 (N_7575,N_7433,N_7277);
and U7576 (N_7576,N_6916,N_7006);
nand U7577 (N_7577,N_6877,N_7427);
or U7578 (N_7578,N_6982,N_7437);
nor U7579 (N_7579,N_7261,N_7472);
nor U7580 (N_7580,N_7077,N_7474);
xor U7581 (N_7581,N_6994,N_7291);
nor U7582 (N_7582,N_7049,N_6900);
or U7583 (N_7583,N_7053,N_7431);
and U7584 (N_7584,N_7027,N_7360);
xor U7585 (N_7585,N_7270,N_7457);
xnor U7586 (N_7586,N_7414,N_7093);
nor U7587 (N_7587,N_7259,N_6886);
nor U7588 (N_7588,N_7453,N_7031);
and U7589 (N_7589,N_7024,N_7058);
xor U7590 (N_7590,N_7145,N_7494);
or U7591 (N_7591,N_7290,N_7226);
nand U7592 (N_7592,N_7383,N_6950);
or U7593 (N_7593,N_7375,N_7147);
xor U7594 (N_7594,N_7304,N_7410);
or U7595 (N_7595,N_7167,N_6979);
and U7596 (N_7596,N_7173,N_7098);
or U7597 (N_7597,N_7177,N_7174);
nand U7598 (N_7598,N_7379,N_7308);
or U7599 (N_7599,N_7471,N_7243);
and U7600 (N_7600,N_6924,N_7060);
nand U7601 (N_7601,N_7142,N_7161);
nand U7602 (N_7602,N_7318,N_7491);
and U7603 (N_7603,N_7233,N_6936);
xor U7604 (N_7604,N_7447,N_6962);
or U7605 (N_7605,N_7402,N_7040);
nor U7606 (N_7606,N_7489,N_7026);
xnor U7607 (N_7607,N_7165,N_6893);
nor U7608 (N_7608,N_7263,N_7253);
and U7609 (N_7609,N_6935,N_7440);
or U7610 (N_7610,N_7179,N_7105);
or U7611 (N_7611,N_7112,N_7374);
nand U7612 (N_7612,N_7497,N_7418);
xnor U7613 (N_7613,N_6945,N_6878);
nand U7614 (N_7614,N_7183,N_7180);
or U7615 (N_7615,N_7313,N_7079);
nand U7616 (N_7616,N_7227,N_7351);
and U7617 (N_7617,N_7047,N_7481);
nor U7618 (N_7618,N_7285,N_7032);
and U7619 (N_7619,N_7062,N_7200);
nor U7620 (N_7620,N_6957,N_6989);
and U7621 (N_7621,N_7081,N_7400);
nand U7622 (N_7622,N_6967,N_7466);
nand U7623 (N_7623,N_7419,N_7335);
xnor U7624 (N_7624,N_6919,N_7122);
and U7625 (N_7625,N_7230,N_7312);
nor U7626 (N_7626,N_7051,N_6929);
or U7627 (N_7627,N_7016,N_7138);
and U7628 (N_7628,N_7170,N_6914);
or U7629 (N_7629,N_7302,N_7307);
xnor U7630 (N_7630,N_7248,N_7151);
nor U7631 (N_7631,N_7292,N_6934);
nor U7632 (N_7632,N_7386,N_6927);
xnor U7633 (N_7633,N_7245,N_7294);
and U7634 (N_7634,N_7368,N_7389);
xnor U7635 (N_7635,N_7413,N_6988);
nand U7636 (N_7636,N_7343,N_7094);
and U7637 (N_7637,N_7241,N_7459);
nand U7638 (N_7638,N_6983,N_7297);
nand U7639 (N_7639,N_7054,N_7340);
or U7640 (N_7640,N_7162,N_6966);
nand U7641 (N_7641,N_7257,N_7251);
xnor U7642 (N_7642,N_7196,N_6951);
or U7643 (N_7643,N_7114,N_6920);
nand U7644 (N_7644,N_6931,N_7063);
or U7645 (N_7645,N_7175,N_7057);
nand U7646 (N_7646,N_6944,N_7279);
and U7647 (N_7647,N_7235,N_7322);
nor U7648 (N_7648,N_7411,N_7163);
nand U7649 (N_7649,N_6970,N_7087);
or U7650 (N_7650,N_7030,N_7467);
xnor U7651 (N_7651,N_7405,N_6963);
nor U7652 (N_7652,N_7017,N_7021);
and U7653 (N_7653,N_7129,N_7320);
xor U7654 (N_7654,N_7028,N_6909);
or U7655 (N_7655,N_7463,N_7325);
or U7656 (N_7656,N_6955,N_7201);
or U7657 (N_7657,N_7218,N_6995);
xor U7658 (N_7658,N_6918,N_7004);
nor U7659 (N_7659,N_7239,N_7102);
xor U7660 (N_7660,N_7446,N_7380);
and U7661 (N_7661,N_7002,N_7267);
nand U7662 (N_7662,N_7190,N_7096);
or U7663 (N_7663,N_7412,N_7237);
nand U7664 (N_7664,N_6997,N_7225);
xor U7665 (N_7665,N_7337,N_7221);
xnor U7666 (N_7666,N_6932,N_7364);
or U7667 (N_7667,N_6958,N_7011);
xor U7668 (N_7668,N_7018,N_7448);
nor U7669 (N_7669,N_7439,N_7013);
xnor U7670 (N_7670,N_7328,N_6896);
nor U7671 (N_7671,N_7224,N_7281);
xnor U7672 (N_7672,N_7269,N_7181);
and U7673 (N_7673,N_6876,N_7369);
xnor U7674 (N_7674,N_7029,N_7042);
and U7675 (N_7675,N_7041,N_6991);
and U7676 (N_7676,N_7432,N_7385);
nor U7677 (N_7677,N_7266,N_7493);
or U7678 (N_7678,N_7387,N_6883);
xnor U7679 (N_7679,N_6943,N_7131);
or U7680 (N_7680,N_7296,N_7347);
or U7681 (N_7681,N_7121,N_6973);
xor U7682 (N_7682,N_7203,N_7265);
nor U7683 (N_7683,N_7367,N_7166);
and U7684 (N_7684,N_7214,N_6949);
nand U7685 (N_7685,N_7341,N_7134);
and U7686 (N_7686,N_7144,N_7480);
or U7687 (N_7687,N_6894,N_7118);
xor U7688 (N_7688,N_6975,N_7186);
or U7689 (N_7689,N_7193,N_7487);
nand U7690 (N_7690,N_7274,N_6980);
nor U7691 (N_7691,N_6985,N_7288);
nand U7692 (N_7692,N_6933,N_6961);
xor U7693 (N_7693,N_7460,N_6939);
nand U7694 (N_7694,N_7485,N_6915);
xnor U7695 (N_7695,N_7059,N_7473);
nor U7696 (N_7696,N_7124,N_7303);
nand U7697 (N_7697,N_6925,N_6905);
nand U7698 (N_7698,N_7377,N_7199);
xor U7699 (N_7699,N_7276,N_6959);
xnor U7700 (N_7700,N_7346,N_7137);
nor U7701 (N_7701,N_7488,N_7363);
and U7702 (N_7702,N_7039,N_6930);
and U7703 (N_7703,N_7306,N_6903);
nand U7704 (N_7704,N_7135,N_7095);
nor U7705 (N_7705,N_7132,N_6917);
nand U7706 (N_7706,N_7490,N_7149);
or U7707 (N_7707,N_7421,N_7005);
xor U7708 (N_7708,N_7468,N_7075);
nand U7709 (N_7709,N_6897,N_7067);
nand U7710 (N_7710,N_7429,N_7212);
nand U7711 (N_7711,N_7050,N_6879);
and U7712 (N_7712,N_7461,N_7436);
nand U7713 (N_7713,N_7172,N_7176);
nand U7714 (N_7714,N_6881,N_6968);
and U7715 (N_7715,N_7260,N_7220);
or U7716 (N_7716,N_7278,N_7256);
nand U7717 (N_7717,N_7345,N_7449);
nand U7718 (N_7718,N_7319,N_7381);
or U7719 (N_7719,N_7475,N_7300);
or U7720 (N_7720,N_6940,N_7085);
nand U7721 (N_7721,N_7188,N_7409);
xor U7722 (N_7722,N_7264,N_7159);
nand U7723 (N_7723,N_7401,N_7358);
xnor U7724 (N_7724,N_7272,N_7074);
and U7725 (N_7725,N_6911,N_7242);
nor U7726 (N_7726,N_7357,N_7089);
xor U7727 (N_7727,N_7110,N_7407);
xnor U7728 (N_7728,N_7109,N_7406);
nor U7729 (N_7729,N_7355,N_7352);
nand U7730 (N_7730,N_7373,N_7090);
xor U7731 (N_7731,N_7106,N_7372);
nor U7732 (N_7732,N_7244,N_6971);
nand U7733 (N_7733,N_7430,N_6946);
nor U7734 (N_7734,N_7020,N_6901);
nand U7735 (N_7735,N_7045,N_7076);
nand U7736 (N_7736,N_6891,N_6993);
nand U7737 (N_7737,N_7185,N_7232);
or U7738 (N_7738,N_7083,N_7139);
nand U7739 (N_7739,N_7157,N_7370);
or U7740 (N_7740,N_7333,N_6986);
nand U7741 (N_7741,N_7293,N_7295);
or U7742 (N_7742,N_7397,N_7426);
nand U7743 (N_7743,N_6947,N_7127);
nor U7744 (N_7744,N_7111,N_6987);
or U7745 (N_7745,N_7498,N_7184);
and U7746 (N_7746,N_7323,N_7178);
and U7747 (N_7747,N_7116,N_7204);
xor U7748 (N_7748,N_6898,N_7254);
nor U7749 (N_7749,N_7014,N_7191);
and U7750 (N_7750,N_7160,N_7391);
nor U7751 (N_7751,N_7327,N_7484);
or U7752 (N_7752,N_6904,N_7025);
xnor U7753 (N_7753,N_7156,N_7255);
nor U7754 (N_7754,N_6977,N_7007);
nand U7755 (N_7755,N_7100,N_6912);
or U7756 (N_7756,N_7465,N_7342);
nor U7757 (N_7757,N_7348,N_7317);
xor U7758 (N_7758,N_7148,N_7286);
or U7759 (N_7759,N_7408,N_7066);
and U7760 (N_7760,N_7384,N_6882);
nor U7761 (N_7761,N_7273,N_7056);
and U7762 (N_7762,N_7223,N_7416);
nor U7763 (N_7763,N_7125,N_7219);
and U7764 (N_7764,N_7169,N_7250);
or U7765 (N_7765,N_6910,N_7428);
and U7766 (N_7766,N_7395,N_7143);
nand U7767 (N_7767,N_7234,N_6974);
xnor U7768 (N_7768,N_7086,N_7376);
nand U7769 (N_7769,N_7052,N_7120);
xor U7770 (N_7770,N_7209,N_7495);
and U7771 (N_7771,N_7339,N_7229);
nor U7772 (N_7772,N_7438,N_7311);
nor U7773 (N_7773,N_6954,N_7398);
and U7774 (N_7774,N_7205,N_6899);
xor U7775 (N_7775,N_7365,N_7080);
nand U7776 (N_7776,N_7073,N_7326);
nor U7777 (N_7777,N_7362,N_7350);
xnor U7778 (N_7778,N_6978,N_7044);
xor U7779 (N_7779,N_7396,N_7470);
xnor U7780 (N_7780,N_6938,N_7211);
xnor U7781 (N_7781,N_6937,N_7123);
nand U7782 (N_7782,N_7349,N_7128);
nand U7783 (N_7783,N_7287,N_7182);
and U7784 (N_7784,N_6884,N_7422);
xnor U7785 (N_7785,N_7482,N_7033);
xor U7786 (N_7786,N_6908,N_7023);
nor U7787 (N_7787,N_7061,N_7207);
nand U7788 (N_7788,N_7310,N_6926);
and U7789 (N_7789,N_7194,N_7009);
nand U7790 (N_7790,N_7231,N_7456);
or U7791 (N_7791,N_7064,N_7126);
and U7792 (N_7792,N_7483,N_7479);
or U7793 (N_7793,N_7070,N_7268);
and U7794 (N_7794,N_7331,N_7477);
xnor U7795 (N_7795,N_7082,N_7150);
nor U7796 (N_7796,N_7280,N_7356);
xor U7797 (N_7797,N_6880,N_6981);
or U7798 (N_7798,N_6952,N_7189);
xor U7799 (N_7799,N_7249,N_7103);
and U7800 (N_7800,N_7198,N_7330);
or U7801 (N_7801,N_6906,N_7071);
or U7802 (N_7802,N_7283,N_7262);
and U7803 (N_7803,N_7035,N_7034);
nand U7804 (N_7804,N_7394,N_7141);
xor U7805 (N_7805,N_7037,N_7450);
nor U7806 (N_7806,N_7499,N_7246);
nand U7807 (N_7807,N_7344,N_7117);
nand U7808 (N_7808,N_7236,N_7038);
xnor U7809 (N_7809,N_6887,N_7442);
and U7810 (N_7810,N_7425,N_7382);
nor U7811 (N_7811,N_7078,N_7099);
nor U7812 (N_7812,N_7476,N_6931);
and U7813 (N_7813,N_7053,N_7442);
nor U7814 (N_7814,N_6896,N_7338);
or U7815 (N_7815,N_6932,N_7424);
nand U7816 (N_7816,N_7164,N_7034);
xnor U7817 (N_7817,N_7315,N_7303);
and U7818 (N_7818,N_7291,N_7008);
or U7819 (N_7819,N_7355,N_7244);
and U7820 (N_7820,N_7426,N_7362);
nor U7821 (N_7821,N_7441,N_7162);
nor U7822 (N_7822,N_7288,N_6961);
nor U7823 (N_7823,N_7070,N_7446);
xnor U7824 (N_7824,N_7198,N_6924);
and U7825 (N_7825,N_7316,N_7012);
and U7826 (N_7826,N_6974,N_7390);
and U7827 (N_7827,N_7266,N_6968);
nand U7828 (N_7828,N_7261,N_7382);
or U7829 (N_7829,N_7419,N_7476);
nand U7830 (N_7830,N_7348,N_7112);
nor U7831 (N_7831,N_7369,N_7078);
nor U7832 (N_7832,N_6929,N_7427);
nand U7833 (N_7833,N_7059,N_7346);
or U7834 (N_7834,N_7184,N_7230);
nand U7835 (N_7835,N_7487,N_7384);
nor U7836 (N_7836,N_7167,N_7299);
nand U7837 (N_7837,N_7499,N_7337);
nor U7838 (N_7838,N_7408,N_7175);
xor U7839 (N_7839,N_6886,N_7131);
nor U7840 (N_7840,N_7425,N_7336);
or U7841 (N_7841,N_7274,N_6984);
xnor U7842 (N_7842,N_7084,N_7271);
and U7843 (N_7843,N_6884,N_7305);
nand U7844 (N_7844,N_7267,N_6932);
nor U7845 (N_7845,N_7465,N_7012);
xnor U7846 (N_7846,N_7463,N_7452);
nor U7847 (N_7847,N_6900,N_7067);
nand U7848 (N_7848,N_7458,N_7431);
nand U7849 (N_7849,N_7290,N_7179);
xnor U7850 (N_7850,N_6936,N_7210);
or U7851 (N_7851,N_7148,N_7060);
and U7852 (N_7852,N_7324,N_7192);
xor U7853 (N_7853,N_7364,N_7306);
xnor U7854 (N_7854,N_7377,N_7072);
xnor U7855 (N_7855,N_7164,N_7395);
nor U7856 (N_7856,N_7189,N_7060);
and U7857 (N_7857,N_6928,N_7132);
or U7858 (N_7858,N_6893,N_7247);
nand U7859 (N_7859,N_7153,N_7374);
and U7860 (N_7860,N_7369,N_6968);
or U7861 (N_7861,N_7294,N_7452);
nor U7862 (N_7862,N_6951,N_7212);
or U7863 (N_7863,N_7490,N_7342);
nor U7864 (N_7864,N_6989,N_7090);
nor U7865 (N_7865,N_6988,N_7287);
xor U7866 (N_7866,N_7013,N_6941);
and U7867 (N_7867,N_7096,N_7434);
xor U7868 (N_7868,N_7468,N_7195);
or U7869 (N_7869,N_7254,N_7299);
nor U7870 (N_7870,N_6964,N_7203);
or U7871 (N_7871,N_7341,N_7333);
xor U7872 (N_7872,N_7216,N_7012);
and U7873 (N_7873,N_7324,N_7401);
nor U7874 (N_7874,N_7146,N_6963);
and U7875 (N_7875,N_6954,N_7026);
xnor U7876 (N_7876,N_7359,N_6984);
and U7877 (N_7877,N_6932,N_7276);
or U7878 (N_7878,N_7080,N_7177);
nand U7879 (N_7879,N_6945,N_6919);
nand U7880 (N_7880,N_7494,N_7439);
and U7881 (N_7881,N_6988,N_7461);
xor U7882 (N_7882,N_7054,N_7472);
or U7883 (N_7883,N_7436,N_7022);
nor U7884 (N_7884,N_7204,N_7469);
xor U7885 (N_7885,N_7364,N_7085);
and U7886 (N_7886,N_7074,N_7327);
and U7887 (N_7887,N_7027,N_7320);
and U7888 (N_7888,N_7192,N_7012);
nand U7889 (N_7889,N_7329,N_7342);
xnor U7890 (N_7890,N_7166,N_7342);
and U7891 (N_7891,N_7467,N_7332);
nor U7892 (N_7892,N_7430,N_7024);
nand U7893 (N_7893,N_7068,N_6975);
and U7894 (N_7894,N_7043,N_7450);
xor U7895 (N_7895,N_7354,N_6965);
nor U7896 (N_7896,N_6938,N_7349);
xnor U7897 (N_7897,N_7119,N_7480);
xnor U7898 (N_7898,N_7153,N_7458);
xnor U7899 (N_7899,N_7332,N_7374);
or U7900 (N_7900,N_6915,N_6963);
nor U7901 (N_7901,N_7271,N_7034);
and U7902 (N_7902,N_7490,N_7202);
and U7903 (N_7903,N_7008,N_7385);
and U7904 (N_7904,N_7087,N_7222);
nor U7905 (N_7905,N_7364,N_6976);
or U7906 (N_7906,N_7319,N_7146);
or U7907 (N_7907,N_7342,N_7324);
nand U7908 (N_7908,N_7263,N_6885);
xnor U7909 (N_7909,N_6906,N_7140);
and U7910 (N_7910,N_7065,N_7184);
nor U7911 (N_7911,N_7050,N_6881);
or U7912 (N_7912,N_7196,N_7186);
nand U7913 (N_7913,N_7469,N_6931);
or U7914 (N_7914,N_7175,N_7297);
nand U7915 (N_7915,N_7014,N_6980);
and U7916 (N_7916,N_6886,N_7233);
and U7917 (N_7917,N_7226,N_7466);
nor U7918 (N_7918,N_7494,N_6900);
xor U7919 (N_7919,N_7335,N_6943);
nor U7920 (N_7920,N_7263,N_7162);
nor U7921 (N_7921,N_7390,N_7105);
and U7922 (N_7922,N_6895,N_7199);
or U7923 (N_7923,N_6885,N_7269);
or U7924 (N_7924,N_7141,N_7358);
xnor U7925 (N_7925,N_7067,N_7219);
and U7926 (N_7926,N_7111,N_7127);
nor U7927 (N_7927,N_7109,N_7227);
xnor U7928 (N_7928,N_7031,N_6973);
nor U7929 (N_7929,N_7418,N_7342);
xnor U7930 (N_7930,N_7318,N_7468);
nand U7931 (N_7931,N_7005,N_7023);
nor U7932 (N_7932,N_7399,N_7320);
nand U7933 (N_7933,N_7194,N_7035);
and U7934 (N_7934,N_7244,N_7266);
nand U7935 (N_7935,N_7171,N_7285);
or U7936 (N_7936,N_7222,N_7321);
nor U7937 (N_7937,N_7154,N_7032);
xnor U7938 (N_7938,N_6884,N_7378);
and U7939 (N_7939,N_6966,N_7440);
xor U7940 (N_7940,N_6917,N_7320);
or U7941 (N_7941,N_7073,N_6882);
or U7942 (N_7942,N_7362,N_7345);
or U7943 (N_7943,N_7390,N_7469);
xnor U7944 (N_7944,N_7452,N_7187);
nand U7945 (N_7945,N_7143,N_7482);
nor U7946 (N_7946,N_6999,N_7218);
xor U7947 (N_7947,N_7479,N_7125);
or U7948 (N_7948,N_7372,N_6990);
xnor U7949 (N_7949,N_7075,N_7487);
nor U7950 (N_7950,N_7471,N_6892);
xor U7951 (N_7951,N_7257,N_7018);
or U7952 (N_7952,N_7014,N_7125);
and U7953 (N_7953,N_7440,N_6888);
or U7954 (N_7954,N_7177,N_6962);
xnor U7955 (N_7955,N_6905,N_7426);
or U7956 (N_7956,N_7132,N_7385);
or U7957 (N_7957,N_6878,N_7048);
nor U7958 (N_7958,N_7147,N_6947);
or U7959 (N_7959,N_6907,N_7464);
and U7960 (N_7960,N_7238,N_7252);
nor U7961 (N_7961,N_6987,N_7475);
nand U7962 (N_7962,N_7412,N_7355);
and U7963 (N_7963,N_7116,N_7280);
and U7964 (N_7964,N_7463,N_7293);
and U7965 (N_7965,N_7149,N_7438);
nand U7966 (N_7966,N_7379,N_6914);
nor U7967 (N_7967,N_7491,N_7053);
or U7968 (N_7968,N_7425,N_7172);
or U7969 (N_7969,N_7205,N_7214);
and U7970 (N_7970,N_7267,N_7010);
xnor U7971 (N_7971,N_7089,N_7464);
or U7972 (N_7972,N_7222,N_7475);
nor U7973 (N_7973,N_7154,N_7494);
xor U7974 (N_7974,N_7497,N_7312);
nor U7975 (N_7975,N_7261,N_7301);
or U7976 (N_7976,N_7289,N_6903);
and U7977 (N_7977,N_6994,N_7334);
xor U7978 (N_7978,N_6964,N_7270);
or U7979 (N_7979,N_7374,N_7464);
or U7980 (N_7980,N_7284,N_6997);
xnor U7981 (N_7981,N_7024,N_7494);
and U7982 (N_7982,N_7451,N_7333);
nor U7983 (N_7983,N_7019,N_7486);
nand U7984 (N_7984,N_7211,N_6934);
nand U7985 (N_7985,N_7153,N_7356);
and U7986 (N_7986,N_6943,N_7123);
and U7987 (N_7987,N_7010,N_7463);
nand U7988 (N_7988,N_7268,N_6985);
nand U7989 (N_7989,N_7435,N_7453);
and U7990 (N_7990,N_6990,N_7310);
nand U7991 (N_7991,N_7430,N_7149);
nand U7992 (N_7992,N_7401,N_7174);
and U7993 (N_7993,N_6942,N_7329);
and U7994 (N_7994,N_7309,N_7457);
xnor U7995 (N_7995,N_7453,N_7343);
and U7996 (N_7996,N_7064,N_7345);
nand U7997 (N_7997,N_7097,N_7023);
or U7998 (N_7998,N_7470,N_6893);
and U7999 (N_7999,N_7272,N_7036);
or U8000 (N_8000,N_7352,N_7273);
and U8001 (N_8001,N_6978,N_7274);
nand U8002 (N_8002,N_7363,N_7077);
nor U8003 (N_8003,N_6949,N_7358);
and U8004 (N_8004,N_7127,N_7465);
or U8005 (N_8005,N_7019,N_7365);
xnor U8006 (N_8006,N_7002,N_6969);
xor U8007 (N_8007,N_6945,N_7037);
and U8008 (N_8008,N_7249,N_7080);
and U8009 (N_8009,N_7001,N_6879);
nand U8010 (N_8010,N_7497,N_6919);
nand U8011 (N_8011,N_7422,N_6977);
and U8012 (N_8012,N_6937,N_6999);
xnor U8013 (N_8013,N_7065,N_7453);
and U8014 (N_8014,N_7054,N_7081);
and U8015 (N_8015,N_6970,N_7025);
nand U8016 (N_8016,N_6892,N_7393);
nor U8017 (N_8017,N_7006,N_7136);
or U8018 (N_8018,N_7437,N_7335);
and U8019 (N_8019,N_7381,N_7359);
xor U8020 (N_8020,N_7021,N_7427);
nor U8021 (N_8021,N_7466,N_7488);
nand U8022 (N_8022,N_6983,N_7462);
xor U8023 (N_8023,N_7370,N_7174);
nor U8024 (N_8024,N_6974,N_7426);
or U8025 (N_8025,N_7469,N_7287);
or U8026 (N_8026,N_7154,N_7196);
or U8027 (N_8027,N_7183,N_7339);
nor U8028 (N_8028,N_7335,N_7363);
nand U8029 (N_8029,N_7298,N_7307);
nand U8030 (N_8030,N_7020,N_6886);
or U8031 (N_8031,N_7410,N_6928);
or U8032 (N_8032,N_7174,N_6954);
nor U8033 (N_8033,N_7028,N_7070);
xnor U8034 (N_8034,N_7079,N_6999);
nand U8035 (N_8035,N_7129,N_6892);
xnor U8036 (N_8036,N_7473,N_7379);
nand U8037 (N_8037,N_6897,N_7006);
or U8038 (N_8038,N_7485,N_6909);
nor U8039 (N_8039,N_6999,N_7068);
or U8040 (N_8040,N_7134,N_7061);
xor U8041 (N_8041,N_7275,N_6934);
and U8042 (N_8042,N_7018,N_7158);
nor U8043 (N_8043,N_6908,N_7358);
or U8044 (N_8044,N_7335,N_6960);
nand U8045 (N_8045,N_7185,N_6924);
nand U8046 (N_8046,N_7379,N_7469);
or U8047 (N_8047,N_7453,N_7315);
nor U8048 (N_8048,N_7111,N_7176);
nor U8049 (N_8049,N_7361,N_6985);
or U8050 (N_8050,N_7110,N_7127);
or U8051 (N_8051,N_7356,N_6952);
and U8052 (N_8052,N_7088,N_6929);
or U8053 (N_8053,N_6941,N_7037);
and U8054 (N_8054,N_7120,N_6926);
or U8055 (N_8055,N_7458,N_6883);
nor U8056 (N_8056,N_7046,N_6937);
xor U8057 (N_8057,N_7127,N_6903);
nand U8058 (N_8058,N_7132,N_7093);
xor U8059 (N_8059,N_7006,N_7097);
nor U8060 (N_8060,N_7348,N_7101);
xnor U8061 (N_8061,N_7456,N_7060);
or U8062 (N_8062,N_7371,N_7435);
nand U8063 (N_8063,N_7326,N_7016);
or U8064 (N_8064,N_7445,N_7165);
xnor U8065 (N_8065,N_7046,N_6989);
or U8066 (N_8066,N_6926,N_7437);
or U8067 (N_8067,N_7362,N_6908);
or U8068 (N_8068,N_7482,N_7407);
nand U8069 (N_8069,N_7389,N_7254);
nand U8070 (N_8070,N_7312,N_7135);
or U8071 (N_8071,N_7433,N_7235);
and U8072 (N_8072,N_7238,N_7415);
and U8073 (N_8073,N_7320,N_7263);
or U8074 (N_8074,N_7170,N_7224);
or U8075 (N_8075,N_6882,N_7433);
nand U8076 (N_8076,N_7168,N_7373);
nand U8077 (N_8077,N_7258,N_7070);
or U8078 (N_8078,N_7222,N_7067);
or U8079 (N_8079,N_7459,N_6911);
nand U8080 (N_8080,N_7384,N_7462);
nand U8081 (N_8081,N_7466,N_7434);
or U8082 (N_8082,N_7242,N_7240);
or U8083 (N_8083,N_7480,N_6938);
xor U8084 (N_8084,N_7425,N_7119);
nand U8085 (N_8085,N_7113,N_7087);
and U8086 (N_8086,N_7299,N_7433);
nor U8087 (N_8087,N_7466,N_6899);
or U8088 (N_8088,N_7061,N_6942);
xnor U8089 (N_8089,N_7154,N_7348);
or U8090 (N_8090,N_7006,N_7171);
nor U8091 (N_8091,N_7248,N_7345);
or U8092 (N_8092,N_7423,N_7146);
or U8093 (N_8093,N_7007,N_7024);
xor U8094 (N_8094,N_7187,N_7113);
and U8095 (N_8095,N_6908,N_7469);
or U8096 (N_8096,N_6953,N_7445);
nand U8097 (N_8097,N_7022,N_6958);
xnor U8098 (N_8098,N_6896,N_7029);
nor U8099 (N_8099,N_7062,N_7170);
nor U8100 (N_8100,N_7203,N_7066);
nand U8101 (N_8101,N_7176,N_7041);
or U8102 (N_8102,N_7066,N_7417);
xnor U8103 (N_8103,N_7031,N_6875);
nor U8104 (N_8104,N_6913,N_6876);
nand U8105 (N_8105,N_7379,N_7055);
and U8106 (N_8106,N_6963,N_7205);
and U8107 (N_8107,N_7487,N_6919);
nor U8108 (N_8108,N_7002,N_7491);
nand U8109 (N_8109,N_6937,N_7251);
nor U8110 (N_8110,N_7265,N_7190);
xor U8111 (N_8111,N_6988,N_7271);
and U8112 (N_8112,N_6992,N_7437);
nor U8113 (N_8113,N_7035,N_7398);
or U8114 (N_8114,N_6951,N_7421);
and U8115 (N_8115,N_6997,N_7497);
or U8116 (N_8116,N_7279,N_7114);
or U8117 (N_8117,N_7273,N_7445);
nor U8118 (N_8118,N_7158,N_6975);
nor U8119 (N_8119,N_6953,N_7165);
xor U8120 (N_8120,N_7111,N_6914);
or U8121 (N_8121,N_7422,N_6925);
or U8122 (N_8122,N_7111,N_7316);
or U8123 (N_8123,N_6996,N_7063);
or U8124 (N_8124,N_7289,N_7373);
nor U8125 (N_8125,N_7737,N_7706);
nand U8126 (N_8126,N_8121,N_7618);
nor U8127 (N_8127,N_7540,N_7928);
nor U8128 (N_8128,N_7527,N_8018);
xnor U8129 (N_8129,N_8037,N_7855);
xor U8130 (N_8130,N_7833,N_7735);
nor U8131 (N_8131,N_8109,N_7890);
xor U8132 (N_8132,N_7940,N_7663);
nand U8133 (N_8133,N_7981,N_7589);
nand U8134 (N_8134,N_7807,N_7953);
xnor U8135 (N_8135,N_7742,N_7688);
xor U8136 (N_8136,N_7858,N_7636);
or U8137 (N_8137,N_7776,N_7613);
nand U8138 (N_8138,N_7673,N_7917);
or U8139 (N_8139,N_7511,N_8074);
nand U8140 (N_8140,N_7767,N_7924);
or U8141 (N_8141,N_8010,N_7604);
nor U8142 (N_8142,N_8106,N_8009);
nor U8143 (N_8143,N_7734,N_7582);
and U8144 (N_8144,N_8052,N_7725);
nand U8145 (N_8145,N_7709,N_7947);
and U8146 (N_8146,N_7643,N_7983);
xor U8147 (N_8147,N_7978,N_7514);
nor U8148 (N_8148,N_7634,N_7930);
or U8149 (N_8149,N_7875,N_7968);
nand U8150 (N_8150,N_7784,N_8093);
and U8151 (N_8151,N_7820,N_7568);
nand U8152 (N_8152,N_7899,N_7842);
nand U8153 (N_8153,N_7547,N_8075);
xor U8154 (N_8154,N_7621,N_7977);
nand U8155 (N_8155,N_7843,N_7641);
xor U8156 (N_8156,N_7707,N_7727);
or U8157 (N_8157,N_7720,N_7874);
xnor U8158 (N_8158,N_7597,N_7608);
nand U8159 (N_8159,N_7505,N_8029);
nand U8160 (N_8160,N_7691,N_7648);
or U8161 (N_8161,N_7835,N_7906);
nor U8162 (N_8162,N_7640,N_8124);
and U8163 (N_8163,N_7609,N_7572);
and U8164 (N_8164,N_7635,N_7620);
nand U8165 (N_8165,N_7837,N_7586);
or U8166 (N_8166,N_8105,N_7852);
nor U8167 (N_8167,N_7984,N_7530);
and U8168 (N_8168,N_7980,N_7740);
nand U8169 (N_8169,N_8058,N_7768);
nor U8170 (N_8170,N_7877,N_7506);
xor U8171 (N_8171,N_7678,N_8080);
nand U8172 (N_8172,N_7779,N_7675);
nand U8173 (N_8173,N_7934,N_8030);
or U8174 (N_8174,N_7670,N_7948);
or U8175 (N_8175,N_7668,N_7769);
or U8176 (N_8176,N_7856,N_8086);
nor U8177 (N_8177,N_7610,N_7908);
nor U8178 (N_8178,N_7646,N_8055);
nand U8179 (N_8179,N_7519,N_7607);
nand U8180 (N_8180,N_7717,N_8116);
xor U8181 (N_8181,N_7799,N_7606);
xnor U8182 (N_8182,N_7937,N_8059);
nand U8183 (N_8183,N_7963,N_7942);
nor U8184 (N_8184,N_7950,N_7927);
nor U8185 (N_8185,N_7793,N_7971);
xor U8186 (N_8186,N_7726,N_7712);
nand U8187 (N_8187,N_7830,N_8017);
xnor U8188 (N_8188,N_7571,N_8011);
nor U8189 (N_8189,N_7790,N_7796);
or U8190 (N_8190,N_7555,N_7987);
nor U8191 (N_8191,N_7680,N_7693);
xnor U8192 (N_8192,N_7681,N_7504);
xor U8193 (N_8193,N_7660,N_7774);
nand U8194 (N_8194,N_7944,N_8005);
and U8195 (N_8195,N_7755,N_7913);
xnor U8196 (N_8196,N_7894,N_7603);
or U8197 (N_8197,N_7638,N_7801);
xnor U8198 (N_8198,N_8061,N_7936);
and U8199 (N_8199,N_7736,N_7600);
or U8200 (N_8200,N_7509,N_7869);
nand U8201 (N_8201,N_7683,N_8047);
or U8202 (N_8202,N_8049,N_7792);
and U8203 (N_8203,N_7554,N_8036);
or U8204 (N_8204,N_7721,N_7876);
and U8205 (N_8205,N_8008,N_8042);
and U8206 (N_8206,N_7901,N_7816);
and U8207 (N_8207,N_7786,N_7914);
xnor U8208 (N_8208,N_7840,N_7757);
and U8209 (N_8209,N_7775,N_7849);
and U8210 (N_8210,N_7538,N_7829);
nor U8211 (N_8211,N_7935,N_7549);
nor U8212 (N_8212,N_8107,N_7574);
xnor U8213 (N_8213,N_7637,N_7836);
xnor U8214 (N_8214,N_7868,N_7897);
nand U8215 (N_8215,N_7803,N_7754);
nor U8216 (N_8216,N_8056,N_7535);
nor U8217 (N_8217,N_7933,N_7871);
xor U8218 (N_8218,N_7850,N_7878);
nand U8219 (N_8219,N_8067,N_7602);
or U8220 (N_8220,N_7999,N_7872);
nand U8221 (N_8221,N_7516,N_7985);
nand U8222 (N_8222,N_7809,N_7748);
and U8223 (N_8223,N_7870,N_7827);
nand U8224 (N_8224,N_8064,N_7806);
nor U8225 (N_8225,N_7524,N_8048);
nand U8226 (N_8226,N_7986,N_7811);
xnor U8227 (N_8227,N_8031,N_7567);
and U8228 (N_8228,N_7605,N_8054);
and U8229 (N_8229,N_7922,N_7818);
or U8230 (N_8230,N_8114,N_8092);
xnor U8231 (N_8231,N_8072,N_7565);
and U8232 (N_8232,N_8083,N_7627);
or U8233 (N_8233,N_7698,N_7629);
nor U8234 (N_8234,N_7665,N_7817);
xor U8235 (N_8235,N_7543,N_7728);
and U8236 (N_8236,N_7961,N_7802);
and U8237 (N_8237,N_7743,N_7882);
nor U8238 (N_8238,N_7791,N_7741);
nand U8239 (N_8239,N_7584,N_8103);
nor U8240 (N_8240,N_7708,N_7886);
or U8241 (N_8241,N_7896,N_7761);
nor U8242 (N_8242,N_8070,N_7911);
or U8243 (N_8243,N_7888,N_7957);
xnor U8244 (N_8244,N_8014,N_7601);
xnor U8245 (N_8245,N_8123,N_7879);
nor U8246 (N_8246,N_7825,N_8004);
or U8247 (N_8247,N_7612,N_8113);
and U8248 (N_8248,N_7510,N_7976);
or U8249 (N_8249,N_7531,N_7501);
or U8250 (N_8250,N_8079,N_7599);
or U8251 (N_8251,N_7580,N_7611);
xnor U8252 (N_8252,N_8046,N_7548);
xor U8253 (N_8253,N_7955,N_7916);
xnor U8254 (N_8254,N_7557,N_7521);
or U8255 (N_8255,N_7639,N_7782);
nor U8256 (N_8256,N_7810,N_7903);
nor U8257 (N_8257,N_7762,N_7772);
nor U8258 (N_8258,N_7552,N_8057);
nor U8259 (N_8259,N_7729,N_7566);
or U8260 (N_8260,N_7625,N_7834);
or U8261 (N_8261,N_7657,N_8087);
or U8262 (N_8262,N_8104,N_7969);
and U8263 (N_8263,N_7518,N_8040);
xnor U8264 (N_8264,N_7528,N_8088);
nand U8265 (N_8265,N_7700,N_7551);
nand U8266 (N_8266,N_7958,N_7997);
or U8267 (N_8267,N_7529,N_7503);
xor U8268 (N_8268,N_8100,N_7919);
or U8269 (N_8269,N_7838,N_7777);
nand U8270 (N_8270,N_8095,N_8015);
xor U8271 (N_8271,N_8089,N_7770);
or U8272 (N_8272,N_7536,N_7560);
nand U8273 (N_8273,N_7576,N_7993);
nor U8274 (N_8274,N_7645,N_7695);
nor U8275 (N_8275,N_7533,N_8021);
and U8276 (N_8276,N_7750,N_8077);
xor U8277 (N_8277,N_7546,N_7841);
and U8278 (N_8278,N_8016,N_7739);
or U8279 (N_8279,N_7656,N_8060);
xnor U8280 (N_8280,N_8084,N_7990);
or U8281 (N_8281,N_7701,N_8020);
and U8282 (N_8282,N_7960,N_7523);
nor U8283 (N_8283,N_8007,N_7705);
nor U8284 (N_8284,N_7598,N_7926);
and U8285 (N_8285,N_7515,N_7884);
and U8286 (N_8286,N_7800,N_7561);
nor U8287 (N_8287,N_8038,N_7915);
xor U8288 (N_8288,N_7594,N_7704);
nor U8289 (N_8289,N_8065,N_7550);
xnor U8290 (N_8290,N_7661,N_8101);
or U8291 (N_8291,N_7655,N_7822);
and U8292 (N_8292,N_7659,N_7780);
nand U8293 (N_8293,N_7692,N_7844);
xnor U8294 (N_8294,N_7889,N_7824);
nand U8295 (N_8295,N_8120,N_8019);
nand U8296 (N_8296,N_7633,N_7732);
and U8297 (N_8297,N_7920,N_7956);
nand U8298 (N_8298,N_7970,N_8000);
xor U8299 (N_8299,N_7859,N_7685);
xor U8300 (N_8300,N_7677,N_7595);
and U8301 (N_8301,N_7626,N_7642);
nand U8302 (N_8302,N_7716,N_7553);
and U8303 (N_8303,N_7781,N_7938);
nor U8304 (N_8304,N_7723,N_7585);
or U8305 (N_8305,N_7587,N_7703);
nor U8306 (N_8306,N_7787,N_7904);
and U8307 (N_8307,N_7860,N_8099);
xnor U8308 (N_8308,N_7764,N_7593);
or U8309 (N_8309,N_7541,N_7672);
xnor U8310 (N_8310,N_7615,N_7885);
nor U8311 (N_8311,N_7722,N_7814);
or U8312 (N_8312,N_7865,N_7733);
nand U8313 (N_8313,N_7846,N_7819);
or U8314 (N_8314,N_7679,N_7813);
xnor U8315 (N_8315,N_7545,N_7851);
or U8316 (N_8316,N_7632,N_8118);
nand U8317 (N_8317,N_7949,N_7715);
and U8318 (N_8318,N_7697,N_7500);
nand U8319 (N_8319,N_7630,N_7873);
and U8320 (N_8320,N_7783,N_7974);
xor U8321 (N_8321,N_8026,N_7893);
nand U8322 (N_8322,N_7578,N_7570);
and U8323 (N_8323,N_7943,N_8003);
or U8324 (N_8324,N_7912,N_7861);
xnor U8325 (N_8325,N_7756,N_8051);
and U8326 (N_8326,N_7828,N_7508);
nor U8327 (N_8327,N_7614,N_7525);
nand U8328 (N_8328,N_8078,N_8012);
or U8329 (N_8329,N_7517,N_7952);
xor U8330 (N_8330,N_7789,N_7684);
xnor U8331 (N_8331,N_7895,N_7752);
nand U8332 (N_8332,N_7946,N_7805);
nand U8333 (N_8333,N_7579,N_7682);
or U8334 (N_8334,N_7988,N_8053);
and U8335 (N_8335,N_7902,N_7959);
nor U8336 (N_8336,N_7651,N_7596);
nand U8337 (N_8337,N_8025,N_8108);
nand U8338 (N_8338,N_7649,N_7972);
or U8339 (N_8339,N_7652,N_7992);
or U8340 (N_8340,N_7713,N_7711);
xor U8341 (N_8341,N_7773,N_7989);
xnor U8342 (N_8342,N_8097,N_8028);
nand U8343 (N_8343,N_7839,N_7590);
nor U8344 (N_8344,N_8071,N_8034);
xnor U8345 (N_8345,N_8094,N_7994);
nand U8346 (N_8346,N_7905,N_8085);
nand U8347 (N_8347,N_7699,N_8066);
nor U8348 (N_8348,N_7512,N_7619);
xnor U8349 (N_8349,N_7965,N_7719);
or U8350 (N_8350,N_7794,N_7520);
nand U8351 (N_8351,N_7746,N_7667);
or U8352 (N_8352,N_8110,N_7866);
or U8353 (N_8353,N_8076,N_7558);
or U8354 (N_8354,N_7798,N_7687);
nor U8355 (N_8355,N_7671,N_7804);
nand U8356 (N_8356,N_7556,N_7867);
or U8357 (N_8357,N_7815,N_7907);
xor U8358 (N_8358,N_7845,N_7666);
xor U8359 (N_8359,N_7542,N_7622);
nand U8360 (N_8360,N_8043,N_7881);
and U8361 (N_8361,N_7653,N_7563);
nand U8362 (N_8362,N_8102,N_8098);
nor U8363 (N_8363,N_7966,N_8033);
and U8364 (N_8364,N_8112,N_7854);
xor U8365 (N_8365,N_7941,N_7945);
xor U8366 (N_8366,N_7591,N_7583);
and U8367 (N_8367,N_7887,N_7778);
and U8368 (N_8368,N_7559,N_7749);
nor U8369 (N_8369,N_7588,N_7996);
xnor U8370 (N_8370,N_7674,N_7647);
nand U8371 (N_8371,N_7724,N_7628);
nor U8372 (N_8372,N_7853,N_7812);
or U8373 (N_8373,N_8050,N_7581);
or U8374 (N_8374,N_7880,N_7502);
xor U8375 (N_8375,N_7891,N_7650);
nand U8376 (N_8376,N_7951,N_7702);
xnor U8377 (N_8377,N_7785,N_7532);
nand U8378 (N_8378,N_7730,N_7537);
nand U8379 (N_8379,N_7522,N_8090);
nor U8380 (N_8380,N_7654,N_7751);
nand U8381 (N_8381,N_7795,N_7689);
xnor U8382 (N_8382,N_7964,N_8032);
or U8383 (N_8383,N_7765,N_7975);
or U8384 (N_8384,N_7967,N_8119);
nor U8385 (N_8385,N_8117,N_8068);
xnor U8386 (N_8386,N_7898,N_8045);
or U8387 (N_8387,N_7760,N_7892);
or U8388 (N_8388,N_7771,N_7939);
or U8389 (N_8389,N_7747,N_7714);
nand U8390 (N_8390,N_7696,N_8096);
and U8391 (N_8391,N_7577,N_7863);
xor U8392 (N_8392,N_7831,N_7564);
or U8393 (N_8393,N_8069,N_7573);
or U8394 (N_8394,N_7932,N_7534);
and U8395 (N_8395,N_8024,N_7797);
nand U8396 (N_8396,N_8062,N_8027);
nand U8397 (N_8397,N_7718,N_7918);
or U8398 (N_8398,N_7826,N_7669);
or U8399 (N_8399,N_7788,N_8111);
or U8400 (N_8400,N_7857,N_7982);
nand U8401 (N_8401,N_7900,N_8081);
xnor U8402 (N_8402,N_7758,N_7623);
xnor U8403 (N_8403,N_7923,N_8002);
nand U8404 (N_8404,N_7562,N_7738);
xnor U8405 (N_8405,N_7929,N_7624);
and U8406 (N_8406,N_8044,N_7998);
nor U8407 (N_8407,N_7847,N_7539);
nand U8408 (N_8408,N_7832,N_7662);
nand U8409 (N_8409,N_7526,N_7823);
nor U8410 (N_8410,N_7763,N_7617);
and U8411 (N_8411,N_7690,N_7694);
and U8412 (N_8412,N_7745,N_7676);
nor U8413 (N_8413,N_7513,N_7864);
nand U8414 (N_8414,N_7808,N_8063);
and U8415 (N_8415,N_7731,N_7883);
xnor U8416 (N_8416,N_8006,N_7686);
xnor U8417 (N_8417,N_7962,N_8001);
xor U8418 (N_8418,N_7664,N_8041);
or U8419 (N_8419,N_7569,N_7931);
nor U8420 (N_8420,N_7862,N_8091);
nor U8421 (N_8421,N_7973,N_7631);
nand U8422 (N_8422,N_7575,N_7925);
or U8423 (N_8423,N_8082,N_8022);
nand U8424 (N_8424,N_8035,N_8115);
and U8425 (N_8425,N_7848,N_8013);
xnor U8426 (N_8426,N_7821,N_7644);
nor U8427 (N_8427,N_7507,N_7744);
nor U8428 (N_8428,N_8023,N_8073);
nand U8429 (N_8429,N_7909,N_7658);
xor U8430 (N_8430,N_8039,N_7710);
nor U8431 (N_8431,N_7995,N_7544);
xor U8432 (N_8432,N_8122,N_7910);
nor U8433 (N_8433,N_7759,N_7753);
xor U8434 (N_8434,N_7921,N_7954);
nand U8435 (N_8435,N_7616,N_7979);
or U8436 (N_8436,N_7991,N_7592);
nand U8437 (N_8437,N_7766,N_7539);
or U8438 (N_8438,N_7598,N_7757);
and U8439 (N_8439,N_7911,N_7591);
or U8440 (N_8440,N_7738,N_7923);
xor U8441 (N_8441,N_7948,N_7965);
nand U8442 (N_8442,N_7967,N_8108);
nor U8443 (N_8443,N_7745,N_8046);
xnor U8444 (N_8444,N_7504,N_7785);
nor U8445 (N_8445,N_7867,N_7690);
or U8446 (N_8446,N_7945,N_7722);
nand U8447 (N_8447,N_8120,N_7538);
nor U8448 (N_8448,N_8096,N_7926);
xnor U8449 (N_8449,N_7854,N_7813);
nor U8450 (N_8450,N_7779,N_7701);
nand U8451 (N_8451,N_7760,N_7834);
xnor U8452 (N_8452,N_7745,N_7539);
nand U8453 (N_8453,N_7562,N_7802);
or U8454 (N_8454,N_7868,N_7558);
or U8455 (N_8455,N_7944,N_7754);
and U8456 (N_8456,N_7693,N_7993);
nor U8457 (N_8457,N_7757,N_7702);
or U8458 (N_8458,N_7535,N_7609);
and U8459 (N_8459,N_7743,N_7973);
or U8460 (N_8460,N_8083,N_8095);
xor U8461 (N_8461,N_7834,N_7927);
xnor U8462 (N_8462,N_7553,N_7696);
or U8463 (N_8463,N_7561,N_7934);
nor U8464 (N_8464,N_7641,N_7783);
and U8465 (N_8465,N_7904,N_7817);
nor U8466 (N_8466,N_8106,N_7517);
nand U8467 (N_8467,N_7764,N_8036);
or U8468 (N_8468,N_7834,N_8041);
or U8469 (N_8469,N_7670,N_7761);
and U8470 (N_8470,N_7599,N_7538);
nand U8471 (N_8471,N_7977,N_7672);
xor U8472 (N_8472,N_7590,N_8043);
and U8473 (N_8473,N_7912,N_8084);
and U8474 (N_8474,N_7610,N_7740);
xor U8475 (N_8475,N_7851,N_7542);
xor U8476 (N_8476,N_7818,N_7600);
or U8477 (N_8477,N_7598,N_7835);
and U8478 (N_8478,N_7811,N_7851);
xor U8479 (N_8479,N_7669,N_7531);
or U8480 (N_8480,N_7513,N_7884);
or U8481 (N_8481,N_8036,N_7906);
nor U8482 (N_8482,N_8119,N_7685);
xnor U8483 (N_8483,N_7996,N_7553);
or U8484 (N_8484,N_7955,N_8087);
nor U8485 (N_8485,N_7885,N_7963);
xor U8486 (N_8486,N_7547,N_7868);
or U8487 (N_8487,N_7639,N_7811);
nor U8488 (N_8488,N_7517,N_7716);
and U8489 (N_8489,N_7887,N_7717);
and U8490 (N_8490,N_7666,N_7524);
nor U8491 (N_8491,N_7865,N_7570);
nor U8492 (N_8492,N_7814,N_7503);
and U8493 (N_8493,N_8122,N_7802);
nor U8494 (N_8494,N_7558,N_7551);
and U8495 (N_8495,N_7880,N_7872);
or U8496 (N_8496,N_7795,N_7666);
nand U8497 (N_8497,N_7617,N_7924);
nor U8498 (N_8498,N_7841,N_8009);
and U8499 (N_8499,N_8106,N_7646);
xnor U8500 (N_8500,N_7543,N_7503);
nor U8501 (N_8501,N_7597,N_7644);
nor U8502 (N_8502,N_7741,N_7700);
nor U8503 (N_8503,N_7945,N_7962);
nand U8504 (N_8504,N_7807,N_7533);
nand U8505 (N_8505,N_8104,N_7708);
and U8506 (N_8506,N_7731,N_7741);
and U8507 (N_8507,N_8086,N_7733);
or U8508 (N_8508,N_7607,N_7689);
or U8509 (N_8509,N_8076,N_7974);
and U8510 (N_8510,N_7978,N_7752);
or U8511 (N_8511,N_7597,N_8123);
nor U8512 (N_8512,N_7706,N_7515);
or U8513 (N_8513,N_7690,N_7509);
xnor U8514 (N_8514,N_7532,N_7825);
nor U8515 (N_8515,N_8066,N_7918);
nor U8516 (N_8516,N_7597,N_7756);
or U8517 (N_8517,N_7853,N_7977);
and U8518 (N_8518,N_7687,N_7979);
nor U8519 (N_8519,N_7600,N_7664);
and U8520 (N_8520,N_7977,N_7574);
nand U8521 (N_8521,N_7869,N_7717);
or U8522 (N_8522,N_7737,N_7661);
and U8523 (N_8523,N_7667,N_7590);
nand U8524 (N_8524,N_8051,N_7624);
nor U8525 (N_8525,N_7954,N_7856);
and U8526 (N_8526,N_7888,N_7541);
xor U8527 (N_8527,N_7916,N_7713);
or U8528 (N_8528,N_7753,N_8027);
xnor U8529 (N_8529,N_7605,N_7835);
xnor U8530 (N_8530,N_7808,N_7513);
nor U8531 (N_8531,N_7519,N_7536);
xnor U8532 (N_8532,N_7550,N_7669);
xor U8533 (N_8533,N_7832,N_7647);
nand U8534 (N_8534,N_7647,N_8062);
and U8535 (N_8535,N_8037,N_7906);
xnor U8536 (N_8536,N_7802,N_7670);
xnor U8537 (N_8537,N_7994,N_8007);
nand U8538 (N_8538,N_7800,N_8051);
and U8539 (N_8539,N_7726,N_7884);
or U8540 (N_8540,N_7587,N_7669);
nor U8541 (N_8541,N_7624,N_7896);
or U8542 (N_8542,N_7679,N_8050);
or U8543 (N_8543,N_7988,N_7954);
and U8544 (N_8544,N_7636,N_8100);
xnor U8545 (N_8545,N_7525,N_7583);
nand U8546 (N_8546,N_7632,N_7742);
and U8547 (N_8547,N_7748,N_8103);
nand U8548 (N_8548,N_7733,N_7906);
nand U8549 (N_8549,N_7647,N_7844);
or U8550 (N_8550,N_7602,N_7625);
nand U8551 (N_8551,N_7936,N_7740);
and U8552 (N_8552,N_7613,N_7952);
and U8553 (N_8553,N_7815,N_7622);
xor U8554 (N_8554,N_8042,N_8079);
xnor U8555 (N_8555,N_7772,N_8073);
or U8556 (N_8556,N_7793,N_7862);
nor U8557 (N_8557,N_7708,N_7929);
or U8558 (N_8558,N_8047,N_7598);
or U8559 (N_8559,N_7956,N_8109);
nor U8560 (N_8560,N_8013,N_7744);
nor U8561 (N_8561,N_7900,N_7574);
and U8562 (N_8562,N_8000,N_8071);
and U8563 (N_8563,N_7841,N_7799);
and U8564 (N_8564,N_7934,N_7576);
nand U8565 (N_8565,N_7534,N_7845);
nand U8566 (N_8566,N_8036,N_7859);
nor U8567 (N_8567,N_7810,N_7935);
nor U8568 (N_8568,N_7554,N_7684);
nand U8569 (N_8569,N_7964,N_7801);
xor U8570 (N_8570,N_7725,N_7521);
or U8571 (N_8571,N_8115,N_7792);
or U8572 (N_8572,N_7947,N_8040);
or U8573 (N_8573,N_7975,N_7775);
nor U8574 (N_8574,N_7554,N_7521);
and U8575 (N_8575,N_7761,N_7955);
nand U8576 (N_8576,N_7555,N_8119);
xnor U8577 (N_8577,N_7894,N_7720);
nand U8578 (N_8578,N_7581,N_7768);
xnor U8579 (N_8579,N_7744,N_7953);
and U8580 (N_8580,N_7780,N_7788);
nor U8581 (N_8581,N_7910,N_8060);
and U8582 (N_8582,N_8065,N_7901);
and U8583 (N_8583,N_7649,N_7980);
nand U8584 (N_8584,N_7650,N_7740);
xor U8585 (N_8585,N_7522,N_7819);
nor U8586 (N_8586,N_7819,N_8124);
nand U8587 (N_8587,N_8080,N_7950);
or U8588 (N_8588,N_8014,N_7854);
xnor U8589 (N_8589,N_7921,N_7618);
or U8590 (N_8590,N_7756,N_7536);
xor U8591 (N_8591,N_7833,N_7696);
xnor U8592 (N_8592,N_7773,N_8095);
xnor U8593 (N_8593,N_7817,N_7797);
nor U8594 (N_8594,N_7525,N_7728);
nand U8595 (N_8595,N_7586,N_7600);
and U8596 (N_8596,N_7809,N_7986);
nor U8597 (N_8597,N_7896,N_7506);
nor U8598 (N_8598,N_7640,N_7520);
and U8599 (N_8599,N_8030,N_7942);
or U8600 (N_8600,N_7562,N_8079);
and U8601 (N_8601,N_7879,N_7925);
and U8602 (N_8602,N_8070,N_7584);
nand U8603 (N_8603,N_7997,N_7609);
nand U8604 (N_8604,N_8117,N_7732);
nor U8605 (N_8605,N_8111,N_8110);
and U8606 (N_8606,N_7763,N_8052);
or U8607 (N_8607,N_7837,N_7972);
xor U8608 (N_8608,N_7945,N_8071);
xor U8609 (N_8609,N_8124,N_8022);
and U8610 (N_8610,N_7910,N_7556);
nand U8611 (N_8611,N_8064,N_8012);
and U8612 (N_8612,N_7606,N_7911);
xnor U8613 (N_8613,N_7620,N_8011);
nor U8614 (N_8614,N_7950,N_7866);
nor U8615 (N_8615,N_7631,N_7873);
xnor U8616 (N_8616,N_7787,N_7574);
xnor U8617 (N_8617,N_7923,N_7758);
xnor U8618 (N_8618,N_7691,N_7658);
or U8619 (N_8619,N_7751,N_7826);
or U8620 (N_8620,N_7729,N_7762);
nor U8621 (N_8621,N_7824,N_7587);
nor U8622 (N_8622,N_7798,N_7645);
xnor U8623 (N_8623,N_7959,N_7834);
or U8624 (N_8624,N_7984,N_7532);
and U8625 (N_8625,N_7881,N_7559);
or U8626 (N_8626,N_7706,N_7842);
nor U8627 (N_8627,N_8119,N_8031);
and U8628 (N_8628,N_7863,N_7636);
nand U8629 (N_8629,N_7780,N_7688);
nand U8630 (N_8630,N_7673,N_8041);
or U8631 (N_8631,N_7989,N_7572);
and U8632 (N_8632,N_7991,N_7625);
nand U8633 (N_8633,N_7872,N_7852);
or U8634 (N_8634,N_7749,N_7964);
and U8635 (N_8635,N_7535,N_7747);
nand U8636 (N_8636,N_8046,N_7901);
nand U8637 (N_8637,N_7929,N_7622);
and U8638 (N_8638,N_7912,N_7818);
nand U8639 (N_8639,N_7758,N_7549);
or U8640 (N_8640,N_7947,N_7724);
and U8641 (N_8641,N_7979,N_7794);
nand U8642 (N_8642,N_8038,N_7734);
nor U8643 (N_8643,N_7992,N_8010);
or U8644 (N_8644,N_7905,N_7952);
xnor U8645 (N_8645,N_7683,N_7704);
and U8646 (N_8646,N_7834,N_7965);
and U8647 (N_8647,N_7530,N_7779);
nor U8648 (N_8648,N_7797,N_7963);
and U8649 (N_8649,N_7873,N_7704);
nor U8650 (N_8650,N_7595,N_7702);
nand U8651 (N_8651,N_7573,N_7913);
xor U8652 (N_8652,N_7905,N_8000);
xnor U8653 (N_8653,N_7797,N_7523);
or U8654 (N_8654,N_7865,N_7993);
nor U8655 (N_8655,N_7924,N_7611);
nand U8656 (N_8656,N_7914,N_8095);
nand U8657 (N_8657,N_8005,N_8119);
nor U8658 (N_8658,N_7942,N_8037);
nand U8659 (N_8659,N_7871,N_7526);
or U8660 (N_8660,N_8108,N_7725);
nor U8661 (N_8661,N_7991,N_7944);
nand U8662 (N_8662,N_7900,N_7867);
or U8663 (N_8663,N_7836,N_8067);
and U8664 (N_8664,N_7787,N_8122);
nand U8665 (N_8665,N_7825,N_7781);
xor U8666 (N_8666,N_7993,N_7899);
xor U8667 (N_8667,N_7933,N_7710);
or U8668 (N_8668,N_7518,N_7804);
or U8669 (N_8669,N_7591,N_7956);
nand U8670 (N_8670,N_7985,N_7912);
and U8671 (N_8671,N_7699,N_7647);
nor U8672 (N_8672,N_7569,N_8110);
or U8673 (N_8673,N_7526,N_7611);
nor U8674 (N_8674,N_7904,N_8110);
nor U8675 (N_8675,N_8017,N_8082);
nand U8676 (N_8676,N_7582,N_7534);
nand U8677 (N_8677,N_7571,N_8124);
or U8678 (N_8678,N_7715,N_7507);
and U8679 (N_8679,N_8096,N_7504);
nand U8680 (N_8680,N_8030,N_7685);
and U8681 (N_8681,N_7724,N_8121);
nor U8682 (N_8682,N_8072,N_7801);
xnor U8683 (N_8683,N_7984,N_7898);
xor U8684 (N_8684,N_7977,N_7630);
or U8685 (N_8685,N_7774,N_7981);
nand U8686 (N_8686,N_7999,N_7743);
xor U8687 (N_8687,N_7966,N_7543);
nor U8688 (N_8688,N_7637,N_7997);
xnor U8689 (N_8689,N_7856,N_7909);
xor U8690 (N_8690,N_7519,N_8022);
xnor U8691 (N_8691,N_7754,N_8037);
and U8692 (N_8692,N_7893,N_8018);
and U8693 (N_8693,N_7950,N_7880);
nor U8694 (N_8694,N_7518,N_7653);
or U8695 (N_8695,N_7978,N_8000);
nand U8696 (N_8696,N_7870,N_7649);
or U8697 (N_8697,N_7716,N_7900);
and U8698 (N_8698,N_8069,N_7999);
nand U8699 (N_8699,N_7772,N_7572);
or U8700 (N_8700,N_8093,N_7725);
nand U8701 (N_8701,N_8070,N_7615);
xor U8702 (N_8702,N_7876,N_7709);
nor U8703 (N_8703,N_7655,N_7787);
xor U8704 (N_8704,N_7513,N_7698);
xor U8705 (N_8705,N_7772,N_7641);
nand U8706 (N_8706,N_7723,N_7921);
and U8707 (N_8707,N_7999,N_7641);
nor U8708 (N_8708,N_7719,N_8022);
xor U8709 (N_8709,N_7655,N_7605);
nand U8710 (N_8710,N_7927,N_8086);
xor U8711 (N_8711,N_7659,N_7906);
or U8712 (N_8712,N_7556,N_7840);
xor U8713 (N_8713,N_7792,N_7602);
and U8714 (N_8714,N_7804,N_7567);
or U8715 (N_8715,N_7750,N_7676);
nor U8716 (N_8716,N_8005,N_7635);
and U8717 (N_8717,N_7524,N_7764);
nor U8718 (N_8718,N_7694,N_7693);
xnor U8719 (N_8719,N_7539,N_7873);
nor U8720 (N_8720,N_7987,N_7967);
and U8721 (N_8721,N_7853,N_7514);
or U8722 (N_8722,N_7833,N_8030);
and U8723 (N_8723,N_8111,N_7513);
and U8724 (N_8724,N_7982,N_7963);
nor U8725 (N_8725,N_7889,N_7988);
nor U8726 (N_8726,N_8065,N_7949);
or U8727 (N_8727,N_7846,N_7677);
nor U8728 (N_8728,N_7806,N_7569);
and U8729 (N_8729,N_8014,N_7762);
or U8730 (N_8730,N_7558,N_7581);
xor U8731 (N_8731,N_7665,N_7893);
and U8732 (N_8732,N_7800,N_7601);
nor U8733 (N_8733,N_7945,N_7694);
and U8734 (N_8734,N_7819,N_8103);
nor U8735 (N_8735,N_7512,N_7681);
and U8736 (N_8736,N_8120,N_7598);
nand U8737 (N_8737,N_7943,N_8118);
or U8738 (N_8738,N_7927,N_7961);
xnor U8739 (N_8739,N_8063,N_8011);
nor U8740 (N_8740,N_7853,N_7564);
nor U8741 (N_8741,N_8011,N_8080);
or U8742 (N_8742,N_7669,N_8109);
or U8743 (N_8743,N_7800,N_7989);
xor U8744 (N_8744,N_7633,N_7562);
and U8745 (N_8745,N_7808,N_7588);
nand U8746 (N_8746,N_7834,N_7615);
xnor U8747 (N_8747,N_7739,N_7720);
nand U8748 (N_8748,N_7648,N_7895);
xnor U8749 (N_8749,N_7956,N_7558);
nor U8750 (N_8750,N_8630,N_8206);
xor U8751 (N_8751,N_8158,N_8136);
or U8752 (N_8752,N_8716,N_8474);
and U8753 (N_8753,N_8594,N_8374);
xor U8754 (N_8754,N_8420,N_8628);
or U8755 (N_8755,N_8208,N_8307);
or U8756 (N_8756,N_8595,N_8584);
nand U8757 (N_8757,N_8293,N_8703);
nor U8758 (N_8758,N_8183,N_8339);
or U8759 (N_8759,N_8521,N_8234);
or U8760 (N_8760,N_8658,N_8333);
nor U8761 (N_8761,N_8318,N_8589);
and U8762 (N_8762,N_8733,N_8670);
nand U8763 (N_8763,N_8164,N_8572);
and U8764 (N_8764,N_8676,N_8639);
xor U8765 (N_8765,N_8140,N_8240);
or U8766 (N_8766,N_8463,N_8461);
nor U8767 (N_8767,N_8260,N_8534);
and U8768 (N_8768,N_8616,N_8338);
and U8769 (N_8769,N_8618,N_8673);
nor U8770 (N_8770,N_8680,N_8490);
nor U8771 (N_8771,N_8558,N_8223);
nand U8772 (N_8772,N_8276,N_8612);
nor U8773 (N_8773,N_8704,N_8373);
nand U8774 (N_8774,N_8249,N_8479);
or U8775 (N_8775,N_8688,N_8398);
xor U8776 (N_8776,N_8404,N_8361);
xnor U8777 (N_8777,N_8453,N_8264);
nor U8778 (N_8778,N_8334,N_8313);
nand U8779 (N_8779,N_8407,N_8605);
nor U8780 (N_8780,N_8391,N_8532);
xor U8781 (N_8781,N_8135,N_8615);
nand U8782 (N_8782,N_8585,N_8459);
and U8783 (N_8783,N_8263,N_8270);
and U8784 (N_8784,N_8405,N_8531);
nand U8785 (N_8785,N_8233,N_8429);
or U8786 (N_8786,N_8443,N_8554);
nand U8787 (N_8787,N_8286,N_8745);
or U8788 (N_8788,N_8440,N_8672);
or U8789 (N_8789,N_8412,N_8288);
and U8790 (N_8790,N_8316,N_8509);
nand U8791 (N_8791,N_8596,N_8343);
nor U8792 (N_8792,N_8312,N_8484);
or U8793 (N_8793,N_8351,N_8458);
or U8794 (N_8794,N_8719,N_8471);
nand U8795 (N_8795,N_8232,N_8542);
or U8796 (N_8796,N_8267,N_8623);
xnor U8797 (N_8797,N_8151,N_8146);
and U8798 (N_8798,N_8631,N_8283);
and U8799 (N_8799,N_8574,N_8408);
nor U8800 (N_8800,N_8721,N_8529);
or U8801 (N_8801,N_8355,N_8185);
and U8802 (N_8802,N_8485,N_8551);
or U8803 (N_8803,N_8147,N_8362);
xnor U8804 (N_8804,N_8156,N_8261);
nand U8805 (N_8805,N_8285,N_8237);
and U8806 (N_8806,N_8674,N_8567);
nand U8807 (N_8807,N_8132,N_8305);
nor U8808 (N_8808,N_8298,N_8488);
xnor U8809 (N_8809,N_8396,N_8495);
or U8810 (N_8810,N_8191,N_8257);
nand U8811 (N_8811,N_8430,N_8535);
or U8812 (N_8812,N_8347,N_8350);
xor U8813 (N_8813,N_8619,N_8138);
or U8814 (N_8814,N_8211,N_8617);
or U8815 (N_8815,N_8235,N_8248);
and U8816 (N_8816,N_8632,N_8527);
nor U8817 (N_8817,N_8737,N_8345);
nand U8818 (N_8818,N_8171,N_8399);
or U8819 (N_8819,N_8653,N_8370);
nand U8820 (N_8820,N_8513,N_8386);
xor U8821 (N_8821,N_8516,N_8626);
and U8822 (N_8822,N_8418,N_8342);
and U8823 (N_8823,N_8281,N_8512);
or U8824 (N_8824,N_8321,N_8473);
and U8825 (N_8825,N_8246,N_8395);
nor U8826 (N_8826,N_8468,N_8256);
and U8827 (N_8827,N_8460,N_8603);
xor U8828 (N_8828,N_8450,N_8215);
nor U8829 (N_8829,N_8387,N_8525);
nand U8830 (N_8830,N_8648,N_8250);
nor U8831 (N_8831,N_8508,N_8413);
and U8832 (N_8832,N_8165,N_8655);
nand U8833 (N_8833,N_8221,N_8252);
nand U8834 (N_8834,N_8462,N_8664);
or U8835 (N_8835,N_8569,N_8131);
or U8836 (N_8836,N_8651,N_8625);
nor U8837 (N_8837,N_8590,N_8269);
nand U8838 (N_8838,N_8524,N_8601);
nor U8839 (N_8839,N_8592,N_8295);
nand U8840 (N_8840,N_8315,N_8394);
nor U8841 (N_8841,N_8292,N_8369);
nand U8842 (N_8842,N_8702,N_8682);
and U8843 (N_8843,N_8685,N_8465);
and U8844 (N_8844,N_8354,N_8402);
or U8845 (N_8845,N_8176,N_8587);
nand U8846 (N_8846,N_8125,N_8480);
or U8847 (N_8847,N_8352,N_8517);
and U8848 (N_8848,N_8547,N_8503);
nand U8849 (N_8849,N_8643,N_8492);
or U8850 (N_8850,N_8228,N_8642);
nor U8851 (N_8851,N_8679,N_8296);
or U8852 (N_8852,N_8698,N_8403);
or U8853 (N_8853,N_8620,N_8466);
or U8854 (N_8854,N_8477,N_8144);
nand U8855 (N_8855,N_8222,N_8677);
nor U8856 (N_8856,N_8259,N_8134);
and U8857 (N_8857,N_8299,N_8725);
nor U8858 (N_8858,N_8734,N_8720);
nor U8859 (N_8859,N_8634,N_8602);
nor U8860 (N_8860,N_8194,N_8749);
xnor U8861 (N_8861,N_8707,N_8491);
nor U8862 (N_8862,N_8543,N_8435);
nand U8863 (N_8863,N_8741,N_8691);
and U8864 (N_8864,N_8559,N_8700);
or U8865 (N_8865,N_8188,N_8470);
or U8866 (N_8866,N_8381,N_8425);
nor U8867 (N_8867,N_8169,N_8364);
nand U8868 (N_8868,N_8278,N_8337);
xor U8869 (N_8869,N_8282,N_8445);
and U8870 (N_8870,N_8715,N_8376);
and U8871 (N_8871,N_8501,N_8444);
and U8872 (N_8872,N_8437,N_8689);
and U8873 (N_8873,N_8732,N_8694);
or U8874 (N_8874,N_8371,N_8476);
or U8875 (N_8875,N_8708,N_8583);
or U8876 (N_8876,N_8469,N_8375);
and U8877 (N_8877,N_8481,N_8379);
or U8878 (N_8878,N_8254,N_8192);
nand U8879 (N_8879,N_8693,N_8726);
xor U8880 (N_8880,N_8552,N_8538);
or U8881 (N_8881,N_8730,N_8314);
and U8882 (N_8882,N_8515,N_8200);
xnor U8883 (N_8883,N_8209,N_8678);
xor U8884 (N_8884,N_8199,N_8238);
or U8885 (N_8885,N_8181,N_8340);
and U8886 (N_8886,N_8377,N_8239);
or U8887 (N_8887,N_8201,N_8217);
nor U8888 (N_8888,N_8638,N_8493);
or U8889 (N_8889,N_8633,N_8563);
nor U8890 (N_8890,N_8177,N_8159);
and U8891 (N_8891,N_8290,N_8436);
and U8892 (N_8892,N_8539,N_8230);
nor U8893 (N_8893,N_8499,N_8581);
and U8894 (N_8894,N_8520,N_8668);
or U8895 (N_8895,N_8519,N_8243);
or U8896 (N_8896,N_8597,N_8184);
xor U8897 (N_8897,N_8706,N_8656);
nor U8898 (N_8898,N_8550,N_8195);
or U8899 (N_8899,N_8294,N_8744);
nor U8900 (N_8900,N_8378,N_8329);
nor U8901 (N_8901,N_8502,N_8448);
nand U8902 (N_8902,N_8203,N_8665);
nand U8903 (N_8903,N_8560,N_8701);
xor U8904 (N_8904,N_8566,N_8526);
nor U8905 (N_8905,N_8747,N_8145);
nand U8906 (N_8906,N_8220,N_8649);
xnor U8907 (N_8907,N_8696,N_8161);
nor U8908 (N_8908,N_8507,N_8360);
and U8909 (N_8909,N_8393,N_8660);
xnor U8910 (N_8910,N_8671,N_8611);
and U8911 (N_8911,N_8735,N_8434);
nor U8912 (N_8912,N_8586,N_8168);
or U8913 (N_8913,N_8728,N_8406);
nand U8914 (N_8914,N_8301,N_8126);
or U8915 (N_8915,N_8478,N_8322);
or U8916 (N_8916,N_8356,N_8722);
xnor U8917 (N_8917,N_8311,N_8142);
nand U8918 (N_8918,N_8363,N_8353);
nor U8919 (N_8919,N_8262,N_8523);
and U8920 (N_8920,N_8729,N_8537);
nand U8921 (N_8921,N_8179,N_8506);
nor U8922 (N_8922,N_8178,N_8302);
nand U8923 (N_8923,N_8505,N_8604);
xnor U8924 (N_8924,N_8546,N_8731);
nor U8925 (N_8925,N_8385,N_8289);
or U8926 (N_8926,N_8280,N_8582);
nor U8927 (N_8927,N_8401,N_8225);
or U8928 (N_8928,N_8323,N_8482);
or U8929 (N_8929,N_8287,N_8175);
or U8930 (N_8930,N_8357,N_8153);
nand U8931 (N_8931,N_8128,N_8723);
xnor U8932 (N_8932,N_8736,N_8576);
nor U8933 (N_8933,N_8562,N_8455);
and U8934 (N_8934,N_8621,N_8389);
xor U8935 (N_8935,N_8167,N_8675);
or U8936 (N_8936,N_8600,N_8160);
or U8937 (N_8937,N_8207,N_8454);
nor U8938 (N_8938,N_8705,N_8711);
xor U8939 (N_8939,N_8666,N_8258);
xnor U8940 (N_8940,N_8533,N_8186);
nor U8941 (N_8941,N_8622,N_8487);
or U8942 (N_8942,N_8300,N_8359);
or U8943 (N_8943,N_8424,N_8226);
and U8944 (N_8944,N_8739,N_8710);
and U8945 (N_8945,N_8555,N_8669);
nor U8946 (N_8946,N_8641,N_8326);
and U8947 (N_8947,N_8661,N_8244);
nor U8948 (N_8948,N_8686,N_8549);
xnor U8949 (N_8949,N_8331,N_8219);
and U8950 (N_8950,N_8580,N_8330);
nor U8951 (N_8951,N_8504,N_8189);
and U8952 (N_8952,N_8273,N_8556);
xnor U8953 (N_8953,N_8697,N_8613);
or U8954 (N_8954,N_8204,N_8266);
and U8955 (N_8955,N_8486,N_8155);
xor U8956 (N_8956,N_8614,N_8748);
or U8957 (N_8957,N_8304,N_8432);
xnor U8958 (N_8958,N_8740,N_8245);
nor U8959 (N_8959,N_8709,N_8646);
and U8960 (N_8960,N_8170,N_8324);
or U8961 (N_8961,N_8599,N_8528);
nand U8962 (N_8962,N_8422,N_8335);
nand U8963 (N_8963,N_8242,N_8724);
nand U8964 (N_8964,N_8428,N_8163);
nand U8965 (N_8965,N_8718,N_8635);
nor U8966 (N_8966,N_8416,N_8452);
nor U8967 (N_8967,N_8187,N_8182);
or U8968 (N_8968,N_8489,N_8570);
and U8969 (N_8969,N_8654,N_8540);
or U8970 (N_8970,N_8588,N_8297);
or U8971 (N_8971,N_8205,N_8557);
nand U8972 (N_8972,N_8341,N_8644);
and U8973 (N_8973,N_8383,N_8475);
and U8974 (N_8974,N_8609,N_8746);
xor U8975 (N_8975,N_8514,N_8277);
xor U8976 (N_8976,N_8196,N_8336);
and U8977 (N_8977,N_8637,N_8141);
and U8978 (N_8978,N_8172,N_8308);
or U8979 (N_8979,N_8571,N_8561);
and U8980 (N_8980,N_8197,N_8662);
xnor U8981 (N_8981,N_8433,N_8446);
or U8982 (N_8982,N_8667,N_8224);
or U8983 (N_8983,N_8231,N_8467);
or U8984 (N_8984,N_8511,N_8421);
nor U8985 (N_8985,N_8607,N_8564);
nand U8986 (N_8986,N_8714,N_8657);
and U8987 (N_8987,N_8143,N_8154);
or U8988 (N_8988,N_8684,N_8149);
nand U8989 (N_8989,N_8227,N_8449);
or U8990 (N_8990,N_8640,N_8247);
nor U8991 (N_8991,N_8652,N_8627);
nand U8992 (N_8992,N_8447,N_8368);
and U8993 (N_8993,N_8742,N_8137);
or U8994 (N_8994,N_8472,N_8522);
nor U8995 (N_8995,N_8390,N_8152);
and U8996 (N_8996,N_8579,N_8738);
nand U8997 (N_8997,N_8423,N_8712);
xor U8998 (N_8998,N_8332,N_8216);
nor U8999 (N_8999,N_8743,N_8442);
xor U9000 (N_9000,N_8415,N_8255);
nor U9001 (N_9001,N_8213,N_8544);
xnor U9002 (N_9002,N_8645,N_8310);
xor U9003 (N_9003,N_8309,N_8148);
xnor U9004 (N_9004,N_8348,N_8210);
nand U9005 (N_9005,N_8411,N_8380);
nor U9006 (N_9006,N_8464,N_8575);
or U9007 (N_9007,N_8218,N_8193);
xnor U9008 (N_9008,N_8229,N_8553);
xnor U9009 (N_9009,N_8241,N_8536);
or U9010 (N_9010,N_8236,N_8496);
and U9011 (N_9011,N_8272,N_8279);
or U9012 (N_9012,N_8659,N_8382);
and U9013 (N_9013,N_8365,N_8275);
or U9014 (N_9014,N_8510,N_8441);
and U9015 (N_9015,N_8268,N_8150);
nand U9016 (N_9016,N_8202,N_8687);
nor U9017 (N_9017,N_8457,N_8212);
nand U9018 (N_9018,N_8577,N_8409);
xor U9019 (N_9019,N_8291,N_8320);
or U9020 (N_9020,N_8568,N_8683);
or U9021 (N_9021,N_8593,N_8419);
or U9022 (N_9022,N_8173,N_8180);
nor U9023 (N_9023,N_8174,N_8573);
xnor U9024 (N_9024,N_8610,N_8699);
nor U9025 (N_9025,N_8157,N_8498);
nand U9026 (N_9026,N_8349,N_8127);
or U9027 (N_9027,N_8133,N_8624);
nand U9028 (N_9028,N_8426,N_8636);
xnor U9029 (N_9029,N_8190,N_8650);
nand U9030 (N_9030,N_8541,N_8451);
or U9031 (N_9031,N_8500,N_8397);
xnor U9032 (N_9032,N_8690,N_8306);
xnor U9033 (N_9033,N_8591,N_8325);
nand U9034 (N_9034,N_8410,N_8497);
nor U9035 (N_9035,N_8372,N_8427);
nor U9036 (N_9036,N_8358,N_8545);
nor U9037 (N_9037,N_8253,N_8548);
nor U9038 (N_9038,N_8392,N_8695);
and U9039 (N_9039,N_8565,N_8274);
nand U9040 (N_9040,N_8327,N_8414);
nor U9041 (N_9041,N_8647,N_8400);
nand U9042 (N_9042,N_8162,N_8578);
nor U9043 (N_9043,N_8328,N_8214);
and U9044 (N_9044,N_8319,N_8317);
nand U9045 (N_9045,N_8494,N_8384);
and U9046 (N_9046,N_8388,N_8129);
and U9047 (N_9047,N_8606,N_8139);
nor U9048 (N_9048,N_8166,N_8598);
xor U9049 (N_9049,N_8367,N_8251);
xor U9050 (N_9050,N_8456,N_8265);
xor U9051 (N_9051,N_8271,N_8284);
or U9052 (N_9052,N_8518,N_8629);
nor U9053 (N_9053,N_8431,N_8692);
and U9054 (N_9054,N_8303,N_8530);
and U9055 (N_9055,N_8727,N_8366);
xnor U9056 (N_9056,N_8344,N_8717);
xnor U9057 (N_9057,N_8130,N_8438);
xnor U9058 (N_9058,N_8346,N_8663);
nor U9059 (N_9059,N_8483,N_8198);
or U9060 (N_9060,N_8608,N_8439);
xor U9061 (N_9061,N_8713,N_8417);
and U9062 (N_9062,N_8681,N_8546);
nand U9063 (N_9063,N_8604,N_8485);
or U9064 (N_9064,N_8686,N_8733);
nand U9065 (N_9065,N_8286,N_8378);
nand U9066 (N_9066,N_8261,N_8612);
nor U9067 (N_9067,N_8682,N_8193);
nand U9068 (N_9068,N_8600,N_8204);
and U9069 (N_9069,N_8196,N_8424);
nor U9070 (N_9070,N_8586,N_8196);
or U9071 (N_9071,N_8364,N_8452);
and U9072 (N_9072,N_8211,N_8563);
nand U9073 (N_9073,N_8703,N_8201);
nand U9074 (N_9074,N_8126,N_8573);
xor U9075 (N_9075,N_8494,N_8173);
and U9076 (N_9076,N_8169,N_8730);
xnor U9077 (N_9077,N_8381,N_8322);
xnor U9078 (N_9078,N_8387,N_8141);
or U9079 (N_9079,N_8605,N_8324);
nand U9080 (N_9080,N_8125,N_8499);
and U9081 (N_9081,N_8384,N_8247);
nand U9082 (N_9082,N_8194,N_8490);
nand U9083 (N_9083,N_8377,N_8743);
xor U9084 (N_9084,N_8457,N_8620);
or U9085 (N_9085,N_8153,N_8282);
or U9086 (N_9086,N_8442,N_8518);
nor U9087 (N_9087,N_8696,N_8190);
nand U9088 (N_9088,N_8443,N_8653);
or U9089 (N_9089,N_8341,N_8618);
and U9090 (N_9090,N_8300,N_8293);
nor U9091 (N_9091,N_8315,N_8254);
and U9092 (N_9092,N_8382,N_8371);
and U9093 (N_9093,N_8546,N_8209);
nor U9094 (N_9094,N_8362,N_8300);
and U9095 (N_9095,N_8679,N_8598);
nor U9096 (N_9096,N_8409,N_8155);
xnor U9097 (N_9097,N_8353,N_8575);
xnor U9098 (N_9098,N_8366,N_8289);
and U9099 (N_9099,N_8218,N_8425);
and U9100 (N_9100,N_8473,N_8208);
and U9101 (N_9101,N_8610,N_8706);
and U9102 (N_9102,N_8286,N_8262);
xnor U9103 (N_9103,N_8219,N_8450);
and U9104 (N_9104,N_8395,N_8262);
or U9105 (N_9105,N_8276,N_8614);
or U9106 (N_9106,N_8511,N_8164);
and U9107 (N_9107,N_8135,N_8374);
and U9108 (N_9108,N_8701,N_8498);
or U9109 (N_9109,N_8322,N_8588);
nor U9110 (N_9110,N_8717,N_8611);
nand U9111 (N_9111,N_8406,N_8287);
and U9112 (N_9112,N_8689,N_8278);
or U9113 (N_9113,N_8306,N_8654);
xnor U9114 (N_9114,N_8323,N_8280);
xnor U9115 (N_9115,N_8220,N_8179);
nand U9116 (N_9116,N_8486,N_8293);
and U9117 (N_9117,N_8159,N_8324);
xor U9118 (N_9118,N_8453,N_8657);
and U9119 (N_9119,N_8518,N_8639);
nand U9120 (N_9120,N_8613,N_8641);
nor U9121 (N_9121,N_8614,N_8304);
nor U9122 (N_9122,N_8211,N_8601);
xnor U9123 (N_9123,N_8608,N_8431);
or U9124 (N_9124,N_8486,N_8221);
and U9125 (N_9125,N_8286,N_8242);
nor U9126 (N_9126,N_8215,N_8237);
xor U9127 (N_9127,N_8255,N_8465);
and U9128 (N_9128,N_8339,N_8153);
xor U9129 (N_9129,N_8393,N_8476);
or U9130 (N_9130,N_8560,N_8136);
xor U9131 (N_9131,N_8466,N_8629);
and U9132 (N_9132,N_8680,N_8551);
nand U9133 (N_9133,N_8215,N_8236);
nor U9134 (N_9134,N_8686,N_8644);
or U9135 (N_9135,N_8488,N_8398);
or U9136 (N_9136,N_8317,N_8325);
or U9137 (N_9137,N_8185,N_8384);
xor U9138 (N_9138,N_8174,N_8500);
and U9139 (N_9139,N_8392,N_8201);
or U9140 (N_9140,N_8434,N_8626);
or U9141 (N_9141,N_8207,N_8522);
and U9142 (N_9142,N_8524,N_8288);
xnor U9143 (N_9143,N_8631,N_8412);
nand U9144 (N_9144,N_8498,N_8465);
and U9145 (N_9145,N_8173,N_8206);
and U9146 (N_9146,N_8201,N_8385);
xnor U9147 (N_9147,N_8477,N_8181);
or U9148 (N_9148,N_8426,N_8665);
xnor U9149 (N_9149,N_8743,N_8258);
and U9150 (N_9150,N_8313,N_8180);
nand U9151 (N_9151,N_8206,N_8686);
xor U9152 (N_9152,N_8567,N_8605);
nand U9153 (N_9153,N_8673,N_8157);
and U9154 (N_9154,N_8285,N_8218);
xnor U9155 (N_9155,N_8731,N_8513);
and U9156 (N_9156,N_8411,N_8651);
and U9157 (N_9157,N_8207,N_8576);
xor U9158 (N_9158,N_8321,N_8570);
xnor U9159 (N_9159,N_8621,N_8252);
xnor U9160 (N_9160,N_8353,N_8554);
and U9161 (N_9161,N_8151,N_8177);
nand U9162 (N_9162,N_8296,N_8216);
and U9163 (N_9163,N_8126,N_8721);
or U9164 (N_9164,N_8737,N_8503);
xor U9165 (N_9165,N_8645,N_8609);
nand U9166 (N_9166,N_8251,N_8359);
and U9167 (N_9167,N_8508,N_8670);
nand U9168 (N_9168,N_8226,N_8353);
or U9169 (N_9169,N_8434,N_8333);
and U9170 (N_9170,N_8462,N_8737);
nor U9171 (N_9171,N_8303,N_8386);
xor U9172 (N_9172,N_8463,N_8288);
nand U9173 (N_9173,N_8141,N_8521);
and U9174 (N_9174,N_8335,N_8480);
and U9175 (N_9175,N_8244,N_8577);
nand U9176 (N_9176,N_8510,N_8169);
xnor U9177 (N_9177,N_8167,N_8171);
and U9178 (N_9178,N_8228,N_8643);
and U9179 (N_9179,N_8467,N_8405);
or U9180 (N_9180,N_8254,N_8151);
or U9181 (N_9181,N_8488,N_8687);
and U9182 (N_9182,N_8497,N_8446);
or U9183 (N_9183,N_8162,N_8689);
and U9184 (N_9184,N_8631,N_8701);
and U9185 (N_9185,N_8739,N_8230);
or U9186 (N_9186,N_8570,N_8271);
nor U9187 (N_9187,N_8476,N_8695);
nand U9188 (N_9188,N_8163,N_8636);
and U9189 (N_9189,N_8656,N_8355);
nor U9190 (N_9190,N_8543,N_8156);
nand U9191 (N_9191,N_8707,N_8455);
and U9192 (N_9192,N_8472,N_8223);
nor U9193 (N_9193,N_8655,N_8421);
nor U9194 (N_9194,N_8447,N_8592);
or U9195 (N_9195,N_8576,N_8252);
nand U9196 (N_9196,N_8142,N_8290);
nand U9197 (N_9197,N_8734,N_8559);
nor U9198 (N_9198,N_8331,N_8537);
nand U9199 (N_9199,N_8413,N_8138);
nor U9200 (N_9200,N_8374,N_8550);
or U9201 (N_9201,N_8565,N_8281);
or U9202 (N_9202,N_8742,N_8194);
nor U9203 (N_9203,N_8360,N_8594);
and U9204 (N_9204,N_8641,N_8352);
xor U9205 (N_9205,N_8349,N_8586);
and U9206 (N_9206,N_8362,N_8184);
or U9207 (N_9207,N_8704,N_8256);
nor U9208 (N_9208,N_8237,N_8454);
or U9209 (N_9209,N_8457,N_8401);
nor U9210 (N_9210,N_8309,N_8158);
nand U9211 (N_9211,N_8526,N_8398);
nor U9212 (N_9212,N_8460,N_8616);
nand U9213 (N_9213,N_8233,N_8625);
nand U9214 (N_9214,N_8176,N_8669);
or U9215 (N_9215,N_8736,N_8173);
and U9216 (N_9216,N_8739,N_8486);
nand U9217 (N_9217,N_8611,N_8366);
nand U9218 (N_9218,N_8163,N_8229);
nor U9219 (N_9219,N_8368,N_8525);
xnor U9220 (N_9220,N_8248,N_8695);
or U9221 (N_9221,N_8415,N_8715);
nand U9222 (N_9222,N_8704,N_8485);
nor U9223 (N_9223,N_8389,N_8211);
nand U9224 (N_9224,N_8366,N_8346);
nor U9225 (N_9225,N_8583,N_8522);
and U9226 (N_9226,N_8455,N_8730);
nand U9227 (N_9227,N_8414,N_8182);
and U9228 (N_9228,N_8663,N_8204);
nand U9229 (N_9229,N_8337,N_8147);
and U9230 (N_9230,N_8515,N_8539);
nand U9231 (N_9231,N_8137,N_8700);
xor U9232 (N_9232,N_8635,N_8641);
and U9233 (N_9233,N_8743,N_8364);
nor U9234 (N_9234,N_8551,N_8508);
nand U9235 (N_9235,N_8398,N_8164);
or U9236 (N_9236,N_8278,N_8199);
or U9237 (N_9237,N_8218,N_8568);
nand U9238 (N_9238,N_8597,N_8319);
nand U9239 (N_9239,N_8529,N_8192);
nand U9240 (N_9240,N_8187,N_8473);
or U9241 (N_9241,N_8137,N_8334);
or U9242 (N_9242,N_8246,N_8410);
and U9243 (N_9243,N_8478,N_8405);
or U9244 (N_9244,N_8222,N_8138);
and U9245 (N_9245,N_8188,N_8694);
xor U9246 (N_9246,N_8419,N_8226);
nand U9247 (N_9247,N_8466,N_8535);
and U9248 (N_9248,N_8674,N_8516);
nand U9249 (N_9249,N_8721,N_8551);
and U9250 (N_9250,N_8586,N_8180);
nor U9251 (N_9251,N_8317,N_8381);
xor U9252 (N_9252,N_8274,N_8735);
or U9253 (N_9253,N_8652,N_8488);
xnor U9254 (N_9254,N_8621,N_8604);
nor U9255 (N_9255,N_8307,N_8278);
or U9256 (N_9256,N_8595,N_8249);
nand U9257 (N_9257,N_8462,N_8264);
nand U9258 (N_9258,N_8166,N_8407);
xnor U9259 (N_9259,N_8737,N_8468);
nand U9260 (N_9260,N_8512,N_8722);
xnor U9261 (N_9261,N_8312,N_8474);
and U9262 (N_9262,N_8637,N_8327);
xor U9263 (N_9263,N_8297,N_8138);
xnor U9264 (N_9264,N_8344,N_8622);
nand U9265 (N_9265,N_8226,N_8429);
and U9266 (N_9266,N_8718,N_8390);
or U9267 (N_9267,N_8488,N_8749);
nand U9268 (N_9268,N_8553,N_8389);
xnor U9269 (N_9269,N_8187,N_8638);
xor U9270 (N_9270,N_8301,N_8509);
or U9271 (N_9271,N_8179,N_8128);
nand U9272 (N_9272,N_8681,N_8250);
nand U9273 (N_9273,N_8414,N_8299);
nand U9274 (N_9274,N_8207,N_8624);
nand U9275 (N_9275,N_8383,N_8148);
and U9276 (N_9276,N_8749,N_8609);
nand U9277 (N_9277,N_8589,N_8196);
nor U9278 (N_9278,N_8744,N_8458);
nor U9279 (N_9279,N_8156,N_8600);
nor U9280 (N_9280,N_8142,N_8522);
nor U9281 (N_9281,N_8180,N_8129);
and U9282 (N_9282,N_8740,N_8405);
or U9283 (N_9283,N_8414,N_8497);
xnor U9284 (N_9284,N_8503,N_8323);
nor U9285 (N_9285,N_8634,N_8329);
xnor U9286 (N_9286,N_8645,N_8615);
nand U9287 (N_9287,N_8489,N_8606);
or U9288 (N_9288,N_8608,N_8536);
or U9289 (N_9289,N_8657,N_8717);
and U9290 (N_9290,N_8428,N_8518);
xnor U9291 (N_9291,N_8668,N_8468);
xor U9292 (N_9292,N_8586,N_8450);
xnor U9293 (N_9293,N_8691,N_8470);
xnor U9294 (N_9294,N_8235,N_8424);
or U9295 (N_9295,N_8382,N_8127);
and U9296 (N_9296,N_8692,N_8604);
xnor U9297 (N_9297,N_8505,N_8331);
and U9298 (N_9298,N_8471,N_8684);
nand U9299 (N_9299,N_8313,N_8418);
and U9300 (N_9300,N_8402,N_8699);
nand U9301 (N_9301,N_8319,N_8397);
nor U9302 (N_9302,N_8177,N_8325);
and U9303 (N_9303,N_8712,N_8278);
nor U9304 (N_9304,N_8541,N_8623);
or U9305 (N_9305,N_8596,N_8234);
nor U9306 (N_9306,N_8550,N_8577);
nand U9307 (N_9307,N_8249,N_8341);
nand U9308 (N_9308,N_8206,N_8158);
nand U9309 (N_9309,N_8272,N_8384);
nor U9310 (N_9310,N_8642,N_8220);
xor U9311 (N_9311,N_8734,N_8642);
nor U9312 (N_9312,N_8744,N_8461);
nand U9313 (N_9313,N_8681,N_8655);
or U9314 (N_9314,N_8674,N_8696);
nor U9315 (N_9315,N_8733,N_8341);
and U9316 (N_9316,N_8235,N_8223);
and U9317 (N_9317,N_8674,N_8366);
and U9318 (N_9318,N_8479,N_8135);
nor U9319 (N_9319,N_8179,N_8515);
nor U9320 (N_9320,N_8417,N_8210);
xnor U9321 (N_9321,N_8493,N_8169);
nand U9322 (N_9322,N_8383,N_8167);
nand U9323 (N_9323,N_8641,N_8575);
nor U9324 (N_9324,N_8422,N_8612);
nand U9325 (N_9325,N_8520,N_8333);
nand U9326 (N_9326,N_8314,N_8217);
or U9327 (N_9327,N_8393,N_8472);
or U9328 (N_9328,N_8469,N_8368);
nor U9329 (N_9329,N_8387,N_8408);
xor U9330 (N_9330,N_8642,N_8428);
and U9331 (N_9331,N_8258,N_8566);
and U9332 (N_9332,N_8204,N_8456);
or U9333 (N_9333,N_8675,N_8653);
xnor U9334 (N_9334,N_8389,N_8735);
or U9335 (N_9335,N_8508,N_8245);
nand U9336 (N_9336,N_8143,N_8263);
nand U9337 (N_9337,N_8260,N_8475);
and U9338 (N_9338,N_8212,N_8564);
nand U9339 (N_9339,N_8165,N_8351);
nor U9340 (N_9340,N_8549,N_8191);
nor U9341 (N_9341,N_8285,N_8307);
nand U9342 (N_9342,N_8558,N_8160);
xor U9343 (N_9343,N_8127,N_8283);
xnor U9344 (N_9344,N_8607,N_8257);
or U9345 (N_9345,N_8148,N_8642);
nor U9346 (N_9346,N_8331,N_8530);
or U9347 (N_9347,N_8490,N_8193);
or U9348 (N_9348,N_8229,N_8156);
xor U9349 (N_9349,N_8229,N_8263);
or U9350 (N_9350,N_8625,N_8133);
nand U9351 (N_9351,N_8581,N_8152);
nand U9352 (N_9352,N_8216,N_8713);
nand U9353 (N_9353,N_8217,N_8613);
or U9354 (N_9354,N_8621,N_8262);
nand U9355 (N_9355,N_8197,N_8183);
nand U9356 (N_9356,N_8712,N_8215);
nand U9357 (N_9357,N_8379,N_8453);
or U9358 (N_9358,N_8632,N_8409);
and U9359 (N_9359,N_8445,N_8578);
or U9360 (N_9360,N_8252,N_8450);
nor U9361 (N_9361,N_8583,N_8731);
nand U9362 (N_9362,N_8493,N_8172);
nand U9363 (N_9363,N_8156,N_8464);
xor U9364 (N_9364,N_8137,N_8267);
xor U9365 (N_9365,N_8522,N_8382);
and U9366 (N_9366,N_8340,N_8728);
xor U9367 (N_9367,N_8205,N_8130);
xnor U9368 (N_9368,N_8132,N_8208);
xnor U9369 (N_9369,N_8425,N_8382);
xor U9370 (N_9370,N_8349,N_8534);
or U9371 (N_9371,N_8567,N_8187);
nor U9372 (N_9372,N_8218,N_8275);
and U9373 (N_9373,N_8188,N_8475);
nand U9374 (N_9374,N_8152,N_8517);
nand U9375 (N_9375,N_9081,N_9204);
nor U9376 (N_9376,N_9140,N_9163);
xnor U9377 (N_9377,N_8927,N_9214);
nor U9378 (N_9378,N_9281,N_8880);
nand U9379 (N_9379,N_8819,N_8989);
nand U9380 (N_9380,N_8978,N_8957);
nor U9381 (N_9381,N_9271,N_9217);
or U9382 (N_9382,N_9187,N_9000);
xnor U9383 (N_9383,N_8904,N_9199);
nand U9384 (N_9384,N_9086,N_8785);
and U9385 (N_9385,N_8805,N_8853);
nand U9386 (N_9386,N_8921,N_9111);
or U9387 (N_9387,N_9243,N_9269);
nand U9388 (N_9388,N_9312,N_9331);
nor U9389 (N_9389,N_8808,N_9150);
and U9390 (N_9390,N_9161,N_9309);
nand U9391 (N_9391,N_9236,N_9045);
or U9392 (N_9392,N_8831,N_8983);
nand U9393 (N_9393,N_9014,N_8855);
and U9394 (N_9394,N_9127,N_8856);
or U9395 (N_9395,N_8999,N_8789);
nand U9396 (N_9396,N_9042,N_8824);
or U9397 (N_9397,N_9213,N_9030);
and U9398 (N_9398,N_8851,N_9036);
xor U9399 (N_9399,N_9316,N_9003);
nor U9400 (N_9400,N_9273,N_9361);
nand U9401 (N_9401,N_9137,N_9308);
nor U9402 (N_9402,N_9135,N_9118);
and U9403 (N_9403,N_9097,N_9073);
xnor U9404 (N_9404,N_9034,N_9181);
xnor U9405 (N_9405,N_8770,N_9363);
and U9406 (N_9406,N_9099,N_8766);
xnor U9407 (N_9407,N_9178,N_8798);
and U9408 (N_9408,N_9151,N_8875);
nor U9409 (N_9409,N_9223,N_8771);
or U9410 (N_9410,N_8852,N_9136);
xor U9411 (N_9411,N_9301,N_9225);
xnor U9412 (N_9412,N_8950,N_9292);
nand U9413 (N_9413,N_8833,N_9129);
xnor U9414 (N_9414,N_8937,N_9249);
nor U9415 (N_9415,N_9252,N_9145);
xor U9416 (N_9416,N_9044,N_8991);
nor U9417 (N_9417,N_8759,N_9186);
or U9418 (N_9418,N_8810,N_9173);
nor U9419 (N_9419,N_9205,N_9152);
and U9420 (N_9420,N_9355,N_8912);
and U9421 (N_9421,N_9048,N_9267);
nand U9422 (N_9422,N_8839,N_9371);
nor U9423 (N_9423,N_8962,N_8955);
and U9424 (N_9424,N_9015,N_9246);
xor U9425 (N_9425,N_8891,N_9056);
nor U9426 (N_9426,N_9133,N_9191);
nor U9427 (N_9427,N_9041,N_9114);
xnor U9428 (N_9428,N_8760,N_8972);
nor U9429 (N_9429,N_9296,N_9354);
nand U9430 (N_9430,N_8842,N_8933);
or U9431 (N_9431,N_9218,N_9280);
nand U9432 (N_9432,N_8920,N_8821);
or U9433 (N_9433,N_8823,N_9113);
nand U9434 (N_9434,N_9166,N_8879);
or U9435 (N_9435,N_9033,N_9234);
nand U9436 (N_9436,N_9294,N_8985);
nor U9437 (N_9437,N_9046,N_8848);
or U9438 (N_9438,N_9334,N_9244);
xnor U9439 (N_9439,N_9324,N_8783);
xnor U9440 (N_9440,N_9260,N_9126);
nor U9441 (N_9441,N_8870,N_9195);
and U9442 (N_9442,N_9369,N_9220);
and U9443 (N_9443,N_8996,N_9255);
nor U9444 (N_9444,N_9071,N_8815);
nor U9445 (N_9445,N_8750,N_9117);
nor U9446 (N_9446,N_9277,N_9091);
or U9447 (N_9447,N_9125,N_9289);
xor U9448 (N_9448,N_9122,N_8993);
and U9449 (N_9449,N_9050,N_9291);
xnor U9450 (N_9450,N_9184,N_8900);
or U9451 (N_9451,N_9176,N_9356);
nand U9452 (N_9452,N_9028,N_9343);
and U9453 (N_9453,N_8780,N_9158);
and U9454 (N_9454,N_9227,N_8782);
xnor U9455 (N_9455,N_8915,N_8752);
or U9456 (N_9456,N_9007,N_8887);
or U9457 (N_9457,N_8896,N_8938);
nand U9458 (N_9458,N_9333,N_8832);
or U9459 (N_9459,N_9221,N_9266);
and U9460 (N_9460,N_9077,N_8926);
nor U9461 (N_9461,N_8930,N_9327);
or U9462 (N_9462,N_8894,N_9299);
or U9463 (N_9463,N_8994,N_8943);
and U9464 (N_9464,N_9265,N_9337);
nor U9465 (N_9465,N_8992,N_9237);
xor U9466 (N_9466,N_8923,N_9283);
nor U9467 (N_9467,N_9105,N_9175);
and U9468 (N_9468,N_9314,N_9310);
xor U9469 (N_9469,N_9021,N_8885);
xnor U9470 (N_9470,N_9057,N_9123);
xnor U9471 (N_9471,N_8827,N_9180);
nand U9472 (N_9472,N_8997,N_9206);
and U9473 (N_9473,N_8814,N_8778);
and U9474 (N_9474,N_8917,N_9160);
or U9475 (N_9475,N_9018,N_9116);
nand U9476 (N_9476,N_9222,N_8871);
or U9477 (N_9477,N_9079,N_9274);
xor U9478 (N_9478,N_8939,N_9335);
nor U9479 (N_9479,N_9275,N_8850);
and U9480 (N_9480,N_9035,N_9229);
nor U9481 (N_9481,N_9322,N_8948);
or U9482 (N_9482,N_8807,N_8854);
or U9483 (N_9483,N_9104,N_9124);
or U9484 (N_9484,N_9142,N_9263);
or U9485 (N_9485,N_9303,N_8818);
nor U9486 (N_9486,N_8811,N_8998);
nor U9487 (N_9487,N_9287,N_8784);
xor U9488 (N_9488,N_8794,N_9169);
xor U9489 (N_9489,N_9276,N_9272);
nor U9490 (N_9490,N_9211,N_8932);
or U9491 (N_9491,N_9207,N_9072);
xnor U9492 (N_9492,N_8906,N_9149);
and U9493 (N_9493,N_9132,N_8796);
or U9494 (N_9494,N_8756,N_8835);
nor U9495 (N_9495,N_8960,N_8914);
and U9496 (N_9496,N_9366,N_8940);
nand U9497 (N_9497,N_9242,N_8929);
nand U9498 (N_9498,N_9198,N_8988);
nand U9499 (N_9499,N_8990,N_9188);
and U9500 (N_9500,N_9351,N_9082);
or U9501 (N_9501,N_8909,N_9216);
xor U9502 (N_9502,N_9112,N_8864);
nand U9503 (N_9503,N_8956,N_9304);
nor U9504 (N_9504,N_8869,N_9202);
nor U9505 (N_9505,N_9367,N_9193);
nand U9506 (N_9506,N_9031,N_9154);
nor U9507 (N_9507,N_8764,N_9254);
xnor U9508 (N_9508,N_8874,N_8945);
nand U9509 (N_9509,N_9360,N_9010);
and U9510 (N_9510,N_9182,N_9087);
nor U9511 (N_9511,N_9336,N_8883);
nand U9512 (N_9512,N_8973,N_8795);
xnor U9513 (N_9513,N_8986,N_9319);
nand U9514 (N_9514,N_9006,N_8836);
or U9515 (N_9515,N_8858,N_9102);
nor U9516 (N_9516,N_9352,N_9159);
and U9517 (N_9517,N_8754,N_9059);
xor U9518 (N_9518,N_9330,N_8918);
nand U9519 (N_9519,N_9210,N_8892);
nand U9520 (N_9520,N_9053,N_9247);
nor U9521 (N_9521,N_8788,N_9374);
nor U9522 (N_9522,N_9344,N_8843);
nand U9523 (N_9523,N_9239,N_8895);
or U9524 (N_9524,N_8804,N_8862);
or U9525 (N_9525,N_9295,N_9224);
nor U9526 (N_9526,N_9095,N_9016);
nor U9527 (N_9527,N_8898,N_9253);
nor U9528 (N_9528,N_9325,N_9342);
and U9529 (N_9529,N_8758,N_8897);
or U9530 (N_9530,N_8961,N_8838);
nor U9531 (N_9531,N_9096,N_8905);
nor U9532 (N_9532,N_9088,N_9185);
nand U9533 (N_9533,N_9215,N_9108);
xor U9534 (N_9534,N_8817,N_9305);
xnor U9535 (N_9535,N_9005,N_9085);
nor U9536 (N_9536,N_9162,N_9084);
nand U9537 (N_9537,N_9340,N_9212);
or U9538 (N_9538,N_9144,N_8801);
and U9539 (N_9539,N_8888,N_8834);
nand U9540 (N_9540,N_9139,N_9128);
xor U9541 (N_9541,N_8837,N_9120);
nor U9542 (N_9542,N_8882,N_9062);
or U9543 (N_9543,N_9165,N_8790);
and U9544 (N_9544,N_9228,N_9157);
or U9545 (N_9545,N_8901,N_8775);
or U9546 (N_9546,N_8907,N_8865);
nor U9547 (N_9547,N_9089,N_8952);
xor U9548 (N_9548,N_8859,N_9365);
or U9549 (N_9549,N_9231,N_9232);
nand U9550 (N_9550,N_9256,N_8987);
and U9551 (N_9551,N_9285,N_9092);
xor U9552 (N_9552,N_9370,N_8968);
nor U9553 (N_9553,N_9315,N_8868);
xor U9554 (N_9554,N_8820,N_9359);
xnor U9555 (N_9555,N_8773,N_9038);
and U9556 (N_9556,N_8899,N_9338);
xnor U9557 (N_9557,N_9197,N_8800);
and U9558 (N_9558,N_8916,N_9290);
and U9559 (N_9559,N_9037,N_8840);
nand U9560 (N_9560,N_9268,N_9278);
xnor U9561 (N_9561,N_9208,N_9357);
and U9562 (N_9562,N_9172,N_8846);
or U9563 (N_9563,N_8867,N_8942);
nor U9564 (N_9564,N_9284,N_9013);
and U9565 (N_9565,N_8826,N_8951);
xor U9566 (N_9566,N_9238,N_9098);
nand U9567 (N_9567,N_9320,N_9350);
nor U9568 (N_9568,N_8753,N_8911);
and U9569 (N_9569,N_9115,N_8975);
and U9570 (N_9570,N_9029,N_8762);
or U9571 (N_9571,N_9332,N_9282);
xor U9572 (N_9572,N_9347,N_8779);
and U9573 (N_9573,N_9027,N_8792);
or U9574 (N_9574,N_9100,N_8847);
nand U9575 (N_9575,N_9341,N_9307);
and U9576 (N_9576,N_8936,N_9131);
xor U9577 (N_9577,N_8849,N_8893);
and U9578 (N_9578,N_8763,N_8980);
or U9579 (N_9579,N_9022,N_9090);
or U9580 (N_9580,N_8953,N_9194);
nor U9581 (N_9581,N_9233,N_9051);
nor U9582 (N_9582,N_9040,N_8949);
xor U9583 (N_9583,N_9043,N_8866);
or U9584 (N_9584,N_8844,N_9329);
or U9585 (N_9585,N_8787,N_9372);
and U9586 (N_9586,N_8863,N_8772);
nor U9587 (N_9587,N_9047,N_9058);
and U9588 (N_9588,N_9346,N_9349);
xor U9589 (N_9589,N_9201,N_8816);
nor U9590 (N_9590,N_9001,N_9074);
nor U9591 (N_9591,N_8793,N_8889);
nand U9592 (N_9592,N_8995,N_9317);
nor U9593 (N_9593,N_9004,N_8884);
nor U9594 (N_9594,N_9203,N_9261);
nand U9595 (N_9595,N_8967,N_8876);
nand U9596 (N_9596,N_9270,N_9017);
nand U9597 (N_9597,N_8881,N_8913);
nand U9598 (N_9598,N_9147,N_9002);
xnor U9599 (N_9599,N_9302,N_8931);
or U9600 (N_9600,N_9311,N_8928);
nor U9601 (N_9601,N_8769,N_9313);
xor U9602 (N_9602,N_8860,N_9138);
nor U9603 (N_9603,N_9141,N_9192);
nor U9604 (N_9604,N_9298,N_9323);
xor U9605 (N_9605,N_8971,N_9107);
nand U9606 (N_9606,N_9300,N_9251);
xnor U9607 (N_9607,N_9258,N_9064);
and U9608 (N_9608,N_9143,N_8755);
nor U9609 (N_9609,N_9167,N_8802);
and U9610 (N_9610,N_9094,N_9293);
and U9611 (N_9611,N_9297,N_9121);
or U9612 (N_9612,N_9235,N_9068);
and U9613 (N_9613,N_9326,N_9364);
xor U9614 (N_9614,N_9262,N_8902);
nor U9615 (N_9615,N_8776,N_8878);
nand U9616 (N_9616,N_8828,N_9019);
xor U9617 (N_9617,N_8829,N_9358);
or U9618 (N_9618,N_9103,N_8944);
nor U9619 (N_9619,N_9279,N_9240);
and U9620 (N_9620,N_9009,N_8903);
nand U9621 (N_9621,N_8922,N_8774);
and U9622 (N_9622,N_9339,N_9134);
xor U9623 (N_9623,N_8803,N_9230);
or U9624 (N_9624,N_8768,N_9259);
nor U9625 (N_9625,N_8965,N_8791);
and U9626 (N_9626,N_8924,N_8761);
and U9627 (N_9627,N_9170,N_9171);
nand U9628 (N_9628,N_9101,N_9264);
nor U9629 (N_9629,N_9373,N_8857);
and U9630 (N_9630,N_8925,N_9250);
or U9631 (N_9631,N_9226,N_9368);
xnor U9632 (N_9632,N_9196,N_8935);
or U9633 (N_9633,N_9061,N_9008);
or U9634 (N_9634,N_9164,N_9023);
nor U9635 (N_9635,N_8958,N_8841);
or U9636 (N_9636,N_8812,N_8877);
nor U9637 (N_9637,N_8830,N_9076);
xnor U9638 (N_9638,N_8934,N_8977);
nor U9639 (N_9639,N_9110,N_9248);
or U9640 (N_9640,N_9179,N_8777);
nor U9641 (N_9641,N_9183,N_8799);
and U9642 (N_9642,N_9348,N_9190);
nor U9643 (N_9643,N_8765,N_9054);
and U9644 (N_9644,N_8966,N_9321);
nand U9645 (N_9645,N_8982,N_8969);
nand U9646 (N_9646,N_9065,N_8974);
xnor U9647 (N_9647,N_9109,N_9024);
and U9648 (N_9648,N_9012,N_8984);
xnor U9649 (N_9649,N_8964,N_9328);
or U9650 (N_9650,N_9168,N_8781);
or U9651 (N_9651,N_9011,N_8947);
and U9652 (N_9652,N_9055,N_8910);
and U9653 (N_9653,N_9070,N_9075);
and U9654 (N_9654,N_9306,N_8872);
xor U9655 (N_9655,N_9245,N_8786);
xor U9656 (N_9656,N_9318,N_8979);
and U9657 (N_9657,N_8886,N_9052);
nand U9658 (N_9658,N_8861,N_9069);
nor U9659 (N_9659,N_8941,N_9288);
or U9660 (N_9660,N_9153,N_8890);
nand U9661 (N_9661,N_9080,N_8970);
and U9662 (N_9662,N_9020,N_8919);
or U9663 (N_9663,N_9067,N_9093);
and U9664 (N_9664,N_8813,N_8845);
nand U9665 (N_9665,N_9119,N_9146);
or U9666 (N_9666,N_9362,N_9200);
xor U9667 (N_9667,N_9066,N_9345);
or U9668 (N_9668,N_9155,N_9060);
nor U9669 (N_9669,N_9049,N_8963);
nand U9670 (N_9670,N_9032,N_9130);
nor U9671 (N_9671,N_8797,N_9025);
nor U9672 (N_9672,N_9286,N_8976);
xnor U9673 (N_9673,N_8822,N_9078);
and U9674 (N_9674,N_9257,N_8981);
and U9675 (N_9675,N_9039,N_9174);
or U9676 (N_9676,N_9353,N_8825);
or U9677 (N_9677,N_8767,N_9083);
and U9678 (N_9678,N_9063,N_9156);
nand U9679 (N_9679,N_9219,N_8954);
nor U9680 (N_9680,N_9106,N_8908);
or U9681 (N_9681,N_9177,N_8959);
xnor U9682 (N_9682,N_9189,N_8873);
nor U9683 (N_9683,N_8809,N_8946);
or U9684 (N_9684,N_9241,N_8806);
or U9685 (N_9685,N_8757,N_9209);
and U9686 (N_9686,N_8751,N_9148);
nor U9687 (N_9687,N_9026,N_8807);
or U9688 (N_9688,N_9224,N_9017);
nor U9689 (N_9689,N_9334,N_8948);
xor U9690 (N_9690,N_9226,N_9022);
or U9691 (N_9691,N_8828,N_9281);
or U9692 (N_9692,N_9144,N_9278);
nor U9693 (N_9693,N_9049,N_8775);
xnor U9694 (N_9694,N_9215,N_9030);
xor U9695 (N_9695,N_8982,N_9356);
xor U9696 (N_9696,N_8914,N_8974);
nor U9697 (N_9697,N_9325,N_9012);
nand U9698 (N_9698,N_9331,N_9107);
nor U9699 (N_9699,N_8782,N_9078);
nor U9700 (N_9700,N_8777,N_9214);
or U9701 (N_9701,N_8852,N_9189);
and U9702 (N_9702,N_8886,N_9292);
xnor U9703 (N_9703,N_9113,N_9149);
xor U9704 (N_9704,N_9178,N_9187);
and U9705 (N_9705,N_8833,N_8924);
xor U9706 (N_9706,N_9326,N_8785);
nand U9707 (N_9707,N_8879,N_9340);
and U9708 (N_9708,N_8943,N_9335);
or U9709 (N_9709,N_8965,N_9200);
nor U9710 (N_9710,N_8955,N_9001);
and U9711 (N_9711,N_8818,N_9021);
or U9712 (N_9712,N_8964,N_9365);
nor U9713 (N_9713,N_8753,N_8898);
and U9714 (N_9714,N_8803,N_8833);
nand U9715 (N_9715,N_9075,N_9184);
xor U9716 (N_9716,N_8809,N_9160);
xnor U9717 (N_9717,N_9203,N_9106);
xor U9718 (N_9718,N_8804,N_9091);
nor U9719 (N_9719,N_9370,N_9097);
nor U9720 (N_9720,N_9098,N_8777);
nor U9721 (N_9721,N_8971,N_9114);
and U9722 (N_9722,N_9321,N_9119);
and U9723 (N_9723,N_9313,N_9083);
nor U9724 (N_9724,N_9035,N_8997);
and U9725 (N_9725,N_8799,N_9275);
nand U9726 (N_9726,N_9228,N_8912);
xnor U9727 (N_9727,N_8777,N_8750);
nor U9728 (N_9728,N_8900,N_8916);
nand U9729 (N_9729,N_9055,N_9294);
and U9730 (N_9730,N_8821,N_9281);
and U9731 (N_9731,N_8832,N_8998);
nor U9732 (N_9732,N_9121,N_9253);
and U9733 (N_9733,N_8990,N_8754);
and U9734 (N_9734,N_8941,N_9268);
or U9735 (N_9735,N_8893,N_8964);
or U9736 (N_9736,N_9113,N_8885);
xnor U9737 (N_9737,N_8830,N_9152);
nor U9738 (N_9738,N_8838,N_8992);
xor U9739 (N_9739,N_9346,N_9344);
nand U9740 (N_9740,N_8959,N_8972);
and U9741 (N_9741,N_9095,N_9017);
and U9742 (N_9742,N_9087,N_8947);
and U9743 (N_9743,N_9307,N_8876);
xor U9744 (N_9744,N_8809,N_9211);
xor U9745 (N_9745,N_8813,N_9262);
and U9746 (N_9746,N_9019,N_9145);
or U9747 (N_9747,N_9290,N_8850);
or U9748 (N_9748,N_8920,N_8795);
nor U9749 (N_9749,N_8775,N_9027);
nor U9750 (N_9750,N_9072,N_8937);
nor U9751 (N_9751,N_9002,N_8916);
xnor U9752 (N_9752,N_8939,N_9098);
and U9753 (N_9753,N_9292,N_9113);
or U9754 (N_9754,N_8775,N_8875);
nor U9755 (N_9755,N_9225,N_9278);
or U9756 (N_9756,N_8837,N_8929);
nor U9757 (N_9757,N_9268,N_9318);
and U9758 (N_9758,N_9045,N_9223);
or U9759 (N_9759,N_8835,N_9147);
nor U9760 (N_9760,N_9143,N_8823);
nand U9761 (N_9761,N_8853,N_9130);
and U9762 (N_9762,N_8942,N_8843);
and U9763 (N_9763,N_9200,N_8960);
xor U9764 (N_9764,N_8839,N_9012);
or U9765 (N_9765,N_9062,N_9092);
and U9766 (N_9766,N_9195,N_9197);
nand U9767 (N_9767,N_9002,N_9155);
nor U9768 (N_9768,N_8914,N_8900);
nor U9769 (N_9769,N_9306,N_9370);
and U9770 (N_9770,N_9258,N_9132);
xnor U9771 (N_9771,N_9056,N_9341);
or U9772 (N_9772,N_8869,N_8972);
or U9773 (N_9773,N_8810,N_9100);
xor U9774 (N_9774,N_8897,N_9245);
and U9775 (N_9775,N_9044,N_8971);
or U9776 (N_9776,N_8925,N_8872);
and U9777 (N_9777,N_9259,N_8982);
nand U9778 (N_9778,N_9198,N_9190);
nor U9779 (N_9779,N_9308,N_9082);
or U9780 (N_9780,N_8959,N_8792);
and U9781 (N_9781,N_9152,N_9019);
or U9782 (N_9782,N_8993,N_9240);
xor U9783 (N_9783,N_9354,N_9224);
or U9784 (N_9784,N_9073,N_9127);
and U9785 (N_9785,N_9174,N_8912);
and U9786 (N_9786,N_9112,N_9097);
nor U9787 (N_9787,N_8938,N_8998);
xnor U9788 (N_9788,N_9130,N_9312);
nor U9789 (N_9789,N_8875,N_9101);
and U9790 (N_9790,N_8802,N_8751);
nand U9791 (N_9791,N_9154,N_8957);
nor U9792 (N_9792,N_9245,N_9182);
and U9793 (N_9793,N_9105,N_8950);
or U9794 (N_9794,N_9232,N_8808);
xnor U9795 (N_9795,N_8794,N_9156);
or U9796 (N_9796,N_9191,N_9005);
xnor U9797 (N_9797,N_8786,N_9116);
nor U9798 (N_9798,N_9307,N_9373);
nor U9799 (N_9799,N_8977,N_9281);
or U9800 (N_9800,N_9246,N_8976);
xor U9801 (N_9801,N_9080,N_8973);
nor U9802 (N_9802,N_9163,N_9109);
or U9803 (N_9803,N_9233,N_9166);
nor U9804 (N_9804,N_9081,N_9271);
xnor U9805 (N_9805,N_8811,N_8992);
and U9806 (N_9806,N_9127,N_9342);
or U9807 (N_9807,N_9181,N_8973);
xnor U9808 (N_9808,N_8909,N_8973);
and U9809 (N_9809,N_9235,N_9345);
xnor U9810 (N_9810,N_9020,N_8965);
xor U9811 (N_9811,N_9062,N_8952);
nor U9812 (N_9812,N_9231,N_9130);
nor U9813 (N_9813,N_9157,N_8860);
and U9814 (N_9814,N_9030,N_9192);
xor U9815 (N_9815,N_8798,N_8857);
nor U9816 (N_9816,N_8928,N_8788);
and U9817 (N_9817,N_9326,N_9208);
and U9818 (N_9818,N_9320,N_8829);
and U9819 (N_9819,N_9252,N_8888);
or U9820 (N_9820,N_8997,N_9069);
xor U9821 (N_9821,N_8815,N_9147);
nor U9822 (N_9822,N_9246,N_9175);
and U9823 (N_9823,N_9266,N_8898);
nand U9824 (N_9824,N_9333,N_9326);
and U9825 (N_9825,N_9227,N_9297);
nor U9826 (N_9826,N_9256,N_8757);
xor U9827 (N_9827,N_9233,N_9068);
xor U9828 (N_9828,N_9058,N_9289);
xor U9829 (N_9829,N_8785,N_9014);
nor U9830 (N_9830,N_8832,N_9131);
nand U9831 (N_9831,N_8914,N_9064);
nor U9832 (N_9832,N_8838,N_9365);
or U9833 (N_9833,N_9329,N_9020);
and U9834 (N_9834,N_8809,N_8938);
or U9835 (N_9835,N_8830,N_8829);
nand U9836 (N_9836,N_8776,N_9302);
xnor U9837 (N_9837,N_9232,N_9096);
xor U9838 (N_9838,N_9246,N_8876);
and U9839 (N_9839,N_9082,N_9056);
nand U9840 (N_9840,N_9010,N_9334);
nand U9841 (N_9841,N_9100,N_9120);
xor U9842 (N_9842,N_8844,N_9369);
xnor U9843 (N_9843,N_8776,N_8962);
xor U9844 (N_9844,N_8843,N_9094);
xor U9845 (N_9845,N_9124,N_9076);
nand U9846 (N_9846,N_8905,N_9068);
or U9847 (N_9847,N_9348,N_9125);
and U9848 (N_9848,N_9353,N_8802);
nand U9849 (N_9849,N_8961,N_9158);
or U9850 (N_9850,N_8993,N_9226);
nor U9851 (N_9851,N_9034,N_9355);
or U9852 (N_9852,N_8822,N_8889);
nor U9853 (N_9853,N_8784,N_8865);
or U9854 (N_9854,N_8826,N_9001);
or U9855 (N_9855,N_9109,N_9198);
nor U9856 (N_9856,N_8818,N_9358);
xnor U9857 (N_9857,N_9294,N_9251);
xor U9858 (N_9858,N_8824,N_9151);
and U9859 (N_9859,N_8756,N_9132);
xnor U9860 (N_9860,N_8880,N_8903);
or U9861 (N_9861,N_8833,N_9161);
nor U9862 (N_9862,N_8945,N_9037);
nor U9863 (N_9863,N_8827,N_8879);
nand U9864 (N_9864,N_8828,N_9282);
and U9865 (N_9865,N_8750,N_8896);
nor U9866 (N_9866,N_8906,N_8771);
and U9867 (N_9867,N_9152,N_9090);
nand U9868 (N_9868,N_8858,N_9056);
nor U9869 (N_9869,N_9282,N_9015);
nand U9870 (N_9870,N_8824,N_8964);
nand U9871 (N_9871,N_8755,N_9067);
xor U9872 (N_9872,N_9365,N_9025);
nand U9873 (N_9873,N_9052,N_9182);
xnor U9874 (N_9874,N_9135,N_8894);
and U9875 (N_9875,N_8955,N_8895);
or U9876 (N_9876,N_9061,N_8818);
or U9877 (N_9877,N_9273,N_9321);
nor U9878 (N_9878,N_9171,N_8952);
and U9879 (N_9879,N_8946,N_9110);
or U9880 (N_9880,N_9259,N_9060);
or U9881 (N_9881,N_9140,N_9038);
xor U9882 (N_9882,N_8964,N_9054);
nand U9883 (N_9883,N_8889,N_9341);
or U9884 (N_9884,N_9182,N_9121);
nor U9885 (N_9885,N_9126,N_9165);
xnor U9886 (N_9886,N_9083,N_8879);
nand U9887 (N_9887,N_8916,N_8845);
and U9888 (N_9888,N_8786,N_9011);
nor U9889 (N_9889,N_8787,N_9101);
and U9890 (N_9890,N_9365,N_9166);
nand U9891 (N_9891,N_9240,N_8965);
nand U9892 (N_9892,N_8948,N_9283);
or U9893 (N_9893,N_8868,N_9150);
nand U9894 (N_9894,N_8767,N_9080);
xnor U9895 (N_9895,N_9076,N_9083);
or U9896 (N_9896,N_9085,N_9247);
xnor U9897 (N_9897,N_8884,N_9070);
xnor U9898 (N_9898,N_8937,N_8900);
nor U9899 (N_9899,N_8813,N_8781);
or U9900 (N_9900,N_8807,N_9110);
and U9901 (N_9901,N_8805,N_9139);
or U9902 (N_9902,N_9012,N_9022);
nor U9903 (N_9903,N_8896,N_9110);
nor U9904 (N_9904,N_9240,N_8903);
xnor U9905 (N_9905,N_9169,N_9203);
nor U9906 (N_9906,N_9349,N_9072);
nor U9907 (N_9907,N_9280,N_8993);
nor U9908 (N_9908,N_9108,N_9332);
xor U9909 (N_9909,N_9218,N_8955);
xor U9910 (N_9910,N_8858,N_8780);
or U9911 (N_9911,N_9325,N_8936);
nand U9912 (N_9912,N_8794,N_8913);
nor U9913 (N_9913,N_8902,N_8949);
or U9914 (N_9914,N_9147,N_8935);
nand U9915 (N_9915,N_8851,N_9277);
or U9916 (N_9916,N_8757,N_8802);
or U9917 (N_9917,N_9035,N_9209);
and U9918 (N_9918,N_8910,N_9295);
nor U9919 (N_9919,N_9210,N_9111);
xnor U9920 (N_9920,N_9219,N_9290);
nor U9921 (N_9921,N_9065,N_9133);
and U9922 (N_9922,N_9079,N_9107);
nand U9923 (N_9923,N_8810,N_9305);
xor U9924 (N_9924,N_9073,N_9024);
or U9925 (N_9925,N_8981,N_9362);
xnor U9926 (N_9926,N_8946,N_9077);
xnor U9927 (N_9927,N_8926,N_8949);
nor U9928 (N_9928,N_8780,N_8758);
nand U9929 (N_9929,N_9300,N_9000);
nand U9930 (N_9930,N_9181,N_9158);
or U9931 (N_9931,N_9152,N_8961);
xor U9932 (N_9932,N_8887,N_8900);
and U9933 (N_9933,N_9127,N_9075);
nand U9934 (N_9934,N_8794,N_9125);
nor U9935 (N_9935,N_8996,N_9182);
and U9936 (N_9936,N_8961,N_8834);
nor U9937 (N_9937,N_8790,N_8774);
nor U9938 (N_9938,N_8791,N_8949);
nand U9939 (N_9939,N_8799,N_8846);
xor U9940 (N_9940,N_9145,N_8812);
or U9941 (N_9941,N_8885,N_9238);
xnor U9942 (N_9942,N_9108,N_9155);
nor U9943 (N_9943,N_8911,N_9035);
or U9944 (N_9944,N_9201,N_9289);
and U9945 (N_9945,N_8782,N_8981);
xor U9946 (N_9946,N_9270,N_8950);
nor U9947 (N_9947,N_9168,N_8950);
xnor U9948 (N_9948,N_9031,N_9098);
nand U9949 (N_9949,N_8902,N_9351);
nor U9950 (N_9950,N_9201,N_8815);
nor U9951 (N_9951,N_8989,N_8786);
nor U9952 (N_9952,N_8972,N_9251);
or U9953 (N_9953,N_9048,N_9158);
nor U9954 (N_9954,N_8875,N_9236);
and U9955 (N_9955,N_9290,N_8885);
or U9956 (N_9956,N_9121,N_8991);
xor U9957 (N_9957,N_8769,N_9070);
xnor U9958 (N_9958,N_9104,N_8800);
xnor U9959 (N_9959,N_8961,N_8778);
nand U9960 (N_9960,N_9316,N_9309);
nor U9961 (N_9961,N_9326,N_8843);
nor U9962 (N_9962,N_8810,N_9012);
nand U9963 (N_9963,N_9324,N_9238);
or U9964 (N_9964,N_9361,N_9238);
nand U9965 (N_9965,N_9106,N_8954);
xnor U9966 (N_9966,N_9217,N_9057);
xnor U9967 (N_9967,N_9147,N_8846);
xor U9968 (N_9968,N_9114,N_9139);
and U9969 (N_9969,N_8849,N_9066);
nor U9970 (N_9970,N_8765,N_9139);
and U9971 (N_9971,N_9059,N_8757);
xor U9972 (N_9972,N_9151,N_8899);
nor U9973 (N_9973,N_8973,N_8862);
or U9974 (N_9974,N_9362,N_8903);
xor U9975 (N_9975,N_9013,N_8908);
nand U9976 (N_9976,N_9139,N_8849);
and U9977 (N_9977,N_8800,N_9164);
nand U9978 (N_9978,N_8782,N_8940);
and U9979 (N_9979,N_9209,N_9144);
xor U9980 (N_9980,N_9232,N_9156);
or U9981 (N_9981,N_8861,N_8802);
and U9982 (N_9982,N_9214,N_8851);
nor U9983 (N_9983,N_9138,N_8931);
nor U9984 (N_9984,N_8945,N_8933);
nor U9985 (N_9985,N_8823,N_8856);
and U9986 (N_9986,N_9005,N_8769);
or U9987 (N_9987,N_9161,N_8958);
xnor U9988 (N_9988,N_8802,N_9276);
nand U9989 (N_9989,N_8938,N_9217);
nand U9990 (N_9990,N_8828,N_9363);
nand U9991 (N_9991,N_9213,N_8781);
nor U9992 (N_9992,N_9255,N_8819);
and U9993 (N_9993,N_9302,N_9197);
and U9994 (N_9994,N_8962,N_8841);
and U9995 (N_9995,N_8816,N_8775);
nand U9996 (N_9996,N_8847,N_9195);
nor U9997 (N_9997,N_8813,N_9324);
or U9998 (N_9998,N_9296,N_9282);
xor U9999 (N_9999,N_9353,N_8954);
and U10000 (N_10000,N_9856,N_9471);
nand U10001 (N_10001,N_9943,N_9530);
nand U10002 (N_10002,N_9861,N_9986);
or U10003 (N_10003,N_9784,N_9953);
nand U10004 (N_10004,N_9996,N_9490);
xnor U10005 (N_10005,N_9540,N_9580);
nand U10006 (N_10006,N_9764,N_9839);
or U10007 (N_10007,N_9698,N_9512);
nand U10008 (N_10008,N_9837,N_9380);
nor U10009 (N_10009,N_9898,N_9911);
and U10010 (N_10010,N_9711,N_9757);
and U10011 (N_10011,N_9554,N_9915);
xnor U10012 (N_10012,N_9716,N_9809);
xor U10013 (N_10013,N_9460,N_9476);
nor U10014 (N_10014,N_9412,N_9690);
nand U10015 (N_10015,N_9655,N_9594);
or U10016 (N_10016,N_9833,N_9922);
xnor U10017 (N_10017,N_9546,N_9989);
nor U10018 (N_10018,N_9563,N_9744);
or U10019 (N_10019,N_9997,N_9397);
xor U10020 (N_10020,N_9959,N_9806);
nor U10021 (N_10021,N_9488,N_9613);
nand U10022 (N_10022,N_9500,N_9936);
or U10023 (N_10023,N_9693,N_9736);
nand U10024 (N_10024,N_9383,N_9468);
and U10025 (N_10025,N_9639,N_9559);
nand U10026 (N_10026,N_9504,N_9623);
and U10027 (N_10027,N_9527,N_9436);
or U10028 (N_10028,N_9450,N_9466);
or U10029 (N_10029,N_9887,N_9393);
and U10030 (N_10030,N_9684,N_9664);
xor U10031 (N_10031,N_9858,N_9726);
nand U10032 (N_10032,N_9657,N_9782);
xnor U10033 (N_10033,N_9987,N_9905);
or U10034 (N_10034,N_9955,N_9823);
xor U10035 (N_10035,N_9973,N_9673);
nor U10036 (N_10036,N_9950,N_9574);
xnor U10037 (N_10037,N_9890,N_9560);
nand U10038 (N_10038,N_9850,N_9398);
nor U10039 (N_10039,N_9451,N_9618);
or U10040 (N_10040,N_9995,N_9854);
nand U10041 (N_10041,N_9982,N_9708);
nand U10042 (N_10042,N_9789,N_9386);
nor U10043 (N_10043,N_9998,N_9941);
and U10044 (N_10044,N_9914,N_9579);
nor U10045 (N_10045,N_9608,N_9881);
nand U10046 (N_10046,N_9805,N_9528);
xor U10047 (N_10047,N_9666,N_9886);
and U10048 (N_10048,N_9503,N_9962);
nand U10049 (N_10049,N_9773,N_9739);
nor U10050 (N_10050,N_9552,N_9536);
nor U10051 (N_10051,N_9831,N_9897);
or U10052 (N_10052,N_9663,N_9958);
or U10053 (N_10053,N_9642,N_9849);
xor U10054 (N_10054,N_9689,N_9867);
or U10055 (N_10055,N_9644,N_9584);
nand U10056 (N_10056,N_9878,N_9427);
nand U10057 (N_10057,N_9767,N_9847);
and U10058 (N_10058,N_9961,N_9990);
or U10059 (N_10059,N_9960,N_9970);
nand U10060 (N_10060,N_9585,N_9769);
nand U10061 (N_10061,N_9686,N_9855);
nand U10062 (N_10062,N_9889,N_9907);
or U10063 (N_10063,N_9649,N_9801);
nor U10064 (N_10064,N_9654,N_9691);
nor U10065 (N_10065,N_9884,N_9851);
xor U10066 (N_10066,N_9414,N_9892);
and U10067 (N_10067,N_9766,N_9821);
and U10068 (N_10068,N_9582,N_9683);
xor U10069 (N_10069,N_9755,N_9695);
nand U10070 (N_10070,N_9944,N_9724);
or U10071 (N_10071,N_9906,N_9830);
nor U10072 (N_10072,N_9675,N_9583);
nand U10073 (N_10073,N_9413,N_9692);
nand U10074 (N_10074,N_9923,N_9635);
and U10075 (N_10075,N_9550,N_9390);
nor U10076 (N_10076,N_9719,N_9824);
xnor U10077 (N_10077,N_9481,N_9566);
nand U10078 (N_10078,N_9632,N_9904);
and U10079 (N_10079,N_9803,N_9981);
nor U10080 (N_10080,N_9571,N_9377);
nor U10081 (N_10081,N_9510,N_9511);
xor U10082 (N_10082,N_9796,N_9533);
and U10083 (N_10083,N_9539,N_9478);
xnor U10084 (N_10084,N_9707,N_9857);
nand U10085 (N_10085,N_9487,N_9624);
xor U10086 (N_10086,N_9388,N_9760);
or U10087 (N_10087,N_9859,N_9843);
xnor U10088 (N_10088,N_9910,N_9799);
xnor U10089 (N_10089,N_9551,N_9865);
or U10090 (N_10090,N_9697,N_9746);
and U10091 (N_10091,N_9917,N_9593);
and U10092 (N_10092,N_9709,N_9677);
xor U10093 (N_10093,N_9676,N_9862);
or U10094 (N_10094,N_9896,N_9971);
nand U10095 (N_10095,N_9699,N_9991);
nor U10096 (N_10096,N_9431,N_9807);
or U10097 (N_10097,N_9758,N_9491);
nand U10098 (N_10098,N_9727,N_9592);
xnor U10099 (N_10099,N_9591,N_9710);
nand U10100 (N_10100,N_9794,N_9756);
nor U10101 (N_10101,N_9834,N_9474);
nor U10102 (N_10102,N_9422,N_9885);
and U10103 (N_10103,N_9828,N_9581);
and U10104 (N_10104,N_9440,N_9389);
nand U10105 (N_10105,N_9542,N_9826);
nor U10106 (N_10106,N_9932,N_9455);
nor U10107 (N_10107,N_9477,N_9660);
or U10108 (N_10108,N_9548,N_9815);
and U10109 (N_10109,N_9507,N_9406);
and U10110 (N_10110,N_9827,N_9588);
xor U10111 (N_10111,N_9547,N_9395);
nand U10112 (N_10112,N_9670,N_9974);
or U10113 (N_10113,N_9420,N_9493);
xnor U10114 (N_10114,N_9903,N_9720);
nand U10115 (N_10115,N_9751,N_9921);
or U10116 (N_10116,N_9852,N_9496);
or U10117 (N_10117,N_9405,N_9901);
or U10118 (N_10118,N_9453,N_9771);
nand U10119 (N_10119,N_9517,N_9653);
or U10120 (N_10120,N_9718,N_9871);
or U10121 (N_10121,N_9965,N_9438);
nand U10122 (N_10122,N_9715,N_9514);
xor U10123 (N_10123,N_9461,N_9387);
nor U10124 (N_10124,N_9629,N_9752);
and U10125 (N_10125,N_9616,N_9534);
nor U10126 (N_10126,N_9628,N_9780);
nor U10127 (N_10127,N_9685,N_9983);
xor U10128 (N_10128,N_9439,N_9734);
and U10129 (N_10129,N_9602,N_9385);
nor U10130 (N_10130,N_9772,N_9521);
and U10131 (N_10131,N_9661,N_9706);
xnor U10132 (N_10132,N_9988,N_9938);
nor U10133 (N_10133,N_9688,N_9515);
xnor U10134 (N_10134,N_9770,N_9577);
nor U10135 (N_10135,N_9721,N_9810);
nor U10136 (N_10136,N_9424,N_9741);
and U10137 (N_10137,N_9786,N_9410);
nor U10138 (N_10138,N_9379,N_9599);
and U10139 (N_10139,N_9381,N_9929);
nand U10140 (N_10140,N_9745,N_9893);
and U10141 (N_10141,N_9646,N_9595);
nand U10142 (N_10142,N_9482,N_9817);
xnor U10143 (N_10143,N_9696,N_9637);
and U10144 (N_10144,N_9924,N_9444);
and U10145 (N_10145,N_9656,N_9658);
and U10146 (N_10146,N_9868,N_9875);
or U10147 (N_10147,N_9747,N_9912);
xor U10148 (N_10148,N_9877,N_9553);
nor U10149 (N_10149,N_9399,N_9494);
or U10150 (N_10150,N_9880,N_9407);
or U10151 (N_10151,N_9732,N_9781);
or U10152 (N_10152,N_9733,N_9568);
nand U10153 (N_10153,N_9625,N_9761);
or U10154 (N_10154,N_9607,N_9798);
or U10155 (N_10155,N_9442,N_9863);
nor U10156 (N_10156,N_9425,N_9452);
and U10157 (N_10157,N_9419,N_9882);
nor U10158 (N_10158,N_9384,N_9870);
or U10159 (N_10159,N_9802,N_9793);
nand U10160 (N_10160,N_9909,N_9565);
nand U10161 (N_10161,N_9788,N_9735);
and U10162 (N_10162,N_9813,N_9722);
xor U10163 (N_10163,N_9952,N_9900);
and U10164 (N_10164,N_9681,N_9648);
nor U10165 (N_10165,N_9475,N_9753);
or U10166 (N_10166,N_9590,N_9489);
xor U10167 (N_10167,N_9940,N_9454);
nor U10168 (N_10168,N_9790,N_9668);
xor U10169 (N_10169,N_9860,N_9768);
or U10170 (N_10170,N_9462,N_9956);
or U10171 (N_10171,N_9509,N_9783);
nand U10172 (N_10172,N_9626,N_9712);
nand U10173 (N_10173,N_9762,N_9469);
xor U10174 (N_10174,N_9416,N_9879);
xor U10175 (N_10175,N_9844,N_9842);
or U10176 (N_10176,N_9894,N_9501);
and U10177 (N_10177,N_9538,N_9423);
nand U10178 (N_10178,N_9957,N_9446);
nor U10179 (N_10179,N_9576,N_9874);
nor U10180 (N_10180,N_9611,N_9967);
xor U10181 (N_10181,N_9409,N_9933);
or U10182 (N_10182,N_9964,N_9949);
xnor U10183 (N_10183,N_9428,N_9603);
xnor U10184 (N_10184,N_9508,N_9759);
nand U10185 (N_10185,N_9787,N_9717);
and U10186 (N_10186,N_9408,N_9627);
nand U10187 (N_10187,N_9415,N_9774);
nor U10188 (N_10188,N_9633,N_9704);
nor U10189 (N_10189,N_9836,N_9640);
nor U10190 (N_10190,N_9433,N_9819);
nand U10191 (N_10191,N_9641,N_9946);
or U10192 (N_10192,N_9978,N_9435);
nand U10193 (N_10193,N_9919,N_9418);
xor U10194 (N_10194,N_9643,N_9445);
nor U10195 (N_10195,N_9524,N_9532);
xor U10196 (N_10196,N_9457,N_9876);
or U10197 (N_10197,N_9825,N_9812);
nand U10198 (N_10198,N_9908,N_9984);
or U10199 (N_10199,N_9700,N_9776);
or U10200 (N_10200,N_9951,N_9662);
and U10201 (N_10201,N_9537,N_9808);
nand U10202 (N_10202,N_9421,N_9572);
or U10203 (N_10203,N_9569,N_9479);
nor U10204 (N_10204,N_9678,N_9969);
and U10205 (N_10205,N_9864,N_9578);
nor U10206 (N_10206,N_9846,N_9609);
and U10207 (N_10207,N_9601,N_9441);
nor U10208 (N_10208,N_9523,N_9895);
xnor U10209 (N_10209,N_9520,N_9672);
or U10210 (N_10210,N_9645,N_9920);
nor U10211 (N_10211,N_9737,N_9561);
and U10212 (N_10212,N_9596,N_9604);
and U10213 (N_10213,N_9480,N_9619);
or U10214 (N_10214,N_9713,N_9531);
xor U10215 (N_10215,N_9615,N_9391);
or U10216 (N_10216,N_9522,N_9667);
xnor U10217 (N_10217,N_9483,N_9979);
xnor U10218 (N_10218,N_9529,N_9394);
or U10219 (N_10219,N_9703,N_9518);
or U10220 (N_10220,N_9541,N_9976);
nand U10221 (N_10221,N_9838,N_9417);
nor U10222 (N_10222,N_9543,N_9647);
xor U10223 (N_10223,N_9738,N_9456);
nand U10224 (N_10224,N_9763,N_9492);
xnor U10225 (N_10225,N_9634,N_9411);
nand U10226 (N_10226,N_9945,N_9994);
nor U10227 (N_10227,N_9785,N_9845);
or U10228 (N_10228,N_9485,N_9972);
xnor U10229 (N_10229,N_9525,N_9883);
nand U10230 (N_10230,N_9954,N_9401);
xor U10231 (N_10231,N_9866,N_9631);
nand U10232 (N_10232,N_9728,N_9557);
nand U10233 (N_10233,N_9535,N_9749);
xnor U10234 (N_10234,N_9621,N_9927);
nand U10235 (N_10235,N_9587,N_9447);
xor U10236 (N_10236,N_9564,N_9832);
xor U10237 (N_10237,N_9396,N_9814);
xor U10238 (N_10238,N_9519,N_9916);
or U10239 (N_10239,N_9651,N_9470);
or U10240 (N_10240,N_9777,N_9443);
and U10241 (N_10241,N_9544,N_9742);
and U10242 (N_10242,N_9975,N_9495);
xor U10243 (N_10243,N_9636,N_9558);
nor U10244 (N_10244,N_9937,N_9376);
or U10245 (N_10245,N_9570,N_9448);
xnor U10246 (N_10246,N_9650,N_9797);
or U10247 (N_10247,N_9723,N_9586);
nand U10248 (N_10248,N_9665,N_9891);
xor U10249 (N_10249,N_9400,N_9502);
nor U10250 (N_10250,N_9968,N_9754);
nand U10251 (N_10251,N_9873,N_9404);
xor U10252 (N_10252,N_9464,N_9942);
xor U10253 (N_10253,N_9597,N_9562);
nor U10254 (N_10254,N_9966,N_9382);
or U10255 (N_10255,N_9606,N_9985);
nor U10256 (N_10256,N_9841,N_9614);
and U10257 (N_10257,N_9934,N_9498);
nand U10258 (N_10258,N_9775,N_9437);
or U10259 (N_10259,N_9638,N_9549);
or U10260 (N_10260,N_9467,N_9714);
and U10261 (N_10261,N_9926,N_9935);
xnor U10262 (N_10262,N_9820,N_9497);
or U10263 (N_10263,N_9499,N_9899);
nor U10264 (N_10264,N_9816,N_9791);
nand U10265 (N_10265,N_9622,N_9913);
nand U10266 (N_10266,N_9853,N_9818);
nand U10267 (N_10267,N_9925,N_9378);
nor U10268 (N_10268,N_9800,N_9573);
or U10269 (N_10269,N_9486,N_9598);
or U10270 (N_10270,N_9947,N_9659);
and U10271 (N_10271,N_9432,N_9556);
xnor U10272 (N_10272,N_9575,N_9620);
or U10273 (N_10273,N_9617,N_9459);
xnor U10274 (N_10274,N_9392,N_9829);
nor U10275 (N_10275,N_9999,N_9931);
nand U10276 (N_10276,N_9682,N_9484);
nand U10277 (N_10277,N_9473,N_9928);
and U10278 (N_10278,N_9822,N_9730);
nor U10279 (N_10279,N_9679,N_9630);
xor U10280 (N_10280,N_9612,N_9993);
nand U10281 (N_10281,N_9701,N_9729);
and U10282 (N_10282,N_9605,N_9930);
nor U10283 (N_10283,N_9600,N_9779);
and U10284 (N_10284,N_9434,N_9429);
and U10285 (N_10285,N_9804,N_9795);
and U10286 (N_10286,N_9505,N_9835);
xnor U10287 (N_10287,N_9743,N_9977);
and U10288 (N_10288,N_9902,N_9702);
xor U10289 (N_10289,N_9992,N_9513);
nor U10290 (N_10290,N_9740,N_9516);
nand U10291 (N_10291,N_9840,N_9725);
nand U10292 (N_10292,N_9567,N_9375);
or U10293 (N_10293,N_9811,N_9506);
and U10294 (N_10294,N_9669,N_9674);
nor U10295 (N_10295,N_9526,N_9750);
nor U10296 (N_10296,N_9430,N_9671);
and U10297 (N_10297,N_9872,N_9545);
or U10298 (N_10298,N_9888,N_9948);
nor U10299 (N_10299,N_9402,N_9472);
nand U10300 (N_10300,N_9748,N_9731);
nand U10301 (N_10301,N_9589,N_9705);
nand U10302 (N_10302,N_9792,N_9458);
nor U10303 (N_10303,N_9963,N_9869);
nor U10304 (N_10304,N_9610,N_9652);
and U10305 (N_10305,N_9687,N_9680);
or U10306 (N_10306,N_9555,N_9918);
xor U10307 (N_10307,N_9426,N_9848);
or U10308 (N_10308,N_9449,N_9463);
nand U10309 (N_10309,N_9694,N_9765);
nor U10310 (N_10310,N_9980,N_9465);
xnor U10311 (N_10311,N_9403,N_9939);
xnor U10312 (N_10312,N_9778,N_9699);
nand U10313 (N_10313,N_9835,N_9970);
and U10314 (N_10314,N_9952,N_9619);
or U10315 (N_10315,N_9403,N_9478);
xor U10316 (N_10316,N_9521,N_9984);
xor U10317 (N_10317,N_9468,N_9530);
nand U10318 (N_10318,N_9601,N_9475);
nand U10319 (N_10319,N_9958,N_9930);
xnor U10320 (N_10320,N_9582,N_9934);
and U10321 (N_10321,N_9806,N_9954);
xor U10322 (N_10322,N_9656,N_9376);
nor U10323 (N_10323,N_9526,N_9687);
xor U10324 (N_10324,N_9830,N_9859);
xor U10325 (N_10325,N_9547,N_9786);
nand U10326 (N_10326,N_9848,N_9634);
nor U10327 (N_10327,N_9985,N_9500);
nor U10328 (N_10328,N_9894,N_9576);
or U10329 (N_10329,N_9669,N_9791);
and U10330 (N_10330,N_9881,N_9499);
nand U10331 (N_10331,N_9543,N_9852);
or U10332 (N_10332,N_9717,N_9506);
nand U10333 (N_10333,N_9647,N_9849);
and U10334 (N_10334,N_9899,N_9498);
xor U10335 (N_10335,N_9600,N_9853);
nor U10336 (N_10336,N_9464,N_9456);
xnor U10337 (N_10337,N_9509,N_9781);
nand U10338 (N_10338,N_9683,N_9871);
and U10339 (N_10339,N_9529,N_9836);
or U10340 (N_10340,N_9747,N_9591);
xor U10341 (N_10341,N_9416,N_9393);
and U10342 (N_10342,N_9908,N_9620);
nand U10343 (N_10343,N_9652,N_9804);
xor U10344 (N_10344,N_9648,N_9412);
xor U10345 (N_10345,N_9882,N_9380);
nand U10346 (N_10346,N_9497,N_9463);
or U10347 (N_10347,N_9524,N_9538);
xnor U10348 (N_10348,N_9858,N_9524);
and U10349 (N_10349,N_9739,N_9806);
nor U10350 (N_10350,N_9787,N_9692);
nand U10351 (N_10351,N_9481,N_9816);
or U10352 (N_10352,N_9859,N_9748);
xnor U10353 (N_10353,N_9413,N_9465);
xnor U10354 (N_10354,N_9514,N_9375);
nor U10355 (N_10355,N_9548,N_9841);
or U10356 (N_10356,N_9992,N_9574);
or U10357 (N_10357,N_9632,N_9564);
nand U10358 (N_10358,N_9659,N_9503);
nor U10359 (N_10359,N_9643,N_9986);
or U10360 (N_10360,N_9509,N_9852);
or U10361 (N_10361,N_9579,N_9483);
xor U10362 (N_10362,N_9830,N_9683);
nor U10363 (N_10363,N_9779,N_9698);
nand U10364 (N_10364,N_9619,N_9447);
nor U10365 (N_10365,N_9509,N_9740);
and U10366 (N_10366,N_9811,N_9680);
and U10367 (N_10367,N_9738,N_9694);
nand U10368 (N_10368,N_9785,N_9810);
nand U10369 (N_10369,N_9931,N_9868);
xor U10370 (N_10370,N_9750,N_9749);
and U10371 (N_10371,N_9673,N_9459);
xnor U10372 (N_10372,N_9845,N_9524);
xor U10373 (N_10373,N_9432,N_9567);
or U10374 (N_10374,N_9431,N_9384);
xor U10375 (N_10375,N_9452,N_9706);
or U10376 (N_10376,N_9810,N_9880);
or U10377 (N_10377,N_9592,N_9416);
or U10378 (N_10378,N_9711,N_9972);
nand U10379 (N_10379,N_9468,N_9829);
nor U10380 (N_10380,N_9876,N_9883);
and U10381 (N_10381,N_9781,N_9965);
nor U10382 (N_10382,N_9418,N_9927);
nor U10383 (N_10383,N_9592,N_9391);
nand U10384 (N_10384,N_9554,N_9519);
or U10385 (N_10385,N_9480,N_9812);
or U10386 (N_10386,N_9706,N_9736);
nand U10387 (N_10387,N_9742,N_9994);
nand U10388 (N_10388,N_9572,N_9547);
nand U10389 (N_10389,N_9839,N_9787);
nor U10390 (N_10390,N_9534,N_9693);
or U10391 (N_10391,N_9829,N_9866);
or U10392 (N_10392,N_9821,N_9758);
xnor U10393 (N_10393,N_9735,N_9499);
and U10394 (N_10394,N_9706,N_9893);
nor U10395 (N_10395,N_9863,N_9801);
xnor U10396 (N_10396,N_9702,N_9641);
xnor U10397 (N_10397,N_9497,N_9383);
nand U10398 (N_10398,N_9805,N_9858);
or U10399 (N_10399,N_9554,N_9599);
nor U10400 (N_10400,N_9856,N_9704);
or U10401 (N_10401,N_9698,N_9997);
nand U10402 (N_10402,N_9801,N_9866);
nor U10403 (N_10403,N_9622,N_9638);
and U10404 (N_10404,N_9684,N_9694);
or U10405 (N_10405,N_9700,N_9612);
and U10406 (N_10406,N_9395,N_9801);
or U10407 (N_10407,N_9735,N_9895);
and U10408 (N_10408,N_9455,N_9829);
nand U10409 (N_10409,N_9662,N_9920);
nor U10410 (N_10410,N_9800,N_9881);
nand U10411 (N_10411,N_9776,N_9427);
and U10412 (N_10412,N_9659,N_9559);
or U10413 (N_10413,N_9808,N_9686);
nand U10414 (N_10414,N_9996,N_9462);
or U10415 (N_10415,N_9624,N_9535);
xor U10416 (N_10416,N_9630,N_9781);
or U10417 (N_10417,N_9608,N_9906);
and U10418 (N_10418,N_9661,N_9834);
nor U10419 (N_10419,N_9918,N_9940);
nor U10420 (N_10420,N_9991,N_9670);
xnor U10421 (N_10421,N_9902,N_9463);
nand U10422 (N_10422,N_9747,N_9768);
nor U10423 (N_10423,N_9711,N_9932);
and U10424 (N_10424,N_9432,N_9499);
nand U10425 (N_10425,N_9876,N_9710);
or U10426 (N_10426,N_9450,N_9724);
or U10427 (N_10427,N_9685,N_9839);
and U10428 (N_10428,N_9973,N_9669);
nand U10429 (N_10429,N_9781,N_9644);
xnor U10430 (N_10430,N_9493,N_9986);
or U10431 (N_10431,N_9607,N_9713);
or U10432 (N_10432,N_9928,N_9803);
nor U10433 (N_10433,N_9685,N_9379);
nand U10434 (N_10434,N_9580,N_9601);
and U10435 (N_10435,N_9454,N_9809);
xnor U10436 (N_10436,N_9521,N_9858);
xor U10437 (N_10437,N_9901,N_9793);
nor U10438 (N_10438,N_9674,N_9762);
nand U10439 (N_10439,N_9768,N_9848);
or U10440 (N_10440,N_9506,N_9723);
xnor U10441 (N_10441,N_9846,N_9608);
xnor U10442 (N_10442,N_9647,N_9678);
nor U10443 (N_10443,N_9587,N_9425);
or U10444 (N_10444,N_9575,N_9857);
nor U10445 (N_10445,N_9518,N_9595);
or U10446 (N_10446,N_9441,N_9814);
nand U10447 (N_10447,N_9889,N_9753);
nand U10448 (N_10448,N_9566,N_9485);
nand U10449 (N_10449,N_9688,N_9966);
or U10450 (N_10450,N_9831,N_9786);
and U10451 (N_10451,N_9637,N_9685);
and U10452 (N_10452,N_9607,N_9410);
nand U10453 (N_10453,N_9626,N_9635);
and U10454 (N_10454,N_9753,N_9767);
nand U10455 (N_10455,N_9431,N_9563);
or U10456 (N_10456,N_9894,N_9593);
nor U10457 (N_10457,N_9626,N_9893);
and U10458 (N_10458,N_9637,N_9930);
nor U10459 (N_10459,N_9765,N_9652);
nand U10460 (N_10460,N_9599,N_9440);
nor U10461 (N_10461,N_9767,N_9866);
nand U10462 (N_10462,N_9998,N_9639);
xor U10463 (N_10463,N_9913,N_9453);
and U10464 (N_10464,N_9783,N_9702);
nor U10465 (N_10465,N_9478,N_9734);
and U10466 (N_10466,N_9914,N_9834);
xnor U10467 (N_10467,N_9889,N_9748);
and U10468 (N_10468,N_9522,N_9849);
nor U10469 (N_10469,N_9723,N_9718);
nor U10470 (N_10470,N_9490,N_9412);
xor U10471 (N_10471,N_9501,N_9755);
or U10472 (N_10472,N_9892,N_9544);
nand U10473 (N_10473,N_9744,N_9980);
nor U10474 (N_10474,N_9711,N_9808);
nand U10475 (N_10475,N_9511,N_9445);
or U10476 (N_10476,N_9801,N_9885);
or U10477 (N_10477,N_9949,N_9494);
xor U10478 (N_10478,N_9942,N_9645);
or U10479 (N_10479,N_9697,N_9382);
nor U10480 (N_10480,N_9387,N_9599);
nand U10481 (N_10481,N_9412,N_9729);
nand U10482 (N_10482,N_9449,N_9785);
nor U10483 (N_10483,N_9525,N_9480);
nand U10484 (N_10484,N_9459,N_9795);
and U10485 (N_10485,N_9492,N_9873);
nand U10486 (N_10486,N_9887,N_9635);
and U10487 (N_10487,N_9591,N_9696);
and U10488 (N_10488,N_9964,N_9529);
or U10489 (N_10489,N_9712,N_9569);
or U10490 (N_10490,N_9393,N_9989);
and U10491 (N_10491,N_9769,N_9715);
nor U10492 (N_10492,N_9856,N_9592);
and U10493 (N_10493,N_9627,N_9772);
and U10494 (N_10494,N_9828,N_9878);
and U10495 (N_10495,N_9718,N_9544);
nand U10496 (N_10496,N_9708,N_9480);
xnor U10497 (N_10497,N_9832,N_9854);
and U10498 (N_10498,N_9577,N_9993);
and U10499 (N_10499,N_9745,N_9943);
nand U10500 (N_10500,N_9831,N_9701);
nand U10501 (N_10501,N_9415,N_9503);
and U10502 (N_10502,N_9901,N_9460);
nand U10503 (N_10503,N_9983,N_9544);
and U10504 (N_10504,N_9901,N_9904);
and U10505 (N_10505,N_9706,N_9725);
and U10506 (N_10506,N_9468,N_9980);
or U10507 (N_10507,N_9735,N_9672);
xnor U10508 (N_10508,N_9906,N_9963);
or U10509 (N_10509,N_9623,N_9990);
and U10510 (N_10510,N_9641,N_9602);
nand U10511 (N_10511,N_9912,N_9545);
nor U10512 (N_10512,N_9754,N_9644);
nand U10513 (N_10513,N_9779,N_9761);
nor U10514 (N_10514,N_9881,N_9651);
nor U10515 (N_10515,N_9507,N_9909);
or U10516 (N_10516,N_9836,N_9923);
xor U10517 (N_10517,N_9716,N_9946);
xnor U10518 (N_10518,N_9984,N_9870);
and U10519 (N_10519,N_9553,N_9597);
xnor U10520 (N_10520,N_9586,N_9674);
xnor U10521 (N_10521,N_9605,N_9541);
xor U10522 (N_10522,N_9473,N_9894);
nor U10523 (N_10523,N_9660,N_9637);
nand U10524 (N_10524,N_9850,N_9524);
or U10525 (N_10525,N_9498,N_9800);
or U10526 (N_10526,N_9863,N_9477);
or U10527 (N_10527,N_9699,N_9595);
and U10528 (N_10528,N_9780,N_9515);
or U10529 (N_10529,N_9649,N_9771);
nand U10530 (N_10530,N_9416,N_9662);
and U10531 (N_10531,N_9623,N_9472);
and U10532 (N_10532,N_9998,N_9709);
and U10533 (N_10533,N_9837,N_9688);
or U10534 (N_10534,N_9956,N_9596);
xor U10535 (N_10535,N_9481,N_9915);
nand U10536 (N_10536,N_9483,N_9426);
nand U10537 (N_10537,N_9965,N_9655);
xnor U10538 (N_10538,N_9624,N_9791);
xnor U10539 (N_10539,N_9744,N_9424);
or U10540 (N_10540,N_9548,N_9956);
and U10541 (N_10541,N_9887,N_9512);
or U10542 (N_10542,N_9394,N_9402);
xor U10543 (N_10543,N_9777,N_9651);
nand U10544 (N_10544,N_9826,N_9743);
nand U10545 (N_10545,N_9489,N_9440);
nand U10546 (N_10546,N_9992,N_9900);
nand U10547 (N_10547,N_9832,N_9437);
nor U10548 (N_10548,N_9651,N_9686);
xnor U10549 (N_10549,N_9674,N_9885);
xor U10550 (N_10550,N_9978,N_9875);
or U10551 (N_10551,N_9849,N_9961);
and U10552 (N_10552,N_9544,N_9895);
nor U10553 (N_10553,N_9936,N_9385);
xor U10554 (N_10554,N_9705,N_9500);
and U10555 (N_10555,N_9497,N_9638);
and U10556 (N_10556,N_9686,N_9930);
nor U10557 (N_10557,N_9782,N_9463);
nand U10558 (N_10558,N_9518,N_9831);
xor U10559 (N_10559,N_9617,N_9712);
or U10560 (N_10560,N_9824,N_9769);
or U10561 (N_10561,N_9715,N_9761);
xnor U10562 (N_10562,N_9815,N_9753);
nor U10563 (N_10563,N_9387,N_9428);
and U10564 (N_10564,N_9866,N_9915);
nand U10565 (N_10565,N_9568,N_9895);
and U10566 (N_10566,N_9996,N_9468);
nand U10567 (N_10567,N_9814,N_9738);
or U10568 (N_10568,N_9866,N_9842);
and U10569 (N_10569,N_9820,N_9875);
and U10570 (N_10570,N_9721,N_9704);
nand U10571 (N_10571,N_9904,N_9558);
nor U10572 (N_10572,N_9482,N_9440);
nand U10573 (N_10573,N_9757,N_9685);
nor U10574 (N_10574,N_9520,N_9455);
xor U10575 (N_10575,N_9428,N_9558);
xor U10576 (N_10576,N_9809,N_9519);
or U10577 (N_10577,N_9738,N_9674);
nand U10578 (N_10578,N_9721,N_9943);
and U10579 (N_10579,N_9595,N_9536);
or U10580 (N_10580,N_9694,N_9896);
and U10581 (N_10581,N_9788,N_9628);
or U10582 (N_10582,N_9744,N_9919);
xor U10583 (N_10583,N_9860,N_9624);
and U10584 (N_10584,N_9485,N_9948);
xnor U10585 (N_10585,N_9773,N_9905);
nor U10586 (N_10586,N_9736,N_9532);
nor U10587 (N_10587,N_9591,N_9493);
xnor U10588 (N_10588,N_9939,N_9585);
nand U10589 (N_10589,N_9804,N_9665);
xor U10590 (N_10590,N_9930,N_9629);
or U10591 (N_10591,N_9419,N_9630);
or U10592 (N_10592,N_9868,N_9558);
xnor U10593 (N_10593,N_9668,N_9706);
nand U10594 (N_10594,N_9808,N_9563);
or U10595 (N_10595,N_9942,N_9421);
and U10596 (N_10596,N_9891,N_9959);
or U10597 (N_10597,N_9729,N_9920);
and U10598 (N_10598,N_9741,N_9597);
nand U10599 (N_10599,N_9974,N_9994);
xnor U10600 (N_10600,N_9537,N_9963);
or U10601 (N_10601,N_9950,N_9912);
or U10602 (N_10602,N_9811,N_9883);
xor U10603 (N_10603,N_9442,N_9640);
or U10604 (N_10604,N_9913,N_9788);
nor U10605 (N_10605,N_9672,N_9578);
and U10606 (N_10606,N_9931,N_9871);
and U10607 (N_10607,N_9995,N_9813);
or U10608 (N_10608,N_9845,N_9620);
nand U10609 (N_10609,N_9969,N_9751);
xor U10610 (N_10610,N_9698,N_9843);
and U10611 (N_10611,N_9844,N_9677);
nor U10612 (N_10612,N_9614,N_9730);
nor U10613 (N_10613,N_9905,N_9849);
and U10614 (N_10614,N_9691,N_9380);
nor U10615 (N_10615,N_9666,N_9474);
nor U10616 (N_10616,N_9955,N_9934);
and U10617 (N_10617,N_9375,N_9467);
nand U10618 (N_10618,N_9641,N_9591);
xnor U10619 (N_10619,N_9375,N_9570);
xnor U10620 (N_10620,N_9571,N_9517);
nand U10621 (N_10621,N_9435,N_9544);
nor U10622 (N_10622,N_9941,N_9503);
xnor U10623 (N_10623,N_9836,N_9567);
or U10624 (N_10624,N_9981,N_9768);
or U10625 (N_10625,N_10552,N_10592);
and U10626 (N_10626,N_10174,N_10134);
xor U10627 (N_10627,N_10195,N_10453);
nor U10628 (N_10628,N_10374,N_10284);
nor U10629 (N_10629,N_10233,N_10491);
nor U10630 (N_10630,N_10367,N_10496);
or U10631 (N_10631,N_10467,N_10069);
xor U10632 (N_10632,N_10021,N_10152);
nand U10633 (N_10633,N_10263,N_10312);
xor U10634 (N_10634,N_10330,N_10487);
or U10635 (N_10635,N_10131,N_10297);
or U10636 (N_10636,N_10031,N_10256);
nand U10637 (N_10637,N_10465,N_10371);
xor U10638 (N_10638,N_10381,N_10214);
xnor U10639 (N_10639,N_10156,N_10614);
xor U10640 (N_10640,N_10389,N_10165);
or U10641 (N_10641,N_10291,N_10412);
xor U10642 (N_10642,N_10114,N_10544);
and U10643 (N_10643,N_10223,N_10117);
xnor U10644 (N_10644,N_10408,N_10012);
xnor U10645 (N_10645,N_10049,N_10455);
xnor U10646 (N_10646,N_10307,N_10621);
and U10647 (N_10647,N_10176,N_10301);
or U10648 (N_10648,N_10331,N_10249);
nor U10649 (N_10649,N_10609,N_10024);
or U10650 (N_10650,N_10622,N_10187);
or U10651 (N_10651,N_10484,N_10155);
or U10652 (N_10652,N_10136,N_10603);
or U10653 (N_10653,N_10497,N_10539);
and U10654 (N_10654,N_10557,N_10063);
nor U10655 (N_10655,N_10146,N_10202);
and U10656 (N_10656,N_10115,N_10343);
or U10657 (N_10657,N_10189,N_10161);
or U10658 (N_10658,N_10243,N_10498);
and U10659 (N_10659,N_10342,N_10066);
or U10660 (N_10660,N_10555,N_10207);
xnor U10661 (N_10661,N_10043,N_10444);
or U10662 (N_10662,N_10507,N_10569);
xor U10663 (N_10663,N_10275,N_10060);
xor U10664 (N_10664,N_10298,N_10001);
and U10665 (N_10665,N_10350,N_10047);
nor U10666 (N_10666,N_10104,N_10011);
xor U10667 (N_10667,N_10283,N_10052);
nand U10668 (N_10668,N_10567,N_10378);
xnor U10669 (N_10669,N_10006,N_10604);
nand U10670 (N_10670,N_10304,N_10272);
and U10671 (N_10671,N_10404,N_10510);
or U10672 (N_10672,N_10356,N_10328);
xnor U10673 (N_10673,N_10322,N_10584);
or U10674 (N_10674,N_10222,N_10113);
xnor U10675 (N_10675,N_10366,N_10396);
nand U10676 (N_10676,N_10565,N_10125);
xor U10677 (N_10677,N_10137,N_10605);
nand U10678 (N_10678,N_10613,N_10421);
and U10679 (N_10679,N_10261,N_10542);
or U10680 (N_10680,N_10418,N_10094);
nor U10681 (N_10681,N_10279,N_10405);
and U10682 (N_10682,N_10167,N_10437);
xor U10683 (N_10683,N_10305,N_10061);
xor U10684 (N_10684,N_10382,N_10074);
or U10685 (N_10685,N_10281,N_10205);
nand U10686 (N_10686,N_10217,N_10116);
and U10687 (N_10687,N_10502,N_10025);
nand U10688 (N_10688,N_10314,N_10320);
or U10689 (N_10689,N_10540,N_10129);
xnor U10690 (N_10690,N_10563,N_10581);
or U10691 (N_10691,N_10135,N_10463);
and U10692 (N_10692,N_10435,N_10461);
nor U10693 (N_10693,N_10282,N_10588);
and U10694 (N_10694,N_10329,N_10144);
or U10695 (N_10695,N_10427,N_10193);
and U10696 (N_10696,N_10485,N_10601);
nor U10697 (N_10697,N_10124,N_10589);
and U10698 (N_10698,N_10000,N_10364);
xor U10699 (N_10699,N_10219,N_10624);
nor U10700 (N_10700,N_10494,N_10492);
or U10701 (N_10701,N_10109,N_10562);
xor U10702 (N_10702,N_10260,N_10310);
and U10703 (N_10703,N_10186,N_10262);
and U10704 (N_10704,N_10376,N_10140);
and U10705 (N_10705,N_10500,N_10442);
xnor U10706 (N_10706,N_10375,N_10379);
nor U10707 (N_10707,N_10248,N_10608);
and U10708 (N_10708,N_10091,N_10058);
nand U10709 (N_10709,N_10531,N_10355);
and U10710 (N_10710,N_10600,N_10577);
nand U10711 (N_10711,N_10230,N_10602);
and U10712 (N_10712,N_10290,N_10570);
and U10713 (N_10713,N_10481,N_10341);
or U10714 (N_10714,N_10332,N_10587);
xnor U10715 (N_10715,N_10623,N_10452);
xnor U10716 (N_10716,N_10572,N_10118);
nand U10717 (N_10717,N_10050,N_10321);
and U10718 (N_10718,N_10126,N_10289);
xor U10719 (N_10719,N_10560,N_10415);
xor U10720 (N_10720,N_10607,N_10299);
nor U10721 (N_10721,N_10468,N_10547);
nor U10722 (N_10722,N_10175,N_10559);
or U10723 (N_10723,N_10130,N_10259);
or U10724 (N_10724,N_10029,N_10111);
and U10725 (N_10725,N_10346,N_10285);
and U10726 (N_10726,N_10534,N_10392);
and U10727 (N_10727,N_10466,N_10288);
and U10728 (N_10728,N_10537,N_10218);
xor U10729 (N_10729,N_10402,N_10151);
or U10730 (N_10730,N_10546,N_10294);
or U10731 (N_10731,N_10267,N_10513);
or U10732 (N_10732,N_10076,N_10070);
and U10733 (N_10733,N_10456,N_10423);
xor U10734 (N_10734,N_10016,N_10480);
nor U10735 (N_10735,N_10286,N_10048);
nand U10736 (N_10736,N_10348,N_10361);
and U10737 (N_10737,N_10514,N_10270);
xnor U10738 (N_10738,N_10169,N_10334);
and U10739 (N_10739,N_10420,N_10578);
or U10740 (N_10740,N_10028,N_10154);
xnor U10741 (N_10741,N_10457,N_10441);
and U10742 (N_10742,N_10393,N_10191);
nand U10743 (N_10743,N_10010,N_10429);
and U10744 (N_10744,N_10178,N_10323);
or U10745 (N_10745,N_10386,N_10422);
nand U10746 (N_10746,N_10065,N_10571);
nor U10747 (N_10747,N_10564,N_10019);
nor U10748 (N_10748,N_10236,N_10073);
xor U10749 (N_10749,N_10524,N_10145);
nor U10750 (N_10750,N_10095,N_10345);
xor U10751 (N_10751,N_10170,N_10293);
or U10752 (N_10752,N_10459,N_10177);
xnor U10753 (N_10753,N_10295,N_10088);
and U10754 (N_10754,N_10265,N_10590);
and U10755 (N_10755,N_10034,N_10264);
or U10756 (N_10756,N_10520,N_10287);
and U10757 (N_10757,N_10159,N_10319);
and U10758 (N_10758,N_10398,N_10042);
and U10759 (N_10759,N_10004,N_10183);
nand U10760 (N_10760,N_10383,N_10394);
or U10761 (N_10761,N_10142,N_10210);
nand U10762 (N_10762,N_10020,N_10399);
or U10763 (N_10763,N_10054,N_10610);
xor U10764 (N_10764,N_10228,N_10072);
and U10765 (N_10765,N_10548,N_10106);
nand U10766 (N_10766,N_10119,N_10045);
or U10767 (N_10767,N_10244,N_10495);
nand U10768 (N_10768,N_10018,N_10414);
nand U10769 (N_10769,N_10164,N_10253);
xnor U10770 (N_10770,N_10273,N_10612);
or U10771 (N_10771,N_10211,N_10445);
xor U10772 (N_10772,N_10450,N_10168);
nor U10773 (N_10773,N_10201,N_10357);
or U10774 (N_10774,N_10204,N_10580);
nor U10775 (N_10775,N_10416,N_10220);
nand U10776 (N_10776,N_10338,N_10464);
or U10777 (N_10777,N_10215,N_10132);
nand U10778 (N_10778,N_10199,N_10092);
nor U10779 (N_10779,N_10369,N_10234);
nand U10780 (N_10780,N_10086,N_10527);
nor U10781 (N_10781,N_10340,N_10009);
xor U10782 (N_10782,N_10121,N_10083);
or U10783 (N_10783,N_10162,N_10311);
and U10784 (N_10784,N_10053,N_10384);
xnor U10785 (N_10785,N_10436,N_10258);
nor U10786 (N_10786,N_10166,N_10120);
xnor U10787 (N_10787,N_10216,N_10254);
nor U10788 (N_10788,N_10352,N_10362);
nor U10789 (N_10789,N_10532,N_10158);
and U10790 (N_10790,N_10595,N_10108);
nand U10791 (N_10791,N_10337,N_10098);
nor U10792 (N_10792,N_10424,N_10551);
or U10793 (N_10793,N_10071,N_10212);
nand U10794 (N_10794,N_10180,N_10105);
or U10795 (N_10795,N_10354,N_10561);
nor U10796 (N_10796,N_10160,N_10093);
nor U10797 (N_10797,N_10472,N_10380);
nor U10798 (N_10798,N_10242,N_10079);
xor U10799 (N_10799,N_10411,N_10333);
nor U10800 (N_10800,N_10078,N_10153);
or U10801 (N_10801,N_10489,N_10451);
nor U10802 (N_10802,N_10476,N_10479);
or U10803 (N_10803,N_10250,N_10470);
and U10804 (N_10804,N_10543,N_10059);
nand U10805 (N_10805,N_10067,N_10017);
nand U10806 (N_10806,N_10505,N_10511);
nor U10807 (N_10807,N_10198,N_10147);
nand U10808 (N_10808,N_10224,N_10276);
xnor U10809 (N_10809,N_10255,N_10473);
and U10810 (N_10810,N_10553,N_10518);
nand U10811 (N_10811,N_10344,N_10475);
nand U10812 (N_10812,N_10454,N_10274);
or U10813 (N_10813,N_10064,N_10426);
and U10814 (N_10814,N_10616,N_10430);
or U10815 (N_10815,N_10406,N_10529);
nor U10816 (N_10816,N_10516,N_10339);
or U10817 (N_10817,N_10133,N_10008);
and U10818 (N_10818,N_10432,N_10315);
or U10819 (N_10819,N_10390,N_10038);
nand U10820 (N_10820,N_10002,N_10122);
or U10821 (N_10821,N_10040,N_10324);
and U10822 (N_10822,N_10309,N_10535);
nand U10823 (N_10823,N_10179,N_10139);
xor U10824 (N_10824,N_10438,N_10317);
nor U10825 (N_10825,N_10280,N_10549);
nor U10826 (N_10826,N_10611,N_10030);
and U10827 (N_10827,N_10128,N_10449);
and U10828 (N_10828,N_10150,N_10512);
or U10829 (N_10829,N_10051,N_10077);
nor U10830 (N_10830,N_10428,N_10431);
xnor U10831 (N_10831,N_10082,N_10231);
or U10832 (N_10832,N_10556,N_10141);
xnor U10833 (N_10833,N_10469,N_10353);
or U10834 (N_10834,N_10593,N_10617);
nand U10835 (N_10835,N_10358,N_10585);
and U10836 (N_10836,N_10530,N_10575);
and U10837 (N_10837,N_10620,N_10599);
nor U10838 (N_10838,N_10081,N_10509);
xor U10839 (N_10839,N_10413,N_10318);
or U10840 (N_10840,N_10172,N_10080);
nand U10841 (N_10841,N_10003,N_10097);
and U10842 (N_10842,N_10084,N_10107);
and U10843 (N_10843,N_10194,N_10127);
and U10844 (N_10844,N_10506,N_10185);
xnor U10845 (N_10845,N_10395,N_10316);
and U10846 (N_10846,N_10359,N_10443);
and U10847 (N_10847,N_10460,N_10574);
or U10848 (N_10848,N_10618,N_10022);
nand U10849 (N_10849,N_10138,N_10591);
xnor U10850 (N_10850,N_10519,N_10397);
and U10851 (N_10851,N_10488,N_10368);
and U10852 (N_10852,N_10410,N_10373);
xor U10853 (N_10853,N_10568,N_10477);
nor U10854 (N_10854,N_10586,N_10268);
or U10855 (N_10855,N_10184,N_10594);
xor U10856 (N_10856,N_10057,N_10583);
or U10857 (N_10857,N_10143,N_10227);
nor U10858 (N_10858,N_10296,N_10278);
nor U10859 (N_10859,N_10090,N_10232);
or U10860 (N_10860,N_10046,N_10388);
xor U10861 (N_10861,N_10112,N_10606);
nor U10862 (N_10862,N_10221,N_10313);
nand U10863 (N_10863,N_10525,N_10271);
xnor U10864 (N_10864,N_10229,N_10521);
and U10865 (N_10865,N_10440,N_10190);
or U10866 (N_10866,N_10303,N_10504);
or U10867 (N_10867,N_10062,N_10566);
nor U10868 (N_10868,N_10385,N_10203);
or U10869 (N_10869,N_10417,N_10173);
xnor U10870 (N_10870,N_10433,N_10099);
or U10871 (N_10871,N_10325,N_10501);
or U10872 (N_10872,N_10035,N_10200);
xor U10873 (N_10873,N_10089,N_10163);
nand U10874 (N_10874,N_10336,N_10157);
nor U10875 (N_10875,N_10188,N_10251);
and U10876 (N_10876,N_10508,N_10209);
or U10877 (N_10877,N_10068,N_10225);
and U10878 (N_10878,N_10598,N_10522);
or U10879 (N_10879,N_10447,N_10370);
nor U10880 (N_10880,N_10013,N_10523);
xor U10881 (N_10881,N_10075,N_10023);
nand U10882 (N_10882,N_10558,N_10409);
nor U10883 (N_10883,N_10087,N_10596);
nor U10884 (N_10884,N_10306,N_10181);
nand U10885 (N_10885,N_10387,N_10434);
or U10886 (N_10886,N_10246,N_10123);
nand U10887 (N_10887,N_10171,N_10041);
xor U10888 (N_10888,N_10100,N_10037);
and U10889 (N_10889,N_10326,N_10372);
and U10890 (N_10890,N_10536,N_10482);
or U10891 (N_10891,N_10597,N_10266);
nand U10892 (N_10892,N_10302,N_10056);
xnor U10893 (N_10893,N_10085,N_10493);
or U10894 (N_10894,N_10550,N_10103);
nor U10895 (N_10895,N_10615,N_10247);
or U10896 (N_10896,N_10446,N_10014);
nand U10897 (N_10897,N_10096,N_10365);
and U10898 (N_10898,N_10226,N_10619);
nor U10899 (N_10899,N_10448,N_10238);
nor U10900 (N_10900,N_10576,N_10538);
or U10901 (N_10901,N_10425,N_10528);
nor U10902 (N_10902,N_10335,N_10478);
nor U10903 (N_10903,N_10292,N_10245);
nand U10904 (N_10904,N_10360,N_10363);
and U10905 (N_10905,N_10327,N_10192);
or U10906 (N_10906,N_10182,N_10015);
nor U10907 (N_10907,N_10486,N_10471);
nand U10908 (N_10908,N_10213,N_10407);
xnor U10909 (N_10909,N_10515,N_10241);
nor U10910 (N_10910,N_10252,N_10517);
nand U10911 (N_10911,N_10027,N_10545);
nor U10912 (N_10912,N_10403,N_10036);
nor U10913 (N_10913,N_10439,N_10462);
nand U10914 (N_10914,N_10401,N_10208);
or U10915 (N_10915,N_10101,N_10582);
xnor U10916 (N_10916,N_10573,N_10039);
nand U10917 (N_10917,N_10490,N_10110);
or U10918 (N_10918,N_10102,N_10308);
nand U10919 (N_10919,N_10377,N_10347);
nand U10920 (N_10920,N_10044,N_10026);
xor U10921 (N_10921,N_10349,N_10474);
nor U10922 (N_10922,N_10033,N_10483);
or U10923 (N_10923,N_10391,N_10351);
nand U10924 (N_10924,N_10032,N_10237);
and U10925 (N_10925,N_10239,N_10240);
nor U10926 (N_10926,N_10007,N_10197);
xor U10927 (N_10927,N_10579,N_10541);
xor U10928 (N_10928,N_10148,N_10257);
xor U10929 (N_10929,N_10458,N_10149);
or U10930 (N_10930,N_10055,N_10206);
or U10931 (N_10931,N_10005,N_10400);
and U10932 (N_10932,N_10554,N_10526);
nand U10933 (N_10933,N_10235,N_10196);
or U10934 (N_10934,N_10277,N_10419);
xor U10935 (N_10935,N_10503,N_10269);
nand U10936 (N_10936,N_10499,N_10300);
or U10937 (N_10937,N_10533,N_10242);
and U10938 (N_10938,N_10096,N_10445);
or U10939 (N_10939,N_10126,N_10249);
xnor U10940 (N_10940,N_10002,N_10605);
nor U10941 (N_10941,N_10424,N_10498);
xor U10942 (N_10942,N_10055,N_10043);
nor U10943 (N_10943,N_10566,N_10025);
xnor U10944 (N_10944,N_10271,N_10326);
nand U10945 (N_10945,N_10013,N_10289);
or U10946 (N_10946,N_10517,N_10612);
and U10947 (N_10947,N_10515,N_10278);
nand U10948 (N_10948,N_10475,N_10511);
or U10949 (N_10949,N_10037,N_10160);
nor U10950 (N_10950,N_10540,N_10080);
or U10951 (N_10951,N_10155,N_10593);
nand U10952 (N_10952,N_10045,N_10025);
or U10953 (N_10953,N_10143,N_10421);
or U10954 (N_10954,N_10374,N_10588);
xnor U10955 (N_10955,N_10453,N_10398);
xor U10956 (N_10956,N_10170,N_10151);
and U10957 (N_10957,N_10267,N_10312);
nand U10958 (N_10958,N_10138,N_10515);
nor U10959 (N_10959,N_10013,N_10253);
nor U10960 (N_10960,N_10323,N_10244);
nand U10961 (N_10961,N_10011,N_10584);
xnor U10962 (N_10962,N_10103,N_10614);
nor U10963 (N_10963,N_10372,N_10381);
and U10964 (N_10964,N_10204,N_10179);
xnor U10965 (N_10965,N_10163,N_10367);
nand U10966 (N_10966,N_10412,N_10338);
or U10967 (N_10967,N_10424,N_10615);
nor U10968 (N_10968,N_10280,N_10199);
xor U10969 (N_10969,N_10398,N_10032);
and U10970 (N_10970,N_10341,N_10302);
or U10971 (N_10971,N_10261,N_10288);
nor U10972 (N_10972,N_10452,N_10151);
or U10973 (N_10973,N_10425,N_10598);
nor U10974 (N_10974,N_10171,N_10057);
and U10975 (N_10975,N_10525,N_10079);
xnor U10976 (N_10976,N_10062,N_10461);
or U10977 (N_10977,N_10100,N_10175);
xnor U10978 (N_10978,N_10500,N_10055);
nor U10979 (N_10979,N_10398,N_10321);
and U10980 (N_10980,N_10459,N_10251);
nor U10981 (N_10981,N_10384,N_10238);
and U10982 (N_10982,N_10494,N_10019);
nand U10983 (N_10983,N_10265,N_10467);
or U10984 (N_10984,N_10613,N_10541);
nor U10985 (N_10985,N_10546,N_10081);
or U10986 (N_10986,N_10566,N_10512);
and U10987 (N_10987,N_10289,N_10302);
or U10988 (N_10988,N_10191,N_10057);
xor U10989 (N_10989,N_10437,N_10604);
xnor U10990 (N_10990,N_10586,N_10000);
nor U10991 (N_10991,N_10252,N_10131);
nor U10992 (N_10992,N_10247,N_10328);
nand U10993 (N_10993,N_10376,N_10433);
nand U10994 (N_10994,N_10004,N_10386);
and U10995 (N_10995,N_10532,N_10266);
nand U10996 (N_10996,N_10263,N_10612);
and U10997 (N_10997,N_10341,N_10088);
nand U10998 (N_10998,N_10470,N_10202);
and U10999 (N_10999,N_10534,N_10524);
and U11000 (N_11000,N_10368,N_10603);
and U11001 (N_11001,N_10399,N_10420);
xor U11002 (N_11002,N_10507,N_10302);
and U11003 (N_11003,N_10501,N_10001);
and U11004 (N_11004,N_10522,N_10615);
or U11005 (N_11005,N_10027,N_10521);
nand U11006 (N_11006,N_10615,N_10596);
xnor U11007 (N_11007,N_10136,N_10122);
or U11008 (N_11008,N_10269,N_10105);
xor U11009 (N_11009,N_10018,N_10245);
nor U11010 (N_11010,N_10206,N_10049);
nand U11011 (N_11011,N_10517,N_10189);
nand U11012 (N_11012,N_10375,N_10089);
or U11013 (N_11013,N_10174,N_10096);
xnor U11014 (N_11014,N_10322,N_10124);
and U11015 (N_11015,N_10043,N_10124);
or U11016 (N_11016,N_10232,N_10144);
or U11017 (N_11017,N_10061,N_10398);
nand U11018 (N_11018,N_10236,N_10281);
nand U11019 (N_11019,N_10007,N_10357);
or U11020 (N_11020,N_10543,N_10100);
or U11021 (N_11021,N_10291,N_10295);
or U11022 (N_11022,N_10560,N_10516);
and U11023 (N_11023,N_10266,N_10039);
or U11024 (N_11024,N_10323,N_10030);
nand U11025 (N_11025,N_10353,N_10381);
nor U11026 (N_11026,N_10188,N_10462);
nand U11027 (N_11027,N_10027,N_10605);
or U11028 (N_11028,N_10533,N_10495);
xnor U11029 (N_11029,N_10068,N_10368);
nor U11030 (N_11030,N_10295,N_10153);
nand U11031 (N_11031,N_10568,N_10308);
or U11032 (N_11032,N_10394,N_10370);
nand U11033 (N_11033,N_10446,N_10111);
nand U11034 (N_11034,N_10413,N_10164);
nor U11035 (N_11035,N_10425,N_10420);
nor U11036 (N_11036,N_10009,N_10507);
or U11037 (N_11037,N_10292,N_10059);
nand U11038 (N_11038,N_10199,N_10513);
nand U11039 (N_11039,N_10079,N_10445);
nand U11040 (N_11040,N_10298,N_10469);
nand U11041 (N_11041,N_10336,N_10360);
or U11042 (N_11042,N_10078,N_10414);
nor U11043 (N_11043,N_10493,N_10510);
and U11044 (N_11044,N_10500,N_10308);
and U11045 (N_11045,N_10391,N_10152);
and U11046 (N_11046,N_10175,N_10243);
nand U11047 (N_11047,N_10599,N_10421);
nor U11048 (N_11048,N_10234,N_10125);
xnor U11049 (N_11049,N_10518,N_10511);
nand U11050 (N_11050,N_10440,N_10341);
nor U11051 (N_11051,N_10097,N_10356);
xnor U11052 (N_11052,N_10511,N_10394);
nand U11053 (N_11053,N_10023,N_10251);
xor U11054 (N_11054,N_10536,N_10499);
nand U11055 (N_11055,N_10485,N_10589);
and U11056 (N_11056,N_10122,N_10462);
xor U11057 (N_11057,N_10161,N_10142);
nand U11058 (N_11058,N_10223,N_10589);
xor U11059 (N_11059,N_10223,N_10324);
nand U11060 (N_11060,N_10260,N_10348);
or U11061 (N_11061,N_10165,N_10429);
nor U11062 (N_11062,N_10036,N_10607);
nor U11063 (N_11063,N_10346,N_10492);
xor U11064 (N_11064,N_10342,N_10295);
and U11065 (N_11065,N_10194,N_10018);
nand U11066 (N_11066,N_10274,N_10559);
xnor U11067 (N_11067,N_10343,N_10580);
xor U11068 (N_11068,N_10098,N_10193);
nor U11069 (N_11069,N_10332,N_10065);
xor U11070 (N_11070,N_10537,N_10480);
xor U11071 (N_11071,N_10240,N_10584);
nand U11072 (N_11072,N_10419,N_10071);
nor U11073 (N_11073,N_10089,N_10403);
or U11074 (N_11074,N_10243,N_10041);
or U11075 (N_11075,N_10543,N_10286);
nand U11076 (N_11076,N_10099,N_10436);
xnor U11077 (N_11077,N_10331,N_10326);
nand U11078 (N_11078,N_10291,N_10466);
and U11079 (N_11079,N_10460,N_10570);
nor U11080 (N_11080,N_10266,N_10359);
or U11081 (N_11081,N_10313,N_10075);
and U11082 (N_11082,N_10183,N_10396);
nor U11083 (N_11083,N_10339,N_10347);
nor U11084 (N_11084,N_10169,N_10430);
or U11085 (N_11085,N_10132,N_10539);
nand U11086 (N_11086,N_10435,N_10174);
nand U11087 (N_11087,N_10502,N_10000);
nand U11088 (N_11088,N_10181,N_10194);
nand U11089 (N_11089,N_10427,N_10064);
xor U11090 (N_11090,N_10394,N_10444);
nand U11091 (N_11091,N_10387,N_10619);
and U11092 (N_11092,N_10167,N_10286);
nand U11093 (N_11093,N_10245,N_10445);
nand U11094 (N_11094,N_10319,N_10258);
or U11095 (N_11095,N_10045,N_10061);
nand U11096 (N_11096,N_10452,N_10210);
and U11097 (N_11097,N_10364,N_10464);
nand U11098 (N_11098,N_10104,N_10595);
nor U11099 (N_11099,N_10277,N_10465);
nand U11100 (N_11100,N_10425,N_10390);
nor U11101 (N_11101,N_10280,N_10346);
nand U11102 (N_11102,N_10044,N_10439);
or U11103 (N_11103,N_10608,N_10572);
nand U11104 (N_11104,N_10367,N_10056);
xor U11105 (N_11105,N_10304,N_10175);
or U11106 (N_11106,N_10239,N_10126);
nor U11107 (N_11107,N_10217,N_10560);
or U11108 (N_11108,N_10598,N_10378);
nand U11109 (N_11109,N_10331,N_10026);
or U11110 (N_11110,N_10446,N_10101);
nand U11111 (N_11111,N_10475,N_10304);
and U11112 (N_11112,N_10549,N_10350);
and U11113 (N_11113,N_10166,N_10153);
and U11114 (N_11114,N_10360,N_10172);
or U11115 (N_11115,N_10065,N_10434);
nor U11116 (N_11116,N_10233,N_10615);
nor U11117 (N_11117,N_10155,N_10430);
and U11118 (N_11118,N_10588,N_10498);
and U11119 (N_11119,N_10127,N_10226);
xor U11120 (N_11120,N_10048,N_10129);
nand U11121 (N_11121,N_10108,N_10443);
or U11122 (N_11122,N_10455,N_10454);
and U11123 (N_11123,N_10064,N_10553);
and U11124 (N_11124,N_10386,N_10501);
xnor U11125 (N_11125,N_10230,N_10084);
and U11126 (N_11126,N_10460,N_10186);
nor U11127 (N_11127,N_10343,N_10420);
and U11128 (N_11128,N_10124,N_10612);
nor U11129 (N_11129,N_10358,N_10551);
nor U11130 (N_11130,N_10599,N_10027);
xor U11131 (N_11131,N_10002,N_10140);
nor U11132 (N_11132,N_10517,N_10122);
and U11133 (N_11133,N_10008,N_10083);
nor U11134 (N_11134,N_10218,N_10456);
nor U11135 (N_11135,N_10547,N_10624);
nand U11136 (N_11136,N_10400,N_10445);
nand U11137 (N_11137,N_10188,N_10147);
xor U11138 (N_11138,N_10579,N_10032);
or U11139 (N_11139,N_10471,N_10075);
or U11140 (N_11140,N_10349,N_10123);
xor U11141 (N_11141,N_10040,N_10104);
xnor U11142 (N_11142,N_10499,N_10594);
nor U11143 (N_11143,N_10169,N_10267);
xnor U11144 (N_11144,N_10216,N_10366);
nor U11145 (N_11145,N_10275,N_10334);
nand U11146 (N_11146,N_10577,N_10173);
nand U11147 (N_11147,N_10497,N_10430);
and U11148 (N_11148,N_10134,N_10561);
xor U11149 (N_11149,N_10008,N_10079);
or U11150 (N_11150,N_10126,N_10180);
and U11151 (N_11151,N_10022,N_10565);
and U11152 (N_11152,N_10347,N_10380);
nand U11153 (N_11153,N_10461,N_10362);
nor U11154 (N_11154,N_10196,N_10367);
or U11155 (N_11155,N_10039,N_10376);
xor U11156 (N_11156,N_10344,N_10260);
or U11157 (N_11157,N_10260,N_10427);
xnor U11158 (N_11158,N_10098,N_10232);
nand U11159 (N_11159,N_10522,N_10502);
nand U11160 (N_11160,N_10136,N_10204);
xor U11161 (N_11161,N_10149,N_10493);
nor U11162 (N_11162,N_10027,N_10179);
nor U11163 (N_11163,N_10519,N_10406);
or U11164 (N_11164,N_10120,N_10320);
nor U11165 (N_11165,N_10407,N_10245);
nor U11166 (N_11166,N_10304,N_10246);
nor U11167 (N_11167,N_10101,N_10518);
nand U11168 (N_11168,N_10005,N_10159);
nand U11169 (N_11169,N_10025,N_10610);
and U11170 (N_11170,N_10470,N_10403);
nand U11171 (N_11171,N_10470,N_10156);
nor U11172 (N_11172,N_10336,N_10522);
nor U11173 (N_11173,N_10463,N_10439);
xnor U11174 (N_11174,N_10403,N_10603);
and U11175 (N_11175,N_10362,N_10569);
nand U11176 (N_11176,N_10464,N_10552);
nor U11177 (N_11177,N_10449,N_10050);
and U11178 (N_11178,N_10083,N_10318);
xnor U11179 (N_11179,N_10225,N_10180);
xor U11180 (N_11180,N_10124,N_10073);
xor U11181 (N_11181,N_10595,N_10375);
xnor U11182 (N_11182,N_10425,N_10401);
and U11183 (N_11183,N_10050,N_10196);
nor U11184 (N_11184,N_10460,N_10274);
nor U11185 (N_11185,N_10301,N_10353);
and U11186 (N_11186,N_10090,N_10380);
nand U11187 (N_11187,N_10021,N_10050);
nand U11188 (N_11188,N_10051,N_10305);
nand U11189 (N_11189,N_10143,N_10471);
and U11190 (N_11190,N_10485,N_10367);
nand U11191 (N_11191,N_10566,N_10465);
or U11192 (N_11192,N_10234,N_10300);
nor U11193 (N_11193,N_10263,N_10602);
and U11194 (N_11194,N_10035,N_10538);
xnor U11195 (N_11195,N_10380,N_10611);
or U11196 (N_11196,N_10476,N_10596);
xor U11197 (N_11197,N_10270,N_10090);
or U11198 (N_11198,N_10284,N_10565);
nand U11199 (N_11199,N_10312,N_10129);
nor U11200 (N_11200,N_10413,N_10368);
nor U11201 (N_11201,N_10576,N_10561);
and U11202 (N_11202,N_10292,N_10503);
and U11203 (N_11203,N_10092,N_10240);
nand U11204 (N_11204,N_10522,N_10589);
xnor U11205 (N_11205,N_10056,N_10528);
and U11206 (N_11206,N_10322,N_10116);
and U11207 (N_11207,N_10384,N_10557);
and U11208 (N_11208,N_10018,N_10169);
and U11209 (N_11209,N_10388,N_10532);
nand U11210 (N_11210,N_10400,N_10394);
xnor U11211 (N_11211,N_10526,N_10509);
and U11212 (N_11212,N_10088,N_10535);
and U11213 (N_11213,N_10348,N_10331);
nor U11214 (N_11214,N_10541,N_10036);
nand U11215 (N_11215,N_10228,N_10094);
nand U11216 (N_11216,N_10066,N_10223);
and U11217 (N_11217,N_10028,N_10504);
nor U11218 (N_11218,N_10515,N_10557);
and U11219 (N_11219,N_10158,N_10617);
nor U11220 (N_11220,N_10349,N_10572);
nor U11221 (N_11221,N_10544,N_10543);
nor U11222 (N_11222,N_10082,N_10204);
and U11223 (N_11223,N_10144,N_10434);
nand U11224 (N_11224,N_10110,N_10279);
and U11225 (N_11225,N_10429,N_10132);
and U11226 (N_11226,N_10373,N_10197);
nor U11227 (N_11227,N_10014,N_10402);
nand U11228 (N_11228,N_10350,N_10364);
or U11229 (N_11229,N_10259,N_10378);
and U11230 (N_11230,N_10456,N_10036);
xor U11231 (N_11231,N_10417,N_10022);
and U11232 (N_11232,N_10106,N_10047);
or U11233 (N_11233,N_10135,N_10338);
nand U11234 (N_11234,N_10468,N_10259);
and U11235 (N_11235,N_10436,N_10231);
and U11236 (N_11236,N_10487,N_10410);
nor U11237 (N_11237,N_10197,N_10012);
nand U11238 (N_11238,N_10470,N_10535);
nand U11239 (N_11239,N_10298,N_10208);
nor U11240 (N_11240,N_10581,N_10514);
nand U11241 (N_11241,N_10272,N_10081);
or U11242 (N_11242,N_10550,N_10105);
nor U11243 (N_11243,N_10594,N_10615);
or U11244 (N_11244,N_10390,N_10593);
and U11245 (N_11245,N_10167,N_10244);
and U11246 (N_11246,N_10143,N_10270);
and U11247 (N_11247,N_10000,N_10167);
nor U11248 (N_11248,N_10399,N_10516);
or U11249 (N_11249,N_10589,N_10508);
nor U11250 (N_11250,N_11130,N_11042);
xnor U11251 (N_11251,N_10791,N_10935);
xnor U11252 (N_11252,N_11020,N_10788);
and U11253 (N_11253,N_11024,N_10975);
or U11254 (N_11254,N_11086,N_10685);
or U11255 (N_11255,N_11058,N_10989);
xnor U11256 (N_11256,N_10814,N_11137);
xor U11257 (N_11257,N_11126,N_11098);
nand U11258 (N_11258,N_10742,N_10886);
nand U11259 (N_11259,N_10993,N_10775);
nand U11260 (N_11260,N_11049,N_10729);
or U11261 (N_11261,N_11139,N_11050);
nand U11262 (N_11262,N_10896,N_10837);
nor U11263 (N_11263,N_11189,N_11048);
and U11264 (N_11264,N_10626,N_11116);
or U11265 (N_11265,N_11009,N_11145);
nor U11266 (N_11266,N_10759,N_11125);
or U11267 (N_11267,N_10924,N_10855);
xnor U11268 (N_11268,N_11207,N_10877);
and U11269 (N_11269,N_11103,N_11008);
and U11270 (N_11270,N_10998,N_10833);
nand U11271 (N_11271,N_11117,N_10981);
nand U11272 (N_11272,N_10789,N_11151);
nor U11273 (N_11273,N_11065,N_10724);
and U11274 (N_11274,N_10779,N_10867);
nor U11275 (N_11275,N_11108,N_11053);
xor U11276 (N_11276,N_10658,N_10909);
xnor U11277 (N_11277,N_11107,N_11224);
nand U11278 (N_11278,N_11032,N_10634);
nand U11279 (N_11279,N_10978,N_10915);
xor U11280 (N_11280,N_11028,N_10891);
nand U11281 (N_11281,N_11027,N_10693);
nand U11282 (N_11282,N_11011,N_11233);
nand U11283 (N_11283,N_10838,N_11242);
or U11284 (N_11284,N_10986,N_10848);
and U11285 (N_11285,N_11182,N_11169);
nand U11286 (N_11286,N_10962,N_11121);
nand U11287 (N_11287,N_10919,N_11093);
nor U11288 (N_11288,N_11101,N_10827);
nand U11289 (N_11289,N_10644,N_11016);
and U11290 (N_11290,N_10763,N_10912);
xnor U11291 (N_11291,N_10799,N_11148);
xor U11292 (N_11292,N_11179,N_11076);
nand U11293 (N_11293,N_10839,N_10632);
xor U11294 (N_11294,N_11160,N_11128);
nand U11295 (N_11295,N_10996,N_10860);
xnor U11296 (N_11296,N_10670,N_10942);
nor U11297 (N_11297,N_10653,N_10890);
or U11298 (N_11298,N_11085,N_10951);
nor U11299 (N_11299,N_10739,N_10790);
nor U11300 (N_11300,N_10657,N_11023);
or U11301 (N_11301,N_10899,N_10692);
or U11302 (N_11302,N_10805,N_11123);
nor U11303 (N_11303,N_10625,N_10948);
nand U11304 (N_11304,N_10917,N_11136);
nor U11305 (N_11305,N_10888,N_10647);
and U11306 (N_11306,N_10894,N_11246);
nor U11307 (N_11307,N_10771,N_11120);
nor U11308 (N_11308,N_11174,N_10711);
nand U11309 (N_11309,N_11010,N_10752);
nand U11310 (N_11310,N_11163,N_10728);
xnor U11311 (N_11311,N_11037,N_11188);
and U11312 (N_11312,N_11102,N_11007);
nand U11313 (N_11313,N_11134,N_11210);
nor U11314 (N_11314,N_10801,N_10684);
xnor U11315 (N_11315,N_10655,N_11190);
and U11316 (N_11316,N_10881,N_10803);
or U11317 (N_11317,N_11018,N_10770);
and U11318 (N_11318,N_10686,N_11031);
or U11319 (N_11319,N_10804,N_11014);
and U11320 (N_11320,N_11083,N_11026);
and U11321 (N_11321,N_11112,N_10941);
xnor U11322 (N_11322,N_10662,N_11132);
or U11323 (N_11323,N_10722,N_10979);
and U11324 (N_11324,N_11054,N_10883);
nand U11325 (N_11325,N_10635,N_10938);
nor U11326 (N_11326,N_10889,N_10636);
and U11327 (N_11327,N_11061,N_11229);
or U11328 (N_11328,N_10781,N_10806);
or U11329 (N_11329,N_10836,N_10908);
or U11330 (N_11330,N_10832,N_10664);
xor U11331 (N_11331,N_10776,N_11115);
xnor U11332 (N_11332,N_10800,N_11232);
nor U11333 (N_11333,N_11200,N_11039);
xnor U11334 (N_11334,N_10842,N_10920);
xnor U11335 (N_11335,N_10822,N_11127);
nor U11336 (N_11336,N_11034,N_11154);
xor U11337 (N_11337,N_10665,N_10965);
and U11338 (N_11338,N_10744,N_11144);
and U11339 (N_11339,N_10694,N_10982);
nor U11340 (N_11340,N_11041,N_10937);
nor U11341 (N_11341,N_11196,N_10817);
xor U11342 (N_11342,N_10631,N_10754);
xor U11343 (N_11343,N_11087,N_11118);
or U11344 (N_11344,N_10733,N_10701);
and U11345 (N_11345,N_10959,N_11149);
xnor U11346 (N_11346,N_10874,N_10892);
or U11347 (N_11347,N_10756,N_10731);
or U11348 (N_11348,N_11161,N_10679);
or U11349 (N_11349,N_10821,N_11124);
xor U11350 (N_11350,N_11077,N_10727);
and U11351 (N_11351,N_11140,N_10847);
nand U11352 (N_11352,N_10830,N_11216);
and U11353 (N_11353,N_10926,N_11156);
or U11354 (N_11354,N_11106,N_10627);
or U11355 (N_11355,N_10708,N_11045);
and U11356 (N_11356,N_11212,N_10649);
nand U11357 (N_11357,N_10699,N_11094);
and U11358 (N_11358,N_10650,N_10871);
xor U11359 (N_11359,N_11135,N_10936);
xnor U11360 (N_11360,N_10939,N_10787);
and U11361 (N_11361,N_11183,N_10835);
and U11362 (N_11362,N_10716,N_10897);
nand U11363 (N_11363,N_10648,N_10854);
nor U11364 (N_11364,N_10947,N_10667);
or U11365 (N_11365,N_11055,N_11243);
nor U11366 (N_11366,N_10726,N_10893);
or U11367 (N_11367,N_10755,N_11066);
and U11368 (N_11368,N_11063,N_10700);
xnor U11369 (N_11369,N_11131,N_10910);
and U11370 (N_11370,N_10849,N_10774);
nand U11371 (N_11371,N_10970,N_11003);
xor U11372 (N_11372,N_10902,N_11095);
and U11373 (N_11373,N_11173,N_10863);
nor U11374 (N_11374,N_10933,N_11238);
nand U11375 (N_11375,N_10639,N_11071);
nand U11376 (N_11376,N_10809,N_10977);
xnor U11377 (N_11377,N_11043,N_10741);
xnor U11378 (N_11378,N_10732,N_11064);
or U11379 (N_11379,N_10630,N_11244);
nor U11380 (N_11380,N_10844,N_10955);
or U11381 (N_11381,N_11180,N_11249);
nand U11382 (N_11382,N_11217,N_10918);
and U11383 (N_11383,N_10845,N_11158);
nor U11384 (N_11384,N_11165,N_10629);
nand U11385 (N_11385,N_10840,N_10654);
and U11386 (N_11386,N_10780,N_11172);
nor U11387 (N_11387,N_10683,N_10834);
nor U11388 (N_11388,N_11138,N_10786);
and U11389 (N_11389,N_11046,N_10905);
and U11390 (N_11390,N_10859,N_11100);
and U11391 (N_11391,N_11241,N_11090);
and U11392 (N_11392,N_10703,N_11060);
nand U11393 (N_11393,N_10702,N_10929);
nand U11394 (N_11394,N_10795,N_10813);
xnor U11395 (N_11395,N_10954,N_11091);
or U11396 (N_11396,N_11030,N_11167);
nor U11397 (N_11397,N_11035,N_11036);
nor U11398 (N_11398,N_11017,N_10802);
and U11399 (N_11399,N_10812,N_10972);
xnor U11400 (N_11400,N_11159,N_10995);
nor U11401 (N_11401,N_10829,N_10769);
or U11402 (N_11402,N_10641,N_11226);
nand U11403 (N_11403,N_11202,N_10946);
and U11404 (N_11404,N_10949,N_11067);
xor U11405 (N_11405,N_11062,N_10705);
nand U11406 (N_11406,N_10669,N_10944);
xor U11407 (N_11407,N_10868,N_10969);
nor U11408 (N_11408,N_10792,N_10778);
xor U11409 (N_11409,N_11203,N_11245);
nor U11410 (N_11410,N_10717,N_10968);
xnor U11411 (N_11411,N_10921,N_10735);
xnor U11412 (N_11412,N_10911,N_10676);
nor U11413 (N_11413,N_11199,N_10927);
or U11414 (N_11414,N_11022,N_10730);
nand U11415 (N_11415,N_11236,N_11015);
and U11416 (N_11416,N_10709,N_10678);
nand U11417 (N_11417,N_10747,N_10850);
or U11418 (N_11418,N_10828,N_11195);
or U11419 (N_11419,N_10913,N_10740);
nor U11420 (N_11420,N_11033,N_10643);
nand U11421 (N_11421,N_10857,N_10956);
nor U11422 (N_11422,N_10876,N_11143);
xor U11423 (N_11423,N_10677,N_11114);
xor U11424 (N_11424,N_11004,N_11038);
xor U11425 (N_11425,N_10807,N_10628);
nor U11426 (N_11426,N_10745,N_11168);
nand U11427 (N_11427,N_10691,N_11092);
or U11428 (N_11428,N_11070,N_10906);
and U11429 (N_11429,N_10777,N_10661);
nand U11430 (N_11430,N_11147,N_11240);
or U11431 (N_11431,N_10818,N_10736);
xnor U11432 (N_11432,N_10698,N_10760);
nand U11433 (N_11433,N_10858,N_10963);
or U11434 (N_11434,N_10922,N_11157);
and U11435 (N_11435,N_10971,N_10994);
or U11436 (N_11436,N_11150,N_10690);
xnor U11437 (N_11437,N_10797,N_11215);
nand U11438 (N_11438,N_11211,N_11084);
xnor U11439 (N_11439,N_11079,N_10875);
and U11440 (N_11440,N_10943,N_11186);
xor U11441 (N_11441,N_10825,N_10682);
and U11442 (N_11442,N_10967,N_10637);
or U11443 (N_11443,N_11142,N_10723);
nand U11444 (N_11444,N_10934,N_10898);
and U11445 (N_11445,N_10880,N_10695);
xor U11446 (N_11446,N_10932,N_10952);
nor U11447 (N_11447,N_10748,N_11237);
and U11448 (N_11448,N_10931,N_10707);
nand U11449 (N_11449,N_10879,N_10687);
or U11450 (N_11450,N_11080,N_11025);
nor U11451 (N_11451,N_10973,N_10900);
nor U11452 (N_11452,N_10988,N_11185);
nor U11453 (N_11453,N_10652,N_11214);
nand U11454 (N_11454,N_10895,N_10642);
or U11455 (N_11455,N_10697,N_10987);
and U11456 (N_11456,N_10816,N_10841);
nand U11457 (N_11457,N_11109,N_11047);
or U11458 (N_11458,N_10758,N_10925);
nor U11459 (N_11459,N_10671,N_10704);
xor U11460 (N_11460,N_11170,N_10718);
and U11461 (N_11461,N_10743,N_11164);
or U11462 (N_11462,N_11073,N_10945);
and U11463 (N_11463,N_11155,N_11228);
nor U11464 (N_11464,N_10864,N_10903);
and U11465 (N_11465,N_11175,N_11088);
xnor U11466 (N_11466,N_10870,N_10793);
nor U11467 (N_11467,N_10784,N_10633);
or U11468 (N_11468,N_11178,N_11122);
or U11469 (N_11469,N_10706,N_11069);
or U11470 (N_11470,N_10976,N_10843);
xor U11471 (N_11471,N_10734,N_10824);
or U11472 (N_11472,N_10980,N_10820);
nor U11473 (N_11473,N_11187,N_10646);
and U11474 (N_11474,N_10861,N_11113);
and U11475 (N_11475,N_10904,N_11052);
nand U11476 (N_11476,N_10940,N_10974);
and U11477 (N_11477,N_10826,N_11005);
xor U11478 (N_11478,N_10680,N_10907);
nor U11479 (N_11479,N_11074,N_10794);
and U11480 (N_11480,N_10985,N_10878);
xnor U11481 (N_11481,N_10992,N_11192);
nor U11482 (N_11482,N_10882,N_11089);
xor U11483 (N_11483,N_10961,N_11230);
or U11484 (N_11484,N_10872,N_11184);
and U11485 (N_11485,N_11248,N_10873);
and U11486 (N_11486,N_10668,N_10715);
nand U11487 (N_11487,N_11097,N_10689);
and U11488 (N_11488,N_11040,N_10983);
nor U11489 (N_11489,N_11082,N_11221);
nor U11490 (N_11490,N_11044,N_10785);
nand U11491 (N_11491,N_10765,N_11153);
nand U11492 (N_11492,N_10656,N_11162);
or U11493 (N_11493,N_10750,N_11078);
or U11494 (N_11494,N_11176,N_10681);
or U11495 (N_11495,N_10865,N_10960);
and U11496 (N_11496,N_10997,N_11218);
nor U11497 (N_11497,N_10966,N_11220);
or U11498 (N_11498,N_11213,N_10764);
or U11499 (N_11499,N_11225,N_11166);
and U11500 (N_11500,N_10749,N_10819);
nand U11501 (N_11501,N_11219,N_10719);
xor U11502 (N_11502,N_10768,N_10757);
and U11503 (N_11503,N_11208,N_11234);
and U11504 (N_11504,N_11068,N_10930);
or U11505 (N_11505,N_10866,N_10957);
xor U11506 (N_11506,N_11209,N_10796);
nand U11507 (N_11507,N_11222,N_11231);
nor U11508 (N_11508,N_11146,N_10991);
or U11509 (N_11509,N_11206,N_11194);
xnor U11510 (N_11510,N_10746,N_10885);
and U11511 (N_11511,N_11099,N_11006);
or U11512 (N_11512,N_10953,N_10713);
nor U11513 (N_11513,N_10811,N_10720);
xnor U11514 (N_11514,N_10710,N_11104);
or U11515 (N_11515,N_10901,N_10810);
or U11516 (N_11516,N_10928,N_11197);
or U11517 (N_11517,N_11205,N_11235);
or U11518 (N_11518,N_10914,N_10767);
or U11519 (N_11519,N_11081,N_10762);
and U11520 (N_11520,N_10651,N_11096);
nand U11521 (N_11521,N_11012,N_11177);
nand U11522 (N_11522,N_10712,N_10846);
nor U11523 (N_11523,N_11002,N_11110);
or U11524 (N_11524,N_11075,N_10660);
or U11525 (N_11525,N_10772,N_10761);
nand U11526 (N_11526,N_11129,N_10673);
and U11527 (N_11527,N_10688,N_10950);
xnor U11528 (N_11528,N_10725,N_11193);
nor U11529 (N_11529,N_10999,N_11227);
nor U11530 (N_11530,N_10659,N_10645);
nand U11531 (N_11531,N_10831,N_10853);
and U11532 (N_11532,N_10958,N_10887);
or U11533 (N_11533,N_10783,N_10852);
nand U11534 (N_11534,N_11223,N_10753);
xor U11535 (N_11535,N_11051,N_10990);
xor U11536 (N_11536,N_10666,N_11204);
and U11537 (N_11537,N_11111,N_10823);
nor U11538 (N_11538,N_10815,N_11201);
xor U11539 (N_11539,N_11105,N_10751);
nand U11540 (N_11540,N_10851,N_11072);
nand U11541 (N_11541,N_10674,N_11056);
nand U11542 (N_11542,N_11059,N_10798);
xor U11543 (N_11543,N_10663,N_10782);
xor U11544 (N_11544,N_11181,N_10672);
and U11545 (N_11545,N_10984,N_11013);
or U11546 (N_11546,N_10737,N_11152);
nand U11547 (N_11547,N_10721,N_10773);
xor U11548 (N_11548,N_10862,N_11133);
xnor U11549 (N_11549,N_10808,N_11029);
and U11550 (N_11550,N_11171,N_11000);
or U11551 (N_11551,N_10869,N_10856);
nor U11552 (N_11552,N_11198,N_11141);
or U11553 (N_11553,N_11239,N_11191);
and U11554 (N_11554,N_11247,N_10884);
nand U11555 (N_11555,N_11019,N_10766);
or U11556 (N_11556,N_10640,N_10696);
and U11557 (N_11557,N_10675,N_11057);
nand U11558 (N_11558,N_11119,N_10964);
xnor U11559 (N_11559,N_10738,N_10714);
nor U11560 (N_11560,N_10923,N_11021);
nand U11561 (N_11561,N_10916,N_10638);
nand U11562 (N_11562,N_11001,N_11030);
xnor U11563 (N_11563,N_10980,N_10763);
and U11564 (N_11564,N_10934,N_11082);
nor U11565 (N_11565,N_10676,N_11011);
and U11566 (N_11566,N_10711,N_10721);
or U11567 (N_11567,N_11180,N_10628);
nor U11568 (N_11568,N_10845,N_10951);
nand U11569 (N_11569,N_10821,N_10807);
and U11570 (N_11570,N_11030,N_10801);
or U11571 (N_11571,N_11132,N_10940);
nor U11572 (N_11572,N_11219,N_11221);
nand U11573 (N_11573,N_11105,N_10677);
xor U11574 (N_11574,N_10786,N_11176);
or U11575 (N_11575,N_11223,N_10904);
nand U11576 (N_11576,N_11172,N_10831);
and U11577 (N_11577,N_11145,N_10750);
or U11578 (N_11578,N_10715,N_10697);
nor U11579 (N_11579,N_10785,N_10849);
or U11580 (N_11580,N_11021,N_10661);
or U11581 (N_11581,N_11042,N_11004);
nand U11582 (N_11582,N_10727,N_11048);
nor U11583 (N_11583,N_11036,N_11163);
nor U11584 (N_11584,N_10727,N_10649);
nand U11585 (N_11585,N_10974,N_10792);
and U11586 (N_11586,N_10711,N_11237);
or U11587 (N_11587,N_10794,N_10886);
xor U11588 (N_11588,N_11211,N_11067);
and U11589 (N_11589,N_11132,N_11177);
nand U11590 (N_11590,N_11240,N_11175);
nand U11591 (N_11591,N_10673,N_10731);
nand U11592 (N_11592,N_11104,N_10636);
xor U11593 (N_11593,N_11024,N_10822);
nor U11594 (N_11594,N_10908,N_11218);
and U11595 (N_11595,N_11050,N_10686);
xor U11596 (N_11596,N_11226,N_10807);
and U11597 (N_11597,N_11115,N_10859);
nor U11598 (N_11598,N_10952,N_11165);
nor U11599 (N_11599,N_10701,N_10817);
and U11600 (N_11600,N_11031,N_10919);
nand U11601 (N_11601,N_10851,N_10809);
xor U11602 (N_11602,N_11018,N_10875);
xnor U11603 (N_11603,N_11230,N_10783);
xor U11604 (N_11604,N_10652,N_11087);
or U11605 (N_11605,N_10871,N_11019);
nor U11606 (N_11606,N_11246,N_10877);
and U11607 (N_11607,N_11172,N_11032);
and U11608 (N_11608,N_10752,N_10853);
nor U11609 (N_11609,N_10784,N_11141);
nor U11610 (N_11610,N_11113,N_11020);
xor U11611 (N_11611,N_10802,N_10996);
nor U11612 (N_11612,N_11168,N_10960);
nor U11613 (N_11613,N_11194,N_11122);
nand U11614 (N_11614,N_10743,N_10874);
nor U11615 (N_11615,N_11022,N_11082);
nor U11616 (N_11616,N_10761,N_10947);
or U11617 (N_11617,N_11070,N_10939);
nand U11618 (N_11618,N_10822,N_11136);
and U11619 (N_11619,N_10811,N_10952);
xnor U11620 (N_11620,N_10883,N_11226);
xor U11621 (N_11621,N_11068,N_11058);
and U11622 (N_11622,N_11195,N_10869);
xnor U11623 (N_11623,N_11118,N_10997);
xnor U11624 (N_11624,N_10981,N_10973);
xnor U11625 (N_11625,N_10712,N_10804);
nand U11626 (N_11626,N_11220,N_10891);
nor U11627 (N_11627,N_10940,N_10844);
nor U11628 (N_11628,N_11135,N_11106);
and U11629 (N_11629,N_11048,N_11139);
nor U11630 (N_11630,N_11212,N_11122);
nand U11631 (N_11631,N_11027,N_10801);
nor U11632 (N_11632,N_11062,N_11196);
and U11633 (N_11633,N_10949,N_11233);
nor U11634 (N_11634,N_11006,N_11151);
or U11635 (N_11635,N_10956,N_11072);
and U11636 (N_11636,N_10869,N_10772);
xor U11637 (N_11637,N_10779,N_10834);
nor U11638 (N_11638,N_10977,N_11107);
or U11639 (N_11639,N_10799,N_10938);
xnor U11640 (N_11640,N_11156,N_11091);
and U11641 (N_11641,N_10970,N_10725);
or U11642 (N_11642,N_10984,N_10849);
and U11643 (N_11643,N_11038,N_10902);
nand U11644 (N_11644,N_10969,N_10913);
nand U11645 (N_11645,N_10768,N_10955);
nand U11646 (N_11646,N_10698,N_10806);
xor U11647 (N_11647,N_11236,N_10922);
nand U11648 (N_11648,N_10996,N_10762);
and U11649 (N_11649,N_10960,N_11172);
nand U11650 (N_11650,N_10993,N_10784);
nand U11651 (N_11651,N_10700,N_11138);
and U11652 (N_11652,N_10868,N_10944);
nor U11653 (N_11653,N_11109,N_11137);
and U11654 (N_11654,N_10864,N_11163);
xor U11655 (N_11655,N_11229,N_11012);
or U11656 (N_11656,N_11017,N_10869);
and U11657 (N_11657,N_10870,N_10713);
or U11658 (N_11658,N_10626,N_10628);
nand U11659 (N_11659,N_10669,N_10886);
and U11660 (N_11660,N_11043,N_11115);
or U11661 (N_11661,N_10992,N_10984);
nand U11662 (N_11662,N_10667,N_11147);
xnor U11663 (N_11663,N_11167,N_10860);
and U11664 (N_11664,N_10914,N_11081);
and U11665 (N_11665,N_10868,N_11011);
nor U11666 (N_11666,N_10723,N_10671);
nand U11667 (N_11667,N_10925,N_10667);
nand U11668 (N_11668,N_11145,N_11010);
xor U11669 (N_11669,N_11194,N_10844);
or U11670 (N_11670,N_10745,N_10927);
and U11671 (N_11671,N_10741,N_11080);
nand U11672 (N_11672,N_10927,N_10877);
xor U11673 (N_11673,N_10900,N_10722);
and U11674 (N_11674,N_11000,N_11110);
or U11675 (N_11675,N_11239,N_11007);
nor U11676 (N_11676,N_10965,N_11179);
nand U11677 (N_11677,N_10747,N_11039);
nand U11678 (N_11678,N_10657,N_10938);
or U11679 (N_11679,N_10657,N_10834);
and U11680 (N_11680,N_10626,N_10653);
or U11681 (N_11681,N_11237,N_11194);
xor U11682 (N_11682,N_11084,N_11119);
and U11683 (N_11683,N_11220,N_10788);
nor U11684 (N_11684,N_10730,N_10751);
nor U11685 (N_11685,N_11246,N_10715);
nor U11686 (N_11686,N_11223,N_10822);
nor U11687 (N_11687,N_10630,N_10922);
and U11688 (N_11688,N_11183,N_11137);
and U11689 (N_11689,N_11004,N_11205);
nand U11690 (N_11690,N_10971,N_10906);
xnor U11691 (N_11691,N_10931,N_11022);
and U11692 (N_11692,N_10656,N_10926);
nand U11693 (N_11693,N_10809,N_10960);
and U11694 (N_11694,N_11157,N_10898);
xnor U11695 (N_11695,N_11125,N_10639);
nor U11696 (N_11696,N_10853,N_10709);
xor U11697 (N_11697,N_11181,N_10849);
or U11698 (N_11698,N_10758,N_10804);
nand U11699 (N_11699,N_10952,N_11127);
nand U11700 (N_11700,N_10739,N_10661);
nor U11701 (N_11701,N_10811,N_10764);
nand U11702 (N_11702,N_11027,N_11091);
nand U11703 (N_11703,N_10917,N_11150);
and U11704 (N_11704,N_10887,N_11031);
nand U11705 (N_11705,N_11043,N_10763);
xor U11706 (N_11706,N_10816,N_11178);
and U11707 (N_11707,N_11069,N_10626);
nor U11708 (N_11708,N_11015,N_11101);
xor U11709 (N_11709,N_11002,N_11232);
and U11710 (N_11710,N_10633,N_11106);
nand U11711 (N_11711,N_10759,N_11180);
nand U11712 (N_11712,N_11100,N_10634);
nand U11713 (N_11713,N_11140,N_11068);
nand U11714 (N_11714,N_10836,N_10634);
or U11715 (N_11715,N_11097,N_10724);
nand U11716 (N_11716,N_11230,N_11179);
xor U11717 (N_11717,N_11245,N_10745);
or U11718 (N_11718,N_11005,N_10968);
and U11719 (N_11719,N_10988,N_10917);
nand U11720 (N_11720,N_10937,N_10846);
or U11721 (N_11721,N_10860,N_10733);
nand U11722 (N_11722,N_10943,N_10917);
or U11723 (N_11723,N_10674,N_10758);
xnor U11724 (N_11724,N_10977,N_11152);
xor U11725 (N_11725,N_11131,N_10927);
xnor U11726 (N_11726,N_11118,N_11190);
or U11727 (N_11727,N_10912,N_11174);
and U11728 (N_11728,N_10958,N_11119);
or U11729 (N_11729,N_11223,N_11210);
nor U11730 (N_11730,N_10636,N_10716);
nand U11731 (N_11731,N_10635,N_10771);
or U11732 (N_11732,N_10767,N_10714);
nor U11733 (N_11733,N_10680,N_11142);
and U11734 (N_11734,N_10632,N_11123);
nand U11735 (N_11735,N_11163,N_11122);
xor U11736 (N_11736,N_10852,N_10706);
or U11737 (N_11737,N_11203,N_11042);
or U11738 (N_11738,N_11105,N_10691);
or U11739 (N_11739,N_10742,N_10896);
nor U11740 (N_11740,N_10866,N_11196);
xnor U11741 (N_11741,N_11162,N_11130);
xor U11742 (N_11742,N_11248,N_10725);
and U11743 (N_11743,N_11116,N_10874);
nand U11744 (N_11744,N_10981,N_11181);
or U11745 (N_11745,N_10880,N_11078);
nor U11746 (N_11746,N_10854,N_11128);
xor U11747 (N_11747,N_10868,N_10972);
xor U11748 (N_11748,N_11070,N_10757);
nand U11749 (N_11749,N_11243,N_10632);
nor U11750 (N_11750,N_10698,N_10865);
and U11751 (N_11751,N_11074,N_10735);
nor U11752 (N_11752,N_11209,N_10686);
or U11753 (N_11753,N_11195,N_11070);
and U11754 (N_11754,N_11174,N_11168);
xor U11755 (N_11755,N_11137,N_11126);
xor U11756 (N_11756,N_10633,N_10805);
nor U11757 (N_11757,N_10745,N_10955);
or U11758 (N_11758,N_11248,N_10705);
xor U11759 (N_11759,N_10944,N_11245);
xnor U11760 (N_11760,N_11025,N_10924);
nand U11761 (N_11761,N_11148,N_10959);
xnor U11762 (N_11762,N_11214,N_11141);
or U11763 (N_11763,N_10900,N_10920);
and U11764 (N_11764,N_11008,N_10900);
and U11765 (N_11765,N_11072,N_10653);
and U11766 (N_11766,N_10773,N_10627);
or U11767 (N_11767,N_10751,N_10944);
or U11768 (N_11768,N_10830,N_11007);
nor U11769 (N_11769,N_11016,N_11003);
nand U11770 (N_11770,N_11125,N_10786);
nand U11771 (N_11771,N_10989,N_11181);
nand U11772 (N_11772,N_11189,N_11179);
nor U11773 (N_11773,N_11025,N_11057);
or U11774 (N_11774,N_10830,N_11206);
nand U11775 (N_11775,N_10874,N_11210);
and U11776 (N_11776,N_11137,N_11020);
and U11777 (N_11777,N_10894,N_10804);
nor U11778 (N_11778,N_10773,N_11125);
or U11779 (N_11779,N_11082,N_10955);
or U11780 (N_11780,N_11047,N_10963);
nor U11781 (N_11781,N_10970,N_11149);
xor U11782 (N_11782,N_10841,N_10638);
or U11783 (N_11783,N_11180,N_10993);
nor U11784 (N_11784,N_10833,N_11028);
nand U11785 (N_11785,N_11116,N_10738);
and U11786 (N_11786,N_11177,N_10890);
and U11787 (N_11787,N_10864,N_10960);
nand U11788 (N_11788,N_10717,N_10890);
or U11789 (N_11789,N_11234,N_11019);
nand U11790 (N_11790,N_10773,N_10778);
or U11791 (N_11791,N_11208,N_11045);
nor U11792 (N_11792,N_11029,N_11159);
nor U11793 (N_11793,N_10893,N_11232);
nand U11794 (N_11794,N_10661,N_10907);
and U11795 (N_11795,N_10668,N_10812);
nand U11796 (N_11796,N_11145,N_11093);
nor U11797 (N_11797,N_10778,N_11096);
or U11798 (N_11798,N_10856,N_11085);
xor U11799 (N_11799,N_10995,N_10870);
nand U11800 (N_11800,N_10753,N_11091);
xnor U11801 (N_11801,N_11199,N_11139);
or U11802 (N_11802,N_10936,N_10654);
nand U11803 (N_11803,N_11187,N_10888);
or U11804 (N_11804,N_10702,N_11128);
nand U11805 (N_11805,N_10707,N_10873);
nor U11806 (N_11806,N_10647,N_10689);
and U11807 (N_11807,N_11214,N_11154);
nand U11808 (N_11808,N_10892,N_10828);
and U11809 (N_11809,N_10631,N_11150);
nand U11810 (N_11810,N_10946,N_10853);
and U11811 (N_11811,N_10712,N_10802);
nand U11812 (N_11812,N_10848,N_10660);
nand U11813 (N_11813,N_11142,N_10996);
nor U11814 (N_11814,N_11007,N_10894);
xnor U11815 (N_11815,N_11098,N_10724);
nor U11816 (N_11816,N_10729,N_10953);
nand U11817 (N_11817,N_10814,N_11154);
xor U11818 (N_11818,N_11049,N_10748);
xor U11819 (N_11819,N_11225,N_11019);
nor U11820 (N_11820,N_11246,N_11044);
nor U11821 (N_11821,N_10941,N_11175);
xor U11822 (N_11822,N_10782,N_10643);
xor U11823 (N_11823,N_10730,N_10728);
and U11824 (N_11824,N_10929,N_11183);
or U11825 (N_11825,N_11002,N_11047);
nor U11826 (N_11826,N_10761,N_10681);
and U11827 (N_11827,N_11157,N_10866);
or U11828 (N_11828,N_11060,N_10893);
or U11829 (N_11829,N_11180,N_10654);
xor U11830 (N_11830,N_10909,N_10646);
and U11831 (N_11831,N_10998,N_10965);
or U11832 (N_11832,N_10792,N_10829);
nand U11833 (N_11833,N_10863,N_10696);
nor U11834 (N_11834,N_11187,N_10751);
nand U11835 (N_11835,N_11086,N_10858);
nor U11836 (N_11836,N_10660,N_10837);
nand U11837 (N_11837,N_10756,N_11232);
nand U11838 (N_11838,N_10627,N_10662);
or U11839 (N_11839,N_10776,N_10675);
nor U11840 (N_11840,N_11176,N_11204);
and U11841 (N_11841,N_10956,N_10853);
and U11842 (N_11842,N_11183,N_10819);
nand U11843 (N_11843,N_10800,N_11125);
and U11844 (N_11844,N_11103,N_11134);
xor U11845 (N_11845,N_11102,N_10685);
nand U11846 (N_11846,N_10912,N_10811);
or U11847 (N_11847,N_10662,N_10636);
and U11848 (N_11848,N_11201,N_10981);
nand U11849 (N_11849,N_11013,N_10788);
nand U11850 (N_11850,N_11149,N_10804);
or U11851 (N_11851,N_10972,N_11067);
nor U11852 (N_11852,N_11162,N_11166);
xnor U11853 (N_11853,N_10937,N_10866);
xnor U11854 (N_11854,N_10769,N_10774);
nand U11855 (N_11855,N_10687,N_10790);
nand U11856 (N_11856,N_10666,N_10931);
and U11857 (N_11857,N_10897,N_11143);
xor U11858 (N_11858,N_11004,N_10637);
xnor U11859 (N_11859,N_10707,N_10998);
nand U11860 (N_11860,N_11140,N_11117);
nand U11861 (N_11861,N_10642,N_10706);
xnor U11862 (N_11862,N_10932,N_10725);
or U11863 (N_11863,N_10860,N_11204);
xor U11864 (N_11864,N_10746,N_11125);
nor U11865 (N_11865,N_10974,N_10626);
xor U11866 (N_11866,N_10984,N_10647);
nand U11867 (N_11867,N_10727,N_10953);
and U11868 (N_11868,N_10689,N_11055);
xnor U11869 (N_11869,N_10647,N_10761);
xor U11870 (N_11870,N_10754,N_10755);
xor U11871 (N_11871,N_11098,N_10828);
or U11872 (N_11872,N_10993,N_11000);
and U11873 (N_11873,N_10961,N_10921);
nand U11874 (N_11874,N_10629,N_10809);
or U11875 (N_11875,N_11394,N_11425);
nand U11876 (N_11876,N_11635,N_11250);
nand U11877 (N_11877,N_11252,N_11561);
nor U11878 (N_11878,N_11779,N_11822);
xnor U11879 (N_11879,N_11507,N_11293);
xor U11880 (N_11880,N_11782,N_11435);
xnor U11881 (N_11881,N_11688,N_11813);
and U11882 (N_11882,N_11473,N_11639);
nor U11883 (N_11883,N_11479,N_11644);
or U11884 (N_11884,N_11572,N_11613);
nand U11885 (N_11885,N_11254,N_11628);
xor U11886 (N_11886,N_11695,N_11570);
nor U11887 (N_11887,N_11777,N_11553);
or U11888 (N_11888,N_11275,N_11843);
xor U11889 (N_11889,N_11804,N_11638);
xnor U11890 (N_11890,N_11640,N_11512);
or U11891 (N_11891,N_11337,N_11461);
and U11892 (N_11892,N_11294,N_11456);
nand U11893 (N_11893,N_11606,N_11513);
and U11894 (N_11894,N_11632,N_11444);
xnor U11895 (N_11895,N_11370,N_11543);
xnor U11896 (N_11896,N_11710,N_11314);
nand U11897 (N_11897,N_11375,N_11298);
nand U11898 (N_11898,N_11812,N_11565);
nand U11899 (N_11899,N_11380,N_11746);
nand U11900 (N_11900,N_11492,N_11788);
nand U11901 (N_11901,N_11851,N_11622);
or U11902 (N_11902,N_11665,N_11516);
and U11903 (N_11903,N_11554,N_11750);
or U11904 (N_11904,N_11366,N_11723);
or U11905 (N_11905,N_11649,N_11608);
nand U11906 (N_11906,N_11534,N_11678);
and U11907 (N_11907,N_11302,N_11864);
nor U11908 (N_11908,N_11433,N_11675);
and U11909 (N_11909,N_11480,N_11481);
nor U11910 (N_11910,N_11815,N_11859);
nand U11911 (N_11911,N_11489,N_11576);
and U11912 (N_11912,N_11288,N_11765);
or U11913 (N_11913,N_11388,N_11797);
nand U11914 (N_11914,N_11369,N_11422);
nand U11915 (N_11915,N_11276,N_11354);
xor U11916 (N_11916,N_11588,N_11420);
nand U11917 (N_11917,N_11630,N_11817);
nand U11918 (N_11918,N_11872,N_11358);
xnor U11919 (N_11919,N_11826,N_11284);
xnor U11920 (N_11920,N_11615,N_11487);
xnor U11921 (N_11921,N_11407,N_11811);
nand U11922 (N_11922,N_11426,N_11263);
and U11923 (N_11923,N_11497,N_11629);
nor U11924 (N_11924,N_11373,N_11621);
nand U11925 (N_11925,N_11566,N_11690);
xnor U11926 (N_11926,N_11315,N_11463);
and U11927 (N_11927,N_11626,N_11620);
and U11928 (N_11928,N_11574,N_11273);
nor U11929 (N_11929,N_11790,N_11436);
xnor U11930 (N_11930,N_11339,N_11671);
nand U11931 (N_11931,N_11267,N_11795);
nor U11932 (N_11932,N_11532,N_11735);
and U11933 (N_11933,N_11274,N_11329);
nor U11934 (N_11934,N_11381,N_11331);
nand U11935 (N_11935,N_11345,N_11474);
nor U11936 (N_11936,N_11453,N_11819);
and U11937 (N_11937,N_11552,N_11696);
nor U11938 (N_11938,N_11564,N_11726);
or U11939 (N_11939,N_11402,N_11711);
nand U11940 (N_11940,N_11482,N_11457);
nor U11941 (N_11941,N_11742,N_11803);
and U11942 (N_11942,N_11837,N_11719);
nand U11943 (N_11943,N_11673,N_11770);
xnor U11944 (N_11944,N_11529,N_11762);
xor U11945 (N_11945,N_11736,N_11739);
xor U11946 (N_11946,N_11538,N_11557);
or U11947 (N_11947,N_11708,N_11292);
or U11948 (N_11948,N_11865,N_11705);
xnor U11949 (N_11949,N_11413,N_11547);
and U11950 (N_11950,N_11862,N_11856);
nor U11951 (N_11951,N_11344,N_11562);
or U11952 (N_11952,N_11443,N_11300);
or U11953 (N_11953,N_11858,N_11698);
and U11954 (N_11954,N_11661,N_11841);
and U11955 (N_11955,N_11336,N_11476);
nand U11956 (N_11956,N_11301,N_11351);
xor U11957 (N_11957,N_11521,N_11289);
or U11958 (N_11958,N_11799,N_11488);
and U11959 (N_11959,N_11801,N_11467);
or U11960 (N_11960,N_11501,N_11663);
or U11961 (N_11961,N_11846,N_11541);
xor U11962 (N_11962,N_11796,N_11597);
xnor U11963 (N_11963,N_11546,N_11328);
or U11964 (N_11964,N_11773,N_11763);
nand U11965 (N_11965,N_11401,N_11802);
nand U11966 (N_11966,N_11352,N_11692);
nor U11967 (N_11967,N_11338,N_11563);
nand U11968 (N_11968,N_11787,N_11262);
xor U11969 (N_11969,N_11485,N_11845);
or U11970 (N_11970,N_11585,N_11537);
or U11971 (N_11971,N_11468,N_11542);
or U11972 (N_11972,N_11737,N_11540);
or U11973 (N_11973,N_11775,N_11764);
and U11974 (N_11974,N_11504,N_11659);
nor U11975 (N_11975,N_11522,N_11636);
xnor U11976 (N_11976,N_11808,N_11399);
or U11977 (N_11977,N_11397,N_11838);
xnor U11978 (N_11978,N_11423,N_11580);
xnor U11979 (N_11979,N_11428,N_11486);
nand U11980 (N_11980,N_11367,N_11560);
xor U11981 (N_11981,N_11475,N_11556);
or U11982 (N_11982,N_11440,N_11449);
xnor U11983 (N_11983,N_11323,N_11596);
nor U11984 (N_11984,N_11438,N_11478);
nand U11985 (N_11985,N_11558,N_11785);
nor U11986 (N_11986,N_11519,N_11283);
and U11987 (N_11987,N_11450,N_11325);
nor U11988 (N_11988,N_11664,N_11748);
nor U11989 (N_11989,N_11469,N_11820);
nor U11990 (N_11990,N_11670,N_11386);
and U11991 (N_11991,N_11306,N_11310);
nand U11992 (N_11992,N_11860,N_11717);
or U11993 (N_11993,N_11729,N_11834);
nand U11994 (N_11994,N_11259,N_11569);
nor U11995 (N_11995,N_11725,N_11627);
xnor U11996 (N_11996,N_11732,N_11681);
nand U11997 (N_11997,N_11674,N_11848);
and U11998 (N_11998,N_11660,N_11322);
or U11999 (N_11999,N_11633,N_11609);
and U12000 (N_12000,N_11330,N_11494);
nand U12001 (N_12001,N_11571,N_11490);
xnor U12002 (N_12002,N_11704,N_11508);
nor U12003 (N_12003,N_11427,N_11421);
nor U12004 (N_12004,N_11411,N_11730);
and U12005 (N_12005,N_11391,N_11677);
nor U12006 (N_12006,N_11409,N_11281);
nor U12007 (N_12007,N_11832,N_11458);
and U12008 (N_12008,N_11577,N_11528);
nor U12009 (N_12009,N_11551,N_11718);
nand U12010 (N_12010,N_11265,N_11805);
or U12011 (N_12011,N_11840,N_11269);
or U12012 (N_12012,N_11405,N_11587);
xor U12013 (N_12013,N_11578,N_11693);
or U12014 (N_12014,N_11784,N_11669);
or U12015 (N_12015,N_11251,N_11774);
or U12016 (N_12016,N_11272,N_11472);
xnor U12017 (N_12017,N_11518,N_11415);
xor U12018 (N_12018,N_11359,N_11642);
nand U12019 (N_12019,N_11349,N_11701);
and U12020 (N_12020,N_11874,N_11548);
nor U12021 (N_12021,N_11745,N_11694);
or U12022 (N_12022,N_11767,N_11744);
xor U12023 (N_12023,N_11786,N_11270);
nor U12024 (N_12024,N_11307,N_11376);
nand U12025 (N_12025,N_11441,N_11549);
or U12026 (N_12026,N_11517,N_11584);
and U12027 (N_12027,N_11364,N_11545);
or U12028 (N_12028,N_11687,N_11643);
or U12029 (N_12029,N_11434,N_11583);
nor U12030 (N_12030,N_11818,N_11477);
and U12031 (N_12031,N_11685,N_11672);
xnor U12032 (N_12032,N_11760,N_11277);
nor U12033 (N_12033,N_11334,N_11430);
and U12034 (N_12034,N_11776,N_11484);
nand U12035 (N_12035,N_11800,N_11618);
xor U12036 (N_12036,N_11503,N_11442);
nor U12037 (N_12037,N_11279,N_11740);
xor U12038 (N_12038,N_11747,N_11839);
or U12039 (N_12039,N_11849,N_11614);
nor U12040 (N_12040,N_11781,N_11523);
nand U12041 (N_12041,N_11362,N_11835);
xor U12042 (N_12042,N_11761,N_11470);
nor U12043 (N_12043,N_11326,N_11731);
or U12044 (N_12044,N_11448,N_11857);
xnor U12045 (N_12045,N_11684,N_11741);
and U12046 (N_12046,N_11390,N_11460);
and U12047 (N_12047,N_11868,N_11495);
xor U12048 (N_12048,N_11424,N_11645);
and U12049 (N_12049,N_11357,N_11828);
nand U12050 (N_12050,N_11810,N_11823);
or U12051 (N_12051,N_11320,N_11291);
nand U12052 (N_12052,N_11637,N_11520);
nand U12053 (N_12053,N_11855,N_11721);
nor U12054 (N_12054,N_11668,N_11256);
nand U12055 (N_12055,N_11707,N_11647);
xor U12056 (N_12056,N_11535,N_11396);
or U12057 (N_12057,N_11612,N_11550);
nor U12058 (N_12058,N_11821,N_11816);
nor U12059 (N_12059,N_11445,N_11371);
nand U12060 (N_12060,N_11733,N_11814);
nor U12061 (N_12061,N_11483,N_11631);
and U12062 (N_12062,N_11738,N_11780);
nand U12063 (N_12063,N_11253,N_11753);
or U12064 (N_12064,N_11335,N_11869);
xnor U12065 (N_12065,N_11379,N_11825);
and U12066 (N_12066,N_11683,N_11806);
and U12067 (N_12067,N_11378,N_11327);
nor U12068 (N_12068,N_11408,N_11383);
and U12069 (N_12069,N_11586,N_11459);
or U12070 (N_12070,N_11317,N_11511);
or U12071 (N_12071,N_11416,N_11316);
or U12072 (N_12072,N_11446,N_11452);
nand U12073 (N_12073,N_11842,N_11703);
and U12074 (N_12074,N_11682,N_11333);
xor U12075 (N_12075,N_11505,N_11527);
or U12076 (N_12076,N_11297,N_11866);
xnor U12077 (N_12077,N_11728,N_11616);
nand U12078 (N_12078,N_11657,N_11400);
nand U12079 (N_12079,N_11533,N_11676);
and U12080 (N_12080,N_11346,N_11686);
xor U12081 (N_12081,N_11266,N_11257);
xor U12082 (N_12082,N_11305,N_11355);
nand U12083 (N_12083,N_11432,N_11361);
nor U12084 (N_12084,N_11623,N_11496);
and U12085 (N_12085,N_11592,N_11713);
nor U12086 (N_12086,N_11395,N_11313);
and U12087 (N_12087,N_11309,N_11798);
or U12088 (N_12088,N_11382,N_11595);
nor U12089 (N_12089,N_11590,N_11743);
and U12090 (N_12090,N_11295,N_11491);
xnor U12091 (N_12091,N_11789,N_11524);
nor U12092 (N_12092,N_11510,N_11699);
nor U12093 (N_12093,N_11599,N_11648);
and U12094 (N_12094,N_11363,N_11619);
nand U12095 (N_12095,N_11844,N_11356);
and U12096 (N_12096,N_11809,N_11304);
or U12097 (N_12097,N_11712,N_11303);
nand U12098 (N_12098,N_11831,N_11418);
nand U12099 (N_12099,N_11385,N_11754);
xnor U12100 (N_12100,N_11836,N_11625);
nor U12101 (N_12101,N_11419,N_11258);
xor U12102 (N_12102,N_11451,N_11853);
nand U12103 (N_12103,N_11567,N_11287);
nand U12104 (N_12104,N_11278,N_11311);
or U12105 (N_12105,N_11611,N_11575);
xor U12106 (N_12106,N_11350,N_11827);
nor U12107 (N_12107,N_11652,N_11598);
xor U12108 (N_12108,N_11689,N_11393);
or U12109 (N_12109,N_11286,N_11493);
nand U12110 (N_12110,N_11404,N_11515);
nand U12111 (N_12111,N_11861,N_11829);
nor U12112 (N_12112,N_11589,N_11332);
or U12113 (N_12113,N_11593,N_11720);
and U12114 (N_12114,N_11617,N_11714);
and U12115 (N_12115,N_11656,N_11471);
or U12116 (N_12116,N_11847,N_11431);
nand U12117 (N_12117,N_11360,N_11414);
xor U12118 (N_12118,N_11771,N_11268);
xor U12119 (N_12119,N_11759,N_11679);
or U12120 (N_12120,N_11260,N_11772);
nor U12121 (N_12121,N_11666,N_11282);
xnor U12122 (N_12122,N_11465,N_11389);
and U12123 (N_12123,N_11667,N_11285);
and U12124 (N_12124,N_11500,N_11755);
nor U12125 (N_12125,N_11769,N_11462);
nor U12126 (N_12126,N_11624,N_11321);
xor U12127 (N_12127,N_11579,N_11498);
and U12128 (N_12128,N_11792,N_11530);
xor U12129 (N_12129,N_11793,N_11850);
and U12130 (N_12130,N_11499,N_11749);
nor U12131 (N_12131,N_11392,N_11417);
nand U12132 (N_12132,N_11766,N_11502);
nor U12133 (N_12133,N_11651,N_11706);
nand U12134 (N_12134,N_11271,N_11568);
xnor U12135 (N_12135,N_11752,N_11873);
nand U12136 (N_12136,N_11634,N_11348);
and U12137 (N_12137,N_11374,N_11715);
or U12138 (N_12138,N_11555,N_11384);
nand U12139 (N_12139,N_11646,N_11783);
and U12140 (N_12140,N_11807,N_11340);
nor U12141 (N_12141,N_11734,N_11824);
or U12142 (N_12142,N_11830,N_11312);
nor U12143 (N_12143,N_11261,N_11264);
nand U12144 (N_12144,N_11758,N_11600);
xnor U12145 (N_12145,N_11724,N_11255);
or U12146 (N_12146,N_11372,N_11854);
or U12147 (N_12147,N_11607,N_11709);
and U12148 (N_12148,N_11654,N_11591);
or U12149 (N_12149,N_11368,N_11347);
and U12150 (N_12150,N_11594,N_11662);
nor U12151 (N_12151,N_11653,N_11602);
nand U12152 (N_12152,N_11406,N_11324);
and U12153 (N_12153,N_11308,N_11455);
nor U12154 (N_12154,N_11655,N_11605);
nand U12155 (N_12155,N_11466,N_11447);
xor U12156 (N_12156,N_11751,N_11641);
xnor U12157 (N_12157,N_11531,N_11365);
or U12158 (N_12158,N_11603,N_11377);
nand U12159 (N_12159,N_11757,N_11871);
nand U12160 (N_12160,N_11778,N_11296);
and U12161 (N_12161,N_11680,N_11768);
and U12162 (N_12162,N_11658,N_11341);
nand U12163 (N_12163,N_11581,N_11722);
nor U12164 (N_12164,N_11299,N_11727);
nor U12165 (N_12165,N_11343,N_11716);
and U12166 (N_12166,N_11691,N_11318);
or U12167 (N_12167,N_11536,N_11387);
or U12168 (N_12168,N_11702,N_11610);
and U12169 (N_12169,N_11506,N_11791);
xor U12170 (N_12170,N_11863,N_11756);
and U12171 (N_12171,N_11700,N_11852);
nand U12172 (N_12172,N_11559,N_11509);
and U12173 (N_12173,N_11403,N_11290);
xnor U12174 (N_12174,N_11867,N_11604);
or U12175 (N_12175,N_11353,N_11601);
nand U12176 (N_12176,N_11464,N_11437);
xor U12177 (N_12177,N_11439,N_11412);
xnor U12178 (N_12178,N_11398,N_11582);
and U12179 (N_12179,N_11342,N_11794);
and U12180 (N_12180,N_11697,N_11514);
nand U12181 (N_12181,N_11525,N_11526);
xnor U12182 (N_12182,N_11544,N_11280);
and U12183 (N_12183,N_11573,N_11319);
or U12184 (N_12184,N_11454,N_11410);
and U12185 (N_12185,N_11833,N_11539);
and U12186 (N_12186,N_11650,N_11870);
and U12187 (N_12187,N_11429,N_11850);
nand U12188 (N_12188,N_11779,N_11377);
nor U12189 (N_12189,N_11742,N_11734);
nand U12190 (N_12190,N_11870,N_11614);
nor U12191 (N_12191,N_11489,N_11797);
or U12192 (N_12192,N_11458,N_11860);
xnor U12193 (N_12193,N_11540,N_11395);
nor U12194 (N_12194,N_11736,N_11409);
xor U12195 (N_12195,N_11715,N_11486);
or U12196 (N_12196,N_11849,N_11610);
nand U12197 (N_12197,N_11752,N_11321);
nand U12198 (N_12198,N_11421,N_11558);
and U12199 (N_12199,N_11862,N_11530);
or U12200 (N_12200,N_11593,N_11677);
nand U12201 (N_12201,N_11324,N_11812);
nand U12202 (N_12202,N_11489,N_11697);
xnor U12203 (N_12203,N_11404,N_11366);
nor U12204 (N_12204,N_11284,N_11329);
xnor U12205 (N_12205,N_11717,N_11585);
nand U12206 (N_12206,N_11688,N_11610);
or U12207 (N_12207,N_11419,N_11310);
xor U12208 (N_12208,N_11824,N_11869);
nor U12209 (N_12209,N_11556,N_11619);
xnor U12210 (N_12210,N_11686,N_11754);
nand U12211 (N_12211,N_11274,N_11332);
xnor U12212 (N_12212,N_11666,N_11706);
and U12213 (N_12213,N_11525,N_11252);
and U12214 (N_12214,N_11781,N_11672);
and U12215 (N_12215,N_11623,N_11329);
and U12216 (N_12216,N_11606,N_11597);
nand U12217 (N_12217,N_11826,N_11611);
and U12218 (N_12218,N_11521,N_11430);
nor U12219 (N_12219,N_11589,N_11378);
nand U12220 (N_12220,N_11665,N_11259);
xnor U12221 (N_12221,N_11311,N_11815);
and U12222 (N_12222,N_11818,N_11589);
xor U12223 (N_12223,N_11470,N_11326);
nor U12224 (N_12224,N_11668,N_11396);
or U12225 (N_12225,N_11835,N_11836);
nand U12226 (N_12226,N_11645,N_11439);
nor U12227 (N_12227,N_11304,N_11406);
and U12228 (N_12228,N_11502,N_11629);
nor U12229 (N_12229,N_11572,N_11677);
xnor U12230 (N_12230,N_11742,N_11453);
xor U12231 (N_12231,N_11487,N_11759);
xnor U12232 (N_12232,N_11402,N_11694);
nor U12233 (N_12233,N_11722,N_11486);
nor U12234 (N_12234,N_11380,N_11366);
xnor U12235 (N_12235,N_11627,N_11528);
or U12236 (N_12236,N_11295,N_11487);
nand U12237 (N_12237,N_11293,N_11528);
nand U12238 (N_12238,N_11801,N_11787);
nor U12239 (N_12239,N_11743,N_11546);
nand U12240 (N_12240,N_11268,N_11574);
xor U12241 (N_12241,N_11841,N_11761);
nor U12242 (N_12242,N_11405,N_11484);
and U12243 (N_12243,N_11776,N_11583);
xnor U12244 (N_12244,N_11638,N_11849);
and U12245 (N_12245,N_11795,N_11666);
nand U12246 (N_12246,N_11283,N_11310);
or U12247 (N_12247,N_11372,N_11406);
nand U12248 (N_12248,N_11714,N_11350);
nand U12249 (N_12249,N_11491,N_11644);
nand U12250 (N_12250,N_11341,N_11315);
or U12251 (N_12251,N_11522,N_11331);
or U12252 (N_12252,N_11430,N_11658);
or U12253 (N_12253,N_11480,N_11666);
or U12254 (N_12254,N_11324,N_11703);
and U12255 (N_12255,N_11447,N_11837);
nand U12256 (N_12256,N_11809,N_11390);
nand U12257 (N_12257,N_11677,N_11514);
and U12258 (N_12258,N_11684,N_11481);
nor U12259 (N_12259,N_11859,N_11487);
or U12260 (N_12260,N_11770,N_11623);
nand U12261 (N_12261,N_11407,N_11721);
nand U12262 (N_12262,N_11643,N_11638);
and U12263 (N_12263,N_11457,N_11845);
xor U12264 (N_12264,N_11593,N_11459);
and U12265 (N_12265,N_11411,N_11613);
nor U12266 (N_12266,N_11474,N_11314);
or U12267 (N_12267,N_11787,N_11487);
nor U12268 (N_12268,N_11580,N_11519);
and U12269 (N_12269,N_11375,N_11852);
or U12270 (N_12270,N_11874,N_11343);
nor U12271 (N_12271,N_11512,N_11846);
or U12272 (N_12272,N_11321,N_11381);
xnor U12273 (N_12273,N_11807,N_11800);
nand U12274 (N_12274,N_11431,N_11349);
and U12275 (N_12275,N_11617,N_11749);
nor U12276 (N_12276,N_11548,N_11860);
xor U12277 (N_12277,N_11652,N_11605);
and U12278 (N_12278,N_11434,N_11771);
and U12279 (N_12279,N_11369,N_11377);
nand U12280 (N_12280,N_11825,N_11404);
nor U12281 (N_12281,N_11482,N_11812);
nand U12282 (N_12282,N_11617,N_11785);
nor U12283 (N_12283,N_11387,N_11825);
nor U12284 (N_12284,N_11447,N_11792);
and U12285 (N_12285,N_11705,N_11340);
xor U12286 (N_12286,N_11266,N_11457);
xnor U12287 (N_12287,N_11755,N_11389);
or U12288 (N_12288,N_11715,N_11797);
and U12289 (N_12289,N_11500,N_11518);
or U12290 (N_12290,N_11504,N_11474);
nor U12291 (N_12291,N_11685,N_11475);
or U12292 (N_12292,N_11658,N_11277);
or U12293 (N_12293,N_11665,N_11296);
and U12294 (N_12294,N_11423,N_11291);
nand U12295 (N_12295,N_11634,N_11668);
and U12296 (N_12296,N_11750,N_11480);
nor U12297 (N_12297,N_11524,N_11777);
xnor U12298 (N_12298,N_11262,N_11567);
nor U12299 (N_12299,N_11851,N_11525);
or U12300 (N_12300,N_11386,N_11335);
and U12301 (N_12301,N_11302,N_11763);
nor U12302 (N_12302,N_11743,N_11628);
nor U12303 (N_12303,N_11855,N_11442);
nor U12304 (N_12304,N_11565,N_11444);
or U12305 (N_12305,N_11303,N_11589);
and U12306 (N_12306,N_11342,N_11617);
nor U12307 (N_12307,N_11833,N_11757);
or U12308 (N_12308,N_11730,N_11573);
and U12309 (N_12309,N_11866,N_11659);
nor U12310 (N_12310,N_11312,N_11448);
xor U12311 (N_12311,N_11383,N_11701);
nor U12312 (N_12312,N_11755,N_11646);
and U12313 (N_12313,N_11324,N_11871);
nor U12314 (N_12314,N_11350,N_11708);
and U12315 (N_12315,N_11684,N_11263);
or U12316 (N_12316,N_11561,N_11635);
nor U12317 (N_12317,N_11430,N_11827);
nor U12318 (N_12318,N_11649,N_11501);
and U12319 (N_12319,N_11727,N_11328);
or U12320 (N_12320,N_11764,N_11835);
or U12321 (N_12321,N_11677,N_11471);
xor U12322 (N_12322,N_11322,N_11330);
nand U12323 (N_12323,N_11561,N_11460);
or U12324 (N_12324,N_11273,N_11526);
and U12325 (N_12325,N_11816,N_11831);
or U12326 (N_12326,N_11275,N_11774);
and U12327 (N_12327,N_11360,N_11511);
xor U12328 (N_12328,N_11261,N_11471);
xor U12329 (N_12329,N_11364,N_11614);
nand U12330 (N_12330,N_11684,N_11566);
and U12331 (N_12331,N_11823,N_11673);
xnor U12332 (N_12332,N_11282,N_11575);
or U12333 (N_12333,N_11580,N_11490);
nand U12334 (N_12334,N_11358,N_11510);
nor U12335 (N_12335,N_11511,N_11272);
nand U12336 (N_12336,N_11774,N_11343);
or U12337 (N_12337,N_11573,N_11724);
nand U12338 (N_12338,N_11415,N_11709);
xnor U12339 (N_12339,N_11400,N_11691);
xor U12340 (N_12340,N_11864,N_11856);
and U12341 (N_12341,N_11314,N_11452);
nand U12342 (N_12342,N_11261,N_11306);
xnor U12343 (N_12343,N_11370,N_11520);
and U12344 (N_12344,N_11360,N_11472);
nor U12345 (N_12345,N_11612,N_11469);
and U12346 (N_12346,N_11386,N_11659);
nor U12347 (N_12347,N_11265,N_11344);
and U12348 (N_12348,N_11541,N_11503);
nand U12349 (N_12349,N_11355,N_11424);
or U12350 (N_12350,N_11598,N_11290);
xor U12351 (N_12351,N_11741,N_11347);
nor U12352 (N_12352,N_11457,N_11313);
xnor U12353 (N_12353,N_11760,N_11322);
nand U12354 (N_12354,N_11317,N_11773);
nor U12355 (N_12355,N_11437,N_11279);
nand U12356 (N_12356,N_11273,N_11590);
or U12357 (N_12357,N_11467,N_11377);
and U12358 (N_12358,N_11798,N_11772);
nor U12359 (N_12359,N_11833,N_11711);
nand U12360 (N_12360,N_11514,N_11434);
nor U12361 (N_12361,N_11700,N_11452);
and U12362 (N_12362,N_11511,N_11429);
nand U12363 (N_12363,N_11392,N_11696);
and U12364 (N_12364,N_11827,N_11250);
and U12365 (N_12365,N_11309,N_11826);
or U12366 (N_12366,N_11507,N_11762);
or U12367 (N_12367,N_11486,N_11558);
or U12368 (N_12368,N_11487,N_11268);
nand U12369 (N_12369,N_11568,N_11474);
nand U12370 (N_12370,N_11406,N_11288);
and U12371 (N_12371,N_11749,N_11299);
nand U12372 (N_12372,N_11339,N_11817);
nor U12373 (N_12373,N_11436,N_11805);
xnor U12374 (N_12374,N_11609,N_11470);
nor U12375 (N_12375,N_11745,N_11575);
nand U12376 (N_12376,N_11521,N_11365);
and U12377 (N_12377,N_11517,N_11659);
nand U12378 (N_12378,N_11740,N_11581);
and U12379 (N_12379,N_11452,N_11668);
nor U12380 (N_12380,N_11287,N_11870);
or U12381 (N_12381,N_11738,N_11284);
xnor U12382 (N_12382,N_11870,N_11491);
xnor U12383 (N_12383,N_11661,N_11276);
or U12384 (N_12384,N_11288,N_11833);
nand U12385 (N_12385,N_11348,N_11813);
nor U12386 (N_12386,N_11376,N_11302);
and U12387 (N_12387,N_11683,N_11314);
nor U12388 (N_12388,N_11271,N_11384);
and U12389 (N_12389,N_11282,N_11777);
and U12390 (N_12390,N_11475,N_11612);
and U12391 (N_12391,N_11656,N_11668);
or U12392 (N_12392,N_11279,N_11254);
xnor U12393 (N_12393,N_11533,N_11466);
nor U12394 (N_12394,N_11475,N_11550);
xnor U12395 (N_12395,N_11568,N_11865);
or U12396 (N_12396,N_11473,N_11601);
and U12397 (N_12397,N_11265,N_11500);
nand U12398 (N_12398,N_11436,N_11526);
nand U12399 (N_12399,N_11583,N_11452);
or U12400 (N_12400,N_11640,N_11676);
nor U12401 (N_12401,N_11300,N_11290);
nand U12402 (N_12402,N_11618,N_11357);
xor U12403 (N_12403,N_11760,N_11337);
or U12404 (N_12404,N_11622,N_11648);
and U12405 (N_12405,N_11774,N_11798);
nor U12406 (N_12406,N_11290,N_11369);
nor U12407 (N_12407,N_11614,N_11505);
and U12408 (N_12408,N_11722,N_11617);
nor U12409 (N_12409,N_11431,N_11725);
or U12410 (N_12410,N_11603,N_11685);
and U12411 (N_12411,N_11422,N_11850);
or U12412 (N_12412,N_11262,N_11758);
nor U12413 (N_12413,N_11469,N_11566);
nor U12414 (N_12414,N_11461,N_11557);
and U12415 (N_12415,N_11660,N_11760);
nand U12416 (N_12416,N_11809,N_11750);
nand U12417 (N_12417,N_11735,N_11826);
or U12418 (N_12418,N_11351,N_11445);
xnor U12419 (N_12419,N_11427,N_11326);
xor U12420 (N_12420,N_11571,N_11300);
xor U12421 (N_12421,N_11553,N_11812);
nor U12422 (N_12422,N_11330,N_11847);
xor U12423 (N_12423,N_11400,N_11591);
and U12424 (N_12424,N_11590,N_11592);
or U12425 (N_12425,N_11385,N_11677);
nor U12426 (N_12426,N_11301,N_11587);
and U12427 (N_12427,N_11273,N_11317);
nor U12428 (N_12428,N_11655,N_11289);
or U12429 (N_12429,N_11453,N_11483);
and U12430 (N_12430,N_11519,N_11429);
xor U12431 (N_12431,N_11625,N_11743);
or U12432 (N_12432,N_11588,N_11483);
and U12433 (N_12433,N_11650,N_11732);
nand U12434 (N_12434,N_11843,N_11477);
nor U12435 (N_12435,N_11722,N_11821);
xor U12436 (N_12436,N_11649,N_11465);
or U12437 (N_12437,N_11718,N_11330);
nor U12438 (N_12438,N_11597,N_11356);
xor U12439 (N_12439,N_11259,N_11326);
and U12440 (N_12440,N_11251,N_11852);
and U12441 (N_12441,N_11488,N_11390);
xor U12442 (N_12442,N_11443,N_11253);
and U12443 (N_12443,N_11624,N_11812);
or U12444 (N_12444,N_11505,N_11477);
nor U12445 (N_12445,N_11499,N_11449);
or U12446 (N_12446,N_11446,N_11349);
nor U12447 (N_12447,N_11281,N_11312);
nand U12448 (N_12448,N_11648,N_11299);
and U12449 (N_12449,N_11677,N_11594);
nor U12450 (N_12450,N_11593,N_11324);
nor U12451 (N_12451,N_11861,N_11567);
or U12452 (N_12452,N_11444,N_11691);
or U12453 (N_12453,N_11788,N_11333);
nand U12454 (N_12454,N_11286,N_11704);
and U12455 (N_12455,N_11305,N_11458);
nor U12456 (N_12456,N_11814,N_11276);
and U12457 (N_12457,N_11557,N_11669);
xor U12458 (N_12458,N_11738,N_11304);
or U12459 (N_12459,N_11325,N_11670);
and U12460 (N_12460,N_11301,N_11300);
or U12461 (N_12461,N_11721,N_11481);
nor U12462 (N_12462,N_11682,N_11504);
xor U12463 (N_12463,N_11535,N_11858);
nand U12464 (N_12464,N_11456,N_11824);
and U12465 (N_12465,N_11848,N_11684);
nand U12466 (N_12466,N_11449,N_11852);
or U12467 (N_12467,N_11525,N_11667);
nor U12468 (N_12468,N_11817,N_11871);
or U12469 (N_12469,N_11415,N_11727);
xnor U12470 (N_12470,N_11395,N_11489);
xnor U12471 (N_12471,N_11842,N_11426);
or U12472 (N_12472,N_11780,N_11834);
xor U12473 (N_12473,N_11682,N_11456);
nand U12474 (N_12474,N_11447,N_11486);
nand U12475 (N_12475,N_11591,N_11252);
and U12476 (N_12476,N_11420,N_11778);
nor U12477 (N_12477,N_11710,N_11569);
nand U12478 (N_12478,N_11308,N_11289);
nand U12479 (N_12479,N_11320,N_11496);
and U12480 (N_12480,N_11497,N_11677);
and U12481 (N_12481,N_11266,N_11645);
xnor U12482 (N_12482,N_11574,N_11402);
nor U12483 (N_12483,N_11391,N_11695);
nor U12484 (N_12484,N_11800,N_11419);
nor U12485 (N_12485,N_11513,N_11461);
and U12486 (N_12486,N_11674,N_11833);
nand U12487 (N_12487,N_11575,N_11497);
xnor U12488 (N_12488,N_11759,N_11660);
nor U12489 (N_12489,N_11262,N_11423);
xnor U12490 (N_12490,N_11270,N_11864);
xnor U12491 (N_12491,N_11862,N_11735);
or U12492 (N_12492,N_11808,N_11434);
xnor U12493 (N_12493,N_11517,N_11464);
xnor U12494 (N_12494,N_11607,N_11829);
and U12495 (N_12495,N_11618,N_11529);
and U12496 (N_12496,N_11321,N_11829);
nor U12497 (N_12497,N_11661,N_11255);
nor U12498 (N_12498,N_11798,N_11691);
nor U12499 (N_12499,N_11332,N_11341);
and U12500 (N_12500,N_12226,N_12407);
xor U12501 (N_12501,N_12095,N_12420);
nor U12502 (N_12502,N_11994,N_12471);
nand U12503 (N_12503,N_12399,N_11881);
xnor U12504 (N_12504,N_12002,N_12227);
and U12505 (N_12505,N_11875,N_11905);
and U12506 (N_12506,N_12311,N_12495);
nand U12507 (N_12507,N_11930,N_12120);
nor U12508 (N_12508,N_12172,N_12127);
nand U12509 (N_12509,N_11947,N_12241);
nor U12510 (N_12510,N_12481,N_12388);
and U12511 (N_12511,N_12493,N_12331);
xnor U12512 (N_12512,N_12079,N_12479);
or U12513 (N_12513,N_12083,N_12422);
nor U12514 (N_12514,N_12237,N_11898);
nor U12515 (N_12515,N_11902,N_12474);
and U12516 (N_12516,N_11979,N_11988);
and U12517 (N_12517,N_12193,N_12393);
nand U12518 (N_12518,N_12443,N_12490);
nand U12519 (N_12519,N_11931,N_12194);
nor U12520 (N_12520,N_12261,N_12013);
and U12521 (N_12521,N_12044,N_11912);
nand U12522 (N_12522,N_12030,N_12449);
xor U12523 (N_12523,N_12370,N_12119);
and U12524 (N_12524,N_12289,N_12483);
nand U12525 (N_12525,N_11993,N_12484);
nand U12526 (N_12526,N_12208,N_12287);
xnor U12527 (N_12527,N_12378,N_11942);
nor U12528 (N_12528,N_12110,N_11906);
or U12529 (N_12529,N_12174,N_11998);
or U12530 (N_12530,N_12494,N_12253);
or U12531 (N_12531,N_12201,N_12229);
xor U12532 (N_12532,N_11933,N_12042);
or U12533 (N_12533,N_12296,N_12077);
nand U12534 (N_12534,N_11914,N_12233);
xnor U12535 (N_12535,N_12255,N_12472);
or U12536 (N_12536,N_11969,N_12459);
nor U12537 (N_12537,N_12272,N_12069);
nor U12538 (N_12538,N_12305,N_12409);
nor U12539 (N_12539,N_12448,N_12021);
xnor U12540 (N_12540,N_12497,N_11965);
or U12541 (N_12541,N_11903,N_12344);
or U12542 (N_12542,N_12076,N_12334);
nor U12543 (N_12543,N_11926,N_12346);
or U12544 (N_12544,N_12178,N_12453);
and U12545 (N_12545,N_11948,N_11911);
nor U12546 (N_12546,N_12267,N_12169);
and U12547 (N_12547,N_12209,N_12088);
nand U12548 (N_12548,N_12298,N_12437);
nor U12549 (N_12549,N_12338,N_12185);
nor U12550 (N_12550,N_12432,N_12245);
nand U12551 (N_12551,N_12089,N_12191);
and U12552 (N_12552,N_12262,N_11985);
nand U12553 (N_12553,N_11953,N_12386);
xnor U12554 (N_12554,N_12286,N_12124);
nor U12555 (N_12555,N_12220,N_12224);
or U12556 (N_12556,N_11888,N_12288);
nand U12557 (N_12557,N_12379,N_12102);
nand U12558 (N_12558,N_12499,N_12452);
and U12559 (N_12559,N_12055,N_11900);
xnor U12560 (N_12560,N_12339,N_12247);
and U12561 (N_12561,N_12009,N_12200);
xor U12562 (N_12562,N_12382,N_11952);
nand U12563 (N_12563,N_12248,N_12160);
and U12564 (N_12564,N_12246,N_12099);
or U12565 (N_12565,N_12072,N_12019);
or U12566 (N_12566,N_12010,N_12403);
and U12567 (N_12567,N_12163,N_12475);
nand U12568 (N_12568,N_12166,N_12284);
nor U12569 (N_12569,N_12151,N_11886);
or U12570 (N_12570,N_12353,N_12275);
nor U12571 (N_12571,N_12056,N_12413);
or U12572 (N_12572,N_12461,N_11890);
and U12573 (N_12573,N_12463,N_12274);
nor U12574 (N_12574,N_12416,N_12478);
xnor U12575 (N_12575,N_11929,N_12427);
nor U12576 (N_12576,N_12325,N_12111);
and U12577 (N_12577,N_11913,N_12024);
nand U12578 (N_12578,N_12423,N_12428);
or U12579 (N_12579,N_12450,N_12492);
and U12580 (N_12580,N_12097,N_12045);
nand U12581 (N_12581,N_12349,N_12431);
nand U12582 (N_12582,N_11996,N_11934);
xnor U12583 (N_12583,N_12332,N_12301);
and U12584 (N_12584,N_12041,N_11995);
nand U12585 (N_12585,N_12051,N_12276);
or U12586 (N_12586,N_12371,N_12036);
and U12587 (N_12587,N_12468,N_12150);
or U12588 (N_12588,N_12299,N_11970);
xnor U12589 (N_12589,N_12436,N_12199);
nand U12590 (N_12590,N_12458,N_12059);
xnor U12591 (N_12591,N_12016,N_12447);
nor U12592 (N_12592,N_11918,N_12093);
xor U12593 (N_12593,N_12176,N_12328);
nor U12594 (N_12594,N_12103,N_12131);
or U12595 (N_12595,N_12361,N_11961);
nor U12596 (N_12596,N_12364,N_12130);
xnor U12597 (N_12597,N_11999,N_12114);
nand U12598 (N_12598,N_11946,N_12306);
xnor U12599 (N_12599,N_12367,N_11981);
nand U12600 (N_12600,N_12467,N_12425);
nor U12601 (N_12601,N_12020,N_12335);
or U12602 (N_12602,N_11925,N_11959);
nor U12603 (N_12603,N_12001,N_11889);
nor U12604 (N_12604,N_12268,N_12142);
or U12605 (N_12605,N_12312,N_12405);
xnor U12606 (N_12606,N_12122,N_12061);
xor U12607 (N_12607,N_12278,N_12085);
or U12608 (N_12608,N_12387,N_12108);
nor U12609 (N_12609,N_11878,N_12090);
and U12610 (N_12610,N_12218,N_12018);
xor U12611 (N_12611,N_11984,N_12139);
or U12612 (N_12612,N_12133,N_12330);
and U12613 (N_12613,N_12071,N_12215);
and U12614 (N_12614,N_12121,N_12424);
xor U12615 (N_12615,N_12357,N_12179);
and U12616 (N_12616,N_12377,N_12207);
and U12617 (N_12617,N_11887,N_11960);
nor U12618 (N_12618,N_12115,N_12234);
nor U12619 (N_12619,N_12113,N_11958);
and U12620 (N_12620,N_12197,N_12080);
and U12621 (N_12621,N_12029,N_12145);
and U12622 (N_12622,N_12400,N_12165);
xnor U12623 (N_12623,N_12318,N_11921);
xor U12624 (N_12624,N_11992,N_12337);
nand U12625 (N_12625,N_12270,N_12012);
or U12626 (N_12626,N_12292,N_12256);
nand U12627 (N_12627,N_11923,N_12170);
nor U12628 (N_12628,N_12317,N_12290);
nor U12629 (N_12629,N_11917,N_12252);
nand U12630 (N_12630,N_12466,N_12273);
nor U12631 (N_12631,N_12496,N_11955);
and U12632 (N_12632,N_11991,N_12281);
nand U12633 (N_12633,N_12392,N_11928);
or U12634 (N_12634,N_12035,N_12190);
nand U12635 (N_12635,N_12203,N_12106);
xor U12636 (N_12636,N_12054,N_12123);
xnor U12637 (N_12637,N_12236,N_12008);
or U12638 (N_12638,N_12310,N_12000);
or U12639 (N_12639,N_12372,N_12143);
nand U12640 (N_12640,N_11980,N_12362);
and U12641 (N_12641,N_12486,N_11972);
nor U12642 (N_12642,N_12212,N_11922);
xor U12643 (N_12643,N_12391,N_12359);
or U12644 (N_12644,N_12049,N_12319);
xnor U12645 (N_12645,N_12415,N_12410);
nor U12646 (N_12646,N_12417,N_12107);
or U12647 (N_12647,N_12438,N_12063);
nor U12648 (N_12648,N_11907,N_12104);
nand U12649 (N_12649,N_12219,N_11943);
xnor U12650 (N_12650,N_12140,N_12375);
and U12651 (N_12651,N_11879,N_12052);
xnor U12652 (N_12652,N_12026,N_11932);
xnor U12653 (N_12653,N_12148,N_12309);
nand U12654 (N_12654,N_12389,N_12263);
or U12655 (N_12655,N_12180,N_12320);
nor U12656 (N_12656,N_12395,N_12304);
nor U12657 (N_12657,N_12451,N_12129);
and U12658 (N_12658,N_11908,N_12360);
nand U12659 (N_12659,N_12098,N_12006);
nand U12660 (N_12660,N_12015,N_12153);
and U12661 (N_12661,N_12092,N_11904);
or U12662 (N_12662,N_12105,N_12348);
xor U12663 (N_12663,N_12068,N_11893);
nor U12664 (N_12664,N_12254,N_12297);
or U12665 (N_12665,N_11973,N_12047);
xnor U12666 (N_12666,N_12198,N_12487);
or U12667 (N_12667,N_12141,N_12161);
xor U12668 (N_12668,N_12135,N_12075);
nand U12669 (N_12669,N_12214,N_11920);
nand U12670 (N_12670,N_12155,N_12316);
xor U12671 (N_12671,N_12308,N_12152);
nand U12672 (N_12672,N_12136,N_12396);
nor U12673 (N_12673,N_12404,N_12390);
xor U12674 (N_12674,N_12154,N_12446);
nand U12675 (N_12675,N_12336,N_12457);
and U12676 (N_12676,N_12017,N_12003);
nand U12677 (N_12677,N_12005,N_12302);
or U12678 (N_12678,N_12096,N_12081);
xnor U12679 (N_12679,N_11990,N_12369);
or U12680 (N_12680,N_12007,N_12421);
and U12681 (N_12681,N_12144,N_11936);
or U12682 (N_12682,N_12473,N_12430);
nand U12683 (N_12683,N_12406,N_12048);
and U12684 (N_12684,N_11891,N_12498);
xnor U12685 (N_12685,N_12147,N_12239);
xor U12686 (N_12686,N_12265,N_11882);
or U12687 (N_12687,N_12283,N_12225);
nand U12688 (N_12688,N_12394,N_11895);
nand U12689 (N_12689,N_12381,N_11940);
and U12690 (N_12690,N_12482,N_11986);
and U12691 (N_12691,N_12285,N_12232);
xnor U12692 (N_12692,N_12192,N_12347);
nor U12693 (N_12693,N_12164,N_12350);
or U12694 (N_12694,N_12258,N_12277);
or U12695 (N_12695,N_11949,N_12175);
nand U12696 (N_12696,N_12053,N_12231);
or U12697 (N_12697,N_12322,N_12132);
and U12698 (N_12698,N_12238,N_12204);
and U12699 (N_12699,N_11899,N_12429);
and U12700 (N_12700,N_12294,N_12167);
xnor U12701 (N_12701,N_12279,N_12128);
and U12702 (N_12702,N_11944,N_12398);
xnor U12703 (N_12703,N_12159,N_11909);
or U12704 (N_12704,N_12078,N_12327);
nand U12705 (N_12705,N_12455,N_11916);
nor U12706 (N_12706,N_12380,N_12066);
nand U12707 (N_12707,N_11915,N_12383);
or U12708 (N_12708,N_12489,N_11924);
xor U12709 (N_12709,N_12038,N_12266);
or U12710 (N_12710,N_12374,N_12456);
xnor U12711 (N_12711,N_12343,N_12345);
and U12712 (N_12712,N_12402,N_11896);
or U12713 (N_12713,N_12210,N_12125);
nand U12714 (N_12714,N_12173,N_12189);
nor U12715 (N_12715,N_12470,N_12216);
nand U12716 (N_12716,N_12363,N_12014);
nand U12717 (N_12717,N_11966,N_12315);
nor U12718 (N_12718,N_12480,N_12100);
nor U12719 (N_12719,N_12454,N_11937);
nor U12720 (N_12720,N_12243,N_11971);
nor U12721 (N_12721,N_12464,N_12050);
xor U12722 (N_12722,N_12117,N_12356);
xnor U12723 (N_12723,N_11987,N_12333);
xnor U12724 (N_12724,N_12476,N_11919);
nand U12725 (N_12725,N_12329,N_12134);
nor U12726 (N_12726,N_12412,N_12181);
nor U12727 (N_12727,N_12168,N_12291);
nand U12728 (N_12728,N_12213,N_12462);
nand U12729 (N_12729,N_12228,N_12477);
nor U12730 (N_12730,N_12032,N_12419);
nand U12731 (N_12731,N_12314,N_12433);
xnor U12732 (N_12732,N_11963,N_12149);
nand U12733 (N_12733,N_11978,N_12058);
and U12734 (N_12734,N_12295,N_12184);
nand U12735 (N_12735,N_12023,N_12313);
nor U12736 (N_12736,N_12376,N_12101);
nor U12737 (N_12737,N_11885,N_12094);
xnor U12738 (N_12738,N_12082,N_12156);
nor U12739 (N_12739,N_12087,N_12465);
nand U12740 (N_12740,N_12358,N_12025);
nand U12741 (N_12741,N_12027,N_12303);
and U12742 (N_12742,N_12355,N_12046);
nand U12743 (N_12743,N_12414,N_12205);
nand U12744 (N_12744,N_11957,N_11939);
nand U12745 (N_12745,N_11983,N_11892);
xor U12746 (N_12746,N_12249,N_12022);
nand U12747 (N_12747,N_12488,N_11938);
or U12748 (N_12748,N_11884,N_12491);
or U12749 (N_12749,N_12091,N_12440);
nand U12750 (N_12750,N_11967,N_12351);
nor U12751 (N_12751,N_12158,N_12401);
and U12752 (N_12752,N_12342,N_12426);
nand U12753 (N_12753,N_12307,N_11877);
or U12754 (N_12754,N_12469,N_12043);
or U12755 (N_12755,N_12251,N_12341);
and U12756 (N_12756,N_12062,N_12031);
xor U12757 (N_12757,N_12385,N_12445);
xor U12758 (N_12758,N_12485,N_12188);
or U12759 (N_12759,N_11880,N_11901);
and U12760 (N_12760,N_12157,N_12171);
xor U12761 (N_12761,N_11897,N_12222);
and U12762 (N_12762,N_12195,N_12418);
and U12763 (N_12763,N_12460,N_12293);
xnor U12764 (N_12764,N_12354,N_12244);
nor U12765 (N_12765,N_11975,N_12271);
nor U12766 (N_12766,N_12242,N_11956);
and U12767 (N_12767,N_12259,N_12250);
xor U12768 (N_12768,N_12408,N_12074);
nand U12769 (N_12769,N_12441,N_12070);
nor U12770 (N_12770,N_12211,N_12444);
xor U12771 (N_12771,N_12177,N_12137);
and U12772 (N_12772,N_12257,N_12202);
and U12773 (N_12773,N_12057,N_11935);
or U12774 (N_12774,N_11894,N_12067);
nand U12775 (N_12775,N_11951,N_12182);
or U12776 (N_12776,N_12240,N_12206);
or U12777 (N_12777,N_12126,N_11964);
nor U12778 (N_12778,N_11982,N_12435);
xnor U12779 (N_12779,N_12028,N_12324);
or U12780 (N_12780,N_11974,N_12065);
xor U12781 (N_12781,N_11977,N_12260);
and U12782 (N_12782,N_11997,N_12384);
nor U12783 (N_12783,N_11910,N_12186);
nor U12784 (N_12784,N_12340,N_12365);
and U12785 (N_12785,N_12280,N_12146);
or U12786 (N_12786,N_12060,N_12040);
nor U12787 (N_12787,N_12033,N_11989);
xor U12788 (N_12788,N_12084,N_12282);
and U12789 (N_12789,N_11927,N_11954);
or U12790 (N_12790,N_12217,N_12323);
nand U12791 (N_12791,N_12411,N_11950);
nor U12792 (N_12792,N_11941,N_12439);
nor U12793 (N_12793,N_12230,N_11976);
nor U12794 (N_12794,N_12434,N_12162);
or U12795 (N_12795,N_12223,N_12235);
or U12796 (N_12796,N_12086,N_12269);
or U12797 (N_12797,N_12187,N_12442);
and U12798 (N_12798,N_12321,N_12366);
nor U12799 (N_12799,N_12368,N_12326);
or U12800 (N_12800,N_12264,N_11962);
nand U12801 (N_12801,N_12109,N_12034);
nand U12802 (N_12802,N_11968,N_11876);
nand U12803 (N_12803,N_12300,N_12112);
xnor U12804 (N_12804,N_12221,N_12073);
nand U12805 (N_12805,N_12118,N_12397);
and U12806 (N_12806,N_12373,N_12196);
nor U12807 (N_12807,N_11883,N_12064);
xnor U12808 (N_12808,N_12004,N_12183);
and U12809 (N_12809,N_12352,N_12116);
nand U12810 (N_12810,N_12039,N_12037);
xor U12811 (N_12811,N_12138,N_12011);
and U12812 (N_12812,N_11945,N_12008);
nor U12813 (N_12813,N_11938,N_12484);
xnor U12814 (N_12814,N_11996,N_12417);
and U12815 (N_12815,N_12247,N_12293);
xor U12816 (N_12816,N_11931,N_12423);
and U12817 (N_12817,N_12220,N_12379);
nor U12818 (N_12818,N_12003,N_12357);
nor U12819 (N_12819,N_12017,N_12230);
or U12820 (N_12820,N_12461,N_12383);
and U12821 (N_12821,N_12129,N_12191);
nand U12822 (N_12822,N_12367,N_12297);
nand U12823 (N_12823,N_12474,N_12002);
xnor U12824 (N_12824,N_12448,N_11983);
xnor U12825 (N_12825,N_12167,N_12010);
nand U12826 (N_12826,N_12287,N_12196);
and U12827 (N_12827,N_12017,N_11964);
and U12828 (N_12828,N_12109,N_12106);
and U12829 (N_12829,N_12286,N_12376);
or U12830 (N_12830,N_12069,N_12182);
nand U12831 (N_12831,N_12371,N_12313);
and U12832 (N_12832,N_12269,N_12125);
or U12833 (N_12833,N_12444,N_12219);
xnor U12834 (N_12834,N_12300,N_12252);
nor U12835 (N_12835,N_12240,N_12440);
nand U12836 (N_12836,N_12162,N_12126);
or U12837 (N_12837,N_11972,N_11988);
nor U12838 (N_12838,N_12326,N_12458);
and U12839 (N_12839,N_12276,N_11957);
nand U12840 (N_12840,N_12263,N_11905);
nand U12841 (N_12841,N_12329,N_11916);
xnor U12842 (N_12842,N_12101,N_12355);
nand U12843 (N_12843,N_12212,N_12434);
and U12844 (N_12844,N_11947,N_12489);
nand U12845 (N_12845,N_11899,N_12318);
xor U12846 (N_12846,N_11987,N_11940);
xnor U12847 (N_12847,N_12097,N_12167);
xor U12848 (N_12848,N_12267,N_12355);
and U12849 (N_12849,N_12294,N_12351);
nand U12850 (N_12850,N_12031,N_12166);
nor U12851 (N_12851,N_12304,N_11936);
xor U12852 (N_12852,N_12358,N_12332);
nor U12853 (N_12853,N_12351,N_11928);
xnor U12854 (N_12854,N_12435,N_12369);
or U12855 (N_12855,N_12179,N_12126);
or U12856 (N_12856,N_12170,N_12239);
or U12857 (N_12857,N_12245,N_12477);
and U12858 (N_12858,N_12466,N_11986);
nor U12859 (N_12859,N_12191,N_11975);
xnor U12860 (N_12860,N_12084,N_11919);
nand U12861 (N_12861,N_12404,N_12155);
nor U12862 (N_12862,N_12168,N_12104);
nor U12863 (N_12863,N_12196,N_11999);
and U12864 (N_12864,N_11975,N_12488);
and U12865 (N_12865,N_12365,N_12277);
nor U12866 (N_12866,N_12410,N_11912);
or U12867 (N_12867,N_12458,N_12309);
nand U12868 (N_12868,N_12174,N_12049);
or U12869 (N_12869,N_11964,N_12223);
nor U12870 (N_12870,N_12173,N_11914);
or U12871 (N_12871,N_12013,N_11989);
or U12872 (N_12872,N_12211,N_12493);
or U12873 (N_12873,N_12234,N_11966);
or U12874 (N_12874,N_11921,N_12343);
and U12875 (N_12875,N_12476,N_12347);
nand U12876 (N_12876,N_12240,N_12244);
xor U12877 (N_12877,N_12393,N_11944);
xnor U12878 (N_12878,N_12445,N_12047);
nand U12879 (N_12879,N_12345,N_12061);
nor U12880 (N_12880,N_12275,N_12197);
nand U12881 (N_12881,N_12284,N_12143);
xnor U12882 (N_12882,N_12205,N_12121);
nand U12883 (N_12883,N_12349,N_12423);
nand U12884 (N_12884,N_12147,N_12203);
or U12885 (N_12885,N_12428,N_11896);
xnor U12886 (N_12886,N_12369,N_11911);
and U12887 (N_12887,N_11996,N_12101);
nor U12888 (N_12888,N_12025,N_12405);
nor U12889 (N_12889,N_12296,N_11991);
or U12890 (N_12890,N_12322,N_11995);
nor U12891 (N_12891,N_12481,N_12246);
and U12892 (N_12892,N_12396,N_12182);
and U12893 (N_12893,N_12330,N_12132);
nand U12894 (N_12894,N_12072,N_12359);
xor U12895 (N_12895,N_12123,N_12184);
nor U12896 (N_12896,N_12377,N_12199);
nand U12897 (N_12897,N_12246,N_12130);
nand U12898 (N_12898,N_12263,N_11933);
or U12899 (N_12899,N_12488,N_12320);
nand U12900 (N_12900,N_12336,N_11925);
and U12901 (N_12901,N_11969,N_12232);
nand U12902 (N_12902,N_12494,N_12419);
xnor U12903 (N_12903,N_11906,N_12035);
xnor U12904 (N_12904,N_12357,N_12476);
xor U12905 (N_12905,N_12326,N_12142);
and U12906 (N_12906,N_12465,N_12216);
and U12907 (N_12907,N_12027,N_12464);
nor U12908 (N_12908,N_11938,N_12117);
xnor U12909 (N_12909,N_12277,N_11998);
or U12910 (N_12910,N_12237,N_12059);
nand U12911 (N_12911,N_12470,N_12455);
or U12912 (N_12912,N_12294,N_12121);
xnor U12913 (N_12913,N_12275,N_12248);
and U12914 (N_12914,N_12310,N_12198);
nor U12915 (N_12915,N_12254,N_12215);
xor U12916 (N_12916,N_12055,N_12421);
or U12917 (N_12917,N_11992,N_12276);
nor U12918 (N_12918,N_12166,N_12438);
xnor U12919 (N_12919,N_12222,N_12213);
nor U12920 (N_12920,N_12310,N_12012);
and U12921 (N_12921,N_12190,N_12223);
and U12922 (N_12922,N_12205,N_12213);
nor U12923 (N_12923,N_12280,N_12401);
xnor U12924 (N_12924,N_12454,N_12125);
or U12925 (N_12925,N_12343,N_12338);
nor U12926 (N_12926,N_11989,N_11900);
and U12927 (N_12927,N_12012,N_12466);
nor U12928 (N_12928,N_11969,N_12456);
nand U12929 (N_12929,N_12312,N_12065);
or U12930 (N_12930,N_11967,N_12189);
xnor U12931 (N_12931,N_11954,N_12147);
xnor U12932 (N_12932,N_12487,N_11888);
or U12933 (N_12933,N_12392,N_12444);
or U12934 (N_12934,N_12246,N_12406);
xnor U12935 (N_12935,N_12421,N_11897);
nand U12936 (N_12936,N_11961,N_12229);
and U12937 (N_12937,N_12180,N_12142);
and U12938 (N_12938,N_12482,N_11922);
and U12939 (N_12939,N_12140,N_12025);
or U12940 (N_12940,N_11903,N_12395);
xnor U12941 (N_12941,N_12013,N_12087);
xnor U12942 (N_12942,N_11981,N_12102);
xor U12943 (N_12943,N_12068,N_11902);
or U12944 (N_12944,N_12400,N_12134);
nand U12945 (N_12945,N_12466,N_12460);
xor U12946 (N_12946,N_11967,N_12408);
nand U12947 (N_12947,N_11904,N_11910);
xor U12948 (N_12948,N_12464,N_12400);
nor U12949 (N_12949,N_12059,N_12321);
and U12950 (N_12950,N_12166,N_11981);
nand U12951 (N_12951,N_12192,N_12362);
xnor U12952 (N_12952,N_12139,N_11952);
or U12953 (N_12953,N_11934,N_12156);
xnor U12954 (N_12954,N_12075,N_12335);
nor U12955 (N_12955,N_11909,N_12012);
or U12956 (N_12956,N_11992,N_12016);
and U12957 (N_12957,N_12358,N_11886);
nand U12958 (N_12958,N_12355,N_12071);
nor U12959 (N_12959,N_11914,N_12014);
or U12960 (N_12960,N_12363,N_12005);
nand U12961 (N_12961,N_11891,N_11898);
and U12962 (N_12962,N_12096,N_12389);
xnor U12963 (N_12963,N_11992,N_12372);
nor U12964 (N_12964,N_11912,N_12246);
nand U12965 (N_12965,N_12149,N_12165);
xor U12966 (N_12966,N_12364,N_11899);
or U12967 (N_12967,N_12389,N_12136);
and U12968 (N_12968,N_12419,N_12432);
and U12969 (N_12969,N_12369,N_11877);
xnor U12970 (N_12970,N_12060,N_12251);
or U12971 (N_12971,N_11920,N_11929);
or U12972 (N_12972,N_12311,N_12444);
or U12973 (N_12973,N_11969,N_12095);
and U12974 (N_12974,N_12192,N_11996);
xnor U12975 (N_12975,N_12464,N_12151);
and U12976 (N_12976,N_12414,N_12379);
or U12977 (N_12977,N_12051,N_12057);
nand U12978 (N_12978,N_11928,N_12144);
or U12979 (N_12979,N_11904,N_11900);
xor U12980 (N_12980,N_12175,N_12319);
and U12981 (N_12981,N_12484,N_12478);
nor U12982 (N_12982,N_12482,N_12379);
nand U12983 (N_12983,N_12110,N_11944);
nand U12984 (N_12984,N_12315,N_12040);
nand U12985 (N_12985,N_12279,N_12186);
nand U12986 (N_12986,N_11906,N_12250);
nand U12987 (N_12987,N_12281,N_12326);
nand U12988 (N_12988,N_12384,N_12118);
xor U12989 (N_12989,N_11922,N_12437);
and U12990 (N_12990,N_12004,N_12223);
nand U12991 (N_12991,N_12400,N_12053);
and U12992 (N_12992,N_12070,N_12002);
nand U12993 (N_12993,N_12412,N_12246);
and U12994 (N_12994,N_12323,N_12249);
or U12995 (N_12995,N_12223,N_11955);
nand U12996 (N_12996,N_12433,N_12311);
and U12997 (N_12997,N_11951,N_12339);
or U12998 (N_12998,N_12074,N_12091);
or U12999 (N_12999,N_12451,N_12326);
nand U13000 (N_13000,N_11884,N_12462);
xnor U13001 (N_13001,N_12239,N_12159);
xor U13002 (N_13002,N_12113,N_12261);
nor U13003 (N_13003,N_11996,N_12193);
nor U13004 (N_13004,N_12199,N_12319);
nor U13005 (N_13005,N_12213,N_12055);
nor U13006 (N_13006,N_12147,N_12218);
nand U13007 (N_13007,N_12377,N_12482);
nor U13008 (N_13008,N_12470,N_12243);
nand U13009 (N_13009,N_12238,N_12269);
and U13010 (N_13010,N_12282,N_11894);
and U13011 (N_13011,N_12124,N_12022);
nand U13012 (N_13012,N_12322,N_12137);
nand U13013 (N_13013,N_12495,N_12034);
or U13014 (N_13014,N_11992,N_12044);
nand U13015 (N_13015,N_12355,N_12386);
or U13016 (N_13016,N_12125,N_12401);
xor U13017 (N_13017,N_12248,N_11880);
or U13018 (N_13018,N_11927,N_12334);
nand U13019 (N_13019,N_12119,N_12395);
nor U13020 (N_13020,N_11987,N_12484);
nand U13021 (N_13021,N_12021,N_12435);
and U13022 (N_13022,N_12174,N_12327);
or U13023 (N_13023,N_11910,N_12488);
and U13024 (N_13024,N_11921,N_12268);
and U13025 (N_13025,N_11935,N_12000);
xor U13026 (N_13026,N_11991,N_11998);
or U13027 (N_13027,N_12042,N_12309);
nor U13028 (N_13028,N_12335,N_12333);
nand U13029 (N_13029,N_12086,N_12442);
xnor U13030 (N_13030,N_12286,N_11950);
and U13031 (N_13031,N_12333,N_12449);
nand U13032 (N_13032,N_12239,N_12336);
xnor U13033 (N_13033,N_12432,N_12467);
nor U13034 (N_13034,N_12003,N_11903);
nor U13035 (N_13035,N_12104,N_12032);
and U13036 (N_13036,N_11978,N_11902);
nand U13037 (N_13037,N_12158,N_12255);
nor U13038 (N_13038,N_12327,N_12266);
xnor U13039 (N_13039,N_11954,N_12267);
xnor U13040 (N_13040,N_12132,N_12402);
and U13041 (N_13041,N_12353,N_11904);
or U13042 (N_13042,N_12272,N_12139);
or U13043 (N_13043,N_12434,N_12177);
or U13044 (N_13044,N_11951,N_11912);
xor U13045 (N_13045,N_11923,N_12428);
and U13046 (N_13046,N_12056,N_11923);
or U13047 (N_13047,N_12276,N_12019);
nand U13048 (N_13048,N_12430,N_12278);
nand U13049 (N_13049,N_11914,N_11995);
nand U13050 (N_13050,N_11904,N_12151);
and U13051 (N_13051,N_12337,N_11909);
nor U13052 (N_13052,N_12254,N_12404);
nand U13053 (N_13053,N_12255,N_12004);
nor U13054 (N_13054,N_11893,N_11933);
or U13055 (N_13055,N_11907,N_12455);
and U13056 (N_13056,N_12129,N_12047);
xnor U13057 (N_13057,N_12310,N_12131);
and U13058 (N_13058,N_11933,N_12053);
or U13059 (N_13059,N_11949,N_12299);
nor U13060 (N_13060,N_12479,N_12395);
or U13061 (N_13061,N_12167,N_11970);
nor U13062 (N_13062,N_12398,N_12062);
or U13063 (N_13063,N_12087,N_12162);
or U13064 (N_13064,N_12082,N_11955);
or U13065 (N_13065,N_12218,N_12405);
nand U13066 (N_13066,N_12434,N_12089);
nor U13067 (N_13067,N_12100,N_11932);
xor U13068 (N_13068,N_12099,N_12160);
or U13069 (N_13069,N_12182,N_12188);
nor U13070 (N_13070,N_12446,N_12431);
or U13071 (N_13071,N_11983,N_12471);
or U13072 (N_13072,N_11923,N_12273);
xnor U13073 (N_13073,N_11898,N_12281);
nand U13074 (N_13074,N_11897,N_11888);
xor U13075 (N_13075,N_12340,N_12293);
xor U13076 (N_13076,N_12250,N_12105);
nor U13077 (N_13077,N_12255,N_12008);
and U13078 (N_13078,N_11987,N_12118);
nor U13079 (N_13079,N_12485,N_12497);
xnor U13080 (N_13080,N_12154,N_12441);
xor U13081 (N_13081,N_12130,N_12234);
or U13082 (N_13082,N_12439,N_11932);
and U13083 (N_13083,N_12008,N_12205);
nand U13084 (N_13084,N_12199,N_12000);
and U13085 (N_13085,N_12234,N_11914);
or U13086 (N_13086,N_11935,N_12201);
xor U13087 (N_13087,N_12266,N_12365);
and U13088 (N_13088,N_11922,N_11889);
or U13089 (N_13089,N_12329,N_12138);
nor U13090 (N_13090,N_11942,N_12283);
xor U13091 (N_13091,N_12118,N_11983);
and U13092 (N_13092,N_12187,N_12377);
nand U13093 (N_13093,N_12213,N_12291);
and U13094 (N_13094,N_12421,N_11983);
nor U13095 (N_13095,N_12233,N_12360);
or U13096 (N_13096,N_11975,N_11876);
nor U13097 (N_13097,N_12042,N_12040);
nor U13098 (N_13098,N_12367,N_12064);
and U13099 (N_13099,N_11897,N_12262);
nor U13100 (N_13100,N_12081,N_12451);
xnor U13101 (N_13101,N_12266,N_11902);
and U13102 (N_13102,N_11947,N_12041);
xor U13103 (N_13103,N_12136,N_12260);
nor U13104 (N_13104,N_12437,N_12292);
nand U13105 (N_13105,N_12115,N_11971);
nand U13106 (N_13106,N_12168,N_12399);
xnor U13107 (N_13107,N_12398,N_12138);
nor U13108 (N_13108,N_12059,N_12345);
xnor U13109 (N_13109,N_12289,N_12085);
nand U13110 (N_13110,N_12484,N_12352);
or U13111 (N_13111,N_12478,N_11976);
nor U13112 (N_13112,N_12395,N_12076);
nand U13113 (N_13113,N_12025,N_12076);
xnor U13114 (N_13114,N_12244,N_12262);
nand U13115 (N_13115,N_11915,N_12163);
or U13116 (N_13116,N_11875,N_12213);
or U13117 (N_13117,N_12415,N_11983);
xnor U13118 (N_13118,N_12256,N_12377);
or U13119 (N_13119,N_12082,N_11926);
nor U13120 (N_13120,N_12144,N_12355);
nand U13121 (N_13121,N_11939,N_12245);
nand U13122 (N_13122,N_12464,N_12036);
xnor U13123 (N_13123,N_12132,N_12323);
and U13124 (N_13124,N_11994,N_12249);
and U13125 (N_13125,N_12929,N_12648);
and U13126 (N_13126,N_12657,N_12667);
and U13127 (N_13127,N_12543,N_12551);
nor U13128 (N_13128,N_12621,N_12526);
nand U13129 (N_13129,N_13073,N_12663);
and U13130 (N_13130,N_12601,N_12606);
or U13131 (N_13131,N_12767,N_13053);
nor U13132 (N_13132,N_13015,N_12576);
and U13133 (N_13133,N_12567,N_12936);
or U13134 (N_13134,N_12997,N_12788);
nand U13135 (N_13135,N_12868,N_12783);
or U13136 (N_13136,N_12636,N_13001);
nor U13137 (N_13137,N_13122,N_12638);
nand U13138 (N_13138,N_13044,N_13049);
and U13139 (N_13139,N_12906,N_12653);
and U13140 (N_13140,N_12772,N_12646);
xor U13141 (N_13141,N_13036,N_12629);
nor U13142 (N_13142,N_12969,N_12747);
and U13143 (N_13143,N_13029,N_12943);
or U13144 (N_13144,N_12872,N_13118);
and U13145 (N_13145,N_12743,N_12907);
and U13146 (N_13146,N_12709,N_13115);
xnor U13147 (N_13147,N_12630,N_12544);
nand U13148 (N_13148,N_13061,N_12804);
nor U13149 (N_13149,N_12990,N_12961);
nor U13150 (N_13150,N_12723,N_12710);
or U13151 (N_13151,N_12904,N_12847);
nand U13152 (N_13152,N_12507,N_12729);
xor U13153 (N_13153,N_13060,N_12587);
and U13154 (N_13154,N_13086,N_12799);
or U13155 (N_13155,N_12958,N_12752);
or U13156 (N_13156,N_12637,N_12983);
nand U13157 (N_13157,N_12859,N_12966);
or U13158 (N_13158,N_13028,N_12921);
and U13159 (N_13159,N_12725,N_13108);
or U13160 (N_13160,N_12550,N_12707);
nand U13161 (N_13161,N_12968,N_12655);
and U13162 (N_13162,N_12843,N_12771);
nor U13163 (N_13163,N_12774,N_12835);
or U13164 (N_13164,N_13035,N_12738);
xnor U13165 (N_13165,N_12863,N_12501);
or U13166 (N_13166,N_12581,N_12886);
nor U13167 (N_13167,N_13100,N_13006);
nor U13168 (N_13168,N_13111,N_13027);
and U13169 (N_13169,N_13120,N_12631);
nand U13170 (N_13170,N_12977,N_12930);
nor U13171 (N_13171,N_13017,N_12684);
xnor U13172 (N_13172,N_12611,N_12866);
or U13173 (N_13173,N_12950,N_13024);
and U13174 (N_13174,N_12882,N_12677);
and U13175 (N_13175,N_12945,N_12937);
nand U13176 (N_13176,N_12589,N_12915);
and U13177 (N_13177,N_12726,N_12632);
and U13178 (N_13178,N_13033,N_12765);
nand U13179 (N_13179,N_12972,N_12787);
or U13180 (N_13180,N_12876,N_12586);
and U13181 (N_13181,N_13000,N_12650);
or U13182 (N_13182,N_12916,N_12923);
nand U13183 (N_13183,N_12640,N_12645);
xnor U13184 (N_13184,N_13034,N_12508);
nand U13185 (N_13185,N_12773,N_12794);
nor U13186 (N_13186,N_12815,N_12880);
nor U13187 (N_13187,N_12885,N_12696);
nor U13188 (N_13188,N_12582,N_12701);
nor U13189 (N_13189,N_12609,N_13025);
or U13190 (N_13190,N_12952,N_12524);
nand U13191 (N_13191,N_12678,N_12911);
xor U13192 (N_13192,N_12846,N_12635);
nand U13193 (N_13193,N_12825,N_13055);
and U13194 (N_13194,N_12509,N_13002);
nand U13195 (N_13195,N_12698,N_12792);
nor U13196 (N_13196,N_12973,N_12728);
nor U13197 (N_13197,N_12626,N_12702);
nor U13198 (N_13198,N_12778,N_12675);
and U13199 (N_13199,N_12775,N_12959);
nor U13200 (N_13200,N_13010,N_12529);
or U13201 (N_13201,N_12548,N_12522);
nor U13202 (N_13202,N_13080,N_12542);
and U13203 (N_13203,N_12855,N_12754);
or U13204 (N_13204,N_12727,N_12612);
xor U13205 (N_13205,N_12895,N_12992);
nor U13206 (N_13206,N_13063,N_12730);
nor U13207 (N_13207,N_13058,N_12713);
xnor U13208 (N_13208,N_12776,N_12742);
nor U13209 (N_13209,N_13030,N_12602);
or U13210 (N_13210,N_12789,N_12506);
or U13211 (N_13211,N_12527,N_12926);
xnor U13212 (N_13212,N_12664,N_12549);
nand U13213 (N_13213,N_13023,N_12830);
nand U13214 (N_13214,N_12692,N_12674);
nand U13215 (N_13215,N_12999,N_12759);
xor U13216 (N_13216,N_12570,N_13075);
nor U13217 (N_13217,N_12914,N_12623);
xnor U13218 (N_13218,N_12736,N_12547);
and U13219 (N_13219,N_13095,N_12735);
nor U13220 (N_13220,N_12853,N_13003);
or U13221 (N_13221,N_13094,N_12532);
xor U13222 (N_13222,N_12962,N_13087);
or U13223 (N_13223,N_12564,N_13059);
and U13224 (N_13224,N_12770,N_12536);
xor U13225 (N_13225,N_13011,N_12947);
nand U13226 (N_13226,N_12644,N_12817);
nand U13227 (N_13227,N_12541,N_12852);
and U13228 (N_13228,N_12714,N_13074);
or U13229 (N_13229,N_12732,N_12545);
xor U13230 (N_13230,N_12615,N_12856);
or U13231 (N_13231,N_12503,N_12669);
and U13232 (N_13232,N_12687,N_12965);
and U13233 (N_13233,N_13048,N_12516);
and U13234 (N_13234,N_12671,N_13052);
or U13235 (N_13235,N_12731,N_12748);
nand U13236 (N_13236,N_12812,N_12610);
or U13237 (N_13237,N_12777,N_12976);
nand U13238 (N_13238,N_12598,N_13121);
or U13239 (N_13239,N_12889,N_13103);
xor U13240 (N_13240,N_12837,N_12809);
or U13241 (N_13241,N_13046,N_12652);
nor U13242 (N_13242,N_12898,N_12569);
nand U13243 (N_13243,N_12672,N_13051);
nand U13244 (N_13244,N_12896,N_12989);
nand U13245 (N_13245,N_12873,N_12520);
and U13246 (N_13246,N_12697,N_12944);
or U13247 (N_13247,N_12917,N_12500);
nand U13248 (N_13248,N_13038,N_13039);
nand U13249 (N_13249,N_13081,N_13040);
nand U13250 (N_13250,N_12991,N_12539);
nand U13251 (N_13251,N_12528,N_12801);
nor U13252 (N_13252,N_12993,N_13005);
and U13253 (N_13253,N_12596,N_12718);
nor U13254 (N_13254,N_13070,N_13014);
and U13255 (N_13255,N_12922,N_12806);
nor U13256 (N_13256,N_12768,N_12888);
nand U13257 (N_13257,N_12786,N_12733);
xnor U13258 (N_13258,N_13007,N_12593);
or U13259 (N_13259,N_12502,N_12592);
nand U13260 (N_13260,N_13101,N_12643);
nor U13261 (N_13261,N_12975,N_12927);
nor U13262 (N_13262,N_12721,N_13114);
xor U13263 (N_13263,N_13096,N_12967);
nand U13264 (N_13264,N_12935,N_12763);
and U13265 (N_13265,N_12960,N_12744);
and U13266 (N_13266,N_13124,N_12505);
and U13267 (N_13267,N_12795,N_12802);
or U13268 (N_13268,N_13112,N_13056);
or U13269 (N_13269,N_13031,N_13082);
nor U13270 (N_13270,N_12893,N_12715);
nor U13271 (N_13271,N_12562,N_12558);
or U13272 (N_13272,N_12790,N_12757);
nand U13273 (N_13273,N_12963,N_13119);
nand U13274 (N_13274,N_12620,N_12689);
nor U13275 (N_13275,N_12591,N_13105);
and U13276 (N_13276,N_13097,N_12634);
xnor U13277 (N_13277,N_12942,N_12600);
or U13278 (N_13278,N_12628,N_12749);
xor U13279 (N_13279,N_12980,N_12836);
xnor U13280 (N_13280,N_13042,N_13085);
nor U13281 (N_13281,N_12690,N_12642);
nand U13282 (N_13282,N_12884,N_13072);
nand U13283 (N_13283,N_13062,N_12537);
nor U13284 (N_13284,N_13107,N_12941);
nand U13285 (N_13285,N_13068,N_12782);
xor U13286 (N_13286,N_12662,N_12595);
xor U13287 (N_13287,N_12946,N_12588);
nand U13288 (N_13288,N_12820,N_12580);
and U13289 (N_13289,N_12761,N_12666);
or U13290 (N_13290,N_12685,N_12828);
and U13291 (N_13291,N_12627,N_12982);
nand U13292 (N_13292,N_12762,N_12574);
nor U13293 (N_13293,N_12780,N_12622);
nor U13294 (N_13294,N_12784,N_12909);
nor U13295 (N_13295,N_12877,N_12779);
nor U13296 (N_13296,N_12954,N_12850);
or U13297 (N_13297,N_12750,N_12682);
nand U13298 (N_13298,N_12938,N_12870);
xor U13299 (N_13299,N_12513,N_12970);
xor U13300 (N_13300,N_12823,N_13021);
or U13301 (N_13301,N_12619,N_12745);
nor U13302 (N_13302,N_12875,N_13009);
and U13303 (N_13303,N_12561,N_12679);
nand U13304 (N_13304,N_12785,N_12974);
nand U13305 (N_13305,N_12614,N_12791);
or U13306 (N_13306,N_13045,N_12881);
xor U13307 (N_13307,N_12816,N_12845);
nand U13308 (N_13308,N_12673,N_12840);
xnor U13309 (N_13309,N_12818,N_13091);
or U13310 (N_13310,N_12981,N_12932);
nor U13311 (N_13311,N_12831,N_12764);
nor U13312 (N_13312,N_12741,N_12552);
xor U13313 (N_13313,N_12533,N_12985);
xor U13314 (N_13314,N_12813,N_12824);
and U13315 (N_13315,N_12902,N_12579);
or U13316 (N_13316,N_13093,N_12555);
xnor U13317 (N_13317,N_12560,N_13104);
nor U13318 (N_13318,N_12940,N_12808);
xnor U13319 (N_13319,N_12572,N_12583);
and U13320 (N_13320,N_12905,N_13019);
nand U13321 (N_13321,N_12769,N_12857);
and U13322 (N_13322,N_12519,N_12793);
nand U13323 (N_13323,N_12703,N_12565);
nand U13324 (N_13324,N_12607,N_12858);
xnor U13325 (N_13325,N_12874,N_12633);
or U13326 (N_13326,N_12971,N_12854);
or U13327 (N_13327,N_12668,N_12918);
xor U13328 (N_13328,N_12624,N_12525);
or U13329 (N_13329,N_13109,N_12901);
nand U13330 (N_13330,N_12807,N_13084);
nor U13331 (N_13331,N_12996,N_12510);
nand U13332 (N_13332,N_12578,N_12604);
nand U13333 (N_13333,N_12821,N_12819);
and U13334 (N_13334,N_13012,N_12694);
nand U13335 (N_13335,N_12867,N_13047);
nor U13336 (N_13336,N_12849,N_12964);
or U13337 (N_13337,N_13050,N_12618);
xnor U13338 (N_13338,N_13013,N_12805);
xor U13339 (N_13339,N_12753,N_12538);
and U13340 (N_13340,N_12546,N_12711);
nand U13341 (N_13341,N_12957,N_13041);
nor U13342 (N_13342,N_12654,N_12851);
xnor U13343 (N_13343,N_12810,N_12512);
nand U13344 (N_13344,N_13004,N_12766);
or U13345 (N_13345,N_12939,N_12660);
or U13346 (N_13346,N_12737,N_12515);
nor U13347 (N_13347,N_12998,N_13099);
nor U13348 (N_13348,N_12878,N_12755);
xor U13349 (N_13349,N_12683,N_12597);
nand U13350 (N_13350,N_12756,N_12594);
and U13351 (N_13351,N_12891,N_12688);
nand U13352 (N_13352,N_12693,N_12920);
nand U13353 (N_13353,N_12613,N_12559);
nor U13354 (N_13354,N_12826,N_12798);
and U13355 (N_13355,N_12900,N_12608);
nand U13356 (N_13356,N_12933,N_13018);
or U13357 (N_13357,N_12625,N_12722);
or U13358 (N_13358,N_12887,N_12861);
and U13359 (N_13359,N_12712,N_13077);
or U13360 (N_13360,N_12871,N_13057);
xor U13361 (N_13361,N_13076,N_12869);
and U13362 (N_13362,N_12862,N_12517);
xnor U13363 (N_13363,N_12986,N_12670);
or U13364 (N_13364,N_12557,N_12563);
or U13365 (N_13365,N_12984,N_13113);
and U13366 (N_13366,N_12739,N_13090);
and U13367 (N_13367,N_13071,N_12720);
xor U13368 (N_13368,N_12554,N_12834);
xnor U13369 (N_13369,N_13066,N_13117);
nor U13370 (N_13370,N_13079,N_12695);
nor U13371 (N_13371,N_12568,N_12751);
and U13372 (N_13372,N_12848,N_12504);
xnor U13373 (N_13373,N_13008,N_13065);
nor U13374 (N_13374,N_12803,N_12955);
and U13375 (N_13375,N_12530,N_12556);
nand U13376 (N_13376,N_13022,N_12708);
nor U13377 (N_13377,N_12704,N_12535);
nand U13378 (N_13378,N_12681,N_12903);
or U13379 (N_13379,N_12924,N_12827);
and U13380 (N_13380,N_12603,N_13043);
and U13381 (N_13381,N_12925,N_12511);
xnor U13382 (N_13382,N_13083,N_12814);
nor U13383 (N_13383,N_12740,N_12978);
xnor U13384 (N_13384,N_12676,N_12716);
nor U13385 (N_13385,N_12760,N_12832);
and U13386 (N_13386,N_12979,N_12647);
and U13387 (N_13387,N_12949,N_12521);
and U13388 (N_13388,N_12995,N_12599);
nor U13389 (N_13389,N_13078,N_13032);
and U13390 (N_13390,N_12822,N_12531);
and U13391 (N_13391,N_12860,N_12724);
nand U13392 (N_13392,N_12894,N_12605);
nand U13393 (N_13393,N_12584,N_12616);
and U13394 (N_13394,N_12910,N_12659);
nor U13395 (N_13395,N_12540,N_12649);
or U13396 (N_13396,N_12841,N_12680);
and U13397 (N_13397,N_13106,N_12706);
nand U13398 (N_13398,N_12956,N_13064);
or U13399 (N_13399,N_12890,N_12717);
and U13400 (N_13400,N_12908,N_12796);
or U13401 (N_13401,N_12691,N_13098);
nor U13402 (N_13402,N_13092,N_13069);
nand U13403 (N_13403,N_12879,N_12577);
nand U13404 (N_13404,N_12700,N_12686);
nor U13405 (N_13405,N_12534,N_12518);
xor U13406 (N_13406,N_12641,N_12590);
nand U13407 (N_13407,N_12864,N_12658);
nor U13408 (N_13408,N_12734,N_12842);
nand U13409 (N_13409,N_13102,N_13067);
nand U13410 (N_13410,N_12951,N_12948);
nand U13411 (N_13411,N_12839,N_12575);
xor U13412 (N_13412,N_13054,N_13020);
nand U13413 (N_13413,N_12987,N_12931);
nor U13414 (N_13414,N_12617,N_13026);
and U13415 (N_13415,N_12953,N_12571);
nor U13416 (N_13416,N_12639,N_12883);
nor U13417 (N_13417,N_12899,N_12838);
xnor U13418 (N_13418,N_12514,N_13037);
and U13419 (N_13419,N_12919,N_12912);
nor U13420 (N_13420,N_13110,N_12800);
nand U13421 (N_13421,N_12797,N_12746);
nor U13422 (N_13422,N_12665,N_12897);
nor U13423 (N_13423,N_12699,N_12566);
and U13424 (N_13424,N_13088,N_12811);
nand U13425 (N_13425,N_12705,N_12833);
or U13426 (N_13426,N_12661,N_12585);
nand U13427 (N_13427,N_12829,N_12934);
xor U13428 (N_13428,N_12988,N_12656);
nand U13429 (N_13429,N_12758,N_12573);
nand U13430 (N_13430,N_13116,N_12844);
and U13431 (N_13431,N_12913,N_12928);
nor U13432 (N_13432,N_12994,N_12892);
nor U13433 (N_13433,N_12719,N_12553);
or U13434 (N_13434,N_13089,N_12523);
nand U13435 (N_13435,N_12651,N_12781);
and U13436 (N_13436,N_13123,N_13016);
or U13437 (N_13437,N_12865,N_12663);
nand U13438 (N_13438,N_12836,N_12511);
nor U13439 (N_13439,N_12506,N_13030);
nand U13440 (N_13440,N_12883,N_12853);
nor U13441 (N_13441,N_12916,N_12925);
nand U13442 (N_13442,N_13124,N_13019);
nand U13443 (N_13443,N_12603,N_12965);
nand U13444 (N_13444,N_12589,N_12956);
xor U13445 (N_13445,N_12996,N_12998);
and U13446 (N_13446,N_12689,N_13018);
xnor U13447 (N_13447,N_12794,N_13121);
or U13448 (N_13448,N_12883,N_12699);
and U13449 (N_13449,N_12872,N_12564);
xnor U13450 (N_13450,N_13009,N_13066);
xor U13451 (N_13451,N_12876,N_12621);
xor U13452 (N_13452,N_12708,N_12518);
and U13453 (N_13453,N_12612,N_12509);
or U13454 (N_13454,N_12546,N_12993);
and U13455 (N_13455,N_12700,N_13121);
nand U13456 (N_13456,N_13000,N_13094);
xnor U13457 (N_13457,N_12538,N_12862);
nor U13458 (N_13458,N_12986,N_13116);
or U13459 (N_13459,N_12986,N_13011);
xnor U13460 (N_13460,N_12521,N_13117);
xnor U13461 (N_13461,N_12850,N_12984);
nand U13462 (N_13462,N_12870,N_12588);
nor U13463 (N_13463,N_12886,N_12822);
or U13464 (N_13464,N_12880,N_12966);
or U13465 (N_13465,N_13116,N_12948);
or U13466 (N_13466,N_12695,N_12597);
nor U13467 (N_13467,N_12831,N_12754);
nor U13468 (N_13468,N_12671,N_13080);
xnor U13469 (N_13469,N_12816,N_12857);
and U13470 (N_13470,N_12906,N_13076);
or U13471 (N_13471,N_12519,N_12837);
xnor U13472 (N_13472,N_12868,N_12672);
xor U13473 (N_13473,N_12922,N_12737);
and U13474 (N_13474,N_13020,N_13090);
nor U13475 (N_13475,N_12769,N_12926);
nor U13476 (N_13476,N_12740,N_12618);
and U13477 (N_13477,N_12844,N_12514);
xor U13478 (N_13478,N_12799,N_12984);
or U13479 (N_13479,N_13055,N_12770);
and U13480 (N_13480,N_12916,N_12573);
xnor U13481 (N_13481,N_12538,N_13080);
or U13482 (N_13482,N_12669,N_12986);
nor U13483 (N_13483,N_12907,N_12801);
nand U13484 (N_13484,N_12720,N_12581);
nand U13485 (N_13485,N_12599,N_12513);
xnor U13486 (N_13486,N_12553,N_12951);
nor U13487 (N_13487,N_13038,N_12667);
or U13488 (N_13488,N_12859,N_12986);
nand U13489 (N_13489,N_13063,N_12654);
nor U13490 (N_13490,N_12852,N_12531);
nand U13491 (N_13491,N_13063,N_12784);
nor U13492 (N_13492,N_12658,N_13070);
nand U13493 (N_13493,N_12561,N_12903);
xnor U13494 (N_13494,N_12786,N_12910);
nor U13495 (N_13495,N_12682,N_12852);
and U13496 (N_13496,N_12652,N_13056);
nand U13497 (N_13497,N_13009,N_13002);
nand U13498 (N_13498,N_12699,N_12748);
nor U13499 (N_13499,N_12814,N_13019);
and U13500 (N_13500,N_12670,N_13053);
nand U13501 (N_13501,N_13096,N_12946);
nor U13502 (N_13502,N_12868,N_12767);
nor U13503 (N_13503,N_13027,N_12902);
nor U13504 (N_13504,N_12920,N_12837);
nand U13505 (N_13505,N_13088,N_13004);
nand U13506 (N_13506,N_12859,N_12642);
nor U13507 (N_13507,N_12771,N_12838);
and U13508 (N_13508,N_12677,N_12824);
xor U13509 (N_13509,N_12738,N_12913);
or U13510 (N_13510,N_12898,N_12704);
xnor U13511 (N_13511,N_12800,N_12539);
nor U13512 (N_13512,N_12681,N_13052);
nor U13513 (N_13513,N_12538,N_13074);
nor U13514 (N_13514,N_12713,N_12604);
and U13515 (N_13515,N_12843,N_12855);
nand U13516 (N_13516,N_12826,N_13009);
and U13517 (N_13517,N_12697,N_12565);
nor U13518 (N_13518,N_12639,N_13061);
and U13519 (N_13519,N_12952,N_12945);
nor U13520 (N_13520,N_12753,N_12912);
nor U13521 (N_13521,N_12690,N_12675);
xnor U13522 (N_13522,N_12719,N_13082);
and U13523 (N_13523,N_12986,N_13094);
and U13524 (N_13524,N_13107,N_12960);
xnor U13525 (N_13525,N_12564,N_13036);
xnor U13526 (N_13526,N_13063,N_12541);
and U13527 (N_13527,N_12621,N_12820);
xnor U13528 (N_13528,N_12920,N_13051);
and U13529 (N_13529,N_13089,N_12602);
nor U13530 (N_13530,N_12632,N_12754);
or U13531 (N_13531,N_12568,N_13028);
nand U13532 (N_13532,N_12840,N_12784);
nand U13533 (N_13533,N_12804,N_12669);
nand U13534 (N_13534,N_12820,N_12527);
nand U13535 (N_13535,N_12761,N_12648);
nand U13536 (N_13536,N_12664,N_12673);
or U13537 (N_13537,N_13109,N_13045);
or U13538 (N_13538,N_12508,N_13007);
xor U13539 (N_13539,N_12631,N_12756);
xnor U13540 (N_13540,N_12545,N_12720);
nor U13541 (N_13541,N_12857,N_13049);
or U13542 (N_13542,N_12718,N_12635);
and U13543 (N_13543,N_13060,N_13071);
and U13544 (N_13544,N_13012,N_13044);
or U13545 (N_13545,N_12513,N_12734);
or U13546 (N_13546,N_12756,N_12879);
nand U13547 (N_13547,N_12618,N_12834);
nor U13548 (N_13548,N_12913,N_13000);
and U13549 (N_13549,N_12735,N_12751);
nand U13550 (N_13550,N_12783,N_13031);
and U13551 (N_13551,N_12744,N_12985);
and U13552 (N_13552,N_12532,N_12753);
and U13553 (N_13553,N_12865,N_12901);
xnor U13554 (N_13554,N_12629,N_12940);
and U13555 (N_13555,N_12578,N_13112);
xor U13556 (N_13556,N_12526,N_13115);
nand U13557 (N_13557,N_13058,N_12799);
xnor U13558 (N_13558,N_13108,N_12973);
xnor U13559 (N_13559,N_12685,N_12695);
and U13560 (N_13560,N_12725,N_12551);
nor U13561 (N_13561,N_12985,N_12785);
nand U13562 (N_13562,N_12792,N_12577);
nor U13563 (N_13563,N_12772,N_12895);
or U13564 (N_13564,N_12776,N_13123);
nand U13565 (N_13565,N_12833,N_12611);
xnor U13566 (N_13566,N_12939,N_12565);
and U13567 (N_13567,N_13053,N_12613);
xor U13568 (N_13568,N_12512,N_13084);
and U13569 (N_13569,N_12751,N_13103);
nand U13570 (N_13570,N_13055,N_12719);
xor U13571 (N_13571,N_12954,N_12757);
or U13572 (N_13572,N_12621,N_12736);
or U13573 (N_13573,N_12897,N_12951);
nand U13574 (N_13574,N_12517,N_12996);
and U13575 (N_13575,N_12521,N_12799);
nand U13576 (N_13576,N_12640,N_12670);
and U13577 (N_13577,N_12957,N_12575);
or U13578 (N_13578,N_12610,N_12865);
nor U13579 (N_13579,N_12792,N_13048);
and U13580 (N_13580,N_12979,N_12940);
nand U13581 (N_13581,N_12703,N_12639);
and U13582 (N_13582,N_12651,N_12913);
xor U13583 (N_13583,N_12949,N_12535);
and U13584 (N_13584,N_12719,N_13014);
and U13585 (N_13585,N_13074,N_12875);
xnor U13586 (N_13586,N_12879,N_12931);
xnor U13587 (N_13587,N_12989,N_13084);
nor U13588 (N_13588,N_12563,N_12797);
nor U13589 (N_13589,N_12957,N_12557);
xor U13590 (N_13590,N_13052,N_12707);
nor U13591 (N_13591,N_12583,N_13027);
nand U13592 (N_13592,N_12568,N_12720);
nor U13593 (N_13593,N_13030,N_12759);
and U13594 (N_13594,N_13083,N_12683);
xor U13595 (N_13595,N_12817,N_12972);
and U13596 (N_13596,N_12628,N_12738);
nand U13597 (N_13597,N_12805,N_12837);
nand U13598 (N_13598,N_12693,N_13060);
xor U13599 (N_13599,N_13109,N_12615);
xnor U13600 (N_13600,N_12561,N_12984);
xor U13601 (N_13601,N_12622,N_12930);
and U13602 (N_13602,N_12614,N_12901);
nand U13603 (N_13603,N_13069,N_12524);
and U13604 (N_13604,N_13056,N_12814);
nand U13605 (N_13605,N_12843,N_12951);
xor U13606 (N_13606,N_13073,N_12955);
xor U13607 (N_13607,N_13027,N_12938);
nor U13608 (N_13608,N_13098,N_12789);
or U13609 (N_13609,N_12762,N_12552);
nand U13610 (N_13610,N_13082,N_12700);
or U13611 (N_13611,N_12752,N_12704);
nor U13612 (N_13612,N_12944,N_12750);
xor U13613 (N_13613,N_13050,N_12547);
xnor U13614 (N_13614,N_12575,N_13017);
xnor U13615 (N_13615,N_12794,N_12744);
nand U13616 (N_13616,N_12512,N_12950);
xnor U13617 (N_13617,N_12632,N_12866);
xnor U13618 (N_13618,N_13070,N_12768);
xor U13619 (N_13619,N_12865,N_12508);
nand U13620 (N_13620,N_12929,N_12819);
nor U13621 (N_13621,N_12503,N_12597);
xor U13622 (N_13622,N_12767,N_12604);
xor U13623 (N_13623,N_12873,N_13025);
nor U13624 (N_13624,N_13123,N_13099);
nand U13625 (N_13625,N_12805,N_12718);
nand U13626 (N_13626,N_12882,N_12964);
nand U13627 (N_13627,N_12880,N_12801);
or U13628 (N_13628,N_12883,N_13098);
xnor U13629 (N_13629,N_12730,N_12672);
nand U13630 (N_13630,N_12704,N_12884);
nor U13631 (N_13631,N_13099,N_12849);
nor U13632 (N_13632,N_12547,N_12713);
xnor U13633 (N_13633,N_12833,N_12940);
and U13634 (N_13634,N_12877,N_12728);
xor U13635 (N_13635,N_12803,N_12562);
or U13636 (N_13636,N_12870,N_12582);
or U13637 (N_13637,N_12941,N_12953);
nor U13638 (N_13638,N_12798,N_12763);
xor U13639 (N_13639,N_12561,N_12587);
nand U13640 (N_13640,N_12892,N_13103);
xnor U13641 (N_13641,N_13025,N_12906);
or U13642 (N_13642,N_12596,N_12637);
or U13643 (N_13643,N_13094,N_12690);
and U13644 (N_13644,N_12520,N_12575);
or U13645 (N_13645,N_12703,N_12704);
nand U13646 (N_13646,N_12583,N_13071);
nor U13647 (N_13647,N_12725,N_12786);
nor U13648 (N_13648,N_12569,N_12672);
xor U13649 (N_13649,N_13063,N_12974);
xnor U13650 (N_13650,N_12989,N_13070);
nand U13651 (N_13651,N_12848,N_12816);
nand U13652 (N_13652,N_12918,N_12598);
xor U13653 (N_13653,N_12656,N_13034);
and U13654 (N_13654,N_12894,N_12798);
nand U13655 (N_13655,N_13019,N_12715);
and U13656 (N_13656,N_12977,N_13020);
xnor U13657 (N_13657,N_12793,N_12695);
xnor U13658 (N_13658,N_12521,N_12831);
or U13659 (N_13659,N_12613,N_12775);
or U13660 (N_13660,N_12503,N_12834);
or U13661 (N_13661,N_12773,N_12953);
nor U13662 (N_13662,N_12609,N_12909);
and U13663 (N_13663,N_12740,N_12591);
xnor U13664 (N_13664,N_13095,N_12824);
xor U13665 (N_13665,N_13078,N_12731);
or U13666 (N_13666,N_12535,N_12741);
and U13667 (N_13667,N_12699,N_12995);
and U13668 (N_13668,N_12913,N_12800);
xnor U13669 (N_13669,N_12713,N_12808);
or U13670 (N_13670,N_12798,N_12707);
nand U13671 (N_13671,N_12702,N_12865);
and U13672 (N_13672,N_12659,N_12941);
or U13673 (N_13673,N_12864,N_12906);
or U13674 (N_13674,N_12507,N_12981);
nand U13675 (N_13675,N_12748,N_12680);
nor U13676 (N_13676,N_12636,N_12776);
or U13677 (N_13677,N_12786,N_12584);
nand U13678 (N_13678,N_12613,N_12574);
or U13679 (N_13679,N_12607,N_12541);
nor U13680 (N_13680,N_12648,N_12540);
or U13681 (N_13681,N_12806,N_12538);
or U13682 (N_13682,N_13117,N_12878);
nand U13683 (N_13683,N_13114,N_12579);
and U13684 (N_13684,N_12998,N_12617);
xnor U13685 (N_13685,N_12718,N_12714);
nand U13686 (N_13686,N_12899,N_13040);
or U13687 (N_13687,N_12550,N_13069);
nand U13688 (N_13688,N_12934,N_12831);
or U13689 (N_13689,N_12535,N_12586);
nor U13690 (N_13690,N_12608,N_12516);
nand U13691 (N_13691,N_12869,N_12779);
and U13692 (N_13692,N_13078,N_13063);
nor U13693 (N_13693,N_12963,N_12686);
nor U13694 (N_13694,N_12510,N_12813);
nor U13695 (N_13695,N_12725,N_12841);
and U13696 (N_13696,N_13087,N_12985);
and U13697 (N_13697,N_12747,N_12611);
nand U13698 (N_13698,N_12910,N_12500);
and U13699 (N_13699,N_13059,N_12866);
xnor U13700 (N_13700,N_12999,N_12905);
nor U13701 (N_13701,N_12995,N_12665);
xnor U13702 (N_13702,N_12539,N_12690);
and U13703 (N_13703,N_12526,N_12840);
xor U13704 (N_13704,N_12653,N_12588);
nand U13705 (N_13705,N_13103,N_13076);
nor U13706 (N_13706,N_12924,N_12563);
nor U13707 (N_13707,N_12774,N_12514);
nor U13708 (N_13708,N_12793,N_13000);
or U13709 (N_13709,N_12883,N_12976);
xor U13710 (N_13710,N_12715,N_13089);
nand U13711 (N_13711,N_12899,N_12888);
or U13712 (N_13712,N_12531,N_12667);
nand U13713 (N_13713,N_12577,N_12872);
or U13714 (N_13714,N_12808,N_12511);
and U13715 (N_13715,N_12624,N_12789);
and U13716 (N_13716,N_12640,N_12720);
and U13717 (N_13717,N_12741,N_12879);
or U13718 (N_13718,N_13116,N_12760);
xor U13719 (N_13719,N_12684,N_12975);
nor U13720 (N_13720,N_12941,N_12546);
xnor U13721 (N_13721,N_12874,N_12989);
nor U13722 (N_13722,N_12869,N_12885);
nor U13723 (N_13723,N_12736,N_13036);
or U13724 (N_13724,N_12973,N_12754);
xnor U13725 (N_13725,N_12852,N_12609);
or U13726 (N_13726,N_12968,N_13051);
and U13727 (N_13727,N_12542,N_13099);
nand U13728 (N_13728,N_12659,N_12798);
or U13729 (N_13729,N_12921,N_13016);
or U13730 (N_13730,N_12552,N_12871);
nor U13731 (N_13731,N_12888,N_12590);
nand U13732 (N_13732,N_12759,N_12791);
and U13733 (N_13733,N_12774,N_12855);
xor U13734 (N_13734,N_12772,N_12826);
xnor U13735 (N_13735,N_12562,N_12542);
xor U13736 (N_13736,N_12681,N_13114);
nor U13737 (N_13737,N_12834,N_12896);
nand U13738 (N_13738,N_12997,N_12514);
xor U13739 (N_13739,N_12784,N_12605);
nand U13740 (N_13740,N_12877,N_12757);
and U13741 (N_13741,N_12549,N_13086);
and U13742 (N_13742,N_12514,N_12582);
nand U13743 (N_13743,N_12979,N_12599);
and U13744 (N_13744,N_12917,N_12676);
nor U13745 (N_13745,N_12718,N_12881);
xor U13746 (N_13746,N_12670,N_12917);
or U13747 (N_13747,N_12678,N_12966);
xor U13748 (N_13748,N_13079,N_12794);
nand U13749 (N_13749,N_12817,N_12872);
or U13750 (N_13750,N_13468,N_13674);
and U13751 (N_13751,N_13205,N_13542);
nor U13752 (N_13752,N_13214,N_13248);
and U13753 (N_13753,N_13316,N_13356);
nor U13754 (N_13754,N_13151,N_13475);
xnor U13755 (N_13755,N_13638,N_13389);
xor U13756 (N_13756,N_13278,N_13559);
nor U13757 (N_13757,N_13155,N_13552);
nor U13758 (N_13758,N_13364,N_13661);
nand U13759 (N_13759,N_13716,N_13259);
and U13760 (N_13760,N_13533,N_13386);
nor U13761 (N_13761,N_13195,N_13613);
nor U13762 (N_13762,N_13376,N_13518);
xnor U13763 (N_13763,N_13403,N_13460);
and U13764 (N_13764,N_13299,N_13422);
nor U13765 (N_13765,N_13623,N_13747);
and U13766 (N_13766,N_13605,N_13597);
nand U13767 (N_13767,N_13304,N_13560);
and U13768 (N_13768,N_13230,N_13586);
or U13769 (N_13769,N_13558,N_13228);
or U13770 (N_13770,N_13235,N_13295);
and U13771 (N_13771,N_13244,N_13440);
nor U13772 (N_13772,N_13175,N_13372);
nor U13773 (N_13773,N_13226,N_13131);
xor U13774 (N_13774,N_13261,N_13222);
and U13775 (N_13775,N_13712,N_13187);
xor U13776 (N_13776,N_13578,N_13240);
and U13777 (N_13777,N_13448,N_13388);
xor U13778 (N_13778,N_13576,N_13333);
nor U13779 (N_13779,N_13251,N_13441);
nand U13780 (N_13780,N_13341,N_13132);
and U13781 (N_13781,N_13434,N_13643);
or U13782 (N_13782,N_13238,N_13503);
nand U13783 (N_13783,N_13289,N_13365);
or U13784 (N_13784,N_13306,N_13508);
and U13785 (N_13785,N_13286,N_13433);
or U13786 (N_13786,N_13413,N_13609);
nor U13787 (N_13787,N_13129,N_13396);
nand U13788 (N_13788,N_13521,N_13621);
xor U13789 (N_13789,N_13672,N_13491);
and U13790 (N_13790,N_13406,N_13449);
or U13791 (N_13791,N_13733,N_13727);
nand U13792 (N_13792,N_13277,N_13344);
and U13793 (N_13793,N_13426,N_13272);
and U13794 (N_13794,N_13375,N_13417);
and U13795 (N_13795,N_13540,N_13152);
or U13796 (N_13796,N_13671,N_13651);
nor U13797 (N_13797,N_13383,N_13711);
and U13798 (N_13798,N_13204,N_13203);
nor U13799 (N_13799,N_13739,N_13557);
and U13800 (N_13800,N_13665,N_13615);
or U13801 (N_13801,N_13703,N_13349);
nor U13802 (N_13802,N_13534,N_13652);
xor U13803 (N_13803,N_13338,N_13469);
nor U13804 (N_13804,N_13271,N_13276);
nand U13805 (N_13805,N_13183,N_13287);
or U13806 (N_13806,N_13630,N_13477);
or U13807 (N_13807,N_13546,N_13258);
nor U13808 (N_13808,N_13218,N_13342);
or U13809 (N_13809,N_13416,N_13685);
nand U13810 (N_13810,N_13208,N_13385);
and U13811 (N_13811,N_13134,N_13487);
nor U13812 (N_13812,N_13328,N_13157);
nor U13813 (N_13813,N_13439,N_13718);
nand U13814 (N_13814,N_13522,N_13331);
and U13815 (N_13815,N_13404,N_13186);
xor U13816 (N_13816,N_13357,N_13162);
xor U13817 (N_13817,N_13516,N_13174);
nor U13818 (N_13818,N_13523,N_13444);
nor U13819 (N_13819,N_13329,N_13141);
xnor U13820 (N_13820,N_13153,N_13177);
or U13821 (N_13821,N_13280,N_13478);
and U13822 (N_13822,N_13352,N_13670);
or U13823 (N_13823,N_13462,N_13721);
nand U13824 (N_13824,N_13362,N_13154);
and U13825 (N_13825,N_13572,N_13749);
or U13826 (N_13826,N_13594,N_13407);
or U13827 (N_13827,N_13683,N_13528);
or U13828 (N_13828,N_13243,N_13506);
nor U13829 (N_13829,N_13419,N_13648);
or U13830 (N_13830,N_13591,N_13150);
nand U13831 (N_13831,N_13346,N_13744);
xor U13832 (N_13832,N_13679,N_13313);
nand U13833 (N_13833,N_13359,N_13464);
nor U13834 (N_13834,N_13392,N_13645);
and U13835 (N_13835,N_13740,N_13178);
xor U13836 (N_13836,N_13361,N_13428);
xnor U13837 (N_13837,N_13380,N_13595);
nor U13838 (N_13838,N_13319,N_13143);
nand U13839 (N_13839,N_13499,N_13147);
or U13840 (N_13840,N_13720,N_13371);
or U13841 (N_13841,N_13476,N_13192);
or U13842 (N_13842,N_13659,N_13320);
or U13843 (N_13843,N_13321,N_13492);
and U13844 (N_13844,N_13411,N_13624);
or U13845 (N_13845,N_13725,N_13505);
or U13846 (N_13846,N_13418,N_13291);
nor U13847 (N_13847,N_13538,N_13577);
xor U13848 (N_13848,N_13254,N_13351);
or U13849 (N_13849,N_13145,N_13582);
nand U13850 (N_13850,N_13260,N_13436);
or U13851 (N_13851,N_13430,N_13710);
nand U13852 (N_13852,N_13590,N_13657);
or U13853 (N_13853,N_13387,N_13736);
or U13854 (N_13854,N_13237,N_13191);
or U13855 (N_13855,N_13457,N_13746);
or U13856 (N_13856,N_13742,N_13539);
nor U13857 (N_13857,N_13748,N_13507);
xnor U13858 (N_13858,N_13250,N_13223);
and U13859 (N_13859,N_13335,N_13513);
nand U13860 (N_13860,N_13379,N_13625);
xor U13861 (N_13861,N_13581,N_13678);
and U13862 (N_13862,N_13398,N_13473);
xor U13863 (N_13863,N_13495,N_13641);
nor U13864 (N_13864,N_13166,N_13239);
xnor U13865 (N_13865,N_13532,N_13544);
or U13866 (N_13866,N_13315,N_13714);
xor U13867 (N_13867,N_13662,N_13587);
xnor U13868 (N_13868,N_13517,N_13241);
nand U13869 (N_13869,N_13179,N_13337);
xnor U13870 (N_13870,N_13451,N_13611);
nor U13871 (N_13871,N_13381,N_13599);
nor U13872 (N_13872,N_13728,N_13137);
nand U13873 (N_13873,N_13202,N_13189);
nand U13874 (N_13874,N_13269,N_13360);
xor U13875 (N_13875,N_13606,N_13181);
or U13876 (N_13876,N_13563,N_13706);
nand U13877 (N_13877,N_13745,N_13246);
xnor U13878 (N_13878,N_13626,N_13501);
and U13879 (N_13879,N_13323,N_13729);
or U13880 (N_13880,N_13281,N_13663);
and U13881 (N_13881,N_13236,N_13160);
or U13882 (N_13882,N_13447,N_13676);
nor U13883 (N_13883,N_13588,N_13694);
nor U13884 (N_13884,N_13571,N_13474);
and U13885 (N_13885,N_13432,N_13301);
nor U13886 (N_13886,N_13410,N_13481);
and U13887 (N_13887,N_13666,N_13322);
nand U13888 (N_13888,N_13483,N_13435);
nand U13889 (N_13889,N_13330,N_13325);
and U13890 (N_13890,N_13128,N_13567);
or U13891 (N_13891,N_13515,N_13391);
nand U13892 (N_13892,N_13705,N_13395);
and U13893 (N_13893,N_13722,N_13732);
or U13894 (N_13894,N_13270,N_13498);
nor U13895 (N_13895,N_13135,N_13427);
nand U13896 (N_13896,N_13194,N_13690);
or U13897 (N_13897,N_13358,N_13536);
nand U13898 (N_13898,N_13514,N_13656);
or U13899 (N_13899,N_13327,N_13632);
and U13900 (N_13900,N_13224,N_13631);
xnor U13901 (N_13901,N_13168,N_13622);
xnor U13902 (N_13902,N_13482,N_13125);
nor U13903 (N_13903,N_13283,N_13456);
nand U13904 (N_13904,N_13575,N_13568);
or U13905 (N_13905,N_13198,N_13212);
and U13906 (N_13906,N_13541,N_13339);
xnor U13907 (N_13907,N_13215,N_13693);
xor U13908 (N_13908,N_13136,N_13555);
or U13909 (N_13909,N_13408,N_13170);
or U13910 (N_13910,N_13138,N_13580);
nor U13911 (N_13911,N_13221,N_13635);
xnor U13912 (N_13912,N_13308,N_13619);
xnor U13913 (N_13913,N_13234,N_13303);
xor U13914 (N_13914,N_13500,N_13616);
xor U13915 (N_13915,N_13696,N_13470);
and U13916 (N_13916,N_13442,N_13188);
nand U13917 (N_13917,N_13680,N_13600);
xnor U13918 (N_13918,N_13553,N_13545);
xor U13919 (N_13919,N_13564,N_13642);
nor U13920 (N_13920,N_13730,N_13159);
nor U13921 (N_13921,N_13264,N_13267);
nor U13922 (N_13922,N_13309,N_13405);
xor U13923 (N_13923,N_13585,N_13658);
xor U13924 (N_13924,N_13378,N_13343);
or U13925 (N_13925,N_13547,N_13247);
and U13926 (N_13926,N_13496,N_13525);
nand U13927 (N_13927,N_13646,N_13377);
nand U13928 (N_13928,N_13190,N_13731);
or U13929 (N_13929,N_13604,N_13139);
nand U13930 (N_13930,N_13163,N_13429);
and U13931 (N_13931,N_13566,N_13282);
and U13932 (N_13932,N_13681,N_13458);
or U13933 (N_13933,N_13737,N_13172);
nand U13934 (N_13934,N_13437,N_13565);
xor U13935 (N_13935,N_13704,N_13726);
nor U13936 (N_13936,N_13471,N_13185);
xor U13937 (N_13937,N_13180,N_13412);
xor U13938 (N_13938,N_13414,N_13312);
nor U13939 (N_13939,N_13164,N_13373);
nor U13940 (N_13940,N_13569,N_13618);
and U13941 (N_13941,N_13452,N_13397);
or U13942 (N_13942,N_13708,N_13682);
xor U13943 (N_13943,N_13400,N_13562);
nor U13944 (N_13944,N_13206,N_13146);
nor U13945 (N_13945,N_13453,N_13715);
nor U13946 (N_13946,N_13573,N_13691);
or U13947 (N_13947,N_13601,N_13142);
xnor U13948 (N_13948,N_13654,N_13574);
or U13949 (N_13949,N_13133,N_13288);
nand U13950 (N_13950,N_13465,N_13485);
or U13951 (N_13951,N_13161,N_13420);
and U13952 (N_13952,N_13265,N_13367);
or U13953 (N_13953,N_13273,N_13274);
xor U13954 (N_13954,N_13700,N_13345);
nand U13955 (N_13955,N_13698,N_13326);
xor U13956 (N_13956,N_13689,N_13374);
and U13957 (N_13957,N_13660,N_13628);
nor U13958 (N_13958,N_13598,N_13310);
or U13959 (N_13959,N_13614,N_13348);
nand U13960 (N_13960,N_13231,N_13617);
or U13961 (N_13961,N_13199,N_13509);
nor U13962 (N_13962,N_13292,N_13561);
or U13963 (N_13963,N_13424,N_13263);
nand U13964 (N_13964,N_13461,N_13233);
or U13965 (N_13965,N_13149,N_13347);
and U13966 (N_13966,N_13255,N_13354);
or U13967 (N_13967,N_13550,N_13519);
nor U13968 (N_13968,N_13423,N_13253);
xor U13969 (N_13969,N_13493,N_13220);
xnor U13970 (N_13970,N_13548,N_13719);
or U13971 (N_13971,N_13445,N_13667);
and U13972 (N_13972,N_13370,N_13596);
nand U13973 (N_13973,N_13664,N_13637);
nand U13974 (N_13974,N_13210,N_13504);
nor U13975 (N_13975,N_13232,N_13511);
nor U13976 (N_13976,N_13402,N_13317);
or U13977 (N_13977,N_13252,N_13684);
xnor U13978 (N_13978,N_13455,N_13620);
or U13979 (N_13979,N_13290,N_13294);
xor U13980 (N_13980,N_13583,N_13543);
or U13981 (N_13981,N_13687,N_13479);
and U13982 (N_13982,N_13285,N_13201);
and U13983 (N_13983,N_13584,N_13697);
or U13984 (N_13984,N_13297,N_13302);
and U13985 (N_13985,N_13130,N_13293);
nand U13986 (N_13986,N_13529,N_13298);
and U13987 (N_13987,N_13366,N_13655);
or U13988 (N_13988,N_13612,N_13401);
nand U13989 (N_13989,N_13421,N_13488);
or U13990 (N_13990,N_13355,N_13490);
nand U13991 (N_13991,N_13296,N_13717);
nor U13992 (N_13992,N_13602,N_13467);
xor U13993 (N_13993,N_13156,N_13211);
and U13994 (N_13994,N_13318,N_13275);
nor U13995 (N_13995,N_13314,N_13394);
xor U13996 (N_13996,N_13535,N_13709);
and U13997 (N_13997,N_13369,N_13551);
or U13998 (N_13998,N_13724,N_13382);
nand U13999 (N_13999,N_13639,N_13673);
or U14000 (N_14000,N_13686,N_13593);
and U14001 (N_14001,N_13677,N_13409);
nor U14002 (N_14002,N_13256,N_13207);
or U14003 (N_14003,N_13171,N_13741);
xor U14004 (N_14004,N_13363,N_13520);
xnor U14005 (N_14005,N_13209,N_13140);
xor U14006 (N_14006,N_13393,N_13549);
nand U14007 (N_14007,N_13443,N_13334);
or U14008 (N_14008,N_13305,N_13459);
and U14009 (N_14009,N_13647,N_13669);
and U14010 (N_14010,N_13350,N_13200);
and U14011 (N_14011,N_13332,N_13300);
and U14012 (N_14012,N_13158,N_13702);
or U14013 (N_14013,N_13148,N_13489);
nor U14014 (N_14014,N_13699,N_13353);
nand U14015 (N_14015,N_13266,N_13307);
and U14016 (N_14016,N_13384,N_13688);
nand U14017 (N_14017,N_13653,N_13390);
and U14018 (N_14018,N_13399,N_13512);
nor U14019 (N_14019,N_13225,N_13668);
and U14020 (N_14020,N_13570,N_13494);
nand U14021 (N_14021,N_13446,N_13324);
or U14022 (N_14022,N_13182,N_13219);
nor U14023 (N_14023,N_13227,N_13636);
and U14024 (N_14024,N_13640,N_13193);
xnor U14025 (N_14025,N_13579,N_13675);
nand U14026 (N_14026,N_13184,N_13216);
xnor U14027 (N_14027,N_13734,N_13425);
and U14028 (N_14028,N_13213,N_13530);
or U14029 (N_14029,N_13268,N_13242);
nor U14030 (N_14030,N_13450,N_13249);
or U14031 (N_14031,N_13486,N_13217);
nor U14032 (N_14032,N_13589,N_13279);
or U14033 (N_14033,N_13634,N_13262);
or U14034 (N_14034,N_13284,N_13603);
nor U14035 (N_14035,N_13510,N_13463);
xnor U14036 (N_14036,N_13497,N_13472);
xnor U14037 (N_14037,N_13176,N_13524);
nand U14038 (N_14038,N_13610,N_13257);
nand U14039 (N_14039,N_13196,N_13415);
nand U14040 (N_14040,N_13738,N_13502);
nor U14041 (N_14041,N_13629,N_13531);
nand U14042 (N_14042,N_13556,N_13340);
or U14043 (N_14043,N_13554,N_13707);
or U14044 (N_14044,N_13311,N_13336);
nor U14045 (N_14045,N_13650,N_13592);
xnor U14046 (N_14046,N_13438,N_13607);
or U14047 (N_14047,N_13197,N_13627);
nand U14048 (N_14048,N_13537,N_13173);
and U14049 (N_14049,N_13431,N_13713);
xor U14050 (N_14050,N_13480,N_13526);
nand U14051 (N_14051,N_13723,N_13165);
or U14052 (N_14052,N_13701,N_13368);
nor U14053 (N_14053,N_13644,N_13169);
nor U14054 (N_14054,N_13692,N_13126);
nand U14055 (N_14055,N_13527,N_13466);
nand U14056 (N_14056,N_13127,N_13608);
nand U14057 (N_14057,N_13695,N_13454);
and U14058 (N_14058,N_13484,N_13735);
or U14059 (N_14059,N_13229,N_13743);
nand U14060 (N_14060,N_13167,N_13245);
and U14061 (N_14061,N_13144,N_13633);
and U14062 (N_14062,N_13649,N_13483);
or U14063 (N_14063,N_13689,N_13351);
and U14064 (N_14064,N_13580,N_13746);
xor U14065 (N_14065,N_13448,N_13402);
nor U14066 (N_14066,N_13154,N_13254);
nand U14067 (N_14067,N_13421,N_13416);
xnor U14068 (N_14068,N_13248,N_13486);
nand U14069 (N_14069,N_13257,N_13485);
xnor U14070 (N_14070,N_13593,N_13199);
nand U14071 (N_14071,N_13697,N_13725);
nand U14072 (N_14072,N_13175,N_13568);
or U14073 (N_14073,N_13220,N_13481);
nand U14074 (N_14074,N_13323,N_13417);
and U14075 (N_14075,N_13692,N_13548);
and U14076 (N_14076,N_13685,N_13292);
and U14077 (N_14077,N_13474,N_13508);
nand U14078 (N_14078,N_13135,N_13276);
xnor U14079 (N_14079,N_13377,N_13340);
nand U14080 (N_14080,N_13739,N_13386);
nand U14081 (N_14081,N_13739,N_13388);
nor U14082 (N_14082,N_13605,N_13370);
nor U14083 (N_14083,N_13215,N_13314);
nand U14084 (N_14084,N_13374,N_13570);
or U14085 (N_14085,N_13386,N_13690);
nand U14086 (N_14086,N_13275,N_13368);
or U14087 (N_14087,N_13574,N_13397);
nand U14088 (N_14088,N_13253,N_13546);
xnor U14089 (N_14089,N_13701,N_13248);
and U14090 (N_14090,N_13170,N_13459);
nor U14091 (N_14091,N_13539,N_13417);
and U14092 (N_14092,N_13429,N_13142);
nand U14093 (N_14093,N_13369,N_13212);
nor U14094 (N_14094,N_13401,N_13364);
or U14095 (N_14095,N_13203,N_13452);
xnor U14096 (N_14096,N_13702,N_13272);
nand U14097 (N_14097,N_13333,N_13727);
xnor U14098 (N_14098,N_13475,N_13665);
nand U14099 (N_14099,N_13560,N_13738);
nor U14100 (N_14100,N_13496,N_13126);
nor U14101 (N_14101,N_13666,N_13496);
and U14102 (N_14102,N_13133,N_13197);
and U14103 (N_14103,N_13572,N_13612);
nor U14104 (N_14104,N_13466,N_13528);
xor U14105 (N_14105,N_13659,N_13127);
nor U14106 (N_14106,N_13128,N_13440);
nand U14107 (N_14107,N_13161,N_13146);
xor U14108 (N_14108,N_13154,N_13266);
nor U14109 (N_14109,N_13619,N_13336);
or U14110 (N_14110,N_13404,N_13486);
nand U14111 (N_14111,N_13679,N_13611);
and U14112 (N_14112,N_13296,N_13436);
xor U14113 (N_14113,N_13326,N_13169);
xor U14114 (N_14114,N_13327,N_13739);
nand U14115 (N_14115,N_13526,N_13140);
nor U14116 (N_14116,N_13746,N_13260);
and U14117 (N_14117,N_13347,N_13586);
or U14118 (N_14118,N_13498,N_13724);
nand U14119 (N_14119,N_13458,N_13187);
xnor U14120 (N_14120,N_13361,N_13368);
and U14121 (N_14121,N_13538,N_13387);
or U14122 (N_14122,N_13413,N_13175);
and U14123 (N_14123,N_13699,N_13712);
and U14124 (N_14124,N_13181,N_13474);
xnor U14125 (N_14125,N_13359,N_13287);
nand U14126 (N_14126,N_13550,N_13688);
or U14127 (N_14127,N_13344,N_13539);
xor U14128 (N_14128,N_13497,N_13708);
and U14129 (N_14129,N_13549,N_13337);
nand U14130 (N_14130,N_13701,N_13287);
and U14131 (N_14131,N_13223,N_13455);
nor U14132 (N_14132,N_13717,N_13567);
or U14133 (N_14133,N_13599,N_13447);
nor U14134 (N_14134,N_13423,N_13574);
xnor U14135 (N_14135,N_13473,N_13382);
nand U14136 (N_14136,N_13153,N_13355);
and U14137 (N_14137,N_13479,N_13670);
and U14138 (N_14138,N_13671,N_13332);
xor U14139 (N_14139,N_13566,N_13338);
nand U14140 (N_14140,N_13409,N_13718);
nor U14141 (N_14141,N_13736,N_13537);
nand U14142 (N_14142,N_13355,N_13359);
and U14143 (N_14143,N_13438,N_13445);
or U14144 (N_14144,N_13549,N_13233);
and U14145 (N_14145,N_13300,N_13546);
xor U14146 (N_14146,N_13222,N_13292);
xor U14147 (N_14147,N_13499,N_13432);
and U14148 (N_14148,N_13612,N_13215);
xor U14149 (N_14149,N_13174,N_13731);
nand U14150 (N_14150,N_13459,N_13251);
or U14151 (N_14151,N_13653,N_13538);
and U14152 (N_14152,N_13522,N_13495);
or U14153 (N_14153,N_13223,N_13635);
and U14154 (N_14154,N_13210,N_13358);
nor U14155 (N_14155,N_13464,N_13234);
nand U14156 (N_14156,N_13266,N_13430);
nor U14157 (N_14157,N_13596,N_13472);
or U14158 (N_14158,N_13739,N_13214);
and U14159 (N_14159,N_13332,N_13337);
and U14160 (N_14160,N_13151,N_13289);
or U14161 (N_14161,N_13261,N_13614);
or U14162 (N_14162,N_13388,N_13368);
xor U14163 (N_14163,N_13227,N_13290);
xor U14164 (N_14164,N_13324,N_13696);
and U14165 (N_14165,N_13514,N_13512);
and U14166 (N_14166,N_13356,N_13261);
and U14167 (N_14167,N_13204,N_13512);
nor U14168 (N_14168,N_13666,N_13321);
nor U14169 (N_14169,N_13328,N_13356);
xnor U14170 (N_14170,N_13662,N_13493);
nor U14171 (N_14171,N_13154,N_13157);
or U14172 (N_14172,N_13411,N_13225);
and U14173 (N_14173,N_13256,N_13161);
and U14174 (N_14174,N_13202,N_13196);
nor U14175 (N_14175,N_13452,N_13569);
nor U14176 (N_14176,N_13673,N_13311);
nor U14177 (N_14177,N_13607,N_13268);
nor U14178 (N_14178,N_13461,N_13522);
xor U14179 (N_14179,N_13288,N_13377);
nor U14180 (N_14180,N_13212,N_13184);
nor U14181 (N_14181,N_13465,N_13333);
nor U14182 (N_14182,N_13606,N_13541);
nor U14183 (N_14183,N_13534,N_13436);
xor U14184 (N_14184,N_13416,N_13383);
or U14185 (N_14185,N_13241,N_13518);
nand U14186 (N_14186,N_13467,N_13435);
and U14187 (N_14187,N_13197,N_13630);
or U14188 (N_14188,N_13354,N_13569);
and U14189 (N_14189,N_13735,N_13416);
or U14190 (N_14190,N_13292,N_13713);
xor U14191 (N_14191,N_13692,N_13728);
and U14192 (N_14192,N_13454,N_13421);
or U14193 (N_14193,N_13470,N_13526);
and U14194 (N_14194,N_13469,N_13242);
and U14195 (N_14195,N_13500,N_13703);
or U14196 (N_14196,N_13745,N_13576);
nand U14197 (N_14197,N_13678,N_13246);
or U14198 (N_14198,N_13268,N_13346);
and U14199 (N_14199,N_13487,N_13581);
nand U14200 (N_14200,N_13359,N_13736);
nand U14201 (N_14201,N_13214,N_13580);
nor U14202 (N_14202,N_13283,N_13152);
and U14203 (N_14203,N_13304,N_13514);
or U14204 (N_14204,N_13385,N_13543);
nor U14205 (N_14205,N_13202,N_13313);
xnor U14206 (N_14206,N_13643,N_13228);
nand U14207 (N_14207,N_13316,N_13386);
nand U14208 (N_14208,N_13334,N_13268);
or U14209 (N_14209,N_13268,N_13612);
nand U14210 (N_14210,N_13177,N_13384);
nand U14211 (N_14211,N_13240,N_13197);
nor U14212 (N_14212,N_13307,N_13669);
nand U14213 (N_14213,N_13270,N_13260);
nor U14214 (N_14214,N_13258,N_13674);
nor U14215 (N_14215,N_13525,N_13277);
nand U14216 (N_14216,N_13150,N_13214);
nand U14217 (N_14217,N_13306,N_13714);
and U14218 (N_14218,N_13483,N_13712);
nor U14219 (N_14219,N_13192,N_13655);
nor U14220 (N_14220,N_13219,N_13373);
or U14221 (N_14221,N_13172,N_13646);
or U14222 (N_14222,N_13149,N_13577);
or U14223 (N_14223,N_13368,N_13591);
nand U14224 (N_14224,N_13488,N_13503);
xnor U14225 (N_14225,N_13678,N_13488);
and U14226 (N_14226,N_13270,N_13658);
nor U14227 (N_14227,N_13159,N_13482);
nand U14228 (N_14228,N_13557,N_13644);
nor U14229 (N_14229,N_13145,N_13130);
and U14230 (N_14230,N_13694,N_13561);
nor U14231 (N_14231,N_13541,N_13465);
xnor U14232 (N_14232,N_13519,N_13489);
nor U14233 (N_14233,N_13175,N_13578);
xnor U14234 (N_14234,N_13676,N_13222);
nand U14235 (N_14235,N_13276,N_13615);
nand U14236 (N_14236,N_13396,N_13519);
or U14237 (N_14237,N_13567,N_13195);
and U14238 (N_14238,N_13691,N_13512);
or U14239 (N_14239,N_13623,N_13269);
or U14240 (N_14240,N_13175,N_13144);
or U14241 (N_14241,N_13199,N_13300);
and U14242 (N_14242,N_13444,N_13651);
and U14243 (N_14243,N_13309,N_13501);
nor U14244 (N_14244,N_13394,N_13292);
and U14245 (N_14245,N_13161,N_13436);
xnor U14246 (N_14246,N_13520,N_13227);
and U14247 (N_14247,N_13493,N_13427);
nand U14248 (N_14248,N_13620,N_13253);
nor U14249 (N_14249,N_13547,N_13208);
nand U14250 (N_14250,N_13556,N_13478);
nand U14251 (N_14251,N_13725,N_13747);
or U14252 (N_14252,N_13214,N_13642);
and U14253 (N_14253,N_13607,N_13348);
and U14254 (N_14254,N_13699,N_13705);
or U14255 (N_14255,N_13524,N_13145);
nor U14256 (N_14256,N_13407,N_13713);
or U14257 (N_14257,N_13550,N_13461);
nor U14258 (N_14258,N_13475,N_13629);
xor U14259 (N_14259,N_13615,N_13176);
and U14260 (N_14260,N_13431,N_13653);
and U14261 (N_14261,N_13262,N_13210);
nand U14262 (N_14262,N_13395,N_13540);
nor U14263 (N_14263,N_13300,N_13251);
or U14264 (N_14264,N_13706,N_13415);
xor U14265 (N_14265,N_13448,N_13709);
nor U14266 (N_14266,N_13536,N_13510);
xnor U14267 (N_14267,N_13127,N_13564);
nand U14268 (N_14268,N_13280,N_13290);
xnor U14269 (N_14269,N_13482,N_13495);
xor U14270 (N_14270,N_13398,N_13732);
nand U14271 (N_14271,N_13636,N_13264);
or U14272 (N_14272,N_13234,N_13516);
and U14273 (N_14273,N_13351,N_13217);
and U14274 (N_14274,N_13219,N_13488);
nand U14275 (N_14275,N_13487,N_13445);
nand U14276 (N_14276,N_13558,N_13522);
xnor U14277 (N_14277,N_13660,N_13548);
and U14278 (N_14278,N_13256,N_13672);
or U14279 (N_14279,N_13563,N_13415);
and U14280 (N_14280,N_13675,N_13165);
nor U14281 (N_14281,N_13488,N_13455);
xor U14282 (N_14282,N_13212,N_13319);
or U14283 (N_14283,N_13550,N_13736);
nor U14284 (N_14284,N_13450,N_13555);
and U14285 (N_14285,N_13371,N_13176);
nor U14286 (N_14286,N_13469,N_13544);
nor U14287 (N_14287,N_13423,N_13707);
nand U14288 (N_14288,N_13427,N_13326);
xnor U14289 (N_14289,N_13567,N_13566);
and U14290 (N_14290,N_13169,N_13408);
and U14291 (N_14291,N_13369,N_13636);
xor U14292 (N_14292,N_13320,N_13189);
xor U14293 (N_14293,N_13366,N_13302);
or U14294 (N_14294,N_13734,N_13467);
or U14295 (N_14295,N_13139,N_13556);
or U14296 (N_14296,N_13248,N_13586);
nand U14297 (N_14297,N_13636,N_13284);
nand U14298 (N_14298,N_13155,N_13218);
nor U14299 (N_14299,N_13349,N_13475);
and U14300 (N_14300,N_13714,N_13587);
or U14301 (N_14301,N_13355,N_13236);
nor U14302 (N_14302,N_13410,N_13744);
or U14303 (N_14303,N_13421,N_13379);
and U14304 (N_14304,N_13276,N_13708);
and U14305 (N_14305,N_13232,N_13312);
and U14306 (N_14306,N_13590,N_13498);
and U14307 (N_14307,N_13188,N_13731);
nor U14308 (N_14308,N_13231,N_13175);
xnor U14309 (N_14309,N_13515,N_13429);
and U14310 (N_14310,N_13628,N_13161);
nand U14311 (N_14311,N_13677,N_13156);
xor U14312 (N_14312,N_13657,N_13616);
nor U14313 (N_14313,N_13507,N_13159);
or U14314 (N_14314,N_13570,N_13138);
xor U14315 (N_14315,N_13232,N_13452);
nor U14316 (N_14316,N_13331,N_13281);
and U14317 (N_14317,N_13291,N_13616);
and U14318 (N_14318,N_13667,N_13354);
xnor U14319 (N_14319,N_13326,N_13685);
xnor U14320 (N_14320,N_13457,N_13235);
nor U14321 (N_14321,N_13190,N_13528);
or U14322 (N_14322,N_13537,N_13552);
and U14323 (N_14323,N_13168,N_13174);
or U14324 (N_14324,N_13653,N_13581);
and U14325 (N_14325,N_13211,N_13244);
and U14326 (N_14326,N_13542,N_13424);
and U14327 (N_14327,N_13149,N_13519);
nand U14328 (N_14328,N_13339,N_13528);
nor U14329 (N_14329,N_13678,N_13212);
nand U14330 (N_14330,N_13259,N_13344);
or U14331 (N_14331,N_13444,N_13707);
nor U14332 (N_14332,N_13519,N_13319);
nor U14333 (N_14333,N_13394,N_13356);
xnor U14334 (N_14334,N_13477,N_13365);
or U14335 (N_14335,N_13303,N_13606);
xnor U14336 (N_14336,N_13273,N_13491);
xnor U14337 (N_14337,N_13502,N_13287);
xnor U14338 (N_14338,N_13149,N_13620);
xnor U14339 (N_14339,N_13178,N_13144);
nor U14340 (N_14340,N_13399,N_13335);
nand U14341 (N_14341,N_13580,N_13445);
and U14342 (N_14342,N_13467,N_13243);
xor U14343 (N_14343,N_13215,N_13323);
or U14344 (N_14344,N_13466,N_13243);
nor U14345 (N_14345,N_13729,N_13170);
xnor U14346 (N_14346,N_13281,N_13520);
and U14347 (N_14347,N_13696,N_13482);
nor U14348 (N_14348,N_13592,N_13224);
xor U14349 (N_14349,N_13239,N_13446);
xnor U14350 (N_14350,N_13355,N_13682);
nand U14351 (N_14351,N_13248,N_13495);
nand U14352 (N_14352,N_13405,N_13300);
or U14353 (N_14353,N_13591,N_13380);
nand U14354 (N_14354,N_13440,N_13494);
nor U14355 (N_14355,N_13171,N_13582);
xor U14356 (N_14356,N_13261,N_13176);
nand U14357 (N_14357,N_13441,N_13544);
nor U14358 (N_14358,N_13620,N_13432);
nand U14359 (N_14359,N_13325,N_13467);
or U14360 (N_14360,N_13228,N_13673);
or U14361 (N_14361,N_13713,N_13731);
nand U14362 (N_14362,N_13666,N_13276);
nor U14363 (N_14363,N_13350,N_13579);
nand U14364 (N_14364,N_13530,N_13432);
or U14365 (N_14365,N_13165,N_13378);
nor U14366 (N_14366,N_13358,N_13405);
or U14367 (N_14367,N_13127,N_13178);
or U14368 (N_14368,N_13280,N_13469);
xor U14369 (N_14369,N_13728,N_13444);
or U14370 (N_14370,N_13233,N_13284);
and U14371 (N_14371,N_13192,N_13397);
nand U14372 (N_14372,N_13218,N_13363);
nand U14373 (N_14373,N_13426,N_13340);
xnor U14374 (N_14374,N_13270,N_13585);
and U14375 (N_14375,N_13767,N_14347);
nor U14376 (N_14376,N_14017,N_14030);
xnor U14377 (N_14377,N_14224,N_14229);
nor U14378 (N_14378,N_14210,N_14329);
or U14379 (N_14379,N_13836,N_13868);
nor U14380 (N_14380,N_14273,N_14248);
xnor U14381 (N_14381,N_13828,N_13958);
xnor U14382 (N_14382,N_13804,N_13844);
nor U14383 (N_14383,N_14254,N_13905);
nor U14384 (N_14384,N_14326,N_14269);
or U14385 (N_14385,N_13816,N_13869);
xnor U14386 (N_14386,N_14071,N_13805);
or U14387 (N_14387,N_13842,N_14135);
and U14388 (N_14388,N_14039,N_14008);
xor U14389 (N_14389,N_14000,N_13809);
nand U14390 (N_14390,N_14307,N_13965);
nor U14391 (N_14391,N_13824,N_14213);
and U14392 (N_14392,N_13875,N_14015);
nor U14393 (N_14393,N_14290,N_14049);
and U14394 (N_14394,N_14227,N_14340);
and U14395 (N_14395,N_14029,N_14374);
xor U14396 (N_14396,N_13991,N_13952);
or U14397 (N_14397,N_13838,N_14116);
or U14398 (N_14398,N_13871,N_13788);
nor U14399 (N_14399,N_14137,N_13873);
or U14400 (N_14400,N_14342,N_13832);
and U14401 (N_14401,N_13922,N_14369);
nor U14402 (N_14402,N_14244,N_13887);
or U14403 (N_14403,N_14159,N_14160);
nor U14404 (N_14404,N_13889,N_14281);
nor U14405 (N_14405,N_14218,N_14051);
and U14406 (N_14406,N_14074,N_13821);
nor U14407 (N_14407,N_13776,N_14279);
nand U14408 (N_14408,N_13961,N_14344);
nand U14409 (N_14409,N_13813,N_13798);
and U14410 (N_14410,N_13935,N_14099);
or U14411 (N_14411,N_14180,N_14197);
or U14412 (N_14412,N_14367,N_14038);
or U14413 (N_14413,N_13855,N_14310);
nand U14414 (N_14414,N_14297,N_14291);
nand U14415 (N_14415,N_14028,N_13764);
nor U14416 (N_14416,N_14263,N_13786);
or U14417 (N_14417,N_14276,N_14035);
nor U14418 (N_14418,N_14102,N_13907);
or U14419 (N_14419,N_14370,N_14122);
and U14420 (N_14420,N_13769,N_13973);
or U14421 (N_14421,N_14270,N_14311);
or U14422 (N_14422,N_14048,N_14104);
xnor U14423 (N_14423,N_14126,N_14255);
and U14424 (N_14424,N_14082,N_13941);
or U14425 (N_14425,N_14075,N_13854);
and U14426 (N_14426,N_14253,N_14094);
nor U14427 (N_14427,N_13981,N_14088);
and U14428 (N_14428,N_14241,N_14046);
nand U14429 (N_14429,N_14106,N_14302);
nand U14430 (N_14430,N_14338,N_14353);
or U14431 (N_14431,N_14292,N_13954);
or U14432 (N_14432,N_13807,N_14019);
or U14433 (N_14433,N_14264,N_14172);
or U14434 (N_14434,N_13841,N_14078);
and U14435 (N_14435,N_14271,N_13818);
nor U14436 (N_14436,N_14181,N_14275);
or U14437 (N_14437,N_13926,N_13983);
and U14438 (N_14438,N_14349,N_14167);
nand U14439 (N_14439,N_14298,N_14343);
or U14440 (N_14440,N_14259,N_14260);
and U14441 (N_14441,N_14330,N_14124);
or U14442 (N_14442,N_14143,N_13874);
nand U14443 (N_14443,N_14251,N_13938);
nand U14444 (N_14444,N_13845,N_14056);
nor U14445 (N_14445,N_14186,N_14339);
nor U14446 (N_14446,N_14320,N_14242);
or U14447 (N_14447,N_14138,N_14054);
and U14448 (N_14448,N_13876,N_13860);
or U14449 (N_14449,N_14042,N_14262);
nor U14450 (N_14450,N_14333,N_14199);
or U14451 (N_14451,N_13903,N_14288);
nor U14452 (N_14452,N_13750,N_13772);
or U14453 (N_14453,N_13985,N_13886);
and U14454 (N_14454,N_13997,N_14196);
nand U14455 (N_14455,N_14324,N_13768);
nand U14456 (N_14456,N_13775,N_13762);
or U14457 (N_14457,N_14007,N_14247);
nor U14458 (N_14458,N_13946,N_14204);
xnor U14459 (N_14459,N_14141,N_14058);
and U14460 (N_14460,N_13917,N_14045);
nand U14461 (N_14461,N_13976,N_14146);
or U14462 (N_14462,N_14136,N_13923);
and U14463 (N_14463,N_13864,N_14068);
or U14464 (N_14464,N_14132,N_13911);
or U14465 (N_14465,N_14328,N_14246);
nor U14466 (N_14466,N_13759,N_13900);
xnor U14467 (N_14467,N_13906,N_13819);
xnor U14468 (N_14468,N_13758,N_13882);
nor U14469 (N_14469,N_14257,N_13793);
xnor U14470 (N_14470,N_14059,N_14177);
and U14471 (N_14471,N_14185,N_14002);
xnor U14472 (N_14472,N_14345,N_14113);
xnor U14473 (N_14473,N_14031,N_14108);
xor U14474 (N_14474,N_13843,N_13833);
nand U14475 (N_14475,N_14100,N_14289);
nor U14476 (N_14476,N_14103,N_13990);
xor U14477 (N_14477,N_13970,N_13972);
nand U14478 (N_14478,N_14063,N_14064);
nand U14479 (N_14479,N_13839,N_13802);
and U14480 (N_14480,N_13901,N_14119);
xnor U14481 (N_14481,N_13784,N_14212);
nor U14482 (N_14482,N_13763,N_14336);
and U14483 (N_14483,N_14304,N_13834);
or U14484 (N_14484,N_14243,N_13924);
nor U14485 (N_14485,N_14157,N_13909);
or U14486 (N_14486,N_13808,N_14107);
and U14487 (N_14487,N_14156,N_13996);
or U14488 (N_14488,N_13969,N_14284);
nor U14489 (N_14489,N_14134,N_13773);
xor U14490 (N_14490,N_14325,N_13879);
xnor U14491 (N_14491,N_14024,N_14140);
nand U14492 (N_14492,N_13994,N_14013);
or U14493 (N_14493,N_13890,N_13934);
nor U14494 (N_14494,N_13937,N_13947);
nor U14495 (N_14495,N_13920,N_14006);
nor U14496 (N_14496,N_13799,N_14076);
nor U14497 (N_14497,N_13811,N_13885);
and U14498 (N_14498,N_13929,N_14321);
nand U14499 (N_14499,N_14331,N_14170);
xnor U14500 (N_14500,N_13883,N_13916);
and U14501 (N_14501,N_13930,N_13984);
and U14502 (N_14502,N_14026,N_13992);
nand U14503 (N_14503,N_14223,N_14267);
nor U14504 (N_14504,N_14111,N_14312);
nor U14505 (N_14505,N_14295,N_14182);
and U14506 (N_14506,N_14372,N_14368);
nand U14507 (N_14507,N_13790,N_14004);
nor U14508 (N_14508,N_13778,N_13982);
nor U14509 (N_14509,N_14183,N_14043);
nor U14510 (N_14510,N_13971,N_14014);
or U14511 (N_14511,N_14057,N_14208);
and U14512 (N_14512,N_14256,N_14358);
nand U14513 (N_14513,N_13943,N_13756);
and U14514 (N_14514,N_14309,N_14294);
nand U14515 (N_14515,N_13777,N_14365);
nor U14516 (N_14516,N_14114,N_14123);
and U14517 (N_14517,N_13977,N_14323);
nor U14518 (N_14518,N_14091,N_14316);
nand U14519 (N_14519,N_14190,N_13761);
nand U14520 (N_14520,N_13921,N_14286);
or U14521 (N_14521,N_14205,N_14098);
nor U14522 (N_14522,N_14125,N_13939);
nor U14523 (N_14523,N_14322,N_13978);
nand U14524 (N_14524,N_14303,N_14228);
or U14525 (N_14525,N_14142,N_14209);
nor U14526 (N_14526,N_13851,N_14360);
nor U14527 (N_14527,N_13820,N_13863);
nor U14528 (N_14528,N_14211,N_13770);
nor U14529 (N_14529,N_14221,N_14010);
or U14530 (N_14530,N_14198,N_14171);
or U14531 (N_14531,N_14089,N_13856);
xnor U14532 (N_14532,N_13914,N_13953);
nand U14533 (N_14533,N_14168,N_14266);
nor U14534 (N_14534,N_13794,N_14249);
xnor U14535 (N_14535,N_13754,N_14052);
nor U14536 (N_14536,N_13835,N_13988);
or U14537 (N_14537,N_13897,N_13968);
and U14538 (N_14538,N_14109,N_14261);
nor U14539 (N_14539,N_14173,N_14258);
xnor U14540 (N_14540,N_14151,N_13960);
nor U14541 (N_14541,N_13959,N_14022);
xor U14542 (N_14542,N_14189,N_13862);
and U14543 (N_14543,N_13827,N_13918);
and U14544 (N_14544,N_14315,N_13803);
nand U14545 (N_14545,N_14359,N_14129);
and U14546 (N_14546,N_14152,N_13814);
and U14547 (N_14547,N_13899,N_14037);
and U14548 (N_14548,N_14373,N_14216);
or U14549 (N_14549,N_14222,N_14131);
nand U14550 (N_14550,N_13936,N_14233);
and U14551 (N_14551,N_14194,N_14300);
nand U14552 (N_14552,N_14225,N_14005);
or U14553 (N_14553,N_14240,N_14206);
nor U14554 (N_14554,N_14293,N_14350);
and U14555 (N_14555,N_13894,N_14097);
xnor U14556 (N_14556,N_14053,N_13751);
nand U14557 (N_14557,N_13755,N_14127);
and U14558 (N_14558,N_14341,N_14238);
xor U14559 (N_14559,N_13986,N_13998);
or U14560 (N_14560,N_13904,N_13902);
nor U14561 (N_14561,N_13915,N_13849);
xnor U14562 (N_14562,N_14226,N_14308);
xnor U14563 (N_14563,N_14093,N_14150);
or U14564 (N_14564,N_14237,N_14067);
nor U14565 (N_14565,N_14083,N_14207);
nand U14566 (N_14566,N_14192,N_14154);
or U14567 (N_14567,N_14317,N_14047);
or U14568 (N_14568,N_13753,N_14214);
nor U14569 (N_14569,N_13928,N_14086);
nor U14570 (N_14570,N_13962,N_13781);
nand U14571 (N_14571,N_13933,N_13927);
and U14572 (N_14572,N_14062,N_13865);
xnor U14573 (N_14573,N_13944,N_13846);
and U14574 (N_14574,N_13980,N_14175);
nor U14575 (N_14575,N_14334,N_13910);
and U14576 (N_14576,N_13795,N_14003);
and U14577 (N_14577,N_13955,N_13791);
or U14578 (N_14578,N_14366,N_13787);
xnor U14579 (N_14579,N_14018,N_14230);
and U14580 (N_14580,N_14169,N_14327);
nor U14581 (N_14581,N_13912,N_14027);
nor U14582 (N_14582,N_14069,N_13806);
nand U14583 (N_14583,N_14278,N_14040);
or U14584 (N_14584,N_14299,N_14332);
nor U14585 (N_14585,N_13950,N_13940);
nand U14586 (N_14586,N_14318,N_13895);
and U14587 (N_14587,N_14050,N_13999);
or U14588 (N_14588,N_14188,N_14176);
and U14589 (N_14589,N_14200,N_14371);
and U14590 (N_14590,N_13866,N_13847);
nand U14591 (N_14591,N_13771,N_14105);
nand U14592 (N_14592,N_14001,N_13780);
and U14593 (N_14593,N_13867,N_13812);
nor U14594 (N_14594,N_13757,N_14118);
xor U14595 (N_14595,N_13957,N_14084);
nor U14596 (N_14596,N_13779,N_13979);
nor U14597 (N_14597,N_13989,N_13966);
or U14598 (N_14598,N_13880,N_14357);
xor U14599 (N_14599,N_13857,N_13942);
or U14600 (N_14600,N_13797,N_14162);
or U14601 (N_14601,N_14265,N_13774);
nand U14602 (N_14602,N_14346,N_14348);
nand U14603 (N_14603,N_14147,N_14215);
nor U14604 (N_14604,N_14178,N_13949);
xor U14605 (N_14605,N_14121,N_14232);
and U14606 (N_14606,N_14077,N_14025);
nand U14607 (N_14607,N_13766,N_14239);
xor U14608 (N_14608,N_14335,N_14148);
or U14609 (N_14609,N_14305,N_14250);
or U14610 (N_14610,N_13858,N_14081);
nor U14611 (N_14611,N_14352,N_14155);
and U14612 (N_14612,N_14234,N_13826);
nor U14613 (N_14613,N_13877,N_14179);
nor U14614 (N_14614,N_14220,N_13878);
or U14615 (N_14615,N_13898,N_14033);
nor U14616 (N_14616,N_13796,N_13987);
nor U14617 (N_14617,N_13872,N_14364);
or U14618 (N_14618,N_13792,N_13861);
xnor U14619 (N_14619,N_13891,N_14306);
nand U14620 (N_14620,N_14149,N_14166);
xor U14621 (N_14621,N_13932,N_14319);
nor U14622 (N_14622,N_13785,N_14079);
nand U14623 (N_14623,N_14296,N_14201);
or U14624 (N_14624,N_14036,N_14041);
nor U14625 (N_14625,N_14301,N_13810);
xor U14626 (N_14626,N_14272,N_14268);
xor U14627 (N_14627,N_13850,N_13964);
nor U14628 (N_14628,N_14161,N_14011);
nand U14629 (N_14629,N_13888,N_14021);
nor U14630 (N_14630,N_14144,N_13760);
nor U14631 (N_14631,N_14202,N_14203);
nand U14632 (N_14632,N_14184,N_13801);
xnor U14633 (N_14633,N_13765,N_14095);
nor U14634 (N_14634,N_14245,N_13995);
nand U14635 (N_14635,N_14066,N_14139);
nand U14636 (N_14636,N_13825,N_13956);
nor U14637 (N_14637,N_14195,N_13919);
and U14638 (N_14638,N_14092,N_14044);
xor U14639 (N_14639,N_13783,N_13945);
xnor U14640 (N_14640,N_13829,N_13967);
or U14641 (N_14641,N_14080,N_13951);
and U14642 (N_14642,N_14012,N_14287);
or U14643 (N_14643,N_14217,N_13974);
nand U14644 (N_14644,N_14055,N_13913);
and U14645 (N_14645,N_14337,N_14280);
and U14646 (N_14646,N_14285,N_14158);
xnor U14647 (N_14647,N_13840,N_14072);
xor U14648 (N_14648,N_14016,N_14362);
nand U14649 (N_14649,N_14023,N_14115);
nor U14650 (N_14650,N_13848,N_14085);
or U14651 (N_14651,N_14060,N_14073);
and U14652 (N_14652,N_13789,N_14165);
and U14653 (N_14653,N_14087,N_14351);
nand U14654 (N_14654,N_13908,N_14363);
and U14655 (N_14655,N_13852,N_13815);
or U14656 (N_14656,N_14130,N_14032);
and U14657 (N_14657,N_13837,N_13822);
nand U14658 (N_14658,N_14193,N_13884);
or U14659 (N_14659,N_14219,N_14117);
nand U14660 (N_14660,N_13892,N_14235);
nor U14661 (N_14661,N_14282,N_14128);
and U14662 (N_14662,N_13752,N_13870);
nand U14663 (N_14663,N_14145,N_14252);
xnor U14664 (N_14664,N_13853,N_13993);
nor U14665 (N_14665,N_14090,N_13896);
nor U14666 (N_14666,N_13800,N_14314);
xor U14667 (N_14667,N_14356,N_13817);
and U14668 (N_14668,N_14355,N_13931);
nand U14669 (N_14669,N_14153,N_14133);
nor U14670 (N_14670,N_14313,N_14163);
nand U14671 (N_14671,N_14070,N_13823);
nand U14672 (N_14672,N_14361,N_14020);
xor U14673 (N_14673,N_14096,N_13782);
nand U14674 (N_14674,N_14187,N_14174);
and U14675 (N_14675,N_14101,N_13830);
and U14676 (N_14676,N_14191,N_13859);
or U14677 (N_14677,N_14034,N_14112);
nor U14678 (N_14678,N_13975,N_14283);
xnor U14679 (N_14679,N_14277,N_14061);
or U14680 (N_14680,N_13831,N_13948);
nand U14681 (N_14681,N_14120,N_13925);
nor U14682 (N_14682,N_13963,N_14236);
xnor U14683 (N_14683,N_14164,N_13893);
nand U14684 (N_14684,N_14354,N_14274);
nor U14685 (N_14685,N_14231,N_13881);
nor U14686 (N_14686,N_14065,N_14009);
nor U14687 (N_14687,N_14110,N_13861);
or U14688 (N_14688,N_14192,N_14112);
nor U14689 (N_14689,N_13972,N_14367);
nand U14690 (N_14690,N_14217,N_13973);
nand U14691 (N_14691,N_13965,N_14304);
and U14692 (N_14692,N_14365,N_14098);
and U14693 (N_14693,N_13825,N_14337);
nor U14694 (N_14694,N_13796,N_14368);
nor U14695 (N_14695,N_13757,N_13996);
nand U14696 (N_14696,N_13859,N_14283);
nor U14697 (N_14697,N_14133,N_14236);
and U14698 (N_14698,N_14298,N_14265);
or U14699 (N_14699,N_14205,N_14115);
xor U14700 (N_14700,N_13771,N_14374);
nand U14701 (N_14701,N_13796,N_14270);
nand U14702 (N_14702,N_13990,N_14211);
or U14703 (N_14703,N_14234,N_13852);
nor U14704 (N_14704,N_13754,N_13931);
nand U14705 (N_14705,N_13831,N_13988);
nor U14706 (N_14706,N_14044,N_14127);
xor U14707 (N_14707,N_14047,N_14280);
xnor U14708 (N_14708,N_14234,N_14016);
xor U14709 (N_14709,N_14322,N_14350);
nor U14710 (N_14710,N_14087,N_14305);
xor U14711 (N_14711,N_14158,N_13941);
xnor U14712 (N_14712,N_13750,N_13909);
nor U14713 (N_14713,N_13998,N_14095);
or U14714 (N_14714,N_14114,N_14275);
nand U14715 (N_14715,N_14271,N_13805);
and U14716 (N_14716,N_13882,N_14132);
nand U14717 (N_14717,N_14006,N_13878);
nor U14718 (N_14718,N_14225,N_14125);
xor U14719 (N_14719,N_14086,N_13967);
nand U14720 (N_14720,N_13923,N_14341);
xor U14721 (N_14721,N_13913,N_14089);
nand U14722 (N_14722,N_13805,N_13924);
nand U14723 (N_14723,N_14364,N_14127);
and U14724 (N_14724,N_13908,N_13865);
and U14725 (N_14725,N_14235,N_14066);
and U14726 (N_14726,N_13998,N_14336);
xnor U14727 (N_14727,N_13780,N_13783);
nand U14728 (N_14728,N_14230,N_13895);
xor U14729 (N_14729,N_14324,N_14127);
xor U14730 (N_14730,N_14259,N_14328);
nor U14731 (N_14731,N_14122,N_13769);
xor U14732 (N_14732,N_14255,N_14004);
or U14733 (N_14733,N_13804,N_14301);
and U14734 (N_14734,N_13997,N_14362);
nor U14735 (N_14735,N_14138,N_14044);
nor U14736 (N_14736,N_14184,N_14269);
nand U14737 (N_14737,N_14353,N_14266);
and U14738 (N_14738,N_13786,N_13775);
nand U14739 (N_14739,N_13815,N_13960);
nor U14740 (N_14740,N_13846,N_14033);
xor U14741 (N_14741,N_14304,N_14043);
and U14742 (N_14742,N_13766,N_14353);
nor U14743 (N_14743,N_14089,N_13993);
nand U14744 (N_14744,N_14242,N_14192);
or U14745 (N_14745,N_13938,N_14016);
nor U14746 (N_14746,N_14050,N_14059);
or U14747 (N_14747,N_13889,N_14186);
and U14748 (N_14748,N_14199,N_13911);
or U14749 (N_14749,N_14303,N_13901);
nand U14750 (N_14750,N_13817,N_14199);
nor U14751 (N_14751,N_13998,N_14263);
nor U14752 (N_14752,N_14268,N_14298);
nor U14753 (N_14753,N_14023,N_14270);
and U14754 (N_14754,N_14043,N_14245);
and U14755 (N_14755,N_14028,N_14048);
nor U14756 (N_14756,N_14154,N_14073);
and U14757 (N_14757,N_14178,N_13775);
nor U14758 (N_14758,N_13886,N_14219);
xor U14759 (N_14759,N_14080,N_14146);
nor U14760 (N_14760,N_14102,N_13801);
and U14761 (N_14761,N_13996,N_14033);
and U14762 (N_14762,N_14251,N_13800);
and U14763 (N_14763,N_14205,N_14211);
xnor U14764 (N_14764,N_14154,N_13891);
nand U14765 (N_14765,N_14280,N_13906);
xor U14766 (N_14766,N_14165,N_13829);
or U14767 (N_14767,N_14053,N_14159);
nand U14768 (N_14768,N_14245,N_14089);
nand U14769 (N_14769,N_14218,N_13934);
nand U14770 (N_14770,N_14014,N_13889);
nor U14771 (N_14771,N_13899,N_13787);
or U14772 (N_14772,N_14160,N_13973);
or U14773 (N_14773,N_14139,N_13878);
nor U14774 (N_14774,N_14189,N_13987);
nor U14775 (N_14775,N_14221,N_13906);
or U14776 (N_14776,N_14085,N_14086);
and U14777 (N_14777,N_14149,N_13767);
and U14778 (N_14778,N_14195,N_13835);
nand U14779 (N_14779,N_13902,N_14115);
xor U14780 (N_14780,N_13884,N_13860);
or U14781 (N_14781,N_14189,N_14268);
xnor U14782 (N_14782,N_13751,N_14339);
or U14783 (N_14783,N_13808,N_14312);
or U14784 (N_14784,N_14249,N_14369);
or U14785 (N_14785,N_14010,N_14277);
or U14786 (N_14786,N_13869,N_14126);
nand U14787 (N_14787,N_13814,N_14226);
nor U14788 (N_14788,N_14077,N_14294);
nor U14789 (N_14789,N_14065,N_13868);
xnor U14790 (N_14790,N_13875,N_14146);
xor U14791 (N_14791,N_14336,N_14355);
nand U14792 (N_14792,N_14247,N_14124);
or U14793 (N_14793,N_13790,N_14355);
nand U14794 (N_14794,N_14112,N_14141);
nand U14795 (N_14795,N_13910,N_13999);
nor U14796 (N_14796,N_14043,N_13934);
nor U14797 (N_14797,N_14364,N_14165);
nand U14798 (N_14798,N_13880,N_14035);
nand U14799 (N_14799,N_14007,N_13758);
and U14800 (N_14800,N_14254,N_14308);
or U14801 (N_14801,N_13880,N_14179);
or U14802 (N_14802,N_13968,N_14289);
nor U14803 (N_14803,N_14072,N_14020);
or U14804 (N_14804,N_14220,N_14222);
nor U14805 (N_14805,N_13798,N_14303);
nor U14806 (N_14806,N_13869,N_14018);
and U14807 (N_14807,N_13890,N_14136);
nand U14808 (N_14808,N_13910,N_14026);
nand U14809 (N_14809,N_14249,N_13958);
or U14810 (N_14810,N_14101,N_14100);
nand U14811 (N_14811,N_14015,N_13823);
xnor U14812 (N_14812,N_13849,N_14326);
nand U14813 (N_14813,N_13928,N_14225);
nor U14814 (N_14814,N_14330,N_14132);
and U14815 (N_14815,N_14081,N_14031);
or U14816 (N_14816,N_14087,N_14335);
xor U14817 (N_14817,N_13988,N_13885);
and U14818 (N_14818,N_14178,N_14177);
and U14819 (N_14819,N_13939,N_14360);
and U14820 (N_14820,N_13755,N_13849);
xor U14821 (N_14821,N_13828,N_14117);
and U14822 (N_14822,N_14196,N_14002);
or U14823 (N_14823,N_13927,N_14117);
nand U14824 (N_14824,N_14252,N_13826);
or U14825 (N_14825,N_14035,N_13953);
nor U14826 (N_14826,N_14027,N_13926);
nor U14827 (N_14827,N_14178,N_13804);
nand U14828 (N_14828,N_14201,N_14171);
nand U14829 (N_14829,N_14215,N_13834);
nor U14830 (N_14830,N_14026,N_13956);
nand U14831 (N_14831,N_14294,N_14183);
and U14832 (N_14832,N_14042,N_14200);
nor U14833 (N_14833,N_13974,N_14179);
or U14834 (N_14834,N_14133,N_14105);
nor U14835 (N_14835,N_14327,N_13795);
and U14836 (N_14836,N_13971,N_13785);
xor U14837 (N_14837,N_13831,N_14022);
and U14838 (N_14838,N_13801,N_14071);
xor U14839 (N_14839,N_14011,N_14019);
xor U14840 (N_14840,N_13911,N_13928);
nor U14841 (N_14841,N_13895,N_14103);
xor U14842 (N_14842,N_14098,N_14008);
nand U14843 (N_14843,N_13899,N_13790);
and U14844 (N_14844,N_13867,N_14322);
xnor U14845 (N_14845,N_14066,N_14330);
xnor U14846 (N_14846,N_14317,N_14044);
xnor U14847 (N_14847,N_14308,N_13915);
nand U14848 (N_14848,N_14284,N_13753);
and U14849 (N_14849,N_14076,N_14308);
or U14850 (N_14850,N_13951,N_13994);
xnor U14851 (N_14851,N_14274,N_13991);
nor U14852 (N_14852,N_14045,N_14009);
or U14853 (N_14853,N_14007,N_14351);
xor U14854 (N_14854,N_13796,N_13988);
xnor U14855 (N_14855,N_14183,N_14058);
nor U14856 (N_14856,N_14286,N_14169);
or U14857 (N_14857,N_13991,N_14155);
or U14858 (N_14858,N_14048,N_14354);
nor U14859 (N_14859,N_14191,N_14054);
nor U14860 (N_14860,N_14354,N_14049);
and U14861 (N_14861,N_13900,N_14149);
and U14862 (N_14862,N_14010,N_13791);
or U14863 (N_14863,N_14192,N_14161);
or U14864 (N_14864,N_14157,N_14096);
and U14865 (N_14865,N_13835,N_14336);
nand U14866 (N_14866,N_14102,N_14288);
nand U14867 (N_14867,N_14044,N_14013);
nand U14868 (N_14868,N_13921,N_13977);
nand U14869 (N_14869,N_14292,N_13764);
xor U14870 (N_14870,N_14144,N_14351);
or U14871 (N_14871,N_13977,N_14032);
or U14872 (N_14872,N_14118,N_13974);
xor U14873 (N_14873,N_14185,N_14253);
xor U14874 (N_14874,N_14326,N_14225);
xnor U14875 (N_14875,N_14322,N_13779);
xor U14876 (N_14876,N_14269,N_13833);
xor U14877 (N_14877,N_14043,N_14339);
nand U14878 (N_14878,N_13777,N_14291);
xnor U14879 (N_14879,N_13924,N_13923);
nor U14880 (N_14880,N_14119,N_14164);
nor U14881 (N_14881,N_14146,N_13780);
nand U14882 (N_14882,N_14294,N_14084);
and U14883 (N_14883,N_13802,N_14236);
nor U14884 (N_14884,N_14029,N_14138);
and U14885 (N_14885,N_13862,N_13786);
and U14886 (N_14886,N_14019,N_14169);
nor U14887 (N_14887,N_13785,N_13964);
xnor U14888 (N_14888,N_14175,N_13893);
or U14889 (N_14889,N_14349,N_14191);
and U14890 (N_14890,N_14332,N_13888);
and U14891 (N_14891,N_14235,N_14028);
and U14892 (N_14892,N_14040,N_14358);
or U14893 (N_14893,N_14045,N_13784);
and U14894 (N_14894,N_13981,N_14101);
xor U14895 (N_14895,N_13771,N_14154);
xor U14896 (N_14896,N_14092,N_14122);
xnor U14897 (N_14897,N_13899,N_14335);
nand U14898 (N_14898,N_13812,N_14210);
nand U14899 (N_14899,N_14110,N_14211);
or U14900 (N_14900,N_14059,N_14280);
or U14901 (N_14901,N_13992,N_14230);
and U14902 (N_14902,N_14165,N_14356);
nand U14903 (N_14903,N_14032,N_14038);
or U14904 (N_14904,N_13895,N_13821);
nor U14905 (N_14905,N_14114,N_14314);
xnor U14906 (N_14906,N_13863,N_14177);
nor U14907 (N_14907,N_14105,N_14172);
and U14908 (N_14908,N_14076,N_13894);
or U14909 (N_14909,N_13881,N_14125);
nor U14910 (N_14910,N_14188,N_13831);
and U14911 (N_14911,N_14337,N_13760);
nor U14912 (N_14912,N_14080,N_13955);
and U14913 (N_14913,N_14280,N_14035);
nand U14914 (N_14914,N_14296,N_14129);
and U14915 (N_14915,N_14106,N_14295);
and U14916 (N_14916,N_14222,N_13790);
nand U14917 (N_14917,N_14070,N_14002);
or U14918 (N_14918,N_14298,N_13986);
xnor U14919 (N_14919,N_14272,N_14093);
xnor U14920 (N_14920,N_13881,N_13790);
and U14921 (N_14921,N_14353,N_13785);
and U14922 (N_14922,N_14264,N_14306);
xor U14923 (N_14923,N_14129,N_13836);
and U14924 (N_14924,N_13877,N_13789);
and U14925 (N_14925,N_14233,N_13827);
nand U14926 (N_14926,N_14236,N_14330);
nand U14927 (N_14927,N_13918,N_13932);
xor U14928 (N_14928,N_13817,N_13840);
nand U14929 (N_14929,N_14175,N_14181);
or U14930 (N_14930,N_13809,N_14094);
nor U14931 (N_14931,N_13996,N_14280);
nand U14932 (N_14932,N_13953,N_14138);
or U14933 (N_14933,N_14323,N_14069);
xnor U14934 (N_14934,N_13765,N_14311);
and U14935 (N_14935,N_14137,N_14301);
nand U14936 (N_14936,N_14010,N_14170);
and U14937 (N_14937,N_14373,N_14168);
nor U14938 (N_14938,N_13845,N_13956);
xnor U14939 (N_14939,N_13836,N_13801);
nand U14940 (N_14940,N_14016,N_14257);
nand U14941 (N_14941,N_14268,N_14256);
xor U14942 (N_14942,N_14250,N_13849);
nor U14943 (N_14943,N_14127,N_14085);
nor U14944 (N_14944,N_13827,N_14138);
nor U14945 (N_14945,N_13823,N_13802);
or U14946 (N_14946,N_14235,N_13799);
and U14947 (N_14947,N_14102,N_14099);
nor U14948 (N_14948,N_14196,N_14303);
and U14949 (N_14949,N_14101,N_13822);
and U14950 (N_14950,N_14211,N_14193);
xnor U14951 (N_14951,N_13874,N_14104);
xor U14952 (N_14952,N_13944,N_14225);
nand U14953 (N_14953,N_14209,N_14201);
xnor U14954 (N_14954,N_13812,N_14156);
or U14955 (N_14955,N_14328,N_14275);
xnor U14956 (N_14956,N_14229,N_14215);
nor U14957 (N_14957,N_13902,N_14190);
or U14958 (N_14958,N_13800,N_14348);
nand U14959 (N_14959,N_14146,N_13909);
nand U14960 (N_14960,N_14117,N_14222);
nor U14961 (N_14961,N_13977,N_14060);
xor U14962 (N_14962,N_14221,N_13982);
or U14963 (N_14963,N_14183,N_14261);
xnor U14964 (N_14964,N_13840,N_14089);
nand U14965 (N_14965,N_13899,N_14248);
and U14966 (N_14966,N_14371,N_14185);
or U14967 (N_14967,N_14247,N_13906);
or U14968 (N_14968,N_14195,N_13766);
and U14969 (N_14969,N_13827,N_14132);
or U14970 (N_14970,N_14246,N_14250);
nor U14971 (N_14971,N_13804,N_14058);
or U14972 (N_14972,N_14134,N_13923);
nor U14973 (N_14973,N_13938,N_14106);
or U14974 (N_14974,N_13753,N_13820);
nand U14975 (N_14975,N_13829,N_13777);
nand U14976 (N_14976,N_14370,N_14247);
xnor U14977 (N_14977,N_13918,N_13831);
or U14978 (N_14978,N_13950,N_14225);
and U14979 (N_14979,N_14236,N_14282);
nand U14980 (N_14980,N_14169,N_14349);
xor U14981 (N_14981,N_14166,N_14023);
nand U14982 (N_14982,N_14308,N_14056);
or U14983 (N_14983,N_13803,N_13967);
nand U14984 (N_14984,N_13948,N_13812);
and U14985 (N_14985,N_13812,N_13834);
nand U14986 (N_14986,N_14183,N_13953);
or U14987 (N_14987,N_14355,N_13876);
nor U14988 (N_14988,N_14221,N_14119);
or U14989 (N_14989,N_14198,N_14141);
and U14990 (N_14990,N_14302,N_13848);
nor U14991 (N_14991,N_14097,N_13915);
and U14992 (N_14992,N_14085,N_14247);
nor U14993 (N_14993,N_13974,N_14258);
nor U14994 (N_14994,N_14207,N_13930);
nand U14995 (N_14995,N_13966,N_13847);
or U14996 (N_14996,N_14029,N_13849);
or U14997 (N_14997,N_13825,N_14010);
nor U14998 (N_14998,N_14033,N_14274);
nand U14999 (N_14999,N_14103,N_14354);
and U15000 (N_15000,N_14827,N_14579);
or U15001 (N_15001,N_14677,N_14481);
xor U15002 (N_15002,N_14713,N_14486);
or U15003 (N_15003,N_14728,N_14989);
xnor U15004 (N_15004,N_14392,N_14779);
xnor U15005 (N_15005,N_14907,N_14516);
nor U15006 (N_15006,N_14709,N_14658);
nand U15007 (N_15007,N_14806,N_14882);
nand U15008 (N_15008,N_14884,N_14825);
nand U15009 (N_15009,N_14740,N_14404);
nor U15010 (N_15010,N_14777,N_14894);
and U15011 (N_15011,N_14477,N_14844);
or U15012 (N_15012,N_14459,N_14536);
and U15013 (N_15013,N_14970,N_14465);
nand U15014 (N_15014,N_14749,N_14457);
nor U15015 (N_15015,N_14968,N_14976);
and U15016 (N_15016,N_14873,N_14429);
and U15017 (N_15017,N_14794,N_14904);
xor U15018 (N_15018,N_14456,N_14801);
or U15019 (N_15019,N_14542,N_14415);
nand U15020 (N_15020,N_14909,N_14550);
nor U15021 (N_15021,N_14831,N_14697);
xor U15022 (N_15022,N_14756,N_14377);
nand U15023 (N_15023,N_14791,N_14863);
nand U15024 (N_15024,N_14645,N_14802);
nand U15025 (N_15025,N_14770,N_14594);
xor U15026 (N_15026,N_14534,N_14785);
and U15027 (N_15027,N_14981,N_14855);
and U15028 (N_15028,N_14955,N_14530);
xnor U15029 (N_15029,N_14793,N_14500);
or U15030 (N_15030,N_14620,N_14463);
and U15031 (N_15031,N_14730,N_14551);
nand U15032 (N_15032,N_14667,N_14553);
nand U15033 (N_15033,N_14973,N_14621);
nor U15034 (N_15034,N_14914,N_14910);
nor U15035 (N_15035,N_14450,N_14480);
nor U15036 (N_15036,N_14874,N_14478);
nand U15037 (N_15037,N_14715,N_14765);
nor U15038 (N_15038,N_14915,N_14647);
and U15039 (N_15039,N_14518,N_14591);
nand U15040 (N_15040,N_14637,N_14517);
nand U15041 (N_15041,N_14528,N_14615);
nand U15042 (N_15042,N_14771,N_14575);
nor U15043 (N_15043,N_14431,N_14501);
and U15044 (N_15044,N_14397,N_14495);
and U15045 (N_15045,N_14767,N_14502);
or U15046 (N_15046,N_14418,N_14674);
and U15047 (N_15047,N_14755,N_14818);
nor U15048 (N_15048,N_14710,N_14650);
or U15049 (N_15049,N_14387,N_14706);
and U15050 (N_15050,N_14483,N_14969);
or U15051 (N_15051,N_14736,N_14399);
or U15052 (N_15052,N_14752,N_14526);
nor U15053 (N_15053,N_14813,N_14744);
nor U15054 (N_15054,N_14971,N_14963);
or U15055 (N_15055,N_14379,N_14659);
xnor U15056 (N_15056,N_14430,N_14701);
and U15057 (N_15057,N_14389,N_14543);
nor U15058 (N_15058,N_14656,N_14671);
and U15059 (N_15059,N_14673,N_14610);
nor U15060 (N_15060,N_14883,N_14845);
nand U15061 (N_15061,N_14695,N_14394);
nor U15062 (N_15062,N_14898,N_14563);
nand U15063 (N_15063,N_14405,N_14408);
nand U15064 (N_15064,N_14796,N_14690);
or U15065 (N_15065,N_14643,N_14789);
or U15066 (N_15066,N_14733,N_14577);
or U15067 (N_15067,N_14631,N_14686);
or U15068 (N_15068,N_14675,N_14788);
xor U15069 (N_15069,N_14750,N_14447);
and U15070 (N_15070,N_14416,N_14716);
and U15071 (N_15071,N_14832,N_14376);
nor U15072 (N_15072,N_14861,N_14602);
xnor U15073 (N_15073,N_14584,N_14539);
xnor U15074 (N_15074,N_14913,N_14614);
and U15075 (N_15075,N_14609,N_14757);
nor U15076 (N_15076,N_14538,N_14804);
nor U15077 (N_15077,N_14922,N_14726);
nand U15078 (N_15078,N_14411,N_14451);
nor U15079 (N_15079,N_14654,N_14762);
nand U15080 (N_15080,N_14952,N_14908);
nor U15081 (N_15081,N_14812,N_14696);
nand U15082 (N_15082,N_14996,N_14928);
xnor U15083 (N_15083,N_14871,N_14878);
and U15084 (N_15084,N_14848,N_14665);
or U15085 (N_15085,N_14475,N_14820);
or U15086 (N_15086,N_14854,N_14759);
and U15087 (N_15087,N_14412,N_14596);
nand U15088 (N_15088,N_14766,N_14717);
nor U15089 (N_15089,N_14433,N_14703);
or U15090 (N_15090,N_14962,N_14428);
xnor U15091 (N_15091,N_14541,N_14881);
or U15092 (N_15092,N_14491,N_14698);
nor U15093 (N_15093,N_14498,N_14509);
and U15094 (N_15094,N_14639,N_14833);
or U15095 (N_15095,N_14395,N_14980);
nor U15096 (N_15096,N_14811,N_14834);
or U15097 (N_15097,N_14626,N_14941);
and U15098 (N_15098,N_14573,N_14920);
xor U15099 (N_15099,N_14660,N_14448);
nand U15100 (N_15100,N_14512,N_14768);
nor U15101 (N_15101,N_14604,N_14571);
nor U15102 (N_15102,N_14522,N_14565);
nor U15103 (N_15103,N_14830,N_14926);
nand U15104 (N_15104,N_14380,N_14747);
nor U15105 (N_15105,N_14829,N_14484);
and U15106 (N_15106,N_14760,N_14781);
nand U15107 (N_15107,N_14548,N_14817);
nor U15108 (N_15108,N_14648,N_14492);
nor U15109 (N_15109,N_14877,N_14819);
and U15110 (N_15110,N_14672,N_14720);
and U15111 (N_15111,N_14807,N_14824);
xnor U15112 (N_15112,N_14646,N_14931);
nor U15113 (N_15113,N_14891,N_14470);
or U15114 (N_15114,N_14959,N_14957);
or U15115 (N_15115,N_14396,N_14381);
and U15116 (N_15116,N_14616,N_14892);
nor U15117 (N_15117,N_14613,N_14511);
and U15118 (N_15118,N_14566,N_14799);
nand U15119 (N_15119,N_14601,N_14642);
xor U15120 (N_15120,N_14978,N_14600);
nand U15121 (N_15121,N_14722,N_14531);
and U15122 (N_15122,N_14684,N_14545);
and U15123 (N_15123,N_14835,N_14840);
and U15124 (N_15124,N_14816,N_14505);
nand U15125 (N_15125,N_14972,N_14544);
xnor U15126 (N_15126,N_14721,N_14977);
nor U15127 (N_15127,N_14960,N_14670);
xor U15128 (N_15128,N_14445,N_14617);
nand U15129 (N_15129,N_14446,N_14514);
or U15130 (N_15130,N_14582,N_14893);
nor U15131 (N_15131,N_14623,N_14921);
or U15132 (N_15132,N_14440,N_14438);
xnor U15133 (N_15133,N_14496,N_14761);
nor U15134 (N_15134,N_14439,N_14632);
xor U15135 (N_15135,N_14669,N_14588);
or U15136 (N_15136,N_14946,N_14435);
and U15137 (N_15137,N_14403,N_14776);
xnor U15138 (N_15138,N_14687,N_14655);
nand U15139 (N_15139,N_14466,N_14856);
and U15140 (N_15140,N_14510,N_14751);
nor U15141 (N_15141,N_14618,N_14723);
and U15142 (N_15142,N_14940,N_14520);
nor U15143 (N_15143,N_14975,N_14585);
and U15144 (N_15144,N_14662,N_14676);
xnor U15145 (N_15145,N_14432,N_14443);
nand U15146 (N_15146,N_14557,N_14853);
nand U15147 (N_15147,N_14912,N_14842);
or U15148 (N_15148,N_14895,N_14993);
nor U15149 (N_15149,N_14508,N_14939);
and U15150 (N_15150,N_14388,N_14590);
nand U15151 (N_15151,N_14803,N_14515);
or U15152 (N_15152,N_14866,N_14783);
nor U15153 (N_15153,N_14763,N_14810);
nor U15154 (N_15154,N_14570,N_14461);
xor U15155 (N_15155,N_14568,N_14727);
nand U15156 (N_15156,N_14964,N_14917);
and U15157 (N_15157,N_14918,N_14990);
nor U15158 (N_15158,N_14692,N_14493);
xnor U15159 (N_15159,N_14619,N_14778);
and U15160 (N_15160,N_14635,N_14537);
and U15161 (N_15161,N_14737,N_14754);
and U15162 (N_15162,N_14562,N_14578);
or U15163 (N_15163,N_14549,N_14400);
xnor U15164 (N_15164,N_14950,N_14985);
and U15165 (N_15165,N_14902,N_14857);
and U15166 (N_15166,N_14540,N_14956);
nand U15167 (N_15167,N_14487,N_14499);
nand U15168 (N_15168,N_14592,N_14407);
xor U15169 (N_15169,N_14906,N_14741);
xor U15170 (N_15170,N_14468,N_14986);
or U15171 (N_15171,N_14524,N_14870);
xnor U15172 (N_15172,N_14953,N_14567);
or U15173 (N_15173,N_14378,N_14471);
nor U15174 (N_15174,N_14688,N_14595);
or U15175 (N_15175,N_14497,N_14982);
and U15176 (N_15176,N_14485,N_14862);
and U15177 (N_15177,N_14561,N_14454);
and U15178 (N_15178,N_14995,N_14734);
xnor U15179 (N_15179,N_14651,N_14879);
or U15180 (N_15180,N_14683,N_14961);
and U15181 (N_15181,N_14663,N_14867);
nor U15182 (N_15182,N_14797,N_14899);
or U15183 (N_15183,N_14814,N_14942);
nand U15184 (N_15184,N_14455,N_14729);
nor U15185 (N_15185,N_14847,N_14398);
or U15186 (N_15186,N_14997,N_14556);
or U15187 (N_15187,N_14503,N_14896);
nor U15188 (N_15188,N_14384,N_14598);
xor U15189 (N_15189,N_14991,N_14605);
nand U15190 (N_15190,N_14574,N_14850);
nor U15191 (N_15191,N_14958,N_14554);
nor U15192 (N_15192,N_14886,N_14712);
and U15193 (N_15193,N_14624,N_14414);
nor U15194 (N_15194,N_14427,N_14386);
or U15195 (N_15195,N_14738,N_14782);
nand U15196 (N_15196,N_14823,N_14519);
and U15197 (N_15197,N_14453,N_14489);
nor U15198 (N_15198,N_14641,N_14979);
xor U15199 (N_15199,N_14535,N_14533);
xnor U15200 (N_15200,N_14800,N_14467);
xnor U15201 (N_15201,N_14589,N_14705);
xnor U15202 (N_15202,N_14586,N_14441);
xor U15203 (N_15203,N_14419,N_14652);
and U15204 (N_15204,N_14420,N_14666);
and U15205 (N_15205,N_14772,N_14406);
nand U15206 (N_15206,N_14924,N_14965);
nor U15207 (N_15207,N_14599,N_14943);
or U15208 (N_15208,N_14880,N_14947);
nand U15209 (N_15209,N_14815,N_14685);
and U15210 (N_15210,N_14790,N_14994);
nand U15211 (N_15211,N_14664,N_14436);
xnor U15212 (N_15212,N_14558,N_14638);
xor U15213 (N_15213,N_14748,N_14935);
nand U15214 (N_15214,N_14402,N_14984);
xor U15215 (N_15215,N_14636,N_14929);
and U15216 (N_15216,N_14699,N_14704);
or U15217 (N_15217,N_14689,N_14858);
xor U15218 (N_15218,N_14821,N_14490);
nand U15219 (N_15219,N_14739,N_14795);
and U15220 (N_15220,N_14462,N_14787);
nand U15221 (N_15221,N_14691,N_14682);
nand U15222 (N_15222,N_14580,N_14869);
nand U15223 (N_15223,N_14808,N_14826);
xnor U15224 (N_15224,N_14967,N_14966);
nor U15225 (N_15225,N_14992,N_14743);
xor U15226 (N_15226,N_14809,N_14385);
nand U15227 (N_15227,N_14547,N_14611);
nand U15228 (N_15228,N_14634,N_14753);
and U15229 (N_15229,N_14426,N_14887);
nand U15230 (N_15230,N_14401,N_14625);
nand U15231 (N_15231,N_14786,N_14775);
nor U15232 (N_15232,N_14383,N_14513);
nand U15233 (N_15233,N_14555,N_14828);
or U15234 (N_15234,N_14629,N_14839);
and U15235 (N_15235,N_14927,N_14872);
and U15236 (N_15236,N_14504,N_14606);
nand U15237 (N_15237,N_14424,N_14597);
nor U15238 (N_15238,N_14938,N_14897);
nand U15239 (N_15239,N_14843,N_14933);
nor U15240 (N_15240,N_14805,N_14476);
nor U15241 (N_15241,N_14937,N_14925);
and U15242 (N_15242,N_14678,N_14627);
nor U15243 (N_15243,N_14668,N_14494);
and U15244 (N_15244,N_14780,N_14849);
and U15245 (N_15245,N_14607,N_14560);
nor U15246 (N_15246,N_14482,N_14564);
xor U15247 (N_15247,N_14630,N_14889);
xor U15248 (N_15248,N_14949,N_14581);
xnor U15249 (N_15249,N_14532,N_14905);
nand U15250 (N_15250,N_14391,N_14507);
or U15251 (N_15251,N_14948,N_14444);
nor U15252 (N_15252,N_14425,N_14774);
xnor U15253 (N_15253,N_14983,N_14934);
nand U15254 (N_15254,N_14393,N_14919);
nor U15255 (N_15255,N_14474,N_14603);
xnor U15256 (N_15256,N_14900,N_14836);
nand U15257 (N_15257,N_14951,N_14552);
xnor U15258 (N_15258,N_14735,N_14527);
or U15259 (N_15259,N_14846,N_14569);
and U15260 (N_15260,N_14657,N_14473);
xnor U15261 (N_15261,N_14523,N_14746);
xor U15262 (N_15262,N_14525,N_14434);
and U15263 (N_15263,N_14864,N_14583);
xor U15264 (N_15264,N_14731,N_14792);
xor U15265 (N_15265,N_14410,N_14479);
or U15266 (N_15266,N_14865,N_14714);
nand U15267 (N_15267,N_14888,N_14608);
nand U15268 (N_15268,N_14382,N_14576);
nor U15269 (N_15269,N_14375,N_14725);
xor U15270 (N_15270,N_14923,N_14472);
nor U15271 (N_15271,N_14851,N_14890);
or U15272 (N_15272,N_14868,N_14679);
and U15273 (N_15273,N_14649,N_14587);
or U15274 (N_15274,N_14708,N_14661);
nor U15275 (N_15275,N_14944,N_14837);
or U15276 (N_15276,N_14521,N_14469);
or U15277 (N_15277,N_14681,N_14593);
and U15278 (N_15278,N_14719,N_14885);
nand U15279 (N_15279,N_14680,N_14745);
xnor U15280 (N_15280,N_14945,N_14572);
nor U15281 (N_15281,N_14622,N_14644);
or U15282 (N_15282,N_14764,N_14449);
xor U15283 (N_15283,N_14653,N_14390);
nand U15284 (N_15284,N_14529,N_14732);
xnor U15285 (N_15285,N_14633,N_14852);
nor U15286 (N_15286,N_14999,N_14488);
or U15287 (N_15287,N_14901,N_14694);
xor U15288 (N_15288,N_14442,N_14936);
nand U15289 (N_15289,N_14930,N_14707);
nor U15290 (N_15290,N_14423,N_14422);
nand U15291 (N_15291,N_14838,N_14464);
or U15292 (N_15292,N_14974,N_14742);
nand U15293 (N_15293,N_14841,N_14987);
and U15294 (N_15294,N_14718,N_14460);
nor U15295 (N_15295,N_14911,N_14758);
xor U15296 (N_15296,N_14546,N_14822);
xnor U15297 (N_15297,N_14437,N_14702);
nand U15298 (N_15298,N_14700,N_14413);
nor U15299 (N_15299,N_14875,N_14417);
or U15300 (N_15300,N_14612,N_14693);
and U15301 (N_15301,N_14773,N_14859);
nand U15302 (N_15302,N_14954,N_14640);
or U15303 (N_15303,N_14724,N_14559);
xnor U15304 (N_15304,N_14421,N_14998);
nor U15305 (N_15305,N_14798,N_14506);
and U15306 (N_15306,N_14711,N_14628);
or U15307 (N_15307,N_14784,N_14860);
nand U15308 (N_15308,N_14932,N_14903);
xor U15309 (N_15309,N_14409,N_14876);
nand U15310 (N_15310,N_14988,N_14769);
or U15311 (N_15311,N_14916,N_14452);
nor U15312 (N_15312,N_14458,N_14410);
nor U15313 (N_15313,N_14588,N_14641);
or U15314 (N_15314,N_14567,N_14906);
xnor U15315 (N_15315,N_14643,N_14717);
xnor U15316 (N_15316,N_14587,N_14390);
or U15317 (N_15317,N_14709,N_14478);
and U15318 (N_15318,N_14967,N_14748);
and U15319 (N_15319,N_14684,N_14619);
and U15320 (N_15320,N_14669,N_14504);
and U15321 (N_15321,N_14580,N_14910);
nor U15322 (N_15322,N_14588,N_14495);
and U15323 (N_15323,N_14904,N_14939);
nand U15324 (N_15324,N_14423,N_14994);
or U15325 (N_15325,N_14583,N_14593);
or U15326 (N_15326,N_14874,N_14655);
and U15327 (N_15327,N_14997,N_14437);
nor U15328 (N_15328,N_14481,N_14759);
nand U15329 (N_15329,N_14613,N_14411);
nand U15330 (N_15330,N_14589,N_14836);
nor U15331 (N_15331,N_14605,N_14407);
nor U15332 (N_15332,N_14709,N_14670);
nand U15333 (N_15333,N_14600,N_14722);
nand U15334 (N_15334,N_14486,N_14620);
nand U15335 (N_15335,N_14829,N_14854);
xnor U15336 (N_15336,N_14646,N_14837);
or U15337 (N_15337,N_14691,N_14584);
nand U15338 (N_15338,N_14978,N_14510);
nand U15339 (N_15339,N_14962,N_14402);
or U15340 (N_15340,N_14901,N_14379);
and U15341 (N_15341,N_14503,N_14981);
or U15342 (N_15342,N_14742,N_14421);
nand U15343 (N_15343,N_14867,N_14565);
or U15344 (N_15344,N_14909,N_14997);
and U15345 (N_15345,N_14850,N_14712);
nor U15346 (N_15346,N_14848,N_14667);
nand U15347 (N_15347,N_14717,N_14701);
or U15348 (N_15348,N_14453,N_14768);
and U15349 (N_15349,N_14552,N_14550);
and U15350 (N_15350,N_14997,N_14778);
or U15351 (N_15351,N_14512,N_14982);
or U15352 (N_15352,N_14861,N_14797);
xnor U15353 (N_15353,N_14806,N_14748);
and U15354 (N_15354,N_14923,N_14753);
and U15355 (N_15355,N_14992,N_14729);
nand U15356 (N_15356,N_14551,N_14891);
and U15357 (N_15357,N_14490,N_14699);
nand U15358 (N_15358,N_14796,N_14893);
xnor U15359 (N_15359,N_14632,N_14547);
xnor U15360 (N_15360,N_14903,N_14642);
nand U15361 (N_15361,N_14569,N_14736);
or U15362 (N_15362,N_14847,N_14627);
nor U15363 (N_15363,N_14861,N_14655);
or U15364 (N_15364,N_14726,N_14871);
nand U15365 (N_15365,N_14666,N_14870);
and U15366 (N_15366,N_14980,N_14623);
nand U15367 (N_15367,N_14927,N_14946);
and U15368 (N_15368,N_14637,N_14987);
nand U15369 (N_15369,N_14682,N_14647);
nand U15370 (N_15370,N_14958,N_14807);
and U15371 (N_15371,N_14428,N_14375);
nor U15372 (N_15372,N_14515,N_14487);
and U15373 (N_15373,N_14647,N_14640);
nor U15374 (N_15374,N_14797,N_14826);
or U15375 (N_15375,N_14953,N_14935);
and U15376 (N_15376,N_14675,N_14453);
nor U15377 (N_15377,N_14614,N_14844);
xnor U15378 (N_15378,N_14729,N_14514);
xnor U15379 (N_15379,N_14386,N_14862);
nor U15380 (N_15380,N_14743,N_14645);
or U15381 (N_15381,N_14559,N_14768);
xor U15382 (N_15382,N_14529,N_14808);
xnor U15383 (N_15383,N_14638,N_14553);
or U15384 (N_15384,N_14968,N_14454);
and U15385 (N_15385,N_14503,N_14409);
nor U15386 (N_15386,N_14896,N_14780);
nor U15387 (N_15387,N_14438,N_14890);
or U15388 (N_15388,N_14642,N_14836);
or U15389 (N_15389,N_14418,N_14513);
and U15390 (N_15390,N_14392,N_14733);
nor U15391 (N_15391,N_14703,N_14705);
and U15392 (N_15392,N_14779,N_14599);
xor U15393 (N_15393,N_14898,N_14427);
xor U15394 (N_15394,N_14685,N_14741);
or U15395 (N_15395,N_14512,N_14523);
nor U15396 (N_15396,N_14407,N_14689);
or U15397 (N_15397,N_14399,N_14409);
nor U15398 (N_15398,N_14727,N_14949);
and U15399 (N_15399,N_14822,N_14621);
or U15400 (N_15400,N_14833,N_14940);
or U15401 (N_15401,N_14721,N_14467);
or U15402 (N_15402,N_14460,N_14511);
or U15403 (N_15403,N_14520,N_14463);
xnor U15404 (N_15404,N_14440,N_14471);
or U15405 (N_15405,N_14887,N_14847);
and U15406 (N_15406,N_14502,N_14975);
or U15407 (N_15407,N_14644,N_14525);
or U15408 (N_15408,N_14464,N_14744);
or U15409 (N_15409,N_14804,N_14796);
nor U15410 (N_15410,N_14843,N_14571);
nor U15411 (N_15411,N_14795,N_14819);
and U15412 (N_15412,N_14829,N_14941);
nand U15413 (N_15413,N_14481,N_14464);
or U15414 (N_15414,N_14790,N_14521);
nand U15415 (N_15415,N_14991,N_14589);
nand U15416 (N_15416,N_14757,N_14655);
or U15417 (N_15417,N_14509,N_14665);
nor U15418 (N_15418,N_14608,N_14501);
or U15419 (N_15419,N_14400,N_14667);
or U15420 (N_15420,N_14546,N_14682);
and U15421 (N_15421,N_14580,N_14883);
nor U15422 (N_15422,N_14589,N_14527);
nor U15423 (N_15423,N_14554,N_14829);
or U15424 (N_15424,N_14990,N_14858);
and U15425 (N_15425,N_14938,N_14598);
or U15426 (N_15426,N_14981,N_14483);
nor U15427 (N_15427,N_14430,N_14633);
or U15428 (N_15428,N_14422,N_14931);
nand U15429 (N_15429,N_14971,N_14847);
and U15430 (N_15430,N_14796,N_14675);
and U15431 (N_15431,N_14547,N_14512);
xor U15432 (N_15432,N_14844,N_14723);
and U15433 (N_15433,N_14610,N_14447);
and U15434 (N_15434,N_14646,N_14579);
nor U15435 (N_15435,N_14611,N_14482);
xnor U15436 (N_15436,N_14499,N_14927);
nand U15437 (N_15437,N_14798,N_14476);
nand U15438 (N_15438,N_14623,N_14381);
or U15439 (N_15439,N_14772,N_14956);
and U15440 (N_15440,N_14876,N_14619);
xor U15441 (N_15441,N_14992,N_14384);
nor U15442 (N_15442,N_14826,N_14789);
nor U15443 (N_15443,N_14590,N_14568);
nand U15444 (N_15444,N_14929,N_14760);
nand U15445 (N_15445,N_14913,N_14819);
nand U15446 (N_15446,N_14808,N_14736);
nor U15447 (N_15447,N_14937,N_14879);
or U15448 (N_15448,N_14686,N_14660);
nor U15449 (N_15449,N_14833,N_14870);
or U15450 (N_15450,N_14704,N_14606);
or U15451 (N_15451,N_14916,N_14789);
and U15452 (N_15452,N_14890,N_14958);
or U15453 (N_15453,N_14605,N_14482);
nand U15454 (N_15454,N_14790,N_14677);
or U15455 (N_15455,N_14924,N_14953);
xnor U15456 (N_15456,N_14655,N_14380);
nor U15457 (N_15457,N_14382,N_14736);
xor U15458 (N_15458,N_14409,N_14885);
nor U15459 (N_15459,N_14749,N_14507);
and U15460 (N_15460,N_14575,N_14507);
nor U15461 (N_15461,N_14982,N_14438);
and U15462 (N_15462,N_14957,N_14518);
nor U15463 (N_15463,N_14818,N_14963);
nand U15464 (N_15464,N_14512,N_14710);
and U15465 (N_15465,N_14563,N_14910);
nor U15466 (N_15466,N_14522,N_14942);
nor U15467 (N_15467,N_14574,N_14381);
or U15468 (N_15468,N_14606,N_14883);
xor U15469 (N_15469,N_14748,N_14884);
nand U15470 (N_15470,N_14813,N_14416);
or U15471 (N_15471,N_14859,N_14789);
or U15472 (N_15472,N_14537,N_14774);
and U15473 (N_15473,N_14381,N_14974);
or U15474 (N_15474,N_14716,N_14517);
nor U15475 (N_15475,N_14485,N_14886);
nor U15476 (N_15476,N_14537,N_14833);
xnor U15477 (N_15477,N_14741,N_14502);
xnor U15478 (N_15478,N_14688,N_14785);
nor U15479 (N_15479,N_14444,N_14647);
nor U15480 (N_15480,N_14499,N_14484);
xor U15481 (N_15481,N_14718,N_14438);
and U15482 (N_15482,N_14762,N_14671);
or U15483 (N_15483,N_14433,N_14731);
and U15484 (N_15484,N_14795,N_14918);
nor U15485 (N_15485,N_14917,N_14644);
and U15486 (N_15486,N_14514,N_14454);
and U15487 (N_15487,N_14883,N_14886);
nor U15488 (N_15488,N_14896,N_14591);
and U15489 (N_15489,N_14383,N_14599);
nand U15490 (N_15490,N_14380,N_14476);
nor U15491 (N_15491,N_14609,N_14825);
or U15492 (N_15492,N_14626,N_14665);
or U15493 (N_15493,N_14521,N_14597);
or U15494 (N_15494,N_14550,N_14418);
and U15495 (N_15495,N_14582,N_14996);
or U15496 (N_15496,N_14969,N_14582);
or U15497 (N_15497,N_14864,N_14607);
and U15498 (N_15498,N_14566,N_14640);
nor U15499 (N_15499,N_14961,N_14859);
and U15500 (N_15500,N_14899,N_14646);
nand U15501 (N_15501,N_14696,N_14906);
or U15502 (N_15502,N_14541,N_14376);
or U15503 (N_15503,N_14440,N_14930);
nor U15504 (N_15504,N_14782,N_14415);
or U15505 (N_15505,N_14473,N_14732);
xnor U15506 (N_15506,N_14486,N_14493);
nand U15507 (N_15507,N_14452,N_14802);
nand U15508 (N_15508,N_14569,N_14428);
nor U15509 (N_15509,N_14866,N_14770);
nor U15510 (N_15510,N_14816,N_14922);
and U15511 (N_15511,N_14980,N_14971);
xor U15512 (N_15512,N_14759,N_14517);
or U15513 (N_15513,N_14927,N_14701);
or U15514 (N_15514,N_14681,N_14777);
nand U15515 (N_15515,N_14828,N_14891);
nand U15516 (N_15516,N_14512,N_14686);
nor U15517 (N_15517,N_14644,N_14697);
nor U15518 (N_15518,N_14526,N_14894);
nand U15519 (N_15519,N_14433,N_14587);
nor U15520 (N_15520,N_14452,N_14998);
and U15521 (N_15521,N_14863,N_14984);
and U15522 (N_15522,N_14507,N_14493);
nor U15523 (N_15523,N_14573,N_14918);
xnor U15524 (N_15524,N_14502,N_14903);
nand U15525 (N_15525,N_14899,N_14613);
nor U15526 (N_15526,N_14467,N_14885);
xnor U15527 (N_15527,N_14714,N_14441);
nor U15528 (N_15528,N_14429,N_14650);
or U15529 (N_15529,N_14448,N_14912);
or U15530 (N_15530,N_14486,N_14871);
nor U15531 (N_15531,N_14953,N_14443);
xor U15532 (N_15532,N_14425,N_14451);
or U15533 (N_15533,N_14860,N_14487);
and U15534 (N_15534,N_14847,N_14493);
and U15535 (N_15535,N_14699,N_14444);
nand U15536 (N_15536,N_14402,N_14488);
and U15537 (N_15537,N_14528,N_14984);
xnor U15538 (N_15538,N_14821,N_14902);
and U15539 (N_15539,N_14458,N_14703);
nor U15540 (N_15540,N_14881,N_14462);
and U15541 (N_15541,N_14660,N_14498);
nand U15542 (N_15542,N_14583,N_14445);
xor U15543 (N_15543,N_14972,N_14963);
nor U15544 (N_15544,N_14835,N_14683);
or U15545 (N_15545,N_14495,N_14823);
nand U15546 (N_15546,N_14997,N_14941);
and U15547 (N_15547,N_14718,N_14636);
nor U15548 (N_15548,N_14926,N_14458);
xnor U15549 (N_15549,N_14543,N_14772);
or U15550 (N_15550,N_14823,N_14720);
and U15551 (N_15551,N_14455,N_14395);
nand U15552 (N_15552,N_14651,N_14687);
xor U15553 (N_15553,N_14425,N_14592);
or U15554 (N_15554,N_14541,N_14679);
xnor U15555 (N_15555,N_14872,N_14520);
xor U15556 (N_15556,N_14896,N_14889);
nor U15557 (N_15557,N_14997,N_14861);
or U15558 (N_15558,N_14667,N_14410);
nor U15559 (N_15559,N_14937,N_14383);
and U15560 (N_15560,N_14704,N_14443);
and U15561 (N_15561,N_14598,N_14555);
nand U15562 (N_15562,N_14878,N_14835);
nor U15563 (N_15563,N_14615,N_14888);
or U15564 (N_15564,N_14389,N_14622);
xnor U15565 (N_15565,N_14690,N_14596);
nand U15566 (N_15566,N_14513,N_14452);
xor U15567 (N_15567,N_14729,N_14581);
and U15568 (N_15568,N_14769,N_14721);
xnor U15569 (N_15569,N_14402,N_14431);
or U15570 (N_15570,N_14377,N_14575);
and U15571 (N_15571,N_14429,N_14958);
xnor U15572 (N_15572,N_14669,N_14478);
nor U15573 (N_15573,N_14997,N_14417);
nand U15574 (N_15574,N_14610,N_14624);
nand U15575 (N_15575,N_14384,N_14982);
nor U15576 (N_15576,N_14559,N_14851);
nor U15577 (N_15577,N_14992,N_14956);
nor U15578 (N_15578,N_14664,N_14521);
or U15579 (N_15579,N_14535,N_14590);
or U15580 (N_15580,N_14686,N_14779);
or U15581 (N_15581,N_14500,N_14593);
nor U15582 (N_15582,N_14657,N_14610);
and U15583 (N_15583,N_14433,N_14733);
xnor U15584 (N_15584,N_14979,N_14801);
nor U15585 (N_15585,N_14980,N_14739);
or U15586 (N_15586,N_14769,N_14798);
nand U15587 (N_15587,N_14460,N_14866);
nor U15588 (N_15588,N_14488,N_14452);
xor U15589 (N_15589,N_14568,N_14483);
xnor U15590 (N_15590,N_14635,N_14888);
or U15591 (N_15591,N_14728,N_14913);
and U15592 (N_15592,N_14742,N_14397);
nand U15593 (N_15593,N_14671,N_14696);
xor U15594 (N_15594,N_14842,N_14546);
and U15595 (N_15595,N_14994,N_14874);
xor U15596 (N_15596,N_14512,N_14428);
xor U15597 (N_15597,N_14709,N_14578);
nor U15598 (N_15598,N_14561,N_14469);
nand U15599 (N_15599,N_14827,N_14443);
and U15600 (N_15600,N_14678,N_14523);
and U15601 (N_15601,N_14664,N_14507);
nor U15602 (N_15602,N_14465,N_14545);
nor U15603 (N_15603,N_14875,N_14939);
and U15604 (N_15604,N_14448,N_14501);
nor U15605 (N_15605,N_14631,N_14974);
or U15606 (N_15606,N_14849,N_14992);
xnor U15607 (N_15607,N_14918,N_14728);
or U15608 (N_15608,N_14520,N_14705);
or U15609 (N_15609,N_14680,N_14779);
nor U15610 (N_15610,N_14738,N_14678);
xnor U15611 (N_15611,N_14485,N_14816);
xor U15612 (N_15612,N_14770,N_14863);
nor U15613 (N_15613,N_14905,N_14577);
or U15614 (N_15614,N_14798,N_14520);
and U15615 (N_15615,N_14661,N_14970);
nor U15616 (N_15616,N_14560,N_14460);
nor U15617 (N_15617,N_14428,N_14658);
and U15618 (N_15618,N_14721,N_14535);
xor U15619 (N_15619,N_14528,N_14679);
and U15620 (N_15620,N_14625,N_14564);
nor U15621 (N_15621,N_14548,N_14450);
and U15622 (N_15622,N_14486,N_14821);
and U15623 (N_15623,N_14929,N_14785);
nor U15624 (N_15624,N_14649,N_14495);
nor U15625 (N_15625,N_15296,N_15616);
nor U15626 (N_15626,N_15354,N_15340);
or U15627 (N_15627,N_15197,N_15112);
nor U15628 (N_15628,N_15143,N_15017);
nand U15629 (N_15629,N_15499,N_15294);
nand U15630 (N_15630,N_15398,N_15267);
xnor U15631 (N_15631,N_15566,N_15129);
xnor U15632 (N_15632,N_15297,N_15302);
nor U15633 (N_15633,N_15490,N_15356);
xnor U15634 (N_15634,N_15567,N_15344);
nor U15635 (N_15635,N_15313,N_15127);
and U15636 (N_15636,N_15259,N_15561);
and U15637 (N_15637,N_15138,N_15236);
nor U15638 (N_15638,N_15170,N_15406);
xor U15639 (N_15639,N_15521,N_15016);
nor U15640 (N_15640,N_15229,N_15169);
or U15641 (N_15641,N_15046,N_15612);
xnor U15642 (N_15642,N_15393,N_15055);
or U15643 (N_15643,N_15115,N_15200);
xnor U15644 (N_15644,N_15492,N_15333);
or U15645 (N_15645,N_15311,N_15149);
or U15646 (N_15646,N_15166,N_15152);
and U15647 (N_15647,N_15537,N_15586);
xor U15648 (N_15648,N_15319,N_15349);
or U15649 (N_15649,N_15188,N_15425);
nand U15650 (N_15650,N_15601,N_15308);
and U15651 (N_15651,N_15044,N_15225);
nor U15652 (N_15652,N_15462,N_15284);
nor U15653 (N_15653,N_15010,N_15325);
xor U15654 (N_15654,N_15584,N_15224);
nand U15655 (N_15655,N_15079,N_15494);
or U15656 (N_15656,N_15565,N_15193);
and U15657 (N_15657,N_15029,N_15518);
xnor U15658 (N_15658,N_15263,N_15108);
and U15659 (N_15659,N_15620,N_15502);
or U15660 (N_15660,N_15126,N_15179);
or U15661 (N_15661,N_15360,N_15542);
nand U15662 (N_15662,N_15597,N_15098);
and U15663 (N_15663,N_15615,N_15417);
and U15664 (N_15664,N_15124,N_15051);
nand U15665 (N_15665,N_15575,N_15275);
nor U15666 (N_15666,N_15345,N_15059);
and U15667 (N_15667,N_15387,N_15441);
xor U15668 (N_15668,N_15581,N_15008);
and U15669 (N_15669,N_15205,N_15142);
and U15670 (N_15670,N_15135,N_15505);
nor U15671 (N_15671,N_15270,N_15107);
nor U15672 (N_15672,N_15524,N_15272);
or U15673 (N_15673,N_15165,N_15426);
nand U15674 (N_15674,N_15181,N_15508);
and U15675 (N_15675,N_15442,N_15621);
xor U15676 (N_15676,N_15266,N_15276);
or U15677 (N_15677,N_15409,N_15289);
nand U15678 (N_15678,N_15128,N_15243);
nor U15679 (N_15679,N_15538,N_15024);
nor U15680 (N_15680,N_15255,N_15322);
nor U15681 (N_15681,N_15549,N_15412);
xnor U15682 (N_15682,N_15609,N_15047);
or U15683 (N_15683,N_15058,N_15240);
nand U15684 (N_15684,N_15156,N_15230);
or U15685 (N_15685,N_15323,N_15336);
xnor U15686 (N_15686,N_15217,N_15591);
nor U15687 (N_15687,N_15429,N_15277);
or U15688 (N_15688,N_15171,N_15174);
xnor U15689 (N_15689,N_15557,N_15421);
xnor U15690 (N_15690,N_15383,N_15301);
xnor U15691 (N_15691,N_15030,N_15032);
nand U15692 (N_15692,N_15511,N_15137);
or U15693 (N_15693,N_15083,N_15530);
nand U15694 (N_15694,N_15448,N_15209);
nor U15695 (N_15695,N_15309,N_15196);
xor U15696 (N_15696,N_15210,N_15062);
nor U15697 (N_15697,N_15465,N_15004);
and U15698 (N_15698,N_15026,N_15592);
xor U15699 (N_15699,N_15324,N_15361);
and U15700 (N_15700,N_15555,N_15221);
or U15701 (N_15701,N_15559,N_15553);
and U15702 (N_15702,N_15624,N_15019);
xor U15703 (N_15703,N_15139,N_15214);
nor U15704 (N_15704,N_15435,N_15326);
nor U15705 (N_15705,N_15509,N_15510);
and U15706 (N_15706,N_15239,N_15121);
or U15707 (N_15707,N_15254,N_15379);
xnor U15708 (N_15708,N_15479,N_15274);
xnor U15709 (N_15709,N_15410,N_15558);
xnor U15710 (N_15710,N_15076,N_15038);
nor U15711 (N_15711,N_15623,N_15212);
xnor U15712 (N_15712,N_15288,N_15613);
and U15713 (N_15713,N_15244,N_15574);
and U15714 (N_15714,N_15560,N_15251);
nor U15715 (N_15715,N_15310,N_15457);
xnor U15716 (N_15716,N_15105,N_15431);
nor U15717 (N_15717,N_15529,N_15416);
or U15718 (N_15718,N_15204,N_15110);
nand U15719 (N_15719,N_15201,N_15271);
or U15720 (N_15720,N_15415,N_15485);
xnor U15721 (N_15721,N_15118,N_15213);
nand U15722 (N_15722,N_15056,N_15388);
xor U15723 (N_15723,N_15473,N_15245);
and U15724 (N_15724,N_15164,N_15475);
nor U15725 (N_15725,N_15268,N_15295);
or U15726 (N_15726,N_15380,N_15516);
nor U15727 (N_15727,N_15596,N_15403);
nor U15728 (N_15728,N_15178,N_15104);
nand U15729 (N_15729,N_15544,N_15235);
xor U15730 (N_15730,N_15595,N_15351);
xnor U15731 (N_15731,N_15015,N_15327);
xnor U15732 (N_15732,N_15283,N_15081);
nand U15733 (N_15733,N_15172,N_15192);
or U15734 (N_15734,N_15452,N_15523);
nor U15735 (N_15735,N_15202,N_15394);
or U15736 (N_15736,N_15419,N_15247);
nor U15737 (N_15737,N_15150,N_15021);
and U15738 (N_15738,N_15552,N_15018);
nor U15739 (N_15739,N_15023,N_15153);
and U15740 (N_15740,N_15378,N_15500);
nand U15741 (N_15741,N_15265,N_15604);
or U15742 (N_15742,N_15374,N_15386);
xor U15743 (N_15743,N_15260,N_15158);
nor U15744 (N_15744,N_15161,N_15232);
xnor U15745 (N_15745,N_15547,N_15446);
or U15746 (N_15746,N_15414,N_15009);
and U15747 (N_15747,N_15183,N_15337);
nor U15748 (N_15748,N_15102,N_15472);
nor U15749 (N_15749,N_15003,N_15256);
nor U15750 (N_15750,N_15582,N_15054);
and U15751 (N_15751,N_15314,N_15321);
nor U15752 (N_15752,N_15618,N_15233);
and U15753 (N_15753,N_15001,N_15238);
xor U15754 (N_15754,N_15608,N_15501);
nor U15755 (N_15755,N_15223,N_15078);
or U15756 (N_15756,N_15532,N_15151);
nand U15757 (N_15757,N_15437,N_15569);
xor U15758 (N_15758,N_15052,N_15159);
nand U15759 (N_15759,N_15610,N_15342);
nor U15760 (N_15760,N_15488,N_15194);
and U15761 (N_15761,N_15384,N_15514);
xor U15762 (N_15762,N_15487,N_15042);
nor U15763 (N_15763,N_15546,N_15136);
or U15764 (N_15764,N_15031,N_15182);
xnor U15765 (N_15765,N_15306,N_15450);
xor U15766 (N_15766,N_15145,N_15113);
or U15767 (N_15767,N_15373,N_15065);
nor U15768 (N_15768,N_15368,N_15504);
nand U15769 (N_15769,N_15400,N_15377);
xnor U15770 (N_15770,N_15167,N_15404);
and U15771 (N_15771,N_15061,N_15594);
or U15772 (N_15772,N_15366,N_15503);
and U15773 (N_15773,N_15035,N_15125);
or U15774 (N_15774,N_15453,N_15341);
nor U15775 (N_15775,N_15449,N_15307);
nand U15776 (N_15776,N_15376,N_15563);
nor U15777 (N_15777,N_15572,N_15067);
and U15778 (N_15778,N_15533,N_15157);
nor U15779 (N_15779,N_15605,N_15428);
or U15780 (N_15780,N_15034,N_15060);
xnor U15781 (N_15781,N_15071,N_15292);
or U15782 (N_15782,N_15474,N_15116);
nand U15783 (N_15783,N_15550,N_15535);
and U15784 (N_15784,N_15362,N_15439);
nor U15785 (N_15785,N_15445,N_15619);
xnor U15786 (N_15786,N_15534,N_15513);
and U15787 (N_15787,N_15028,N_15000);
or U15788 (N_15788,N_15423,N_15576);
nand U15789 (N_15789,N_15334,N_15543);
xor U15790 (N_15790,N_15607,N_15068);
or U15791 (N_15791,N_15617,N_15131);
nor U15792 (N_15792,N_15208,N_15285);
xor U15793 (N_15793,N_15303,N_15525);
and U15794 (N_15794,N_15231,N_15287);
nand U15795 (N_15795,N_15427,N_15057);
xnor U15796 (N_15796,N_15072,N_15162);
and U15797 (N_15797,N_15541,N_15467);
or U15798 (N_15798,N_15216,N_15461);
or U15799 (N_15799,N_15082,N_15536);
or U15800 (N_15800,N_15471,N_15364);
or U15801 (N_15801,N_15358,N_15025);
or U15802 (N_15802,N_15154,N_15352);
nand U15803 (N_15803,N_15290,N_15433);
xor U15804 (N_15804,N_15237,N_15088);
nor U15805 (N_15805,N_15049,N_15579);
nor U15806 (N_15806,N_15005,N_15495);
nor U15807 (N_15807,N_15073,N_15329);
or U15808 (N_15808,N_15335,N_15583);
or U15809 (N_15809,N_15053,N_15163);
xor U15810 (N_15810,N_15177,N_15087);
nor U15811 (N_15811,N_15248,N_15228);
and U15812 (N_15812,N_15033,N_15482);
and U15813 (N_15813,N_15041,N_15347);
or U15814 (N_15814,N_15093,N_15346);
xor U15815 (N_15815,N_15070,N_15548);
or U15816 (N_15816,N_15084,N_15522);
nor U15817 (N_15817,N_15278,N_15066);
or U15818 (N_15818,N_15382,N_15585);
and U15819 (N_15819,N_15220,N_15027);
nand U15820 (N_15820,N_15211,N_15578);
and U15821 (N_15821,N_15614,N_15189);
or U15822 (N_15822,N_15350,N_15593);
xor U15823 (N_15823,N_15381,N_15043);
nand U15824 (N_15824,N_15447,N_15074);
or U15825 (N_15825,N_15440,N_15249);
or U15826 (N_15826,N_15551,N_15463);
nand U15827 (N_15827,N_15097,N_15198);
nand U15828 (N_15828,N_15117,N_15391);
and U15829 (N_15829,N_15257,N_15246);
nand U15830 (N_15830,N_15119,N_15286);
and U15831 (N_15831,N_15291,N_15353);
or U15832 (N_15832,N_15497,N_15133);
nor U15833 (N_15833,N_15491,N_15064);
xor U15834 (N_15834,N_15106,N_15422);
and U15835 (N_15835,N_15395,N_15280);
nor U15836 (N_15836,N_15480,N_15101);
nand U15837 (N_15837,N_15331,N_15191);
nor U15838 (N_15838,N_15262,N_15040);
and U15839 (N_15839,N_15526,N_15587);
nand U15840 (N_15840,N_15570,N_15436);
and U15841 (N_15841,N_15556,N_15180);
xnor U15842 (N_15842,N_15468,N_15269);
or U15843 (N_15843,N_15554,N_15493);
or U15844 (N_15844,N_15094,N_15090);
nor U15845 (N_15845,N_15506,N_15222);
nand U15846 (N_15846,N_15517,N_15199);
or U15847 (N_15847,N_15375,N_15226);
nor U15848 (N_15848,N_15515,N_15122);
nand U15849 (N_15849,N_15092,N_15011);
and U15850 (N_15850,N_15564,N_15185);
or U15851 (N_15851,N_15372,N_15397);
nand U15852 (N_15852,N_15464,N_15568);
or U15853 (N_15853,N_15218,N_15330);
nand U15854 (N_15854,N_15173,N_15466);
xnor U15855 (N_15855,N_15519,N_15147);
nor U15856 (N_15856,N_15408,N_15577);
xnor U15857 (N_15857,N_15022,N_15316);
and U15858 (N_15858,N_15469,N_15120);
nand U15859 (N_15859,N_15187,N_15545);
xnor U15860 (N_15860,N_15432,N_15063);
nor U15861 (N_15861,N_15273,N_15370);
and U15862 (N_15862,N_15085,N_15075);
and U15863 (N_15863,N_15298,N_15571);
nor U15864 (N_15864,N_15328,N_15250);
xor U15865 (N_15865,N_15012,N_15091);
nor U15866 (N_15866,N_15455,N_15389);
nor U15867 (N_15867,N_15014,N_15252);
or U15868 (N_15868,N_15606,N_15281);
or U15869 (N_15869,N_15589,N_15603);
xor U15870 (N_15870,N_15095,N_15176);
nor U15871 (N_15871,N_15103,N_15300);
nand U15872 (N_15872,N_15484,N_15407);
nor U15873 (N_15873,N_15434,N_15206);
xor U15874 (N_15874,N_15369,N_15343);
nand U15875 (N_15875,N_15454,N_15520);
nand U15876 (N_15876,N_15600,N_15020);
nor U15877 (N_15877,N_15320,N_15599);
xnor U15878 (N_15878,N_15175,N_15168);
nand U15879 (N_15879,N_15392,N_15512);
nor U15880 (N_15880,N_15590,N_15007);
nand U15881 (N_15881,N_15402,N_15481);
nand U15882 (N_15882,N_15050,N_15299);
or U15883 (N_15883,N_15258,N_15588);
nor U15884 (N_15884,N_15317,N_15477);
nor U15885 (N_15885,N_15456,N_15048);
nand U15886 (N_15886,N_15315,N_15451);
and U15887 (N_15887,N_15045,N_15365);
and U15888 (N_15888,N_15359,N_15155);
xnor U15889 (N_15889,N_15305,N_15332);
xnor U15890 (N_15890,N_15195,N_15486);
or U15891 (N_15891,N_15443,N_15099);
or U15892 (N_15892,N_15219,N_15390);
or U15893 (N_15893,N_15489,N_15227);
nand U15894 (N_15894,N_15430,N_15241);
nand U15895 (N_15895,N_15242,N_15215);
nor U15896 (N_15896,N_15496,N_15363);
nor U15897 (N_15897,N_15186,N_15540);
xnor U15898 (N_15898,N_15203,N_15413);
nor U15899 (N_15899,N_15405,N_15318);
nor U15900 (N_15900,N_15411,N_15140);
or U15901 (N_15901,N_15483,N_15562);
nand U15902 (N_15902,N_15144,N_15111);
or U15903 (N_15903,N_15385,N_15253);
or U15904 (N_15904,N_15123,N_15598);
nand U15905 (N_15905,N_15424,N_15077);
nand U15906 (N_15906,N_15234,N_15148);
or U15907 (N_15907,N_15531,N_15438);
nor U15908 (N_15908,N_15507,N_15036);
and U15909 (N_15909,N_15355,N_15312);
and U15910 (N_15910,N_15527,N_15611);
nor U15911 (N_15911,N_15371,N_15539);
nand U15912 (N_15912,N_15080,N_15089);
nor U15913 (N_15913,N_15130,N_15207);
or U15914 (N_15914,N_15348,N_15013);
xor U15915 (N_15915,N_15134,N_15339);
or U15916 (N_15916,N_15420,N_15293);
nand U15917 (N_15917,N_15114,N_15037);
nand U15918 (N_15918,N_15498,N_15086);
nor U15919 (N_15919,N_15418,N_15458);
xnor U15920 (N_15920,N_15160,N_15580);
nor U15921 (N_15921,N_15146,N_15282);
xnor U15922 (N_15922,N_15190,N_15460);
nand U15923 (N_15923,N_15141,N_15357);
and U15924 (N_15924,N_15602,N_15264);
nand U15925 (N_15925,N_15096,N_15367);
xor U15926 (N_15926,N_15399,N_15002);
xnor U15927 (N_15927,N_15261,N_15470);
nand U15928 (N_15928,N_15622,N_15069);
nand U15929 (N_15929,N_15184,N_15109);
xor U15930 (N_15930,N_15401,N_15478);
nand U15931 (N_15931,N_15039,N_15396);
nand U15932 (N_15932,N_15459,N_15444);
and U15933 (N_15933,N_15338,N_15573);
xnor U15934 (N_15934,N_15132,N_15100);
nor U15935 (N_15935,N_15304,N_15279);
or U15936 (N_15936,N_15006,N_15476);
nand U15937 (N_15937,N_15528,N_15624);
xnor U15938 (N_15938,N_15086,N_15100);
or U15939 (N_15939,N_15304,N_15102);
xnor U15940 (N_15940,N_15317,N_15172);
or U15941 (N_15941,N_15122,N_15321);
nor U15942 (N_15942,N_15566,N_15393);
nand U15943 (N_15943,N_15557,N_15414);
xnor U15944 (N_15944,N_15169,N_15523);
and U15945 (N_15945,N_15084,N_15441);
or U15946 (N_15946,N_15028,N_15374);
nand U15947 (N_15947,N_15037,N_15094);
nand U15948 (N_15948,N_15122,N_15065);
nand U15949 (N_15949,N_15529,N_15541);
nor U15950 (N_15950,N_15030,N_15451);
nand U15951 (N_15951,N_15550,N_15266);
nand U15952 (N_15952,N_15603,N_15458);
or U15953 (N_15953,N_15446,N_15475);
xor U15954 (N_15954,N_15380,N_15572);
and U15955 (N_15955,N_15390,N_15584);
and U15956 (N_15956,N_15062,N_15519);
or U15957 (N_15957,N_15005,N_15370);
nand U15958 (N_15958,N_15367,N_15209);
nor U15959 (N_15959,N_15052,N_15519);
xnor U15960 (N_15960,N_15007,N_15463);
nand U15961 (N_15961,N_15501,N_15399);
and U15962 (N_15962,N_15405,N_15511);
and U15963 (N_15963,N_15029,N_15037);
nand U15964 (N_15964,N_15058,N_15408);
nor U15965 (N_15965,N_15238,N_15397);
nand U15966 (N_15966,N_15579,N_15465);
and U15967 (N_15967,N_15616,N_15211);
and U15968 (N_15968,N_15536,N_15013);
nor U15969 (N_15969,N_15231,N_15479);
and U15970 (N_15970,N_15089,N_15470);
xnor U15971 (N_15971,N_15532,N_15482);
nand U15972 (N_15972,N_15115,N_15541);
or U15973 (N_15973,N_15182,N_15268);
or U15974 (N_15974,N_15180,N_15066);
or U15975 (N_15975,N_15375,N_15154);
xor U15976 (N_15976,N_15400,N_15095);
nand U15977 (N_15977,N_15321,N_15474);
nand U15978 (N_15978,N_15555,N_15334);
or U15979 (N_15979,N_15001,N_15179);
or U15980 (N_15980,N_15111,N_15509);
and U15981 (N_15981,N_15443,N_15327);
or U15982 (N_15982,N_15341,N_15528);
nand U15983 (N_15983,N_15123,N_15125);
and U15984 (N_15984,N_15222,N_15439);
or U15985 (N_15985,N_15316,N_15452);
xnor U15986 (N_15986,N_15204,N_15315);
and U15987 (N_15987,N_15081,N_15426);
xnor U15988 (N_15988,N_15571,N_15465);
nor U15989 (N_15989,N_15052,N_15049);
or U15990 (N_15990,N_15214,N_15579);
xnor U15991 (N_15991,N_15478,N_15137);
nor U15992 (N_15992,N_15036,N_15443);
nand U15993 (N_15993,N_15295,N_15497);
and U15994 (N_15994,N_15172,N_15339);
nor U15995 (N_15995,N_15301,N_15106);
xnor U15996 (N_15996,N_15349,N_15604);
nor U15997 (N_15997,N_15095,N_15111);
xnor U15998 (N_15998,N_15404,N_15313);
xnor U15999 (N_15999,N_15613,N_15083);
and U16000 (N_16000,N_15348,N_15293);
nor U16001 (N_16001,N_15389,N_15192);
and U16002 (N_16002,N_15299,N_15153);
xnor U16003 (N_16003,N_15251,N_15367);
and U16004 (N_16004,N_15570,N_15372);
or U16005 (N_16005,N_15179,N_15216);
xnor U16006 (N_16006,N_15051,N_15497);
nor U16007 (N_16007,N_15361,N_15614);
or U16008 (N_16008,N_15576,N_15493);
xor U16009 (N_16009,N_15487,N_15171);
nor U16010 (N_16010,N_15241,N_15535);
and U16011 (N_16011,N_15422,N_15334);
and U16012 (N_16012,N_15248,N_15043);
nand U16013 (N_16013,N_15574,N_15429);
nand U16014 (N_16014,N_15614,N_15278);
xor U16015 (N_16015,N_15171,N_15048);
xnor U16016 (N_16016,N_15580,N_15561);
nor U16017 (N_16017,N_15566,N_15098);
xnor U16018 (N_16018,N_15504,N_15430);
and U16019 (N_16019,N_15037,N_15013);
and U16020 (N_16020,N_15034,N_15602);
and U16021 (N_16021,N_15029,N_15200);
or U16022 (N_16022,N_15128,N_15051);
nor U16023 (N_16023,N_15568,N_15173);
and U16024 (N_16024,N_15258,N_15414);
nor U16025 (N_16025,N_15360,N_15350);
xor U16026 (N_16026,N_15225,N_15600);
xor U16027 (N_16027,N_15364,N_15441);
xnor U16028 (N_16028,N_15320,N_15153);
xnor U16029 (N_16029,N_15271,N_15296);
xnor U16030 (N_16030,N_15330,N_15612);
and U16031 (N_16031,N_15353,N_15341);
nor U16032 (N_16032,N_15160,N_15342);
xor U16033 (N_16033,N_15187,N_15304);
nand U16034 (N_16034,N_15539,N_15353);
nand U16035 (N_16035,N_15410,N_15600);
nor U16036 (N_16036,N_15139,N_15288);
and U16037 (N_16037,N_15185,N_15179);
xor U16038 (N_16038,N_15562,N_15089);
xnor U16039 (N_16039,N_15353,N_15420);
xor U16040 (N_16040,N_15277,N_15128);
xor U16041 (N_16041,N_15564,N_15191);
or U16042 (N_16042,N_15505,N_15086);
nor U16043 (N_16043,N_15127,N_15106);
and U16044 (N_16044,N_15222,N_15556);
or U16045 (N_16045,N_15288,N_15360);
xor U16046 (N_16046,N_15409,N_15314);
nand U16047 (N_16047,N_15475,N_15577);
and U16048 (N_16048,N_15521,N_15443);
nor U16049 (N_16049,N_15307,N_15612);
nor U16050 (N_16050,N_15425,N_15445);
nand U16051 (N_16051,N_15436,N_15604);
xor U16052 (N_16052,N_15366,N_15118);
and U16053 (N_16053,N_15312,N_15328);
or U16054 (N_16054,N_15268,N_15118);
nor U16055 (N_16055,N_15578,N_15074);
xor U16056 (N_16056,N_15608,N_15437);
xor U16057 (N_16057,N_15274,N_15397);
and U16058 (N_16058,N_15457,N_15602);
or U16059 (N_16059,N_15615,N_15325);
and U16060 (N_16060,N_15418,N_15222);
or U16061 (N_16061,N_15391,N_15434);
nor U16062 (N_16062,N_15044,N_15366);
nor U16063 (N_16063,N_15154,N_15577);
or U16064 (N_16064,N_15285,N_15540);
nand U16065 (N_16065,N_15218,N_15451);
or U16066 (N_16066,N_15524,N_15082);
nor U16067 (N_16067,N_15485,N_15301);
xnor U16068 (N_16068,N_15033,N_15301);
or U16069 (N_16069,N_15192,N_15007);
nor U16070 (N_16070,N_15188,N_15179);
and U16071 (N_16071,N_15471,N_15124);
or U16072 (N_16072,N_15307,N_15158);
xnor U16073 (N_16073,N_15369,N_15550);
or U16074 (N_16074,N_15439,N_15265);
xor U16075 (N_16075,N_15132,N_15174);
xnor U16076 (N_16076,N_15527,N_15364);
and U16077 (N_16077,N_15498,N_15510);
and U16078 (N_16078,N_15530,N_15004);
nor U16079 (N_16079,N_15064,N_15136);
and U16080 (N_16080,N_15010,N_15623);
nor U16081 (N_16081,N_15579,N_15274);
xor U16082 (N_16082,N_15566,N_15172);
nand U16083 (N_16083,N_15130,N_15342);
or U16084 (N_16084,N_15067,N_15384);
and U16085 (N_16085,N_15209,N_15208);
or U16086 (N_16086,N_15481,N_15081);
or U16087 (N_16087,N_15016,N_15158);
xnor U16088 (N_16088,N_15006,N_15479);
xor U16089 (N_16089,N_15222,N_15207);
or U16090 (N_16090,N_15019,N_15190);
or U16091 (N_16091,N_15402,N_15462);
or U16092 (N_16092,N_15150,N_15158);
nand U16093 (N_16093,N_15565,N_15479);
nand U16094 (N_16094,N_15478,N_15139);
nand U16095 (N_16095,N_15501,N_15078);
and U16096 (N_16096,N_15600,N_15505);
and U16097 (N_16097,N_15218,N_15515);
xor U16098 (N_16098,N_15004,N_15195);
or U16099 (N_16099,N_15142,N_15469);
nor U16100 (N_16100,N_15602,N_15350);
xor U16101 (N_16101,N_15382,N_15410);
nand U16102 (N_16102,N_15069,N_15307);
nor U16103 (N_16103,N_15389,N_15330);
or U16104 (N_16104,N_15264,N_15020);
or U16105 (N_16105,N_15406,N_15108);
nor U16106 (N_16106,N_15421,N_15364);
nor U16107 (N_16107,N_15239,N_15387);
nor U16108 (N_16108,N_15413,N_15284);
or U16109 (N_16109,N_15416,N_15309);
xor U16110 (N_16110,N_15345,N_15513);
nand U16111 (N_16111,N_15282,N_15546);
and U16112 (N_16112,N_15479,N_15578);
or U16113 (N_16113,N_15515,N_15288);
or U16114 (N_16114,N_15049,N_15428);
xnor U16115 (N_16115,N_15339,N_15200);
nand U16116 (N_16116,N_15295,N_15504);
nand U16117 (N_16117,N_15383,N_15083);
and U16118 (N_16118,N_15425,N_15272);
or U16119 (N_16119,N_15312,N_15204);
xnor U16120 (N_16120,N_15511,N_15317);
nor U16121 (N_16121,N_15169,N_15109);
or U16122 (N_16122,N_15437,N_15533);
xnor U16123 (N_16123,N_15461,N_15145);
nor U16124 (N_16124,N_15592,N_15170);
or U16125 (N_16125,N_15345,N_15025);
xor U16126 (N_16126,N_15211,N_15366);
nand U16127 (N_16127,N_15285,N_15199);
xor U16128 (N_16128,N_15011,N_15127);
nand U16129 (N_16129,N_15117,N_15387);
nand U16130 (N_16130,N_15123,N_15199);
and U16131 (N_16131,N_15053,N_15076);
or U16132 (N_16132,N_15586,N_15421);
xor U16133 (N_16133,N_15399,N_15136);
or U16134 (N_16134,N_15376,N_15289);
and U16135 (N_16135,N_15210,N_15419);
or U16136 (N_16136,N_15026,N_15237);
xor U16137 (N_16137,N_15446,N_15077);
or U16138 (N_16138,N_15316,N_15128);
xor U16139 (N_16139,N_15137,N_15524);
nand U16140 (N_16140,N_15111,N_15551);
and U16141 (N_16141,N_15105,N_15429);
and U16142 (N_16142,N_15199,N_15128);
or U16143 (N_16143,N_15521,N_15065);
nor U16144 (N_16144,N_15045,N_15011);
and U16145 (N_16145,N_15023,N_15078);
and U16146 (N_16146,N_15190,N_15433);
nand U16147 (N_16147,N_15593,N_15239);
nand U16148 (N_16148,N_15533,N_15209);
nand U16149 (N_16149,N_15251,N_15579);
xor U16150 (N_16150,N_15020,N_15565);
nor U16151 (N_16151,N_15190,N_15081);
xnor U16152 (N_16152,N_15459,N_15411);
nor U16153 (N_16153,N_15488,N_15468);
and U16154 (N_16154,N_15043,N_15546);
xor U16155 (N_16155,N_15234,N_15492);
nor U16156 (N_16156,N_15507,N_15486);
and U16157 (N_16157,N_15198,N_15584);
and U16158 (N_16158,N_15059,N_15616);
nand U16159 (N_16159,N_15285,N_15216);
and U16160 (N_16160,N_15347,N_15241);
and U16161 (N_16161,N_15456,N_15619);
nand U16162 (N_16162,N_15137,N_15127);
nor U16163 (N_16163,N_15535,N_15490);
xor U16164 (N_16164,N_15097,N_15374);
or U16165 (N_16165,N_15468,N_15028);
or U16166 (N_16166,N_15224,N_15354);
or U16167 (N_16167,N_15532,N_15084);
xnor U16168 (N_16168,N_15325,N_15173);
xor U16169 (N_16169,N_15505,N_15552);
or U16170 (N_16170,N_15567,N_15008);
xor U16171 (N_16171,N_15193,N_15057);
or U16172 (N_16172,N_15183,N_15388);
or U16173 (N_16173,N_15575,N_15449);
or U16174 (N_16174,N_15148,N_15223);
or U16175 (N_16175,N_15305,N_15510);
or U16176 (N_16176,N_15310,N_15196);
and U16177 (N_16177,N_15242,N_15216);
nand U16178 (N_16178,N_15185,N_15093);
nand U16179 (N_16179,N_15327,N_15253);
nand U16180 (N_16180,N_15276,N_15264);
and U16181 (N_16181,N_15389,N_15493);
xor U16182 (N_16182,N_15156,N_15034);
xnor U16183 (N_16183,N_15506,N_15510);
nor U16184 (N_16184,N_15392,N_15203);
nand U16185 (N_16185,N_15351,N_15303);
nor U16186 (N_16186,N_15060,N_15360);
or U16187 (N_16187,N_15605,N_15159);
nor U16188 (N_16188,N_15156,N_15570);
or U16189 (N_16189,N_15338,N_15172);
or U16190 (N_16190,N_15558,N_15136);
xnor U16191 (N_16191,N_15511,N_15589);
or U16192 (N_16192,N_15077,N_15540);
nor U16193 (N_16193,N_15240,N_15216);
nand U16194 (N_16194,N_15169,N_15083);
and U16195 (N_16195,N_15064,N_15409);
xnor U16196 (N_16196,N_15062,N_15487);
xnor U16197 (N_16197,N_15256,N_15054);
xor U16198 (N_16198,N_15046,N_15578);
xor U16199 (N_16199,N_15253,N_15196);
or U16200 (N_16200,N_15001,N_15190);
xor U16201 (N_16201,N_15240,N_15357);
and U16202 (N_16202,N_15285,N_15103);
or U16203 (N_16203,N_15602,N_15423);
or U16204 (N_16204,N_15073,N_15029);
nor U16205 (N_16205,N_15486,N_15318);
nand U16206 (N_16206,N_15144,N_15461);
or U16207 (N_16207,N_15295,N_15058);
nor U16208 (N_16208,N_15407,N_15223);
nand U16209 (N_16209,N_15526,N_15330);
or U16210 (N_16210,N_15535,N_15099);
xnor U16211 (N_16211,N_15554,N_15292);
and U16212 (N_16212,N_15393,N_15251);
nand U16213 (N_16213,N_15621,N_15174);
or U16214 (N_16214,N_15523,N_15571);
nand U16215 (N_16215,N_15136,N_15077);
and U16216 (N_16216,N_15613,N_15450);
and U16217 (N_16217,N_15518,N_15345);
or U16218 (N_16218,N_15171,N_15009);
or U16219 (N_16219,N_15237,N_15421);
xnor U16220 (N_16220,N_15261,N_15378);
or U16221 (N_16221,N_15132,N_15041);
or U16222 (N_16222,N_15274,N_15432);
xnor U16223 (N_16223,N_15260,N_15145);
xnor U16224 (N_16224,N_15170,N_15519);
nor U16225 (N_16225,N_15548,N_15210);
or U16226 (N_16226,N_15516,N_15318);
nor U16227 (N_16227,N_15403,N_15394);
xor U16228 (N_16228,N_15532,N_15242);
nand U16229 (N_16229,N_15480,N_15183);
nor U16230 (N_16230,N_15449,N_15619);
and U16231 (N_16231,N_15177,N_15615);
xnor U16232 (N_16232,N_15099,N_15437);
xor U16233 (N_16233,N_15457,N_15216);
or U16234 (N_16234,N_15087,N_15576);
or U16235 (N_16235,N_15004,N_15016);
xnor U16236 (N_16236,N_15254,N_15412);
and U16237 (N_16237,N_15214,N_15194);
or U16238 (N_16238,N_15088,N_15261);
nand U16239 (N_16239,N_15094,N_15124);
nand U16240 (N_16240,N_15301,N_15193);
xor U16241 (N_16241,N_15472,N_15145);
xnor U16242 (N_16242,N_15498,N_15499);
and U16243 (N_16243,N_15519,N_15404);
and U16244 (N_16244,N_15479,N_15158);
nor U16245 (N_16245,N_15396,N_15584);
and U16246 (N_16246,N_15368,N_15439);
nor U16247 (N_16247,N_15542,N_15318);
xnor U16248 (N_16248,N_15189,N_15384);
xor U16249 (N_16249,N_15593,N_15540);
nand U16250 (N_16250,N_15704,N_15715);
xnor U16251 (N_16251,N_15727,N_16110);
and U16252 (N_16252,N_15854,N_15833);
xor U16253 (N_16253,N_16175,N_15733);
nor U16254 (N_16254,N_16040,N_16094);
nand U16255 (N_16255,N_15716,N_16112);
and U16256 (N_16256,N_15776,N_15708);
and U16257 (N_16257,N_15674,N_15763);
xnor U16258 (N_16258,N_15686,N_16236);
nand U16259 (N_16259,N_15948,N_16188);
nand U16260 (N_16260,N_15749,N_16027);
or U16261 (N_16261,N_15880,N_15933);
or U16262 (N_16262,N_15697,N_15847);
or U16263 (N_16263,N_16105,N_15921);
xor U16264 (N_16264,N_15844,N_16136);
nor U16265 (N_16265,N_16121,N_16157);
and U16266 (N_16266,N_15789,N_16051);
xor U16267 (N_16267,N_16178,N_16182);
xnor U16268 (N_16268,N_15748,N_16088);
nor U16269 (N_16269,N_16035,N_16099);
nand U16270 (N_16270,N_16216,N_15871);
and U16271 (N_16271,N_15744,N_15852);
xnor U16272 (N_16272,N_16210,N_15754);
and U16273 (N_16273,N_16108,N_16229);
xnor U16274 (N_16274,N_16010,N_15953);
or U16275 (N_16275,N_16167,N_16185);
nor U16276 (N_16276,N_15839,N_16041);
nor U16277 (N_16277,N_15809,N_16195);
nor U16278 (N_16278,N_16119,N_15894);
nand U16279 (N_16279,N_16064,N_16181);
xnor U16280 (N_16280,N_15978,N_15658);
nand U16281 (N_16281,N_16179,N_15807);
xnor U16282 (N_16282,N_16173,N_15627);
nor U16283 (N_16283,N_16084,N_15856);
xor U16284 (N_16284,N_15737,N_15756);
xnor U16285 (N_16285,N_16044,N_15974);
and U16286 (N_16286,N_16004,N_16144);
and U16287 (N_16287,N_15814,N_15739);
nor U16288 (N_16288,N_15977,N_15904);
and U16289 (N_16289,N_16221,N_16159);
or U16290 (N_16290,N_16102,N_15734);
or U16291 (N_16291,N_16196,N_15677);
nor U16292 (N_16292,N_16039,N_16218);
or U16293 (N_16293,N_15946,N_15652);
nor U16294 (N_16294,N_15960,N_16097);
or U16295 (N_16295,N_15730,N_15656);
nand U16296 (N_16296,N_15801,N_15817);
or U16297 (N_16297,N_16042,N_16015);
nor U16298 (N_16298,N_15812,N_15689);
xor U16299 (N_16299,N_15701,N_15661);
nor U16300 (N_16300,N_16202,N_16007);
or U16301 (N_16301,N_15911,N_15797);
xnor U16302 (N_16302,N_15944,N_15965);
xnor U16303 (N_16303,N_15855,N_15712);
and U16304 (N_16304,N_15806,N_15980);
nor U16305 (N_16305,N_15741,N_15825);
nor U16306 (N_16306,N_15631,N_15897);
nor U16307 (N_16307,N_15872,N_16036);
or U16308 (N_16308,N_16057,N_16049);
nor U16309 (N_16309,N_15875,N_16190);
nand U16310 (N_16310,N_15784,N_16245);
xor U16311 (N_16311,N_15829,N_15939);
xnor U16312 (N_16312,N_15992,N_15673);
nor U16313 (N_16313,N_15775,N_16000);
and U16314 (N_16314,N_15705,N_15752);
xor U16315 (N_16315,N_15821,N_16061);
nor U16316 (N_16316,N_15832,N_15930);
and U16317 (N_16317,N_16138,N_15934);
and U16318 (N_16318,N_16031,N_15685);
and U16319 (N_16319,N_16169,N_16212);
or U16320 (N_16320,N_16087,N_16028);
or U16321 (N_16321,N_15907,N_15771);
xor U16322 (N_16322,N_16063,N_15638);
nor U16323 (N_16323,N_16209,N_16006);
xnor U16324 (N_16324,N_15909,N_16075);
nand U16325 (N_16325,N_16106,N_16111);
nor U16326 (N_16326,N_15700,N_15867);
xor U16327 (N_16327,N_16052,N_15824);
or U16328 (N_16328,N_16226,N_16002);
nand U16329 (N_16329,N_15710,N_16153);
nand U16330 (N_16330,N_15850,N_15794);
nand U16331 (N_16331,N_16020,N_15728);
xor U16332 (N_16332,N_16001,N_16215);
nor U16333 (N_16333,N_16205,N_16095);
xnor U16334 (N_16334,N_15740,N_15684);
or U16335 (N_16335,N_15866,N_16204);
nor U16336 (N_16336,N_15681,N_16140);
nand U16337 (N_16337,N_15757,N_16082);
nand U16338 (N_16338,N_16141,N_16053);
nor U16339 (N_16339,N_16171,N_16032);
and U16340 (N_16340,N_16076,N_15888);
nor U16341 (N_16341,N_15891,N_16176);
and U16342 (N_16342,N_15780,N_15896);
nor U16343 (N_16343,N_15670,N_15663);
xnor U16344 (N_16344,N_15859,N_16223);
xor U16345 (N_16345,N_15901,N_15922);
and U16346 (N_16346,N_15947,N_16071);
and U16347 (N_16347,N_15800,N_16249);
nor U16348 (N_16348,N_15957,N_15840);
or U16349 (N_16349,N_16241,N_15761);
xor U16350 (N_16350,N_16239,N_16164);
and U16351 (N_16351,N_16243,N_15906);
xor U16352 (N_16352,N_16078,N_15795);
xnor U16353 (N_16353,N_16127,N_16101);
or U16354 (N_16354,N_15869,N_15952);
and U16355 (N_16355,N_16151,N_15975);
nor U16356 (N_16356,N_16107,N_16191);
nor U16357 (N_16357,N_16069,N_15818);
and U16358 (N_16358,N_15815,N_15675);
nor U16359 (N_16359,N_15945,N_15767);
and U16360 (N_16360,N_15713,N_15924);
nand U16361 (N_16361,N_16056,N_16012);
or U16362 (N_16362,N_16149,N_15643);
nor U16363 (N_16363,N_15903,N_16129);
nand U16364 (N_16364,N_16005,N_15830);
and U16365 (N_16365,N_16174,N_15936);
xor U16366 (N_16366,N_15654,N_15963);
nand U16367 (N_16367,N_16059,N_16026);
nor U16368 (N_16368,N_15991,N_15885);
nor U16369 (N_16369,N_15826,N_16100);
and U16370 (N_16370,N_15802,N_16222);
xor U16371 (N_16371,N_16208,N_15692);
or U16372 (N_16372,N_15782,N_15861);
xor U16373 (N_16373,N_16065,N_16085);
nor U16374 (N_16374,N_16183,N_15942);
nand U16375 (N_16375,N_16003,N_15785);
nand U16376 (N_16376,N_15647,N_15923);
and U16377 (N_16377,N_15683,N_15706);
or U16378 (N_16378,N_16091,N_15990);
or U16379 (N_16379,N_15941,N_15786);
nor U16380 (N_16380,N_16192,N_15864);
nand U16381 (N_16381,N_15926,N_15645);
xor U16382 (N_16382,N_15770,N_16077);
nand U16383 (N_16383,N_16023,N_16083);
nand U16384 (N_16384,N_16067,N_15717);
nand U16385 (N_16385,N_16139,N_15849);
xor U16386 (N_16386,N_15696,N_15816);
nand U16387 (N_16387,N_16013,N_16214);
and U16388 (N_16388,N_16156,N_15790);
and U16389 (N_16389,N_15777,N_16206);
nor U16390 (N_16390,N_16184,N_15639);
or U16391 (N_16391,N_16131,N_15759);
and U16392 (N_16392,N_15862,N_15900);
nor U16393 (N_16393,N_16201,N_15693);
nor U16394 (N_16394,N_15707,N_15913);
xnor U16395 (N_16395,N_16019,N_15860);
and U16396 (N_16396,N_15640,N_15884);
nor U16397 (N_16397,N_15838,N_16117);
xor U16398 (N_16398,N_15822,N_16120);
or U16399 (N_16399,N_15938,N_16114);
nor U16400 (N_16400,N_16034,N_15986);
nor U16401 (N_16401,N_15653,N_16062);
xor U16402 (N_16402,N_16038,N_16021);
nor U16403 (N_16403,N_15742,N_16242);
nor U16404 (N_16404,N_15961,N_15720);
nor U16405 (N_16405,N_16194,N_15955);
nand U16406 (N_16406,N_15718,N_16207);
nor U16407 (N_16407,N_15778,N_15917);
nor U16408 (N_16408,N_15949,N_15711);
and U16409 (N_16409,N_16103,N_15665);
or U16410 (N_16410,N_15971,N_15798);
and U16411 (N_16411,N_16160,N_15695);
or U16412 (N_16412,N_15803,N_15820);
and U16413 (N_16413,N_15646,N_16022);
nor U16414 (N_16414,N_15632,N_16043);
or U16415 (N_16415,N_16066,N_15687);
nor U16416 (N_16416,N_16161,N_15962);
nand U16417 (N_16417,N_15732,N_15726);
xnor U16418 (N_16418,N_15811,N_16168);
and U16419 (N_16419,N_15679,N_15671);
nor U16420 (N_16420,N_15912,N_15808);
nand U16421 (N_16421,N_16247,N_15951);
or U16422 (N_16422,N_16096,N_15662);
xor U16423 (N_16423,N_15743,N_15878);
or U16424 (N_16424,N_15877,N_15976);
xor U16425 (N_16425,N_16165,N_16033);
xnor U16426 (N_16426,N_16074,N_16118);
xor U16427 (N_16427,N_16073,N_15845);
and U16428 (N_16428,N_15981,N_15625);
xor U16429 (N_16429,N_16092,N_15998);
and U16430 (N_16430,N_15967,N_16227);
nand U16431 (N_16431,N_15937,N_15731);
nor U16432 (N_16432,N_16220,N_15724);
nor U16433 (N_16433,N_16014,N_15905);
and U16434 (N_16434,N_16130,N_15642);
xor U16435 (N_16435,N_16152,N_15881);
nor U16436 (N_16436,N_15870,N_15753);
nor U16437 (N_16437,N_15667,N_15769);
xor U16438 (N_16438,N_15851,N_16011);
nand U16439 (N_16439,N_16234,N_15766);
xnor U16440 (N_16440,N_16050,N_15659);
or U16441 (N_16441,N_16081,N_16128);
nor U16442 (N_16442,N_15651,N_16232);
nor U16443 (N_16443,N_16186,N_15982);
or U16444 (N_16444,N_15865,N_16045);
or U16445 (N_16445,N_15846,N_16104);
nor U16446 (N_16446,N_15672,N_16070);
and U16447 (N_16447,N_15993,N_16122);
xor U16448 (N_16448,N_15630,N_15968);
xor U16449 (N_16449,N_16172,N_15994);
and U16450 (N_16450,N_16046,N_15764);
xnor U16451 (N_16451,N_16158,N_16155);
xor U16452 (N_16452,N_15755,N_15823);
and U16453 (N_16453,N_15781,N_15956);
nand U16454 (N_16454,N_16029,N_15751);
nand U16455 (N_16455,N_15902,N_15633);
nor U16456 (N_16456,N_15736,N_15792);
xnor U16457 (N_16457,N_15669,N_16123);
nor U16458 (N_16458,N_16219,N_15635);
nand U16459 (N_16459,N_16008,N_16217);
or U16460 (N_16460,N_15799,N_15834);
nand U16461 (N_16461,N_15779,N_16170);
or U16462 (N_16462,N_16054,N_15721);
or U16463 (N_16463,N_15626,N_15893);
or U16464 (N_16464,N_16133,N_16132);
xnor U16465 (N_16465,N_15837,N_15719);
nand U16466 (N_16466,N_15868,N_15762);
and U16467 (N_16467,N_16142,N_15698);
xnor U16468 (N_16468,N_15848,N_16124);
nand U16469 (N_16469,N_15882,N_15746);
and U16470 (N_16470,N_16233,N_15649);
xor U16471 (N_16471,N_15887,N_15788);
xnor U16472 (N_16472,N_15666,N_15995);
nor U16473 (N_16473,N_15931,N_15916);
xor U16474 (N_16474,N_16089,N_15898);
nand U16475 (N_16475,N_15908,N_15929);
xnor U16476 (N_16476,N_16193,N_16009);
nor U16477 (N_16477,N_16072,N_16163);
and U16478 (N_16478,N_16187,N_15804);
or U16479 (N_16479,N_16109,N_15973);
nor U16480 (N_16480,N_16150,N_15835);
and U16481 (N_16481,N_16199,N_15932);
nor U16482 (N_16482,N_15954,N_15876);
xor U16483 (N_16483,N_15950,N_15983);
and U16484 (N_16484,N_16248,N_16162);
nor U16485 (N_16485,N_16225,N_15783);
and U16486 (N_16486,N_16017,N_15879);
and U16487 (N_16487,N_15873,N_15919);
or U16488 (N_16488,N_15972,N_15883);
nand U16489 (N_16489,N_15765,N_15690);
nor U16490 (N_16490,N_15745,N_16115);
xnor U16491 (N_16491,N_16025,N_15676);
nor U16492 (N_16492,N_16198,N_15958);
or U16493 (N_16493,N_16180,N_15680);
and U16494 (N_16494,N_16211,N_16228);
xor U16495 (N_16495,N_15940,N_15858);
nor U16496 (N_16496,N_15655,N_15996);
and U16497 (N_16497,N_15819,N_15969);
nand U16498 (N_16498,N_15747,N_15691);
or U16499 (N_16499,N_15889,N_15703);
xnor U16500 (N_16500,N_15979,N_15644);
or U16501 (N_16501,N_15637,N_15660);
nor U16502 (N_16502,N_16098,N_15657);
or U16503 (N_16503,N_16018,N_15629);
xnor U16504 (N_16504,N_16030,N_16024);
nand U16505 (N_16505,N_15970,N_15964);
nand U16506 (N_16506,N_15828,N_15628);
nand U16507 (N_16507,N_15650,N_16135);
or U16508 (N_16508,N_15925,N_15668);
or U16509 (N_16509,N_15805,N_15714);
nand U16510 (N_16510,N_15648,N_16224);
xor U16511 (N_16511,N_15920,N_16055);
nand U16512 (N_16512,N_15989,N_15895);
xnor U16513 (N_16513,N_16086,N_15738);
and U16514 (N_16514,N_15966,N_16189);
nor U16515 (N_16515,N_16240,N_16203);
xnor U16516 (N_16516,N_16137,N_15999);
nor U16517 (N_16517,N_15723,N_15943);
and U16518 (N_16518,N_15773,N_15664);
nand U16519 (N_16519,N_15796,N_16200);
nor U16520 (N_16520,N_16093,N_15699);
xor U16521 (N_16521,N_15910,N_15694);
nor U16522 (N_16522,N_15793,N_16048);
or U16523 (N_16523,N_16079,N_15750);
or U16524 (N_16524,N_15890,N_16238);
nor U16525 (N_16525,N_16090,N_15915);
nand U16526 (N_16526,N_15857,N_15702);
nand U16527 (N_16527,N_15843,N_15641);
nor U16528 (N_16528,N_15688,N_15886);
and U16529 (N_16529,N_16197,N_16231);
nor U16530 (N_16530,N_16166,N_15831);
or U16531 (N_16531,N_16235,N_15935);
nor U16532 (N_16532,N_15827,N_15959);
xor U16533 (N_16533,N_15787,N_16125);
or U16534 (N_16534,N_15634,N_16047);
nor U16535 (N_16535,N_16113,N_15841);
nor U16536 (N_16536,N_15853,N_15874);
nand U16537 (N_16537,N_15774,N_15928);
nand U16538 (N_16538,N_16145,N_16080);
nand U16539 (N_16539,N_15772,N_15636);
xnor U16540 (N_16540,N_16237,N_15987);
nor U16541 (N_16541,N_15918,N_15813);
or U16542 (N_16542,N_15914,N_15892);
and U16543 (N_16543,N_15682,N_16154);
nand U16544 (N_16544,N_15836,N_16148);
nand U16545 (N_16545,N_16146,N_16230);
and U16546 (N_16546,N_15722,N_16058);
nand U16547 (N_16547,N_15729,N_15984);
nor U16548 (N_16548,N_15927,N_15768);
nor U16549 (N_16549,N_15899,N_16116);
xor U16550 (N_16550,N_15997,N_15985);
xnor U16551 (N_16551,N_15842,N_15758);
and U16552 (N_16552,N_16037,N_15791);
nor U16553 (N_16553,N_15725,N_16244);
nand U16554 (N_16554,N_15810,N_16177);
nand U16555 (N_16555,N_16143,N_15988);
nand U16556 (N_16556,N_16246,N_16126);
xor U16557 (N_16557,N_16016,N_15678);
and U16558 (N_16558,N_16213,N_16068);
and U16559 (N_16559,N_16147,N_16060);
xor U16560 (N_16560,N_15863,N_15709);
and U16561 (N_16561,N_16134,N_15735);
xor U16562 (N_16562,N_15760,N_15953);
nand U16563 (N_16563,N_15714,N_15666);
and U16564 (N_16564,N_16188,N_16055);
xnor U16565 (N_16565,N_16139,N_15658);
and U16566 (N_16566,N_16230,N_16080);
and U16567 (N_16567,N_15636,N_15860);
xor U16568 (N_16568,N_16090,N_16007);
and U16569 (N_16569,N_16013,N_16244);
and U16570 (N_16570,N_16022,N_15783);
xnor U16571 (N_16571,N_15718,N_15746);
and U16572 (N_16572,N_16171,N_15879);
xor U16573 (N_16573,N_15656,N_15735);
nand U16574 (N_16574,N_15774,N_16144);
nand U16575 (N_16575,N_15923,N_15896);
and U16576 (N_16576,N_15999,N_16028);
and U16577 (N_16577,N_15692,N_16059);
nor U16578 (N_16578,N_16170,N_15688);
nand U16579 (N_16579,N_15636,N_15683);
or U16580 (N_16580,N_15923,N_15707);
nand U16581 (N_16581,N_15940,N_15765);
nand U16582 (N_16582,N_16184,N_15919);
xor U16583 (N_16583,N_15755,N_16106);
nand U16584 (N_16584,N_16171,N_16204);
nor U16585 (N_16585,N_16020,N_15792);
or U16586 (N_16586,N_16154,N_16095);
or U16587 (N_16587,N_15686,N_16242);
or U16588 (N_16588,N_16194,N_16186);
xor U16589 (N_16589,N_15957,N_15694);
nand U16590 (N_16590,N_15978,N_15888);
or U16591 (N_16591,N_15970,N_16046);
and U16592 (N_16592,N_16161,N_15783);
or U16593 (N_16593,N_15768,N_15733);
nand U16594 (N_16594,N_16015,N_16016);
and U16595 (N_16595,N_15732,N_16044);
xor U16596 (N_16596,N_15674,N_15950);
or U16597 (N_16597,N_16002,N_15954);
or U16598 (N_16598,N_15828,N_16014);
nor U16599 (N_16599,N_15748,N_15673);
xnor U16600 (N_16600,N_16037,N_15994);
nor U16601 (N_16601,N_15834,N_15808);
nor U16602 (N_16602,N_15818,N_15913);
or U16603 (N_16603,N_16248,N_15968);
nand U16604 (N_16604,N_15910,N_15828);
nor U16605 (N_16605,N_16213,N_16243);
and U16606 (N_16606,N_15968,N_16243);
or U16607 (N_16607,N_16124,N_16247);
or U16608 (N_16608,N_16161,N_15817);
nand U16609 (N_16609,N_16066,N_15733);
or U16610 (N_16610,N_16034,N_16213);
xor U16611 (N_16611,N_16084,N_15632);
and U16612 (N_16612,N_16038,N_16049);
nor U16613 (N_16613,N_15652,N_16112);
or U16614 (N_16614,N_16041,N_15683);
nand U16615 (N_16615,N_16102,N_16172);
or U16616 (N_16616,N_15865,N_15805);
nand U16617 (N_16617,N_16145,N_16037);
nor U16618 (N_16618,N_16092,N_15837);
nand U16619 (N_16619,N_15653,N_15797);
nand U16620 (N_16620,N_15984,N_15665);
or U16621 (N_16621,N_16031,N_15672);
nor U16622 (N_16622,N_15952,N_15873);
nor U16623 (N_16623,N_15726,N_15759);
nand U16624 (N_16624,N_15649,N_16047);
nor U16625 (N_16625,N_16133,N_15930);
and U16626 (N_16626,N_15633,N_16043);
xor U16627 (N_16627,N_15870,N_16033);
nor U16628 (N_16628,N_16040,N_15722);
or U16629 (N_16629,N_15969,N_15893);
or U16630 (N_16630,N_16051,N_16205);
and U16631 (N_16631,N_16023,N_16183);
xnor U16632 (N_16632,N_16004,N_15858);
or U16633 (N_16633,N_15910,N_16202);
nor U16634 (N_16634,N_15645,N_15712);
nor U16635 (N_16635,N_16145,N_15759);
and U16636 (N_16636,N_16162,N_16031);
nor U16637 (N_16637,N_16142,N_16000);
nand U16638 (N_16638,N_15695,N_16200);
and U16639 (N_16639,N_16166,N_15670);
xnor U16640 (N_16640,N_15780,N_16110);
nor U16641 (N_16641,N_16113,N_16225);
nand U16642 (N_16642,N_15989,N_15710);
nor U16643 (N_16643,N_15656,N_16183);
and U16644 (N_16644,N_15874,N_15977);
xor U16645 (N_16645,N_15712,N_16165);
and U16646 (N_16646,N_15658,N_16042);
and U16647 (N_16647,N_15680,N_15991);
nor U16648 (N_16648,N_15919,N_16219);
nand U16649 (N_16649,N_16227,N_15700);
or U16650 (N_16650,N_16031,N_15859);
or U16651 (N_16651,N_16194,N_16115);
nand U16652 (N_16652,N_16045,N_16024);
and U16653 (N_16653,N_15928,N_15838);
nor U16654 (N_16654,N_16053,N_15770);
xor U16655 (N_16655,N_16085,N_16049);
and U16656 (N_16656,N_16197,N_15965);
nor U16657 (N_16657,N_15786,N_16057);
and U16658 (N_16658,N_15732,N_15693);
and U16659 (N_16659,N_15804,N_15770);
xor U16660 (N_16660,N_16212,N_16028);
or U16661 (N_16661,N_15670,N_15743);
xnor U16662 (N_16662,N_16005,N_16127);
nand U16663 (N_16663,N_15691,N_15744);
nand U16664 (N_16664,N_15697,N_16156);
or U16665 (N_16665,N_15686,N_15680);
nor U16666 (N_16666,N_15852,N_16215);
and U16667 (N_16667,N_15962,N_16082);
or U16668 (N_16668,N_16086,N_16020);
and U16669 (N_16669,N_15986,N_16030);
nor U16670 (N_16670,N_16005,N_16032);
and U16671 (N_16671,N_16160,N_16132);
or U16672 (N_16672,N_15731,N_16173);
or U16673 (N_16673,N_16141,N_15833);
nand U16674 (N_16674,N_16021,N_15830);
or U16675 (N_16675,N_16198,N_15693);
and U16676 (N_16676,N_15780,N_15753);
and U16677 (N_16677,N_15796,N_16169);
and U16678 (N_16678,N_15951,N_16087);
or U16679 (N_16679,N_15877,N_15918);
and U16680 (N_16680,N_16022,N_15664);
nor U16681 (N_16681,N_15865,N_16107);
xnor U16682 (N_16682,N_15625,N_16161);
or U16683 (N_16683,N_16069,N_16080);
or U16684 (N_16684,N_16183,N_15922);
xnor U16685 (N_16685,N_16206,N_16122);
nand U16686 (N_16686,N_15688,N_15888);
nor U16687 (N_16687,N_15955,N_16221);
nand U16688 (N_16688,N_15916,N_15848);
nand U16689 (N_16689,N_15853,N_16232);
and U16690 (N_16690,N_15818,N_15729);
nor U16691 (N_16691,N_15947,N_16025);
nor U16692 (N_16692,N_15668,N_15722);
or U16693 (N_16693,N_15986,N_15936);
or U16694 (N_16694,N_16075,N_15716);
nor U16695 (N_16695,N_15663,N_15989);
and U16696 (N_16696,N_15912,N_15640);
and U16697 (N_16697,N_15927,N_16216);
nand U16698 (N_16698,N_15947,N_16085);
or U16699 (N_16699,N_16225,N_15713);
and U16700 (N_16700,N_16167,N_16130);
nor U16701 (N_16701,N_15739,N_15974);
nand U16702 (N_16702,N_15806,N_15901);
xor U16703 (N_16703,N_15896,N_16242);
or U16704 (N_16704,N_16143,N_16066);
nand U16705 (N_16705,N_16197,N_16009);
xor U16706 (N_16706,N_16050,N_15958);
and U16707 (N_16707,N_16028,N_15836);
nand U16708 (N_16708,N_15949,N_15645);
xnor U16709 (N_16709,N_16118,N_16148);
or U16710 (N_16710,N_16081,N_16206);
xnor U16711 (N_16711,N_16226,N_15905);
nor U16712 (N_16712,N_16234,N_16114);
nor U16713 (N_16713,N_16028,N_16057);
or U16714 (N_16714,N_15852,N_15807);
nor U16715 (N_16715,N_15768,N_16140);
nor U16716 (N_16716,N_15698,N_15682);
and U16717 (N_16717,N_16160,N_15828);
xor U16718 (N_16718,N_15996,N_15808);
nand U16719 (N_16719,N_16071,N_16105);
nor U16720 (N_16720,N_15975,N_15631);
or U16721 (N_16721,N_15671,N_16102);
xor U16722 (N_16722,N_15658,N_16039);
nor U16723 (N_16723,N_16132,N_16073);
xor U16724 (N_16724,N_16043,N_16128);
nor U16725 (N_16725,N_15907,N_16050);
and U16726 (N_16726,N_15861,N_16237);
and U16727 (N_16727,N_15934,N_15740);
or U16728 (N_16728,N_16011,N_15642);
or U16729 (N_16729,N_16020,N_15884);
and U16730 (N_16730,N_16131,N_16205);
nor U16731 (N_16731,N_15900,N_15845);
and U16732 (N_16732,N_16062,N_15853);
xnor U16733 (N_16733,N_15765,N_16188);
or U16734 (N_16734,N_16208,N_15847);
xor U16735 (N_16735,N_15702,N_16190);
xor U16736 (N_16736,N_15675,N_16168);
nor U16737 (N_16737,N_16009,N_15920);
or U16738 (N_16738,N_15754,N_16188);
nor U16739 (N_16739,N_15693,N_15789);
xor U16740 (N_16740,N_15691,N_16087);
and U16741 (N_16741,N_16040,N_15823);
xnor U16742 (N_16742,N_15808,N_15767);
or U16743 (N_16743,N_16179,N_16229);
xor U16744 (N_16744,N_16195,N_15905);
nand U16745 (N_16745,N_16200,N_16211);
nor U16746 (N_16746,N_16031,N_15908);
or U16747 (N_16747,N_15770,N_15856);
nor U16748 (N_16748,N_15825,N_16146);
and U16749 (N_16749,N_15965,N_16168);
nand U16750 (N_16750,N_15820,N_15728);
nor U16751 (N_16751,N_15789,N_15634);
nand U16752 (N_16752,N_16082,N_16054);
nand U16753 (N_16753,N_16047,N_15911);
xnor U16754 (N_16754,N_15791,N_15981);
xnor U16755 (N_16755,N_16089,N_16204);
nor U16756 (N_16756,N_15972,N_15965);
or U16757 (N_16757,N_15706,N_15809);
nand U16758 (N_16758,N_15963,N_15877);
nor U16759 (N_16759,N_15965,N_16201);
nor U16760 (N_16760,N_16180,N_16137);
or U16761 (N_16761,N_16150,N_15964);
xor U16762 (N_16762,N_15805,N_16194);
nand U16763 (N_16763,N_15793,N_16015);
nand U16764 (N_16764,N_16060,N_15930);
nor U16765 (N_16765,N_15929,N_15803);
nand U16766 (N_16766,N_15635,N_16245);
xor U16767 (N_16767,N_16233,N_16042);
nor U16768 (N_16768,N_15978,N_16164);
nand U16769 (N_16769,N_16172,N_15637);
xor U16770 (N_16770,N_16158,N_15827);
or U16771 (N_16771,N_16070,N_15711);
and U16772 (N_16772,N_15724,N_16166);
xnor U16773 (N_16773,N_16243,N_16228);
and U16774 (N_16774,N_16010,N_15820);
nor U16775 (N_16775,N_16109,N_15901);
or U16776 (N_16776,N_16111,N_15984);
nand U16777 (N_16777,N_15892,N_15860);
or U16778 (N_16778,N_15662,N_15729);
nor U16779 (N_16779,N_16172,N_15950);
and U16780 (N_16780,N_15708,N_16025);
nor U16781 (N_16781,N_15877,N_15957);
nor U16782 (N_16782,N_15843,N_16140);
and U16783 (N_16783,N_16064,N_16069);
and U16784 (N_16784,N_15825,N_15908);
and U16785 (N_16785,N_16092,N_16183);
and U16786 (N_16786,N_15929,N_16145);
or U16787 (N_16787,N_15684,N_15950);
or U16788 (N_16788,N_16164,N_16234);
nand U16789 (N_16789,N_15963,N_15959);
or U16790 (N_16790,N_16212,N_16211);
xor U16791 (N_16791,N_15904,N_16197);
nor U16792 (N_16792,N_16209,N_15676);
xor U16793 (N_16793,N_15707,N_15636);
or U16794 (N_16794,N_16008,N_15666);
xnor U16795 (N_16795,N_15987,N_16056);
nand U16796 (N_16796,N_16066,N_15819);
or U16797 (N_16797,N_15944,N_16171);
nand U16798 (N_16798,N_15915,N_15771);
xnor U16799 (N_16799,N_15789,N_16099);
nand U16800 (N_16800,N_15986,N_16023);
nand U16801 (N_16801,N_15850,N_16134);
nand U16802 (N_16802,N_16239,N_16135);
and U16803 (N_16803,N_15890,N_15769);
or U16804 (N_16804,N_15682,N_15838);
and U16805 (N_16805,N_15949,N_16065);
or U16806 (N_16806,N_15849,N_16138);
and U16807 (N_16807,N_15651,N_16096);
or U16808 (N_16808,N_15720,N_15854);
nand U16809 (N_16809,N_16089,N_16117);
xnor U16810 (N_16810,N_15870,N_15983);
and U16811 (N_16811,N_16105,N_16149);
or U16812 (N_16812,N_16170,N_15786);
xnor U16813 (N_16813,N_15652,N_15667);
nand U16814 (N_16814,N_15904,N_15678);
nand U16815 (N_16815,N_15885,N_16108);
or U16816 (N_16816,N_16083,N_16032);
nor U16817 (N_16817,N_15812,N_16010);
nand U16818 (N_16818,N_15641,N_15826);
or U16819 (N_16819,N_16208,N_15686);
xor U16820 (N_16820,N_16081,N_15843);
or U16821 (N_16821,N_16046,N_15741);
or U16822 (N_16822,N_15828,N_16184);
nor U16823 (N_16823,N_16209,N_15965);
or U16824 (N_16824,N_16021,N_16095);
and U16825 (N_16825,N_15895,N_15730);
and U16826 (N_16826,N_15903,N_16174);
nor U16827 (N_16827,N_15791,N_15820);
nand U16828 (N_16828,N_15994,N_15715);
xnor U16829 (N_16829,N_15780,N_15845);
xor U16830 (N_16830,N_16241,N_15878);
or U16831 (N_16831,N_16087,N_15826);
or U16832 (N_16832,N_16092,N_16081);
or U16833 (N_16833,N_16167,N_16236);
xor U16834 (N_16834,N_15748,N_15675);
and U16835 (N_16835,N_15635,N_15734);
nand U16836 (N_16836,N_15777,N_16167);
or U16837 (N_16837,N_15940,N_15991);
and U16838 (N_16838,N_15712,N_15675);
nand U16839 (N_16839,N_16135,N_16057);
or U16840 (N_16840,N_16026,N_16173);
and U16841 (N_16841,N_16151,N_15901);
or U16842 (N_16842,N_15680,N_16135);
xnor U16843 (N_16843,N_15670,N_15640);
and U16844 (N_16844,N_15679,N_15697);
nor U16845 (N_16845,N_15763,N_16188);
nor U16846 (N_16846,N_15667,N_16055);
or U16847 (N_16847,N_16085,N_16215);
nand U16848 (N_16848,N_15637,N_15858);
nand U16849 (N_16849,N_15694,N_15708);
and U16850 (N_16850,N_15648,N_15674);
or U16851 (N_16851,N_16247,N_15908);
or U16852 (N_16852,N_15808,N_16142);
nand U16853 (N_16853,N_16096,N_15970);
xnor U16854 (N_16854,N_15881,N_15762);
nand U16855 (N_16855,N_16074,N_15856);
or U16856 (N_16856,N_15985,N_15780);
xor U16857 (N_16857,N_16062,N_15877);
or U16858 (N_16858,N_15745,N_15814);
nand U16859 (N_16859,N_15786,N_16159);
nor U16860 (N_16860,N_15626,N_15882);
and U16861 (N_16861,N_15995,N_16191);
and U16862 (N_16862,N_15889,N_15835);
or U16863 (N_16863,N_16213,N_16208);
and U16864 (N_16864,N_16046,N_15762);
nor U16865 (N_16865,N_15828,N_16244);
nand U16866 (N_16866,N_16111,N_15939);
or U16867 (N_16867,N_16021,N_16066);
nor U16868 (N_16868,N_15783,N_15683);
or U16869 (N_16869,N_16058,N_15674);
nand U16870 (N_16870,N_16048,N_16100);
xnor U16871 (N_16871,N_15676,N_16184);
xnor U16872 (N_16872,N_16151,N_16138);
and U16873 (N_16873,N_15766,N_16173);
and U16874 (N_16874,N_15933,N_16061);
or U16875 (N_16875,N_16873,N_16575);
and U16876 (N_16876,N_16831,N_16471);
xnor U16877 (N_16877,N_16441,N_16447);
nor U16878 (N_16878,N_16334,N_16439);
and U16879 (N_16879,N_16299,N_16607);
nor U16880 (N_16880,N_16353,N_16642);
and U16881 (N_16881,N_16786,N_16468);
and U16882 (N_16882,N_16292,N_16511);
or U16883 (N_16883,N_16584,N_16836);
nor U16884 (N_16884,N_16290,N_16323);
and U16885 (N_16885,N_16291,N_16378);
xor U16886 (N_16886,N_16658,N_16677);
or U16887 (N_16887,N_16636,N_16619);
or U16888 (N_16888,N_16683,N_16525);
xnor U16889 (N_16889,N_16773,N_16874);
nand U16890 (N_16890,N_16557,N_16304);
and U16891 (N_16891,N_16380,N_16802);
nor U16892 (N_16892,N_16665,N_16676);
xor U16893 (N_16893,N_16377,N_16365);
or U16894 (N_16894,N_16777,N_16261);
or U16895 (N_16895,N_16765,N_16253);
or U16896 (N_16896,N_16706,N_16598);
and U16897 (N_16897,N_16685,N_16474);
or U16898 (N_16898,N_16274,N_16537);
and U16899 (N_16899,N_16805,N_16398);
nand U16900 (N_16900,N_16281,N_16479);
or U16901 (N_16901,N_16345,N_16858);
nor U16902 (N_16902,N_16548,N_16846);
and U16903 (N_16903,N_16824,N_16724);
nand U16904 (N_16904,N_16670,N_16250);
nand U16905 (N_16905,N_16652,N_16576);
nand U16906 (N_16906,N_16404,N_16754);
and U16907 (N_16907,N_16579,N_16632);
xnor U16908 (N_16908,N_16317,N_16593);
or U16909 (N_16909,N_16708,N_16432);
or U16910 (N_16910,N_16461,N_16637);
and U16911 (N_16911,N_16798,N_16507);
nand U16912 (N_16912,N_16610,N_16395);
or U16913 (N_16913,N_16739,N_16302);
nor U16914 (N_16914,N_16324,N_16341);
nand U16915 (N_16915,N_16280,N_16311);
nor U16916 (N_16916,N_16418,N_16329);
xor U16917 (N_16917,N_16847,N_16767);
xor U16918 (N_16918,N_16499,N_16622);
xnor U16919 (N_16919,N_16809,N_16297);
and U16920 (N_16920,N_16743,N_16258);
nand U16921 (N_16921,N_16456,N_16806);
nand U16922 (N_16922,N_16675,N_16366);
or U16923 (N_16923,N_16449,N_16348);
xor U16924 (N_16924,N_16803,N_16408);
nor U16925 (N_16925,N_16394,N_16497);
xor U16926 (N_16926,N_16626,N_16662);
or U16927 (N_16927,N_16428,N_16691);
nand U16928 (N_16928,N_16382,N_16533);
xor U16929 (N_16929,N_16480,N_16780);
nand U16930 (N_16930,N_16571,N_16519);
and U16931 (N_16931,N_16860,N_16407);
nor U16932 (N_16932,N_16271,N_16655);
and U16933 (N_16933,N_16262,N_16793);
xor U16934 (N_16934,N_16726,N_16856);
xor U16935 (N_16935,N_16732,N_16494);
xor U16936 (N_16936,N_16750,N_16761);
xnor U16937 (N_16937,N_16355,N_16707);
nand U16938 (N_16938,N_16633,N_16473);
or U16939 (N_16939,N_16838,N_16276);
xnor U16940 (N_16940,N_16427,N_16293);
or U16941 (N_16941,N_16429,N_16544);
xor U16942 (N_16942,N_16866,N_16784);
nand U16943 (N_16943,N_16360,N_16747);
nor U16944 (N_16944,N_16603,N_16712);
and U16945 (N_16945,N_16681,N_16412);
and U16946 (N_16946,N_16554,N_16451);
nand U16947 (N_16947,N_16472,N_16864);
or U16948 (N_16948,N_16374,N_16556);
or U16949 (N_16949,N_16401,N_16616);
nor U16950 (N_16950,N_16434,N_16645);
xor U16951 (N_16951,N_16347,N_16498);
and U16952 (N_16952,N_16352,N_16789);
xor U16953 (N_16953,N_16346,N_16267);
or U16954 (N_16954,N_16564,N_16390);
and U16955 (N_16955,N_16755,N_16410);
and U16956 (N_16956,N_16463,N_16791);
or U16957 (N_16957,N_16693,N_16697);
nor U16958 (N_16958,N_16667,N_16825);
xor U16959 (N_16959,N_16844,N_16771);
nand U16960 (N_16960,N_16335,N_16698);
nand U16961 (N_16961,N_16344,N_16857);
xor U16962 (N_16962,N_16621,N_16251);
or U16963 (N_16963,N_16617,N_16478);
and U16964 (N_16964,N_16597,N_16464);
and U16965 (N_16965,N_16490,N_16289);
xnor U16966 (N_16966,N_16336,N_16592);
nand U16967 (N_16967,N_16295,N_16254);
xnor U16968 (N_16968,N_16406,N_16466);
xor U16969 (N_16969,N_16322,N_16285);
nand U16970 (N_16970,N_16435,N_16531);
nor U16971 (N_16971,N_16550,N_16298);
xor U16972 (N_16972,N_16587,N_16259);
and U16973 (N_16973,N_16651,N_16327);
or U16974 (N_16974,N_16692,N_16385);
or U16975 (N_16975,N_16294,N_16438);
nand U16976 (N_16976,N_16872,N_16588);
xor U16977 (N_16977,N_16837,N_16530);
nand U16978 (N_16978,N_16419,N_16284);
nand U16979 (N_16979,N_16397,N_16462);
nand U16980 (N_16980,N_16255,N_16672);
nor U16981 (N_16981,N_16359,N_16339);
and U16982 (N_16982,N_16300,N_16371);
xor U16983 (N_16983,N_16850,N_16534);
nand U16984 (N_16984,N_16721,N_16423);
or U16985 (N_16985,N_16639,N_16442);
nor U16986 (N_16986,N_16606,N_16361);
and U16987 (N_16987,N_16528,N_16331);
or U16988 (N_16988,N_16287,N_16605);
nor U16989 (N_16989,N_16833,N_16391);
xor U16990 (N_16990,N_16379,N_16723);
nor U16991 (N_16991,N_16759,N_16745);
nor U16992 (N_16992,N_16868,N_16792);
nand U16993 (N_16993,N_16728,N_16363);
nor U16994 (N_16994,N_16565,N_16520);
and U16995 (N_16995,N_16711,N_16653);
and U16996 (N_16996,N_16426,N_16646);
or U16997 (N_16997,N_16535,N_16826);
nand U16998 (N_16998,N_16774,N_16573);
nand U16999 (N_16999,N_16853,N_16599);
nand U17000 (N_17000,N_16720,N_16492);
xor U17001 (N_17001,N_16443,N_16278);
xnor U17002 (N_17002,N_16370,N_16594);
or U17003 (N_17003,N_16785,N_16614);
or U17004 (N_17004,N_16562,N_16421);
nor U17005 (N_17005,N_16811,N_16738);
nor U17006 (N_17006,N_16638,N_16779);
and U17007 (N_17007,N_16744,N_16608);
and U17008 (N_17008,N_16263,N_16736);
nand U17009 (N_17009,N_16612,N_16558);
nor U17010 (N_17010,N_16387,N_16756);
nor U17011 (N_17011,N_16431,N_16867);
nand U17012 (N_17012,N_16735,N_16265);
or U17013 (N_17013,N_16787,N_16264);
nand U17014 (N_17014,N_16402,N_16269);
or U17015 (N_17015,N_16839,N_16581);
xnor U17016 (N_17016,N_16318,N_16815);
nor U17017 (N_17017,N_16440,N_16372);
nor U17018 (N_17018,N_16524,N_16635);
xor U17019 (N_17019,N_16338,N_16748);
nand U17020 (N_17020,N_16800,N_16521);
nor U17021 (N_17021,N_16852,N_16515);
nor U17022 (N_17022,N_16770,N_16717);
nand U17023 (N_17023,N_16673,N_16527);
or U17024 (N_17024,N_16325,N_16600);
and U17025 (N_17025,N_16489,N_16319);
or U17026 (N_17026,N_16381,N_16545);
xor U17027 (N_17027,N_16386,N_16816);
and U17028 (N_17028,N_16714,N_16812);
or U17029 (N_17029,N_16580,N_16817);
nor U17030 (N_17030,N_16790,N_16769);
nor U17031 (N_17031,N_16666,N_16749);
or U17032 (N_17032,N_16611,N_16475);
and U17033 (N_17033,N_16567,N_16768);
and U17034 (N_17034,N_16668,N_16843);
or U17035 (N_17035,N_16574,N_16517);
nand U17036 (N_17036,N_16848,N_16446);
nor U17037 (N_17037,N_16482,N_16448);
nor U17038 (N_17038,N_16303,N_16296);
nand U17039 (N_17039,N_16582,N_16585);
nor U17040 (N_17040,N_16686,N_16312);
or U17041 (N_17041,N_16591,N_16861);
and U17042 (N_17042,N_16827,N_16467);
or U17043 (N_17043,N_16804,N_16518);
xnor U17044 (N_17044,N_16357,N_16742);
nand U17045 (N_17045,N_16551,N_16595);
nand U17046 (N_17046,N_16716,N_16604);
nor U17047 (N_17047,N_16602,N_16737);
and U17048 (N_17048,N_16457,N_16454);
and U17049 (N_17049,N_16763,N_16384);
and U17050 (N_17050,N_16659,N_16413);
nor U17051 (N_17051,N_16859,N_16409);
or U17052 (N_17052,N_16752,N_16851);
nor U17053 (N_17053,N_16627,N_16741);
or U17054 (N_17054,N_16425,N_16829);
nor U17055 (N_17055,N_16620,N_16758);
or U17056 (N_17056,N_16730,N_16561);
and U17057 (N_17057,N_16333,N_16649);
nor U17058 (N_17058,N_16354,N_16506);
or U17059 (N_17059,N_16688,N_16753);
and U17060 (N_17060,N_16689,N_16559);
nor U17061 (N_17061,N_16678,N_16500);
and U17062 (N_17062,N_16465,N_16332);
nor U17063 (N_17063,N_16514,N_16705);
xnor U17064 (N_17064,N_16775,N_16664);
or U17065 (N_17065,N_16648,N_16808);
xor U17066 (N_17066,N_16650,N_16256);
and U17067 (N_17067,N_16855,N_16504);
nand U17068 (N_17068,N_16729,N_16420);
and U17069 (N_17069,N_16814,N_16657);
and U17070 (N_17070,N_16863,N_16268);
or U17071 (N_17071,N_16283,N_16687);
and U17072 (N_17072,N_16546,N_16563);
nand U17073 (N_17073,N_16695,N_16656);
and U17074 (N_17074,N_16794,N_16453);
xnor U17075 (N_17075,N_16640,N_16356);
nand U17076 (N_17076,N_16388,N_16376);
or U17077 (N_17077,N_16772,N_16424);
nand U17078 (N_17078,N_16654,N_16330);
xor U17079 (N_17079,N_16845,N_16694);
and U17080 (N_17080,N_16358,N_16870);
nor U17081 (N_17081,N_16310,N_16275);
nor U17082 (N_17082,N_16552,N_16458);
and U17083 (N_17083,N_16415,N_16841);
and U17084 (N_17084,N_16306,N_16822);
xor U17085 (N_17085,N_16375,N_16628);
nor U17086 (N_17086,N_16586,N_16510);
nor U17087 (N_17087,N_16549,N_16350);
and U17088 (N_17088,N_16286,N_16630);
nor U17089 (N_17089,N_16734,N_16799);
nor U17090 (N_17090,N_16618,N_16495);
nand U17091 (N_17091,N_16340,N_16301);
and U17092 (N_17092,N_16647,N_16342);
nand U17093 (N_17093,N_16279,N_16543);
nand U17094 (N_17094,N_16444,N_16437);
or U17095 (N_17095,N_16733,N_16682);
xor U17096 (N_17096,N_16710,N_16541);
xor U17097 (N_17097,N_16288,N_16487);
or U17098 (N_17098,N_16625,N_16555);
xor U17099 (N_17099,N_16349,N_16272);
xnor U17100 (N_17100,N_16417,N_16400);
xnor U17101 (N_17101,N_16623,N_16849);
xnor U17102 (N_17102,N_16674,N_16485);
nand U17103 (N_17103,N_16644,N_16782);
and U17104 (N_17104,N_16493,N_16613);
nor U17105 (N_17105,N_16315,N_16491);
nand U17106 (N_17106,N_16871,N_16522);
and U17107 (N_17107,N_16718,N_16422);
and U17108 (N_17108,N_16513,N_16641);
and U17109 (N_17109,N_16307,N_16788);
nor U17110 (N_17110,N_16796,N_16389);
and U17111 (N_17111,N_16508,N_16835);
xnor U17112 (N_17112,N_16807,N_16722);
xor U17113 (N_17113,N_16516,N_16416);
nor U17114 (N_17114,N_16542,N_16309);
nor U17115 (N_17115,N_16455,N_16411);
xor U17116 (N_17116,N_16813,N_16572);
or U17117 (N_17117,N_16368,N_16660);
and U17118 (N_17118,N_16501,N_16696);
and U17119 (N_17119,N_16452,N_16529);
or U17120 (N_17120,N_16713,N_16364);
nand U17121 (N_17121,N_16430,N_16578);
nor U17122 (N_17122,N_16631,N_16776);
or U17123 (N_17123,N_16690,N_16823);
xnor U17124 (N_17124,N_16308,N_16526);
or U17125 (N_17125,N_16820,N_16781);
or U17126 (N_17126,N_16362,N_16762);
nor U17127 (N_17127,N_16797,N_16684);
or U17128 (N_17128,N_16252,N_16760);
nor U17129 (N_17129,N_16680,N_16320);
or U17130 (N_17130,N_16373,N_16570);
nand U17131 (N_17131,N_16701,N_16405);
nor U17132 (N_17132,N_16764,N_16343);
xnor U17133 (N_17133,N_16488,N_16709);
xor U17134 (N_17134,N_16821,N_16832);
or U17135 (N_17135,N_16643,N_16509);
nand U17136 (N_17136,N_16547,N_16316);
nor U17137 (N_17137,N_16477,N_16450);
xnor U17138 (N_17138,N_16273,N_16679);
xnor U17139 (N_17139,N_16393,N_16321);
or U17140 (N_17140,N_16369,N_16609);
or U17141 (N_17141,N_16536,N_16566);
nor U17142 (N_17142,N_16476,N_16260);
nand U17143 (N_17143,N_16663,N_16337);
xor U17144 (N_17144,N_16740,N_16532);
nand U17145 (N_17145,N_16433,N_16396);
or U17146 (N_17146,N_16795,N_16810);
and U17147 (N_17147,N_16801,N_16589);
xnor U17148 (N_17148,N_16703,N_16481);
nand U17149 (N_17149,N_16624,N_16560);
nor U17150 (N_17150,N_16569,N_16746);
and U17151 (N_17151,N_16751,N_16469);
or U17152 (N_17152,N_16470,N_16270);
nand U17153 (N_17153,N_16725,N_16326);
or U17154 (N_17154,N_16601,N_16818);
or U17155 (N_17155,N_16834,N_16577);
nand U17156 (N_17156,N_16266,N_16778);
xor U17157 (N_17157,N_16828,N_16634);
or U17158 (N_17158,N_16328,N_16671);
and U17159 (N_17159,N_16783,N_16483);
or U17160 (N_17160,N_16819,N_16757);
nor U17161 (N_17161,N_16539,N_16719);
nand U17162 (N_17162,N_16661,N_16862);
xor U17163 (N_17163,N_16854,N_16445);
or U17164 (N_17164,N_16596,N_16367);
and U17165 (N_17165,N_16282,N_16484);
nand U17166 (N_17166,N_16731,N_16700);
xor U17167 (N_17167,N_16496,N_16590);
xor U17168 (N_17168,N_16314,N_16540);
nor U17169 (N_17169,N_16583,N_16383);
and U17170 (N_17170,N_16277,N_16715);
xor U17171 (N_17171,N_16842,N_16436);
nor U17172 (N_17172,N_16392,N_16869);
nand U17173 (N_17173,N_16257,N_16615);
and U17174 (N_17174,N_16313,N_16727);
nand U17175 (N_17175,N_16704,N_16865);
nand U17176 (N_17176,N_16512,N_16460);
nor U17177 (N_17177,N_16414,N_16699);
nor U17178 (N_17178,N_16399,N_16305);
and U17179 (N_17179,N_16766,N_16502);
nand U17180 (N_17180,N_16486,N_16568);
xnor U17181 (N_17181,N_16840,N_16403);
nor U17182 (N_17182,N_16351,N_16503);
or U17183 (N_17183,N_16538,N_16505);
or U17184 (N_17184,N_16629,N_16669);
xor U17185 (N_17185,N_16553,N_16702);
and U17186 (N_17186,N_16459,N_16830);
nor U17187 (N_17187,N_16523,N_16504);
nand U17188 (N_17188,N_16261,N_16272);
xor U17189 (N_17189,N_16417,N_16450);
xor U17190 (N_17190,N_16582,N_16618);
nor U17191 (N_17191,N_16563,N_16278);
and U17192 (N_17192,N_16442,N_16428);
and U17193 (N_17193,N_16843,N_16296);
nand U17194 (N_17194,N_16330,N_16359);
xnor U17195 (N_17195,N_16376,N_16841);
or U17196 (N_17196,N_16366,N_16867);
nor U17197 (N_17197,N_16298,N_16611);
nor U17198 (N_17198,N_16821,N_16275);
xor U17199 (N_17199,N_16347,N_16424);
or U17200 (N_17200,N_16510,N_16661);
and U17201 (N_17201,N_16682,N_16418);
xnor U17202 (N_17202,N_16601,N_16586);
xnor U17203 (N_17203,N_16827,N_16452);
or U17204 (N_17204,N_16581,N_16448);
xor U17205 (N_17205,N_16265,N_16675);
nand U17206 (N_17206,N_16669,N_16642);
nor U17207 (N_17207,N_16824,N_16638);
nand U17208 (N_17208,N_16591,N_16669);
xor U17209 (N_17209,N_16520,N_16439);
and U17210 (N_17210,N_16722,N_16543);
nand U17211 (N_17211,N_16850,N_16844);
nor U17212 (N_17212,N_16811,N_16671);
nand U17213 (N_17213,N_16559,N_16775);
nand U17214 (N_17214,N_16372,N_16374);
nor U17215 (N_17215,N_16643,N_16566);
nor U17216 (N_17216,N_16366,N_16385);
or U17217 (N_17217,N_16763,N_16812);
nand U17218 (N_17218,N_16610,N_16553);
nand U17219 (N_17219,N_16771,N_16316);
nand U17220 (N_17220,N_16602,N_16756);
or U17221 (N_17221,N_16528,N_16447);
and U17222 (N_17222,N_16780,N_16680);
nand U17223 (N_17223,N_16425,N_16428);
xnor U17224 (N_17224,N_16572,N_16652);
nand U17225 (N_17225,N_16294,N_16606);
nor U17226 (N_17226,N_16293,N_16579);
and U17227 (N_17227,N_16579,N_16482);
and U17228 (N_17228,N_16656,N_16852);
xor U17229 (N_17229,N_16786,N_16371);
or U17230 (N_17230,N_16630,N_16842);
and U17231 (N_17231,N_16718,N_16418);
and U17232 (N_17232,N_16653,N_16608);
and U17233 (N_17233,N_16663,N_16855);
nand U17234 (N_17234,N_16806,N_16515);
nor U17235 (N_17235,N_16823,N_16857);
xnor U17236 (N_17236,N_16797,N_16867);
or U17237 (N_17237,N_16768,N_16314);
xnor U17238 (N_17238,N_16784,N_16562);
xnor U17239 (N_17239,N_16578,N_16674);
and U17240 (N_17240,N_16627,N_16467);
and U17241 (N_17241,N_16612,N_16520);
nor U17242 (N_17242,N_16609,N_16536);
xor U17243 (N_17243,N_16567,N_16653);
xor U17244 (N_17244,N_16571,N_16266);
or U17245 (N_17245,N_16294,N_16445);
xnor U17246 (N_17246,N_16810,N_16302);
nor U17247 (N_17247,N_16759,N_16675);
and U17248 (N_17248,N_16803,N_16812);
and U17249 (N_17249,N_16677,N_16583);
nand U17250 (N_17250,N_16615,N_16688);
and U17251 (N_17251,N_16318,N_16763);
or U17252 (N_17252,N_16758,N_16851);
nor U17253 (N_17253,N_16453,N_16437);
nor U17254 (N_17254,N_16295,N_16410);
nor U17255 (N_17255,N_16659,N_16767);
and U17256 (N_17256,N_16621,N_16391);
or U17257 (N_17257,N_16517,N_16582);
or U17258 (N_17258,N_16806,N_16470);
and U17259 (N_17259,N_16866,N_16654);
xnor U17260 (N_17260,N_16314,N_16508);
or U17261 (N_17261,N_16456,N_16561);
or U17262 (N_17262,N_16570,N_16567);
xnor U17263 (N_17263,N_16375,N_16873);
xor U17264 (N_17264,N_16629,N_16446);
nor U17265 (N_17265,N_16298,N_16333);
nor U17266 (N_17266,N_16787,N_16495);
or U17267 (N_17267,N_16547,N_16527);
nand U17268 (N_17268,N_16851,N_16674);
xnor U17269 (N_17269,N_16831,N_16353);
or U17270 (N_17270,N_16650,N_16750);
xnor U17271 (N_17271,N_16288,N_16419);
nor U17272 (N_17272,N_16586,N_16298);
nor U17273 (N_17273,N_16705,N_16261);
and U17274 (N_17274,N_16360,N_16479);
and U17275 (N_17275,N_16721,N_16419);
xnor U17276 (N_17276,N_16678,N_16727);
nor U17277 (N_17277,N_16402,N_16845);
or U17278 (N_17278,N_16799,N_16352);
xnor U17279 (N_17279,N_16520,N_16257);
and U17280 (N_17280,N_16803,N_16662);
xnor U17281 (N_17281,N_16410,N_16412);
or U17282 (N_17282,N_16639,N_16419);
nor U17283 (N_17283,N_16554,N_16853);
and U17284 (N_17284,N_16600,N_16558);
nand U17285 (N_17285,N_16848,N_16498);
or U17286 (N_17286,N_16682,N_16689);
xor U17287 (N_17287,N_16791,N_16347);
nand U17288 (N_17288,N_16493,N_16772);
nand U17289 (N_17289,N_16691,N_16457);
nand U17290 (N_17290,N_16321,N_16534);
nor U17291 (N_17291,N_16524,N_16645);
and U17292 (N_17292,N_16802,N_16453);
or U17293 (N_17293,N_16467,N_16837);
xnor U17294 (N_17294,N_16518,N_16568);
nand U17295 (N_17295,N_16715,N_16760);
and U17296 (N_17296,N_16580,N_16359);
xor U17297 (N_17297,N_16784,N_16554);
and U17298 (N_17298,N_16677,N_16471);
or U17299 (N_17299,N_16286,N_16695);
or U17300 (N_17300,N_16792,N_16766);
or U17301 (N_17301,N_16485,N_16330);
nand U17302 (N_17302,N_16503,N_16417);
and U17303 (N_17303,N_16540,N_16357);
and U17304 (N_17304,N_16759,N_16848);
and U17305 (N_17305,N_16718,N_16397);
nor U17306 (N_17306,N_16533,N_16601);
or U17307 (N_17307,N_16628,N_16382);
or U17308 (N_17308,N_16446,N_16424);
xor U17309 (N_17309,N_16255,N_16687);
nor U17310 (N_17310,N_16779,N_16750);
xnor U17311 (N_17311,N_16703,N_16544);
nand U17312 (N_17312,N_16367,N_16322);
or U17313 (N_17313,N_16706,N_16731);
nand U17314 (N_17314,N_16828,N_16504);
nand U17315 (N_17315,N_16438,N_16545);
and U17316 (N_17316,N_16334,N_16413);
nand U17317 (N_17317,N_16507,N_16597);
nor U17318 (N_17318,N_16489,N_16583);
nand U17319 (N_17319,N_16555,N_16492);
xor U17320 (N_17320,N_16665,N_16343);
xnor U17321 (N_17321,N_16514,N_16578);
nand U17322 (N_17322,N_16431,N_16534);
nand U17323 (N_17323,N_16713,N_16645);
xor U17324 (N_17324,N_16643,N_16456);
nand U17325 (N_17325,N_16656,N_16427);
xor U17326 (N_17326,N_16874,N_16619);
nand U17327 (N_17327,N_16754,N_16846);
or U17328 (N_17328,N_16480,N_16328);
nand U17329 (N_17329,N_16560,N_16563);
nand U17330 (N_17330,N_16700,N_16417);
nand U17331 (N_17331,N_16278,N_16489);
and U17332 (N_17332,N_16799,N_16836);
or U17333 (N_17333,N_16454,N_16279);
nand U17334 (N_17334,N_16304,N_16458);
nand U17335 (N_17335,N_16579,N_16652);
nand U17336 (N_17336,N_16605,N_16277);
or U17337 (N_17337,N_16602,N_16377);
or U17338 (N_17338,N_16379,N_16430);
or U17339 (N_17339,N_16771,N_16608);
or U17340 (N_17340,N_16544,N_16345);
and U17341 (N_17341,N_16569,N_16471);
and U17342 (N_17342,N_16374,N_16756);
and U17343 (N_17343,N_16518,N_16695);
xnor U17344 (N_17344,N_16296,N_16385);
nor U17345 (N_17345,N_16438,N_16744);
nand U17346 (N_17346,N_16822,N_16655);
nand U17347 (N_17347,N_16466,N_16252);
or U17348 (N_17348,N_16363,N_16836);
xor U17349 (N_17349,N_16657,N_16815);
xnor U17350 (N_17350,N_16679,N_16393);
or U17351 (N_17351,N_16492,N_16787);
or U17352 (N_17352,N_16389,N_16285);
xor U17353 (N_17353,N_16404,N_16689);
nor U17354 (N_17354,N_16284,N_16739);
or U17355 (N_17355,N_16429,N_16499);
xnor U17356 (N_17356,N_16480,N_16397);
or U17357 (N_17357,N_16360,N_16539);
or U17358 (N_17358,N_16777,N_16613);
and U17359 (N_17359,N_16578,N_16571);
or U17360 (N_17360,N_16748,N_16402);
nor U17361 (N_17361,N_16346,N_16790);
nand U17362 (N_17362,N_16354,N_16687);
or U17363 (N_17363,N_16522,N_16872);
nand U17364 (N_17364,N_16512,N_16414);
and U17365 (N_17365,N_16362,N_16257);
nor U17366 (N_17366,N_16666,N_16815);
or U17367 (N_17367,N_16769,N_16399);
and U17368 (N_17368,N_16267,N_16460);
nor U17369 (N_17369,N_16298,N_16794);
and U17370 (N_17370,N_16829,N_16691);
nor U17371 (N_17371,N_16411,N_16668);
xnor U17372 (N_17372,N_16855,N_16868);
nand U17373 (N_17373,N_16342,N_16437);
and U17374 (N_17374,N_16828,N_16493);
and U17375 (N_17375,N_16271,N_16429);
nor U17376 (N_17376,N_16627,N_16515);
or U17377 (N_17377,N_16844,N_16359);
nor U17378 (N_17378,N_16670,N_16428);
or U17379 (N_17379,N_16522,N_16678);
or U17380 (N_17380,N_16304,N_16589);
xnor U17381 (N_17381,N_16525,N_16756);
xnor U17382 (N_17382,N_16260,N_16533);
nor U17383 (N_17383,N_16667,N_16551);
nor U17384 (N_17384,N_16779,N_16587);
and U17385 (N_17385,N_16774,N_16554);
nand U17386 (N_17386,N_16402,N_16420);
or U17387 (N_17387,N_16353,N_16666);
xor U17388 (N_17388,N_16496,N_16664);
or U17389 (N_17389,N_16851,N_16565);
and U17390 (N_17390,N_16728,N_16488);
nor U17391 (N_17391,N_16396,N_16825);
nor U17392 (N_17392,N_16558,N_16502);
nor U17393 (N_17393,N_16508,N_16316);
or U17394 (N_17394,N_16821,N_16765);
nand U17395 (N_17395,N_16403,N_16606);
nand U17396 (N_17396,N_16484,N_16812);
nor U17397 (N_17397,N_16312,N_16306);
or U17398 (N_17398,N_16578,N_16368);
nor U17399 (N_17399,N_16688,N_16405);
or U17400 (N_17400,N_16278,N_16326);
nand U17401 (N_17401,N_16558,N_16287);
xor U17402 (N_17402,N_16369,N_16810);
nand U17403 (N_17403,N_16340,N_16325);
xor U17404 (N_17404,N_16368,N_16540);
or U17405 (N_17405,N_16650,N_16266);
xor U17406 (N_17406,N_16620,N_16606);
xnor U17407 (N_17407,N_16489,N_16810);
xnor U17408 (N_17408,N_16484,N_16768);
nor U17409 (N_17409,N_16366,N_16739);
xor U17410 (N_17410,N_16750,N_16489);
xor U17411 (N_17411,N_16576,N_16452);
or U17412 (N_17412,N_16265,N_16493);
nor U17413 (N_17413,N_16505,N_16265);
or U17414 (N_17414,N_16849,N_16669);
nand U17415 (N_17415,N_16835,N_16473);
nand U17416 (N_17416,N_16257,N_16306);
or U17417 (N_17417,N_16414,N_16261);
nand U17418 (N_17418,N_16777,N_16516);
or U17419 (N_17419,N_16822,N_16253);
nor U17420 (N_17420,N_16463,N_16339);
xnor U17421 (N_17421,N_16622,N_16740);
xor U17422 (N_17422,N_16564,N_16813);
and U17423 (N_17423,N_16475,N_16497);
and U17424 (N_17424,N_16650,N_16580);
nor U17425 (N_17425,N_16470,N_16291);
xor U17426 (N_17426,N_16295,N_16623);
and U17427 (N_17427,N_16591,N_16619);
nor U17428 (N_17428,N_16652,N_16669);
nor U17429 (N_17429,N_16410,N_16262);
xor U17430 (N_17430,N_16746,N_16315);
nor U17431 (N_17431,N_16765,N_16489);
nand U17432 (N_17432,N_16317,N_16769);
and U17433 (N_17433,N_16301,N_16819);
nand U17434 (N_17434,N_16315,N_16268);
nand U17435 (N_17435,N_16511,N_16393);
or U17436 (N_17436,N_16747,N_16536);
and U17437 (N_17437,N_16872,N_16342);
nor U17438 (N_17438,N_16512,N_16549);
nand U17439 (N_17439,N_16767,N_16608);
xor U17440 (N_17440,N_16645,N_16512);
or U17441 (N_17441,N_16560,N_16857);
nand U17442 (N_17442,N_16461,N_16381);
nor U17443 (N_17443,N_16534,N_16794);
or U17444 (N_17444,N_16378,N_16580);
nand U17445 (N_17445,N_16613,N_16840);
xnor U17446 (N_17446,N_16780,N_16354);
xnor U17447 (N_17447,N_16584,N_16598);
or U17448 (N_17448,N_16438,N_16665);
nor U17449 (N_17449,N_16264,N_16556);
nand U17450 (N_17450,N_16382,N_16732);
nand U17451 (N_17451,N_16769,N_16668);
xnor U17452 (N_17452,N_16467,N_16826);
and U17453 (N_17453,N_16316,N_16697);
xnor U17454 (N_17454,N_16273,N_16659);
nand U17455 (N_17455,N_16451,N_16659);
nand U17456 (N_17456,N_16605,N_16656);
xor U17457 (N_17457,N_16532,N_16555);
xor U17458 (N_17458,N_16566,N_16327);
nor U17459 (N_17459,N_16356,N_16564);
nand U17460 (N_17460,N_16655,N_16411);
xnor U17461 (N_17461,N_16422,N_16814);
and U17462 (N_17462,N_16737,N_16698);
nor U17463 (N_17463,N_16684,N_16497);
xnor U17464 (N_17464,N_16360,N_16536);
nand U17465 (N_17465,N_16385,N_16684);
and U17466 (N_17466,N_16694,N_16346);
nand U17467 (N_17467,N_16534,N_16319);
nand U17468 (N_17468,N_16690,N_16551);
nor U17469 (N_17469,N_16819,N_16476);
or U17470 (N_17470,N_16557,N_16861);
xnor U17471 (N_17471,N_16798,N_16824);
xor U17472 (N_17472,N_16731,N_16604);
nand U17473 (N_17473,N_16591,N_16823);
nand U17474 (N_17474,N_16404,N_16512);
xor U17475 (N_17475,N_16732,N_16260);
xnor U17476 (N_17476,N_16455,N_16553);
and U17477 (N_17477,N_16680,N_16768);
nand U17478 (N_17478,N_16523,N_16501);
or U17479 (N_17479,N_16671,N_16685);
or U17480 (N_17480,N_16599,N_16739);
or U17481 (N_17481,N_16738,N_16418);
nor U17482 (N_17482,N_16705,N_16831);
xnor U17483 (N_17483,N_16341,N_16588);
and U17484 (N_17484,N_16712,N_16780);
or U17485 (N_17485,N_16604,N_16538);
nor U17486 (N_17486,N_16763,N_16696);
nor U17487 (N_17487,N_16719,N_16414);
nand U17488 (N_17488,N_16484,N_16413);
nand U17489 (N_17489,N_16864,N_16439);
nand U17490 (N_17490,N_16458,N_16447);
nor U17491 (N_17491,N_16325,N_16491);
or U17492 (N_17492,N_16398,N_16724);
or U17493 (N_17493,N_16598,N_16459);
nor U17494 (N_17494,N_16785,N_16681);
or U17495 (N_17495,N_16476,N_16568);
and U17496 (N_17496,N_16475,N_16253);
nor U17497 (N_17497,N_16709,N_16378);
and U17498 (N_17498,N_16326,N_16268);
and U17499 (N_17499,N_16423,N_16837);
and U17500 (N_17500,N_17320,N_17488);
and U17501 (N_17501,N_17353,N_16988);
and U17502 (N_17502,N_17202,N_17229);
or U17503 (N_17503,N_17096,N_17107);
nand U17504 (N_17504,N_17355,N_17310);
and U17505 (N_17505,N_16875,N_17257);
xnor U17506 (N_17506,N_17497,N_17483);
and U17507 (N_17507,N_17236,N_17116);
nor U17508 (N_17508,N_16883,N_16998);
and U17509 (N_17509,N_17030,N_17144);
nand U17510 (N_17510,N_16910,N_17270);
nand U17511 (N_17511,N_17370,N_17165);
nor U17512 (N_17512,N_17239,N_17232);
or U17513 (N_17513,N_17474,N_17324);
nand U17514 (N_17514,N_17237,N_17117);
or U17515 (N_17515,N_17036,N_17003);
and U17516 (N_17516,N_17216,N_16878);
and U17517 (N_17517,N_17098,N_17214);
nor U17518 (N_17518,N_16944,N_17449);
nor U17519 (N_17519,N_16924,N_17146);
nand U17520 (N_17520,N_17022,N_17460);
nor U17521 (N_17521,N_16876,N_17073);
and U17522 (N_17522,N_17447,N_16982);
xnor U17523 (N_17523,N_16949,N_17392);
and U17524 (N_17524,N_17225,N_17046);
or U17525 (N_17525,N_17391,N_17372);
nor U17526 (N_17526,N_17135,N_17095);
and U17527 (N_17527,N_17057,N_17174);
and U17528 (N_17528,N_17430,N_17331);
nand U17529 (N_17529,N_17045,N_17345);
and U17530 (N_17530,N_16970,N_16922);
nor U17531 (N_17531,N_17489,N_17050);
xor U17532 (N_17532,N_16972,N_17175);
nor U17533 (N_17533,N_17443,N_17452);
xnor U17534 (N_17534,N_17246,N_17111);
nand U17535 (N_17535,N_16997,N_17312);
or U17536 (N_17536,N_17192,N_17496);
or U17537 (N_17537,N_16955,N_17256);
or U17538 (N_17538,N_17186,N_17089);
xor U17539 (N_17539,N_17173,N_17351);
or U17540 (N_17540,N_17131,N_17434);
and U17541 (N_17541,N_17197,N_17487);
nand U17542 (N_17542,N_17087,N_17259);
nor U17543 (N_17543,N_17486,N_17380);
and U17544 (N_17544,N_17228,N_17008);
or U17545 (N_17545,N_17491,N_17100);
and U17546 (N_17546,N_16945,N_17226);
and U17547 (N_17547,N_17335,N_17262);
and U17548 (N_17548,N_17442,N_17207);
nand U17549 (N_17549,N_17278,N_17342);
xor U17550 (N_17550,N_17381,N_17025);
and U17551 (N_17551,N_17122,N_17357);
nor U17552 (N_17552,N_17356,N_17439);
and U17553 (N_17553,N_17401,N_17332);
and U17554 (N_17554,N_17164,N_17119);
nor U17555 (N_17555,N_17285,N_16999);
or U17556 (N_17556,N_17410,N_17161);
nand U17557 (N_17557,N_17105,N_17420);
nand U17558 (N_17558,N_17037,N_17294);
and U17559 (N_17559,N_17437,N_17080);
xor U17560 (N_17560,N_16879,N_16920);
nand U17561 (N_17561,N_17133,N_17495);
or U17562 (N_17562,N_17147,N_16965);
and U17563 (N_17563,N_16952,N_17140);
xnor U17564 (N_17564,N_17307,N_16925);
nor U17565 (N_17565,N_17063,N_17354);
xor U17566 (N_17566,N_16917,N_17168);
and U17567 (N_17567,N_17267,N_17183);
or U17568 (N_17568,N_17315,N_16967);
and U17569 (N_17569,N_17016,N_17428);
nand U17570 (N_17570,N_17170,N_17438);
or U17571 (N_17571,N_17377,N_17029);
nand U17572 (N_17572,N_17464,N_17473);
or U17573 (N_17573,N_17479,N_16994);
and U17574 (N_17574,N_17276,N_17244);
xor U17575 (N_17575,N_17293,N_16977);
or U17576 (N_17576,N_17426,N_17220);
xor U17577 (N_17577,N_17419,N_16960);
and U17578 (N_17578,N_16905,N_17284);
nor U17579 (N_17579,N_17169,N_17329);
and U17580 (N_17580,N_17039,N_17212);
nor U17581 (N_17581,N_17137,N_17180);
and U17582 (N_17582,N_16969,N_17264);
xor U17583 (N_17583,N_16934,N_16880);
xor U17584 (N_17584,N_17006,N_17453);
nor U17585 (N_17585,N_17138,N_16913);
xor U17586 (N_17586,N_17408,N_16906);
nor U17587 (N_17587,N_17435,N_17166);
nand U17588 (N_17588,N_17152,N_17070);
nor U17589 (N_17589,N_17384,N_17027);
xnor U17590 (N_17590,N_17076,N_17248);
nand U17591 (N_17591,N_17485,N_17313);
xor U17592 (N_17592,N_16961,N_17040);
and U17593 (N_17593,N_17160,N_17238);
and U17594 (N_17594,N_17374,N_17201);
and U17595 (N_17595,N_16963,N_17364);
and U17596 (N_17596,N_16891,N_16939);
xor U17597 (N_17597,N_17305,N_17456);
nor U17598 (N_17598,N_17243,N_17362);
and U17599 (N_17599,N_17360,N_17348);
or U17600 (N_17600,N_17155,N_17013);
and U17601 (N_17601,N_17405,N_17081);
nand U17602 (N_17602,N_17101,N_17072);
and U17603 (N_17603,N_17218,N_17298);
nand U17604 (N_17604,N_17498,N_16940);
or U17605 (N_17605,N_17465,N_17162);
xor U17606 (N_17606,N_17467,N_17071);
xor U17607 (N_17607,N_17157,N_17363);
nor U17608 (N_17608,N_17154,N_17476);
nor U17609 (N_17609,N_16989,N_17454);
nand U17610 (N_17610,N_17250,N_17399);
xnor U17611 (N_17611,N_17222,N_17121);
or U17612 (N_17612,N_17376,N_17459);
xor U17613 (N_17613,N_17407,N_17334);
or U17614 (N_17614,N_17110,N_16936);
xnor U17615 (N_17615,N_16975,N_17083);
nand U17616 (N_17616,N_17432,N_16964);
nor U17617 (N_17617,N_17205,N_17130);
xor U17618 (N_17618,N_17273,N_17242);
or U17619 (N_17619,N_17049,N_17388);
nand U17620 (N_17620,N_17200,N_16895);
and U17621 (N_17621,N_17328,N_17058);
nand U17622 (N_17622,N_17134,N_17463);
xnor U17623 (N_17623,N_17472,N_17382);
xor U17624 (N_17624,N_16896,N_17330);
and U17625 (N_17625,N_17427,N_16902);
nand U17626 (N_17626,N_17224,N_17021);
or U17627 (N_17627,N_17387,N_17094);
and U17628 (N_17628,N_17493,N_16962);
or U17629 (N_17629,N_17118,N_17153);
xnor U17630 (N_17630,N_17340,N_16912);
xnor U17631 (N_17631,N_17150,N_17227);
nand U17632 (N_17632,N_17196,N_16976);
or U17633 (N_17633,N_17249,N_17104);
or U17634 (N_17634,N_17404,N_17341);
and U17635 (N_17635,N_16956,N_17167);
or U17636 (N_17636,N_17423,N_17048);
nand U17637 (N_17637,N_17182,N_17367);
or U17638 (N_17638,N_17457,N_16980);
nor U17639 (N_17639,N_17261,N_17028);
xnor U17640 (N_17640,N_16946,N_17309);
nand U17641 (N_17641,N_17127,N_16968);
nand U17642 (N_17642,N_17093,N_17041);
and U17643 (N_17643,N_17255,N_17068);
nor U17644 (N_17644,N_17191,N_17319);
nor U17645 (N_17645,N_17327,N_17424);
nor U17646 (N_17646,N_16888,N_17017);
or U17647 (N_17647,N_17390,N_16979);
nor U17648 (N_17648,N_17217,N_17106);
nand U17649 (N_17649,N_16993,N_16973);
or U17650 (N_17650,N_17215,N_17316);
nor U17651 (N_17651,N_16890,N_16915);
nand U17652 (N_17652,N_16914,N_16935);
nand U17653 (N_17653,N_17422,N_16899);
nor U17654 (N_17654,N_17339,N_17014);
and U17655 (N_17655,N_17378,N_16941);
xnor U17656 (N_17656,N_17231,N_17299);
xor U17657 (N_17657,N_17252,N_17136);
nand U17658 (N_17658,N_16938,N_17281);
and U17659 (N_17659,N_17296,N_16974);
or U17660 (N_17660,N_17338,N_16921);
nand U17661 (N_17661,N_17251,N_17078);
nor U17662 (N_17662,N_17203,N_17254);
and U17663 (N_17663,N_17300,N_17455);
xor U17664 (N_17664,N_17142,N_17047);
xor U17665 (N_17665,N_17084,N_16923);
or U17666 (N_17666,N_17322,N_17086);
nand U17667 (N_17667,N_17051,N_17092);
and U17668 (N_17668,N_17337,N_17269);
and U17669 (N_17669,N_17002,N_17120);
or U17670 (N_17670,N_16893,N_16919);
or U17671 (N_17671,N_17394,N_17159);
nor U17672 (N_17672,N_17326,N_17210);
and U17673 (N_17673,N_17074,N_17241);
nand U17674 (N_17674,N_17035,N_17425);
and U17675 (N_17675,N_17245,N_17235);
nand U17676 (N_17676,N_17409,N_16995);
or U17677 (N_17677,N_16886,N_17209);
or U17678 (N_17678,N_16918,N_17445);
xnor U17679 (N_17679,N_17321,N_17414);
nor U17680 (N_17680,N_16987,N_17302);
xor U17681 (N_17681,N_17283,N_17373);
or U17682 (N_17682,N_17184,N_16996);
nor U17683 (N_17683,N_17151,N_17415);
or U17684 (N_17684,N_17303,N_16898);
or U17685 (N_17685,N_17194,N_17469);
xor U17686 (N_17686,N_16904,N_17274);
xnor U17687 (N_17687,N_16981,N_17477);
nor U17688 (N_17688,N_17441,N_16985);
and U17689 (N_17689,N_17004,N_17075);
and U17690 (N_17690,N_17123,N_17032);
or U17691 (N_17691,N_16885,N_17350);
nor U17692 (N_17692,N_17352,N_17369);
nor U17693 (N_17693,N_16966,N_17471);
or U17694 (N_17694,N_17065,N_17462);
or U17695 (N_17695,N_17097,N_17343);
nor U17696 (N_17696,N_16986,N_17336);
and U17697 (N_17697,N_17204,N_17188);
nand U17698 (N_17698,N_17418,N_17010);
or U17699 (N_17699,N_17124,N_17451);
nand U17700 (N_17700,N_17126,N_17190);
nand U17701 (N_17701,N_17024,N_17481);
or U17702 (N_17702,N_16881,N_17208);
xnor U17703 (N_17703,N_17125,N_17213);
xnor U17704 (N_17704,N_17280,N_17450);
xnor U17705 (N_17705,N_17007,N_17411);
or U17706 (N_17706,N_16901,N_17088);
xor U17707 (N_17707,N_16884,N_17143);
xnor U17708 (N_17708,N_16889,N_17011);
nand U17709 (N_17709,N_17042,N_17279);
nand U17710 (N_17710,N_17193,N_17026);
xor U17711 (N_17711,N_17091,N_17272);
nand U17712 (N_17712,N_16957,N_16947);
and U17713 (N_17713,N_17234,N_17402);
or U17714 (N_17714,N_17053,N_17385);
nand U17715 (N_17715,N_17361,N_16950);
nand U17716 (N_17716,N_17292,N_17109);
nor U17717 (N_17717,N_17240,N_17230);
nand U17718 (N_17718,N_17141,N_17233);
and U17719 (N_17719,N_17023,N_17311);
xor U17720 (N_17720,N_17349,N_16943);
and U17721 (N_17721,N_17440,N_17368);
nor U17722 (N_17722,N_17031,N_17055);
and U17723 (N_17723,N_17397,N_17478);
and U17724 (N_17724,N_17172,N_17325);
nand U17725 (N_17725,N_17206,N_17366);
nand U17726 (N_17726,N_17358,N_17066);
nor U17727 (N_17727,N_16877,N_17494);
nand U17728 (N_17728,N_16984,N_17112);
nand U17729 (N_17729,N_17379,N_17223);
nor U17730 (N_17730,N_17199,N_17038);
and U17731 (N_17731,N_17114,N_17108);
and U17732 (N_17732,N_16992,N_16927);
nand U17733 (N_17733,N_17344,N_17412);
and U17734 (N_17734,N_17054,N_16908);
nand U17735 (N_17735,N_17490,N_17413);
nand U17736 (N_17736,N_17012,N_17492);
nor U17737 (N_17737,N_17461,N_17444);
nand U17738 (N_17738,N_17482,N_17468);
and U17739 (N_17739,N_17018,N_16911);
xnor U17740 (N_17740,N_17431,N_17033);
xnor U17741 (N_17741,N_17019,N_17346);
xnor U17742 (N_17742,N_17306,N_17365);
xor U17743 (N_17743,N_16892,N_17288);
xor U17744 (N_17744,N_17317,N_17132);
nand U17745 (N_17745,N_17034,N_17102);
and U17746 (N_17746,N_17148,N_17056);
nand U17747 (N_17747,N_17158,N_17177);
and U17748 (N_17748,N_16907,N_17043);
nand U17749 (N_17749,N_17416,N_17044);
nor U17750 (N_17750,N_17258,N_17001);
xor U17751 (N_17751,N_17189,N_17287);
nand U17752 (N_17752,N_16929,N_16937);
nand U17753 (N_17753,N_17145,N_16951);
nor U17754 (N_17754,N_17052,N_17069);
nand U17755 (N_17755,N_17386,N_17389);
and U17756 (N_17756,N_17400,N_17181);
or U17757 (N_17757,N_17297,N_16954);
or U17758 (N_17758,N_17266,N_17253);
nand U17759 (N_17759,N_17176,N_17171);
or U17760 (N_17760,N_17128,N_16983);
nand U17761 (N_17761,N_16928,N_16971);
nor U17762 (N_17762,N_16942,N_17185);
xnor U17763 (N_17763,N_17403,N_17020);
or U17764 (N_17764,N_16931,N_17286);
nand U17765 (N_17765,N_17000,N_17064);
nor U17766 (N_17766,N_17301,N_17077);
or U17767 (N_17767,N_17448,N_17009);
and U17768 (N_17768,N_17271,N_16903);
xor U17769 (N_17769,N_17395,N_17082);
nor U17770 (N_17770,N_17219,N_17421);
nand U17771 (N_17771,N_17396,N_17277);
nor U17772 (N_17772,N_17398,N_16958);
or U17773 (N_17773,N_17067,N_16894);
xor U17774 (N_17774,N_17383,N_17178);
nor U17775 (N_17775,N_17475,N_17371);
nor U17776 (N_17776,N_16882,N_17260);
nand U17777 (N_17777,N_17062,N_17393);
nor U17778 (N_17778,N_17484,N_17433);
xnor U17779 (N_17779,N_16916,N_17221);
nand U17780 (N_17780,N_17458,N_17113);
xnor U17781 (N_17781,N_17195,N_17211);
xor U17782 (N_17782,N_17359,N_17247);
nand U17783 (N_17783,N_17295,N_17265);
and U17784 (N_17784,N_17275,N_17470);
and U17785 (N_17785,N_17347,N_17061);
and U17786 (N_17786,N_17187,N_17406);
or U17787 (N_17787,N_17268,N_16930);
and U17788 (N_17788,N_17198,N_17060);
nand U17789 (N_17789,N_16909,N_17429);
xnor U17790 (N_17790,N_16900,N_17291);
xor U17791 (N_17791,N_16990,N_16959);
nand U17792 (N_17792,N_17480,N_17059);
xor U17793 (N_17793,N_17156,N_17282);
or U17794 (N_17794,N_17304,N_17466);
nand U17795 (N_17795,N_17129,N_16978);
nor U17796 (N_17796,N_17318,N_17417);
nand U17797 (N_17797,N_17308,N_17179);
or U17798 (N_17798,N_16991,N_16926);
nor U17799 (N_17799,N_17323,N_17289);
nor U17800 (N_17800,N_17499,N_17090);
nand U17801 (N_17801,N_17099,N_17446);
nand U17802 (N_17802,N_17263,N_17015);
nor U17803 (N_17803,N_16932,N_17103);
and U17804 (N_17804,N_17333,N_16933);
or U17805 (N_17805,N_17436,N_17290);
and U17806 (N_17806,N_16897,N_17314);
and U17807 (N_17807,N_16948,N_17139);
nand U17808 (N_17808,N_17163,N_17005);
nor U17809 (N_17809,N_17375,N_17149);
or U17810 (N_17810,N_17115,N_17079);
nor U17811 (N_17811,N_16887,N_16953);
or U17812 (N_17812,N_17085,N_17291);
or U17813 (N_17813,N_17445,N_17229);
and U17814 (N_17814,N_17215,N_17192);
and U17815 (N_17815,N_17395,N_16978);
nor U17816 (N_17816,N_17145,N_17056);
xor U17817 (N_17817,N_17175,N_17191);
nand U17818 (N_17818,N_16976,N_16975);
xor U17819 (N_17819,N_16891,N_16953);
and U17820 (N_17820,N_17246,N_17033);
and U17821 (N_17821,N_16950,N_16933);
xor U17822 (N_17822,N_17460,N_16939);
nand U17823 (N_17823,N_17439,N_17170);
or U17824 (N_17824,N_17350,N_17424);
xor U17825 (N_17825,N_17232,N_17178);
and U17826 (N_17826,N_16960,N_16943);
or U17827 (N_17827,N_17017,N_17472);
or U17828 (N_17828,N_17388,N_17019);
and U17829 (N_17829,N_17060,N_17015);
or U17830 (N_17830,N_17435,N_17492);
nor U17831 (N_17831,N_16928,N_17264);
or U17832 (N_17832,N_16917,N_17052);
xnor U17833 (N_17833,N_17227,N_17055);
nand U17834 (N_17834,N_16974,N_17280);
nor U17835 (N_17835,N_17098,N_17107);
xor U17836 (N_17836,N_17299,N_17377);
or U17837 (N_17837,N_17029,N_16936);
xnor U17838 (N_17838,N_17329,N_17373);
nand U17839 (N_17839,N_17302,N_17282);
nand U17840 (N_17840,N_17445,N_17105);
and U17841 (N_17841,N_17418,N_16915);
and U17842 (N_17842,N_16964,N_17239);
and U17843 (N_17843,N_17221,N_17282);
nor U17844 (N_17844,N_17004,N_17475);
and U17845 (N_17845,N_17082,N_16967);
and U17846 (N_17846,N_16937,N_17259);
xor U17847 (N_17847,N_17006,N_17174);
xor U17848 (N_17848,N_16946,N_17221);
or U17849 (N_17849,N_17019,N_17130);
nor U17850 (N_17850,N_17108,N_17467);
and U17851 (N_17851,N_17336,N_16939);
and U17852 (N_17852,N_17159,N_17161);
and U17853 (N_17853,N_17190,N_16892);
or U17854 (N_17854,N_17321,N_17315);
nand U17855 (N_17855,N_17398,N_17325);
and U17856 (N_17856,N_16974,N_17427);
and U17857 (N_17857,N_17242,N_17488);
or U17858 (N_17858,N_17466,N_17063);
xor U17859 (N_17859,N_17470,N_17294);
or U17860 (N_17860,N_16913,N_17095);
and U17861 (N_17861,N_17349,N_17485);
xnor U17862 (N_17862,N_17054,N_17129);
xor U17863 (N_17863,N_16996,N_17478);
or U17864 (N_17864,N_17045,N_17316);
and U17865 (N_17865,N_17032,N_17252);
and U17866 (N_17866,N_17139,N_16994);
nand U17867 (N_17867,N_17448,N_17039);
nor U17868 (N_17868,N_17050,N_17081);
xor U17869 (N_17869,N_17190,N_17290);
and U17870 (N_17870,N_16891,N_17325);
nand U17871 (N_17871,N_17304,N_16892);
xor U17872 (N_17872,N_17237,N_16971);
nor U17873 (N_17873,N_17086,N_17177);
xor U17874 (N_17874,N_17032,N_17231);
xnor U17875 (N_17875,N_17486,N_17370);
xnor U17876 (N_17876,N_16987,N_17487);
or U17877 (N_17877,N_17301,N_17441);
nand U17878 (N_17878,N_17245,N_17287);
and U17879 (N_17879,N_17220,N_16926);
or U17880 (N_17880,N_17452,N_17498);
nand U17881 (N_17881,N_17185,N_17026);
nor U17882 (N_17882,N_17017,N_17256);
nor U17883 (N_17883,N_17223,N_17368);
and U17884 (N_17884,N_17447,N_16965);
nor U17885 (N_17885,N_17134,N_17269);
or U17886 (N_17886,N_17075,N_17168);
and U17887 (N_17887,N_16984,N_17006);
nand U17888 (N_17888,N_16970,N_16897);
or U17889 (N_17889,N_17212,N_17210);
or U17890 (N_17890,N_17395,N_17038);
nor U17891 (N_17891,N_17124,N_17420);
nor U17892 (N_17892,N_17177,N_17330);
or U17893 (N_17893,N_17293,N_17359);
or U17894 (N_17894,N_16927,N_17119);
nor U17895 (N_17895,N_17168,N_16925);
and U17896 (N_17896,N_17499,N_17486);
or U17897 (N_17897,N_17092,N_17352);
or U17898 (N_17898,N_16984,N_17353);
nand U17899 (N_17899,N_17203,N_17418);
nand U17900 (N_17900,N_17435,N_17447);
nand U17901 (N_17901,N_17298,N_17052);
nand U17902 (N_17902,N_17245,N_17283);
or U17903 (N_17903,N_17182,N_17099);
nor U17904 (N_17904,N_17291,N_17325);
or U17905 (N_17905,N_16986,N_17140);
xor U17906 (N_17906,N_16920,N_17295);
nand U17907 (N_17907,N_17249,N_17338);
nor U17908 (N_17908,N_17247,N_17204);
xor U17909 (N_17909,N_16997,N_17141);
xor U17910 (N_17910,N_16947,N_17300);
and U17911 (N_17911,N_17400,N_17066);
xnor U17912 (N_17912,N_17198,N_17126);
and U17913 (N_17913,N_17407,N_17283);
nand U17914 (N_17914,N_17321,N_17292);
nand U17915 (N_17915,N_16875,N_16970);
nand U17916 (N_17916,N_17319,N_17189);
nor U17917 (N_17917,N_17425,N_17082);
and U17918 (N_17918,N_17494,N_17310);
xnor U17919 (N_17919,N_16898,N_17460);
and U17920 (N_17920,N_17140,N_17125);
nor U17921 (N_17921,N_16890,N_17181);
nor U17922 (N_17922,N_17010,N_17367);
nand U17923 (N_17923,N_17324,N_17071);
nand U17924 (N_17924,N_17498,N_16978);
nand U17925 (N_17925,N_17109,N_16967);
xnor U17926 (N_17926,N_16904,N_17344);
and U17927 (N_17927,N_17015,N_17456);
nor U17928 (N_17928,N_17193,N_17466);
or U17929 (N_17929,N_17400,N_16963);
nor U17930 (N_17930,N_17202,N_16898);
nor U17931 (N_17931,N_17258,N_17262);
nor U17932 (N_17932,N_17267,N_17211);
and U17933 (N_17933,N_16926,N_17457);
nor U17934 (N_17934,N_17432,N_17282);
nand U17935 (N_17935,N_17263,N_16886);
xor U17936 (N_17936,N_17300,N_17197);
nand U17937 (N_17937,N_17231,N_17256);
or U17938 (N_17938,N_17282,N_17174);
nand U17939 (N_17939,N_17358,N_16952);
xnor U17940 (N_17940,N_17242,N_17393);
or U17941 (N_17941,N_17211,N_17247);
nor U17942 (N_17942,N_17211,N_17202);
xnor U17943 (N_17943,N_16992,N_17234);
nor U17944 (N_17944,N_17474,N_16883);
nand U17945 (N_17945,N_17245,N_16927);
xor U17946 (N_17946,N_17046,N_17127);
nand U17947 (N_17947,N_17218,N_17159);
nor U17948 (N_17948,N_17498,N_17014);
nand U17949 (N_17949,N_17023,N_17042);
or U17950 (N_17950,N_17107,N_17380);
or U17951 (N_17951,N_17009,N_17233);
and U17952 (N_17952,N_17331,N_17008);
nor U17953 (N_17953,N_17043,N_17027);
or U17954 (N_17954,N_17290,N_17480);
or U17955 (N_17955,N_17246,N_16922);
nand U17956 (N_17956,N_17050,N_16875);
and U17957 (N_17957,N_17385,N_16935);
and U17958 (N_17958,N_17099,N_17413);
or U17959 (N_17959,N_17266,N_17103);
nor U17960 (N_17960,N_17297,N_17175);
xor U17961 (N_17961,N_17429,N_16918);
nor U17962 (N_17962,N_16909,N_17307);
or U17963 (N_17963,N_17053,N_17340);
and U17964 (N_17964,N_17016,N_16875);
or U17965 (N_17965,N_17463,N_16885);
or U17966 (N_17966,N_17036,N_17394);
and U17967 (N_17967,N_17211,N_17341);
nand U17968 (N_17968,N_16885,N_17007);
and U17969 (N_17969,N_16877,N_17215);
xnor U17970 (N_17970,N_17189,N_17472);
nor U17971 (N_17971,N_17392,N_17403);
nand U17972 (N_17972,N_16979,N_17469);
or U17973 (N_17973,N_17213,N_17272);
or U17974 (N_17974,N_16948,N_17414);
and U17975 (N_17975,N_16890,N_17234);
xor U17976 (N_17976,N_17268,N_17223);
xnor U17977 (N_17977,N_17451,N_17409);
xor U17978 (N_17978,N_17447,N_17365);
nand U17979 (N_17979,N_17129,N_17000);
or U17980 (N_17980,N_17168,N_17280);
or U17981 (N_17981,N_16994,N_17488);
nand U17982 (N_17982,N_17315,N_17039);
or U17983 (N_17983,N_17359,N_16930);
nor U17984 (N_17984,N_17255,N_17242);
nor U17985 (N_17985,N_17435,N_17305);
xnor U17986 (N_17986,N_17402,N_17476);
and U17987 (N_17987,N_17204,N_16912);
xor U17988 (N_17988,N_17383,N_16922);
or U17989 (N_17989,N_16947,N_17172);
nor U17990 (N_17990,N_17464,N_17381);
nor U17991 (N_17991,N_17456,N_16939);
xnor U17992 (N_17992,N_17168,N_16984);
xor U17993 (N_17993,N_17148,N_17207);
or U17994 (N_17994,N_17446,N_17307);
or U17995 (N_17995,N_17150,N_17372);
nor U17996 (N_17996,N_16960,N_17183);
nand U17997 (N_17997,N_17324,N_16896);
or U17998 (N_17998,N_17234,N_17467);
xnor U17999 (N_17999,N_17057,N_17273);
xor U18000 (N_18000,N_17235,N_17417);
xor U18001 (N_18001,N_16992,N_16953);
nor U18002 (N_18002,N_16984,N_16881);
nor U18003 (N_18003,N_17171,N_16937);
nor U18004 (N_18004,N_17479,N_17092);
nor U18005 (N_18005,N_16993,N_17181);
nand U18006 (N_18006,N_17485,N_16892);
xnor U18007 (N_18007,N_17450,N_17438);
nand U18008 (N_18008,N_16954,N_17027);
nand U18009 (N_18009,N_17264,N_16937);
or U18010 (N_18010,N_16956,N_17494);
nor U18011 (N_18011,N_17306,N_16887);
or U18012 (N_18012,N_16957,N_17311);
xnor U18013 (N_18013,N_16972,N_17321);
nor U18014 (N_18014,N_17226,N_16929);
nand U18015 (N_18015,N_17413,N_17164);
xor U18016 (N_18016,N_16939,N_17127);
or U18017 (N_18017,N_16918,N_17351);
and U18018 (N_18018,N_17458,N_17313);
and U18019 (N_18019,N_17480,N_17250);
xnor U18020 (N_18020,N_17428,N_17112);
or U18021 (N_18021,N_16956,N_16959);
or U18022 (N_18022,N_17370,N_17081);
or U18023 (N_18023,N_17087,N_17171);
and U18024 (N_18024,N_17225,N_17217);
and U18025 (N_18025,N_17135,N_16939);
xor U18026 (N_18026,N_17478,N_16928);
xnor U18027 (N_18027,N_17050,N_16915);
xor U18028 (N_18028,N_16909,N_17028);
nor U18029 (N_18029,N_17155,N_16917);
xor U18030 (N_18030,N_17192,N_17155);
or U18031 (N_18031,N_17415,N_16976);
or U18032 (N_18032,N_17185,N_17114);
xor U18033 (N_18033,N_17406,N_16915);
or U18034 (N_18034,N_17072,N_17106);
nand U18035 (N_18035,N_17139,N_16953);
nand U18036 (N_18036,N_17237,N_16882);
nand U18037 (N_18037,N_17103,N_16877);
or U18038 (N_18038,N_17301,N_17305);
or U18039 (N_18039,N_17067,N_17489);
nand U18040 (N_18040,N_17090,N_17036);
and U18041 (N_18041,N_17139,N_17039);
xnor U18042 (N_18042,N_17005,N_17052);
or U18043 (N_18043,N_17358,N_17086);
xor U18044 (N_18044,N_17228,N_17420);
nand U18045 (N_18045,N_17045,N_17429);
nand U18046 (N_18046,N_17001,N_17328);
nand U18047 (N_18047,N_17065,N_17070);
xnor U18048 (N_18048,N_16944,N_17161);
nor U18049 (N_18049,N_17324,N_17024);
or U18050 (N_18050,N_17462,N_17370);
or U18051 (N_18051,N_17254,N_17303);
or U18052 (N_18052,N_17333,N_17298);
or U18053 (N_18053,N_16939,N_17060);
nand U18054 (N_18054,N_17272,N_16977);
or U18055 (N_18055,N_17288,N_16903);
nand U18056 (N_18056,N_17209,N_17249);
nor U18057 (N_18057,N_17181,N_17477);
or U18058 (N_18058,N_17287,N_17425);
and U18059 (N_18059,N_17260,N_17203);
nor U18060 (N_18060,N_17286,N_17342);
or U18061 (N_18061,N_17435,N_17381);
xor U18062 (N_18062,N_17401,N_17304);
xnor U18063 (N_18063,N_17098,N_17000);
xnor U18064 (N_18064,N_16895,N_17461);
and U18065 (N_18065,N_17028,N_17035);
nand U18066 (N_18066,N_16928,N_17429);
and U18067 (N_18067,N_16914,N_17162);
and U18068 (N_18068,N_17353,N_17434);
xor U18069 (N_18069,N_17234,N_17045);
nor U18070 (N_18070,N_17127,N_17426);
xnor U18071 (N_18071,N_17253,N_17280);
and U18072 (N_18072,N_16897,N_17116);
nand U18073 (N_18073,N_17220,N_17264);
and U18074 (N_18074,N_17340,N_17387);
nand U18075 (N_18075,N_16949,N_17297);
xnor U18076 (N_18076,N_17086,N_17347);
nor U18077 (N_18077,N_17260,N_17181);
nand U18078 (N_18078,N_17444,N_17117);
nand U18079 (N_18079,N_16961,N_17162);
nand U18080 (N_18080,N_16960,N_17155);
or U18081 (N_18081,N_17135,N_16910);
xnor U18082 (N_18082,N_17392,N_17070);
or U18083 (N_18083,N_16985,N_17045);
and U18084 (N_18084,N_17096,N_16925);
nand U18085 (N_18085,N_17004,N_17284);
nor U18086 (N_18086,N_17422,N_17273);
xor U18087 (N_18087,N_17339,N_17384);
nand U18088 (N_18088,N_16986,N_17213);
xnor U18089 (N_18089,N_17458,N_17166);
nor U18090 (N_18090,N_17039,N_17241);
nand U18091 (N_18091,N_17239,N_17151);
and U18092 (N_18092,N_17389,N_17113);
xor U18093 (N_18093,N_17063,N_17368);
nor U18094 (N_18094,N_17439,N_16940);
nand U18095 (N_18095,N_17478,N_17449);
or U18096 (N_18096,N_16892,N_17105);
or U18097 (N_18097,N_17247,N_17038);
and U18098 (N_18098,N_16882,N_17407);
and U18099 (N_18099,N_16946,N_17370);
xor U18100 (N_18100,N_17063,N_17169);
xor U18101 (N_18101,N_17465,N_17072);
nand U18102 (N_18102,N_17180,N_17057);
nand U18103 (N_18103,N_17189,N_17229);
xnor U18104 (N_18104,N_17004,N_16951);
nor U18105 (N_18105,N_17053,N_16892);
nor U18106 (N_18106,N_16996,N_17036);
and U18107 (N_18107,N_17358,N_17444);
or U18108 (N_18108,N_16876,N_17045);
or U18109 (N_18109,N_17047,N_17095);
nand U18110 (N_18110,N_17383,N_17278);
or U18111 (N_18111,N_17484,N_17256);
nor U18112 (N_18112,N_17206,N_17322);
xor U18113 (N_18113,N_17295,N_16921);
nand U18114 (N_18114,N_17064,N_17037);
nor U18115 (N_18115,N_17000,N_17204);
and U18116 (N_18116,N_17412,N_17335);
nor U18117 (N_18117,N_17072,N_17438);
nor U18118 (N_18118,N_17131,N_17071);
nor U18119 (N_18119,N_17166,N_17223);
nand U18120 (N_18120,N_16967,N_17252);
and U18121 (N_18121,N_16877,N_17379);
or U18122 (N_18122,N_17008,N_16986);
and U18123 (N_18123,N_17454,N_16988);
xnor U18124 (N_18124,N_17268,N_16959);
nor U18125 (N_18125,N_18063,N_18046);
nor U18126 (N_18126,N_17675,N_17619);
xnor U18127 (N_18127,N_18079,N_17722);
and U18128 (N_18128,N_17660,N_17543);
nand U18129 (N_18129,N_17756,N_17652);
nand U18130 (N_18130,N_17970,N_17538);
or U18131 (N_18131,N_17642,N_18039);
or U18132 (N_18132,N_17672,N_18003);
xnor U18133 (N_18133,N_17686,N_17841);
and U18134 (N_18134,N_18076,N_18037);
nor U18135 (N_18135,N_17731,N_17522);
or U18136 (N_18136,N_17968,N_18027);
or U18137 (N_18137,N_18070,N_17744);
xor U18138 (N_18138,N_17516,N_17935);
nand U18139 (N_18139,N_17825,N_17567);
nor U18140 (N_18140,N_17762,N_17618);
nor U18141 (N_18141,N_18058,N_18098);
and U18142 (N_18142,N_17990,N_17822);
or U18143 (N_18143,N_17526,N_17565);
and U18144 (N_18144,N_17629,N_17859);
and U18145 (N_18145,N_17942,N_17773);
nand U18146 (N_18146,N_17662,N_17930);
nand U18147 (N_18147,N_17816,N_17668);
nand U18148 (N_18148,N_17853,N_17902);
nor U18149 (N_18149,N_17546,N_17913);
xnor U18150 (N_18150,N_17715,N_17589);
or U18151 (N_18151,N_17533,N_18056);
or U18152 (N_18152,N_17626,N_17614);
xor U18153 (N_18153,N_17885,N_17837);
nand U18154 (N_18154,N_17509,N_17803);
and U18155 (N_18155,N_18018,N_17698);
xnor U18156 (N_18156,N_17949,N_17860);
xnor U18157 (N_18157,N_17922,N_18089);
xnor U18158 (N_18158,N_17702,N_17513);
xnor U18159 (N_18159,N_17824,N_17745);
or U18160 (N_18160,N_17600,N_17800);
and U18161 (N_18161,N_17937,N_17836);
xnor U18162 (N_18162,N_17921,N_18095);
or U18163 (N_18163,N_17880,N_17839);
nor U18164 (N_18164,N_18080,N_17601);
or U18165 (N_18165,N_18114,N_17973);
or U18166 (N_18166,N_18028,N_17764);
or U18167 (N_18167,N_18106,N_17569);
and U18168 (N_18168,N_17563,N_18066);
and U18169 (N_18169,N_17624,N_17786);
nand U18170 (N_18170,N_17977,N_17527);
nor U18171 (N_18171,N_17828,N_18074);
or U18172 (N_18172,N_17594,N_18030);
xor U18173 (N_18173,N_17713,N_18062);
xor U18174 (N_18174,N_17988,N_17732);
nor U18175 (N_18175,N_17950,N_17632);
nand U18176 (N_18176,N_18049,N_18118);
nand U18177 (N_18177,N_17669,N_17793);
nand U18178 (N_18178,N_17718,N_17573);
and U18179 (N_18179,N_18085,N_18024);
or U18180 (N_18180,N_17708,N_18059);
and U18181 (N_18181,N_18048,N_17939);
nor U18182 (N_18182,N_17647,N_17821);
xor U18183 (N_18183,N_17597,N_17808);
or U18184 (N_18184,N_17879,N_17650);
xor U18185 (N_18185,N_18105,N_17651);
xor U18186 (N_18186,N_17654,N_17925);
xnor U18187 (N_18187,N_17893,N_17799);
xor U18188 (N_18188,N_18026,N_17905);
nor U18189 (N_18189,N_17842,N_17831);
nor U18190 (N_18190,N_17891,N_17749);
or U18191 (N_18191,N_17870,N_17814);
and U18192 (N_18192,N_17792,N_18022);
or U18193 (N_18193,N_17911,N_18033);
xnor U18194 (N_18194,N_17646,N_17528);
nor U18195 (N_18195,N_17941,N_17603);
nor U18196 (N_18196,N_17738,N_17863);
or U18197 (N_18197,N_17735,N_18086);
or U18198 (N_18198,N_17906,N_17625);
or U18199 (N_18199,N_18064,N_17709);
nor U18200 (N_18200,N_17572,N_17818);
and U18201 (N_18201,N_17975,N_17953);
xnor U18202 (N_18202,N_17524,N_17641);
xor U18203 (N_18203,N_17701,N_18023);
nand U18204 (N_18204,N_17697,N_17734);
and U18205 (N_18205,N_17720,N_17552);
nand U18206 (N_18206,N_17932,N_17856);
and U18207 (N_18207,N_17653,N_17520);
and U18208 (N_18208,N_17986,N_17785);
nor U18209 (N_18209,N_17826,N_17894);
xor U18210 (N_18210,N_18120,N_17789);
and U18211 (N_18211,N_17500,N_18099);
xnor U18212 (N_18212,N_17918,N_17945);
xor U18213 (N_18213,N_17804,N_17574);
nor U18214 (N_18214,N_18044,N_17717);
xnor U18215 (N_18215,N_17768,N_17840);
nor U18216 (N_18216,N_17907,N_18013);
or U18217 (N_18217,N_17562,N_17959);
nor U18218 (N_18218,N_17501,N_17615);
and U18219 (N_18219,N_17750,N_17983);
xor U18220 (N_18220,N_18014,N_17888);
xnor U18221 (N_18221,N_18020,N_17895);
xnor U18222 (N_18222,N_17802,N_17725);
nand U18223 (N_18223,N_18052,N_17924);
and U18224 (N_18224,N_17743,N_17502);
xnor U18225 (N_18225,N_17636,N_17577);
xor U18226 (N_18226,N_18008,N_17820);
xnor U18227 (N_18227,N_17693,N_17705);
xnor U18228 (N_18228,N_17515,N_17628);
xnor U18229 (N_18229,N_17663,N_17833);
xor U18230 (N_18230,N_17790,N_18097);
nor U18231 (N_18231,N_17873,N_17881);
nor U18232 (N_18232,N_18112,N_17747);
or U18233 (N_18233,N_17736,N_17550);
or U18234 (N_18234,N_17598,N_17557);
xnor U18235 (N_18235,N_17759,N_17781);
nand U18236 (N_18236,N_17690,N_18035);
nand U18237 (N_18237,N_17882,N_17523);
nand U18238 (N_18238,N_17613,N_18122);
nor U18239 (N_18239,N_17834,N_17583);
nor U18240 (N_18240,N_17761,N_17637);
nor U18241 (N_18241,N_17706,N_17716);
nand U18242 (N_18242,N_18111,N_17537);
or U18243 (N_18243,N_17956,N_17580);
nor U18244 (N_18244,N_17723,N_17846);
nor U18245 (N_18245,N_17805,N_18040);
nor U18246 (N_18246,N_17691,N_17696);
xor U18247 (N_18247,N_17612,N_17605);
and U18248 (N_18248,N_17724,N_17769);
or U18249 (N_18249,N_17689,N_17687);
xnor U18250 (N_18250,N_17917,N_17938);
nor U18251 (N_18251,N_17964,N_18081);
nand U18252 (N_18252,N_17585,N_17763);
nand U18253 (N_18253,N_18042,N_17634);
xor U18254 (N_18254,N_17620,N_18088);
xor U18255 (N_18255,N_17780,N_18041);
and U18256 (N_18256,N_17511,N_17984);
nor U18257 (N_18257,N_17962,N_17829);
nor U18258 (N_18258,N_17517,N_17965);
xnor U18259 (N_18259,N_17510,N_17684);
and U18260 (N_18260,N_17755,N_17754);
nand U18261 (N_18261,N_17643,N_18007);
or U18262 (N_18262,N_17599,N_17787);
and U18263 (N_18263,N_17621,N_17532);
and U18264 (N_18264,N_17765,N_17928);
and U18265 (N_18265,N_17794,N_17998);
or U18266 (N_18266,N_17685,N_17807);
nand U18267 (N_18267,N_17877,N_17823);
xor U18268 (N_18268,N_17994,N_17946);
and U18269 (N_18269,N_17919,N_17931);
and U18270 (N_18270,N_18082,N_18104);
xor U18271 (N_18271,N_17929,N_17608);
xor U18272 (N_18272,N_18102,N_17832);
nand U18273 (N_18273,N_18060,N_17779);
nor U18274 (N_18274,N_17817,N_17739);
and U18275 (N_18275,N_17887,N_18107);
nand U18276 (N_18276,N_17700,N_17561);
or U18277 (N_18277,N_17575,N_17933);
nor U18278 (N_18278,N_17954,N_17982);
or U18279 (N_18279,N_17976,N_17967);
xnor U18280 (N_18280,N_17665,N_17566);
nand U18281 (N_18281,N_18121,N_17812);
nor U18282 (N_18282,N_17943,N_17506);
and U18283 (N_18283,N_17751,N_17910);
nand U18284 (N_18284,N_18077,N_18015);
xor U18285 (N_18285,N_17867,N_17661);
nand U18286 (N_18286,N_17627,N_18025);
nor U18287 (N_18287,N_17896,N_17886);
nor U18288 (N_18288,N_17596,N_17568);
xor U18289 (N_18289,N_17541,N_17678);
xor U18290 (N_18290,N_17767,N_17852);
and U18291 (N_18291,N_17850,N_17948);
and U18292 (N_18292,N_17923,N_17649);
or U18293 (N_18293,N_17507,N_17656);
xnor U18294 (N_18294,N_17901,N_18010);
nand U18295 (N_18295,N_17578,N_18031);
nand U18296 (N_18296,N_17971,N_18053);
or U18297 (N_18297,N_18054,N_17554);
or U18298 (N_18298,N_17677,N_17866);
xnor U18299 (N_18299,N_17726,N_17940);
xor U18300 (N_18300,N_18071,N_17843);
and U18301 (N_18301,N_18115,N_17536);
and U18302 (N_18302,N_17904,N_17679);
nand U18303 (N_18303,N_17555,N_17581);
and U18304 (N_18304,N_17875,N_17991);
or U18305 (N_18305,N_17707,N_17584);
xnor U18306 (N_18306,N_18075,N_17878);
and U18307 (N_18307,N_17951,N_17947);
nor U18308 (N_18308,N_17771,N_17784);
nor U18309 (N_18309,N_17512,N_18043);
xor U18310 (N_18310,N_17861,N_17996);
nor U18311 (N_18311,N_17728,N_17957);
or U18312 (N_18312,N_17611,N_17748);
nor U18313 (N_18313,N_18055,N_17576);
or U18314 (N_18314,N_17635,N_17559);
nand U18315 (N_18315,N_17908,N_18061);
or U18316 (N_18316,N_17876,N_18032);
or U18317 (N_18317,N_17903,N_17884);
and U18318 (N_18318,N_17556,N_17809);
nor U18319 (N_18319,N_18038,N_17855);
nand U18320 (N_18320,N_18029,N_17871);
and U18321 (N_18321,N_17892,N_17529);
nand U18322 (N_18322,N_17609,N_17733);
and U18323 (N_18323,N_17710,N_17737);
xnor U18324 (N_18324,N_17631,N_18057);
xor U18325 (N_18325,N_17796,N_17999);
nand U18326 (N_18326,N_17980,N_17992);
nand U18327 (N_18327,N_17838,N_17978);
and U18328 (N_18328,N_17934,N_17997);
nor U18329 (N_18329,N_18069,N_17508);
nor U18330 (N_18330,N_17848,N_18017);
or U18331 (N_18331,N_17570,N_17798);
or U18332 (N_18332,N_17530,N_18051);
xor U18333 (N_18333,N_18002,N_17847);
and U18334 (N_18334,N_18109,N_17757);
nand U18335 (N_18335,N_17727,N_17670);
xor U18336 (N_18336,N_17741,N_17633);
nor U18337 (N_18337,N_17606,N_17595);
nand U18338 (N_18338,N_17858,N_17591);
or U18339 (N_18339,N_18065,N_17760);
nor U18340 (N_18340,N_17810,N_18011);
or U18341 (N_18341,N_17806,N_17827);
nor U18342 (N_18342,N_18016,N_17699);
and U18343 (N_18343,N_17682,N_17897);
nand U18344 (N_18344,N_17545,N_17914);
nand U18345 (N_18345,N_17961,N_17658);
or U18346 (N_18346,N_17915,N_17638);
nor U18347 (N_18347,N_17695,N_17503);
nor U18348 (N_18348,N_17872,N_17645);
and U18349 (N_18349,N_17714,N_17582);
and U18350 (N_18350,N_18119,N_18034);
xnor U18351 (N_18351,N_17519,N_17776);
and U18352 (N_18352,N_17927,N_17955);
xor U18353 (N_18353,N_18117,N_17740);
nor U18354 (N_18354,N_17518,N_17666);
nand U18355 (N_18355,N_18068,N_18084);
xnor U18356 (N_18356,N_18019,N_17900);
xnor U18357 (N_18357,N_17766,N_17674);
or U18358 (N_18358,N_17788,N_18000);
or U18359 (N_18359,N_17644,N_17610);
or U18360 (N_18360,N_18078,N_17680);
xnor U18361 (N_18361,N_17630,N_17958);
nand U18362 (N_18362,N_17936,N_17558);
xnor U18363 (N_18363,N_17553,N_17874);
or U18364 (N_18364,N_17694,N_17664);
and U18365 (N_18365,N_17719,N_17534);
xor U18366 (N_18366,N_17571,N_17989);
or U18367 (N_18367,N_17602,N_18021);
nor U18368 (N_18368,N_17819,N_18100);
or U18369 (N_18369,N_17623,N_18091);
nor U18370 (N_18370,N_17542,N_17688);
and U18371 (N_18371,N_17981,N_17505);
nand U18372 (N_18372,N_17549,N_17772);
nand U18373 (N_18373,N_17590,N_18103);
nand U18374 (N_18374,N_17778,N_17648);
nand U18375 (N_18375,N_18036,N_17579);
or U18376 (N_18376,N_17865,N_17960);
or U18377 (N_18377,N_17588,N_17616);
xnor U18378 (N_18378,N_17681,N_17862);
and U18379 (N_18379,N_18093,N_17711);
or U18380 (N_18380,N_17531,N_17774);
nor U18381 (N_18381,N_17974,N_18108);
nand U18382 (N_18382,N_17544,N_17801);
nand U18383 (N_18383,N_17547,N_18047);
xnor U18384 (N_18384,N_18096,N_17758);
and U18385 (N_18385,N_17795,N_17592);
xor U18386 (N_18386,N_18083,N_17514);
and U18387 (N_18387,N_18045,N_17972);
nor U18388 (N_18388,N_17667,N_17746);
and U18389 (N_18389,N_17985,N_17551);
nand U18390 (N_18390,N_17890,N_17849);
or U18391 (N_18391,N_17909,N_17920);
nor U18392 (N_18392,N_17966,N_17963);
nand U18393 (N_18393,N_17521,N_17564);
xor U18394 (N_18394,N_17987,N_17639);
xor U18395 (N_18395,N_17811,N_17535);
nand U18396 (N_18396,N_17504,N_17593);
nor U18397 (N_18397,N_17889,N_17604);
nand U18398 (N_18398,N_18123,N_17560);
nand U18399 (N_18399,N_17993,N_17813);
nor U18400 (N_18400,N_17844,N_17883);
xnor U18401 (N_18401,N_18113,N_18073);
nor U18402 (N_18402,N_17797,N_17815);
or U18403 (N_18403,N_18090,N_17912);
nand U18404 (N_18404,N_17657,N_17712);
or U18405 (N_18405,N_17587,N_17869);
nand U18406 (N_18406,N_18009,N_17659);
or U18407 (N_18407,N_17979,N_17539);
nor U18408 (N_18408,N_18124,N_17622);
and U18409 (N_18409,N_17777,N_18050);
nor U18410 (N_18410,N_17525,N_18116);
nand U18411 (N_18411,N_18072,N_18067);
nand U18412 (N_18412,N_17730,N_18005);
nor U18413 (N_18413,N_17721,N_17729);
nand U18414 (N_18414,N_17782,N_17830);
and U18415 (N_18415,N_17916,N_18087);
and U18416 (N_18416,N_17752,N_17775);
and U18417 (N_18417,N_17791,N_17692);
and U18418 (N_18418,N_18094,N_18001);
and U18419 (N_18419,N_18110,N_17753);
nand U18420 (N_18420,N_17969,N_17704);
and U18421 (N_18421,N_17864,N_17548);
and U18422 (N_18422,N_17640,N_17926);
or U18423 (N_18423,N_17835,N_18006);
or U18424 (N_18424,N_17944,N_17952);
and U18425 (N_18425,N_17671,N_18101);
nor U18426 (N_18426,N_17898,N_17783);
nor U18427 (N_18427,N_18004,N_17995);
or U18428 (N_18428,N_17676,N_17857);
xnor U18429 (N_18429,N_17683,N_17868);
nor U18430 (N_18430,N_17586,N_17851);
nand U18431 (N_18431,N_17655,N_18012);
and U18432 (N_18432,N_17617,N_17899);
or U18433 (N_18433,N_17845,N_17607);
nor U18434 (N_18434,N_17540,N_17854);
xor U18435 (N_18435,N_17703,N_18092);
or U18436 (N_18436,N_17673,N_17742);
nor U18437 (N_18437,N_17770,N_18122);
or U18438 (N_18438,N_17570,N_18097);
or U18439 (N_18439,N_17723,N_17571);
nand U18440 (N_18440,N_17546,N_17957);
nor U18441 (N_18441,N_17893,N_17785);
or U18442 (N_18442,N_17671,N_18110);
nor U18443 (N_18443,N_17854,N_17913);
nand U18444 (N_18444,N_17971,N_17814);
and U18445 (N_18445,N_17607,N_17990);
nor U18446 (N_18446,N_17885,N_17612);
and U18447 (N_18447,N_17963,N_17854);
nand U18448 (N_18448,N_17620,N_17583);
xor U18449 (N_18449,N_17547,N_17749);
nor U18450 (N_18450,N_17668,N_18026);
xor U18451 (N_18451,N_17880,N_17998);
nor U18452 (N_18452,N_18094,N_17863);
nand U18453 (N_18453,N_17916,N_17637);
xor U18454 (N_18454,N_17633,N_17810);
nand U18455 (N_18455,N_17955,N_17560);
nand U18456 (N_18456,N_17621,N_17835);
or U18457 (N_18457,N_17765,N_17709);
and U18458 (N_18458,N_17920,N_18115);
nor U18459 (N_18459,N_17627,N_17840);
xnor U18460 (N_18460,N_17650,N_17839);
xnor U18461 (N_18461,N_17953,N_17540);
xor U18462 (N_18462,N_17659,N_17733);
xnor U18463 (N_18463,N_18042,N_17598);
nand U18464 (N_18464,N_17740,N_18017);
nor U18465 (N_18465,N_18019,N_17604);
or U18466 (N_18466,N_17817,N_17780);
and U18467 (N_18467,N_17544,N_17907);
and U18468 (N_18468,N_18113,N_17653);
or U18469 (N_18469,N_18022,N_17944);
or U18470 (N_18470,N_17830,N_17640);
or U18471 (N_18471,N_17725,N_17683);
nand U18472 (N_18472,N_17598,N_17621);
nand U18473 (N_18473,N_17888,N_17663);
or U18474 (N_18474,N_17971,N_18123);
xor U18475 (N_18475,N_17505,N_17594);
nand U18476 (N_18476,N_17840,N_17928);
or U18477 (N_18477,N_17839,N_18019);
nand U18478 (N_18478,N_17928,N_17897);
and U18479 (N_18479,N_17765,N_17869);
xnor U18480 (N_18480,N_17622,N_18087);
nand U18481 (N_18481,N_17788,N_17508);
xnor U18482 (N_18482,N_17656,N_17872);
or U18483 (N_18483,N_18096,N_17909);
nor U18484 (N_18484,N_17643,N_18119);
and U18485 (N_18485,N_17813,N_17548);
or U18486 (N_18486,N_17787,N_18060);
nand U18487 (N_18487,N_17864,N_18079);
nor U18488 (N_18488,N_17671,N_17500);
xor U18489 (N_18489,N_17533,N_17954);
nand U18490 (N_18490,N_18000,N_17597);
xor U18491 (N_18491,N_18124,N_17704);
or U18492 (N_18492,N_17578,N_17862);
nand U18493 (N_18493,N_18005,N_17598);
xor U18494 (N_18494,N_17809,N_17950);
nor U18495 (N_18495,N_17740,N_18042);
xor U18496 (N_18496,N_17996,N_17732);
nand U18497 (N_18497,N_17889,N_18123);
or U18498 (N_18498,N_17967,N_18066);
nand U18499 (N_18499,N_17861,N_17648);
nand U18500 (N_18500,N_17797,N_17878);
nor U18501 (N_18501,N_17656,N_17628);
nor U18502 (N_18502,N_17563,N_17613);
and U18503 (N_18503,N_18068,N_17833);
or U18504 (N_18504,N_17572,N_17582);
and U18505 (N_18505,N_18031,N_17884);
xnor U18506 (N_18506,N_17520,N_17780);
nor U18507 (N_18507,N_17889,N_18111);
or U18508 (N_18508,N_17581,N_17619);
and U18509 (N_18509,N_17996,N_17871);
nor U18510 (N_18510,N_17530,N_18019);
and U18511 (N_18511,N_17751,N_17913);
xor U18512 (N_18512,N_18077,N_17945);
or U18513 (N_18513,N_17645,N_17896);
and U18514 (N_18514,N_18122,N_17729);
xnor U18515 (N_18515,N_17785,N_18113);
nand U18516 (N_18516,N_17889,N_17855);
xnor U18517 (N_18517,N_17846,N_17549);
nand U18518 (N_18518,N_17871,N_17975);
nor U18519 (N_18519,N_17521,N_18052);
xnor U18520 (N_18520,N_17701,N_18095);
xnor U18521 (N_18521,N_17761,N_17918);
xor U18522 (N_18522,N_18026,N_17897);
and U18523 (N_18523,N_18092,N_17949);
nand U18524 (N_18524,N_17692,N_17697);
nor U18525 (N_18525,N_17712,N_17590);
or U18526 (N_18526,N_17640,N_17869);
nor U18527 (N_18527,N_18044,N_17647);
xnor U18528 (N_18528,N_17913,N_17656);
and U18529 (N_18529,N_17775,N_18009);
and U18530 (N_18530,N_17619,N_17964);
xnor U18531 (N_18531,N_17820,N_17697);
nor U18532 (N_18532,N_17524,N_17942);
and U18533 (N_18533,N_18062,N_18034);
nor U18534 (N_18534,N_18054,N_18074);
xor U18535 (N_18535,N_17681,N_17502);
and U18536 (N_18536,N_17658,N_17828);
nand U18537 (N_18537,N_17583,N_17655);
and U18538 (N_18538,N_17837,N_17932);
nand U18539 (N_18539,N_17500,N_18069);
nand U18540 (N_18540,N_17934,N_17684);
nor U18541 (N_18541,N_17913,N_17621);
nor U18542 (N_18542,N_17622,N_17511);
nand U18543 (N_18543,N_18040,N_17990);
or U18544 (N_18544,N_17662,N_17594);
xnor U18545 (N_18545,N_17987,N_17703);
or U18546 (N_18546,N_17967,N_17665);
or U18547 (N_18547,N_17783,N_17507);
xnor U18548 (N_18548,N_17594,N_17937);
and U18549 (N_18549,N_17757,N_17840);
xnor U18550 (N_18550,N_17963,N_17814);
nor U18551 (N_18551,N_17855,N_18074);
xor U18552 (N_18552,N_17876,N_17829);
or U18553 (N_18553,N_17947,N_17910);
nor U18554 (N_18554,N_17862,N_17984);
nor U18555 (N_18555,N_17797,N_17604);
or U18556 (N_18556,N_17759,N_18047);
or U18557 (N_18557,N_18104,N_17874);
or U18558 (N_18558,N_17668,N_17838);
xor U18559 (N_18559,N_17850,N_17572);
and U18560 (N_18560,N_17559,N_17981);
or U18561 (N_18561,N_18121,N_17683);
xnor U18562 (N_18562,N_17862,N_17831);
and U18563 (N_18563,N_17628,N_17627);
and U18564 (N_18564,N_17932,N_17915);
nor U18565 (N_18565,N_18064,N_17687);
nand U18566 (N_18566,N_17941,N_17751);
nand U18567 (N_18567,N_17719,N_17715);
or U18568 (N_18568,N_17733,N_17740);
or U18569 (N_18569,N_17735,N_17900);
or U18570 (N_18570,N_18053,N_18001);
xnor U18571 (N_18571,N_17763,N_17826);
xor U18572 (N_18572,N_17960,N_18033);
xor U18573 (N_18573,N_18003,N_17799);
nor U18574 (N_18574,N_17945,N_18092);
nor U18575 (N_18575,N_17819,N_17776);
nand U18576 (N_18576,N_17845,N_17506);
nor U18577 (N_18577,N_17922,N_18024);
xor U18578 (N_18578,N_17553,N_17558);
and U18579 (N_18579,N_17866,N_17891);
and U18580 (N_18580,N_17863,N_17509);
or U18581 (N_18581,N_17643,N_17895);
xor U18582 (N_18582,N_17963,N_17987);
nand U18583 (N_18583,N_17590,N_17611);
and U18584 (N_18584,N_17561,N_17523);
xor U18585 (N_18585,N_17993,N_17554);
nand U18586 (N_18586,N_18037,N_17856);
xnor U18587 (N_18587,N_17765,N_17699);
or U18588 (N_18588,N_17547,N_17832);
nor U18589 (N_18589,N_18083,N_17621);
nor U18590 (N_18590,N_18048,N_17812);
nor U18591 (N_18591,N_18028,N_17686);
and U18592 (N_18592,N_17569,N_17506);
and U18593 (N_18593,N_17598,N_18068);
nand U18594 (N_18594,N_17940,N_18009);
and U18595 (N_18595,N_17673,N_17547);
nand U18596 (N_18596,N_17632,N_18088);
xor U18597 (N_18597,N_17781,N_18059);
or U18598 (N_18598,N_17780,N_18045);
nand U18599 (N_18599,N_17642,N_17693);
nand U18600 (N_18600,N_17976,N_17941);
nand U18601 (N_18601,N_17921,N_17666);
nand U18602 (N_18602,N_17953,N_17695);
nand U18603 (N_18603,N_18099,N_18029);
and U18604 (N_18604,N_17790,N_17591);
and U18605 (N_18605,N_17798,N_17616);
and U18606 (N_18606,N_17544,N_17596);
nor U18607 (N_18607,N_17809,N_17840);
and U18608 (N_18608,N_17959,N_17966);
nand U18609 (N_18609,N_17743,N_18105);
xnor U18610 (N_18610,N_17709,N_17652);
nor U18611 (N_18611,N_17789,N_17933);
and U18612 (N_18612,N_17913,N_17800);
nor U18613 (N_18613,N_17664,N_18073);
or U18614 (N_18614,N_17802,N_17931);
or U18615 (N_18615,N_17983,N_17650);
nand U18616 (N_18616,N_17844,N_18084);
or U18617 (N_18617,N_17971,N_17994);
nor U18618 (N_18618,N_17620,N_18020);
xnor U18619 (N_18619,N_17901,N_17842);
nand U18620 (N_18620,N_17952,N_17576);
xor U18621 (N_18621,N_17748,N_17910);
or U18622 (N_18622,N_18059,N_17645);
xnor U18623 (N_18623,N_17770,N_17562);
nor U18624 (N_18624,N_17602,N_17758);
nor U18625 (N_18625,N_17828,N_17957);
xnor U18626 (N_18626,N_17585,N_17717);
and U18627 (N_18627,N_17921,N_17934);
or U18628 (N_18628,N_17664,N_17848);
and U18629 (N_18629,N_17651,N_17865);
or U18630 (N_18630,N_17839,N_17797);
and U18631 (N_18631,N_17830,N_18068);
or U18632 (N_18632,N_18102,N_17700);
or U18633 (N_18633,N_17685,N_17665);
xor U18634 (N_18634,N_17845,N_17985);
and U18635 (N_18635,N_18023,N_17845);
xnor U18636 (N_18636,N_17642,N_17767);
and U18637 (N_18637,N_18016,N_17915);
nand U18638 (N_18638,N_17579,N_17512);
or U18639 (N_18639,N_17975,N_17915);
or U18640 (N_18640,N_17926,N_17838);
nor U18641 (N_18641,N_17867,N_17922);
and U18642 (N_18642,N_18064,N_17739);
nand U18643 (N_18643,N_17789,N_17519);
xor U18644 (N_18644,N_17976,N_17741);
xnor U18645 (N_18645,N_17838,N_18077);
nand U18646 (N_18646,N_17501,N_17587);
nor U18647 (N_18647,N_18091,N_17689);
nand U18648 (N_18648,N_17640,N_17836);
nor U18649 (N_18649,N_17617,N_18060);
nand U18650 (N_18650,N_18025,N_17761);
and U18651 (N_18651,N_17947,N_17908);
nand U18652 (N_18652,N_18113,N_17721);
or U18653 (N_18653,N_17649,N_17632);
nand U18654 (N_18654,N_17706,N_17595);
or U18655 (N_18655,N_17731,N_17975);
or U18656 (N_18656,N_17831,N_17856);
or U18657 (N_18657,N_18007,N_17933);
nand U18658 (N_18658,N_17992,N_17539);
xnor U18659 (N_18659,N_17779,N_17540);
nand U18660 (N_18660,N_17613,N_17797);
or U18661 (N_18661,N_17891,N_17992);
and U18662 (N_18662,N_17583,N_17953);
and U18663 (N_18663,N_18076,N_17967);
and U18664 (N_18664,N_17992,N_17803);
nand U18665 (N_18665,N_17574,N_17547);
or U18666 (N_18666,N_18124,N_18112);
and U18667 (N_18667,N_17576,N_17893);
nor U18668 (N_18668,N_17636,N_17980);
nand U18669 (N_18669,N_17958,N_18055);
xnor U18670 (N_18670,N_18086,N_18087);
nand U18671 (N_18671,N_18064,N_17879);
xor U18672 (N_18672,N_18119,N_17886);
nor U18673 (N_18673,N_17653,N_17803);
xnor U18674 (N_18674,N_18052,N_17913);
nand U18675 (N_18675,N_17553,N_17892);
xnor U18676 (N_18676,N_17827,N_17650);
nor U18677 (N_18677,N_17901,N_17880);
nand U18678 (N_18678,N_17948,N_17789);
nand U18679 (N_18679,N_17743,N_18031);
or U18680 (N_18680,N_17918,N_17851);
nor U18681 (N_18681,N_17753,N_17931);
nor U18682 (N_18682,N_17650,N_17752);
nor U18683 (N_18683,N_17780,N_17939);
or U18684 (N_18684,N_17749,N_18108);
nand U18685 (N_18685,N_17680,N_17583);
or U18686 (N_18686,N_17819,N_18096);
xor U18687 (N_18687,N_17994,N_17884);
and U18688 (N_18688,N_17523,N_17788);
and U18689 (N_18689,N_18067,N_17720);
nor U18690 (N_18690,N_17703,N_17701);
xor U18691 (N_18691,N_17725,N_17958);
or U18692 (N_18692,N_17546,N_17708);
or U18693 (N_18693,N_17958,N_17667);
xor U18694 (N_18694,N_17527,N_17775);
xnor U18695 (N_18695,N_17854,N_17896);
nor U18696 (N_18696,N_17883,N_17884);
xnor U18697 (N_18697,N_17802,N_18001);
nor U18698 (N_18698,N_17873,N_17714);
or U18699 (N_18699,N_17895,N_17979);
or U18700 (N_18700,N_18056,N_17947);
nand U18701 (N_18701,N_17514,N_17832);
or U18702 (N_18702,N_18092,N_18048);
nand U18703 (N_18703,N_18013,N_17894);
and U18704 (N_18704,N_17772,N_17900);
and U18705 (N_18705,N_17557,N_17834);
nor U18706 (N_18706,N_17604,N_17531);
xnor U18707 (N_18707,N_17875,N_17735);
or U18708 (N_18708,N_17830,N_17927);
or U18709 (N_18709,N_18115,N_17657);
nor U18710 (N_18710,N_17544,N_17763);
or U18711 (N_18711,N_17605,N_18111);
and U18712 (N_18712,N_17527,N_18057);
or U18713 (N_18713,N_17628,N_17977);
nand U18714 (N_18714,N_18047,N_17866);
and U18715 (N_18715,N_18006,N_17577);
and U18716 (N_18716,N_17524,N_17972);
nand U18717 (N_18717,N_17603,N_18014);
nor U18718 (N_18718,N_17968,N_17646);
nor U18719 (N_18719,N_17635,N_17983);
nand U18720 (N_18720,N_17941,N_18034);
or U18721 (N_18721,N_18071,N_17718);
xnor U18722 (N_18722,N_17625,N_17981);
or U18723 (N_18723,N_17869,N_18006);
or U18724 (N_18724,N_18044,N_17874);
xor U18725 (N_18725,N_17524,N_17985);
and U18726 (N_18726,N_17983,N_17737);
xor U18727 (N_18727,N_17990,N_17592);
nand U18728 (N_18728,N_17686,N_17613);
and U18729 (N_18729,N_17878,N_17771);
or U18730 (N_18730,N_17802,N_17538);
nand U18731 (N_18731,N_17812,N_17887);
or U18732 (N_18732,N_17985,N_17878);
or U18733 (N_18733,N_17912,N_18030);
nor U18734 (N_18734,N_17911,N_18040);
or U18735 (N_18735,N_17879,N_17630);
nor U18736 (N_18736,N_17525,N_17836);
xnor U18737 (N_18737,N_17615,N_18108);
nor U18738 (N_18738,N_17705,N_17756);
or U18739 (N_18739,N_17879,N_18114);
or U18740 (N_18740,N_17780,N_17504);
and U18741 (N_18741,N_17616,N_17550);
or U18742 (N_18742,N_18047,N_17781);
xor U18743 (N_18743,N_18119,N_18025);
and U18744 (N_18744,N_17986,N_17764);
and U18745 (N_18745,N_17687,N_17908);
xor U18746 (N_18746,N_18024,N_18102);
nor U18747 (N_18747,N_18068,N_17872);
xor U18748 (N_18748,N_17958,N_17895);
nor U18749 (N_18749,N_17962,N_17876);
or U18750 (N_18750,N_18463,N_18459);
and U18751 (N_18751,N_18294,N_18267);
and U18752 (N_18752,N_18297,N_18602);
and U18753 (N_18753,N_18533,N_18171);
and U18754 (N_18754,N_18206,N_18411);
and U18755 (N_18755,N_18486,N_18214);
xnor U18756 (N_18756,N_18188,N_18429);
nor U18757 (N_18757,N_18296,N_18230);
xor U18758 (N_18758,N_18657,N_18387);
nor U18759 (N_18759,N_18271,N_18458);
nand U18760 (N_18760,N_18719,N_18205);
and U18761 (N_18761,N_18419,N_18558);
or U18762 (N_18762,N_18652,N_18312);
and U18763 (N_18763,N_18606,N_18338);
xnor U18764 (N_18764,N_18432,N_18410);
nor U18765 (N_18765,N_18450,N_18368);
and U18766 (N_18766,N_18344,N_18495);
nor U18767 (N_18767,N_18726,N_18663);
or U18768 (N_18768,N_18137,N_18731);
xnor U18769 (N_18769,N_18521,N_18646);
xor U18770 (N_18770,N_18715,N_18626);
or U18771 (N_18771,N_18132,N_18594);
and U18772 (N_18772,N_18467,N_18499);
xnor U18773 (N_18773,N_18728,N_18209);
xor U18774 (N_18774,N_18423,N_18538);
nor U18775 (N_18775,N_18156,N_18404);
xnor U18776 (N_18776,N_18660,N_18196);
and U18777 (N_18777,N_18211,N_18185);
xnor U18778 (N_18778,N_18367,N_18142);
xnor U18779 (N_18779,N_18697,N_18397);
or U18780 (N_18780,N_18222,N_18690);
nor U18781 (N_18781,N_18330,N_18381);
or U18782 (N_18782,N_18317,N_18568);
nand U18783 (N_18783,N_18565,N_18596);
or U18784 (N_18784,N_18694,N_18143);
xnor U18785 (N_18785,N_18258,N_18454);
nor U18786 (N_18786,N_18168,N_18549);
nor U18787 (N_18787,N_18709,N_18203);
xnor U18788 (N_18788,N_18527,N_18712);
and U18789 (N_18789,N_18217,N_18255);
or U18790 (N_18790,N_18377,N_18581);
xnor U18791 (N_18791,N_18640,N_18334);
or U18792 (N_18792,N_18193,N_18714);
or U18793 (N_18793,N_18266,N_18451);
or U18794 (N_18794,N_18460,N_18508);
nor U18795 (N_18795,N_18559,N_18433);
nor U18796 (N_18796,N_18474,N_18325);
xor U18797 (N_18797,N_18625,N_18311);
xnor U18798 (N_18798,N_18286,N_18413);
and U18799 (N_18799,N_18337,N_18277);
or U18800 (N_18800,N_18611,N_18219);
nor U18801 (N_18801,N_18524,N_18208);
nor U18802 (N_18802,N_18420,N_18724);
and U18803 (N_18803,N_18250,N_18529);
xnor U18804 (N_18804,N_18424,N_18456);
nand U18805 (N_18805,N_18160,N_18479);
and U18806 (N_18806,N_18354,N_18335);
and U18807 (N_18807,N_18446,N_18287);
or U18808 (N_18808,N_18157,N_18293);
nor U18809 (N_18809,N_18617,N_18200);
nand U18810 (N_18810,N_18722,N_18585);
and U18811 (N_18811,N_18707,N_18537);
nand U18812 (N_18812,N_18621,N_18434);
nand U18813 (N_18813,N_18542,N_18484);
and U18814 (N_18814,N_18682,N_18135);
nor U18815 (N_18815,N_18476,N_18572);
or U18816 (N_18816,N_18318,N_18610);
nor U18817 (N_18817,N_18609,N_18139);
nand U18818 (N_18818,N_18373,N_18147);
or U18819 (N_18819,N_18361,N_18667);
xor U18820 (N_18820,N_18738,N_18349);
and U18821 (N_18821,N_18741,N_18642);
and U18822 (N_18822,N_18195,N_18341);
and U18823 (N_18823,N_18322,N_18548);
xnor U18824 (N_18824,N_18336,N_18645);
or U18825 (N_18825,N_18704,N_18408);
nand U18826 (N_18826,N_18540,N_18298);
and U18827 (N_18827,N_18723,N_18145);
xnor U18828 (N_18828,N_18278,N_18234);
nor U18829 (N_18829,N_18551,N_18409);
and U18830 (N_18830,N_18616,N_18695);
nand U18831 (N_18831,N_18422,N_18439);
and U18832 (N_18832,N_18735,N_18496);
or U18833 (N_18833,N_18184,N_18612);
nand U18834 (N_18834,N_18315,N_18442);
nor U18835 (N_18835,N_18369,N_18281);
nand U18836 (N_18836,N_18687,N_18473);
xnor U18837 (N_18837,N_18681,N_18493);
or U18838 (N_18838,N_18632,N_18162);
nand U18839 (N_18839,N_18482,N_18194);
nand U18840 (N_18840,N_18169,N_18659);
and U18841 (N_18841,N_18586,N_18597);
nor U18842 (N_18842,N_18375,N_18212);
nor U18843 (N_18843,N_18165,N_18290);
or U18844 (N_18844,N_18563,N_18418);
nand U18845 (N_18845,N_18522,N_18417);
nor U18846 (N_18846,N_18327,N_18405);
xnor U18847 (N_18847,N_18589,N_18452);
and U18848 (N_18848,N_18173,N_18428);
or U18849 (N_18849,N_18183,N_18300);
xnor U18850 (N_18850,N_18187,N_18591);
xnor U18851 (N_18851,N_18430,N_18272);
nand U18852 (N_18852,N_18498,N_18393);
nand U18853 (N_18853,N_18357,N_18435);
nand U18854 (N_18854,N_18680,N_18636);
xnor U18855 (N_18855,N_18264,N_18649);
nor U18856 (N_18856,N_18265,N_18643);
xnor U18857 (N_18857,N_18233,N_18555);
and U18858 (N_18858,N_18530,N_18191);
or U18859 (N_18859,N_18363,N_18678);
xnor U18860 (N_18860,N_18566,N_18666);
nor U18861 (N_18861,N_18746,N_18416);
xnor U18862 (N_18862,N_18438,N_18148);
nand U18863 (N_18863,N_18398,N_18468);
nand U18864 (N_18864,N_18273,N_18362);
nor U18865 (N_18865,N_18204,N_18425);
nand U18866 (N_18866,N_18466,N_18261);
or U18867 (N_18867,N_18729,N_18154);
or U18868 (N_18868,N_18257,N_18447);
nor U18869 (N_18869,N_18130,N_18231);
nor U18870 (N_18870,N_18440,N_18494);
and U18871 (N_18871,N_18742,N_18736);
nor U18872 (N_18872,N_18518,N_18703);
or U18873 (N_18873,N_18553,N_18243);
nor U18874 (N_18874,N_18492,N_18622);
and U18875 (N_18875,N_18749,N_18370);
nand U18876 (N_18876,N_18406,N_18569);
xor U18877 (N_18877,N_18544,N_18613);
and U18878 (N_18878,N_18331,N_18730);
or U18879 (N_18879,N_18477,N_18615);
xor U18880 (N_18880,N_18587,N_18455);
or U18881 (N_18881,N_18737,N_18633);
nand U18882 (N_18882,N_18342,N_18166);
xor U18883 (N_18883,N_18202,N_18299);
nor U18884 (N_18884,N_18592,N_18603);
nand U18885 (N_18885,N_18270,N_18326);
nand U18886 (N_18886,N_18391,N_18229);
and U18887 (N_18887,N_18465,N_18235);
or U18888 (N_18888,N_18283,N_18339);
nand U18889 (N_18889,N_18532,N_18745);
nor U18890 (N_18890,N_18483,N_18675);
nand U18891 (N_18891,N_18249,N_18668);
or U18892 (N_18892,N_18576,N_18547);
xnor U18893 (N_18893,N_18153,N_18520);
or U18894 (N_18894,N_18348,N_18708);
xor U18895 (N_18895,N_18535,N_18321);
nor U18896 (N_18896,N_18172,N_18316);
nand U18897 (N_18897,N_18443,N_18323);
nand U18898 (N_18898,N_18351,N_18329);
nor U18899 (N_18899,N_18614,N_18671);
or U18900 (N_18900,N_18526,N_18554);
and U18901 (N_18901,N_18181,N_18138);
nand U18902 (N_18902,N_18517,N_18259);
xnor U18903 (N_18903,N_18140,N_18502);
xor U18904 (N_18904,N_18689,N_18644);
xnor U18905 (N_18905,N_18155,N_18634);
or U18906 (N_18906,N_18346,N_18402);
or U18907 (N_18907,N_18670,N_18599);
nand U18908 (N_18908,N_18485,N_18292);
and U18909 (N_18909,N_18504,N_18464);
nor U18910 (N_18910,N_18178,N_18552);
or U18911 (N_18911,N_18304,N_18305);
and U18912 (N_18912,N_18125,N_18262);
nand U18913 (N_18913,N_18503,N_18141);
nor U18914 (N_18914,N_18706,N_18475);
nor U18915 (N_18915,N_18340,N_18618);
nor U18916 (N_18916,N_18276,N_18225);
or U18917 (N_18917,N_18511,N_18491);
xor U18918 (N_18918,N_18515,N_18574);
nand U18919 (N_18919,N_18620,N_18371);
or U18920 (N_18920,N_18389,N_18638);
xor U18921 (N_18921,N_18177,N_18306);
xnor U18922 (N_18922,N_18658,N_18543);
and U18923 (N_18923,N_18151,N_18175);
xor U18924 (N_18924,N_18573,N_18718);
nand U18925 (N_18925,N_18131,N_18673);
nor U18926 (N_18926,N_18421,N_18500);
and U18927 (N_18927,N_18747,N_18698);
nand U18928 (N_18928,N_18725,N_18583);
or U18929 (N_18929,N_18386,N_18244);
or U18930 (N_18930,N_18268,N_18720);
and U18931 (N_18931,N_18541,N_18732);
nor U18932 (N_18932,N_18415,N_18358);
nor U18933 (N_18933,N_18693,N_18469);
nor U18934 (N_18934,N_18164,N_18174);
or U18935 (N_18935,N_18711,N_18134);
or U18936 (N_18936,N_18545,N_18279);
nand U18937 (N_18937,N_18282,N_18702);
and U18938 (N_18938,N_18701,N_18528);
or U18939 (N_18939,N_18669,N_18700);
nor U18940 (N_18940,N_18685,N_18241);
nand U18941 (N_18941,N_18383,N_18260);
xnor U18942 (N_18942,N_18601,N_18256);
and U18943 (N_18943,N_18355,N_18733);
or U18944 (N_18944,N_18637,N_18691);
or U18945 (N_18945,N_18710,N_18328);
xnor U18946 (N_18946,N_18240,N_18320);
nor U18947 (N_18947,N_18656,N_18744);
and U18948 (N_18948,N_18186,N_18376);
xnor U18949 (N_18949,N_18679,N_18713);
nand U18950 (N_18950,N_18721,N_18239);
xnor U18951 (N_18951,N_18575,N_18523);
nand U18952 (N_18952,N_18630,N_18384);
nor U18953 (N_18953,N_18136,N_18197);
nand U18954 (N_18954,N_18407,N_18253);
xor U18955 (N_18955,N_18692,N_18146);
and U18956 (N_18956,N_18686,N_18133);
nand U18957 (N_18957,N_18561,N_18490);
xor U18958 (N_18958,N_18635,N_18359);
nor U18959 (N_18959,N_18269,N_18683);
nand U18960 (N_18960,N_18248,N_18274);
xor U18961 (N_18961,N_18623,N_18309);
and U18962 (N_18962,N_18457,N_18441);
nand U18963 (N_18963,N_18661,N_18489);
nor U18964 (N_18964,N_18696,N_18647);
xnor U18965 (N_18965,N_18727,N_18513);
or U18966 (N_18966,N_18471,N_18608);
and U18967 (N_18967,N_18598,N_18578);
and U18968 (N_18968,N_18674,N_18705);
nor U18969 (N_18969,N_18449,N_18295);
and U18970 (N_18970,N_18159,N_18629);
xor U18971 (N_18971,N_18519,N_18288);
xor U18972 (N_18972,N_18247,N_18487);
nand U18973 (N_18973,N_18396,N_18444);
nor U18974 (N_18974,N_18560,N_18382);
nand U18975 (N_18975,N_18158,N_18388);
nand U18976 (N_18976,N_18639,N_18472);
nor U18977 (N_18977,N_18365,N_18672);
nor U18978 (N_18978,N_18514,N_18333);
nand U18979 (N_18979,N_18478,N_18161);
nand U18980 (N_18980,N_18564,N_18650);
xnor U18981 (N_18981,N_18403,N_18289);
xnor U18982 (N_18982,N_18182,N_18536);
and U18983 (N_18983,N_18717,N_18462);
nand U18984 (N_18984,N_18607,N_18655);
or U18985 (N_18985,N_18374,N_18648);
or U18986 (N_18986,N_18412,N_18176);
and U18987 (N_18987,N_18347,N_18242);
or U18988 (N_18988,N_18284,N_18167);
nand U18989 (N_18989,N_18525,N_18604);
or U18990 (N_18990,N_18512,N_18127);
and U18991 (N_18991,N_18509,N_18236);
or U18992 (N_18992,N_18343,N_18199);
xnor U18993 (N_18993,N_18345,N_18567);
or U18994 (N_18994,N_18350,N_18470);
or U18995 (N_18995,N_18220,N_18189);
nand U18996 (N_18996,N_18232,N_18152);
xnor U18997 (N_18997,N_18590,N_18307);
or U18998 (N_18998,N_18605,N_18356);
and U18999 (N_18999,N_18314,N_18228);
nor U19000 (N_19000,N_18180,N_18400);
nor U19001 (N_19001,N_18739,N_18263);
nand U19002 (N_19002,N_18352,N_18399);
or U19003 (N_19003,N_18332,N_18431);
or U19004 (N_19004,N_18394,N_18252);
nand U19005 (N_19005,N_18207,N_18748);
and U19006 (N_19006,N_18510,N_18372);
nor U19007 (N_19007,N_18595,N_18251);
nand U19008 (N_19008,N_18302,N_18366);
and U19009 (N_19009,N_18481,N_18224);
and U19010 (N_19010,N_18353,N_18128);
nand U19011 (N_19011,N_18392,N_18505);
and U19012 (N_19012,N_18593,N_18577);
xor U19013 (N_19013,N_18201,N_18740);
nor U19014 (N_19014,N_18324,N_18488);
nand U19015 (N_19015,N_18507,N_18743);
xor U19016 (N_19016,N_18582,N_18624);
or U19017 (N_19017,N_18215,N_18301);
nand U19018 (N_19018,N_18557,N_18437);
nand U19019 (N_19019,N_18600,N_18227);
xnor U19020 (N_19020,N_18380,N_18144);
and U19021 (N_19021,N_18534,N_18226);
nand U19022 (N_19022,N_18414,N_18190);
or U19023 (N_19023,N_18150,N_18651);
nor U19024 (N_19024,N_18163,N_18285);
nand U19025 (N_19025,N_18641,N_18308);
nand U19026 (N_19026,N_18291,N_18379);
and U19027 (N_19027,N_18631,N_18676);
or U19028 (N_19028,N_18303,N_18313);
xor U19029 (N_19029,N_18584,N_18360);
and U19030 (N_19030,N_18436,N_18480);
and U19031 (N_19031,N_18516,N_18179);
nand U19032 (N_19032,N_18531,N_18506);
or U19033 (N_19033,N_18218,N_18385);
nand U19034 (N_19034,N_18654,N_18129);
and U19035 (N_19035,N_18310,N_18223);
xnor U19036 (N_19036,N_18580,N_18588);
xnor U19037 (N_19037,N_18254,N_18395);
or U19038 (N_19038,N_18628,N_18448);
nor U19039 (N_19039,N_18237,N_18539);
nor U19040 (N_19040,N_18501,N_18497);
and U19041 (N_19041,N_18149,N_18550);
xor U19042 (N_19042,N_18245,N_18378);
nand U19043 (N_19043,N_18546,N_18579);
nand U19044 (N_19044,N_18126,N_18390);
xnor U19045 (N_19045,N_18556,N_18664);
xnor U19046 (N_19046,N_18619,N_18662);
and U19047 (N_19047,N_18213,N_18453);
and U19048 (N_19048,N_18562,N_18570);
or U19049 (N_19049,N_18216,N_18699);
or U19050 (N_19050,N_18677,N_18734);
xor U19051 (N_19051,N_18627,N_18170);
and U19052 (N_19052,N_18364,N_18716);
nor U19053 (N_19053,N_18445,N_18238);
xnor U19054 (N_19054,N_18280,N_18684);
nor U19055 (N_19055,N_18653,N_18319);
nand U19056 (N_19056,N_18275,N_18461);
or U19057 (N_19057,N_18192,N_18210);
xor U19058 (N_19058,N_18198,N_18427);
or U19059 (N_19059,N_18688,N_18571);
or U19060 (N_19060,N_18665,N_18401);
or U19061 (N_19061,N_18221,N_18246);
nor U19062 (N_19062,N_18426,N_18631);
xnor U19063 (N_19063,N_18408,N_18736);
nand U19064 (N_19064,N_18290,N_18709);
nand U19065 (N_19065,N_18680,N_18612);
nand U19066 (N_19066,N_18607,N_18589);
xnor U19067 (N_19067,N_18719,N_18401);
nand U19068 (N_19068,N_18685,N_18199);
and U19069 (N_19069,N_18279,N_18723);
and U19070 (N_19070,N_18274,N_18140);
nor U19071 (N_19071,N_18175,N_18350);
xnor U19072 (N_19072,N_18516,N_18608);
nor U19073 (N_19073,N_18693,N_18560);
and U19074 (N_19074,N_18503,N_18427);
and U19075 (N_19075,N_18157,N_18447);
xnor U19076 (N_19076,N_18336,N_18383);
nand U19077 (N_19077,N_18166,N_18726);
nor U19078 (N_19078,N_18664,N_18475);
or U19079 (N_19079,N_18286,N_18328);
and U19080 (N_19080,N_18649,N_18580);
xor U19081 (N_19081,N_18642,N_18510);
or U19082 (N_19082,N_18652,N_18537);
nand U19083 (N_19083,N_18145,N_18604);
or U19084 (N_19084,N_18253,N_18443);
or U19085 (N_19085,N_18302,N_18360);
and U19086 (N_19086,N_18310,N_18451);
and U19087 (N_19087,N_18637,N_18509);
nor U19088 (N_19088,N_18194,N_18236);
and U19089 (N_19089,N_18345,N_18277);
or U19090 (N_19090,N_18265,N_18168);
or U19091 (N_19091,N_18722,N_18592);
nor U19092 (N_19092,N_18303,N_18133);
or U19093 (N_19093,N_18181,N_18639);
or U19094 (N_19094,N_18193,N_18598);
nand U19095 (N_19095,N_18510,N_18268);
nand U19096 (N_19096,N_18337,N_18210);
nor U19097 (N_19097,N_18508,N_18345);
nand U19098 (N_19098,N_18472,N_18431);
nand U19099 (N_19099,N_18263,N_18611);
or U19100 (N_19100,N_18410,N_18208);
xnor U19101 (N_19101,N_18640,N_18208);
nand U19102 (N_19102,N_18608,N_18566);
nand U19103 (N_19103,N_18568,N_18550);
or U19104 (N_19104,N_18151,N_18447);
or U19105 (N_19105,N_18447,N_18540);
xor U19106 (N_19106,N_18254,N_18732);
or U19107 (N_19107,N_18443,N_18246);
or U19108 (N_19108,N_18441,N_18315);
or U19109 (N_19109,N_18361,N_18592);
nor U19110 (N_19110,N_18259,N_18279);
xnor U19111 (N_19111,N_18598,N_18601);
or U19112 (N_19112,N_18375,N_18522);
or U19113 (N_19113,N_18412,N_18346);
xnor U19114 (N_19114,N_18154,N_18479);
and U19115 (N_19115,N_18297,N_18591);
nor U19116 (N_19116,N_18536,N_18717);
or U19117 (N_19117,N_18671,N_18709);
nand U19118 (N_19118,N_18563,N_18665);
nor U19119 (N_19119,N_18247,N_18161);
xnor U19120 (N_19120,N_18396,N_18745);
xor U19121 (N_19121,N_18445,N_18314);
and U19122 (N_19122,N_18614,N_18374);
xnor U19123 (N_19123,N_18437,N_18652);
and U19124 (N_19124,N_18454,N_18477);
and U19125 (N_19125,N_18698,N_18460);
nand U19126 (N_19126,N_18711,N_18228);
or U19127 (N_19127,N_18134,N_18513);
or U19128 (N_19128,N_18574,N_18203);
or U19129 (N_19129,N_18430,N_18426);
nor U19130 (N_19130,N_18470,N_18339);
nand U19131 (N_19131,N_18450,N_18165);
xnor U19132 (N_19132,N_18386,N_18639);
nor U19133 (N_19133,N_18255,N_18717);
xor U19134 (N_19134,N_18549,N_18695);
or U19135 (N_19135,N_18629,N_18509);
nor U19136 (N_19136,N_18458,N_18494);
xor U19137 (N_19137,N_18625,N_18207);
nand U19138 (N_19138,N_18715,N_18718);
or U19139 (N_19139,N_18404,N_18561);
or U19140 (N_19140,N_18638,N_18199);
nand U19141 (N_19141,N_18162,N_18595);
nand U19142 (N_19142,N_18453,N_18547);
nand U19143 (N_19143,N_18575,N_18196);
nor U19144 (N_19144,N_18561,N_18192);
and U19145 (N_19145,N_18299,N_18562);
or U19146 (N_19146,N_18300,N_18438);
nand U19147 (N_19147,N_18240,N_18350);
xor U19148 (N_19148,N_18369,N_18246);
or U19149 (N_19149,N_18271,N_18616);
nand U19150 (N_19150,N_18172,N_18590);
xor U19151 (N_19151,N_18665,N_18323);
or U19152 (N_19152,N_18211,N_18182);
nor U19153 (N_19153,N_18440,N_18253);
and U19154 (N_19154,N_18306,N_18372);
and U19155 (N_19155,N_18735,N_18420);
and U19156 (N_19156,N_18229,N_18176);
nor U19157 (N_19157,N_18232,N_18658);
xnor U19158 (N_19158,N_18604,N_18340);
xor U19159 (N_19159,N_18286,N_18412);
or U19160 (N_19160,N_18454,N_18585);
or U19161 (N_19161,N_18271,N_18363);
nor U19162 (N_19162,N_18206,N_18139);
or U19163 (N_19163,N_18698,N_18694);
nand U19164 (N_19164,N_18451,N_18676);
nand U19165 (N_19165,N_18272,N_18424);
xor U19166 (N_19166,N_18282,N_18474);
and U19167 (N_19167,N_18285,N_18435);
nand U19168 (N_19168,N_18423,N_18330);
nor U19169 (N_19169,N_18594,N_18643);
nor U19170 (N_19170,N_18536,N_18430);
and U19171 (N_19171,N_18504,N_18377);
nand U19172 (N_19172,N_18587,N_18362);
or U19173 (N_19173,N_18260,N_18268);
or U19174 (N_19174,N_18474,N_18442);
and U19175 (N_19175,N_18466,N_18293);
nor U19176 (N_19176,N_18325,N_18612);
xor U19177 (N_19177,N_18402,N_18707);
or U19178 (N_19178,N_18487,N_18211);
and U19179 (N_19179,N_18483,N_18663);
or U19180 (N_19180,N_18411,N_18143);
nor U19181 (N_19181,N_18464,N_18312);
nor U19182 (N_19182,N_18264,N_18141);
and U19183 (N_19183,N_18226,N_18680);
or U19184 (N_19184,N_18182,N_18399);
xor U19185 (N_19185,N_18194,N_18715);
xnor U19186 (N_19186,N_18545,N_18374);
nor U19187 (N_19187,N_18470,N_18216);
nand U19188 (N_19188,N_18502,N_18421);
or U19189 (N_19189,N_18231,N_18673);
or U19190 (N_19190,N_18432,N_18344);
xor U19191 (N_19191,N_18701,N_18613);
nand U19192 (N_19192,N_18497,N_18270);
or U19193 (N_19193,N_18527,N_18742);
nor U19194 (N_19194,N_18355,N_18519);
xnor U19195 (N_19195,N_18257,N_18406);
xnor U19196 (N_19196,N_18570,N_18165);
nor U19197 (N_19197,N_18718,N_18393);
xnor U19198 (N_19198,N_18466,N_18528);
or U19199 (N_19199,N_18734,N_18499);
and U19200 (N_19200,N_18225,N_18350);
and U19201 (N_19201,N_18195,N_18233);
or U19202 (N_19202,N_18679,N_18600);
and U19203 (N_19203,N_18199,N_18185);
xor U19204 (N_19204,N_18264,N_18535);
xor U19205 (N_19205,N_18317,N_18708);
or U19206 (N_19206,N_18374,N_18233);
nor U19207 (N_19207,N_18580,N_18560);
or U19208 (N_19208,N_18355,N_18326);
nor U19209 (N_19209,N_18541,N_18564);
nand U19210 (N_19210,N_18500,N_18221);
and U19211 (N_19211,N_18456,N_18406);
or U19212 (N_19212,N_18629,N_18590);
nor U19213 (N_19213,N_18483,N_18422);
nor U19214 (N_19214,N_18300,N_18678);
nor U19215 (N_19215,N_18401,N_18227);
and U19216 (N_19216,N_18554,N_18396);
nand U19217 (N_19217,N_18276,N_18317);
xnor U19218 (N_19218,N_18554,N_18571);
xnor U19219 (N_19219,N_18469,N_18316);
xnor U19220 (N_19220,N_18677,N_18571);
nand U19221 (N_19221,N_18155,N_18571);
xnor U19222 (N_19222,N_18634,N_18546);
nand U19223 (N_19223,N_18256,N_18554);
nor U19224 (N_19224,N_18163,N_18262);
nor U19225 (N_19225,N_18490,N_18269);
xor U19226 (N_19226,N_18154,N_18146);
nor U19227 (N_19227,N_18171,N_18133);
xnor U19228 (N_19228,N_18736,N_18542);
nor U19229 (N_19229,N_18273,N_18384);
xor U19230 (N_19230,N_18467,N_18732);
and U19231 (N_19231,N_18695,N_18151);
nor U19232 (N_19232,N_18228,N_18743);
nand U19233 (N_19233,N_18551,N_18554);
xor U19234 (N_19234,N_18476,N_18632);
and U19235 (N_19235,N_18256,N_18723);
nor U19236 (N_19236,N_18459,N_18138);
nor U19237 (N_19237,N_18620,N_18706);
nand U19238 (N_19238,N_18339,N_18668);
or U19239 (N_19239,N_18562,N_18542);
and U19240 (N_19240,N_18672,N_18610);
or U19241 (N_19241,N_18737,N_18653);
and U19242 (N_19242,N_18597,N_18698);
or U19243 (N_19243,N_18595,N_18692);
xor U19244 (N_19244,N_18706,N_18177);
xnor U19245 (N_19245,N_18170,N_18485);
nand U19246 (N_19246,N_18732,N_18488);
nor U19247 (N_19247,N_18657,N_18267);
nor U19248 (N_19248,N_18745,N_18630);
nor U19249 (N_19249,N_18300,N_18593);
nor U19250 (N_19250,N_18356,N_18674);
xnor U19251 (N_19251,N_18283,N_18194);
and U19252 (N_19252,N_18663,N_18582);
xnor U19253 (N_19253,N_18700,N_18336);
and U19254 (N_19254,N_18323,N_18605);
or U19255 (N_19255,N_18639,N_18152);
xor U19256 (N_19256,N_18509,N_18660);
xnor U19257 (N_19257,N_18580,N_18245);
and U19258 (N_19258,N_18581,N_18156);
nand U19259 (N_19259,N_18473,N_18409);
xor U19260 (N_19260,N_18432,N_18640);
nand U19261 (N_19261,N_18504,N_18311);
nand U19262 (N_19262,N_18163,N_18324);
xor U19263 (N_19263,N_18548,N_18160);
and U19264 (N_19264,N_18219,N_18413);
or U19265 (N_19265,N_18196,N_18420);
xnor U19266 (N_19266,N_18624,N_18438);
xor U19267 (N_19267,N_18592,N_18746);
and U19268 (N_19268,N_18540,N_18547);
nand U19269 (N_19269,N_18369,N_18127);
or U19270 (N_19270,N_18192,N_18201);
nand U19271 (N_19271,N_18549,N_18232);
xnor U19272 (N_19272,N_18222,N_18199);
and U19273 (N_19273,N_18238,N_18716);
nand U19274 (N_19274,N_18706,N_18672);
nor U19275 (N_19275,N_18715,N_18477);
nand U19276 (N_19276,N_18742,N_18382);
nor U19277 (N_19277,N_18541,N_18276);
nor U19278 (N_19278,N_18272,N_18305);
xor U19279 (N_19279,N_18526,N_18471);
nand U19280 (N_19280,N_18494,N_18639);
xnor U19281 (N_19281,N_18522,N_18326);
and U19282 (N_19282,N_18409,N_18258);
nand U19283 (N_19283,N_18359,N_18302);
nor U19284 (N_19284,N_18326,N_18289);
xor U19285 (N_19285,N_18663,N_18576);
nand U19286 (N_19286,N_18153,N_18189);
nor U19287 (N_19287,N_18497,N_18350);
nand U19288 (N_19288,N_18518,N_18264);
or U19289 (N_19289,N_18495,N_18467);
nand U19290 (N_19290,N_18682,N_18673);
xor U19291 (N_19291,N_18416,N_18373);
nor U19292 (N_19292,N_18473,N_18630);
and U19293 (N_19293,N_18738,N_18674);
and U19294 (N_19294,N_18711,N_18678);
nor U19295 (N_19295,N_18579,N_18175);
nand U19296 (N_19296,N_18204,N_18621);
nor U19297 (N_19297,N_18151,N_18448);
and U19298 (N_19298,N_18217,N_18293);
nand U19299 (N_19299,N_18491,N_18721);
nor U19300 (N_19300,N_18713,N_18449);
nor U19301 (N_19301,N_18641,N_18269);
and U19302 (N_19302,N_18711,N_18278);
or U19303 (N_19303,N_18616,N_18391);
nor U19304 (N_19304,N_18368,N_18605);
and U19305 (N_19305,N_18320,N_18206);
or U19306 (N_19306,N_18323,N_18387);
xnor U19307 (N_19307,N_18747,N_18201);
nor U19308 (N_19308,N_18417,N_18157);
xnor U19309 (N_19309,N_18135,N_18397);
xnor U19310 (N_19310,N_18398,N_18220);
or U19311 (N_19311,N_18675,N_18281);
nand U19312 (N_19312,N_18671,N_18394);
nor U19313 (N_19313,N_18557,N_18443);
and U19314 (N_19314,N_18642,N_18676);
xnor U19315 (N_19315,N_18135,N_18186);
or U19316 (N_19316,N_18469,N_18166);
and U19317 (N_19317,N_18689,N_18288);
nor U19318 (N_19318,N_18331,N_18266);
nand U19319 (N_19319,N_18160,N_18376);
and U19320 (N_19320,N_18476,N_18352);
nand U19321 (N_19321,N_18191,N_18331);
nor U19322 (N_19322,N_18563,N_18663);
xnor U19323 (N_19323,N_18345,N_18695);
xor U19324 (N_19324,N_18244,N_18745);
or U19325 (N_19325,N_18585,N_18199);
nand U19326 (N_19326,N_18194,N_18207);
or U19327 (N_19327,N_18732,N_18412);
nor U19328 (N_19328,N_18430,N_18244);
xor U19329 (N_19329,N_18274,N_18563);
and U19330 (N_19330,N_18362,N_18304);
and U19331 (N_19331,N_18429,N_18709);
or U19332 (N_19332,N_18544,N_18694);
and U19333 (N_19333,N_18138,N_18478);
and U19334 (N_19334,N_18366,N_18185);
nor U19335 (N_19335,N_18530,N_18192);
and U19336 (N_19336,N_18178,N_18218);
nor U19337 (N_19337,N_18374,N_18338);
and U19338 (N_19338,N_18277,N_18736);
xnor U19339 (N_19339,N_18180,N_18399);
or U19340 (N_19340,N_18347,N_18639);
nand U19341 (N_19341,N_18298,N_18658);
and U19342 (N_19342,N_18480,N_18721);
nand U19343 (N_19343,N_18541,N_18181);
or U19344 (N_19344,N_18515,N_18342);
nand U19345 (N_19345,N_18184,N_18319);
xnor U19346 (N_19346,N_18208,N_18688);
nand U19347 (N_19347,N_18188,N_18348);
and U19348 (N_19348,N_18293,N_18269);
xnor U19349 (N_19349,N_18250,N_18588);
nand U19350 (N_19350,N_18458,N_18619);
or U19351 (N_19351,N_18468,N_18559);
xor U19352 (N_19352,N_18739,N_18564);
xnor U19353 (N_19353,N_18168,N_18614);
xnor U19354 (N_19354,N_18388,N_18651);
nor U19355 (N_19355,N_18728,N_18318);
or U19356 (N_19356,N_18399,N_18670);
and U19357 (N_19357,N_18696,N_18195);
and U19358 (N_19358,N_18690,N_18525);
and U19359 (N_19359,N_18411,N_18407);
nor U19360 (N_19360,N_18432,N_18126);
nor U19361 (N_19361,N_18525,N_18423);
and U19362 (N_19362,N_18376,N_18573);
xnor U19363 (N_19363,N_18724,N_18693);
nand U19364 (N_19364,N_18605,N_18654);
and U19365 (N_19365,N_18630,N_18549);
nand U19366 (N_19366,N_18570,N_18600);
and U19367 (N_19367,N_18493,N_18723);
and U19368 (N_19368,N_18494,N_18170);
or U19369 (N_19369,N_18167,N_18249);
and U19370 (N_19370,N_18266,N_18613);
xnor U19371 (N_19371,N_18333,N_18259);
and U19372 (N_19372,N_18567,N_18184);
nand U19373 (N_19373,N_18492,N_18377);
or U19374 (N_19374,N_18501,N_18363);
nor U19375 (N_19375,N_19072,N_18773);
or U19376 (N_19376,N_18936,N_19358);
xnor U19377 (N_19377,N_19241,N_18981);
or U19378 (N_19378,N_19347,N_18763);
nor U19379 (N_19379,N_19034,N_18872);
nor U19380 (N_19380,N_19143,N_19321);
and U19381 (N_19381,N_19018,N_19170);
and U19382 (N_19382,N_18991,N_19368);
nand U19383 (N_19383,N_19312,N_18964);
nor U19384 (N_19384,N_19235,N_19144);
and U19385 (N_19385,N_19129,N_19017);
and U19386 (N_19386,N_18977,N_19046);
or U19387 (N_19387,N_19128,N_19298);
or U19388 (N_19388,N_19247,N_18846);
xor U19389 (N_19389,N_18770,N_18783);
nand U19390 (N_19390,N_19112,N_19103);
nand U19391 (N_19391,N_19373,N_18759);
nor U19392 (N_19392,N_19332,N_19336);
xnor U19393 (N_19393,N_18864,N_19165);
nor U19394 (N_19394,N_18778,N_19113);
nor U19395 (N_19395,N_19300,N_19320);
nand U19396 (N_19396,N_18942,N_19331);
or U19397 (N_19397,N_19201,N_19360);
xnor U19398 (N_19398,N_18824,N_19123);
nor U19399 (N_19399,N_18779,N_19028);
xor U19400 (N_19400,N_19345,N_19319);
or U19401 (N_19401,N_19192,N_19293);
xor U19402 (N_19402,N_18948,N_18762);
and U19403 (N_19403,N_19288,N_18971);
nand U19404 (N_19404,N_19096,N_18951);
xor U19405 (N_19405,N_18842,N_19250);
nand U19406 (N_19406,N_18799,N_19349);
or U19407 (N_19407,N_18758,N_18999);
nand U19408 (N_19408,N_18751,N_19278);
xnor U19409 (N_19409,N_19374,N_19085);
and U19410 (N_19410,N_19295,N_18768);
nor U19411 (N_19411,N_19038,N_19063);
nor U19412 (N_19412,N_18774,N_18818);
xor U19413 (N_19413,N_19140,N_18823);
nand U19414 (N_19414,N_19111,N_18884);
and U19415 (N_19415,N_19037,N_19322);
nand U19416 (N_19416,N_19166,N_18767);
nand U19417 (N_19417,N_18754,N_18932);
xnor U19418 (N_19418,N_19266,N_18979);
nand U19419 (N_19419,N_18902,N_18817);
and U19420 (N_19420,N_19045,N_18944);
nor U19421 (N_19421,N_18895,N_19048);
and U19422 (N_19422,N_18809,N_19154);
nor U19423 (N_19423,N_19093,N_19196);
and U19424 (N_19424,N_19204,N_19245);
nand U19425 (N_19425,N_19229,N_18924);
nand U19426 (N_19426,N_18963,N_18943);
and U19427 (N_19427,N_19198,N_19289);
or U19428 (N_19428,N_19000,N_19348);
xnor U19429 (N_19429,N_19011,N_19359);
nor U19430 (N_19430,N_19306,N_18791);
nand U19431 (N_19431,N_18833,N_18968);
or U19432 (N_19432,N_18998,N_19127);
xnor U19433 (N_19433,N_19267,N_18929);
and U19434 (N_19434,N_18966,N_18816);
xnor U19435 (N_19435,N_19148,N_19286);
nor U19436 (N_19436,N_19107,N_19169);
xor U19437 (N_19437,N_18920,N_19133);
xnor U19438 (N_19438,N_18992,N_19016);
nand U19439 (N_19439,N_18852,N_19279);
or U19440 (N_19440,N_19032,N_19095);
xnor U19441 (N_19441,N_19369,N_18813);
nand U19442 (N_19442,N_19262,N_18826);
or U19443 (N_19443,N_18910,N_19182);
and U19444 (N_19444,N_19013,N_19342);
and U19445 (N_19445,N_19294,N_18873);
or U19446 (N_19446,N_19364,N_19179);
nor U19447 (N_19447,N_18757,N_18851);
nor U19448 (N_19448,N_18837,N_19118);
xor U19449 (N_19449,N_19268,N_19310);
nor U19450 (N_19450,N_19053,N_18875);
nor U19451 (N_19451,N_19339,N_18900);
nand U19452 (N_19452,N_19015,N_19173);
xnor U19453 (N_19453,N_18814,N_18939);
and U19454 (N_19454,N_19365,N_18993);
nor U19455 (N_19455,N_18804,N_19010);
nand U19456 (N_19456,N_18752,N_18806);
and U19457 (N_19457,N_18792,N_19197);
xnor U19458 (N_19458,N_19226,N_18810);
nand U19459 (N_19459,N_18937,N_19067);
nor U19460 (N_19460,N_19051,N_18974);
or U19461 (N_19461,N_18927,N_18881);
nand U19462 (N_19462,N_18844,N_18866);
xor U19463 (N_19463,N_19090,N_19005);
or U19464 (N_19464,N_18775,N_19210);
nor U19465 (N_19465,N_19185,N_18784);
and U19466 (N_19466,N_19263,N_18938);
and U19467 (N_19467,N_19184,N_18893);
nand U19468 (N_19468,N_19305,N_18917);
or U19469 (N_19469,N_19270,N_19271);
and U19470 (N_19470,N_18878,N_18946);
nand U19471 (N_19471,N_18961,N_19340);
and U19472 (N_19472,N_19054,N_19157);
or U19473 (N_19473,N_18795,N_18868);
xor U19474 (N_19474,N_19042,N_19071);
nor U19475 (N_19475,N_18840,N_18984);
nand U19476 (N_19476,N_19134,N_18827);
xnor U19477 (N_19477,N_19175,N_18997);
nand U19478 (N_19478,N_19301,N_18959);
xor U19479 (N_19479,N_19341,N_19007);
nand U19480 (N_19480,N_18887,N_18975);
nand U19481 (N_19481,N_19338,N_19035);
xor U19482 (N_19482,N_19138,N_19215);
xnor U19483 (N_19483,N_19174,N_18780);
nand U19484 (N_19484,N_18858,N_19002);
or U19485 (N_19485,N_19292,N_18908);
nor U19486 (N_19486,N_18801,N_19323);
and U19487 (N_19487,N_18967,N_19132);
and U19488 (N_19488,N_19328,N_19163);
nor U19489 (N_19489,N_19052,N_18987);
or U19490 (N_19490,N_19251,N_19239);
nand U19491 (N_19491,N_19216,N_18996);
xor U19492 (N_19492,N_18947,N_19199);
xnor U19493 (N_19493,N_18867,N_19167);
and U19494 (N_19494,N_19104,N_18808);
nor U19495 (N_19495,N_19337,N_18901);
nand U19496 (N_19496,N_18822,N_18834);
nor U19497 (N_19497,N_19207,N_19187);
nand U19498 (N_19498,N_19205,N_18897);
nor U19499 (N_19499,N_19194,N_18886);
and U19500 (N_19500,N_18850,N_19316);
or U19501 (N_19501,N_19022,N_19209);
nand U19502 (N_19502,N_18956,N_19073);
and U19503 (N_19503,N_18843,N_18853);
nor U19504 (N_19504,N_18894,N_19162);
or U19505 (N_19505,N_19047,N_19080);
xnor U19506 (N_19506,N_19109,N_19367);
xnor U19507 (N_19507,N_19152,N_19308);
xor U19508 (N_19508,N_19146,N_19353);
nor U19509 (N_19509,N_18880,N_19177);
xor U19510 (N_19510,N_19257,N_18877);
and U19511 (N_19511,N_18766,N_18906);
xnor U19512 (N_19512,N_19275,N_18849);
nand U19513 (N_19513,N_19325,N_18941);
xnor U19514 (N_19514,N_18934,N_18945);
nor U19515 (N_19515,N_18835,N_19131);
nand U19516 (N_19516,N_19222,N_18848);
or U19517 (N_19517,N_18865,N_18776);
and U19518 (N_19518,N_19105,N_19290);
or U19519 (N_19519,N_19237,N_19108);
xnor U19520 (N_19520,N_19183,N_19062);
nor U19521 (N_19521,N_18800,N_19168);
or U19522 (N_19522,N_18830,N_19036);
and U19523 (N_19523,N_18916,N_19003);
nor U19524 (N_19524,N_19001,N_19049);
nor U19525 (N_19525,N_18811,N_19137);
nor U19526 (N_19526,N_19069,N_18871);
or U19527 (N_19527,N_19252,N_19091);
nand U19528 (N_19528,N_18957,N_19060);
or U19529 (N_19529,N_19055,N_19160);
and U19530 (N_19530,N_18876,N_19248);
or U19531 (N_19531,N_19351,N_19021);
or U19532 (N_19532,N_18790,N_19097);
or U19533 (N_19533,N_19086,N_18860);
xor U19534 (N_19534,N_19343,N_19302);
nor U19535 (N_19535,N_19064,N_19020);
xor U19536 (N_19536,N_19119,N_19297);
nand U19537 (N_19537,N_18986,N_19050);
and U19538 (N_19538,N_19335,N_19125);
and U19539 (N_19539,N_18892,N_19158);
xor U19540 (N_19540,N_18962,N_18976);
or U19541 (N_19541,N_19024,N_19083);
and U19542 (N_19542,N_19202,N_19188);
and U19543 (N_19543,N_19136,N_19027);
and U19544 (N_19544,N_18952,N_18965);
xor U19545 (N_19545,N_18926,N_19200);
nor U19546 (N_19546,N_19043,N_18782);
nand U19547 (N_19547,N_19161,N_19078);
and U19548 (N_19548,N_19004,N_19372);
nor U19549 (N_19549,N_18930,N_18898);
or U19550 (N_19550,N_19232,N_18983);
nor U19551 (N_19551,N_18950,N_19041);
or U19552 (N_19552,N_18879,N_19285);
and U19553 (N_19553,N_19361,N_19317);
nand U19554 (N_19554,N_18777,N_19178);
nor U19555 (N_19555,N_19159,N_19324);
nor U19556 (N_19556,N_18863,N_19044);
nor U19557 (N_19557,N_19012,N_19203);
xor U19558 (N_19558,N_18911,N_19130);
xnor U19559 (N_19559,N_19371,N_18785);
xnor U19560 (N_19560,N_18969,N_18885);
xor U19561 (N_19561,N_19304,N_19150);
xor U19562 (N_19562,N_19244,N_18995);
and U19563 (N_19563,N_19327,N_19224);
xnor U19564 (N_19564,N_18793,N_18953);
or U19565 (N_19565,N_18903,N_19121);
nor U19566 (N_19566,N_18954,N_19234);
xor U19567 (N_19567,N_19075,N_19307);
and U19568 (N_19568,N_18819,N_19076);
nand U19569 (N_19569,N_19274,N_19070);
nor U19570 (N_19570,N_19287,N_18909);
nor U19571 (N_19571,N_19106,N_19040);
nor U19572 (N_19572,N_19029,N_18781);
xnor U19573 (N_19573,N_18980,N_19124);
and U19574 (N_19574,N_18803,N_19217);
nand U19575 (N_19575,N_19366,N_19259);
or U19576 (N_19576,N_18847,N_18854);
xor U19577 (N_19577,N_19296,N_19284);
nand U19578 (N_19578,N_19115,N_19006);
nand U19579 (N_19579,N_19151,N_19065);
or U19580 (N_19580,N_19212,N_19068);
or U19581 (N_19581,N_19147,N_19344);
nand U19582 (N_19582,N_18805,N_18859);
or U19583 (N_19583,N_18841,N_19171);
nand U19584 (N_19584,N_18789,N_19329);
xor U19585 (N_19585,N_19087,N_19219);
nor U19586 (N_19586,N_18925,N_19238);
nand U19587 (N_19587,N_18772,N_19153);
or U19588 (N_19588,N_18845,N_19280);
xor U19589 (N_19589,N_18891,N_18982);
or U19590 (N_19590,N_19370,N_19145);
nand U19591 (N_19591,N_18988,N_19318);
or U19592 (N_19592,N_19311,N_19357);
nor U19593 (N_19593,N_18883,N_19142);
nand U19594 (N_19594,N_18755,N_19180);
and U19595 (N_19595,N_18828,N_18855);
nand U19596 (N_19596,N_19117,N_19026);
nand U19597 (N_19597,N_18882,N_19155);
nand U19598 (N_19598,N_19314,N_19208);
xor U19599 (N_19599,N_18921,N_18861);
nor U19600 (N_19600,N_18821,N_19057);
xor U19601 (N_19601,N_18890,N_19030);
xor U19602 (N_19602,N_18958,N_19084);
or U19603 (N_19603,N_18857,N_18912);
nor U19604 (N_19604,N_18940,N_18896);
xor U19605 (N_19605,N_19309,N_18972);
nor U19606 (N_19606,N_18933,N_18862);
nand U19607 (N_19607,N_18838,N_19223);
or U19608 (N_19608,N_19242,N_18787);
nand U19609 (N_19609,N_18960,N_18753);
nand U19610 (N_19610,N_19092,N_19291);
or U19611 (N_19611,N_18904,N_19008);
nor U19612 (N_19612,N_19066,N_19258);
or U19613 (N_19613,N_19355,N_19077);
or U19614 (N_19614,N_19099,N_19326);
or U19615 (N_19615,N_19236,N_19214);
nor U19616 (N_19616,N_18764,N_19283);
or U19617 (N_19617,N_19277,N_18989);
and U19618 (N_19618,N_19061,N_19303);
or U19619 (N_19619,N_19126,N_19135);
nor U19620 (N_19620,N_19120,N_19354);
and U19621 (N_19621,N_19356,N_19246);
and U19622 (N_19622,N_18915,N_19033);
and U19623 (N_19623,N_18802,N_18907);
nor U19624 (N_19624,N_18990,N_18870);
xor U19625 (N_19625,N_19082,N_19272);
xor U19626 (N_19626,N_18831,N_18836);
xnor U19627 (N_19627,N_19114,N_18928);
nor U19628 (N_19628,N_19141,N_18978);
and U19629 (N_19629,N_19228,N_18913);
xor U19630 (N_19630,N_19352,N_18922);
or U19631 (N_19631,N_19206,N_19330);
xnor U19632 (N_19632,N_18949,N_19273);
or U19633 (N_19633,N_19265,N_18985);
xor U19634 (N_19634,N_19009,N_19260);
xnor U19635 (N_19635,N_18935,N_18869);
xor U19636 (N_19636,N_19088,N_19213);
and U19637 (N_19637,N_19313,N_19102);
nand U19638 (N_19638,N_19233,N_19346);
and U19639 (N_19639,N_18765,N_18905);
nor U19640 (N_19640,N_19264,N_19193);
or U19641 (N_19641,N_19195,N_19282);
nor U19642 (N_19642,N_19094,N_19190);
xnor U19643 (N_19643,N_18919,N_18761);
nor U19644 (N_19644,N_18756,N_19172);
nor U19645 (N_19645,N_18825,N_19059);
nand U19646 (N_19646,N_19220,N_19315);
nor U19647 (N_19647,N_19249,N_19019);
nand U19648 (N_19648,N_19254,N_19081);
nand U19649 (N_19649,N_19110,N_18786);
and U19650 (N_19650,N_19230,N_19281);
nand U19651 (N_19651,N_19074,N_18856);
nor U19652 (N_19652,N_19299,N_18788);
and U19653 (N_19653,N_18955,N_19014);
or U19654 (N_19654,N_19243,N_19149);
xor U19655 (N_19655,N_18839,N_18829);
nand U19656 (N_19656,N_19218,N_19101);
and U19657 (N_19657,N_18970,N_19276);
or U19658 (N_19658,N_19079,N_18931);
nor U19659 (N_19659,N_18973,N_18820);
nor U19660 (N_19660,N_18769,N_19122);
nand U19661 (N_19661,N_19253,N_19025);
xor U19662 (N_19662,N_19221,N_18918);
nor U19663 (N_19663,N_18923,N_18888);
nand U19664 (N_19664,N_19098,N_19227);
and U19665 (N_19665,N_18815,N_18914);
xor U19666 (N_19666,N_19191,N_19363);
and U19667 (N_19667,N_19181,N_19362);
nand U19668 (N_19668,N_19211,N_19031);
xor U19669 (N_19669,N_19176,N_19164);
nand U19670 (N_19670,N_18796,N_19116);
xor U19671 (N_19671,N_18889,N_19058);
xor U19672 (N_19672,N_18832,N_19269);
nor U19673 (N_19673,N_19189,N_18994);
and U19674 (N_19674,N_18798,N_18807);
or U19675 (N_19675,N_19156,N_19089);
nand U19676 (N_19676,N_19256,N_19333);
nand U19677 (N_19677,N_18750,N_18874);
nand U19678 (N_19678,N_19261,N_19231);
nand U19679 (N_19679,N_18812,N_19334);
nor U19680 (N_19680,N_18797,N_19139);
nand U19681 (N_19681,N_19350,N_19240);
nor U19682 (N_19682,N_19255,N_19023);
nor U19683 (N_19683,N_18899,N_18771);
nor U19684 (N_19684,N_19100,N_18794);
or U19685 (N_19685,N_19186,N_19039);
xnor U19686 (N_19686,N_19225,N_18760);
nand U19687 (N_19687,N_19056,N_18860);
nand U19688 (N_19688,N_19121,N_19221);
nor U19689 (N_19689,N_18817,N_19334);
or U19690 (N_19690,N_19049,N_19005);
nor U19691 (N_19691,N_18937,N_18876);
nand U19692 (N_19692,N_19220,N_19351);
and U19693 (N_19693,N_18813,N_19302);
nand U19694 (N_19694,N_19368,N_18950);
and U19695 (N_19695,N_18819,N_19055);
and U19696 (N_19696,N_18811,N_18981);
nand U19697 (N_19697,N_19267,N_18888);
or U19698 (N_19698,N_18946,N_18910);
or U19699 (N_19699,N_19013,N_19207);
or U19700 (N_19700,N_18869,N_19257);
xnor U19701 (N_19701,N_18876,N_19355);
nor U19702 (N_19702,N_19234,N_18942);
or U19703 (N_19703,N_18900,N_18766);
nor U19704 (N_19704,N_19043,N_18788);
or U19705 (N_19705,N_19348,N_19074);
or U19706 (N_19706,N_18991,N_18963);
nor U19707 (N_19707,N_19157,N_18925);
nand U19708 (N_19708,N_18772,N_18924);
xor U19709 (N_19709,N_18974,N_18755);
nor U19710 (N_19710,N_18972,N_18803);
nand U19711 (N_19711,N_18755,N_19348);
xnor U19712 (N_19712,N_18760,N_18778);
and U19713 (N_19713,N_19366,N_19288);
and U19714 (N_19714,N_18777,N_19074);
nand U19715 (N_19715,N_19250,N_19057);
xor U19716 (N_19716,N_19042,N_19080);
nand U19717 (N_19717,N_19028,N_19158);
nand U19718 (N_19718,N_18907,N_19046);
nor U19719 (N_19719,N_19080,N_19210);
nand U19720 (N_19720,N_19205,N_18791);
nor U19721 (N_19721,N_18941,N_18966);
nand U19722 (N_19722,N_19358,N_18879);
nor U19723 (N_19723,N_18797,N_18874);
xor U19724 (N_19724,N_19125,N_18885);
nand U19725 (N_19725,N_18793,N_18832);
xor U19726 (N_19726,N_18930,N_19352);
xor U19727 (N_19727,N_18922,N_19065);
xor U19728 (N_19728,N_18765,N_18962);
and U19729 (N_19729,N_19337,N_18892);
and U19730 (N_19730,N_18759,N_18945);
nor U19731 (N_19731,N_18753,N_19277);
xnor U19732 (N_19732,N_19296,N_18800);
or U19733 (N_19733,N_18983,N_19318);
nand U19734 (N_19734,N_19225,N_19234);
and U19735 (N_19735,N_19182,N_19194);
and U19736 (N_19736,N_19374,N_19218);
and U19737 (N_19737,N_19050,N_18797);
xor U19738 (N_19738,N_18998,N_19247);
or U19739 (N_19739,N_19143,N_19148);
and U19740 (N_19740,N_18761,N_19361);
xnor U19741 (N_19741,N_18947,N_19283);
nor U19742 (N_19742,N_19184,N_18834);
and U19743 (N_19743,N_18778,N_19089);
xnor U19744 (N_19744,N_18776,N_19310);
and U19745 (N_19745,N_19248,N_19042);
and U19746 (N_19746,N_18962,N_18773);
and U19747 (N_19747,N_19165,N_18839);
and U19748 (N_19748,N_18801,N_19331);
xnor U19749 (N_19749,N_18930,N_18952);
nor U19750 (N_19750,N_18757,N_19097);
xnor U19751 (N_19751,N_18932,N_19242);
nor U19752 (N_19752,N_19374,N_19055);
or U19753 (N_19753,N_19305,N_19236);
and U19754 (N_19754,N_18899,N_19324);
nand U19755 (N_19755,N_19325,N_18776);
xor U19756 (N_19756,N_19119,N_19363);
xnor U19757 (N_19757,N_18979,N_19342);
and U19758 (N_19758,N_19008,N_19115);
nand U19759 (N_19759,N_19038,N_18998);
or U19760 (N_19760,N_18912,N_19020);
nor U19761 (N_19761,N_18832,N_18787);
nand U19762 (N_19762,N_19148,N_19185);
nand U19763 (N_19763,N_18777,N_19344);
xor U19764 (N_19764,N_19014,N_19021);
or U19765 (N_19765,N_19111,N_19082);
nor U19766 (N_19766,N_19077,N_19283);
nand U19767 (N_19767,N_19032,N_19184);
nand U19768 (N_19768,N_18834,N_19054);
nand U19769 (N_19769,N_19107,N_19256);
nor U19770 (N_19770,N_19016,N_18983);
or U19771 (N_19771,N_19091,N_19261);
or U19772 (N_19772,N_18757,N_18767);
xor U19773 (N_19773,N_18813,N_19191);
xnor U19774 (N_19774,N_19200,N_19350);
xor U19775 (N_19775,N_19111,N_19190);
nor U19776 (N_19776,N_19192,N_19077);
and U19777 (N_19777,N_19163,N_18896);
or U19778 (N_19778,N_18946,N_19193);
xor U19779 (N_19779,N_18876,N_19033);
nand U19780 (N_19780,N_18909,N_18974);
nor U19781 (N_19781,N_18783,N_19164);
nand U19782 (N_19782,N_19371,N_19303);
nor U19783 (N_19783,N_19215,N_18941);
or U19784 (N_19784,N_19145,N_19277);
nand U19785 (N_19785,N_18993,N_19081);
nand U19786 (N_19786,N_18956,N_18999);
xor U19787 (N_19787,N_18877,N_18802);
xor U19788 (N_19788,N_19123,N_18859);
nor U19789 (N_19789,N_18913,N_19172);
and U19790 (N_19790,N_19263,N_19034);
xor U19791 (N_19791,N_18772,N_19038);
or U19792 (N_19792,N_18857,N_19051);
and U19793 (N_19793,N_19075,N_18873);
or U19794 (N_19794,N_18759,N_19043);
or U19795 (N_19795,N_19227,N_18751);
and U19796 (N_19796,N_19218,N_18875);
nor U19797 (N_19797,N_19208,N_18855);
nand U19798 (N_19798,N_18835,N_18912);
or U19799 (N_19799,N_19198,N_18775);
xor U19800 (N_19800,N_19340,N_18939);
or U19801 (N_19801,N_19218,N_18893);
xor U19802 (N_19802,N_19180,N_19274);
or U19803 (N_19803,N_19171,N_19225);
nor U19804 (N_19804,N_19166,N_19136);
and U19805 (N_19805,N_19298,N_18777);
nor U19806 (N_19806,N_19052,N_19214);
nand U19807 (N_19807,N_19015,N_19098);
nand U19808 (N_19808,N_19163,N_19345);
and U19809 (N_19809,N_19174,N_18918);
and U19810 (N_19810,N_19252,N_19103);
and U19811 (N_19811,N_18891,N_18981);
and U19812 (N_19812,N_18853,N_19044);
xor U19813 (N_19813,N_18774,N_19354);
xnor U19814 (N_19814,N_19229,N_19236);
nand U19815 (N_19815,N_19369,N_18891);
nand U19816 (N_19816,N_18820,N_18762);
nand U19817 (N_19817,N_19279,N_19274);
xor U19818 (N_19818,N_18885,N_19019);
and U19819 (N_19819,N_18998,N_18803);
nand U19820 (N_19820,N_18859,N_18806);
nor U19821 (N_19821,N_19336,N_18906);
nor U19822 (N_19822,N_19098,N_19060);
xor U19823 (N_19823,N_19085,N_18874);
or U19824 (N_19824,N_18868,N_19332);
or U19825 (N_19825,N_19189,N_18993);
nand U19826 (N_19826,N_18956,N_18757);
and U19827 (N_19827,N_19208,N_19003);
and U19828 (N_19828,N_19200,N_19033);
and U19829 (N_19829,N_19136,N_19087);
nand U19830 (N_19830,N_19312,N_18762);
nand U19831 (N_19831,N_18752,N_18783);
nor U19832 (N_19832,N_19247,N_19045);
and U19833 (N_19833,N_18896,N_18760);
nand U19834 (N_19834,N_18822,N_19169);
and U19835 (N_19835,N_18781,N_19061);
nand U19836 (N_19836,N_19340,N_18806);
nand U19837 (N_19837,N_19275,N_19022);
and U19838 (N_19838,N_19032,N_18840);
or U19839 (N_19839,N_19092,N_18968);
xor U19840 (N_19840,N_18814,N_18947);
nand U19841 (N_19841,N_19109,N_18991);
or U19842 (N_19842,N_19182,N_18826);
and U19843 (N_19843,N_18954,N_19073);
and U19844 (N_19844,N_19227,N_19269);
or U19845 (N_19845,N_19189,N_19230);
and U19846 (N_19846,N_18769,N_19055);
nand U19847 (N_19847,N_19364,N_18889);
nor U19848 (N_19848,N_18754,N_19322);
and U19849 (N_19849,N_18792,N_18811);
and U19850 (N_19850,N_18786,N_19081);
nand U19851 (N_19851,N_18835,N_18960);
or U19852 (N_19852,N_18786,N_19193);
nor U19853 (N_19853,N_19317,N_19088);
and U19854 (N_19854,N_19124,N_19283);
xnor U19855 (N_19855,N_19229,N_19053);
nand U19856 (N_19856,N_19166,N_18871);
or U19857 (N_19857,N_19213,N_19262);
or U19858 (N_19858,N_18831,N_19330);
or U19859 (N_19859,N_19230,N_19114);
xnor U19860 (N_19860,N_18952,N_19325);
and U19861 (N_19861,N_19105,N_19269);
nor U19862 (N_19862,N_19286,N_18839);
or U19863 (N_19863,N_19091,N_18834);
xor U19864 (N_19864,N_19258,N_18858);
xor U19865 (N_19865,N_19036,N_18786);
or U19866 (N_19866,N_19089,N_19073);
and U19867 (N_19867,N_19278,N_19339);
nor U19868 (N_19868,N_19066,N_19094);
nor U19869 (N_19869,N_19127,N_19006);
nand U19870 (N_19870,N_19259,N_18889);
and U19871 (N_19871,N_19182,N_19227);
or U19872 (N_19872,N_18984,N_19263);
or U19873 (N_19873,N_18760,N_18941);
xnor U19874 (N_19874,N_19021,N_19331);
xnor U19875 (N_19875,N_18879,N_18751);
or U19876 (N_19876,N_18903,N_19373);
nor U19877 (N_19877,N_19211,N_19001);
nand U19878 (N_19878,N_19154,N_19361);
nand U19879 (N_19879,N_19102,N_18910);
or U19880 (N_19880,N_19137,N_19101);
and U19881 (N_19881,N_19286,N_19082);
or U19882 (N_19882,N_18922,N_19055);
xor U19883 (N_19883,N_18816,N_19317);
nand U19884 (N_19884,N_19205,N_19275);
and U19885 (N_19885,N_18927,N_18940);
xnor U19886 (N_19886,N_18952,N_18905);
and U19887 (N_19887,N_18774,N_19215);
xor U19888 (N_19888,N_18942,N_19335);
xnor U19889 (N_19889,N_19008,N_18951);
nor U19890 (N_19890,N_19166,N_19232);
nor U19891 (N_19891,N_19299,N_19075);
or U19892 (N_19892,N_19031,N_19135);
nand U19893 (N_19893,N_19062,N_19015);
nand U19894 (N_19894,N_18827,N_19341);
and U19895 (N_19895,N_18792,N_18997);
and U19896 (N_19896,N_19222,N_19112);
and U19897 (N_19897,N_19307,N_18832);
nand U19898 (N_19898,N_19371,N_18823);
nand U19899 (N_19899,N_19058,N_19002);
nand U19900 (N_19900,N_18777,N_18835);
or U19901 (N_19901,N_18835,N_19330);
nand U19902 (N_19902,N_18929,N_18790);
or U19903 (N_19903,N_18946,N_18876);
or U19904 (N_19904,N_19373,N_18973);
nor U19905 (N_19905,N_18780,N_19055);
or U19906 (N_19906,N_18916,N_18965);
or U19907 (N_19907,N_18795,N_18936);
xor U19908 (N_19908,N_19227,N_19019);
nor U19909 (N_19909,N_19213,N_19169);
xor U19910 (N_19910,N_18895,N_19142);
xnor U19911 (N_19911,N_19197,N_19044);
nor U19912 (N_19912,N_18868,N_18781);
nor U19913 (N_19913,N_18776,N_18882);
nor U19914 (N_19914,N_19016,N_19155);
or U19915 (N_19915,N_18824,N_18892);
nand U19916 (N_19916,N_18878,N_19022);
and U19917 (N_19917,N_19130,N_19242);
xor U19918 (N_19918,N_18823,N_18817);
xnor U19919 (N_19919,N_18790,N_18966);
xor U19920 (N_19920,N_18953,N_18946);
or U19921 (N_19921,N_19330,N_18907);
xor U19922 (N_19922,N_19025,N_19055);
nor U19923 (N_19923,N_18892,N_18760);
nor U19924 (N_19924,N_18844,N_18878);
or U19925 (N_19925,N_19316,N_18929);
nor U19926 (N_19926,N_19050,N_18928);
or U19927 (N_19927,N_18939,N_19055);
and U19928 (N_19928,N_18754,N_19171);
nand U19929 (N_19929,N_19275,N_18922);
or U19930 (N_19930,N_19245,N_18991);
nand U19931 (N_19931,N_19280,N_19033);
or U19932 (N_19932,N_19207,N_18965);
and U19933 (N_19933,N_19133,N_19090);
xnor U19934 (N_19934,N_19330,N_19271);
nor U19935 (N_19935,N_18886,N_18958);
and U19936 (N_19936,N_19348,N_19061);
or U19937 (N_19937,N_19368,N_19196);
and U19938 (N_19938,N_19096,N_19163);
xor U19939 (N_19939,N_19373,N_19237);
nor U19940 (N_19940,N_19211,N_19068);
nor U19941 (N_19941,N_18769,N_18974);
nor U19942 (N_19942,N_19064,N_19074);
nand U19943 (N_19943,N_19216,N_19044);
or U19944 (N_19944,N_19044,N_19204);
or U19945 (N_19945,N_18785,N_19342);
and U19946 (N_19946,N_18790,N_18779);
and U19947 (N_19947,N_19157,N_19194);
or U19948 (N_19948,N_18900,N_19209);
and U19949 (N_19949,N_19333,N_19307);
or U19950 (N_19950,N_18787,N_18895);
xor U19951 (N_19951,N_18926,N_19351);
and U19952 (N_19952,N_19042,N_19298);
or U19953 (N_19953,N_19203,N_19051);
xnor U19954 (N_19954,N_18754,N_19114);
or U19955 (N_19955,N_18796,N_19329);
and U19956 (N_19956,N_19354,N_18807);
and U19957 (N_19957,N_18805,N_18961);
nor U19958 (N_19958,N_19021,N_19215);
and U19959 (N_19959,N_19087,N_19225);
xnor U19960 (N_19960,N_19326,N_19141);
nand U19961 (N_19961,N_19035,N_19000);
xnor U19962 (N_19962,N_18915,N_19349);
nor U19963 (N_19963,N_18804,N_19121);
and U19964 (N_19964,N_19315,N_19178);
and U19965 (N_19965,N_19003,N_18763);
nor U19966 (N_19966,N_18831,N_19231);
and U19967 (N_19967,N_18880,N_19305);
xor U19968 (N_19968,N_18961,N_18938);
nand U19969 (N_19969,N_19334,N_19145);
nand U19970 (N_19970,N_18846,N_19253);
nor U19971 (N_19971,N_19018,N_18904);
xor U19972 (N_19972,N_18867,N_19365);
and U19973 (N_19973,N_18837,N_19198);
xnor U19974 (N_19974,N_18890,N_18871);
or U19975 (N_19975,N_19371,N_19272);
nor U19976 (N_19976,N_19253,N_18971);
and U19977 (N_19977,N_18783,N_19313);
nor U19978 (N_19978,N_19176,N_18941);
or U19979 (N_19979,N_19066,N_19296);
and U19980 (N_19980,N_18951,N_19226);
nor U19981 (N_19981,N_19090,N_18814);
nor U19982 (N_19982,N_19221,N_19241);
xnor U19983 (N_19983,N_18773,N_19036);
nand U19984 (N_19984,N_18895,N_18906);
nand U19985 (N_19985,N_18916,N_18959);
nor U19986 (N_19986,N_18873,N_18940);
xnor U19987 (N_19987,N_19210,N_18861);
xor U19988 (N_19988,N_18754,N_18873);
and U19989 (N_19989,N_19333,N_18881);
nor U19990 (N_19990,N_19074,N_19042);
nor U19991 (N_19991,N_18903,N_19131);
nand U19992 (N_19992,N_19217,N_18849);
and U19993 (N_19993,N_19099,N_19035);
xor U19994 (N_19994,N_19373,N_18929);
nor U19995 (N_19995,N_18958,N_19318);
and U19996 (N_19996,N_19294,N_19352);
or U19997 (N_19997,N_19281,N_19325);
xnor U19998 (N_19998,N_19121,N_19109);
and U19999 (N_19999,N_19101,N_19225);
or U20000 (N_20000,N_19967,N_19397);
or U20001 (N_20001,N_19625,N_19880);
and U20002 (N_20002,N_19960,N_19556);
nor U20003 (N_20003,N_19451,N_19863);
nor U20004 (N_20004,N_19641,N_19929);
xor U20005 (N_20005,N_19998,N_19564);
xnor U20006 (N_20006,N_19622,N_19777);
or U20007 (N_20007,N_19817,N_19485);
xnor U20008 (N_20008,N_19944,N_19838);
nand U20009 (N_20009,N_19923,N_19444);
or U20010 (N_20010,N_19673,N_19710);
or U20011 (N_20011,N_19836,N_19523);
and U20012 (N_20012,N_19380,N_19391);
or U20013 (N_20013,N_19878,N_19437);
and U20014 (N_20014,N_19434,N_19683);
and U20015 (N_20015,N_19847,N_19720);
or U20016 (N_20016,N_19974,N_19454);
nand U20017 (N_20017,N_19565,N_19729);
or U20018 (N_20018,N_19956,N_19870);
and U20019 (N_20019,N_19694,N_19616);
xor U20020 (N_20020,N_19389,N_19457);
nor U20021 (N_20021,N_19471,N_19696);
and U20022 (N_20022,N_19644,N_19885);
or U20023 (N_20023,N_19855,N_19468);
nor U20024 (N_20024,N_19558,N_19527);
xnor U20025 (N_20025,N_19590,N_19536);
nor U20026 (N_20026,N_19497,N_19733);
and U20027 (N_20027,N_19445,N_19781);
nor U20028 (N_20028,N_19830,N_19927);
or U20029 (N_20029,N_19749,N_19959);
or U20030 (N_20030,N_19902,N_19428);
nand U20031 (N_20031,N_19766,N_19841);
and U20032 (N_20032,N_19946,N_19779);
xor U20033 (N_20033,N_19893,N_19985);
xor U20034 (N_20034,N_19381,N_19645);
nor U20035 (N_20035,N_19414,N_19996);
and U20036 (N_20036,N_19529,N_19966);
nor U20037 (N_20037,N_19816,N_19795);
or U20038 (N_20038,N_19970,N_19842);
and U20039 (N_20039,N_19657,N_19859);
nor U20040 (N_20040,N_19964,N_19499);
or U20041 (N_20041,N_19890,N_19634);
xor U20042 (N_20042,N_19753,N_19759);
or U20043 (N_20043,N_19768,N_19783);
nor U20044 (N_20044,N_19422,N_19624);
or U20045 (N_20045,N_19578,N_19399);
or U20046 (N_20046,N_19375,N_19747);
nand U20047 (N_20047,N_19839,N_19463);
or U20048 (N_20048,N_19488,N_19544);
nand U20049 (N_20049,N_19767,N_19543);
and U20050 (N_20050,N_19501,N_19689);
and U20051 (N_20051,N_19553,N_19631);
xnor U20052 (N_20052,N_19494,N_19411);
nand U20053 (N_20053,N_19953,N_19522);
nor U20054 (N_20054,N_19933,N_19937);
xnor U20055 (N_20055,N_19828,N_19732);
and U20056 (N_20056,N_19586,N_19498);
xor U20057 (N_20057,N_19585,N_19947);
nor U20058 (N_20058,N_19789,N_19515);
and U20059 (N_20059,N_19794,N_19793);
nor U20060 (N_20060,N_19980,N_19452);
or U20061 (N_20061,N_19849,N_19396);
and U20062 (N_20062,N_19466,N_19999);
and U20063 (N_20063,N_19879,N_19672);
nor U20064 (N_20064,N_19521,N_19442);
or U20065 (N_20065,N_19853,N_19909);
or U20066 (N_20066,N_19745,N_19426);
and U20067 (N_20067,N_19539,N_19739);
and U20068 (N_20068,N_19635,N_19924);
and U20069 (N_20069,N_19742,N_19570);
nor U20070 (N_20070,N_19934,N_19675);
or U20071 (N_20071,N_19713,N_19928);
nand U20072 (N_20072,N_19740,N_19984);
or U20073 (N_20073,N_19888,N_19982);
or U20074 (N_20074,N_19626,N_19693);
or U20075 (N_20075,N_19652,N_19404);
nand U20076 (N_20076,N_19801,N_19674);
nand U20077 (N_20077,N_19392,N_19459);
and U20078 (N_20078,N_19528,N_19531);
and U20079 (N_20079,N_19701,N_19555);
xnor U20080 (N_20080,N_19702,N_19919);
xnor U20081 (N_20081,N_19524,N_19416);
and U20082 (N_20082,N_19989,N_19541);
xnor U20083 (N_20083,N_19566,N_19867);
nor U20084 (N_20084,N_19695,N_19957);
or U20085 (N_20085,N_19512,N_19639);
nor U20086 (N_20086,N_19886,N_19548);
or U20087 (N_20087,N_19951,N_19973);
or U20088 (N_20088,N_19856,N_19925);
or U20089 (N_20089,N_19771,N_19874);
xor U20090 (N_20090,N_19606,N_19889);
nor U20091 (N_20091,N_19756,N_19572);
and U20092 (N_20092,N_19716,N_19509);
xnor U20093 (N_20093,N_19400,N_19687);
and U20094 (N_20094,N_19845,N_19976);
nand U20095 (N_20095,N_19386,N_19833);
xor U20096 (N_20096,N_19475,N_19642);
nor U20097 (N_20097,N_19649,N_19752);
nand U20098 (N_20098,N_19637,N_19792);
or U20099 (N_20099,N_19419,N_19580);
xor U20100 (N_20100,N_19587,N_19723);
and U20101 (N_20101,N_19395,N_19782);
xnor U20102 (N_20102,N_19837,N_19791);
or U20103 (N_20103,N_19881,N_19812);
nand U20104 (N_20104,N_19744,N_19787);
or U20105 (N_20105,N_19772,N_19507);
nand U20106 (N_20106,N_19861,N_19907);
or U20107 (N_20107,N_19872,N_19832);
or U20108 (N_20108,N_19605,N_19715);
nor U20109 (N_20109,N_19731,N_19894);
nand U20110 (N_20110,N_19986,N_19458);
and U20111 (N_20111,N_19711,N_19895);
xnor U20112 (N_20112,N_19981,N_19450);
nand U20113 (N_20113,N_19987,N_19417);
and U20114 (N_20114,N_19538,N_19576);
nor U20115 (N_20115,N_19574,N_19579);
or U20116 (N_20116,N_19557,N_19656);
nor U20117 (N_20117,N_19505,N_19518);
nor U20118 (N_20118,N_19807,N_19394);
or U20119 (N_20119,N_19776,N_19633);
nand U20120 (N_20120,N_19608,N_19799);
xnor U20121 (N_20121,N_19903,N_19599);
nor U20122 (N_20122,N_19931,N_19537);
or U20123 (N_20123,N_19685,N_19869);
xnor U20124 (N_20124,N_19597,N_19915);
nor U20125 (N_20125,N_19949,N_19769);
or U20126 (N_20126,N_19737,N_19940);
nor U20127 (N_20127,N_19975,N_19554);
nand U20128 (N_20128,N_19628,N_19567);
nand U20129 (N_20129,N_19592,N_19961);
and U20130 (N_20130,N_19669,N_19495);
nor U20131 (N_20131,N_19821,N_19601);
or U20132 (N_20132,N_19593,N_19905);
nor U20133 (N_20133,N_19440,N_19629);
or U20134 (N_20134,N_19800,N_19992);
or U20135 (N_20135,N_19577,N_19467);
nand U20136 (N_20136,N_19377,N_19668);
or U20137 (N_20137,N_19661,N_19460);
and U20138 (N_20138,N_19952,N_19950);
nor U20139 (N_20139,N_19469,N_19493);
nor U20140 (N_20140,N_19690,N_19398);
and U20141 (N_20141,N_19736,N_19848);
nand U20142 (N_20142,N_19532,N_19560);
and U20143 (N_20143,N_19654,N_19826);
nand U20144 (N_20144,N_19912,N_19921);
xor U20145 (N_20145,N_19431,N_19814);
xor U20146 (N_20146,N_19670,N_19384);
nor U20147 (N_20147,N_19806,N_19840);
or U20148 (N_20148,N_19824,N_19650);
and U20149 (N_20149,N_19676,N_19802);
xnor U20150 (N_20150,N_19433,N_19376);
xor U20151 (N_20151,N_19705,N_19803);
nor U20152 (N_20152,N_19750,N_19805);
nand U20153 (N_20153,N_19871,N_19990);
or U20154 (N_20154,N_19862,N_19591);
or U20155 (N_20155,N_19948,N_19575);
xnor U20156 (N_20156,N_19427,N_19546);
xor U20157 (N_20157,N_19425,N_19598);
nor U20158 (N_20158,N_19790,N_19913);
nand U20159 (N_20159,N_19446,N_19712);
xnor U20160 (N_20160,N_19755,N_19653);
or U20161 (N_20161,N_19611,N_19876);
nor U20162 (N_20162,N_19412,N_19686);
xor U20163 (N_20163,N_19390,N_19595);
xnor U20164 (N_20164,N_19786,N_19504);
nor U20165 (N_20165,N_19873,N_19588);
and U20166 (N_20166,N_19762,N_19514);
xnor U20167 (N_20167,N_19378,N_19822);
or U20168 (N_20168,N_19922,N_19691);
and U20169 (N_20169,N_19938,N_19834);
nor U20170 (N_20170,N_19542,N_19612);
xnor U20171 (N_20171,N_19811,N_19735);
xnor U20172 (N_20172,N_19969,N_19835);
or U20173 (N_20173,N_19582,N_19549);
xnor U20174 (N_20174,N_19725,N_19743);
and U20175 (N_20175,N_19774,N_19977);
nor U20176 (N_20176,N_19804,N_19808);
xnor U20177 (N_20177,N_19489,N_19480);
nand U20178 (N_20178,N_19552,N_19569);
nor U20179 (N_20179,N_19526,N_19844);
or U20180 (N_20180,N_19638,N_19813);
and U20181 (N_20181,N_19778,N_19954);
and U20182 (N_20182,N_19614,N_19684);
xnor U20183 (N_20183,N_19430,N_19410);
nand U20184 (N_20184,N_19420,N_19540);
and U20185 (N_20185,N_19917,N_19864);
or U20186 (N_20186,N_19519,N_19746);
nand U20187 (N_20187,N_19882,N_19476);
nand U20188 (N_20188,N_19447,N_19810);
and U20189 (N_20189,N_19827,N_19697);
or U20190 (N_20190,N_19916,N_19854);
nor U20191 (N_20191,N_19939,N_19408);
xnor U20192 (N_20192,N_19911,N_19456);
xor U20193 (N_20193,N_19520,N_19850);
xor U20194 (N_20194,N_19918,N_19496);
xnor U20195 (N_20195,N_19765,N_19525);
or U20196 (N_20196,N_19926,N_19455);
or U20197 (N_20197,N_19534,N_19500);
or U20198 (N_20198,N_19698,N_19892);
nand U20199 (N_20199,N_19868,N_19491);
or U20200 (N_20200,N_19754,N_19535);
xnor U20201 (N_20201,N_19993,N_19995);
nand U20202 (N_20202,N_19941,N_19620);
or U20203 (N_20203,N_19678,N_19908);
nor U20204 (N_20204,N_19852,N_19680);
nand U20205 (N_20205,N_19511,N_19465);
and U20206 (N_20206,N_19618,N_19730);
nor U20207 (N_20207,N_19393,N_19659);
or U20208 (N_20208,N_19714,N_19449);
or U20209 (N_20209,N_19600,N_19884);
nand U20210 (N_20210,N_19462,N_19559);
nand U20211 (N_20211,N_19617,N_19677);
nand U20212 (N_20212,N_19978,N_19760);
xor U20213 (N_20213,N_19971,N_19708);
or U20214 (N_20214,N_19589,N_19453);
or U20215 (N_20215,N_19757,N_19784);
and U20216 (N_20216,N_19407,N_19662);
xnor U20217 (N_20217,N_19843,N_19432);
or U20218 (N_20218,N_19809,N_19798);
nor U20219 (N_20219,N_19610,N_19415);
and U20220 (N_20220,N_19481,N_19761);
xnor U20221 (N_20221,N_19726,N_19464);
nor U20222 (N_20222,N_19722,N_19516);
and U20223 (N_20223,N_19718,N_19914);
nand U20224 (N_20224,N_19621,N_19936);
nor U20225 (N_20225,N_19763,N_19551);
and U20226 (N_20226,N_19994,N_19887);
nand U20227 (N_20227,N_19997,N_19477);
xnor U20228 (N_20228,N_19866,N_19490);
and U20229 (N_20229,N_19510,N_19797);
xnor U20230 (N_20230,N_19898,N_19545);
or U20231 (N_20231,N_19547,N_19663);
nand U20232 (N_20232,N_19820,N_19968);
and U20233 (N_20233,N_19506,N_19823);
or U20234 (N_20234,N_19727,N_19796);
nor U20235 (N_20235,N_19602,N_19901);
xnor U20236 (N_20236,N_19865,N_19831);
or U20237 (N_20237,N_19571,N_19508);
or U20238 (N_20238,N_19671,N_19615);
nand U20239 (N_20239,N_19474,N_19891);
or U20240 (N_20240,N_19770,N_19709);
nand U20241 (N_20241,N_19648,N_19443);
nor U20242 (N_20242,N_19719,N_19403);
xnor U20243 (N_20243,N_19603,N_19660);
xnor U20244 (N_20244,N_19988,N_19703);
nand U20245 (N_20245,N_19435,N_19818);
or U20246 (N_20246,N_19906,N_19651);
nor U20247 (N_20247,N_19857,N_19900);
and U20248 (N_20248,N_19563,N_19627);
nand U20249 (N_20249,N_19406,N_19897);
nand U20250 (N_20250,N_19502,N_19942);
nand U20251 (N_20251,N_19423,N_19581);
nor U20252 (N_20252,N_19724,N_19382);
and U20253 (N_20253,N_19533,N_19643);
or U20254 (N_20254,N_19679,N_19647);
nor U20255 (N_20255,N_19875,N_19387);
or U20256 (N_20256,N_19486,N_19619);
nor U20257 (N_20257,N_19983,N_19472);
nor U20258 (N_20258,N_19943,N_19932);
nor U20259 (N_20259,N_19402,N_19965);
and U20260 (N_20260,N_19513,N_19667);
or U20261 (N_20261,N_19448,N_19479);
and U20262 (N_20262,N_19860,N_19487);
or U20263 (N_20263,N_19955,N_19707);
nor U20264 (N_20264,N_19630,N_19883);
nor U20265 (N_20265,N_19930,N_19562);
nand U20266 (N_20266,N_19728,N_19979);
nand U20267 (N_20267,N_19473,N_19609);
nand U20268 (N_20268,N_19483,N_19482);
or U20269 (N_20269,N_19851,N_19636);
nand U20270 (N_20270,N_19904,N_19706);
xor U20271 (N_20271,N_19388,N_19785);
and U20272 (N_20272,N_19734,N_19401);
nor U20273 (N_20273,N_19846,N_19741);
and U20274 (N_20274,N_19607,N_19681);
nand U20275 (N_20275,N_19613,N_19478);
xor U20276 (N_20276,N_19492,N_19583);
or U20277 (N_20277,N_19640,N_19775);
xnor U20278 (N_20278,N_19920,N_19688);
nor U20279 (N_20279,N_19829,N_19963);
or U20280 (N_20280,N_19436,N_19704);
nor U20281 (N_20281,N_19413,N_19385);
or U20282 (N_20282,N_19584,N_19383);
and U20283 (N_20283,N_19819,N_19935);
nand U20284 (N_20284,N_19899,N_19604);
xnor U20285 (N_20285,N_19470,N_19858);
nor U20286 (N_20286,N_19646,N_19738);
nand U20287 (N_20287,N_19568,N_19910);
xor U20288 (N_20288,N_19517,N_19632);
xor U20289 (N_20289,N_19825,N_19962);
xnor U20290 (N_20290,N_19405,N_19991);
nor U20291 (N_20291,N_19665,N_19379);
nand U20292 (N_20292,N_19972,N_19484);
xor U20293 (N_20293,N_19788,N_19748);
nand U20294 (N_20294,N_19896,N_19550);
and U20295 (N_20295,N_19429,N_19945);
nand U20296 (N_20296,N_19421,N_19700);
or U20297 (N_20297,N_19441,N_19424);
xor U20298 (N_20298,N_19780,N_19764);
and U20299 (N_20299,N_19717,N_19596);
and U20300 (N_20300,N_19958,N_19815);
nor U20301 (N_20301,N_19439,N_19658);
nand U20302 (N_20302,N_19877,N_19594);
or U20303 (N_20303,N_19666,N_19530);
xor U20304 (N_20304,N_19438,N_19461);
or U20305 (N_20305,N_19573,N_19664);
xnor U20306 (N_20306,N_19561,N_19773);
or U20307 (N_20307,N_19758,N_19418);
nor U20308 (N_20308,N_19692,N_19682);
xnor U20309 (N_20309,N_19721,N_19751);
or U20310 (N_20310,N_19409,N_19699);
nor U20311 (N_20311,N_19503,N_19655);
or U20312 (N_20312,N_19623,N_19746);
or U20313 (N_20313,N_19902,N_19606);
xnor U20314 (N_20314,N_19737,N_19709);
and U20315 (N_20315,N_19393,N_19864);
nand U20316 (N_20316,N_19614,N_19679);
nor U20317 (N_20317,N_19795,N_19907);
nand U20318 (N_20318,N_19903,N_19945);
and U20319 (N_20319,N_19774,N_19619);
and U20320 (N_20320,N_19746,N_19592);
nor U20321 (N_20321,N_19585,N_19626);
nand U20322 (N_20322,N_19606,N_19958);
nand U20323 (N_20323,N_19915,N_19415);
nand U20324 (N_20324,N_19865,N_19545);
or U20325 (N_20325,N_19544,N_19715);
nand U20326 (N_20326,N_19517,N_19549);
or U20327 (N_20327,N_19694,N_19605);
xnor U20328 (N_20328,N_19947,N_19873);
nor U20329 (N_20329,N_19379,N_19568);
or U20330 (N_20330,N_19891,N_19477);
and U20331 (N_20331,N_19778,N_19390);
and U20332 (N_20332,N_19707,N_19795);
nor U20333 (N_20333,N_19415,N_19560);
and U20334 (N_20334,N_19401,N_19837);
or U20335 (N_20335,N_19553,N_19634);
xor U20336 (N_20336,N_19981,N_19924);
xor U20337 (N_20337,N_19380,N_19738);
nor U20338 (N_20338,N_19901,N_19789);
xnor U20339 (N_20339,N_19525,N_19993);
nand U20340 (N_20340,N_19391,N_19920);
nand U20341 (N_20341,N_19649,N_19467);
and U20342 (N_20342,N_19711,N_19800);
xnor U20343 (N_20343,N_19554,N_19497);
xor U20344 (N_20344,N_19449,N_19765);
nand U20345 (N_20345,N_19652,N_19562);
xor U20346 (N_20346,N_19869,N_19978);
or U20347 (N_20347,N_19850,N_19598);
and U20348 (N_20348,N_19407,N_19891);
and U20349 (N_20349,N_19393,N_19828);
xnor U20350 (N_20350,N_19553,N_19513);
nand U20351 (N_20351,N_19675,N_19407);
or U20352 (N_20352,N_19607,N_19771);
or U20353 (N_20353,N_19477,N_19722);
xnor U20354 (N_20354,N_19931,N_19568);
xnor U20355 (N_20355,N_19762,N_19755);
xor U20356 (N_20356,N_19713,N_19602);
or U20357 (N_20357,N_19538,N_19678);
nand U20358 (N_20358,N_19690,N_19384);
nand U20359 (N_20359,N_19804,N_19687);
or U20360 (N_20360,N_19447,N_19700);
nand U20361 (N_20361,N_19391,N_19914);
or U20362 (N_20362,N_19517,N_19725);
xor U20363 (N_20363,N_19861,N_19615);
or U20364 (N_20364,N_19821,N_19607);
and U20365 (N_20365,N_19877,N_19646);
or U20366 (N_20366,N_19594,N_19752);
nand U20367 (N_20367,N_19870,N_19785);
xor U20368 (N_20368,N_19659,N_19480);
xnor U20369 (N_20369,N_19883,N_19390);
nand U20370 (N_20370,N_19387,N_19642);
xor U20371 (N_20371,N_19481,N_19569);
nand U20372 (N_20372,N_19666,N_19706);
nand U20373 (N_20373,N_19955,N_19928);
xor U20374 (N_20374,N_19791,N_19803);
or U20375 (N_20375,N_19874,N_19535);
or U20376 (N_20376,N_19402,N_19592);
nor U20377 (N_20377,N_19701,N_19620);
xor U20378 (N_20378,N_19746,N_19699);
xnor U20379 (N_20379,N_19839,N_19931);
nor U20380 (N_20380,N_19516,N_19904);
nand U20381 (N_20381,N_19471,N_19567);
and U20382 (N_20382,N_19895,N_19639);
xor U20383 (N_20383,N_19800,N_19827);
and U20384 (N_20384,N_19477,N_19403);
nand U20385 (N_20385,N_19747,N_19824);
nand U20386 (N_20386,N_19469,N_19999);
nand U20387 (N_20387,N_19922,N_19520);
and U20388 (N_20388,N_19881,N_19566);
and U20389 (N_20389,N_19511,N_19654);
or U20390 (N_20390,N_19870,N_19832);
and U20391 (N_20391,N_19388,N_19857);
or U20392 (N_20392,N_19633,N_19848);
nand U20393 (N_20393,N_19532,N_19397);
or U20394 (N_20394,N_19875,N_19619);
nand U20395 (N_20395,N_19755,N_19840);
nor U20396 (N_20396,N_19793,N_19704);
and U20397 (N_20397,N_19500,N_19473);
nor U20398 (N_20398,N_19922,N_19854);
nand U20399 (N_20399,N_19714,N_19993);
and U20400 (N_20400,N_19686,N_19731);
and U20401 (N_20401,N_19472,N_19810);
nand U20402 (N_20402,N_19903,N_19449);
or U20403 (N_20403,N_19555,N_19581);
and U20404 (N_20404,N_19616,N_19732);
nand U20405 (N_20405,N_19521,N_19947);
nor U20406 (N_20406,N_19446,N_19407);
nand U20407 (N_20407,N_19848,N_19755);
and U20408 (N_20408,N_19916,N_19973);
nor U20409 (N_20409,N_19819,N_19411);
nor U20410 (N_20410,N_19989,N_19489);
xor U20411 (N_20411,N_19498,N_19801);
xor U20412 (N_20412,N_19584,N_19947);
or U20413 (N_20413,N_19413,N_19751);
and U20414 (N_20414,N_19569,N_19841);
and U20415 (N_20415,N_19827,N_19704);
xor U20416 (N_20416,N_19416,N_19736);
nor U20417 (N_20417,N_19582,N_19579);
nand U20418 (N_20418,N_19630,N_19488);
nor U20419 (N_20419,N_19867,N_19643);
xor U20420 (N_20420,N_19768,N_19845);
and U20421 (N_20421,N_19937,N_19573);
nor U20422 (N_20422,N_19726,N_19943);
and U20423 (N_20423,N_19810,N_19785);
or U20424 (N_20424,N_19757,N_19681);
or U20425 (N_20425,N_19896,N_19824);
or U20426 (N_20426,N_19902,N_19888);
and U20427 (N_20427,N_19563,N_19928);
xor U20428 (N_20428,N_19547,N_19863);
and U20429 (N_20429,N_19866,N_19826);
nor U20430 (N_20430,N_19911,N_19766);
and U20431 (N_20431,N_19505,N_19803);
or U20432 (N_20432,N_19402,N_19808);
xnor U20433 (N_20433,N_19803,N_19531);
and U20434 (N_20434,N_19469,N_19870);
and U20435 (N_20435,N_19536,N_19527);
and U20436 (N_20436,N_19969,N_19597);
xnor U20437 (N_20437,N_19410,N_19479);
and U20438 (N_20438,N_19951,N_19744);
xnor U20439 (N_20439,N_19904,N_19391);
xnor U20440 (N_20440,N_19477,N_19815);
xnor U20441 (N_20441,N_19663,N_19582);
xnor U20442 (N_20442,N_19442,N_19526);
xor U20443 (N_20443,N_19439,N_19710);
nor U20444 (N_20444,N_19563,N_19888);
nand U20445 (N_20445,N_19540,N_19729);
and U20446 (N_20446,N_19749,N_19812);
or U20447 (N_20447,N_19985,N_19548);
and U20448 (N_20448,N_19701,N_19763);
or U20449 (N_20449,N_19676,N_19928);
xnor U20450 (N_20450,N_19717,N_19563);
xnor U20451 (N_20451,N_19912,N_19498);
or U20452 (N_20452,N_19768,N_19667);
or U20453 (N_20453,N_19564,N_19681);
nand U20454 (N_20454,N_19510,N_19646);
xor U20455 (N_20455,N_19751,N_19397);
or U20456 (N_20456,N_19495,N_19770);
nand U20457 (N_20457,N_19624,N_19941);
nor U20458 (N_20458,N_19476,N_19407);
nand U20459 (N_20459,N_19838,N_19697);
xor U20460 (N_20460,N_19842,N_19421);
xor U20461 (N_20461,N_19864,N_19663);
and U20462 (N_20462,N_19419,N_19727);
or U20463 (N_20463,N_19683,N_19573);
nor U20464 (N_20464,N_19430,N_19774);
nor U20465 (N_20465,N_19905,N_19540);
or U20466 (N_20466,N_19654,N_19424);
or U20467 (N_20467,N_19953,N_19430);
and U20468 (N_20468,N_19958,N_19670);
nand U20469 (N_20469,N_19762,N_19768);
and U20470 (N_20470,N_19390,N_19986);
nand U20471 (N_20471,N_19619,N_19869);
or U20472 (N_20472,N_19871,N_19379);
nand U20473 (N_20473,N_19922,N_19562);
nor U20474 (N_20474,N_19652,N_19561);
xnor U20475 (N_20475,N_19758,N_19985);
or U20476 (N_20476,N_19815,N_19502);
and U20477 (N_20477,N_19383,N_19921);
and U20478 (N_20478,N_19492,N_19458);
xor U20479 (N_20479,N_19703,N_19456);
or U20480 (N_20480,N_19449,N_19528);
and U20481 (N_20481,N_19773,N_19641);
and U20482 (N_20482,N_19871,N_19680);
nand U20483 (N_20483,N_19480,N_19721);
nand U20484 (N_20484,N_19847,N_19514);
nand U20485 (N_20485,N_19795,N_19614);
nor U20486 (N_20486,N_19818,N_19731);
xor U20487 (N_20487,N_19515,N_19992);
nor U20488 (N_20488,N_19557,N_19404);
and U20489 (N_20489,N_19861,N_19501);
nor U20490 (N_20490,N_19385,N_19414);
or U20491 (N_20491,N_19564,N_19914);
and U20492 (N_20492,N_19802,N_19533);
xnor U20493 (N_20493,N_19727,N_19827);
nand U20494 (N_20494,N_19743,N_19666);
or U20495 (N_20495,N_19555,N_19434);
nand U20496 (N_20496,N_19976,N_19567);
or U20497 (N_20497,N_19387,N_19771);
nor U20498 (N_20498,N_19533,N_19916);
or U20499 (N_20499,N_19394,N_19522);
nand U20500 (N_20500,N_19744,N_19749);
or U20501 (N_20501,N_19501,N_19789);
and U20502 (N_20502,N_19601,N_19404);
nand U20503 (N_20503,N_19496,N_19624);
and U20504 (N_20504,N_19949,N_19517);
nand U20505 (N_20505,N_19595,N_19627);
nor U20506 (N_20506,N_19690,N_19387);
nand U20507 (N_20507,N_19532,N_19753);
or U20508 (N_20508,N_19740,N_19819);
nand U20509 (N_20509,N_19495,N_19794);
xnor U20510 (N_20510,N_19419,N_19476);
and U20511 (N_20511,N_19765,N_19615);
and U20512 (N_20512,N_19602,N_19617);
and U20513 (N_20513,N_19476,N_19980);
nor U20514 (N_20514,N_19487,N_19575);
xnor U20515 (N_20515,N_19470,N_19575);
nor U20516 (N_20516,N_19637,N_19516);
nand U20517 (N_20517,N_19578,N_19949);
or U20518 (N_20518,N_19482,N_19939);
nor U20519 (N_20519,N_19499,N_19874);
nand U20520 (N_20520,N_19488,N_19642);
nor U20521 (N_20521,N_19880,N_19375);
nor U20522 (N_20522,N_19899,N_19742);
nor U20523 (N_20523,N_19921,N_19970);
or U20524 (N_20524,N_19606,N_19974);
xnor U20525 (N_20525,N_19596,N_19386);
xnor U20526 (N_20526,N_19775,N_19784);
xnor U20527 (N_20527,N_19845,N_19571);
and U20528 (N_20528,N_19910,N_19415);
or U20529 (N_20529,N_19626,N_19508);
and U20530 (N_20530,N_19527,N_19509);
xnor U20531 (N_20531,N_19502,N_19425);
and U20532 (N_20532,N_19609,N_19918);
nand U20533 (N_20533,N_19946,N_19428);
nor U20534 (N_20534,N_19580,N_19520);
xor U20535 (N_20535,N_19612,N_19510);
xor U20536 (N_20536,N_19961,N_19385);
nand U20537 (N_20537,N_19942,N_19604);
and U20538 (N_20538,N_19762,N_19509);
nand U20539 (N_20539,N_19994,N_19750);
nand U20540 (N_20540,N_19864,N_19816);
nand U20541 (N_20541,N_19870,N_19866);
xnor U20542 (N_20542,N_19397,N_19549);
or U20543 (N_20543,N_19996,N_19802);
nand U20544 (N_20544,N_19482,N_19936);
nor U20545 (N_20545,N_19994,N_19433);
and U20546 (N_20546,N_19659,N_19567);
nand U20547 (N_20547,N_19615,N_19914);
xor U20548 (N_20548,N_19691,N_19451);
and U20549 (N_20549,N_19668,N_19388);
nor U20550 (N_20550,N_19565,N_19925);
or U20551 (N_20551,N_19973,N_19467);
nand U20552 (N_20552,N_19916,N_19867);
or U20553 (N_20553,N_19715,N_19914);
nand U20554 (N_20554,N_19654,N_19737);
nand U20555 (N_20555,N_19752,N_19546);
or U20556 (N_20556,N_19523,N_19961);
or U20557 (N_20557,N_19573,N_19420);
and U20558 (N_20558,N_19962,N_19651);
or U20559 (N_20559,N_19974,N_19657);
nand U20560 (N_20560,N_19986,N_19782);
nor U20561 (N_20561,N_19905,N_19509);
nand U20562 (N_20562,N_19971,N_19620);
nand U20563 (N_20563,N_19706,N_19874);
nor U20564 (N_20564,N_19931,N_19587);
nor U20565 (N_20565,N_19882,N_19810);
nand U20566 (N_20566,N_19649,N_19819);
nor U20567 (N_20567,N_19725,N_19797);
nand U20568 (N_20568,N_19694,N_19894);
xnor U20569 (N_20569,N_19776,N_19660);
nand U20570 (N_20570,N_19774,N_19662);
or U20571 (N_20571,N_19793,N_19719);
xor U20572 (N_20572,N_19389,N_19918);
nand U20573 (N_20573,N_19467,N_19717);
nand U20574 (N_20574,N_19659,N_19813);
and U20575 (N_20575,N_19546,N_19767);
and U20576 (N_20576,N_19765,N_19855);
and U20577 (N_20577,N_19969,N_19844);
or U20578 (N_20578,N_19690,N_19842);
nor U20579 (N_20579,N_19686,N_19571);
xor U20580 (N_20580,N_19859,N_19634);
nand U20581 (N_20581,N_19915,N_19649);
nor U20582 (N_20582,N_19392,N_19430);
xor U20583 (N_20583,N_19661,N_19813);
xor U20584 (N_20584,N_19841,N_19906);
nand U20585 (N_20585,N_19673,N_19860);
nor U20586 (N_20586,N_19704,N_19798);
nor U20587 (N_20587,N_19927,N_19876);
or U20588 (N_20588,N_19654,N_19506);
nand U20589 (N_20589,N_19656,N_19779);
or U20590 (N_20590,N_19705,N_19753);
or U20591 (N_20591,N_19833,N_19498);
or U20592 (N_20592,N_19551,N_19492);
nor U20593 (N_20593,N_19930,N_19552);
xnor U20594 (N_20594,N_19497,N_19931);
and U20595 (N_20595,N_19669,N_19610);
nor U20596 (N_20596,N_19648,N_19500);
xor U20597 (N_20597,N_19864,N_19762);
nand U20598 (N_20598,N_19831,N_19778);
nor U20599 (N_20599,N_19891,N_19659);
and U20600 (N_20600,N_19810,N_19874);
nor U20601 (N_20601,N_19536,N_19480);
xor U20602 (N_20602,N_19930,N_19595);
nand U20603 (N_20603,N_19739,N_19945);
and U20604 (N_20604,N_19912,N_19540);
xor U20605 (N_20605,N_19449,N_19503);
nand U20606 (N_20606,N_19619,N_19908);
nor U20607 (N_20607,N_19699,N_19766);
or U20608 (N_20608,N_19792,N_19919);
or U20609 (N_20609,N_19608,N_19864);
or U20610 (N_20610,N_19594,N_19510);
nand U20611 (N_20611,N_19899,N_19854);
xor U20612 (N_20612,N_19436,N_19634);
xnor U20613 (N_20613,N_19897,N_19973);
and U20614 (N_20614,N_19609,N_19448);
xor U20615 (N_20615,N_19831,N_19539);
or U20616 (N_20616,N_19388,N_19606);
or U20617 (N_20617,N_19796,N_19613);
and U20618 (N_20618,N_19728,N_19887);
and U20619 (N_20619,N_19626,N_19419);
or U20620 (N_20620,N_19834,N_19455);
xnor U20621 (N_20621,N_19569,N_19881);
or U20622 (N_20622,N_19596,N_19870);
xnor U20623 (N_20623,N_19479,N_19519);
and U20624 (N_20624,N_19958,N_19960);
and U20625 (N_20625,N_20317,N_20293);
xnor U20626 (N_20626,N_20273,N_20426);
or U20627 (N_20627,N_20479,N_20063);
nand U20628 (N_20628,N_20603,N_20262);
or U20629 (N_20629,N_20578,N_20309);
xnor U20630 (N_20630,N_20566,N_20192);
or U20631 (N_20631,N_20606,N_20605);
or U20632 (N_20632,N_20441,N_20181);
xor U20633 (N_20633,N_20624,N_20581);
and U20634 (N_20634,N_20058,N_20199);
nand U20635 (N_20635,N_20448,N_20536);
nor U20636 (N_20636,N_20220,N_20380);
nand U20637 (N_20637,N_20543,N_20169);
nor U20638 (N_20638,N_20240,N_20583);
xor U20639 (N_20639,N_20195,N_20138);
xor U20640 (N_20640,N_20517,N_20456);
xnor U20641 (N_20641,N_20412,N_20491);
and U20642 (N_20642,N_20197,N_20164);
or U20643 (N_20643,N_20613,N_20446);
nand U20644 (N_20644,N_20304,N_20533);
nor U20645 (N_20645,N_20361,N_20442);
or U20646 (N_20646,N_20364,N_20184);
nand U20647 (N_20647,N_20486,N_20104);
and U20648 (N_20648,N_20525,N_20359);
or U20649 (N_20649,N_20400,N_20302);
or U20650 (N_20650,N_20529,N_20259);
nand U20651 (N_20651,N_20389,N_20383);
and U20652 (N_20652,N_20424,N_20026);
xnor U20653 (N_20653,N_20055,N_20590);
nor U20654 (N_20654,N_20177,N_20205);
or U20655 (N_20655,N_20072,N_20222);
or U20656 (N_20656,N_20241,N_20315);
xnor U20657 (N_20657,N_20621,N_20268);
xnor U20658 (N_20658,N_20478,N_20593);
nand U20659 (N_20659,N_20041,N_20530);
xnor U20660 (N_20660,N_20167,N_20194);
nor U20661 (N_20661,N_20556,N_20498);
xnor U20662 (N_20662,N_20013,N_20191);
and U20663 (N_20663,N_20172,N_20185);
and U20664 (N_20664,N_20298,N_20406);
and U20665 (N_20665,N_20054,N_20272);
or U20666 (N_20666,N_20126,N_20562);
or U20667 (N_20667,N_20559,N_20497);
nor U20668 (N_20668,N_20086,N_20170);
nor U20669 (N_20669,N_20074,N_20457);
xnor U20670 (N_20670,N_20029,N_20413);
nand U20671 (N_20671,N_20065,N_20001);
nor U20672 (N_20672,N_20504,N_20542);
and U20673 (N_20673,N_20596,N_20320);
and U20674 (N_20674,N_20440,N_20186);
xor U20675 (N_20675,N_20057,N_20375);
or U20676 (N_20676,N_20474,N_20467);
and U20677 (N_20677,N_20119,N_20537);
nor U20678 (N_20678,N_20544,N_20291);
xor U20679 (N_20679,N_20116,N_20101);
nor U20680 (N_20680,N_20419,N_20196);
nor U20681 (N_20681,N_20469,N_20601);
nor U20682 (N_20682,N_20278,N_20096);
nor U20683 (N_20683,N_20373,N_20303);
xor U20684 (N_20684,N_20025,N_20264);
or U20685 (N_20685,N_20352,N_20234);
xor U20686 (N_20686,N_20447,N_20430);
or U20687 (N_20687,N_20095,N_20108);
xnor U20688 (N_20688,N_20127,N_20082);
nor U20689 (N_20689,N_20396,N_20214);
or U20690 (N_20690,N_20425,N_20168);
nor U20691 (N_20691,N_20011,N_20161);
or U20692 (N_20692,N_20511,N_20592);
nand U20693 (N_20693,N_20023,N_20397);
nand U20694 (N_20694,N_20554,N_20573);
nand U20695 (N_20695,N_20120,N_20618);
nand U20696 (N_20696,N_20549,N_20114);
nor U20697 (N_20697,N_20137,N_20337);
nand U20698 (N_20698,N_20156,N_20575);
nand U20699 (N_20699,N_20421,N_20134);
and U20700 (N_20700,N_20338,N_20062);
xor U20701 (N_20701,N_20034,N_20374);
xnor U20702 (N_20702,N_20051,N_20102);
and U20703 (N_20703,N_20064,N_20030);
nand U20704 (N_20704,N_20093,N_20180);
or U20705 (N_20705,N_20388,N_20219);
or U20706 (N_20706,N_20476,N_20382);
nor U20707 (N_20707,N_20094,N_20407);
and U20708 (N_20708,N_20007,N_20404);
nor U20709 (N_20709,N_20551,N_20092);
xor U20710 (N_20710,N_20574,N_20558);
and U20711 (N_20711,N_20144,N_20132);
nand U20712 (N_20712,N_20066,N_20341);
nor U20713 (N_20713,N_20089,N_20468);
and U20714 (N_20714,N_20021,N_20279);
or U20715 (N_20715,N_20059,N_20330);
xor U20716 (N_20716,N_20378,N_20349);
or U20717 (N_20717,N_20067,N_20075);
and U20718 (N_20718,N_20410,N_20472);
and U20719 (N_20719,N_20294,N_20557);
nand U20720 (N_20720,N_20282,N_20595);
nor U20721 (N_20721,N_20078,N_20500);
or U20722 (N_20722,N_20107,N_20157);
or U20723 (N_20723,N_20516,N_20518);
nor U20724 (N_20724,N_20515,N_20376);
nand U20725 (N_20725,N_20141,N_20236);
or U20726 (N_20726,N_20610,N_20598);
nand U20727 (N_20727,N_20117,N_20328);
nor U20728 (N_20728,N_20193,N_20182);
and U20729 (N_20729,N_20130,N_20512);
nor U20730 (N_20730,N_20466,N_20582);
or U20731 (N_20731,N_20552,N_20296);
xor U20732 (N_20732,N_20343,N_20122);
nand U20733 (N_20733,N_20276,N_20189);
xor U20734 (N_20734,N_20564,N_20420);
or U20735 (N_20735,N_20316,N_20586);
or U20736 (N_20736,N_20414,N_20048);
nor U20737 (N_20737,N_20149,N_20019);
xor U20738 (N_20738,N_20534,N_20002);
and U20739 (N_20739,N_20571,N_20381);
and U20740 (N_20740,N_20232,N_20434);
nand U20741 (N_20741,N_20079,N_20403);
xor U20742 (N_20742,N_20335,N_20576);
nor U20743 (N_20743,N_20611,N_20427);
nand U20744 (N_20744,N_20190,N_20523);
and U20745 (N_20745,N_20269,N_20162);
nor U20746 (N_20746,N_20555,N_20198);
and U20747 (N_20747,N_20077,N_20379);
nand U20748 (N_20748,N_20047,N_20188);
or U20749 (N_20749,N_20433,N_20550);
nor U20750 (N_20750,N_20546,N_20115);
xnor U20751 (N_20751,N_20024,N_20033);
nor U20752 (N_20752,N_20401,N_20422);
and U20753 (N_20753,N_20267,N_20501);
or U20754 (N_20754,N_20052,N_20437);
nor U20755 (N_20755,N_20154,N_20612);
xnor U20756 (N_20756,N_20076,N_20588);
nor U20757 (N_20757,N_20431,N_20284);
or U20758 (N_20758,N_20449,N_20111);
nand U20759 (N_20759,N_20208,N_20443);
nor U20760 (N_20760,N_20288,N_20247);
nor U20761 (N_20761,N_20570,N_20087);
xor U20762 (N_20762,N_20372,N_20020);
and U20763 (N_20763,N_20031,N_20258);
and U20764 (N_20764,N_20540,N_20508);
nand U20765 (N_20765,N_20455,N_20106);
or U20766 (N_20766,N_20461,N_20333);
xor U20767 (N_20767,N_20251,N_20158);
or U20768 (N_20768,N_20432,N_20027);
nor U20769 (N_20769,N_20535,N_20473);
nand U20770 (N_20770,N_20602,N_20248);
or U20771 (N_20771,N_20580,N_20323);
or U20772 (N_20772,N_20069,N_20332);
xnor U20773 (N_20773,N_20460,N_20049);
nor U20774 (N_20774,N_20140,N_20287);
or U20775 (N_20775,N_20006,N_20538);
or U20776 (N_20776,N_20070,N_20056);
xor U20777 (N_20777,N_20520,N_20398);
or U20778 (N_20778,N_20040,N_20622);
xnor U20779 (N_20779,N_20166,N_20326);
or U20780 (N_20780,N_20308,N_20037);
nor U20781 (N_20781,N_20113,N_20297);
or U20782 (N_20782,N_20017,N_20289);
and U20783 (N_20783,N_20014,N_20039);
xor U20784 (N_20784,N_20483,N_20444);
or U20785 (N_20785,N_20405,N_20475);
nor U20786 (N_20786,N_20274,N_20100);
and U20787 (N_20787,N_20271,N_20159);
or U20788 (N_20788,N_20081,N_20452);
and U20789 (N_20789,N_20213,N_20435);
nor U20790 (N_20790,N_20152,N_20585);
nor U20791 (N_20791,N_20347,N_20480);
xor U20792 (N_20792,N_20139,N_20165);
or U20793 (N_20793,N_20045,N_20035);
nand U20794 (N_20794,N_20459,N_20324);
or U20795 (N_20795,N_20136,N_20354);
nor U20796 (N_20796,N_20489,N_20155);
nor U20797 (N_20797,N_20123,N_20385);
xor U20798 (N_20798,N_20371,N_20173);
or U20799 (N_20799,N_20229,N_20547);
and U20800 (N_20800,N_20509,N_20228);
or U20801 (N_20801,N_20344,N_20362);
and U20802 (N_20802,N_20356,N_20176);
or U20803 (N_20803,N_20519,N_20569);
nand U20804 (N_20804,N_20608,N_20567);
nor U20805 (N_20805,N_20129,N_20250);
and U20806 (N_20806,N_20242,N_20615);
nor U20807 (N_20807,N_20524,N_20607);
nor U20808 (N_20808,N_20125,N_20060);
xnor U20809 (N_20809,N_20098,N_20178);
and U20810 (N_20810,N_20390,N_20015);
or U20811 (N_20811,N_20620,N_20312);
and U20812 (N_20812,N_20409,N_20563);
xor U20813 (N_20813,N_20490,N_20348);
nand U20814 (N_20814,N_20256,N_20143);
or U20815 (N_20815,N_20481,N_20553);
xnor U20816 (N_20816,N_20285,N_20392);
or U20817 (N_20817,N_20128,N_20541);
and U20818 (N_20818,N_20604,N_20526);
and U20819 (N_20819,N_20280,N_20445);
or U20820 (N_20820,N_20391,N_20522);
or U20821 (N_20821,N_20150,N_20206);
and U20822 (N_20822,N_20204,N_20277);
and U20823 (N_20823,N_20350,N_20616);
nand U20824 (N_20824,N_20623,N_20145);
xor U20825 (N_20825,N_20153,N_20022);
or U20826 (N_20826,N_20151,N_20210);
or U20827 (N_20827,N_20417,N_20450);
nand U20828 (N_20828,N_20216,N_20253);
nand U20829 (N_20829,N_20009,N_20503);
nand U20830 (N_20830,N_20463,N_20233);
nand U20831 (N_20831,N_20411,N_20482);
or U20832 (N_20832,N_20261,N_20163);
nor U20833 (N_20833,N_20046,N_20451);
or U20834 (N_20834,N_20103,N_20209);
or U20835 (N_20835,N_20387,N_20485);
nand U20836 (N_20836,N_20532,N_20314);
nand U20837 (N_20837,N_20471,N_20599);
xor U20838 (N_20838,N_20146,N_20345);
nand U20839 (N_20839,N_20200,N_20299);
nor U20840 (N_20840,N_20275,N_20281);
and U20841 (N_20841,N_20004,N_20311);
and U20842 (N_20842,N_20353,N_20148);
and U20843 (N_20843,N_20318,N_20321);
nand U20844 (N_20844,N_20028,N_20121);
xnor U20845 (N_20845,N_20370,N_20357);
and U20846 (N_20846,N_20589,N_20230);
and U20847 (N_20847,N_20044,N_20408);
nand U20848 (N_20848,N_20591,N_20428);
xnor U20849 (N_20849,N_20218,N_20458);
and U20850 (N_20850,N_20005,N_20331);
or U20851 (N_20851,N_20239,N_20394);
and U20852 (N_20852,N_20179,N_20513);
nand U20853 (N_20853,N_20355,N_20010);
xor U20854 (N_20854,N_20085,N_20249);
nand U20855 (N_20855,N_20212,N_20000);
or U20856 (N_20856,N_20470,N_20322);
xnor U20857 (N_20857,N_20091,N_20496);
nor U20858 (N_20858,N_20099,N_20012);
nor U20859 (N_20859,N_20484,N_20568);
nand U20860 (N_20860,N_20584,N_20477);
nand U20861 (N_20861,N_20386,N_20502);
nor U20862 (N_20862,N_20528,N_20109);
nand U20863 (N_20863,N_20142,N_20243);
xnor U20864 (N_20864,N_20393,N_20307);
or U20865 (N_20865,N_20226,N_20487);
nor U20866 (N_20866,N_20488,N_20237);
nand U20867 (N_20867,N_20300,N_20083);
nand U20868 (N_20868,N_20325,N_20292);
nand U20869 (N_20869,N_20263,N_20061);
and U20870 (N_20870,N_20118,N_20018);
nand U20871 (N_20871,N_20224,N_20254);
nor U20872 (N_20872,N_20171,N_20495);
and U20873 (N_20873,N_20211,N_20436);
nand U20874 (N_20874,N_20016,N_20053);
nand U20875 (N_20875,N_20160,N_20560);
nand U20876 (N_20876,N_20175,N_20244);
and U20877 (N_20877,N_20071,N_20358);
or U20878 (N_20878,N_20295,N_20365);
and U20879 (N_20879,N_20223,N_20133);
and U20880 (N_20880,N_20453,N_20003);
xor U20881 (N_20881,N_20238,N_20465);
nor U20882 (N_20882,N_20423,N_20201);
and U20883 (N_20883,N_20462,N_20346);
and U20884 (N_20884,N_20492,N_20565);
nor U20885 (N_20885,N_20245,N_20493);
nor U20886 (N_20886,N_20494,N_20454);
nand U20887 (N_20887,N_20609,N_20231);
nand U20888 (N_20888,N_20217,N_20531);
nand U20889 (N_20889,N_20418,N_20614);
xor U20890 (N_20890,N_20283,N_20183);
xor U20891 (N_20891,N_20579,N_20438);
and U20892 (N_20892,N_20577,N_20131);
and U20893 (N_20893,N_20395,N_20510);
or U20894 (N_20894,N_20306,N_20305);
nand U20895 (N_20895,N_20050,N_20545);
nor U20896 (N_20896,N_20360,N_20548);
xnor U20897 (N_20897,N_20600,N_20561);
or U20898 (N_20898,N_20594,N_20084);
nor U20899 (N_20899,N_20068,N_20363);
nand U20900 (N_20900,N_20110,N_20038);
or U20901 (N_20901,N_20135,N_20339);
xor U20902 (N_20902,N_20439,N_20416);
xnor U20903 (N_20903,N_20260,N_20507);
xor U20904 (N_20904,N_20527,N_20539);
xnor U20905 (N_20905,N_20225,N_20246);
nor U20906 (N_20906,N_20080,N_20334);
xor U20907 (N_20907,N_20402,N_20310);
nor U20908 (N_20908,N_20257,N_20215);
xor U20909 (N_20909,N_20266,N_20174);
nor U20910 (N_20910,N_20032,N_20366);
or U20911 (N_20911,N_20572,N_20270);
and U20912 (N_20912,N_20255,N_20368);
nand U20913 (N_20913,N_20384,N_20342);
xnor U20914 (N_20914,N_20351,N_20290);
nor U20915 (N_20915,N_20203,N_20505);
and U20916 (N_20916,N_20301,N_20008);
and U20917 (N_20917,N_20235,N_20327);
nand U20918 (N_20918,N_20521,N_20036);
or U20919 (N_20919,N_20252,N_20090);
and U20920 (N_20920,N_20415,N_20313);
or U20921 (N_20921,N_20202,N_20597);
or U20922 (N_20922,N_20429,N_20336);
or U20923 (N_20923,N_20042,N_20187);
xor U20924 (N_20924,N_20506,N_20043);
or U20925 (N_20925,N_20587,N_20464);
nand U20926 (N_20926,N_20097,N_20367);
and U20927 (N_20927,N_20105,N_20227);
nor U20928 (N_20928,N_20619,N_20369);
or U20929 (N_20929,N_20073,N_20221);
or U20930 (N_20930,N_20207,N_20124);
nand U20931 (N_20931,N_20514,N_20329);
nor U20932 (N_20932,N_20147,N_20377);
nor U20933 (N_20933,N_20286,N_20088);
nor U20934 (N_20934,N_20112,N_20319);
or U20935 (N_20935,N_20399,N_20340);
or U20936 (N_20936,N_20499,N_20265);
xor U20937 (N_20937,N_20617,N_20132);
or U20938 (N_20938,N_20304,N_20559);
nor U20939 (N_20939,N_20293,N_20472);
or U20940 (N_20940,N_20591,N_20376);
xnor U20941 (N_20941,N_20551,N_20460);
and U20942 (N_20942,N_20021,N_20473);
and U20943 (N_20943,N_20445,N_20036);
xnor U20944 (N_20944,N_20331,N_20603);
nand U20945 (N_20945,N_20033,N_20582);
nor U20946 (N_20946,N_20534,N_20522);
nor U20947 (N_20947,N_20258,N_20491);
or U20948 (N_20948,N_20591,N_20382);
nand U20949 (N_20949,N_20231,N_20472);
xor U20950 (N_20950,N_20427,N_20090);
and U20951 (N_20951,N_20605,N_20236);
nand U20952 (N_20952,N_20192,N_20502);
or U20953 (N_20953,N_20232,N_20066);
nor U20954 (N_20954,N_20536,N_20328);
nor U20955 (N_20955,N_20542,N_20318);
nand U20956 (N_20956,N_20294,N_20224);
and U20957 (N_20957,N_20050,N_20475);
nor U20958 (N_20958,N_20065,N_20175);
and U20959 (N_20959,N_20434,N_20167);
xor U20960 (N_20960,N_20549,N_20066);
nand U20961 (N_20961,N_20502,N_20414);
nor U20962 (N_20962,N_20134,N_20382);
and U20963 (N_20963,N_20427,N_20573);
nor U20964 (N_20964,N_20021,N_20563);
or U20965 (N_20965,N_20180,N_20416);
or U20966 (N_20966,N_20029,N_20060);
nor U20967 (N_20967,N_20118,N_20355);
nor U20968 (N_20968,N_20387,N_20616);
xnor U20969 (N_20969,N_20303,N_20112);
xnor U20970 (N_20970,N_20393,N_20355);
nand U20971 (N_20971,N_20545,N_20616);
nor U20972 (N_20972,N_20533,N_20459);
and U20973 (N_20973,N_20565,N_20303);
xnor U20974 (N_20974,N_20086,N_20063);
xor U20975 (N_20975,N_20329,N_20558);
nand U20976 (N_20976,N_20182,N_20587);
nand U20977 (N_20977,N_20200,N_20510);
and U20978 (N_20978,N_20555,N_20115);
or U20979 (N_20979,N_20389,N_20165);
nand U20980 (N_20980,N_20019,N_20568);
nor U20981 (N_20981,N_20132,N_20414);
xor U20982 (N_20982,N_20564,N_20092);
xor U20983 (N_20983,N_20524,N_20509);
and U20984 (N_20984,N_20581,N_20140);
or U20985 (N_20985,N_20333,N_20020);
or U20986 (N_20986,N_20084,N_20288);
nor U20987 (N_20987,N_20095,N_20342);
nor U20988 (N_20988,N_20492,N_20150);
nand U20989 (N_20989,N_20362,N_20169);
nand U20990 (N_20990,N_20133,N_20013);
nor U20991 (N_20991,N_20122,N_20524);
or U20992 (N_20992,N_20035,N_20332);
or U20993 (N_20993,N_20370,N_20226);
and U20994 (N_20994,N_20158,N_20231);
nor U20995 (N_20995,N_20576,N_20402);
nor U20996 (N_20996,N_20077,N_20410);
and U20997 (N_20997,N_20228,N_20317);
xnor U20998 (N_20998,N_20070,N_20113);
nand U20999 (N_20999,N_20341,N_20503);
and U21000 (N_21000,N_20230,N_20170);
nor U21001 (N_21001,N_20046,N_20475);
xnor U21002 (N_21002,N_20135,N_20201);
nand U21003 (N_21003,N_20441,N_20419);
nor U21004 (N_21004,N_20125,N_20430);
xor U21005 (N_21005,N_20052,N_20297);
and U21006 (N_21006,N_20361,N_20149);
nand U21007 (N_21007,N_20151,N_20478);
and U21008 (N_21008,N_20054,N_20121);
nor U21009 (N_21009,N_20376,N_20121);
xor U21010 (N_21010,N_20504,N_20404);
or U21011 (N_21011,N_20092,N_20485);
nand U21012 (N_21012,N_20457,N_20558);
xor U21013 (N_21013,N_20084,N_20249);
or U21014 (N_21014,N_20559,N_20220);
or U21015 (N_21015,N_20033,N_20222);
xor U21016 (N_21016,N_20401,N_20001);
nor U21017 (N_21017,N_20168,N_20253);
nor U21018 (N_21018,N_20135,N_20073);
xnor U21019 (N_21019,N_20021,N_20312);
nand U21020 (N_21020,N_20515,N_20447);
and U21021 (N_21021,N_20552,N_20069);
nor U21022 (N_21022,N_20545,N_20128);
nand U21023 (N_21023,N_20167,N_20473);
nor U21024 (N_21024,N_20251,N_20342);
xor U21025 (N_21025,N_20459,N_20152);
and U21026 (N_21026,N_20616,N_20528);
nand U21027 (N_21027,N_20378,N_20609);
and U21028 (N_21028,N_20220,N_20574);
xor U21029 (N_21029,N_20094,N_20305);
xor U21030 (N_21030,N_20349,N_20259);
nor U21031 (N_21031,N_20488,N_20263);
and U21032 (N_21032,N_20264,N_20323);
xnor U21033 (N_21033,N_20478,N_20378);
and U21034 (N_21034,N_20530,N_20439);
or U21035 (N_21035,N_20523,N_20480);
or U21036 (N_21036,N_20358,N_20150);
and U21037 (N_21037,N_20326,N_20075);
nor U21038 (N_21038,N_20456,N_20207);
nand U21039 (N_21039,N_20255,N_20147);
nand U21040 (N_21040,N_20436,N_20520);
xor U21041 (N_21041,N_20542,N_20445);
or U21042 (N_21042,N_20128,N_20611);
nor U21043 (N_21043,N_20470,N_20432);
nand U21044 (N_21044,N_20506,N_20124);
xor U21045 (N_21045,N_20524,N_20602);
nor U21046 (N_21046,N_20499,N_20565);
xor U21047 (N_21047,N_20118,N_20579);
nand U21048 (N_21048,N_20409,N_20025);
nor U21049 (N_21049,N_20248,N_20123);
nand U21050 (N_21050,N_20189,N_20449);
or U21051 (N_21051,N_20238,N_20295);
nand U21052 (N_21052,N_20192,N_20363);
nand U21053 (N_21053,N_20063,N_20202);
nor U21054 (N_21054,N_20242,N_20624);
nand U21055 (N_21055,N_20577,N_20207);
xor U21056 (N_21056,N_20258,N_20020);
nor U21057 (N_21057,N_20411,N_20421);
xnor U21058 (N_21058,N_20389,N_20449);
nor U21059 (N_21059,N_20520,N_20111);
and U21060 (N_21060,N_20330,N_20453);
nand U21061 (N_21061,N_20527,N_20477);
and U21062 (N_21062,N_20239,N_20042);
xnor U21063 (N_21063,N_20169,N_20618);
and U21064 (N_21064,N_20479,N_20611);
nor U21065 (N_21065,N_20172,N_20453);
xnor U21066 (N_21066,N_20430,N_20037);
nand U21067 (N_21067,N_20418,N_20379);
or U21068 (N_21068,N_20569,N_20516);
or U21069 (N_21069,N_20127,N_20201);
nor U21070 (N_21070,N_20135,N_20443);
and U21071 (N_21071,N_20336,N_20351);
or U21072 (N_21072,N_20493,N_20527);
nor U21073 (N_21073,N_20126,N_20621);
nor U21074 (N_21074,N_20389,N_20603);
or U21075 (N_21075,N_20334,N_20242);
nand U21076 (N_21076,N_20444,N_20347);
nand U21077 (N_21077,N_20224,N_20475);
nand U21078 (N_21078,N_20000,N_20335);
and U21079 (N_21079,N_20353,N_20540);
or U21080 (N_21080,N_20426,N_20542);
or U21081 (N_21081,N_20217,N_20149);
nand U21082 (N_21082,N_20402,N_20317);
xor U21083 (N_21083,N_20260,N_20158);
or U21084 (N_21084,N_20167,N_20413);
nor U21085 (N_21085,N_20571,N_20032);
nor U21086 (N_21086,N_20585,N_20073);
or U21087 (N_21087,N_20622,N_20421);
nand U21088 (N_21088,N_20177,N_20470);
and U21089 (N_21089,N_20612,N_20187);
nor U21090 (N_21090,N_20133,N_20232);
nand U21091 (N_21091,N_20292,N_20564);
xor U21092 (N_21092,N_20533,N_20239);
and U21093 (N_21093,N_20466,N_20538);
xor U21094 (N_21094,N_20537,N_20496);
nand U21095 (N_21095,N_20301,N_20150);
nand U21096 (N_21096,N_20440,N_20581);
nor U21097 (N_21097,N_20264,N_20455);
nor U21098 (N_21098,N_20458,N_20564);
xor U21099 (N_21099,N_20121,N_20296);
and U21100 (N_21100,N_20583,N_20565);
nor U21101 (N_21101,N_20187,N_20221);
nor U21102 (N_21102,N_20601,N_20543);
nor U21103 (N_21103,N_20390,N_20167);
nor U21104 (N_21104,N_20307,N_20179);
and U21105 (N_21105,N_20588,N_20368);
or U21106 (N_21106,N_20378,N_20104);
xnor U21107 (N_21107,N_20531,N_20610);
nor U21108 (N_21108,N_20554,N_20131);
nand U21109 (N_21109,N_20491,N_20116);
or U21110 (N_21110,N_20208,N_20454);
and U21111 (N_21111,N_20464,N_20003);
or U21112 (N_21112,N_20204,N_20449);
or U21113 (N_21113,N_20469,N_20619);
and U21114 (N_21114,N_20606,N_20231);
nand U21115 (N_21115,N_20058,N_20230);
xor U21116 (N_21116,N_20078,N_20325);
xnor U21117 (N_21117,N_20099,N_20224);
and U21118 (N_21118,N_20473,N_20261);
or U21119 (N_21119,N_20456,N_20430);
nor U21120 (N_21120,N_20056,N_20425);
or U21121 (N_21121,N_20501,N_20402);
xnor U21122 (N_21122,N_20582,N_20429);
nor U21123 (N_21123,N_20499,N_20329);
or U21124 (N_21124,N_20236,N_20427);
nor U21125 (N_21125,N_20288,N_20545);
nand U21126 (N_21126,N_20094,N_20612);
and U21127 (N_21127,N_20075,N_20251);
and U21128 (N_21128,N_20260,N_20194);
or U21129 (N_21129,N_20496,N_20369);
nand U21130 (N_21130,N_20226,N_20293);
and U21131 (N_21131,N_20204,N_20467);
xnor U21132 (N_21132,N_20271,N_20116);
and U21133 (N_21133,N_20110,N_20232);
xor U21134 (N_21134,N_20576,N_20437);
or U21135 (N_21135,N_20136,N_20219);
and U21136 (N_21136,N_20209,N_20068);
nor U21137 (N_21137,N_20502,N_20196);
and U21138 (N_21138,N_20479,N_20245);
nor U21139 (N_21139,N_20517,N_20292);
nor U21140 (N_21140,N_20483,N_20127);
or U21141 (N_21141,N_20532,N_20493);
nor U21142 (N_21142,N_20493,N_20470);
nand U21143 (N_21143,N_20322,N_20328);
or U21144 (N_21144,N_20160,N_20460);
nor U21145 (N_21145,N_20481,N_20199);
or U21146 (N_21146,N_20307,N_20291);
xor U21147 (N_21147,N_20293,N_20352);
and U21148 (N_21148,N_20430,N_20584);
and U21149 (N_21149,N_20589,N_20499);
nor U21150 (N_21150,N_20160,N_20056);
nor U21151 (N_21151,N_20150,N_20347);
and U21152 (N_21152,N_20394,N_20428);
xor U21153 (N_21153,N_20326,N_20404);
and U21154 (N_21154,N_20299,N_20091);
xnor U21155 (N_21155,N_20168,N_20538);
nor U21156 (N_21156,N_20403,N_20597);
xor U21157 (N_21157,N_20599,N_20401);
nand U21158 (N_21158,N_20063,N_20079);
xor U21159 (N_21159,N_20470,N_20403);
xnor U21160 (N_21160,N_20345,N_20384);
xnor U21161 (N_21161,N_20346,N_20620);
nor U21162 (N_21162,N_20238,N_20222);
and U21163 (N_21163,N_20030,N_20503);
or U21164 (N_21164,N_20555,N_20546);
nor U21165 (N_21165,N_20169,N_20505);
nand U21166 (N_21166,N_20544,N_20594);
xor U21167 (N_21167,N_20383,N_20098);
or U21168 (N_21168,N_20022,N_20288);
xnor U21169 (N_21169,N_20325,N_20168);
xnor U21170 (N_21170,N_20480,N_20078);
and U21171 (N_21171,N_20311,N_20516);
or U21172 (N_21172,N_20364,N_20252);
nor U21173 (N_21173,N_20374,N_20587);
xor U21174 (N_21174,N_20358,N_20113);
nor U21175 (N_21175,N_20549,N_20446);
and U21176 (N_21176,N_20072,N_20300);
nand U21177 (N_21177,N_20249,N_20623);
and U21178 (N_21178,N_20226,N_20054);
or U21179 (N_21179,N_20563,N_20425);
xor U21180 (N_21180,N_20456,N_20129);
nor U21181 (N_21181,N_20005,N_20624);
nand U21182 (N_21182,N_20203,N_20124);
or U21183 (N_21183,N_20245,N_20489);
and U21184 (N_21184,N_20541,N_20420);
nor U21185 (N_21185,N_20114,N_20141);
xor U21186 (N_21186,N_20331,N_20037);
nor U21187 (N_21187,N_20131,N_20063);
nand U21188 (N_21188,N_20064,N_20374);
or U21189 (N_21189,N_20073,N_20443);
nor U21190 (N_21190,N_20161,N_20129);
or U21191 (N_21191,N_20126,N_20369);
xor U21192 (N_21192,N_20424,N_20086);
and U21193 (N_21193,N_20393,N_20102);
nand U21194 (N_21194,N_20152,N_20148);
and U21195 (N_21195,N_20029,N_20548);
and U21196 (N_21196,N_20094,N_20365);
xnor U21197 (N_21197,N_20350,N_20100);
nor U21198 (N_21198,N_20568,N_20004);
xnor U21199 (N_21199,N_20304,N_20024);
and U21200 (N_21200,N_20268,N_20136);
xnor U21201 (N_21201,N_20255,N_20173);
xnor U21202 (N_21202,N_20000,N_20033);
nor U21203 (N_21203,N_20013,N_20157);
and U21204 (N_21204,N_20095,N_20125);
and U21205 (N_21205,N_20546,N_20046);
nor U21206 (N_21206,N_20056,N_20314);
and U21207 (N_21207,N_20495,N_20488);
nor U21208 (N_21208,N_20382,N_20027);
nor U21209 (N_21209,N_20222,N_20265);
nor U21210 (N_21210,N_20298,N_20262);
or U21211 (N_21211,N_20399,N_20584);
or U21212 (N_21212,N_20326,N_20256);
xor U21213 (N_21213,N_20168,N_20303);
and U21214 (N_21214,N_20069,N_20041);
xnor U21215 (N_21215,N_20357,N_20388);
and U21216 (N_21216,N_20468,N_20084);
or U21217 (N_21217,N_20264,N_20305);
nand U21218 (N_21218,N_20587,N_20019);
xnor U21219 (N_21219,N_20609,N_20124);
xnor U21220 (N_21220,N_20341,N_20486);
or U21221 (N_21221,N_20576,N_20173);
nand U21222 (N_21222,N_20003,N_20554);
or U21223 (N_21223,N_20278,N_20567);
and U21224 (N_21224,N_20546,N_20464);
nand U21225 (N_21225,N_20254,N_20080);
nand U21226 (N_21226,N_20231,N_20589);
and U21227 (N_21227,N_20008,N_20116);
nor U21228 (N_21228,N_20049,N_20553);
nor U21229 (N_21229,N_20047,N_20048);
nand U21230 (N_21230,N_20015,N_20373);
xnor U21231 (N_21231,N_20189,N_20298);
nor U21232 (N_21232,N_20057,N_20271);
xnor U21233 (N_21233,N_20266,N_20471);
nand U21234 (N_21234,N_20103,N_20398);
nand U21235 (N_21235,N_20174,N_20463);
xnor U21236 (N_21236,N_20135,N_20205);
or U21237 (N_21237,N_20117,N_20131);
or U21238 (N_21238,N_20210,N_20522);
xnor U21239 (N_21239,N_20241,N_20344);
or U21240 (N_21240,N_20390,N_20042);
nor U21241 (N_21241,N_20451,N_20285);
and U21242 (N_21242,N_20061,N_20615);
nand U21243 (N_21243,N_20502,N_20439);
nor U21244 (N_21244,N_20198,N_20266);
nand U21245 (N_21245,N_20414,N_20549);
nor U21246 (N_21246,N_20411,N_20358);
or U21247 (N_21247,N_20275,N_20228);
nand U21248 (N_21248,N_20360,N_20219);
or U21249 (N_21249,N_20359,N_20198);
and U21250 (N_21250,N_20686,N_21093);
and U21251 (N_21251,N_21176,N_21145);
xnor U21252 (N_21252,N_20870,N_21162);
and U21253 (N_21253,N_20945,N_20850);
nor U21254 (N_21254,N_20944,N_21121);
and U21255 (N_21255,N_21197,N_21230);
and U21256 (N_21256,N_21248,N_21092);
xor U21257 (N_21257,N_21052,N_20625);
xnor U21258 (N_21258,N_20931,N_20940);
nor U21259 (N_21259,N_20888,N_20834);
xor U21260 (N_21260,N_20833,N_20878);
nand U21261 (N_21261,N_20797,N_20664);
and U21262 (N_21262,N_21185,N_21165);
or U21263 (N_21263,N_20887,N_20800);
nand U21264 (N_21264,N_21013,N_21178);
or U21265 (N_21265,N_20723,N_21099);
nor U21266 (N_21266,N_21048,N_20710);
and U21267 (N_21267,N_20985,N_20875);
nand U21268 (N_21268,N_21078,N_20802);
and U21269 (N_21269,N_21058,N_21017);
nor U21270 (N_21270,N_20793,N_20928);
or U21271 (N_21271,N_21049,N_20938);
nand U21272 (N_21272,N_21210,N_20704);
nor U21273 (N_21273,N_20974,N_20726);
and U21274 (N_21274,N_20993,N_21135);
nand U21275 (N_21275,N_21232,N_20656);
nand U21276 (N_21276,N_20912,N_20829);
and U21277 (N_21277,N_20825,N_21103);
and U21278 (N_21278,N_20730,N_20702);
or U21279 (N_21279,N_21195,N_21066);
nand U21280 (N_21280,N_20916,N_21198);
and U21281 (N_21281,N_20741,N_21130);
nand U21282 (N_21282,N_21073,N_20860);
nand U21283 (N_21283,N_21149,N_20873);
xor U21284 (N_21284,N_20655,N_21204);
nand U21285 (N_21285,N_20679,N_21116);
xnor U21286 (N_21286,N_20922,N_21004);
nand U21287 (N_21287,N_21079,N_21085);
xnor U21288 (N_21288,N_20995,N_20771);
nor U21289 (N_21289,N_20958,N_20661);
xor U21290 (N_21290,N_20663,N_20971);
or U21291 (N_21291,N_20999,N_20708);
nand U21292 (N_21292,N_21148,N_20847);
xnor U21293 (N_21293,N_21194,N_20784);
or U21294 (N_21294,N_20743,N_20735);
or U21295 (N_21295,N_21213,N_21106);
nor U21296 (N_21296,N_20918,N_21137);
or U21297 (N_21297,N_21018,N_21244);
and U21298 (N_21298,N_20991,N_20738);
xnor U21299 (N_21299,N_20909,N_21247);
and U21300 (N_21300,N_20676,N_20646);
xor U21301 (N_21301,N_20897,N_20841);
and U21302 (N_21302,N_20953,N_20721);
nor U21303 (N_21303,N_20798,N_20920);
nor U21304 (N_21304,N_20924,N_20748);
xor U21305 (N_21305,N_20654,N_20633);
xnor U21306 (N_21306,N_21161,N_20967);
or U21307 (N_21307,N_20822,N_20816);
nand U21308 (N_21308,N_20826,N_20719);
nor U21309 (N_21309,N_20840,N_20705);
or U21310 (N_21310,N_21228,N_20947);
nor U21311 (N_21311,N_20858,N_20683);
and U21312 (N_21312,N_21038,N_21104);
nand U21313 (N_21313,N_21168,N_20791);
nor U21314 (N_21314,N_20803,N_21007);
nor U21315 (N_21315,N_21188,N_20965);
or U21316 (N_21316,N_20998,N_21061);
xor U21317 (N_21317,N_20961,N_20765);
or U21318 (N_21318,N_20864,N_20757);
nand U21319 (N_21319,N_21006,N_20786);
nor U21320 (N_21320,N_21109,N_21229);
or U21321 (N_21321,N_21179,N_20720);
or U21322 (N_21322,N_21154,N_20950);
xor U21323 (N_21323,N_21216,N_21059);
nor U21324 (N_21324,N_20976,N_21095);
nor U21325 (N_21325,N_20811,N_20706);
nand U21326 (N_21326,N_20694,N_20750);
nor U21327 (N_21327,N_20648,N_20792);
or U21328 (N_21328,N_20913,N_20684);
nand U21329 (N_21329,N_21167,N_20713);
nand U21330 (N_21330,N_21050,N_21112);
nand U21331 (N_21331,N_21123,N_21016);
nand U21332 (N_21332,N_20707,N_20796);
nand U21333 (N_21333,N_20914,N_20886);
or U21334 (N_21334,N_21060,N_20749);
and U21335 (N_21335,N_20740,N_20855);
or U21336 (N_21336,N_21243,N_20894);
nand U21337 (N_21337,N_20690,N_21136);
or U21338 (N_21338,N_20682,N_20666);
or U21339 (N_21339,N_21002,N_21055);
and U21340 (N_21340,N_20910,N_21040);
nand U21341 (N_21341,N_21105,N_21011);
nor U21342 (N_21342,N_20815,N_20762);
or U21343 (N_21343,N_21029,N_20980);
nand U21344 (N_21344,N_21172,N_21070);
or U21345 (N_21345,N_20760,N_21037);
and U21346 (N_21346,N_20700,N_20634);
and U21347 (N_21347,N_20722,N_21034);
nor U21348 (N_21348,N_21027,N_20814);
nor U21349 (N_21349,N_21242,N_21126);
and U21350 (N_21350,N_20647,N_20709);
xor U21351 (N_21351,N_20691,N_21031);
nor U21352 (N_21352,N_20836,N_20687);
xnor U21353 (N_21353,N_20729,N_20837);
nor U21354 (N_21354,N_20899,N_20832);
nand U21355 (N_21355,N_20667,N_20978);
or U21356 (N_21356,N_20772,N_21199);
or U21357 (N_21357,N_20775,N_21140);
nor U21358 (N_21358,N_20672,N_21118);
and U21359 (N_21359,N_21019,N_20898);
and U21360 (N_21360,N_20879,N_20992);
xor U21361 (N_21361,N_21152,N_20778);
and U21362 (N_21362,N_20665,N_21009);
xor U21363 (N_21363,N_21045,N_20652);
nand U21364 (N_21364,N_20970,N_21206);
nand U21365 (N_21365,N_21226,N_20804);
and U21366 (N_21366,N_20906,N_20675);
and U21367 (N_21367,N_20968,N_21169);
and U21368 (N_21368,N_20880,N_20662);
nand U21369 (N_21369,N_21205,N_21245);
nor U21370 (N_21370,N_20745,N_20859);
nor U21371 (N_21371,N_21182,N_20979);
nor U21372 (N_21372,N_21097,N_21053);
and U21373 (N_21373,N_21107,N_20857);
nor U21374 (N_21374,N_20724,N_21012);
nor U21375 (N_21375,N_21150,N_20787);
and U21376 (N_21376,N_21224,N_21076);
nor U21377 (N_21377,N_21151,N_20636);
nand U21378 (N_21378,N_21193,N_20923);
xnor U21379 (N_21379,N_20669,N_21187);
or U21380 (N_21380,N_21124,N_21100);
nor U21381 (N_21381,N_21227,N_21025);
xnor U21382 (N_21382,N_20812,N_21147);
nand U21383 (N_21383,N_21131,N_20890);
and U21384 (N_21384,N_20751,N_20739);
nor U21385 (N_21385,N_20981,N_21087);
nor U21386 (N_21386,N_21033,N_21177);
and U21387 (N_21387,N_21222,N_20703);
nand U21388 (N_21388,N_21217,N_20766);
or U21389 (N_21389,N_20865,N_21207);
and U21390 (N_21390,N_21200,N_20761);
nor U21391 (N_21391,N_20695,N_20863);
or U21392 (N_21392,N_20728,N_21115);
xor U21393 (N_21393,N_20810,N_21164);
nand U21394 (N_21394,N_20753,N_20642);
nand U21395 (N_21395,N_20711,N_20900);
nor U21396 (N_21396,N_20698,N_20884);
nor U21397 (N_21397,N_20885,N_20649);
or U21398 (N_21398,N_20877,N_20824);
and U21399 (N_21399,N_21234,N_20628);
nand U21400 (N_21400,N_21237,N_20932);
and U21401 (N_21401,N_20997,N_21241);
or U21402 (N_21402,N_20936,N_21111);
nor U21403 (N_21403,N_21190,N_20807);
xnor U21404 (N_21404,N_21035,N_21056);
xor U21405 (N_21405,N_21156,N_20795);
and U21406 (N_21406,N_20955,N_21067);
nand U21407 (N_21407,N_20972,N_20645);
nor U21408 (N_21408,N_21240,N_20629);
and U21409 (N_21409,N_20754,N_21189);
nor U21410 (N_21410,N_20853,N_21080);
xnor U21411 (N_21411,N_21163,N_20638);
xnor U21412 (N_21412,N_20756,N_21125);
nand U21413 (N_21413,N_20821,N_20809);
and U21414 (N_21414,N_21015,N_21122);
and U21415 (N_21415,N_20986,N_20854);
nand U21416 (N_21416,N_20930,N_20843);
and U21417 (N_21417,N_20882,N_21082);
nand U21418 (N_21418,N_21220,N_20902);
nor U21419 (N_21419,N_21218,N_21026);
nand U21420 (N_21420,N_20927,N_20874);
and U21421 (N_21421,N_21246,N_20963);
or U21422 (N_21422,N_21142,N_21180);
xor U21423 (N_21423,N_21249,N_20966);
or U21424 (N_21424,N_20996,N_21157);
xnor U21425 (N_21425,N_20929,N_20658);
or U21426 (N_21426,N_21223,N_20635);
and U21427 (N_21427,N_20678,N_21021);
xor U21428 (N_21428,N_21098,N_20969);
xor U21429 (N_21429,N_20769,N_21030);
nor U21430 (N_21430,N_20881,N_20794);
nand U21431 (N_21431,N_20827,N_20785);
and U21432 (N_21432,N_21202,N_21215);
nand U21433 (N_21433,N_20670,N_20933);
nor U21434 (N_21434,N_20712,N_21214);
xor U21435 (N_21435,N_21022,N_21139);
nor U21436 (N_21436,N_20718,N_20637);
xor U21437 (N_21437,N_20975,N_20901);
xor U21438 (N_21438,N_20697,N_20790);
xnor U21439 (N_21439,N_20768,N_21032);
and U21440 (N_21440,N_20941,N_21014);
nor U21441 (N_21441,N_20988,N_20752);
or U21442 (N_21442,N_21181,N_21094);
nor U21443 (N_21443,N_20959,N_20872);
xnor U21444 (N_21444,N_21236,N_20942);
or U21445 (N_21445,N_21054,N_20773);
or U21446 (N_21446,N_20759,N_20747);
nor U21447 (N_21447,N_20852,N_20957);
nand U21448 (N_21448,N_20630,N_20977);
xor U21449 (N_21449,N_21064,N_20781);
nor U21450 (N_21450,N_20917,N_21127);
xor U21451 (N_21451,N_21192,N_21075);
nor U21452 (N_21452,N_20962,N_21089);
xor U21453 (N_21453,N_21144,N_20671);
xnor U21454 (N_21454,N_20892,N_20650);
and U21455 (N_21455,N_20819,N_21166);
nand U21456 (N_21456,N_20674,N_20788);
and U21457 (N_21457,N_20736,N_21024);
nor U21458 (N_21458,N_21117,N_20844);
nand U21459 (N_21459,N_20935,N_21065);
or U21460 (N_21460,N_21047,N_21084);
nand U21461 (N_21461,N_20767,N_20848);
or U21462 (N_21462,N_21114,N_20943);
nand U21463 (N_21463,N_20701,N_20763);
and U21464 (N_21464,N_21128,N_21201);
xor U21465 (N_21465,N_20956,N_21069);
xnor U21466 (N_21466,N_20934,N_21183);
nor U21467 (N_21467,N_20983,N_20777);
nor U21468 (N_21468,N_20716,N_21233);
xnor U21469 (N_21469,N_21071,N_21175);
xnor U21470 (N_21470,N_20861,N_20994);
and U21471 (N_21471,N_21096,N_20733);
nor U21472 (N_21472,N_21208,N_21063);
nor U21473 (N_21473,N_20799,N_20820);
and U21474 (N_21474,N_21134,N_20937);
or U21475 (N_21475,N_21196,N_21143);
nor U21476 (N_21476,N_21043,N_21209);
nand U21477 (N_21477,N_21219,N_20903);
nor U21478 (N_21478,N_20990,N_20867);
xor U21479 (N_21479,N_20908,N_20987);
and U21480 (N_21480,N_20641,N_20808);
and U21481 (N_21481,N_20727,N_20868);
nor U21482 (N_21482,N_20849,N_21008);
or U21483 (N_21483,N_21184,N_21235);
nand U21484 (N_21484,N_20689,N_20776);
nand U21485 (N_21485,N_20869,N_20742);
or U21486 (N_21486,N_20926,N_20725);
and U21487 (N_21487,N_20846,N_21138);
xor U21488 (N_21488,N_20925,N_21155);
nor U21489 (N_21489,N_20831,N_21203);
xor U21490 (N_21490,N_21120,N_21173);
nor U21491 (N_21491,N_20696,N_20905);
nor U21492 (N_21492,N_21086,N_20680);
xor U21493 (N_21493,N_20866,N_20659);
xnor U21494 (N_21494,N_20673,N_20813);
xor U21495 (N_21495,N_21191,N_20984);
xnor U21496 (N_21496,N_21113,N_20835);
nand U21497 (N_21497,N_21081,N_20737);
xor U21498 (N_21498,N_20838,N_20677);
xor U21499 (N_21499,N_21005,N_20895);
or U21500 (N_21500,N_21010,N_20871);
nand U21501 (N_21501,N_20732,N_21090);
and U21502 (N_21502,N_21101,N_20949);
nand U21503 (N_21503,N_21231,N_20845);
nand U21504 (N_21504,N_21171,N_20627);
nor U21505 (N_21505,N_21102,N_20692);
and U21506 (N_21506,N_21141,N_20982);
nand U21507 (N_21507,N_21119,N_20688);
nand U21508 (N_21508,N_21074,N_20717);
nor U21509 (N_21509,N_21046,N_20911);
xnor U21510 (N_21510,N_20631,N_20699);
or U21511 (N_21511,N_21036,N_21091);
and U21512 (N_21512,N_20904,N_20806);
or U21513 (N_21513,N_20889,N_21153);
xor U21514 (N_21514,N_20842,N_20746);
nor U21515 (N_21515,N_20693,N_20644);
nand U21516 (N_21516,N_21000,N_20668);
and U21517 (N_21517,N_20764,N_20660);
xor U21518 (N_21518,N_21044,N_20960);
and U21519 (N_21519,N_20755,N_21211);
and U21520 (N_21520,N_20973,N_20734);
xor U21521 (N_21521,N_20839,N_21001);
or U21522 (N_21522,N_20681,N_20939);
or U21523 (N_21523,N_20639,N_20801);
or U21524 (N_21524,N_21129,N_20640);
xnor U21525 (N_21525,N_20657,N_20632);
nor U21526 (N_21526,N_21068,N_21003);
or U21527 (N_21527,N_21186,N_20653);
xor U21528 (N_21528,N_20651,N_21028);
xnor U21529 (N_21529,N_20783,N_20893);
or U21530 (N_21530,N_21023,N_20805);
nor U21531 (N_21531,N_21158,N_20714);
or U21532 (N_21532,N_20946,N_21221);
nor U21533 (N_21533,N_20758,N_21160);
or U21534 (N_21534,N_20876,N_20818);
xnor U21535 (N_21535,N_21132,N_21083);
and U21536 (N_21536,N_21077,N_20685);
or U21537 (N_21537,N_21042,N_21238);
xor U21538 (N_21538,N_20780,N_21057);
nor U21539 (N_21539,N_21212,N_21170);
xnor U21540 (N_21540,N_21088,N_21108);
or U21541 (N_21541,N_21110,N_21225);
nor U21542 (N_21542,N_20948,N_20919);
xor U21543 (N_21543,N_20823,N_20921);
nand U21544 (N_21544,N_21039,N_20883);
xor U21545 (N_21545,N_20907,N_21041);
nand U21546 (N_21546,N_20731,N_21072);
xor U21547 (N_21547,N_20830,N_20851);
nor U21548 (N_21548,N_21159,N_20782);
xor U21549 (N_21549,N_20915,N_20779);
or U21550 (N_21550,N_20952,N_20817);
and U21551 (N_21551,N_20774,N_21062);
xnor U21552 (N_21552,N_21020,N_20715);
and U21553 (N_21553,N_20862,N_20828);
and U21554 (N_21554,N_21239,N_20964);
or U21555 (N_21555,N_21146,N_21051);
and U21556 (N_21556,N_20770,N_21133);
and U21557 (N_21557,N_20856,N_20626);
nand U21558 (N_21558,N_20891,N_20951);
nand U21559 (N_21559,N_20789,N_20954);
or U21560 (N_21560,N_20643,N_21174);
and U21561 (N_21561,N_20896,N_20989);
nor U21562 (N_21562,N_20744,N_21072);
or U21563 (N_21563,N_20689,N_20944);
nor U21564 (N_21564,N_21218,N_20889);
or U21565 (N_21565,N_20762,N_20657);
nand U21566 (N_21566,N_21249,N_20688);
or U21567 (N_21567,N_20812,N_20975);
xor U21568 (N_21568,N_21053,N_21201);
and U21569 (N_21569,N_21168,N_21037);
nand U21570 (N_21570,N_21181,N_20870);
nand U21571 (N_21571,N_21151,N_20920);
xor U21572 (N_21572,N_20907,N_20999);
and U21573 (N_21573,N_20814,N_20997);
and U21574 (N_21574,N_21210,N_21109);
or U21575 (N_21575,N_20962,N_21149);
nand U21576 (N_21576,N_20679,N_21141);
and U21577 (N_21577,N_20825,N_20974);
nor U21578 (N_21578,N_20955,N_20635);
xnor U21579 (N_21579,N_20741,N_20787);
and U21580 (N_21580,N_21094,N_20969);
or U21581 (N_21581,N_20749,N_21242);
and U21582 (N_21582,N_20831,N_20822);
xor U21583 (N_21583,N_20650,N_20757);
nand U21584 (N_21584,N_20867,N_20712);
nor U21585 (N_21585,N_20723,N_20673);
nor U21586 (N_21586,N_21138,N_21195);
nand U21587 (N_21587,N_20664,N_21237);
xnor U21588 (N_21588,N_20775,N_21124);
nand U21589 (N_21589,N_20742,N_20953);
and U21590 (N_21590,N_20634,N_20766);
xnor U21591 (N_21591,N_21138,N_20805);
xnor U21592 (N_21592,N_20988,N_21184);
and U21593 (N_21593,N_21083,N_21158);
nand U21594 (N_21594,N_20855,N_21226);
nor U21595 (N_21595,N_20676,N_20675);
nand U21596 (N_21596,N_21104,N_20931);
nor U21597 (N_21597,N_21133,N_20756);
xor U21598 (N_21598,N_20952,N_20680);
and U21599 (N_21599,N_20906,N_20841);
and U21600 (N_21600,N_20815,N_21215);
nor U21601 (N_21601,N_20730,N_20706);
nor U21602 (N_21602,N_21166,N_21158);
nor U21603 (N_21603,N_21109,N_20957);
xnor U21604 (N_21604,N_21080,N_20907);
nand U21605 (N_21605,N_20788,N_21200);
xor U21606 (N_21606,N_21195,N_20938);
or U21607 (N_21607,N_20976,N_20873);
or U21608 (N_21608,N_21185,N_21052);
xnor U21609 (N_21609,N_20711,N_21209);
or U21610 (N_21610,N_21052,N_20950);
or U21611 (N_21611,N_21239,N_21187);
or U21612 (N_21612,N_21168,N_20763);
or U21613 (N_21613,N_20922,N_21138);
or U21614 (N_21614,N_20765,N_21152);
xor U21615 (N_21615,N_20722,N_21145);
or U21616 (N_21616,N_20821,N_20969);
or U21617 (N_21617,N_20706,N_20777);
and U21618 (N_21618,N_21225,N_20955);
nand U21619 (N_21619,N_20724,N_21241);
nand U21620 (N_21620,N_20878,N_20724);
and U21621 (N_21621,N_20825,N_20803);
nor U21622 (N_21622,N_21105,N_20687);
or U21623 (N_21623,N_20653,N_21113);
and U21624 (N_21624,N_20943,N_21146);
nand U21625 (N_21625,N_21207,N_21036);
xor U21626 (N_21626,N_20718,N_20649);
nor U21627 (N_21627,N_20641,N_20864);
nor U21628 (N_21628,N_21230,N_21214);
or U21629 (N_21629,N_20939,N_20831);
and U21630 (N_21630,N_21208,N_21177);
xor U21631 (N_21631,N_20781,N_21094);
nor U21632 (N_21632,N_21057,N_20740);
nand U21633 (N_21633,N_20913,N_20724);
and U21634 (N_21634,N_20768,N_20637);
xnor U21635 (N_21635,N_20817,N_21202);
nor U21636 (N_21636,N_20635,N_20669);
nand U21637 (N_21637,N_20678,N_21079);
nor U21638 (N_21638,N_20771,N_20702);
xor U21639 (N_21639,N_20795,N_20990);
and U21640 (N_21640,N_21183,N_20650);
and U21641 (N_21641,N_20670,N_21144);
xor U21642 (N_21642,N_21207,N_20915);
nand U21643 (N_21643,N_20724,N_21147);
xor U21644 (N_21644,N_20816,N_20946);
nor U21645 (N_21645,N_21123,N_20967);
or U21646 (N_21646,N_20647,N_20714);
nand U21647 (N_21647,N_20715,N_20916);
xnor U21648 (N_21648,N_20772,N_20864);
nor U21649 (N_21649,N_20872,N_20794);
xor U21650 (N_21650,N_21244,N_21023);
nand U21651 (N_21651,N_20759,N_20654);
or U21652 (N_21652,N_20831,N_21130);
xor U21653 (N_21653,N_20792,N_20890);
xnor U21654 (N_21654,N_21023,N_20979);
xnor U21655 (N_21655,N_21203,N_21201);
nand U21656 (N_21656,N_21058,N_20695);
or U21657 (N_21657,N_20846,N_20843);
and U21658 (N_21658,N_21117,N_21002);
and U21659 (N_21659,N_21024,N_21243);
or U21660 (N_21660,N_20846,N_20823);
and U21661 (N_21661,N_21056,N_20786);
nor U21662 (N_21662,N_21016,N_21205);
nor U21663 (N_21663,N_20802,N_21211);
xor U21664 (N_21664,N_21134,N_20946);
nor U21665 (N_21665,N_21001,N_20690);
nor U21666 (N_21666,N_21020,N_21172);
and U21667 (N_21667,N_20823,N_20859);
xnor U21668 (N_21668,N_21042,N_20977);
xnor U21669 (N_21669,N_20663,N_20857);
and U21670 (N_21670,N_21208,N_21220);
nand U21671 (N_21671,N_20673,N_20920);
xnor U21672 (N_21672,N_21108,N_21064);
or U21673 (N_21673,N_21089,N_20933);
and U21674 (N_21674,N_20783,N_20895);
nor U21675 (N_21675,N_20668,N_20749);
nand U21676 (N_21676,N_21042,N_21001);
nor U21677 (N_21677,N_21009,N_21192);
xor U21678 (N_21678,N_21161,N_20947);
or U21679 (N_21679,N_20752,N_21097);
nor U21680 (N_21680,N_20680,N_21234);
nand U21681 (N_21681,N_21034,N_21113);
and U21682 (N_21682,N_20808,N_20662);
xor U21683 (N_21683,N_21108,N_20948);
or U21684 (N_21684,N_20675,N_21189);
nand U21685 (N_21685,N_20846,N_20729);
and U21686 (N_21686,N_20661,N_20778);
or U21687 (N_21687,N_20905,N_20924);
or U21688 (N_21688,N_20924,N_20846);
nand U21689 (N_21689,N_21057,N_21244);
xor U21690 (N_21690,N_20696,N_20686);
nand U21691 (N_21691,N_20787,N_20627);
xor U21692 (N_21692,N_20668,N_20876);
nor U21693 (N_21693,N_20670,N_21214);
xnor U21694 (N_21694,N_20655,N_20934);
xor U21695 (N_21695,N_21151,N_20940);
nor U21696 (N_21696,N_21083,N_20643);
and U21697 (N_21697,N_21109,N_20680);
nor U21698 (N_21698,N_20948,N_20966);
or U21699 (N_21699,N_20820,N_21235);
or U21700 (N_21700,N_21082,N_20744);
xor U21701 (N_21701,N_20953,N_20681);
and U21702 (N_21702,N_20962,N_21071);
or U21703 (N_21703,N_20828,N_21063);
nand U21704 (N_21704,N_20668,N_21071);
xor U21705 (N_21705,N_21167,N_21181);
nor U21706 (N_21706,N_20785,N_21136);
and U21707 (N_21707,N_20837,N_21105);
xor U21708 (N_21708,N_20735,N_20789);
nor U21709 (N_21709,N_20934,N_20843);
xnor U21710 (N_21710,N_20723,N_20746);
or U21711 (N_21711,N_20929,N_20963);
and U21712 (N_21712,N_20829,N_20659);
nand U21713 (N_21713,N_20899,N_20803);
xor U21714 (N_21714,N_20744,N_21034);
or U21715 (N_21715,N_20747,N_21156);
and U21716 (N_21716,N_21213,N_20959);
nand U21717 (N_21717,N_21019,N_21065);
or U21718 (N_21718,N_20707,N_20868);
or U21719 (N_21719,N_20628,N_21152);
or U21720 (N_21720,N_20950,N_20842);
xnor U21721 (N_21721,N_20769,N_21052);
or U21722 (N_21722,N_21020,N_21174);
or U21723 (N_21723,N_20741,N_20819);
nor U21724 (N_21724,N_20862,N_20713);
nor U21725 (N_21725,N_20997,N_21103);
xnor U21726 (N_21726,N_20974,N_20921);
nand U21727 (N_21727,N_20881,N_20637);
nand U21728 (N_21728,N_20824,N_21117);
xor U21729 (N_21729,N_20887,N_21045);
or U21730 (N_21730,N_20892,N_21160);
or U21731 (N_21731,N_20634,N_21151);
nand U21732 (N_21732,N_21234,N_20898);
nand U21733 (N_21733,N_21095,N_21072);
and U21734 (N_21734,N_20967,N_20862);
nand U21735 (N_21735,N_21237,N_20682);
nor U21736 (N_21736,N_20901,N_20721);
xnor U21737 (N_21737,N_20794,N_20946);
xnor U21738 (N_21738,N_20751,N_21233);
or U21739 (N_21739,N_20965,N_20845);
xor U21740 (N_21740,N_20695,N_21169);
and U21741 (N_21741,N_21119,N_21233);
nor U21742 (N_21742,N_20958,N_21065);
or U21743 (N_21743,N_20642,N_20888);
nor U21744 (N_21744,N_20690,N_21075);
nor U21745 (N_21745,N_20795,N_21042);
or U21746 (N_21746,N_21051,N_20978);
and U21747 (N_21747,N_20828,N_20919);
or U21748 (N_21748,N_20803,N_20751);
xnor U21749 (N_21749,N_20799,N_21098);
or U21750 (N_21750,N_21012,N_21204);
nand U21751 (N_21751,N_21092,N_20983);
or U21752 (N_21752,N_21066,N_20848);
xor U21753 (N_21753,N_21234,N_20961);
xor U21754 (N_21754,N_20856,N_20686);
nor U21755 (N_21755,N_21151,N_21080);
nor U21756 (N_21756,N_20731,N_20867);
or U21757 (N_21757,N_21058,N_21072);
xnor U21758 (N_21758,N_20996,N_20715);
xnor U21759 (N_21759,N_20924,N_20973);
nor U21760 (N_21760,N_20882,N_20685);
and U21761 (N_21761,N_20898,N_20628);
nand U21762 (N_21762,N_20685,N_20997);
or U21763 (N_21763,N_20775,N_20930);
xnor U21764 (N_21764,N_20689,N_20884);
and U21765 (N_21765,N_21040,N_20723);
and U21766 (N_21766,N_20942,N_21229);
or U21767 (N_21767,N_20776,N_21207);
or U21768 (N_21768,N_20662,N_21183);
or U21769 (N_21769,N_21095,N_20782);
or U21770 (N_21770,N_20948,N_21227);
or U21771 (N_21771,N_21095,N_21138);
nor U21772 (N_21772,N_20957,N_20657);
xor U21773 (N_21773,N_21169,N_20818);
nor U21774 (N_21774,N_21136,N_20960);
nor U21775 (N_21775,N_20930,N_21228);
nand U21776 (N_21776,N_21091,N_20797);
or U21777 (N_21777,N_20666,N_20881);
and U21778 (N_21778,N_20653,N_20956);
xor U21779 (N_21779,N_21237,N_20803);
xor U21780 (N_21780,N_21069,N_21022);
or U21781 (N_21781,N_21157,N_20899);
nor U21782 (N_21782,N_21236,N_20744);
xnor U21783 (N_21783,N_20989,N_21116);
nor U21784 (N_21784,N_21243,N_20759);
xnor U21785 (N_21785,N_21100,N_21106);
nand U21786 (N_21786,N_21249,N_20788);
xnor U21787 (N_21787,N_20850,N_20893);
nand U21788 (N_21788,N_20649,N_21212);
nor U21789 (N_21789,N_21082,N_21073);
nand U21790 (N_21790,N_20843,N_21228);
xnor U21791 (N_21791,N_20945,N_21222);
nand U21792 (N_21792,N_20747,N_20694);
xor U21793 (N_21793,N_20976,N_20999);
nor U21794 (N_21794,N_21073,N_20953);
and U21795 (N_21795,N_20799,N_21139);
or U21796 (N_21796,N_20831,N_20784);
nand U21797 (N_21797,N_21037,N_20836);
and U21798 (N_21798,N_21021,N_20872);
nor U21799 (N_21799,N_21042,N_21105);
nand U21800 (N_21800,N_20828,N_20825);
and U21801 (N_21801,N_20789,N_20668);
and U21802 (N_21802,N_21027,N_21083);
or U21803 (N_21803,N_21022,N_21125);
or U21804 (N_21804,N_20753,N_21163);
xor U21805 (N_21805,N_20818,N_21229);
nand U21806 (N_21806,N_20700,N_20639);
nand U21807 (N_21807,N_20933,N_21037);
nor U21808 (N_21808,N_21018,N_21058);
and U21809 (N_21809,N_21130,N_21071);
xnor U21810 (N_21810,N_21016,N_20777);
or U21811 (N_21811,N_20853,N_20739);
nand U21812 (N_21812,N_21159,N_20766);
and U21813 (N_21813,N_20941,N_21237);
and U21814 (N_21814,N_20989,N_21141);
xnor U21815 (N_21815,N_21081,N_20770);
or U21816 (N_21816,N_20708,N_20808);
xnor U21817 (N_21817,N_20697,N_20747);
nand U21818 (N_21818,N_21067,N_20721);
nand U21819 (N_21819,N_21122,N_20628);
or U21820 (N_21820,N_20956,N_21158);
or U21821 (N_21821,N_20809,N_20769);
and U21822 (N_21822,N_21134,N_21167);
nand U21823 (N_21823,N_20948,N_21011);
xor U21824 (N_21824,N_20705,N_21122);
xor U21825 (N_21825,N_20810,N_20966);
nor U21826 (N_21826,N_20949,N_21177);
xnor U21827 (N_21827,N_20835,N_21002);
nor U21828 (N_21828,N_20954,N_20769);
nand U21829 (N_21829,N_20630,N_21185);
and U21830 (N_21830,N_21159,N_20762);
and U21831 (N_21831,N_20767,N_20830);
or U21832 (N_21832,N_21128,N_21247);
xnor U21833 (N_21833,N_20776,N_21190);
nand U21834 (N_21834,N_20861,N_21046);
nor U21835 (N_21835,N_21016,N_21121);
or U21836 (N_21836,N_20767,N_21153);
and U21837 (N_21837,N_20855,N_20907);
nor U21838 (N_21838,N_21151,N_20786);
xnor U21839 (N_21839,N_21241,N_20898);
nor U21840 (N_21840,N_20842,N_20784);
or U21841 (N_21841,N_21036,N_20630);
xnor U21842 (N_21842,N_20889,N_21170);
xor U21843 (N_21843,N_20919,N_20652);
xnor U21844 (N_21844,N_20664,N_20807);
nand U21845 (N_21845,N_21143,N_20643);
or U21846 (N_21846,N_21002,N_20826);
nand U21847 (N_21847,N_20881,N_20765);
and U21848 (N_21848,N_20898,N_21195);
xor U21849 (N_21849,N_20742,N_20960);
and U21850 (N_21850,N_20813,N_20959);
nor U21851 (N_21851,N_21070,N_21059);
and U21852 (N_21852,N_20849,N_21201);
xor U21853 (N_21853,N_20841,N_20826);
or U21854 (N_21854,N_21179,N_20864);
nor U21855 (N_21855,N_20814,N_21041);
and U21856 (N_21856,N_21092,N_21159);
or U21857 (N_21857,N_21032,N_20985);
nand U21858 (N_21858,N_21011,N_21209);
or U21859 (N_21859,N_20688,N_21172);
nand U21860 (N_21860,N_20777,N_21162);
or U21861 (N_21861,N_20765,N_20969);
and U21862 (N_21862,N_20820,N_20664);
or U21863 (N_21863,N_20866,N_21191);
xor U21864 (N_21864,N_20942,N_20752);
xnor U21865 (N_21865,N_20988,N_20751);
xor U21866 (N_21866,N_20930,N_20778);
xor U21867 (N_21867,N_21179,N_20847);
and U21868 (N_21868,N_20929,N_20715);
nand U21869 (N_21869,N_21076,N_20996);
nor U21870 (N_21870,N_20794,N_20833);
or U21871 (N_21871,N_20715,N_20828);
and U21872 (N_21872,N_20704,N_20936);
or U21873 (N_21873,N_20852,N_21019);
or U21874 (N_21874,N_21198,N_20883);
nor U21875 (N_21875,N_21424,N_21508);
or U21876 (N_21876,N_21739,N_21314);
and U21877 (N_21877,N_21454,N_21404);
or U21878 (N_21878,N_21851,N_21864);
or U21879 (N_21879,N_21538,N_21728);
nand U21880 (N_21880,N_21437,N_21641);
and U21881 (N_21881,N_21661,N_21348);
or U21882 (N_21882,N_21727,N_21825);
and U21883 (N_21883,N_21572,N_21828);
or U21884 (N_21884,N_21465,N_21292);
xnor U21885 (N_21885,N_21276,N_21750);
xnor U21886 (N_21886,N_21430,N_21627);
and U21887 (N_21887,N_21724,N_21257);
nor U21888 (N_21888,N_21767,N_21329);
xor U21889 (N_21889,N_21312,N_21849);
and U21890 (N_21890,N_21815,N_21592);
nor U21891 (N_21891,N_21487,N_21673);
nor U21892 (N_21892,N_21746,N_21281);
or U21893 (N_21893,N_21555,N_21376);
and U21894 (N_21894,N_21391,N_21480);
or U21895 (N_21895,N_21874,N_21269);
nand U21896 (N_21896,N_21556,N_21524);
or U21897 (N_21897,N_21714,N_21854);
xor U21898 (N_21898,N_21637,N_21725);
or U21899 (N_21899,N_21837,N_21692);
and U21900 (N_21900,N_21558,N_21716);
nor U21901 (N_21901,N_21542,N_21321);
nor U21902 (N_21902,N_21742,N_21327);
xnor U21903 (N_21903,N_21510,N_21835);
nor U21904 (N_21904,N_21826,N_21493);
or U21905 (N_21905,N_21683,N_21316);
nand U21906 (N_21906,N_21722,N_21472);
or U21907 (N_21907,N_21405,N_21460);
nor U21908 (N_21908,N_21775,N_21806);
and U21909 (N_21909,N_21288,N_21611);
nor U21910 (N_21910,N_21559,N_21586);
nor U21911 (N_21911,N_21766,N_21579);
nor U21912 (N_21912,N_21740,N_21400);
nor U21913 (N_21913,N_21505,N_21615);
or U21914 (N_21914,N_21810,N_21318);
nand U21915 (N_21915,N_21383,N_21761);
nand U21916 (N_21916,N_21477,N_21525);
xor U21917 (N_21917,N_21549,N_21395);
or U21918 (N_21918,N_21475,N_21413);
nor U21919 (N_21919,N_21319,N_21596);
or U21920 (N_21920,N_21499,N_21646);
nor U21921 (N_21921,N_21676,N_21602);
xnor U21922 (N_21922,N_21358,N_21462);
nor U21923 (N_21923,N_21565,N_21614);
nand U21924 (N_21924,N_21420,N_21467);
or U21925 (N_21925,N_21363,N_21260);
and U21926 (N_21926,N_21494,N_21832);
nand U21927 (N_21927,N_21600,N_21871);
or U21928 (N_21928,N_21675,N_21546);
nand U21929 (N_21929,N_21790,N_21474);
and U21930 (N_21930,N_21526,N_21456);
nand U21931 (N_21931,N_21299,N_21293);
nor U21932 (N_21932,N_21561,N_21416);
nand U21933 (N_21933,N_21492,N_21337);
or U21934 (N_21934,N_21311,N_21515);
xnor U21935 (N_21935,N_21469,N_21660);
nand U21936 (N_21936,N_21710,N_21721);
xor U21937 (N_21937,N_21489,N_21829);
nor U21938 (N_21938,N_21305,N_21712);
and U21939 (N_21939,N_21709,N_21744);
or U21940 (N_21940,N_21265,N_21693);
nor U21941 (N_21941,N_21354,N_21645);
nor U21942 (N_21942,N_21754,N_21352);
or U21943 (N_21943,N_21623,N_21488);
xor U21944 (N_21944,N_21659,N_21313);
nor U21945 (N_21945,N_21575,N_21523);
or U21946 (N_21946,N_21678,N_21844);
or U21947 (N_21947,N_21333,N_21426);
or U21948 (N_21948,N_21450,N_21407);
xor U21949 (N_21949,N_21422,N_21583);
nand U21950 (N_21950,N_21514,N_21254);
or U21951 (N_21951,N_21268,N_21504);
nor U21952 (N_21952,N_21326,N_21440);
xnor U21953 (N_21953,N_21862,N_21340);
nor U21954 (N_21954,N_21394,N_21274);
nor U21955 (N_21955,N_21848,N_21509);
nor U21956 (N_21956,N_21774,N_21713);
xor U21957 (N_21957,N_21624,N_21258);
and U21958 (N_21958,N_21473,N_21808);
nor U21959 (N_21959,N_21418,N_21735);
nand U21960 (N_21960,N_21399,N_21593);
xnor U21961 (N_21961,N_21591,N_21415);
nand U21962 (N_21962,N_21367,N_21671);
nand U21963 (N_21963,N_21631,N_21870);
or U21964 (N_21964,N_21822,N_21670);
xor U21965 (N_21965,N_21279,N_21522);
nor U21966 (N_21966,N_21451,N_21382);
and U21967 (N_21967,N_21397,N_21763);
nor U21968 (N_21968,N_21696,N_21401);
or U21969 (N_21969,N_21599,N_21873);
xnor U21970 (N_21970,N_21361,N_21642);
and U21971 (N_21971,N_21629,N_21362);
nor U21972 (N_21972,N_21668,N_21393);
nand U21973 (N_21973,N_21616,N_21366);
nand U21974 (N_21974,N_21702,N_21604);
and U21975 (N_21975,N_21785,N_21334);
and U21976 (N_21976,N_21536,N_21286);
and U21977 (N_21977,N_21574,N_21685);
nor U21978 (N_21978,N_21632,N_21356);
or U21979 (N_21979,N_21272,N_21264);
nor U21980 (N_21980,N_21866,N_21807);
nand U21981 (N_21981,N_21689,N_21765);
xnor U21982 (N_21982,N_21533,N_21283);
or U21983 (N_21983,N_21700,N_21789);
and U21984 (N_21984,N_21381,N_21601);
nand U21985 (N_21985,N_21364,N_21349);
or U21986 (N_21986,N_21438,N_21375);
and U21987 (N_21987,N_21799,N_21298);
xnor U21988 (N_21988,N_21845,N_21309);
xnor U21989 (N_21989,N_21506,N_21762);
or U21990 (N_21990,N_21324,N_21501);
nor U21991 (N_21991,N_21651,N_21733);
and U21992 (N_21992,N_21609,N_21541);
or U21993 (N_21993,N_21530,N_21436);
xor U21994 (N_21994,N_21461,N_21804);
nor U21995 (N_21995,N_21567,N_21476);
and U21996 (N_21996,N_21824,N_21408);
nand U21997 (N_21997,N_21372,N_21729);
nand U21998 (N_21998,N_21607,N_21540);
and U21999 (N_21999,N_21385,N_21441);
nand U22000 (N_22000,N_21453,N_21731);
xnor U22001 (N_22001,N_21872,N_21396);
xnor U22002 (N_22002,N_21781,N_21369);
nor U22003 (N_22003,N_21296,N_21386);
nor U22004 (N_22004,N_21784,N_21277);
and U22005 (N_22005,N_21650,N_21672);
nand U22006 (N_22006,N_21705,N_21719);
xor U22007 (N_22007,N_21270,N_21791);
or U22008 (N_22008,N_21306,N_21847);
nor U22009 (N_22009,N_21378,N_21534);
xor U22010 (N_22010,N_21447,N_21425);
or U22011 (N_22011,N_21374,N_21764);
nor U22012 (N_22012,N_21535,N_21332);
and U22013 (N_22013,N_21410,N_21390);
and U22014 (N_22014,N_21503,N_21406);
and U22015 (N_22015,N_21626,N_21730);
and U22016 (N_22016,N_21756,N_21863);
or U22017 (N_22017,N_21585,N_21662);
or U22018 (N_22018,N_21582,N_21708);
nand U22019 (N_22019,N_21328,N_21339);
nor U22020 (N_22020,N_21745,N_21442);
and U22021 (N_22021,N_21697,N_21776);
xor U22022 (N_22022,N_21619,N_21285);
or U22023 (N_22023,N_21545,N_21654);
or U22024 (N_22024,N_21387,N_21857);
nand U22025 (N_22025,N_21649,N_21786);
and U22026 (N_22026,N_21679,N_21794);
and U22027 (N_22027,N_21581,N_21695);
xnor U22028 (N_22028,N_21603,N_21351);
or U22029 (N_22029,N_21652,N_21573);
and U22030 (N_22030,N_21830,N_21818);
xor U22031 (N_22031,N_21335,N_21833);
nor U22032 (N_22032,N_21497,N_21723);
xnor U22033 (N_22033,N_21342,N_21428);
nor U22034 (N_22034,N_21443,N_21256);
and U22035 (N_22035,N_21297,N_21295);
nor U22036 (N_22036,N_21373,N_21528);
and U22037 (N_22037,N_21330,N_21531);
nand U22038 (N_22038,N_21344,N_21663);
or U22039 (N_22039,N_21562,N_21800);
nand U22040 (N_22040,N_21552,N_21606);
or U22041 (N_22041,N_21628,N_21414);
or U22042 (N_22042,N_21360,N_21821);
and U22043 (N_22043,N_21856,N_21273);
nand U22044 (N_22044,N_21741,N_21421);
xnor U22045 (N_22045,N_21669,N_21736);
or U22046 (N_22046,N_21483,N_21639);
nand U22047 (N_22047,N_21777,N_21834);
xor U22048 (N_22048,N_21432,N_21551);
nor U22049 (N_22049,N_21468,N_21691);
or U22050 (N_22050,N_21634,N_21304);
xnor U22051 (N_22051,N_21282,N_21434);
xor U22052 (N_22052,N_21655,N_21294);
or U22053 (N_22053,N_21613,N_21353);
nor U22054 (N_22054,N_21518,N_21417);
nand U22055 (N_22055,N_21588,N_21457);
nand U22056 (N_22056,N_21809,N_21263);
and U22057 (N_22057,N_21760,N_21560);
and U22058 (N_22058,N_21435,N_21635);
and U22059 (N_22059,N_21271,N_21841);
nor U22060 (N_22060,N_21496,N_21563);
and U22061 (N_22061,N_21771,N_21865);
or U22062 (N_22062,N_21644,N_21411);
and U22063 (N_22063,N_21684,N_21618);
xor U22064 (N_22064,N_21287,N_21544);
xor U22065 (N_22065,N_21711,N_21755);
nand U22066 (N_22066,N_21507,N_21554);
nand U22067 (N_22067,N_21796,N_21255);
xnor U22068 (N_22068,N_21699,N_21734);
and U22069 (N_22069,N_21550,N_21814);
or U22070 (N_22070,N_21801,N_21738);
nand U22071 (N_22071,N_21365,N_21860);
and U22072 (N_22072,N_21512,N_21732);
and U22073 (N_22073,N_21433,N_21783);
nand U22074 (N_22074,N_21840,N_21617);
nand U22075 (N_22075,N_21491,N_21647);
xor U22076 (N_22076,N_21769,N_21412);
or U22077 (N_22077,N_21812,N_21278);
nor U22078 (N_22078,N_21869,N_21470);
nand U22079 (N_22079,N_21357,N_21802);
or U22080 (N_22080,N_21547,N_21368);
and U22081 (N_22081,N_21584,N_21701);
and U22082 (N_22082,N_21868,N_21466);
nand U22083 (N_22083,N_21490,N_21388);
and U22084 (N_22084,N_21429,N_21570);
and U22085 (N_22085,N_21608,N_21553);
nor U22086 (N_22086,N_21343,N_21817);
nand U22087 (N_22087,N_21392,N_21770);
nor U22088 (N_22088,N_21532,N_21568);
nor U22089 (N_22089,N_21855,N_21737);
nand U22090 (N_22090,N_21300,N_21636);
and U22091 (N_22091,N_21747,N_21569);
and U22092 (N_22092,N_21743,N_21423);
and U22093 (N_22093,N_21773,N_21682);
nor U22094 (N_22094,N_21315,N_21605);
nor U22095 (N_22095,N_21638,N_21498);
and U22096 (N_22096,N_21816,N_21753);
xnor U22097 (N_22097,N_21621,N_21548);
nand U22098 (N_22098,N_21325,N_21748);
and U22099 (N_22099,N_21464,N_21726);
or U22100 (N_22100,N_21500,N_21686);
nor U22101 (N_22101,N_21658,N_21266);
and U22102 (N_22102,N_21543,N_21839);
xor U22103 (N_22103,N_21620,N_21813);
xnor U22104 (N_22104,N_21398,N_21843);
and U22105 (N_22105,N_21580,N_21595);
xor U22106 (N_22106,N_21805,N_21317);
nand U22107 (N_22107,N_21610,N_21502);
nand U22108 (N_22108,N_21811,N_21694);
nor U22109 (N_22109,N_21290,N_21322);
or U22110 (N_22110,N_21370,N_21846);
nand U22111 (N_22111,N_21384,N_21347);
and U22112 (N_22112,N_21752,N_21867);
and U22113 (N_22113,N_21439,N_21749);
and U22114 (N_22114,N_21706,N_21681);
nor U22115 (N_22115,N_21403,N_21704);
xor U22116 (N_22116,N_21590,N_21788);
or U22117 (N_22117,N_21690,N_21341);
nor U22118 (N_22118,N_21516,N_21519);
or U22119 (N_22119,N_21720,N_21838);
or U22120 (N_22120,N_21823,N_21267);
xor U22121 (N_22121,N_21566,N_21350);
nor U22122 (N_22122,N_21657,N_21836);
xnor U22123 (N_22123,N_21853,N_21779);
nand U22124 (N_22124,N_21444,N_21448);
xor U22125 (N_22125,N_21301,N_21571);
xor U22126 (N_22126,N_21751,N_21331);
and U22127 (N_22127,N_21782,N_21759);
and U22128 (N_22128,N_21557,N_21346);
and U22129 (N_22129,N_21797,N_21643);
xor U22130 (N_22130,N_21481,N_21778);
or U22131 (N_22131,N_21633,N_21455);
nand U22132 (N_22132,N_21513,N_21787);
nand U22133 (N_22133,N_21803,N_21259);
nor U22134 (N_22134,N_21576,N_21380);
nor U22135 (N_22135,N_21355,N_21589);
nand U22136 (N_22136,N_21819,N_21597);
and U22137 (N_22137,N_21289,N_21667);
nor U22138 (N_22138,N_21688,N_21291);
nand U22139 (N_22139,N_21640,N_21484);
and U22140 (N_22140,N_21598,N_21338);
or U22141 (N_22141,N_21310,N_21587);
or U22142 (N_22142,N_21261,N_21303);
and U22143 (N_22143,N_21486,N_21861);
nand U22144 (N_22144,N_21594,N_21427);
and U22145 (N_22145,N_21336,N_21648);
or U22146 (N_22146,N_21452,N_21419);
nand U22147 (N_22147,N_21798,N_21389);
nor U22148 (N_22148,N_21768,N_21379);
xor U22149 (N_22149,N_21793,N_21717);
nor U22150 (N_22150,N_21377,N_21320);
xor U22151 (N_22151,N_21666,N_21792);
nor U22152 (N_22152,N_21520,N_21539);
or U22153 (N_22153,N_21458,N_21529);
xor U22154 (N_22154,N_21485,N_21402);
or U22155 (N_22155,N_21831,N_21253);
xor U22156 (N_22156,N_21459,N_21850);
or U22157 (N_22157,N_21827,N_21517);
and U22158 (N_22158,N_21859,N_21284);
nor U22159 (N_22159,N_21680,N_21511);
and U22160 (N_22160,N_21307,N_21622);
nor U22161 (N_22161,N_21479,N_21446);
or U22162 (N_22162,N_21302,N_21262);
nor U22163 (N_22163,N_21674,N_21758);
nor U22164 (N_22164,N_21323,N_21842);
and U22165 (N_22165,N_21478,N_21772);
nor U22166 (N_22166,N_21409,N_21858);
nand U22167 (N_22167,N_21820,N_21578);
or U22168 (N_22168,N_21653,N_21482);
or U22169 (N_22169,N_21521,N_21715);
xor U22170 (N_22170,N_21564,N_21780);
nand U22171 (N_22171,N_21698,N_21431);
xor U22172 (N_22172,N_21250,N_21577);
xor U22173 (N_22173,N_21449,N_21630);
nor U22174 (N_22174,N_21252,N_21275);
nor U22175 (N_22175,N_21371,N_21665);
nor U22176 (N_22176,N_21677,N_21852);
and U22177 (N_22177,N_21280,N_21308);
or U22178 (N_22178,N_21463,N_21359);
and U22179 (N_22179,N_21345,N_21625);
and U22180 (N_22180,N_21495,N_21795);
and U22181 (N_22181,N_21707,N_21251);
xnor U22182 (N_22182,N_21718,N_21445);
xor U22183 (N_22183,N_21664,N_21757);
and U22184 (N_22184,N_21527,N_21687);
nand U22185 (N_22185,N_21471,N_21537);
nand U22186 (N_22186,N_21656,N_21612);
xnor U22187 (N_22187,N_21703,N_21400);
xnor U22188 (N_22188,N_21494,N_21258);
xnor U22189 (N_22189,N_21495,N_21386);
and U22190 (N_22190,N_21365,N_21375);
or U22191 (N_22191,N_21289,N_21744);
xnor U22192 (N_22192,N_21302,N_21454);
nor U22193 (N_22193,N_21461,N_21281);
and U22194 (N_22194,N_21512,N_21488);
or U22195 (N_22195,N_21628,N_21512);
and U22196 (N_22196,N_21404,N_21277);
xnor U22197 (N_22197,N_21804,N_21671);
or U22198 (N_22198,N_21529,N_21322);
nor U22199 (N_22199,N_21634,N_21671);
and U22200 (N_22200,N_21757,N_21855);
nor U22201 (N_22201,N_21734,N_21463);
or U22202 (N_22202,N_21649,N_21788);
or U22203 (N_22203,N_21748,N_21668);
xor U22204 (N_22204,N_21659,N_21268);
nor U22205 (N_22205,N_21506,N_21355);
xor U22206 (N_22206,N_21598,N_21600);
or U22207 (N_22207,N_21832,N_21492);
nor U22208 (N_22208,N_21256,N_21280);
xnor U22209 (N_22209,N_21819,N_21727);
and U22210 (N_22210,N_21607,N_21730);
nor U22211 (N_22211,N_21475,N_21570);
nor U22212 (N_22212,N_21837,N_21612);
nand U22213 (N_22213,N_21489,N_21747);
nor U22214 (N_22214,N_21387,N_21615);
nor U22215 (N_22215,N_21430,N_21421);
nor U22216 (N_22216,N_21421,N_21870);
nand U22217 (N_22217,N_21336,N_21385);
nand U22218 (N_22218,N_21363,N_21861);
nand U22219 (N_22219,N_21622,N_21428);
nor U22220 (N_22220,N_21557,N_21345);
and U22221 (N_22221,N_21485,N_21686);
nor U22222 (N_22222,N_21349,N_21831);
xnor U22223 (N_22223,N_21529,N_21747);
xnor U22224 (N_22224,N_21706,N_21533);
nand U22225 (N_22225,N_21688,N_21528);
or U22226 (N_22226,N_21479,N_21679);
nor U22227 (N_22227,N_21263,N_21824);
xnor U22228 (N_22228,N_21598,N_21343);
or U22229 (N_22229,N_21312,N_21764);
nor U22230 (N_22230,N_21765,N_21561);
nand U22231 (N_22231,N_21557,N_21469);
nor U22232 (N_22232,N_21294,N_21257);
or U22233 (N_22233,N_21581,N_21557);
nand U22234 (N_22234,N_21669,N_21695);
or U22235 (N_22235,N_21515,N_21548);
nor U22236 (N_22236,N_21548,N_21281);
and U22237 (N_22237,N_21608,N_21470);
nor U22238 (N_22238,N_21603,N_21796);
or U22239 (N_22239,N_21589,N_21662);
or U22240 (N_22240,N_21544,N_21790);
nor U22241 (N_22241,N_21357,N_21678);
or U22242 (N_22242,N_21463,N_21445);
and U22243 (N_22243,N_21544,N_21668);
and U22244 (N_22244,N_21311,N_21324);
or U22245 (N_22245,N_21718,N_21339);
nor U22246 (N_22246,N_21800,N_21873);
nand U22247 (N_22247,N_21549,N_21811);
nor U22248 (N_22248,N_21828,N_21582);
nand U22249 (N_22249,N_21372,N_21571);
nand U22250 (N_22250,N_21559,N_21439);
nor U22251 (N_22251,N_21859,N_21319);
and U22252 (N_22252,N_21265,N_21318);
and U22253 (N_22253,N_21628,N_21339);
and U22254 (N_22254,N_21406,N_21665);
nor U22255 (N_22255,N_21853,N_21673);
and U22256 (N_22256,N_21742,N_21281);
nand U22257 (N_22257,N_21552,N_21484);
xnor U22258 (N_22258,N_21583,N_21742);
nand U22259 (N_22259,N_21411,N_21754);
and U22260 (N_22260,N_21721,N_21446);
xor U22261 (N_22261,N_21724,N_21328);
xor U22262 (N_22262,N_21669,N_21581);
or U22263 (N_22263,N_21697,N_21835);
xor U22264 (N_22264,N_21692,N_21762);
xor U22265 (N_22265,N_21812,N_21492);
or U22266 (N_22266,N_21720,N_21400);
xor U22267 (N_22267,N_21290,N_21608);
nor U22268 (N_22268,N_21335,N_21502);
or U22269 (N_22269,N_21435,N_21694);
xnor U22270 (N_22270,N_21686,N_21789);
nor U22271 (N_22271,N_21786,N_21533);
and U22272 (N_22272,N_21550,N_21594);
xor U22273 (N_22273,N_21805,N_21388);
xor U22274 (N_22274,N_21462,N_21781);
xnor U22275 (N_22275,N_21357,N_21371);
nand U22276 (N_22276,N_21715,N_21739);
xnor U22277 (N_22277,N_21657,N_21819);
nor U22278 (N_22278,N_21504,N_21839);
nor U22279 (N_22279,N_21856,N_21554);
and U22280 (N_22280,N_21808,N_21404);
xor U22281 (N_22281,N_21714,N_21759);
nor U22282 (N_22282,N_21291,N_21486);
nor U22283 (N_22283,N_21362,N_21427);
xor U22284 (N_22284,N_21414,N_21816);
nor U22285 (N_22285,N_21738,N_21283);
nand U22286 (N_22286,N_21727,N_21738);
nand U22287 (N_22287,N_21598,N_21400);
nor U22288 (N_22288,N_21565,N_21667);
nor U22289 (N_22289,N_21390,N_21815);
or U22290 (N_22290,N_21691,N_21671);
and U22291 (N_22291,N_21654,N_21406);
or U22292 (N_22292,N_21300,N_21319);
nand U22293 (N_22293,N_21345,N_21683);
and U22294 (N_22294,N_21556,N_21571);
or U22295 (N_22295,N_21485,N_21569);
or U22296 (N_22296,N_21334,N_21389);
or U22297 (N_22297,N_21869,N_21505);
and U22298 (N_22298,N_21690,N_21834);
nand U22299 (N_22299,N_21332,N_21814);
xnor U22300 (N_22300,N_21531,N_21556);
nand U22301 (N_22301,N_21515,N_21354);
xnor U22302 (N_22302,N_21420,N_21663);
or U22303 (N_22303,N_21613,N_21359);
nor U22304 (N_22304,N_21791,N_21798);
nor U22305 (N_22305,N_21327,N_21672);
nand U22306 (N_22306,N_21533,N_21787);
or U22307 (N_22307,N_21280,N_21550);
nor U22308 (N_22308,N_21805,N_21841);
nor U22309 (N_22309,N_21632,N_21836);
xor U22310 (N_22310,N_21858,N_21794);
or U22311 (N_22311,N_21844,N_21416);
xor U22312 (N_22312,N_21711,N_21642);
and U22313 (N_22313,N_21612,N_21680);
nand U22314 (N_22314,N_21538,N_21793);
xor U22315 (N_22315,N_21505,N_21378);
or U22316 (N_22316,N_21764,N_21825);
or U22317 (N_22317,N_21622,N_21660);
and U22318 (N_22318,N_21445,N_21586);
nand U22319 (N_22319,N_21572,N_21472);
or U22320 (N_22320,N_21678,N_21748);
xor U22321 (N_22321,N_21720,N_21325);
nor U22322 (N_22322,N_21289,N_21595);
nand U22323 (N_22323,N_21545,N_21404);
and U22324 (N_22324,N_21374,N_21254);
xor U22325 (N_22325,N_21651,N_21375);
or U22326 (N_22326,N_21325,N_21333);
or U22327 (N_22327,N_21597,N_21530);
nand U22328 (N_22328,N_21800,N_21586);
xor U22329 (N_22329,N_21359,N_21451);
and U22330 (N_22330,N_21256,N_21775);
nand U22331 (N_22331,N_21600,N_21558);
or U22332 (N_22332,N_21573,N_21343);
and U22333 (N_22333,N_21628,N_21409);
nand U22334 (N_22334,N_21278,N_21808);
and U22335 (N_22335,N_21848,N_21707);
nor U22336 (N_22336,N_21809,N_21771);
nor U22337 (N_22337,N_21647,N_21456);
or U22338 (N_22338,N_21299,N_21708);
or U22339 (N_22339,N_21561,N_21531);
xnor U22340 (N_22340,N_21491,N_21591);
nand U22341 (N_22341,N_21869,N_21670);
or U22342 (N_22342,N_21463,N_21378);
nor U22343 (N_22343,N_21533,N_21296);
and U22344 (N_22344,N_21371,N_21646);
nor U22345 (N_22345,N_21714,N_21393);
nand U22346 (N_22346,N_21691,N_21571);
and U22347 (N_22347,N_21675,N_21416);
nor U22348 (N_22348,N_21344,N_21673);
and U22349 (N_22349,N_21555,N_21398);
nor U22350 (N_22350,N_21678,N_21626);
or U22351 (N_22351,N_21610,N_21793);
xnor U22352 (N_22352,N_21351,N_21856);
xnor U22353 (N_22353,N_21462,N_21828);
nand U22354 (N_22354,N_21276,N_21303);
and U22355 (N_22355,N_21556,N_21563);
nand U22356 (N_22356,N_21320,N_21636);
nor U22357 (N_22357,N_21426,N_21704);
xor U22358 (N_22358,N_21509,N_21318);
or U22359 (N_22359,N_21806,N_21504);
nor U22360 (N_22360,N_21823,N_21818);
and U22361 (N_22361,N_21722,N_21661);
and U22362 (N_22362,N_21546,N_21463);
and U22363 (N_22363,N_21522,N_21782);
xor U22364 (N_22364,N_21573,N_21607);
nand U22365 (N_22365,N_21776,N_21595);
nor U22366 (N_22366,N_21482,N_21782);
nor U22367 (N_22367,N_21845,N_21545);
nand U22368 (N_22368,N_21720,N_21411);
nor U22369 (N_22369,N_21529,N_21422);
nand U22370 (N_22370,N_21679,N_21598);
or U22371 (N_22371,N_21448,N_21331);
and U22372 (N_22372,N_21372,N_21423);
nor U22373 (N_22373,N_21499,N_21354);
and U22374 (N_22374,N_21810,N_21631);
or U22375 (N_22375,N_21599,N_21290);
or U22376 (N_22376,N_21693,N_21298);
and U22377 (N_22377,N_21566,N_21253);
xnor U22378 (N_22378,N_21459,N_21718);
nand U22379 (N_22379,N_21742,N_21778);
and U22380 (N_22380,N_21822,N_21699);
and U22381 (N_22381,N_21759,N_21763);
nor U22382 (N_22382,N_21696,N_21393);
and U22383 (N_22383,N_21851,N_21707);
or U22384 (N_22384,N_21782,N_21558);
nor U22385 (N_22385,N_21778,N_21781);
xnor U22386 (N_22386,N_21357,N_21255);
and U22387 (N_22387,N_21472,N_21369);
nand U22388 (N_22388,N_21733,N_21712);
nand U22389 (N_22389,N_21404,N_21587);
nor U22390 (N_22390,N_21652,N_21829);
or U22391 (N_22391,N_21490,N_21863);
nand U22392 (N_22392,N_21778,N_21871);
nand U22393 (N_22393,N_21525,N_21330);
and U22394 (N_22394,N_21717,N_21519);
nor U22395 (N_22395,N_21553,N_21286);
and U22396 (N_22396,N_21873,N_21814);
xor U22397 (N_22397,N_21722,N_21510);
or U22398 (N_22398,N_21800,N_21637);
xor U22399 (N_22399,N_21445,N_21438);
nor U22400 (N_22400,N_21745,N_21646);
nor U22401 (N_22401,N_21481,N_21869);
nand U22402 (N_22402,N_21742,N_21458);
or U22403 (N_22403,N_21873,N_21743);
xnor U22404 (N_22404,N_21670,N_21459);
nor U22405 (N_22405,N_21626,N_21497);
xor U22406 (N_22406,N_21489,N_21758);
or U22407 (N_22407,N_21526,N_21564);
nor U22408 (N_22408,N_21487,N_21413);
nand U22409 (N_22409,N_21637,N_21862);
or U22410 (N_22410,N_21379,N_21709);
and U22411 (N_22411,N_21666,N_21771);
and U22412 (N_22412,N_21468,N_21313);
xnor U22413 (N_22413,N_21523,N_21689);
and U22414 (N_22414,N_21356,N_21709);
or U22415 (N_22415,N_21435,N_21356);
nand U22416 (N_22416,N_21429,N_21517);
nor U22417 (N_22417,N_21580,N_21545);
nor U22418 (N_22418,N_21592,N_21498);
xnor U22419 (N_22419,N_21374,N_21689);
or U22420 (N_22420,N_21686,N_21513);
nand U22421 (N_22421,N_21702,N_21425);
xnor U22422 (N_22422,N_21413,N_21511);
and U22423 (N_22423,N_21383,N_21837);
nand U22424 (N_22424,N_21652,N_21286);
and U22425 (N_22425,N_21577,N_21461);
nor U22426 (N_22426,N_21514,N_21263);
and U22427 (N_22427,N_21550,N_21390);
nor U22428 (N_22428,N_21641,N_21420);
and U22429 (N_22429,N_21257,N_21469);
and U22430 (N_22430,N_21775,N_21460);
or U22431 (N_22431,N_21676,N_21750);
xor U22432 (N_22432,N_21620,N_21522);
nand U22433 (N_22433,N_21551,N_21575);
xnor U22434 (N_22434,N_21693,N_21382);
nand U22435 (N_22435,N_21281,N_21328);
or U22436 (N_22436,N_21864,N_21431);
or U22437 (N_22437,N_21381,N_21315);
nand U22438 (N_22438,N_21808,N_21256);
nand U22439 (N_22439,N_21811,N_21403);
nor U22440 (N_22440,N_21653,N_21605);
nor U22441 (N_22441,N_21370,N_21643);
and U22442 (N_22442,N_21703,N_21756);
and U22443 (N_22443,N_21538,N_21535);
nor U22444 (N_22444,N_21408,N_21715);
nor U22445 (N_22445,N_21632,N_21526);
nand U22446 (N_22446,N_21760,N_21693);
xnor U22447 (N_22447,N_21672,N_21759);
nor U22448 (N_22448,N_21616,N_21737);
or U22449 (N_22449,N_21601,N_21839);
nand U22450 (N_22450,N_21547,N_21683);
xnor U22451 (N_22451,N_21593,N_21864);
nor U22452 (N_22452,N_21825,N_21385);
or U22453 (N_22453,N_21361,N_21282);
nor U22454 (N_22454,N_21796,N_21805);
and U22455 (N_22455,N_21604,N_21375);
nand U22456 (N_22456,N_21596,N_21822);
and U22457 (N_22457,N_21702,N_21469);
and U22458 (N_22458,N_21576,N_21652);
nand U22459 (N_22459,N_21633,N_21413);
or U22460 (N_22460,N_21521,N_21408);
xnor U22461 (N_22461,N_21614,N_21587);
nand U22462 (N_22462,N_21741,N_21292);
and U22463 (N_22463,N_21364,N_21290);
xor U22464 (N_22464,N_21727,N_21441);
or U22465 (N_22465,N_21860,N_21506);
xnor U22466 (N_22466,N_21623,N_21272);
and U22467 (N_22467,N_21847,N_21671);
nand U22468 (N_22468,N_21362,N_21797);
nor U22469 (N_22469,N_21811,N_21253);
nor U22470 (N_22470,N_21806,N_21739);
and U22471 (N_22471,N_21564,N_21654);
xnor U22472 (N_22472,N_21634,N_21641);
nor U22473 (N_22473,N_21270,N_21483);
and U22474 (N_22474,N_21479,N_21782);
or U22475 (N_22475,N_21779,N_21717);
xor U22476 (N_22476,N_21304,N_21476);
xnor U22477 (N_22477,N_21443,N_21730);
nand U22478 (N_22478,N_21568,N_21735);
nor U22479 (N_22479,N_21402,N_21328);
and U22480 (N_22480,N_21435,N_21436);
nand U22481 (N_22481,N_21506,N_21294);
or U22482 (N_22482,N_21302,N_21736);
xor U22483 (N_22483,N_21639,N_21474);
and U22484 (N_22484,N_21254,N_21763);
xor U22485 (N_22485,N_21865,N_21677);
and U22486 (N_22486,N_21405,N_21766);
xnor U22487 (N_22487,N_21606,N_21833);
and U22488 (N_22488,N_21636,N_21539);
and U22489 (N_22489,N_21579,N_21742);
or U22490 (N_22490,N_21350,N_21300);
and U22491 (N_22491,N_21433,N_21754);
or U22492 (N_22492,N_21693,N_21857);
or U22493 (N_22493,N_21578,N_21795);
xnor U22494 (N_22494,N_21864,N_21632);
xnor U22495 (N_22495,N_21540,N_21711);
nand U22496 (N_22496,N_21799,N_21584);
or U22497 (N_22497,N_21510,N_21688);
and U22498 (N_22498,N_21874,N_21451);
or U22499 (N_22499,N_21364,N_21824);
xor U22500 (N_22500,N_21961,N_22006);
xnor U22501 (N_22501,N_22204,N_21931);
or U22502 (N_22502,N_22441,N_21957);
and U22503 (N_22503,N_22299,N_22057);
nand U22504 (N_22504,N_22402,N_22121);
and U22505 (N_22505,N_22021,N_22040);
xnor U22506 (N_22506,N_22349,N_22265);
xnor U22507 (N_22507,N_22080,N_22115);
xnor U22508 (N_22508,N_22301,N_21956);
nor U22509 (N_22509,N_22059,N_22109);
nand U22510 (N_22510,N_21968,N_21910);
nor U22511 (N_22511,N_22172,N_22048);
nor U22512 (N_22512,N_22184,N_22353);
nor U22513 (N_22513,N_22027,N_22091);
xor U22514 (N_22514,N_22014,N_22208);
nand U22515 (N_22515,N_22219,N_22403);
nor U22516 (N_22516,N_22147,N_22134);
nor U22517 (N_22517,N_22036,N_21877);
xnor U22518 (N_22518,N_22264,N_22022);
nand U22519 (N_22519,N_22181,N_22360);
or U22520 (N_22520,N_21890,N_22466);
xnor U22521 (N_22521,N_22187,N_22019);
and U22522 (N_22522,N_22170,N_21976);
and U22523 (N_22523,N_21982,N_22231);
and U22524 (N_22524,N_22042,N_22128);
and U22525 (N_22525,N_22224,N_22162);
nor U22526 (N_22526,N_22285,N_22207);
xnor U22527 (N_22527,N_22126,N_21886);
nand U22528 (N_22528,N_22029,N_22391);
or U22529 (N_22529,N_22442,N_22116);
nor U22530 (N_22530,N_22125,N_22364);
nand U22531 (N_22531,N_22337,N_22223);
or U22532 (N_22532,N_21879,N_22098);
or U22533 (N_22533,N_22387,N_22086);
and U22534 (N_22534,N_22497,N_22405);
xnor U22535 (N_22535,N_21889,N_21917);
nand U22536 (N_22536,N_22076,N_22038);
nor U22537 (N_22537,N_22238,N_22350);
nand U22538 (N_22538,N_21993,N_22220);
nor U22539 (N_22539,N_21951,N_22490);
and U22540 (N_22540,N_21875,N_22093);
nand U22541 (N_22541,N_22439,N_22020);
nand U22542 (N_22542,N_22133,N_22335);
nand U22543 (N_22543,N_22061,N_22448);
xor U22544 (N_22544,N_21958,N_22324);
nor U22545 (N_22545,N_22176,N_22169);
nor U22546 (N_22546,N_22232,N_22499);
nor U22547 (N_22547,N_22105,N_22461);
xor U22548 (N_22548,N_22140,N_22248);
xor U22549 (N_22549,N_22124,N_22357);
or U22550 (N_22550,N_22097,N_21934);
or U22551 (N_22551,N_22111,N_21992);
or U22552 (N_22552,N_22395,N_22090);
xnor U22553 (N_22553,N_22137,N_21905);
xnor U22554 (N_22554,N_22339,N_22287);
or U22555 (N_22555,N_22229,N_22319);
nand U22556 (N_22556,N_22127,N_22000);
nor U22557 (N_22557,N_21983,N_21988);
or U22558 (N_22558,N_22320,N_21935);
nor U22559 (N_22559,N_22252,N_21954);
or U22560 (N_22560,N_21895,N_22347);
or U22561 (N_22561,N_22321,N_22253);
xnor U22562 (N_22562,N_21939,N_22274);
or U22563 (N_22563,N_22263,N_22377);
nor U22564 (N_22564,N_22278,N_22492);
and U22565 (N_22565,N_22008,N_22420);
or U22566 (N_22566,N_22180,N_22283);
xor U22567 (N_22567,N_22362,N_22393);
or U22568 (N_22568,N_22414,N_21928);
xor U22569 (N_22569,N_22119,N_22191);
xnor U22570 (N_22570,N_22049,N_22400);
or U22571 (N_22571,N_22483,N_22454);
xor U22572 (N_22572,N_22182,N_21906);
or U22573 (N_22573,N_22135,N_21930);
nand U22574 (N_22574,N_22277,N_22205);
nor U22575 (N_22575,N_22068,N_22446);
and U22576 (N_22576,N_22469,N_22046);
nor U22577 (N_22577,N_22388,N_21994);
and U22578 (N_22578,N_22150,N_22236);
nand U22579 (N_22579,N_22235,N_22072);
nand U22580 (N_22580,N_21972,N_22409);
nand U22581 (N_22581,N_21977,N_22112);
nand U22582 (N_22582,N_22331,N_22160);
or U22583 (N_22583,N_22254,N_21911);
nor U22584 (N_22584,N_22437,N_22241);
xor U22585 (N_22585,N_22142,N_22450);
nand U22586 (N_22586,N_22206,N_22078);
xnor U22587 (N_22587,N_22089,N_22193);
or U22588 (N_22588,N_22230,N_22455);
and U22589 (N_22589,N_22416,N_21902);
nand U22590 (N_22590,N_22177,N_21880);
nand U22591 (N_22591,N_22404,N_22002);
nor U22592 (N_22592,N_22034,N_21967);
or U22593 (N_22593,N_22067,N_22183);
and U22594 (N_22594,N_21900,N_22026);
nor U22595 (N_22595,N_22330,N_21922);
or U22596 (N_22596,N_22408,N_22296);
and U22597 (N_22597,N_22394,N_22381);
nand U22598 (N_22598,N_22424,N_22294);
or U22599 (N_22599,N_21901,N_22120);
xnor U22600 (N_22600,N_22435,N_22227);
nand U22601 (N_22601,N_22210,N_21876);
nand U22602 (N_22602,N_21903,N_21947);
nor U22603 (N_22603,N_22380,N_22188);
nor U22604 (N_22604,N_22173,N_21920);
xor U22605 (N_22605,N_21986,N_22001);
nand U22606 (N_22606,N_22488,N_22348);
and U22607 (N_22607,N_21999,N_22043);
xor U22608 (N_22608,N_21897,N_22412);
nand U22609 (N_22609,N_22203,N_21949);
or U22610 (N_22610,N_21887,N_22275);
and U22611 (N_22611,N_22298,N_22444);
nor U22612 (N_22612,N_22246,N_22312);
or U22613 (N_22613,N_22386,N_22302);
or U22614 (N_22614,N_22392,N_22131);
nor U22615 (N_22615,N_22256,N_21884);
xnor U22616 (N_22616,N_22481,N_22062);
nor U22617 (N_22617,N_21925,N_22005);
nor U22618 (N_22618,N_22028,N_22269);
xnor U22619 (N_22619,N_21883,N_22212);
nor U22620 (N_22620,N_22175,N_22385);
nand U22621 (N_22621,N_22276,N_22372);
xor U22622 (N_22622,N_22174,N_22165);
nor U22623 (N_22623,N_22477,N_21996);
nand U22624 (N_22624,N_22251,N_22167);
xnor U22625 (N_22625,N_22015,N_22398);
and U22626 (N_22626,N_22399,N_21978);
xnor U22627 (N_22627,N_21963,N_22250);
xor U22628 (N_22628,N_21918,N_22103);
nor U22629 (N_22629,N_22009,N_21981);
nand U22630 (N_22630,N_22132,N_22311);
and U22631 (N_22631,N_21893,N_22157);
nand U22632 (N_22632,N_22375,N_22194);
nor U22633 (N_22633,N_22260,N_21938);
xnor U22634 (N_22634,N_22305,N_22138);
nand U22635 (N_22635,N_22280,N_22092);
or U22636 (N_22636,N_22214,N_22082);
and U22637 (N_22637,N_21975,N_22159);
nor U22638 (N_22638,N_22318,N_22139);
or U22639 (N_22639,N_21950,N_22069);
xor U22640 (N_22640,N_22491,N_22085);
xnor U22641 (N_22641,N_22423,N_22289);
or U22642 (N_22642,N_22432,N_22270);
nor U22643 (N_22643,N_22343,N_21984);
and U22644 (N_22644,N_22051,N_22401);
or U22645 (N_22645,N_22024,N_22242);
nor U22646 (N_22646,N_22104,N_22056);
xor U22647 (N_22647,N_22023,N_22498);
nand U22648 (N_22648,N_21899,N_22178);
xor U22649 (N_22649,N_22267,N_22351);
nor U22650 (N_22650,N_22415,N_22145);
xnor U22651 (N_22651,N_22130,N_22475);
nand U22652 (N_22652,N_22255,N_21885);
nor U22653 (N_22653,N_22443,N_22050);
nor U22654 (N_22654,N_22007,N_22272);
nand U22655 (N_22655,N_22243,N_21881);
or U22656 (N_22656,N_22213,N_22419);
nor U22657 (N_22657,N_21964,N_22179);
xor U22658 (N_22658,N_22326,N_22379);
and U22659 (N_22659,N_22334,N_21944);
xnor U22660 (N_22660,N_22281,N_22070);
nor U22661 (N_22661,N_21985,N_22237);
and U22662 (N_22662,N_22291,N_22407);
xnor U22663 (N_22663,N_22114,N_22101);
xnor U22664 (N_22664,N_21973,N_22382);
and U22665 (N_22665,N_22218,N_22100);
or U22666 (N_22666,N_22390,N_22313);
nand U22667 (N_22667,N_22164,N_22452);
and U22668 (N_22668,N_22003,N_22447);
nand U22669 (N_22669,N_22356,N_22035);
nand U22670 (N_22670,N_22368,N_22290);
nor U22671 (N_22671,N_21894,N_22359);
nor U22672 (N_22672,N_22077,N_22032);
and U22673 (N_22673,N_22096,N_22457);
nand U22674 (N_22674,N_22438,N_21966);
or U22675 (N_22675,N_22411,N_22480);
xnor U22676 (N_22676,N_22456,N_22118);
xnor U22677 (N_22677,N_22149,N_22016);
nand U22678 (N_22678,N_22462,N_22471);
nand U22679 (N_22679,N_22433,N_21990);
nand U22680 (N_22680,N_22155,N_22216);
xnor U22681 (N_22681,N_22463,N_22106);
or U22682 (N_22682,N_22249,N_22425);
nor U22683 (N_22683,N_22123,N_22327);
nor U22684 (N_22684,N_22322,N_22054);
and U22685 (N_22685,N_21927,N_21896);
or U22686 (N_22686,N_22282,N_22095);
nor U22687 (N_22687,N_21960,N_22371);
xnor U22688 (N_22688,N_22310,N_22245);
xor U22689 (N_22689,N_22010,N_22148);
or U22690 (N_22690,N_21914,N_22358);
xor U22691 (N_22691,N_22222,N_22033);
and U22692 (N_22692,N_22374,N_21924);
nor U22693 (N_22693,N_22268,N_21882);
nor U22694 (N_22694,N_22279,N_22239);
and U22695 (N_22695,N_21912,N_22081);
and U22696 (N_22696,N_22211,N_21941);
or U22697 (N_22697,N_21898,N_22485);
nand U22698 (N_22698,N_22189,N_22384);
or U22699 (N_22699,N_21913,N_21892);
nor U22700 (N_22700,N_22489,N_22151);
and U22701 (N_22701,N_21904,N_22293);
xor U22702 (N_22702,N_22474,N_22261);
or U22703 (N_22703,N_22426,N_22493);
xor U22704 (N_22704,N_22292,N_22304);
xor U22705 (N_22705,N_21971,N_22300);
or U22706 (N_22706,N_22262,N_22284);
nand U22707 (N_22707,N_21915,N_22185);
xor U22708 (N_22708,N_22041,N_22200);
or U22709 (N_22709,N_22136,N_22389);
and U22710 (N_22710,N_22030,N_21936);
and U22711 (N_22711,N_22060,N_22018);
and U22712 (N_22712,N_22053,N_22445);
nor U22713 (N_22713,N_21891,N_22113);
or U22714 (N_22714,N_21995,N_22044);
xor U22715 (N_22715,N_22378,N_22328);
xor U22716 (N_22716,N_22234,N_22064);
xor U22717 (N_22717,N_22266,N_22017);
nor U22718 (N_22718,N_21945,N_22325);
nor U22719 (N_22719,N_22141,N_22215);
xnor U22720 (N_22720,N_22197,N_22440);
xnor U22721 (N_22721,N_22465,N_21991);
nor U22722 (N_22722,N_22217,N_22484);
nor U22723 (N_22723,N_21955,N_22468);
or U22724 (N_22724,N_22088,N_22244);
nor U22725 (N_22725,N_21969,N_21998);
nand U22726 (N_22726,N_22476,N_22354);
and U22727 (N_22727,N_22171,N_22233);
or U22728 (N_22728,N_22195,N_22075);
and U22729 (N_22729,N_22110,N_22122);
or U22730 (N_22730,N_22323,N_22058);
nor U22731 (N_22731,N_22158,N_22434);
and U22732 (N_22732,N_22094,N_22099);
nand U22733 (N_22733,N_22117,N_22315);
xor U22734 (N_22734,N_22365,N_22190);
xnor U22735 (N_22735,N_21929,N_21989);
nand U22736 (N_22736,N_22288,N_22161);
nor U22737 (N_22737,N_22079,N_22317);
nand U22738 (N_22738,N_21923,N_22453);
or U22739 (N_22739,N_21942,N_22329);
nor U22740 (N_22740,N_21953,N_22429);
xor U22741 (N_22741,N_22352,N_22168);
nand U22742 (N_22742,N_22369,N_21919);
nor U22743 (N_22743,N_22199,N_22494);
and U22744 (N_22744,N_22039,N_22073);
nor U22745 (N_22745,N_22376,N_22449);
xor U22746 (N_22746,N_22346,N_22472);
and U22747 (N_22747,N_22355,N_22473);
or U22748 (N_22748,N_22406,N_22209);
xnor U22749 (N_22749,N_21921,N_22226);
nor U22750 (N_22750,N_22108,N_22083);
or U22751 (N_22751,N_21937,N_22436);
xnor U22752 (N_22752,N_22367,N_22340);
nor U22753 (N_22753,N_22052,N_21962);
nor U22754 (N_22754,N_22063,N_21909);
and U22755 (N_22755,N_22308,N_22186);
nand U22756 (N_22756,N_22306,N_22427);
and U22757 (N_22757,N_22045,N_22166);
and U22758 (N_22758,N_22011,N_22307);
and U22759 (N_22759,N_22153,N_22418);
nor U22760 (N_22760,N_22156,N_22336);
nand U22761 (N_22761,N_22065,N_21952);
nand U22762 (N_22762,N_22240,N_21965);
and U22763 (N_22763,N_22397,N_22102);
nand U22764 (N_22764,N_22370,N_22482);
nor U22765 (N_22765,N_22192,N_21908);
and U22766 (N_22766,N_21997,N_21888);
and U22767 (N_22767,N_22273,N_22202);
or U22768 (N_22768,N_21959,N_22004);
nor U22769 (N_22769,N_22459,N_22417);
xnor U22770 (N_22770,N_22496,N_21987);
nor U22771 (N_22771,N_22198,N_22146);
nor U22772 (N_22772,N_22344,N_22413);
nor U22773 (N_22773,N_22295,N_22458);
nor U22774 (N_22774,N_22366,N_22373);
xnor U22775 (N_22775,N_21916,N_22163);
xnor U22776 (N_22776,N_22196,N_22012);
nor U22777 (N_22777,N_22037,N_21878);
or U22778 (N_22778,N_22055,N_22286);
or U22779 (N_22779,N_22410,N_22479);
xor U22780 (N_22780,N_22345,N_22152);
or U22781 (N_22781,N_22396,N_22074);
nand U22782 (N_22782,N_21980,N_22470);
or U22783 (N_22783,N_22129,N_22271);
nor U22784 (N_22784,N_22460,N_21943);
nand U22785 (N_22785,N_22467,N_21979);
or U22786 (N_22786,N_22333,N_22143);
nor U22787 (N_22787,N_22297,N_22428);
xnor U22788 (N_22788,N_22144,N_22478);
nor U22789 (N_22789,N_22495,N_22430);
and U22790 (N_22790,N_22383,N_21932);
and U22791 (N_22791,N_22087,N_22341);
nor U22792 (N_22792,N_22259,N_22486);
nand U22793 (N_22793,N_22332,N_22228);
nand U22794 (N_22794,N_22316,N_22309);
nand U22795 (N_22795,N_22487,N_21948);
nand U22796 (N_22796,N_22013,N_22225);
nor U22797 (N_22797,N_22047,N_22247);
nor U22798 (N_22798,N_22342,N_21907);
nand U22799 (N_22799,N_22464,N_22257);
xor U22800 (N_22800,N_22025,N_22031);
and U22801 (N_22801,N_22422,N_22154);
xnor U22802 (N_22802,N_21933,N_22338);
and U22803 (N_22803,N_22451,N_21974);
and U22804 (N_22804,N_22107,N_21940);
nor U22805 (N_22805,N_21970,N_21926);
or U22806 (N_22806,N_22361,N_22084);
xor U22807 (N_22807,N_22314,N_22221);
or U22808 (N_22808,N_22431,N_22363);
and U22809 (N_22809,N_21946,N_22303);
nand U22810 (N_22810,N_22258,N_22201);
and U22811 (N_22811,N_22071,N_22421);
xnor U22812 (N_22812,N_22066,N_22305);
xnor U22813 (N_22813,N_22380,N_22335);
and U22814 (N_22814,N_21980,N_22417);
and U22815 (N_22815,N_22236,N_22415);
and U22816 (N_22816,N_22070,N_22078);
or U22817 (N_22817,N_21951,N_22155);
nor U22818 (N_22818,N_22327,N_22342);
nor U22819 (N_22819,N_22061,N_22020);
nor U22820 (N_22820,N_22012,N_22106);
nand U22821 (N_22821,N_22095,N_22322);
or U22822 (N_22822,N_22334,N_21904);
nor U22823 (N_22823,N_22358,N_22239);
nor U22824 (N_22824,N_22469,N_22223);
nor U22825 (N_22825,N_21941,N_22222);
and U22826 (N_22826,N_21917,N_22427);
and U22827 (N_22827,N_22225,N_22455);
nor U22828 (N_22828,N_22050,N_22216);
or U22829 (N_22829,N_22496,N_21996);
or U22830 (N_22830,N_22323,N_22245);
or U22831 (N_22831,N_21959,N_22135);
xor U22832 (N_22832,N_22065,N_22415);
or U22833 (N_22833,N_22483,N_22247);
xor U22834 (N_22834,N_22305,N_22292);
xor U22835 (N_22835,N_22395,N_22109);
or U22836 (N_22836,N_22466,N_22272);
and U22837 (N_22837,N_22199,N_22314);
or U22838 (N_22838,N_21929,N_22167);
nand U22839 (N_22839,N_22138,N_21931);
nor U22840 (N_22840,N_21934,N_22358);
or U22841 (N_22841,N_22046,N_22254);
or U22842 (N_22842,N_21929,N_21962);
or U22843 (N_22843,N_22142,N_22024);
and U22844 (N_22844,N_22134,N_22360);
and U22845 (N_22845,N_22150,N_22477);
xnor U22846 (N_22846,N_21938,N_22336);
nand U22847 (N_22847,N_21886,N_21883);
or U22848 (N_22848,N_22468,N_22338);
xor U22849 (N_22849,N_21962,N_22075);
xnor U22850 (N_22850,N_22407,N_22303);
nand U22851 (N_22851,N_22261,N_22251);
nand U22852 (N_22852,N_22257,N_22169);
nand U22853 (N_22853,N_22265,N_21977);
nand U22854 (N_22854,N_22192,N_21915);
nand U22855 (N_22855,N_22066,N_21965);
and U22856 (N_22856,N_22078,N_22088);
nor U22857 (N_22857,N_22444,N_21996);
and U22858 (N_22858,N_22481,N_21906);
and U22859 (N_22859,N_21997,N_21957);
nor U22860 (N_22860,N_22136,N_22210);
nand U22861 (N_22861,N_21945,N_21960);
and U22862 (N_22862,N_22216,N_21988);
or U22863 (N_22863,N_22283,N_22314);
and U22864 (N_22864,N_22358,N_21899);
nor U22865 (N_22865,N_22277,N_21923);
nor U22866 (N_22866,N_22027,N_22033);
nor U22867 (N_22867,N_22139,N_22249);
xnor U22868 (N_22868,N_21955,N_22247);
xor U22869 (N_22869,N_22457,N_22056);
nand U22870 (N_22870,N_22149,N_22039);
or U22871 (N_22871,N_22161,N_21949);
and U22872 (N_22872,N_22238,N_22250);
nor U22873 (N_22873,N_22103,N_22456);
xnor U22874 (N_22874,N_22378,N_21961);
or U22875 (N_22875,N_22480,N_22043);
nor U22876 (N_22876,N_22263,N_22176);
nor U22877 (N_22877,N_22089,N_21970);
and U22878 (N_22878,N_22067,N_22203);
xor U22879 (N_22879,N_22407,N_22016);
xor U22880 (N_22880,N_22498,N_21982);
or U22881 (N_22881,N_22103,N_22256);
nor U22882 (N_22882,N_22104,N_22237);
or U22883 (N_22883,N_22214,N_21983);
nor U22884 (N_22884,N_22425,N_22332);
or U22885 (N_22885,N_22128,N_22377);
and U22886 (N_22886,N_22167,N_22239);
or U22887 (N_22887,N_21972,N_21960);
xnor U22888 (N_22888,N_22051,N_22069);
xnor U22889 (N_22889,N_22391,N_22212);
nor U22890 (N_22890,N_22354,N_22339);
nor U22891 (N_22891,N_22027,N_22422);
or U22892 (N_22892,N_22285,N_22427);
nand U22893 (N_22893,N_22074,N_22433);
nand U22894 (N_22894,N_22410,N_21931);
nand U22895 (N_22895,N_22215,N_22388);
xor U22896 (N_22896,N_21986,N_22301);
nor U22897 (N_22897,N_22264,N_22140);
nand U22898 (N_22898,N_22269,N_22362);
nand U22899 (N_22899,N_22184,N_22481);
nand U22900 (N_22900,N_22364,N_22255);
xor U22901 (N_22901,N_21955,N_22081);
nand U22902 (N_22902,N_22169,N_21884);
xnor U22903 (N_22903,N_22016,N_22163);
nor U22904 (N_22904,N_22144,N_22484);
and U22905 (N_22905,N_22358,N_22376);
xnor U22906 (N_22906,N_22081,N_22405);
or U22907 (N_22907,N_22238,N_21903);
and U22908 (N_22908,N_22103,N_21903);
or U22909 (N_22909,N_22031,N_22480);
or U22910 (N_22910,N_22174,N_22387);
nand U22911 (N_22911,N_21989,N_21955);
nand U22912 (N_22912,N_22055,N_22019);
xor U22913 (N_22913,N_21973,N_22143);
nand U22914 (N_22914,N_22234,N_22127);
nand U22915 (N_22915,N_22266,N_22400);
nor U22916 (N_22916,N_22187,N_22067);
xnor U22917 (N_22917,N_21898,N_21949);
or U22918 (N_22918,N_22292,N_22310);
nor U22919 (N_22919,N_22033,N_21915);
xor U22920 (N_22920,N_22330,N_22395);
and U22921 (N_22921,N_22135,N_22498);
and U22922 (N_22922,N_22368,N_22258);
nand U22923 (N_22923,N_22267,N_22389);
or U22924 (N_22924,N_22031,N_21963);
nand U22925 (N_22925,N_22062,N_22307);
and U22926 (N_22926,N_22165,N_22300);
or U22927 (N_22927,N_22210,N_22223);
and U22928 (N_22928,N_21985,N_22343);
nand U22929 (N_22929,N_22160,N_22493);
nor U22930 (N_22930,N_22426,N_22390);
xnor U22931 (N_22931,N_22021,N_21894);
xnor U22932 (N_22932,N_22375,N_22096);
and U22933 (N_22933,N_22009,N_21889);
xnor U22934 (N_22934,N_22458,N_22187);
nor U22935 (N_22935,N_22488,N_22005);
nor U22936 (N_22936,N_22055,N_22049);
xnor U22937 (N_22937,N_21923,N_22009);
or U22938 (N_22938,N_22443,N_22447);
or U22939 (N_22939,N_22128,N_21883);
and U22940 (N_22940,N_21875,N_22098);
nand U22941 (N_22941,N_22406,N_21947);
xnor U22942 (N_22942,N_22098,N_22244);
xnor U22943 (N_22943,N_22129,N_22482);
xnor U22944 (N_22944,N_22245,N_22451);
nor U22945 (N_22945,N_22106,N_22370);
or U22946 (N_22946,N_22258,N_22353);
nor U22947 (N_22947,N_22490,N_22330);
nand U22948 (N_22948,N_22349,N_22210);
or U22949 (N_22949,N_22211,N_22309);
nor U22950 (N_22950,N_22222,N_22131);
nor U22951 (N_22951,N_22062,N_21946);
xor U22952 (N_22952,N_22224,N_22463);
nand U22953 (N_22953,N_22009,N_21885);
xor U22954 (N_22954,N_22265,N_22407);
or U22955 (N_22955,N_21925,N_22003);
nand U22956 (N_22956,N_21908,N_22438);
xor U22957 (N_22957,N_21949,N_22370);
nand U22958 (N_22958,N_21984,N_22014);
and U22959 (N_22959,N_22315,N_22067);
xnor U22960 (N_22960,N_22070,N_22386);
xor U22961 (N_22961,N_22050,N_22278);
nand U22962 (N_22962,N_22288,N_21998);
or U22963 (N_22963,N_22380,N_22466);
nor U22964 (N_22964,N_22252,N_22099);
nor U22965 (N_22965,N_22285,N_22435);
nand U22966 (N_22966,N_22318,N_22264);
and U22967 (N_22967,N_22195,N_22388);
and U22968 (N_22968,N_22088,N_22030);
xnor U22969 (N_22969,N_22348,N_22394);
xor U22970 (N_22970,N_22377,N_22208);
and U22971 (N_22971,N_22250,N_22043);
nor U22972 (N_22972,N_22280,N_22418);
nand U22973 (N_22973,N_21886,N_22356);
xnor U22974 (N_22974,N_22232,N_22344);
and U22975 (N_22975,N_21936,N_22235);
and U22976 (N_22976,N_21956,N_22335);
nand U22977 (N_22977,N_22076,N_22469);
or U22978 (N_22978,N_22138,N_22112);
xor U22979 (N_22979,N_22460,N_22215);
nor U22980 (N_22980,N_22289,N_21953);
xor U22981 (N_22981,N_22023,N_21984);
or U22982 (N_22982,N_22182,N_22456);
xor U22983 (N_22983,N_22185,N_22453);
nand U22984 (N_22984,N_22144,N_22272);
or U22985 (N_22985,N_22168,N_21977);
and U22986 (N_22986,N_22158,N_22485);
or U22987 (N_22987,N_22145,N_22479);
and U22988 (N_22988,N_22061,N_22250);
or U22989 (N_22989,N_22395,N_22268);
or U22990 (N_22990,N_22220,N_22128);
nor U22991 (N_22991,N_22275,N_22071);
nand U22992 (N_22992,N_22495,N_21963);
nor U22993 (N_22993,N_22340,N_22365);
nor U22994 (N_22994,N_22037,N_22332);
nor U22995 (N_22995,N_22185,N_21885);
xor U22996 (N_22996,N_22208,N_22146);
and U22997 (N_22997,N_22384,N_22194);
or U22998 (N_22998,N_22359,N_22293);
nand U22999 (N_22999,N_22141,N_22409);
and U23000 (N_23000,N_22380,N_22427);
xor U23001 (N_23001,N_22338,N_21951);
xnor U23002 (N_23002,N_22020,N_22113);
xor U23003 (N_23003,N_22304,N_22051);
nor U23004 (N_23004,N_22445,N_22098);
nand U23005 (N_23005,N_22032,N_22196);
nor U23006 (N_23006,N_21958,N_22365);
nand U23007 (N_23007,N_22060,N_22117);
nor U23008 (N_23008,N_22026,N_22123);
nand U23009 (N_23009,N_22004,N_22019);
xor U23010 (N_23010,N_22482,N_22179);
and U23011 (N_23011,N_21903,N_22381);
xnor U23012 (N_23012,N_22257,N_22435);
nor U23013 (N_23013,N_22210,N_22380);
nor U23014 (N_23014,N_22208,N_21966);
and U23015 (N_23015,N_22026,N_22266);
xnor U23016 (N_23016,N_22029,N_22483);
xor U23017 (N_23017,N_22187,N_21954);
and U23018 (N_23018,N_22127,N_22071);
nor U23019 (N_23019,N_21901,N_22205);
nand U23020 (N_23020,N_21882,N_21935);
xnor U23021 (N_23021,N_21881,N_22027);
nand U23022 (N_23022,N_22292,N_22495);
nand U23023 (N_23023,N_22009,N_22006);
or U23024 (N_23024,N_22096,N_22265);
xor U23025 (N_23025,N_22454,N_22452);
or U23026 (N_23026,N_21980,N_22170);
or U23027 (N_23027,N_22017,N_21915);
nand U23028 (N_23028,N_22343,N_22231);
nand U23029 (N_23029,N_21924,N_22150);
or U23030 (N_23030,N_22337,N_22438);
and U23031 (N_23031,N_22014,N_22402);
or U23032 (N_23032,N_22123,N_22028);
or U23033 (N_23033,N_22151,N_22302);
and U23034 (N_23034,N_21887,N_22115);
xnor U23035 (N_23035,N_22192,N_22213);
and U23036 (N_23036,N_22411,N_21915);
xnor U23037 (N_23037,N_22382,N_22206);
xnor U23038 (N_23038,N_22445,N_22185);
and U23039 (N_23039,N_22099,N_21915);
xor U23040 (N_23040,N_22375,N_22370);
xnor U23041 (N_23041,N_22344,N_22058);
xnor U23042 (N_23042,N_21988,N_22156);
nand U23043 (N_23043,N_22314,N_22467);
xor U23044 (N_23044,N_22172,N_22060);
and U23045 (N_23045,N_22038,N_21892);
nand U23046 (N_23046,N_22464,N_22282);
xor U23047 (N_23047,N_22065,N_22126);
and U23048 (N_23048,N_22309,N_22248);
or U23049 (N_23049,N_22286,N_22433);
nor U23050 (N_23050,N_22418,N_22395);
and U23051 (N_23051,N_22424,N_22285);
nor U23052 (N_23052,N_22331,N_22403);
xor U23053 (N_23053,N_22021,N_22088);
nand U23054 (N_23054,N_21982,N_21976);
and U23055 (N_23055,N_22164,N_22290);
nand U23056 (N_23056,N_22394,N_22237);
and U23057 (N_23057,N_21943,N_21895);
and U23058 (N_23058,N_22232,N_21946);
nor U23059 (N_23059,N_22237,N_21877);
nor U23060 (N_23060,N_22228,N_22462);
and U23061 (N_23061,N_22435,N_21922);
nor U23062 (N_23062,N_22171,N_22142);
nand U23063 (N_23063,N_22456,N_22320);
nand U23064 (N_23064,N_21959,N_22060);
or U23065 (N_23065,N_22390,N_22392);
xor U23066 (N_23066,N_22157,N_21878);
or U23067 (N_23067,N_22177,N_22404);
and U23068 (N_23068,N_21930,N_22069);
nand U23069 (N_23069,N_22345,N_21883);
or U23070 (N_23070,N_22381,N_21924);
or U23071 (N_23071,N_22329,N_22375);
nand U23072 (N_23072,N_22335,N_22303);
xor U23073 (N_23073,N_22457,N_22114);
nand U23074 (N_23074,N_21897,N_22298);
or U23075 (N_23075,N_22286,N_21884);
nor U23076 (N_23076,N_22139,N_22272);
xnor U23077 (N_23077,N_22440,N_22131);
or U23078 (N_23078,N_22243,N_22345);
xnor U23079 (N_23079,N_21913,N_22334);
nor U23080 (N_23080,N_21990,N_21943);
or U23081 (N_23081,N_22060,N_22209);
nor U23082 (N_23082,N_22369,N_22432);
nor U23083 (N_23083,N_22307,N_22416);
nor U23084 (N_23084,N_22355,N_21907);
or U23085 (N_23085,N_22372,N_22358);
nand U23086 (N_23086,N_22122,N_22215);
nor U23087 (N_23087,N_22110,N_22444);
xnor U23088 (N_23088,N_22074,N_22398);
nand U23089 (N_23089,N_22328,N_22094);
or U23090 (N_23090,N_22370,N_21960);
and U23091 (N_23091,N_22404,N_22057);
xor U23092 (N_23092,N_22085,N_22069);
nand U23093 (N_23093,N_21892,N_22134);
nand U23094 (N_23094,N_22226,N_22164);
or U23095 (N_23095,N_22037,N_22138);
nand U23096 (N_23096,N_22126,N_21920);
and U23097 (N_23097,N_21907,N_22161);
nor U23098 (N_23098,N_21926,N_22490);
and U23099 (N_23099,N_22488,N_22027);
nor U23100 (N_23100,N_22205,N_21984);
nor U23101 (N_23101,N_22046,N_22149);
xor U23102 (N_23102,N_22078,N_22185);
nand U23103 (N_23103,N_22225,N_22199);
or U23104 (N_23104,N_22451,N_22141);
nand U23105 (N_23105,N_22198,N_22160);
nand U23106 (N_23106,N_22033,N_22307);
xnor U23107 (N_23107,N_22188,N_22172);
and U23108 (N_23108,N_22483,N_22206);
nand U23109 (N_23109,N_22326,N_22392);
nand U23110 (N_23110,N_22363,N_22025);
xnor U23111 (N_23111,N_22428,N_22113);
and U23112 (N_23112,N_22186,N_21951);
nor U23113 (N_23113,N_22328,N_22355);
and U23114 (N_23114,N_22277,N_22062);
or U23115 (N_23115,N_22415,N_22283);
nand U23116 (N_23116,N_21876,N_21968);
nor U23117 (N_23117,N_22349,N_22444);
nor U23118 (N_23118,N_22135,N_22286);
and U23119 (N_23119,N_22368,N_22064);
or U23120 (N_23120,N_22251,N_22213);
nand U23121 (N_23121,N_22320,N_22005);
nand U23122 (N_23122,N_22106,N_22364);
and U23123 (N_23123,N_22083,N_22439);
and U23124 (N_23124,N_21979,N_21877);
nor U23125 (N_23125,N_23053,N_22724);
xor U23126 (N_23126,N_22711,N_22956);
nand U23127 (N_23127,N_22675,N_22510);
or U23128 (N_23128,N_23123,N_22502);
xnor U23129 (N_23129,N_22640,N_23052);
and U23130 (N_23130,N_22784,N_22573);
nor U23131 (N_23131,N_22868,N_22607);
nand U23132 (N_23132,N_23096,N_22568);
xnor U23133 (N_23133,N_22951,N_23028);
nor U23134 (N_23134,N_22958,N_22516);
nor U23135 (N_23135,N_22959,N_22507);
nor U23136 (N_23136,N_22637,N_23080);
nand U23137 (N_23137,N_22582,N_22955);
xor U23138 (N_23138,N_22830,N_22985);
nor U23139 (N_23139,N_22878,N_22850);
nand U23140 (N_23140,N_22741,N_22973);
nand U23141 (N_23141,N_22964,N_22677);
xnor U23142 (N_23142,N_23104,N_22936);
nand U23143 (N_23143,N_22528,N_22881);
nand U23144 (N_23144,N_22639,N_22605);
nor U23145 (N_23145,N_23010,N_22836);
nor U23146 (N_23146,N_22511,N_23050);
xnor U23147 (N_23147,N_22932,N_22734);
and U23148 (N_23148,N_22522,N_22901);
or U23149 (N_23149,N_22898,N_22740);
xnor U23150 (N_23150,N_22861,N_23007);
nand U23151 (N_23151,N_22949,N_22902);
or U23152 (N_23152,N_22681,N_22565);
and U23153 (N_23153,N_22738,N_22648);
and U23154 (N_23154,N_22783,N_22655);
xnor U23155 (N_23155,N_23030,N_23069);
nand U23156 (N_23156,N_22524,N_22937);
nor U23157 (N_23157,N_22555,N_22925);
nand U23158 (N_23158,N_22508,N_22723);
nor U23159 (N_23159,N_22853,N_22796);
nand U23160 (N_23160,N_22577,N_22722);
nand U23161 (N_23161,N_22774,N_22550);
or U23162 (N_23162,N_22644,N_22874);
or U23163 (N_23163,N_22893,N_22814);
xor U23164 (N_23164,N_23061,N_22781);
or U23165 (N_23165,N_22755,N_22752);
nand U23166 (N_23166,N_22993,N_22915);
and U23167 (N_23167,N_22700,N_22883);
xnor U23168 (N_23168,N_22650,N_22616);
nand U23169 (N_23169,N_23040,N_22547);
or U23170 (N_23170,N_22967,N_22660);
nand U23171 (N_23171,N_22886,N_23015);
nor U23172 (N_23172,N_22795,N_23094);
nand U23173 (N_23173,N_22669,N_22745);
nor U23174 (N_23174,N_23012,N_23115);
nand U23175 (N_23175,N_22743,N_22584);
or U23176 (N_23176,N_23033,N_23017);
and U23177 (N_23177,N_22979,N_22569);
nor U23178 (N_23178,N_22978,N_22908);
nor U23179 (N_23179,N_22788,N_22835);
nor U23180 (N_23180,N_22939,N_22710);
and U23181 (N_23181,N_22517,N_22884);
nand U23182 (N_23182,N_22633,N_23026);
nand U23183 (N_23183,N_23065,N_22818);
and U23184 (N_23184,N_22732,N_22802);
xnor U23185 (N_23185,N_22930,N_23064);
xnor U23186 (N_23186,N_22894,N_23071);
xor U23187 (N_23187,N_22923,N_22667);
nor U23188 (N_23188,N_23109,N_22841);
nand U23189 (N_23189,N_22576,N_22594);
xnor U23190 (N_23190,N_22540,N_22578);
nor U23191 (N_23191,N_22621,N_23066);
nor U23192 (N_23192,N_22614,N_22909);
or U23193 (N_23193,N_22876,N_22572);
or U23194 (N_23194,N_22513,N_22651);
xnor U23195 (N_23195,N_22847,N_22845);
or U23196 (N_23196,N_23077,N_23035);
xnor U23197 (N_23197,N_22623,N_22636);
xor U23198 (N_23198,N_22707,N_22635);
nor U23199 (N_23199,N_22778,N_23022);
nand U23200 (N_23200,N_22982,N_22823);
and U23201 (N_23201,N_22684,N_22629);
or U23202 (N_23202,N_22599,N_22529);
or U23203 (N_23203,N_22759,N_22805);
nor U23204 (N_23204,N_22856,N_22574);
xnor U23205 (N_23205,N_23042,N_22882);
nand U23206 (N_23206,N_22996,N_22604);
and U23207 (N_23207,N_22934,N_22679);
xnor U23208 (N_23208,N_22963,N_22981);
nand U23209 (N_23209,N_22763,N_22945);
nand U23210 (N_23210,N_22606,N_22666);
nor U23211 (N_23211,N_23034,N_22846);
or U23212 (N_23212,N_22548,N_23073);
nor U23213 (N_23213,N_22833,N_22962);
nor U23214 (N_23214,N_22900,N_22747);
xnor U23215 (N_23215,N_23114,N_22736);
nand U23216 (N_23216,N_23044,N_23072);
xnor U23217 (N_23217,N_23113,N_22709);
xor U23218 (N_23218,N_23037,N_22543);
nor U23219 (N_23219,N_22843,N_22652);
and U23220 (N_23220,N_22720,N_22779);
or U23221 (N_23221,N_23041,N_23106);
xnor U23222 (N_23222,N_22770,N_22941);
xor U23223 (N_23223,N_22698,N_22873);
nand U23224 (N_23224,N_22597,N_23031);
and U23225 (N_23225,N_22702,N_22626);
nand U23226 (N_23226,N_22521,N_23048);
or U23227 (N_23227,N_22602,N_22704);
or U23228 (N_23228,N_22974,N_22505);
nand U23229 (N_23229,N_22831,N_22731);
nand U23230 (N_23230,N_22773,N_23057);
nand U23231 (N_23231,N_22609,N_23056);
or U23232 (N_23232,N_22880,N_22822);
or U23233 (N_23233,N_22891,N_22813);
or U23234 (N_23234,N_22857,N_22598);
nor U23235 (N_23235,N_22791,N_22559);
or U23236 (N_23236,N_22950,N_22819);
or U23237 (N_23237,N_22921,N_22536);
or U23238 (N_23238,N_22997,N_22692);
nand U23239 (N_23239,N_22627,N_22662);
xnor U23240 (N_23240,N_22775,N_22638);
or U23241 (N_23241,N_22571,N_22674);
or U23242 (N_23242,N_23009,N_22793);
xnor U23243 (N_23243,N_22794,N_22533);
and U23244 (N_23244,N_22917,N_22649);
and U23245 (N_23245,N_22527,N_22608);
nor U23246 (N_23246,N_22879,N_22977);
nand U23247 (N_23247,N_22514,N_22885);
or U23248 (N_23248,N_22988,N_22557);
xnor U23249 (N_23249,N_22531,N_23084);
nor U23250 (N_23250,N_22506,N_22929);
nand U23251 (N_23251,N_22984,N_22926);
xor U23252 (N_23252,N_22986,N_22672);
and U23253 (N_23253,N_23002,N_23068);
nor U23254 (N_23254,N_22686,N_22854);
nand U23255 (N_23255,N_22817,N_22657);
or U23256 (N_23256,N_23027,N_22969);
and U23257 (N_23257,N_22685,N_22535);
or U23258 (N_23258,N_23117,N_22612);
xor U23259 (N_23259,N_22632,N_22566);
xor U23260 (N_23260,N_22983,N_22855);
or U23261 (N_23261,N_22806,N_22613);
and U23262 (N_23262,N_22716,N_23105);
nand U23263 (N_23263,N_23029,N_22552);
xnor U23264 (N_23264,N_23032,N_22664);
nor U23265 (N_23265,N_22532,N_22503);
nor U23266 (N_23266,N_22634,N_22696);
xnor U23267 (N_23267,N_22954,N_22782);
xnor U23268 (N_23268,N_23036,N_22920);
nand U23269 (N_23269,N_22739,N_22590);
and U23270 (N_23270,N_22897,N_22714);
or U23271 (N_23271,N_23110,N_22860);
or U23272 (N_23272,N_22512,N_23008);
nor U23273 (N_23273,N_22694,N_23023);
nor U23274 (N_23274,N_22980,N_22848);
or U23275 (N_23275,N_22768,N_22811);
and U23276 (N_23276,N_23119,N_22538);
or U23277 (N_23277,N_22944,N_22927);
nor U23278 (N_23278,N_22907,N_22742);
and U23279 (N_23279,N_23067,N_22683);
nor U23280 (N_23280,N_22526,N_22849);
nor U23281 (N_23281,N_23098,N_22721);
or U23282 (N_23282,N_22658,N_22999);
and U23283 (N_23283,N_22591,N_22654);
and U23284 (N_23284,N_22541,N_22595);
or U23285 (N_23285,N_23003,N_22834);
nor U23286 (N_23286,N_22760,N_22546);
nor U23287 (N_23287,N_22726,N_22539);
and U23288 (N_23288,N_22500,N_22922);
and U23289 (N_23289,N_22947,N_22942);
and U23290 (N_23290,N_22906,N_23018);
nor U23291 (N_23291,N_22887,N_22646);
nor U23292 (N_23292,N_22787,N_23059);
nand U23293 (N_23293,N_22754,N_22912);
nand U23294 (N_23294,N_23045,N_22560);
or U23295 (N_23295,N_22682,N_22617);
xnor U23296 (N_23296,N_22765,N_22970);
nand U23297 (N_23297,N_22790,N_22735);
nor U23298 (N_23298,N_22693,N_22890);
xor U23299 (N_23299,N_22810,N_22771);
nand U23300 (N_23300,N_22837,N_22989);
nand U23301 (N_23301,N_22689,N_22673);
or U23302 (N_23302,N_22931,N_23097);
xnor U23303 (N_23303,N_23107,N_23047);
or U23304 (N_23304,N_23016,N_22867);
or U23305 (N_23305,N_22807,N_22842);
nor U23306 (N_23306,N_22777,N_22799);
and U23307 (N_23307,N_22618,N_22896);
nand U23308 (N_23308,N_22668,N_22611);
nor U23309 (N_23309,N_22892,N_22757);
or U23310 (N_23310,N_22780,N_22518);
or U23311 (N_23311,N_22859,N_22852);
nor U23312 (N_23312,N_22728,N_22976);
and U23313 (N_23313,N_23020,N_23049);
nor U23314 (N_23314,N_23075,N_23006);
xnor U23315 (N_23315,N_22916,N_23090);
xnor U23316 (N_23316,N_22801,N_22899);
and U23317 (N_23317,N_22975,N_22504);
nand U23318 (N_23318,N_22792,N_22808);
or U23319 (N_23319,N_22653,N_23078);
nand U23320 (N_23320,N_22838,N_22515);
nor U23321 (N_23321,N_22620,N_22863);
nor U23322 (N_23322,N_23005,N_22812);
xor U23323 (N_23323,N_22905,N_22554);
and U23324 (N_23324,N_22940,N_22756);
nor U23325 (N_23325,N_23122,N_22966);
nor U23326 (N_23326,N_22601,N_22889);
and U23327 (N_23327,N_22641,N_22706);
xnor U23328 (N_23328,N_22676,N_22913);
or U23329 (N_23329,N_22776,N_22864);
xnor U23330 (N_23330,N_22866,N_22764);
nor U23331 (N_23331,N_23051,N_22659);
xnor U23332 (N_23332,N_22705,N_22615);
nor U23333 (N_23333,N_23063,N_22625);
and U23334 (N_23334,N_23121,N_22558);
nor U23335 (N_23335,N_22961,N_22816);
xor U23336 (N_23336,N_22581,N_22647);
and U23337 (N_23337,N_22671,N_22772);
or U23338 (N_23338,N_23120,N_23085);
and U23339 (N_23339,N_23014,N_22583);
nand U23340 (N_23340,N_22895,N_23000);
nand U23341 (N_23341,N_22832,N_22730);
and U23342 (N_23342,N_22592,N_22827);
and U23343 (N_23343,N_23103,N_22957);
nor U23344 (N_23344,N_22691,N_22797);
nor U23345 (N_23345,N_22865,N_22642);
and U23346 (N_23346,N_22990,N_22717);
nand U23347 (N_23347,N_22914,N_22858);
xnor U23348 (N_23348,N_22600,N_22871);
nor U23349 (N_23349,N_22828,N_23100);
or U23350 (N_23350,N_22545,N_22713);
nor U23351 (N_23351,N_22924,N_22580);
nor U23352 (N_23352,N_23091,N_22687);
xor U23353 (N_23353,N_22809,N_22656);
xnor U23354 (N_23354,N_22938,N_23102);
nand U23355 (N_23355,N_22537,N_22839);
nand U23356 (N_23356,N_23024,N_23039);
nand U23357 (N_23357,N_22619,N_22870);
nor U23358 (N_23358,N_22544,N_22994);
and U23359 (N_23359,N_22948,N_23038);
nor U23360 (N_23360,N_22570,N_22844);
and U23361 (N_23361,N_22520,N_23019);
nor U23362 (N_23362,N_23083,N_22690);
xnor U23363 (N_23363,N_22821,N_22987);
nand U23364 (N_23364,N_23013,N_22998);
and U23365 (N_23365,N_22911,N_22587);
nor U23366 (N_23366,N_22610,N_22824);
nand U23367 (N_23367,N_22829,N_22820);
nor U23368 (N_23368,N_22919,N_22953);
xor U23369 (N_23369,N_22737,N_22593);
nor U23370 (N_23370,N_22585,N_23004);
and U23371 (N_23371,N_23011,N_22542);
or U23372 (N_23372,N_23116,N_22563);
xor U23373 (N_23373,N_22769,N_23118);
and U23374 (N_23374,N_23086,N_22525);
or U23375 (N_23375,N_22753,N_23055);
or U23376 (N_23376,N_22789,N_22729);
xor U23377 (N_23377,N_22697,N_22579);
nor U23378 (N_23378,N_22553,N_22556);
and U23379 (N_23379,N_22971,N_22751);
nand U23380 (N_23380,N_22869,N_22715);
and U23381 (N_23381,N_22523,N_22851);
nand U23382 (N_23382,N_22630,N_22875);
nor U23383 (N_23383,N_22663,N_23070);
nand U23384 (N_23384,N_23088,N_23099);
and U23385 (N_23385,N_22804,N_23111);
and U23386 (N_23386,N_22519,N_22534);
and U23387 (N_23387,N_22586,N_22965);
and U23388 (N_23388,N_23060,N_23043);
nand U23389 (N_23389,N_22725,N_22840);
xnor U23390 (N_23390,N_22701,N_23054);
and U23391 (N_23391,N_22678,N_22815);
or U23392 (N_23392,N_22631,N_23058);
xnor U23393 (N_23393,N_22643,N_22935);
or U23394 (N_23394,N_22567,N_22718);
and U23395 (N_23395,N_22798,N_22972);
or U23396 (N_23396,N_23021,N_22800);
or U23397 (N_23397,N_22603,N_22952);
nand U23398 (N_23398,N_22624,N_22501);
nand U23399 (N_23399,N_22622,N_23124);
xor U23400 (N_23400,N_22786,N_22562);
nor U23401 (N_23401,N_23101,N_22670);
xnor U23402 (N_23402,N_22995,N_23046);
nor U23403 (N_23403,N_22733,N_22762);
nand U23404 (N_23404,N_23001,N_22928);
or U23405 (N_23405,N_22645,N_22744);
nor U23406 (N_23406,N_23093,N_22589);
nor U23407 (N_23407,N_22767,N_22749);
xnor U23408 (N_23408,N_22877,N_23062);
nand U23409 (N_23409,N_22564,N_22596);
xnor U23410 (N_23410,N_22943,N_22761);
or U23411 (N_23411,N_22712,N_22991);
or U23412 (N_23412,N_22933,N_22661);
and U23413 (N_23413,N_22530,N_23082);
and U23414 (N_23414,N_22551,N_22727);
and U23415 (N_23415,N_22708,N_23089);
nand U23416 (N_23416,N_22750,N_22918);
nand U23417 (N_23417,N_22888,N_22748);
nand U23418 (N_23418,N_22680,N_22960);
nand U23419 (N_23419,N_23095,N_22509);
xor U23420 (N_23420,N_22992,N_22910);
nand U23421 (N_23421,N_23074,N_22588);
or U23422 (N_23422,N_23079,N_22758);
and U23423 (N_23423,N_22549,N_23081);
or U23424 (N_23424,N_22703,N_23108);
and U23425 (N_23425,N_23092,N_22826);
nor U23426 (N_23426,N_22561,N_22688);
and U23427 (N_23427,N_23112,N_23025);
or U23428 (N_23428,N_22968,N_22575);
or U23429 (N_23429,N_22903,N_22628);
nor U23430 (N_23430,N_22719,N_23076);
or U23431 (N_23431,N_22665,N_22785);
or U23432 (N_23432,N_22695,N_22803);
nand U23433 (N_23433,N_22746,N_22946);
nand U23434 (N_23434,N_22825,N_22766);
xor U23435 (N_23435,N_22699,N_23087);
nand U23436 (N_23436,N_22904,N_22862);
or U23437 (N_23437,N_22872,N_22600);
nor U23438 (N_23438,N_22821,N_22549);
and U23439 (N_23439,N_22673,N_23106);
xor U23440 (N_23440,N_22672,N_22507);
or U23441 (N_23441,N_22669,N_22889);
or U23442 (N_23442,N_22524,N_22832);
nand U23443 (N_23443,N_23114,N_22825);
nor U23444 (N_23444,N_22671,N_23078);
and U23445 (N_23445,N_22740,N_22624);
and U23446 (N_23446,N_22760,N_22713);
xnor U23447 (N_23447,N_22580,N_22991);
or U23448 (N_23448,N_22554,N_23010);
nand U23449 (N_23449,N_22589,N_22947);
xnor U23450 (N_23450,N_22779,N_22598);
nor U23451 (N_23451,N_22574,N_22851);
nor U23452 (N_23452,N_22537,N_23005);
nand U23453 (N_23453,N_22715,N_22758);
or U23454 (N_23454,N_23054,N_23100);
nand U23455 (N_23455,N_22942,N_23119);
or U23456 (N_23456,N_22813,N_22647);
nand U23457 (N_23457,N_23048,N_23019);
and U23458 (N_23458,N_22688,N_22525);
nor U23459 (N_23459,N_22819,N_22615);
nor U23460 (N_23460,N_23074,N_22537);
xor U23461 (N_23461,N_22579,N_23005);
xor U23462 (N_23462,N_22954,N_22993);
nand U23463 (N_23463,N_22562,N_23059);
or U23464 (N_23464,N_22813,N_22913);
xor U23465 (N_23465,N_22720,N_22937);
nand U23466 (N_23466,N_22729,N_22812);
and U23467 (N_23467,N_22615,N_22648);
nand U23468 (N_23468,N_22615,N_22574);
and U23469 (N_23469,N_22800,N_22649);
or U23470 (N_23470,N_23080,N_22562);
and U23471 (N_23471,N_23021,N_23085);
or U23472 (N_23472,N_22894,N_22757);
nand U23473 (N_23473,N_22760,N_22522);
nor U23474 (N_23474,N_22645,N_23085);
nand U23475 (N_23475,N_22851,N_22818);
and U23476 (N_23476,N_22970,N_22636);
and U23477 (N_23477,N_22591,N_22864);
nor U23478 (N_23478,N_23008,N_23079);
nor U23479 (N_23479,N_22727,N_22703);
xor U23480 (N_23480,N_23096,N_22558);
or U23481 (N_23481,N_22829,N_22554);
or U23482 (N_23482,N_22613,N_22778);
and U23483 (N_23483,N_22550,N_22871);
nand U23484 (N_23484,N_23026,N_22854);
xor U23485 (N_23485,N_22835,N_22749);
or U23486 (N_23486,N_22997,N_22831);
or U23487 (N_23487,N_22678,N_23085);
and U23488 (N_23488,N_22887,N_22663);
nor U23489 (N_23489,N_23000,N_22994);
nor U23490 (N_23490,N_22625,N_22728);
xor U23491 (N_23491,N_22699,N_22781);
xor U23492 (N_23492,N_23011,N_22640);
nand U23493 (N_23493,N_22881,N_22507);
xnor U23494 (N_23494,N_22566,N_23094);
nand U23495 (N_23495,N_22774,N_22773);
nand U23496 (N_23496,N_22925,N_22641);
nand U23497 (N_23497,N_23095,N_22872);
or U23498 (N_23498,N_22729,N_22945);
and U23499 (N_23499,N_22958,N_22734);
xnor U23500 (N_23500,N_22600,N_23064);
nand U23501 (N_23501,N_23106,N_22604);
or U23502 (N_23502,N_22740,N_23036);
xnor U23503 (N_23503,N_22586,N_22835);
xor U23504 (N_23504,N_22706,N_22766);
nor U23505 (N_23505,N_23023,N_22843);
nor U23506 (N_23506,N_22740,N_22958);
nor U23507 (N_23507,N_22686,N_22889);
xor U23508 (N_23508,N_22535,N_22788);
nand U23509 (N_23509,N_22543,N_22963);
nand U23510 (N_23510,N_22643,N_22783);
xor U23511 (N_23511,N_22694,N_22912);
xnor U23512 (N_23512,N_22574,N_22772);
nor U23513 (N_23513,N_22592,N_22697);
xnor U23514 (N_23514,N_23119,N_22722);
xnor U23515 (N_23515,N_22953,N_22948);
nor U23516 (N_23516,N_22971,N_22506);
or U23517 (N_23517,N_22850,N_22572);
xnor U23518 (N_23518,N_22607,N_23060);
or U23519 (N_23519,N_22928,N_22511);
xor U23520 (N_23520,N_22737,N_22801);
and U23521 (N_23521,N_22790,N_22785);
or U23522 (N_23522,N_23041,N_22688);
nor U23523 (N_23523,N_22510,N_22978);
and U23524 (N_23524,N_22506,N_22595);
nand U23525 (N_23525,N_22568,N_23121);
nor U23526 (N_23526,N_22768,N_23097);
and U23527 (N_23527,N_22837,N_22794);
xor U23528 (N_23528,N_22526,N_23078);
and U23529 (N_23529,N_22621,N_22925);
and U23530 (N_23530,N_22672,N_23124);
and U23531 (N_23531,N_22861,N_23086);
nor U23532 (N_23532,N_22645,N_22702);
xnor U23533 (N_23533,N_22772,N_22512);
and U23534 (N_23534,N_22565,N_23077);
nand U23535 (N_23535,N_23005,N_22681);
xor U23536 (N_23536,N_23092,N_22583);
or U23537 (N_23537,N_22832,N_23071);
nand U23538 (N_23538,N_22986,N_23113);
or U23539 (N_23539,N_22881,N_23005);
nand U23540 (N_23540,N_22625,N_22586);
nand U23541 (N_23541,N_23119,N_23071);
or U23542 (N_23542,N_22980,N_22669);
or U23543 (N_23543,N_22760,N_22796);
nand U23544 (N_23544,N_23012,N_22957);
and U23545 (N_23545,N_22685,N_23043);
nand U23546 (N_23546,N_22933,N_22797);
xor U23547 (N_23547,N_22821,N_22581);
nand U23548 (N_23548,N_22922,N_22726);
nor U23549 (N_23549,N_22779,N_22687);
or U23550 (N_23550,N_23068,N_22846);
nand U23551 (N_23551,N_22810,N_22870);
or U23552 (N_23552,N_22662,N_22716);
or U23553 (N_23553,N_23044,N_22623);
or U23554 (N_23554,N_23079,N_23058);
nor U23555 (N_23555,N_22997,N_23071);
nor U23556 (N_23556,N_22678,N_22707);
xnor U23557 (N_23557,N_22773,N_22597);
and U23558 (N_23558,N_22828,N_22944);
and U23559 (N_23559,N_22665,N_22948);
xor U23560 (N_23560,N_23051,N_22993);
nor U23561 (N_23561,N_22984,N_22961);
nor U23562 (N_23562,N_23100,N_22767);
or U23563 (N_23563,N_22678,N_22508);
and U23564 (N_23564,N_22515,N_22900);
nor U23565 (N_23565,N_22575,N_22830);
or U23566 (N_23566,N_22543,N_22555);
nor U23567 (N_23567,N_22590,N_22740);
or U23568 (N_23568,N_23011,N_22509);
xnor U23569 (N_23569,N_22891,N_23105);
nand U23570 (N_23570,N_23074,N_22734);
or U23571 (N_23571,N_22768,N_22935);
nor U23572 (N_23572,N_23053,N_22532);
nand U23573 (N_23573,N_22687,N_22549);
and U23574 (N_23574,N_23088,N_23096);
nand U23575 (N_23575,N_22693,N_22560);
nand U23576 (N_23576,N_23115,N_22535);
nor U23577 (N_23577,N_23114,N_22916);
xnor U23578 (N_23578,N_22840,N_22993);
xnor U23579 (N_23579,N_22699,N_23037);
or U23580 (N_23580,N_22776,N_22995);
nor U23581 (N_23581,N_22870,N_23108);
nor U23582 (N_23582,N_22848,N_22873);
nand U23583 (N_23583,N_22956,N_22600);
xnor U23584 (N_23584,N_23027,N_22703);
nor U23585 (N_23585,N_22691,N_22803);
xor U23586 (N_23586,N_22713,N_22765);
nor U23587 (N_23587,N_22628,N_22961);
or U23588 (N_23588,N_22861,N_22737);
nor U23589 (N_23589,N_22774,N_22917);
xnor U23590 (N_23590,N_23033,N_22820);
nand U23591 (N_23591,N_22766,N_22542);
or U23592 (N_23592,N_22809,N_22913);
nor U23593 (N_23593,N_22880,N_22976);
and U23594 (N_23594,N_23036,N_23019);
nand U23595 (N_23595,N_23085,N_22530);
xor U23596 (N_23596,N_22857,N_22522);
nand U23597 (N_23597,N_22640,N_22627);
xnor U23598 (N_23598,N_22728,N_23009);
xor U23599 (N_23599,N_22889,N_22764);
nor U23600 (N_23600,N_23108,N_22942);
xnor U23601 (N_23601,N_22759,N_22591);
or U23602 (N_23602,N_22934,N_22965);
nand U23603 (N_23603,N_22645,N_23070);
and U23604 (N_23604,N_22770,N_22884);
nor U23605 (N_23605,N_23037,N_22807);
or U23606 (N_23606,N_22679,N_22660);
nand U23607 (N_23607,N_22608,N_22681);
or U23608 (N_23608,N_22613,N_23034);
xnor U23609 (N_23609,N_22880,N_22742);
nand U23610 (N_23610,N_23048,N_22533);
xor U23611 (N_23611,N_22800,N_22903);
and U23612 (N_23612,N_22546,N_22619);
and U23613 (N_23613,N_22553,N_22967);
nand U23614 (N_23614,N_23011,N_22827);
nor U23615 (N_23615,N_22531,N_22715);
nor U23616 (N_23616,N_22935,N_22564);
and U23617 (N_23617,N_22665,N_22624);
nand U23618 (N_23618,N_22663,N_22966);
nor U23619 (N_23619,N_22771,N_22532);
nor U23620 (N_23620,N_22538,N_22995);
nor U23621 (N_23621,N_22655,N_22699);
and U23622 (N_23622,N_22940,N_22988);
and U23623 (N_23623,N_22553,N_22785);
nand U23624 (N_23624,N_22735,N_22802);
nor U23625 (N_23625,N_22734,N_22963);
nor U23626 (N_23626,N_22900,N_22643);
nand U23627 (N_23627,N_23012,N_23082);
nor U23628 (N_23628,N_22861,N_22546);
and U23629 (N_23629,N_22916,N_22899);
or U23630 (N_23630,N_22821,N_22722);
xnor U23631 (N_23631,N_23106,N_22945);
xnor U23632 (N_23632,N_22770,N_23112);
and U23633 (N_23633,N_23087,N_23026);
nand U23634 (N_23634,N_23116,N_22501);
and U23635 (N_23635,N_22682,N_22837);
or U23636 (N_23636,N_22598,N_22624);
xor U23637 (N_23637,N_22873,N_22978);
and U23638 (N_23638,N_22633,N_22797);
and U23639 (N_23639,N_22742,N_22735);
and U23640 (N_23640,N_22617,N_22905);
and U23641 (N_23641,N_22725,N_22620);
nor U23642 (N_23642,N_22889,N_22769);
nor U23643 (N_23643,N_23075,N_22828);
nor U23644 (N_23644,N_22581,N_22827);
and U23645 (N_23645,N_23123,N_23028);
nand U23646 (N_23646,N_22518,N_23020);
nor U23647 (N_23647,N_22978,N_23076);
nand U23648 (N_23648,N_23008,N_22810);
or U23649 (N_23649,N_23067,N_23075);
xor U23650 (N_23650,N_22955,N_22604);
xnor U23651 (N_23651,N_22867,N_22728);
or U23652 (N_23652,N_22883,N_23099);
xor U23653 (N_23653,N_22599,N_22678);
nor U23654 (N_23654,N_22799,N_22534);
nor U23655 (N_23655,N_23124,N_22816);
nor U23656 (N_23656,N_22858,N_22957);
and U23657 (N_23657,N_22543,N_22613);
nor U23658 (N_23658,N_22708,N_22884);
nand U23659 (N_23659,N_22990,N_23009);
or U23660 (N_23660,N_22765,N_23008);
and U23661 (N_23661,N_22731,N_22985);
nor U23662 (N_23662,N_23112,N_22871);
and U23663 (N_23663,N_22951,N_23122);
and U23664 (N_23664,N_22817,N_22611);
nor U23665 (N_23665,N_22576,N_23007);
nand U23666 (N_23666,N_23059,N_22917);
and U23667 (N_23667,N_22716,N_22981);
nand U23668 (N_23668,N_22658,N_22979);
or U23669 (N_23669,N_22924,N_23003);
or U23670 (N_23670,N_23058,N_22811);
nand U23671 (N_23671,N_22826,N_22865);
or U23672 (N_23672,N_22588,N_23079);
nand U23673 (N_23673,N_22979,N_23061);
and U23674 (N_23674,N_22704,N_23094);
nor U23675 (N_23675,N_23024,N_22852);
xnor U23676 (N_23676,N_23051,N_22897);
nand U23677 (N_23677,N_22830,N_22995);
nor U23678 (N_23678,N_22841,N_22684);
or U23679 (N_23679,N_22536,N_22971);
nand U23680 (N_23680,N_22961,N_22922);
xor U23681 (N_23681,N_22859,N_23002);
and U23682 (N_23682,N_22736,N_22863);
nor U23683 (N_23683,N_22666,N_22635);
xnor U23684 (N_23684,N_22864,N_22799);
xnor U23685 (N_23685,N_23069,N_22569);
or U23686 (N_23686,N_22673,N_22720);
nor U23687 (N_23687,N_22881,N_23064);
xnor U23688 (N_23688,N_23106,N_22828);
and U23689 (N_23689,N_22799,N_23084);
or U23690 (N_23690,N_23107,N_22538);
xnor U23691 (N_23691,N_22862,N_23008);
and U23692 (N_23692,N_22840,N_22724);
xor U23693 (N_23693,N_23121,N_23070);
xor U23694 (N_23694,N_22694,N_22948);
xnor U23695 (N_23695,N_22884,N_22632);
nor U23696 (N_23696,N_23117,N_22514);
xnor U23697 (N_23697,N_22520,N_22787);
and U23698 (N_23698,N_22996,N_22598);
and U23699 (N_23699,N_22936,N_23012);
or U23700 (N_23700,N_22979,N_22649);
nand U23701 (N_23701,N_23091,N_23009);
nand U23702 (N_23702,N_22761,N_22800);
nor U23703 (N_23703,N_22911,N_22702);
or U23704 (N_23704,N_23077,N_22688);
or U23705 (N_23705,N_22940,N_23122);
nand U23706 (N_23706,N_22970,N_23020);
nand U23707 (N_23707,N_22925,N_22524);
or U23708 (N_23708,N_22996,N_22621);
or U23709 (N_23709,N_22642,N_23052);
nor U23710 (N_23710,N_22576,N_22525);
nand U23711 (N_23711,N_22900,N_22546);
nor U23712 (N_23712,N_23068,N_22924);
xor U23713 (N_23713,N_22571,N_22572);
nor U23714 (N_23714,N_22565,N_22615);
or U23715 (N_23715,N_22509,N_22582);
xnor U23716 (N_23716,N_23013,N_22756);
nand U23717 (N_23717,N_22933,N_23006);
xnor U23718 (N_23718,N_22651,N_22796);
xor U23719 (N_23719,N_23113,N_22818);
xnor U23720 (N_23720,N_23017,N_22620);
or U23721 (N_23721,N_22698,N_22676);
or U23722 (N_23722,N_23078,N_22525);
and U23723 (N_23723,N_22706,N_23118);
and U23724 (N_23724,N_22938,N_22640);
or U23725 (N_23725,N_22794,N_22871);
or U23726 (N_23726,N_22520,N_23033);
and U23727 (N_23727,N_23117,N_22943);
xor U23728 (N_23728,N_22557,N_22620);
or U23729 (N_23729,N_23075,N_22621);
or U23730 (N_23730,N_22609,N_22528);
xnor U23731 (N_23731,N_23033,N_22841);
or U23732 (N_23732,N_22553,N_23045);
or U23733 (N_23733,N_22604,N_23101);
nor U23734 (N_23734,N_23043,N_22540);
xor U23735 (N_23735,N_22745,N_22842);
xnor U23736 (N_23736,N_22912,N_22798);
or U23737 (N_23737,N_22709,N_22972);
xor U23738 (N_23738,N_22653,N_23091);
xor U23739 (N_23739,N_23037,N_22733);
or U23740 (N_23740,N_22955,N_22949);
or U23741 (N_23741,N_23087,N_22685);
and U23742 (N_23742,N_23113,N_22922);
or U23743 (N_23743,N_22775,N_22951);
or U23744 (N_23744,N_22908,N_22989);
or U23745 (N_23745,N_22626,N_22739);
or U23746 (N_23746,N_22676,N_22969);
nand U23747 (N_23747,N_22552,N_23116);
and U23748 (N_23748,N_22935,N_22850);
and U23749 (N_23749,N_22548,N_23100);
or U23750 (N_23750,N_23417,N_23257);
and U23751 (N_23751,N_23696,N_23463);
nor U23752 (N_23752,N_23333,N_23379);
nor U23753 (N_23753,N_23337,N_23433);
nor U23754 (N_23754,N_23564,N_23625);
nor U23755 (N_23755,N_23423,N_23161);
nor U23756 (N_23756,N_23348,N_23632);
nand U23757 (N_23757,N_23542,N_23387);
or U23758 (N_23758,N_23631,N_23197);
nor U23759 (N_23759,N_23363,N_23732);
xnor U23760 (N_23760,N_23331,N_23521);
and U23761 (N_23761,N_23226,N_23309);
xnor U23762 (N_23762,N_23425,N_23687);
xor U23763 (N_23763,N_23454,N_23413);
nor U23764 (N_23764,N_23541,N_23357);
or U23765 (N_23765,N_23483,N_23138);
or U23766 (N_23766,N_23285,N_23234);
nand U23767 (N_23767,N_23182,N_23551);
or U23768 (N_23768,N_23730,N_23432);
and U23769 (N_23769,N_23271,N_23195);
or U23770 (N_23770,N_23633,N_23262);
and U23771 (N_23771,N_23471,N_23382);
nand U23772 (N_23772,N_23470,N_23737);
xnor U23773 (N_23773,N_23573,N_23278);
xor U23774 (N_23774,N_23735,N_23682);
xor U23775 (N_23775,N_23476,N_23544);
xnor U23776 (N_23776,N_23281,N_23220);
and U23777 (N_23777,N_23604,N_23709);
or U23778 (N_23778,N_23509,N_23608);
xor U23779 (N_23779,N_23702,N_23232);
nand U23780 (N_23780,N_23666,N_23670);
nand U23781 (N_23781,N_23508,N_23402);
xnor U23782 (N_23782,N_23334,N_23660);
and U23783 (N_23783,N_23571,N_23319);
xnor U23784 (N_23784,N_23200,N_23500);
xnor U23785 (N_23785,N_23684,N_23364);
xnor U23786 (N_23786,N_23403,N_23704);
or U23787 (N_23787,N_23170,N_23388);
and U23788 (N_23788,N_23540,N_23489);
or U23789 (N_23789,N_23506,N_23229);
nand U23790 (N_23790,N_23661,N_23318);
and U23791 (N_23791,N_23261,N_23703);
or U23792 (N_23792,N_23437,N_23241);
nor U23793 (N_23793,N_23305,N_23194);
and U23794 (N_23794,N_23673,N_23301);
and U23795 (N_23795,N_23743,N_23649);
or U23796 (N_23796,N_23204,N_23466);
and U23797 (N_23797,N_23383,N_23130);
and U23798 (N_23798,N_23600,N_23510);
nand U23799 (N_23799,N_23662,N_23280);
or U23800 (N_23800,N_23745,N_23712);
and U23801 (N_23801,N_23239,N_23727);
nand U23802 (N_23802,N_23157,N_23208);
xor U23803 (N_23803,N_23595,N_23691);
or U23804 (N_23804,N_23493,N_23519);
xnor U23805 (N_23805,N_23332,N_23537);
nand U23806 (N_23806,N_23697,N_23335);
xnor U23807 (N_23807,N_23457,N_23160);
nand U23808 (N_23808,N_23135,N_23602);
nand U23809 (N_23809,N_23645,N_23336);
and U23810 (N_23810,N_23441,N_23327);
xor U23811 (N_23811,N_23590,N_23439);
nor U23812 (N_23812,N_23680,N_23693);
and U23813 (N_23813,N_23251,N_23249);
or U23814 (N_23814,N_23260,N_23446);
nor U23815 (N_23815,N_23424,N_23214);
xor U23816 (N_23816,N_23284,N_23530);
and U23817 (N_23817,N_23412,N_23555);
nand U23818 (N_23818,N_23415,N_23283);
nor U23819 (N_23819,N_23607,N_23381);
nor U23820 (N_23820,N_23270,N_23448);
and U23821 (N_23821,N_23450,N_23287);
xor U23822 (N_23822,N_23611,N_23567);
or U23823 (N_23823,N_23527,N_23654);
xnor U23824 (N_23824,N_23218,N_23546);
xnor U23825 (N_23825,N_23517,N_23198);
or U23826 (N_23826,N_23726,N_23346);
nand U23827 (N_23827,N_23344,N_23235);
xnor U23828 (N_23828,N_23236,N_23657);
and U23829 (N_23829,N_23137,N_23139);
xor U23830 (N_23830,N_23177,N_23227);
nor U23831 (N_23831,N_23626,N_23132);
or U23832 (N_23832,N_23591,N_23614);
nor U23833 (N_23833,N_23409,N_23186);
or U23834 (N_23834,N_23523,N_23487);
nand U23835 (N_23835,N_23584,N_23349);
or U23836 (N_23836,N_23223,N_23185);
nand U23837 (N_23837,N_23390,N_23520);
nand U23838 (N_23838,N_23462,N_23216);
or U23839 (N_23839,N_23438,N_23242);
nor U23840 (N_23840,N_23534,N_23414);
or U23841 (N_23841,N_23453,N_23426);
and U23842 (N_23842,N_23651,N_23685);
and U23843 (N_23843,N_23589,N_23265);
nor U23844 (N_23844,N_23557,N_23295);
and U23845 (N_23845,N_23686,N_23293);
nand U23846 (N_23846,N_23711,N_23360);
or U23847 (N_23847,N_23716,N_23428);
nand U23848 (N_23848,N_23744,N_23164);
xor U23849 (N_23849,N_23165,N_23386);
nor U23850 (N_23850,N_23345,N_23581);
and U23851 (N_23851,N_23738,N_23543);
and U23852 (N_23852,N_23374,N_23436);
or U23853 (N_23853,N_23376,N_23256);
and U23854 (N_23854,N_23692,N_23134);
xor U23855 (N_23855,N_23701,N_23695);
nor U23856 (N_23856,N_23275,N_23313);
xor U23857 (N_23857,N_23554,N_23449);
and U23858 (N_23858,N_23330,N_23230);
nor U23859 (N_23859,N_23320,N_23396);
nand U23860 (N_23860,N_23443,N_23529);
nor U23861 (N_23861,N_23380,N_23365);
xor U23862 (N_23862,N_23733,N_23372);
or U23863 (N_23863,N_23707,N_23391);
nand U23864 (N_23864,N_23142,N_23596);
nor U23865 (N_23865,N_23511,N_23178);
nand U23866 (N_23866,N_23491,N_23621);
nor U23867 (N_23867,N_23585,N_23741);
nand U23868 (N_23868,N_23310,N_23538);
nand U23869 (N_23869,N_23269,N_23407);
or U23870 (N_23870,N_23141,N_23484);
xnor U23871 (N_23871,N_23525,N_23634);
or U23872 (N_23872,N_23617,N_23153);
nand U23873 (N_23873,N_23311,N_23723);
xnor U23874 (N_23874,N_23665,N_23427);
xor U23875 (N_23875,N_23445,N_23576);
nand U23876 (N_23876,N_23146,N_23338);
nor U23877 (N_23877,N_23329,N_23627);
nor U23878 (N_23878,N_23145,N_23266);
or U23879 (N_23879,N_23368,N_23370);
xnor U23880 (N_23880,N_23210,N_23375);
or U23881 (N_23881,N_23276,N_23340);
nand U23882 (N_23882,N_23347,N_23440);
or U23883 (N_23883,N_23480,N_23312);
or U23884 (N_23884,N_23181,N_23469);
xor U23885 (N_23885,N_23549,N_23400);
or U23886 (N_23886,N_23558,N_23688);
and U23887 (N_23887,N_23361,N_23201);
or U23888 (N_23888,N_23486,N_23175);
or U23889 (N_23889,N_23434,N_23147);
and U23890 (N_23890,N_23568,N_23352);
and U23891 (N_23891,N_23189,N_23638);
nor U23892 (N_23892,N_23129,N_23421);
nand U23893 (N_23893,N_23292,N_23563);
xnor U23894 (N_23894,N_23255,N_23490);
xor U23895 (N_23895,N_23667,N_23213);
and U23896 (N_23896,N_23501,N_23675);
nand U23897 (N_23897,N_23233,N_23565);
and U23898 (N_23898,N_23246,N_23622);
nor U23899 (N_23899,N_23158,N_23636);
xor U23900 (N_23900,N_23353,N_23315);
nand U23901 (N_23901,N_23384,N_23629);
or U23902 (N_23902,N_23492,N_23222);
or U23903 (N_23903,N_23259,N_23288);
or U23904 (N_23904,N_23274,N_23663);
xor U23905 (N_23905,N_23190,N_23533);
and U23906 (N_23906,N_23588,N_23184);
nor U23907 (N_23907,N_23307,N_23286);
nor U23908 (N_23908,N_23273,N_23304);
xnor U23909 (N_23909,N_23465,N_23643);
xnor U23910 (N_23910,N_23512,N_23639);
nor U23911 (N_23911,N_23362,N_23640);
xor U23912 (N_23912,N_23624,N_23513);
and U23913 (N_23913,N_23650,N_23444);
and U23914 (N_23914,N_23211,N_23290);
and U23915 (N_23915,N_23479,N_23623);
nand U23916 (N_23916,N_23430,N_23408);
nor U23917 (N_23917,N_23299,N_23397);
xnor U23918 (N_23918,N_23166,N_23528);
nor U23919 (N_23919,N_23628,N_23455);
and U23920 (N_23920,N_23326,N_23221);
xor U23921 (N_23921,N_23597,N_23570);
and U23922 (N_23922,N_23442,N_23272);
xor U23923 (N_23923,N_23503,N_23323);
nor U23924 (N_23924,N_23258,N_23163);
nand U23925 (N_23925,N_23725,N_23676);
xnor U23926 (N_23926,N_23172,N_23136);
and U23927 (N_23927,N_23267,N_23196);
or U23928 (N_23928,N_23277,N_23392);
and U23929 (N_23929,N_23524,N_23206);
nor U23930 (N_23930,N_23722,N_23395);
nand U23931 (N_23931,N_23168,N_23366);
or U23932 (N_23932,N_23404,N_23742);
nor U23933 (N_23933,N_23244,N_23672);
nand U23934 (N_23934,N_23664,N_23658);
nand U23935 (N_23935,N_23612,N_23642);
or U23936 (N_23936,N_23322,N_23193);
nor U23937 (N_23937,N_23593,N_23599);
nor U23938 (N_23938,N_23736,N_23248);
nor U23939 (N_23939,N_23720,N_23202);
xnor U23940 (N_23940,N_23561,N_23250);
xnor U23941 (N_23941,N_23552,N_23389);
nor U23942 (N_23942,N_23747,N_23418);
or U23943 (N_23943,N_23497,N_23681);
or U23944 (N_23944,N_23653,N_23156);
or U23945 (N_23945,N_23126,N_23183);
and U23946 (N_23946,N_23398,N_23580);
or U23947 (N_23947,N_23212,N_23586);
nor U23948 (N_23948,N_23566,N_23149);
nor U23949 (N_23949,N_23171,N_23646);
or U23950 (N_23950,N_23494,N_23191);
and U23951 (N_23951,N_23203,N_23536);
and U23952 (N_23952,N_23671,N_23679);
or U23953 (N_23953,N_23648,N_23475);
xnor U23954 (N_23954,N_23488,N_23637);
or U23955 (N_23955,N_23620,N_23578);
or U23956 (N_23956,N_23710,N_23616);
or U23957 (N_23957,N_23678,N_23668);
or U23958 (N_23958,N_23207,N_23209);
or U23959 (N_23959,N_23459,N_23263);
nor U23960 (N_23960,N_23504,N_23467);
nor U23961 (N_23961,N_23308,N_23472);
nand U23962 (N_23962,N_23302,N_23174);
nand U23963 (N_23963,N_23297,N_23169);
xor U23964 (N_23964,N_23393,N_23447);
and U23965 (N_23965,N_23708,N_23435);
xnor U23966 (N_23966,N_23458,N_23609);
nand U23967 (N_23967,N_23635,N_23594);
and U23968 (N_23968,N_23245,N_23495);
nor U23969 (N_23969,N_23575,N_23300);
xor U23970 (N_23970,N_23547,N_23545);
nand U23971 (N_23971,N_23582,N_23539);
and U23972 (N_23972,N_23477,N_23577);
or U23973 (N_23973,N_23401,N_23705);
nand U23974 (N_23974,N_23531,N_23507);
nor U23975 (N_23975,N_23535,N_23592);
nand U23976 (N_23976,N_23151,N_23155);
xor U23977 (N_23977,N_23188,N_23740);
and U23978 (N_23978,N_23548,N_23152);
or U23979 (N_23979,N_23268,N_23369);
xnor U23980 (N_23980,N_23606,N_23598);
or U23981 (N_23981,N_23176,N_23502);
nand U23982 (N_23982,N_23394,N_23748);
nand U23983 (N_23983,N_23526,N_23131);
xnor U23984 (N_23984,N_23619,N_23127);
or U23985 (N_23985,N_23514,N_23410);
nor U23986 (N_23986,N_23464,N_23367);
and U23987 (N_23987,N_23583,N_23419);
nor U23988 (N_23988,N_23719,N_23144);
xnor U23989 (N_23989,N_23699,N_23734);
nand U23990 (N_23990,N_23405,N_23133);
nand U23991 (N_23991,N_23238,N_23496);
nand U23992 (N_23992,N_23505,N_23339);
xor U23993 (N_23993,N_23731,N_23532);
and U23994 (N_23994,N_23150,N_23677);
or U23995 (N_23995,N_23406,N_23187);
or U23996 (N_23996,N_23247,N_23478);
xnor U23997 (N_23997,N_23644,N_23473);
nand U23998 (N_23998,N_23159,N_23219);
or U23999 (N_23999,N_23615,N_23328);
xnor U24000 (N_24000,N_23253,N_23714);
nand U24001 (N_24001,N_23377,N_23314);
or U24002 (N_24002,N_23237,N_23556);
nor U24003 (N_24003,N_23498,N_23350);
nor U24004 (N_24004,N_23515,N_23729);
or U24005 (N_24005,N_23516,N_23356);
and U24006 (N_24006,N_23264,N_23562);
nor U24007 (N_24007,N_23282,N_23354);
and U24008 (N_24008,N_23154,N_23343);
xnor U24009 (N_24009,N_23140,N_23294);
and U24010 (N_24010,N_23579,N_23358);
nor U24011 (N_24011,N_23572,N_23630);
and U24012 (N_24012,N_23205,N_23179);
nand U24013 (N_24013,N_23128,N_23451);
nor U24014 (N_24014,N_23618,N_23173);
xor U24015 (N_24015,N_23610,N_23698);
and U24016 (N_24016,N_23228,N_23192);
or U24017 (N_24017,N_23669,N_23303);
or U24018 (N_24018,N_23298,N_23291);
or U24019 (N_24019,N_23550,N_23605);
or U24020 (N_24020,N_23252,N_23706);
nand U24021 (N_24021,N_23746,N_23215);
nor U24022 (N_24022,N_23167,N_23721);
and U24023 (N_24023,N_23431,N_23199);
nor U24024 (N_24024,N_23143,N_23321);
or U24025 (N_24025,N_23656,N_23341);
xor U24026 (N_24026,N_23689,N_23385);
nor U24027 (N_24027,N_23728,N_23217);
nor U24028 (N_24028,N_23652,N_23713);
and U24029 (N_24029,N_23231,N_23317);
xnor U24030 (N_24030,N_23422,N_23162);
xnor U24031 (N_24031,N_23522,N_23456);
nand U24032 (N_24032,N_23518,N_23243);
nand U24033 (N_24033,N_23420,N_23460);
xor U24034 (N_24034,N_23461,N_23254);
xor U24035 (N_24035,N_23683,N_23749);
xnor U24036 (N_24036,N_23411,N_23371);
nand U24037 (N_24037,N_23481,N_23342);
or U24038 (N_24038,N_23724,N_23378);
and U24039 (N_24039,N_23373,N_23125);
and U24040 (N_24040,N_23452,N_23659);
or U24041 (N_24041,N_23148,N_23324);
and U24042 (N_24042,N_23482,N_23224);
nor U24043 (N_24043,N_23474,N_23306);
and U24044 (N_24044,N_23718,N_23655);
and U24045 (N_24045,N_23296,N_23700);
or U24046 (N_24046,N_23553,N_23351);
and U24047 (N_24047,N_23499,N_23574);
nor U24048 (N_24048,N_23316,N_23674);
nand U24049 (N_24049,N_23429,N_23240);
and U24050 (N_24050,N_23601,N_23569);
xor U24051 (N_24051,N_23641,N_23355);
nor U24052 (N_24052,N_23225,N_23416);
nor U24053 (N_24053,N_23180,N_23325);
nand U24054 (N_24054,N_23559,N_23289);
nand U24055 (N_24055,N_23399,N_23613);
and U24056 (N_24056,N_23587,N_23279);
xnor U24057 (N_24057,N_23694,N_23647);
xnor U24058 (N_24058,N_23485,N_23468);
nand U24059 (N_24059,N_23717,N_23359);
or U24060 (N_24060,N_23560,N_23715);
and U24061 (N_24061,N_23690,N_23739);
nand U24062 (N_24062,N_23603,N_23218);
xnor U24063 (N_24063,N_23725,N_23330);
nor U24064 (N_24064,N_23334,N_23224);
nor U24065 (N_24065,N_23561,N_23652);
and U24066 (N_24066,N_23439,N_23139);
and U24067 (N_24067,N_23301,N_23305);
or U24068 (N_24068,N_23467,N_23430);
xor U24069 (N_24069,N_23300,N_23447);
and U24070 (N_24070,N_23727,N_23479);
or U24071 (N_24071,N_23354,N_23238);
nor U24072 (N_24072,N_23672,N_23701);
nor U24073 (N_24073,N_23482,N_23151);
nand U24074 (N_24074,N_23339,N_23693);
or U24075 (N_24075,N_23398,N_23331);
nand U24076 (N_24076,N_23584,N_23744);
nor U24077 (N_24077,N_23687,N_23476);
xnor U24078 (N_24078,N_23356,N_23255);
or U24079 (N_24079,N_23617,N_23414);
xor U24080 (N_24080,N_23323,N_23368);
nand U24081 (N_24081,N_23480,N_23587);
xor U24082 (N_24082,N_23611,N_23159);
or U24083 (N_24083,N_23732,N_23514);
and U24084 (N_24084,N_23399,N_23489);
or U24085 (N_24085,N_23395,N_23719);
xor U24086 (N_24086,N_23134,N_23641);
or U24087 (N_24087,N_23160,N_23552);
and U24088 (N_24088,N_23429,N_23250);
nor U24089 (N_24089,N_23257,N_23584);
or U24090 (N_24090,N_23320,N_23330);
nor U24091 (N_24091,N_23415,N_23692);
nor U24092 (N_24092,N_23284,N_23203);
nand U24093 (N_24093,N_23216,N_23626);
or U24094 (N_24094,N_23503,N_23382);
or U24095 (N_24095,N_23472,N_23352);
nand U24096 (N_24096,N_23564,N_23308);
or U24097 (N_24097,N_23215,N_23503);
nand U24098 (N_24098,N_23559,N_23743);
nand U24099 (N_24099,N_23462,N_23341);
nand U24100 (N_24100,N_23281,N_23435);
xor U24101 (N_24101,N_23422,N_23164);
or U24102 (N_24102,N_23362,N_23150);
or U24103 (N_24103,N_23704,N_23564);
nor U24104 (N_24104,N_23209,N_23642);
nand U24105 (N_24105,N_23477,N_23657);
xnor U24106 (N_24106,N_23736,N_23498);
nor U24107 (N_24107,N_23571,N_23200);
or U24108 (N_24108,N_23430,N_23149);
or U24109 (N_24109,N_23245,N_23415);
xnor U24110 (N_24110,N_23131,N_23192);
nor U24111 (N_24111,N_23306,N_23522);
xor U24112 (N_24112,N_23500,N_23483);
nand U24113 (N_24113,N_23534,N_23284);
or U24114 (N_24114,N_23500,N_23687);
xor U24115 (N_24115,N_23415,N_23473);
and U24116 (N_24116,N_23518,N_23460);
or U24117 (N_24117,N_23667,N_23316);
xnor U24118 (N_24118,N_23172,N_23333);
nand U24119 (N_24119,N_23494,N_23206);
nand U24120 (N_24120,N_23604,N_23154);
nand U24121 (N_24121,N_23349,N_23380);
and U24122 (N_24122,N_23638,N_23630);
nor U24123 (N_24123,N_23697,N_23255);
and U24124 (N_24124,N_23603,N_23501);
and U24125 (N_24125,N_23608,N_23717);
nand U24126 (N_24126,N_23281,N_23249);
nand U24127 (N_24127,N_23402,N_23694);
nand U24128 (N_24128,N_23614,N_23191);
nand U24129 (N_24129,N_23228,N_23579);
nor U24130 (N_24130,N_23702,N_23705);
nor U24131 (N_24131,N_23630,N_23186);
xor U24132 (N_24132,N_23323,N_23272);
nand U24133 (N_24133,N_23267,N_23240);
and U24134 (N_24134,N_23607,N_23727);
and U24135 (N_24135,N_23609,N_23444);
xor U24136 (N_24136,N_23628,N_23427);
nand U24137 (N_24137,N_23385,N_23199);
xnor U24138 (N_24138,N_23381,N_23741);
nor U24139 (N_24139,N_23292,N_23585);
xor U24140 (N_24140,N_23419,N_23718);
and U24141 (N_24141,N_23182,N_23492);
nor U24142 (N_24142,N_23297,N_23210);
xnor U24143 (N_24143,N_23736,N_23429);
xnor U24144 (N_24144,N_23661,N_23239);
and U24145 (N_24145,N_23550,N_23399);
nor U24146 (N_24146,N_23312,N_23180);
and U24147 (N_24147,N_23693,N_23151);
xor U24148 (N_24148,N_23680,N_23398);
xnor U24149 (N_24149,N_23231,N_23742);
nand U24150 (N_24150,N_23490,N_23391);
and U24151 (N_24151,N_23161,N_23488);
and U24152 (N_24152,N_23531,N_23250);
or U24153 (N_24153,N_23155,N_23361);
xnor U24154 (N_24154,N_23331,N_23485);
and U24155 (N_24155,N_23713,N_23536);
nor U24156 (N_24156,N_23625,N_23389);
nand U24157 (N_24157,N_23720,N_23144);
and U24158 (N_24158,N_23716,N_23722);
or U24159 (N_24159,N_23671,N_23477);
nand U24160 (N_24160,N_23352,N_23195);
nor U24161 (N_24161,N_23304,N_23383);
xor U24162 (N_24162,N_23219,N_23671);
and U24163 (N_24163,N_23208,N_23368);
and U24164 (N_24164,N_23498,N_23324);
nand U24165 (N_24165,N_23621,N_23192);
nor U24166 (N_24166,N_23678,N_23574);
and U24167 (N_24167,N_23359,N_23455);
nor U24168 (N_24168,N_23647,N_23158);
xnor U24169 (N_24169,N_23428,N_23425);
xor U24170 (N_24170,N_23728,N_23691);
and U24171 (N_24171,N_23572,N_23736);
and U24172 (N_24172,N_23586,N_23407);
or U24173 (N_24173,N_23467,N_23639);
nor U24174 (N_24174,N_23247,N_23642);
nand U24175 (N_24175,N_23144,N_23600);
and U24176 (N_24176,N_23460,N_23649);
nand U24177 (N_24177,N_23521,N_23214);
xnor U24178 (N_24178,N_23700,N_23462);
and U24179 (N_24179,N_23521,N_23438);
and U24180 (N_24180,N_23389,N_23460);
nor U24181 (N_24181,N_23134,N_23282);
xor U24182 (N_24182,N_23140,N_23551);
and U24183 (N_24183,N_23465,N_23471);
and U24184 (N_24184,N_23154,N_23570);
or U24185 (N_24185,N_23216,N_23292);
nand U24186 (N_24186,N_23653,N_23464);
and U24187 (N_24187,N_23387,N_23718);
xor U24188 (N_24188,N_23275,N_23498);
xor U24189 (N_24189,N_23587,N_23260);
xnor U24190 (N_24190,N_23322,N_23416);
nand U24191 (N_24191,N_23255,N_23334);
nor U24192 (N_24192,N_23151,N_23347);
nor U24193 (N_24193,N_23195,N_23447);
xnor U24194 (N_24194,N_23627,N_23715);
nor U24195 (N_24195,N_23479,N_23322);
or U24196 (N_24196,N_23610,N_23375);
xor U24197 (N_24197,N_23676,N_23514);
xor U24198 (N_24198,N_23410,N_23166);
nand U24199 (N_24199,N_23359,N_23742);
nor U24200 (N_24200,N_23587,N_23253);
nand U24201 (N_24201,N_23691,N_23542);
and U24202 (N_24202,N_23181,N_23689);
or U24203 (N_24203,N_23349,N_23669);
nor U24204 (N_24204,N_23629,N_23734);
xnor U24205 (N_24205,N_23618,N_23716);
nor U24206 (N_24206,N_23341,N_23336);
nand U24207 (N_24207,N_23593,N_23217);
or U24208 (N_24208,N_23598,N_23707);
xor U24209 (N_24209,N_23545,N_23155);
and U24210 (N_24210,N_23285,N_23483);
xor U24211 (N_24211,N_23257,N_23714);
nand U24212 (N_24212,N_23468,N_23448);
or U24213 (N_24213,N_23171,N_23654);
nand U24214 (N_24214,N_23705,N_23471);
xor U24215 (N_24215,N_23281,N_23512);
or U24216 (N_24216,N_23509,N_23219);
or U24217 (N_24217,N_23175,N_23417);
or U24218 (N_24218,N_23578,N_23336);
xnor U24219 (N_24219,N_23596,N_23324);
nor U24220 (N_24220,N_23450,N_23748);
and U24221 (N_24221,N_23618,N_23622);
xor U24222 (N_24222,N_23713,N_23600);
nand U24223 (N_24223,N_23528,N_23162);
xnor U24224 (N_24224,N_23342,N_23353);
xor U24225 (N_24225,N_23716,N_23126);
and U24226 (N_24226,N_23686,N_23314);
or U24227 (N_24227,N_23427,N_23130);
and U24228 (N_24228,N_23633,N_23727);
nand U24229 (N_24229,N_23430,N_23730);
xnor U24230 (N_24230,N_23265,N_23190);
nand U24231 (N_24231,N_23670,N_23194);
nand U24232 (N_24232,N_23544,N_23206);
nor U24233 (N_24233,N_23244,N_23534);
and U24234 (N_24234,N_23371,N_23240);
or U24235 (N_24235,N_23573,N_23667);
nand U24236 (N_24236,N_23347,N_23740);
nand U24237 (N_24237,N_23187,N_23264);
and U24238 (N_24238,N_23361,N_23298);
nand U24239 (N_24239,N_23377,N_23297);
xnor U24240 (N_24240,N_23344,N_23589);
xor U24241 (N_24241,N_23494,N_23468);
and U24242 (N_24242,N_23746,N_23180);
xor U24243 (N_24243,N_23476,N_23490);
xor U24244 (N_24244,N_23330,N_23525);
nand U24245 (N_24245,N_23324,N_23656);
nand U24246 (N_24246,N_23499,N_23539);
nand U24247 (N_24247,N_23524,N_23231);
nor U24248 (N_24248,N_23219,N_23729);
and U24249 (N_24249,N_23253,N_23462);
nand U24250 (N_24250,N_23283,N_23460);
and U24251 (N_24251,N_23628,N_23226);
xor U24252 (N_24252,N_23156,N_23229);
nand U24253 (N_24253,N_23186,N_23724);
or U24254 (N_24254,N_23490,N_23486);
nand U24255 (N_24255,N_23531,N_23413);
nor U24256 (N_24256,N_23265,N_23378);
nand U24257 (N_24257,N_23641,N_23460);
xnor U24258 (N_24258,N_23158,N_23717);
nand U24259 (N_24259,N_23467,N_23572);
nor U24260 (N_24260,N_23460,N_23717);
and U24261 (N_24261,N_23397,N_23240);
nand U24262 (N_24262,N_23483,N_23364);
or U24263 (N_24263,N_23505,N_23642);
xnor U24264 (N_24264,N_23354,N_23385);
nor U24265 (N_24265,N_23257,N_23736);
xor U24266 (N_24266,N_23168,N_23470);
xor U24267 (N_24267,N_23233,N_23390);
xnor U24268 (N_24268,N_23749,N_23725);
and U24269 (N_24269,N_23443,N_23392);
nor U24270 (N_24270,N_23612,N_23524);
or U24271 (N_24271,N_23240,N_23501);
nand U24272 (N_24272,N_23532,N_23435);
nor U24273 (N_24273,N_23280,N_23636);
nor U24274 (N_24274,N_23257,N_23613);
and U24275 (N_24275,N_23126,N_23251);
nor U24276 (N_24276,N_23251,N_23500);
xor U24277 (N_24277,N_23581,N_23609);
nor U24278 (N_24278,N_23190,N_23312);
xnor U24279 (N_24279,N_23725,N_23700);
nand U24280 (N_24280,N_23748,N_23565);
xnor U24281 (N_24281,N_23149,N_23335);
nor U24282 (N_24282,N_23546,N_23177);
nor U24283 (N_24283,N_23737,N_23391);
or U24284 (N_24284,N_23575,N_23680);
xor U24285 (N_24285,N_23315,N_23206);
xor U24286 (N_24286,N_23370,N_23576);
xnor U24287 (N_24287,N_23541,N_23299);
or U24288 (N_24288,N_23657,N_23305);
xnor U24289 (N_24289,N_23606,N_23584);
and U24290 (N_24290,N_23422,N_23191);
and U24291 (N_24291,N_23429,N_23698);
or U24292 (N_24292,N_23689,N_23224);
xnor U24293 (N_24293,N_23379,N_23145);
xnor U24294 (N_24294,N_23146,N_23286);
or U24295 (N_24295,N_23402,N_23256);
nor U24296 (N_24296,N_23481,N_23646);
nor U24297 (N_24297,N_23618,N_23319);
xor U24298 (N_24298,N_23660,N_23332);
nand U24299 (N_24299,N_23483,N_23613);
nor U24300 (N_24300,N_23377,N_23714);
or U24301 (N_24301,N_23171,N_23454);
nor U24302 (N_24302,N_23271,N_23444);
xor U24303 (N_24303,N_23304,N_23465);
xor U24304 (N_24304,N_23598,N_23384);
or U24305 (N_24305,N_23261,N_23151);
or U24306 (N_24306,N_23688,N_23639);
nand U24307 (N_24307,N_23657,N_23532);
nor U24308 (N_24308,N_23204,N_23725);
or U24309 (N_24309,N_23605,N_23604);
nor U24310 (N_24310,N_23719,N_23542);
and U24311 (N_24311,N_23612,N_23510);
nor U24312 (N_24312,N_23366,N_23667);
or U24313 (N_24313,N_23356,N_23543);
xor U24314 (N_24314,N_23600,N_23213);
xnor U24315 (N_24315,N_23226,N_23159);
and U24316 (N_24316,N_23474,N_23642);
xnor U24317 (N_24317,N_23593,N_23304);
nor U24318 (N_24318,N_23173,N_23614);
or U24319 (N_24319,N_23424,N_23194);
or U24320 (N_24320,N_23259,N_23509);
or U24321 (N_24321,N_23297,N_23678);
or U24322 (N_24322,N_23334,N_23155);
nand U24323 (N_24323,N_23423,N_23163);
nand U24324 (N_24324,N_23303,N_23621);
nor U24325 (N_24325,N_23571,N_23185);
nor U24326 (N_24326,N_23607,N_23402);
nor U24327 (N_24327,N_23454,N_23221);
nor U24328 (N_24328,N_23660,N_23280);
or U24329 (N_24329,N_23408,N_23490);
nor U24330 (N_24330,N_23265,N_23632);
or U24331 (N_24331,N_23723,N_23161);
and U24332 (N_24332,N_23386,N_23553);
xnor U24333 (N_24333,N_23564,N_23547);
or U24334 (N_24334,N_23290,N_23665);
xor U24335 (N_24335,N_23136,N_23492);
xnor U24336 (N_24336,N_23192,N_23212);
nor U24337 (N_24337,N_23319,N_23473);
nand U24338 (N_24338,N_23639,N_23286);
nand U24339 (N_24339,N_23175,N_23312);
xor U24340 (N_24340,N_23432,N_23163);
xnor U24341 (N_24341,N_23242,N_23277);
or U24342 (N_24342,N_23298,N_23645);
and U24343 (N_24343,N_23676,N_23334);
or U24344 (N_24344,N_23314,N_23376);
and U24345 (N_24345,N_23354,N_23689);
nand U24346 (N_24346,N_23625,N_23301);
or U24347 (N_24347,N_23136,N_23688);
nand U24348 (N_24348,N_23555,N_23650);
and U24349 (N_24349,N_23347,N_23570);
and U24350 (N_24350,N_23622,N_23652);
nand U24351 (N_24351,N_23586,N_23690);
xor U24352 (N_24352,N_23202,N_23443);
xnor U24353 (N_24353,N_23471,N_23601);
nor U24354 (N_24354,N_23624,N_23255);
nand U24355 (N_24355,N_23375,N_23595);
nand U24356 (N_24356,N_23528,N_23510);
nand U24357 (N_24357,N_23741,N_23147);
and U24358 (N_24358,N_23432,N_23178);
and U24359 (N_24359,N_23403,N_23505);
nor U24360 (N_24360,N_23567,N_23433);
nor U24361 (N_24361,N_23275,N_23207);
and U24362 (N_24362,N_23184,N_23372);
or U24363 (N_24363,N_23650,N_23237);
xor U24364 (N_24364,N_23474,N_23713);
xnor U24365 (N_24365,N_23272,N_23590);
xnor U24366 (N_24366,N_23480,N_23155);
or U24367 (N_24367,N_23749,N_23672);
nand U24368 (N_24368,N_23475,N_23733);
nor U24369 (N_24369,N_23350,N_23712);
nor U24370 (N_24370,N_23708,N_23507);
nor U24371 (N_24371,N_23138,N_23308);
and U24372 (N_24372,N_23223,N_23557);
or U24373 (N_24373,N_23342,N_23627);
nor U24374 (N_24374,N_23406,N_23615);
xor U24375 (N_24375,N_24033,N_23798);
and U24376 (N_24376,N_23916,N_24130);
nor U24377 (N_24377,N_24270,N_23860);
or U24378 (N_24378,N_23779,N_24068);
or U24379 (N_24379,N_24345,N_23787);
nand U24380 (N_24380,N_24312,N_24063);
or U24381 (N_24381,N_24263,N_24249);
nor U24382 (N_24382,N_23876,N_24005);
nor U24383 (N_24383,N_24031,N_24067);
and U24384 (N_24384,N_24051,N_24281);
and U24385 (N_24385,N_24247,N_23941);
nand U24386 (N_24386,N_24208,N_24344);
and U24387 (N_24387,N_24305,N_24350);
or U24388 (N_24388,N_24003,N_23968);
and U24389 (N_24389,N_23899,N_24369);
nor U24390 (N_24390,N_23750,N_24191);
and U24391 (N_24391,N_23915,N_24091);
or U24392 (N_24392,N_23835,N_23818);
xor U24393 (N_24393,N_23811,N_24084);
nor U24394 (N_24394,N_23874,N_24101);
or U24395 (N_24395,N_24062,N_24254);
nor U24396 (N_24396,N_24296,N_24334);
and U24397 (N_24397,N_23998,N_23971);
xnor U24398 (N_24398,N_24363,N_24374);
and U24399 (N_24399,N_24212,N_23973);
nand U24400 (N_24400,N_23913,N_23910);
nor U24401 (N_24401,N_23946,N_24326);
nor U24402 (N_24402,N_23900,N_23799);
nand U24403 (N_24403,N_24322,N_24144);
nand U24404 (N_24404,N_23948,N_24172);
nand U24405 (N_24405,N_24268,N_24100);
nand U24406 (N_24406,N_23830,N_24006);
xnor U24407 (N_24407,N_24331,N_24008);
nand U24408 (N_24408,N_23982,N_23942);
nand U24409 (N_24409,N_23791,N_24346);
and U24410 (N_24410,N_24114,N_24129);
and U24411 (N_24411,N_23962,N_23834);
or U24412 (N_24412,N_24229,N_23863);
nor U24413 (N_24413,N_24121,N_24293);
and U24414 (N_24414,N_24216,N_24366);
and U24415 (N_24415,N_24037,N_24330);
xor U24416 (N_24416,N_24164,N_23979);
and U24417 (N_24417,N_24324,N_24097);
and U24418 (N_24418,N_24303,N_24160);
xor U24419 (N_24419,N_24079,N_23788);
xnor U24420 (N_24420,N_23757,N_24320);
and U24421 (N_24421,N_24155,N_24302);
xor U24422 (N_24422,N_24170,N_24333);
and U24423 (N_24423,N_23786,N_24244);
xnor U24424 (N_24424,N_23954,N_24047);
nor U24425 (N_24425,N_23872,N_24016);
xor U24426 (N_24426,N_24274,N_24202);
and U24427 (N_24427,N_24359,N_23967);
nand U24428 (N_24428,N_24360,N_24046);
xnor U24429 (N_24429,N_23988,N_24245);
or U24430 (N_24430,N_23930,N_23777);
or U24431 (N_24431,N_23985,N_24197);
and U24432 (N_24432,N_23851,N_24113);
xor U24433 (N_24433,N_24195,N_24089);
nor U24434 (N_24434,N_24027,N_24070);
xor U24435 (N_24435,N_24073,N_23976);
nor U24436 (N_24436,N_24233,N_23986);
and U24437 (N_24437,N_23867,N_24120);
nand U24438 (N_24438,N_24077,N_24314);
nor U24439 (N_24439,N_23782,N_24099);
xnor U24440 (N_24440,N_24282,N_24013);
nand U24441 (N_24441,N_23886,N_24280);
or U24442 (N_24442,N_23908,N_23810);
or U24443 (N_24443,N_24294,N_23881);
and U24444 (N_24444,N_24125,N_24078);
nor U24445 (N_24445,N_23990,N_24140);
and U24446 (N_24446,N_24339,N_23878);
nor U24447 (N_24447,N_24038,N_23822);
nand U24448 (N_24448,N_23964,N_23829);
nand U24449 (N_24449,N_24204,N_24055);
and U24450 (N_24450,N_24227,N_24104);
nand U24451 (N_24451,N_24112,N_23925);
nand U24452 (N_24452,N_23963,N_23958);
or U24453 (N_24453,N_24040,N_24087);
nor U24454 (N_24454,N_23953,N_23823);
nand U24455 (N_24455,N_24116,N_23924);
nand U24456 (N_24456,N_24139,N_24048);
nand U24457 (N_24457,N_23855,N_23914);
and U24458 (N_24458,N_24081,N_23879);
or U24459 (N_24459,N_24222,N_24169);
and U24460 (N_24460,N_23767,N_24021);
and U24461 (N_24461,N_24343,N_24163);
nand U24462 (N_24462,N_23871,N_24029);
nand U24463 (N_24463,N_24161,N_24011);
xnor U24464 (N_24464,N_24026,N_23923);
nand U24465 (N_24465,N_24355,N_24138);
or U24466 (N_24466,N_24236,N_23949);
nand U24467 (N_24467,N_24133,N_23935);
xnor U24468 (N_24468,N_23850,N_23761);
nand U24469 (N_24469,N_24368,N_24143);
and U24470 (N_24470,N_23995,N_24150);
xnor U24471 (N_24471,N_24209,N_24024);
nor U24472 (N_24472,N_24336,N_23909);
or U24473 (N_24473,N_23778,N_24083);
or U24474 (N_24474,N_24354,N_24171);
nand U24475 (N_24475,N_24182,N_23877);
xor U24476 (N_24476,N_23784,N_23919);
or U24477 (N_24477,N_24168,N_23845);
xnor U24478 (N_24478,N_23852,N_24030);
and U24479 (N_24479,N_23992,N_24177);
and U24480 (N_24480,N_23857,N_24127);
or U24481 (N_24481,N_24072,N_23898);
nand U24482 (N_24482,N_23794,N_24064);
xor U24483 (N_24483,N_23795,N_24190);
xnor U24484 (N_24484,N_23831,N_23756);
xnor U24485 (N_24485,N_24325,N_24053);
or U24486 (N_24486,N_24123,N_24242);
xnor U24487 (N_24487,N_23906,N_24102);
xnor U24488 (N_24488,N_24307,N_24225);
or U24489 (N_24489,N_23827,N_24337);
xnor U24490 (N_24490,N_24318,N_23796);
or U24491 (N_24491,N_24019,N_24020);
nand U24492 (N_24492,N_24291,N_24352);
xor U24493 (N_24493,N_24295,N_24213);
or U24494 (N_24494,N_24128,N_23844);
or U24495 (N_24495,N_24057,N_24141);
nand U24496 (N_24496,N_24007,N_23896);
nand U24497 (N_24497,N_24338,N_24036);
or U24498 (N_24498,N_24181,N_23956);
or U24499 (N_24499,N_23918,N_24306);
xnor U24500 (N_24500,N_24285,N_24124);
nor U24501 (N_24501,N_24149,N_23917);
or U24502 (N_24502,N_24224,N_24223);
xnor U24503 (N_24503,N_24267,N_24371);
nor U24504 (N_24504,N_24329,N_24252);
nand U24505 (N_24505,N_24148,N_24273);
xnor U24506 (N_24506,N_23974,N_23864);
nor U24507 (N_24507,N_24134,N_24237);
and U24508 (N_24508,N_24132,N_23836);
or U24509 (N_24509,N_24238,N_24012);
and U24510 (N_24510,N_24235,N_23858);
nand U24511 (N_24511,N_24241,N_24226);
or U24512 (N_24512,N_24275,N_24341);
or U24513 (N_24513,N_24323,N_23873);
nand U24514 (N_24514,N_24042,N_24327);
and U24515 (N_24515,N_24370,N_23933);
nor U24516 (N_24516,N_23965,N_24188);
or U24517 (N_24517,N_24239,N_24192);
and U24518 (N_24518,N_23907,N_24175);
xnor U24519 (N_24519,N_24255,N_23989);
nand U24520 (N_24520,N_24248,N_23849);
xnor U24521 (N_24521,N_23947,N_23856);
nand U24522 (N_24522,N_24156,N_24157);
nand U24523 (N_24523,N_23943,N_23981);
nand U24524 (N_24524,N_23800,N_24362);
nand U24525 (N_24525,N_23870,N_24196);
nor U24526 (N_24526,N_23921,N_24054);
and U24527 (N_24527,N_24317,N_23770);
or U24528 (N_24528,N_23833,N_24018);
nand U24529 (N_24529,N_23821,N_24108);
and U24530 (N_24530,N_24032,N_23848);
nor U24531 (N_24531,N_24186,N_23893);
nand U24532 (N_24532,N_23901,N_24279);
nand U24533 (N_24533,N_23785,N_24076);
and U24534 (N_24534,N_24290,N_23753);
xor U24535 (N_24535,N_23838,N_23868);
nor U24536 (N_24536,N_23996,N_23765);
and U24537 (N_24537,N_23837,N_24219);
or U24538 (N_24538,N_23861,N_24050);
nand U24539 (N_24539,N_23847,N_23820);
nand U24540 (N_24540,N_24304,N_23842);
nand U24541 (N_24541,N_24301,N_24211);
and U24542 (N_24542,N_24059,N_24085);
nor U24543 (N_24543,N_23824,N_23752);
or U24544 (N_24544,N_23984,N_23945);
and U24545 (N_24545,N_24271,N_23926);
xor U24546 (N_24546,N_24287,N_23865);
xnor U24547 (N_24547,N_24142,N_24234);
and U24548 (N_24548,N_24174,N_23997);
and U24549 (N_24549,N_24357,N_24066);
xnor U24550 (N_24550,N_23773,N_24300);
nor U24551 (N_24551,N_23903,N_24074);
nand U24552 (N_24552,N_24253,N_24086);
xor U24553 (N_24553,N_23939,N_24151);
and U24554 (N_24554,N_24146,N_24361);
and U24555 (N_24555,N_23980,N_23790);
xnor U24556 (N_24556,N_24372,N_23781);
xor U24557 (N_24557,N_23772,N_23931);
xor U24558 (N_24558,N_23952,N_24183);
and U24559 (N_24559,N_24122,N_23969);
and U24560 (N_24560,N_24356,N_24289);
nor U24561 (N_24561,N_24058,N_24264);
nor U24562 (N_24562,N_24060,N_23920);
nor U24563 (N_24563,N_24299,N_23755);
or U24564 (N_24564,N_24319,N_24269);
nand U24565 (N_24565,N_24115,N_23819);
xor U24566 (N_24566,N_24035,N_23922);
and U24567 (N_24567,N_24257,N_23936);
xnor U24568 (N_24568,N_24367,N_23768);
or U24569 (N_24569,N_24278,N_24292);
nand U24570 (N_24570,N_24109,N_23760);
and U24571 (N_24571,N_24093,N_24272);
or U24572 (N_24572,N_23802,N_23832);
and U24573 (N_24573,N_23854,N_24111);
nor U24574 (N_24574,N_23816,N_23940);
or U24575 (N_24575,N_23763,N_24052);
nand U24576 (N_24576,N_24259,N_23828);
nor U24577 (N_24577,N_23972,N_24193);
nand U24578 (N_24578,N_24201,N_24205);
or U24579 (N_24579,N_24098,N_24265);
or U24580 (N_24580,N_24117,N_24045);
nand U24581 (N_24581,N_24199,N_23804);
xnor U24582 (N_24582,N_24136,N_23806);
and U24583 (N_24583,N_23991,N_24167);
or U24584 (N_24584,N_23937,N_24313);
and U24585 (N_24585,N_24198,N_23966);
nor U24586 (N_24586,N_24080,N_23888);
nand U24587 (N_24587,N_24034,N_24044);
and U24588 (N_24588,N_24075,N_23875);
nor U24589 (N_24589,N_24258,N_23843);
or U24590 (N_24590,N_24173,N_24315);
or U24591 (N_24591,N_24043,N_23902);
or U24592 (N_24592,N_23957,N_24332);
xor U24593 (N_24593,N_24022,N_24004);
nand U24594 (N_24594,N_23780,N_24110);
and U24595 (N_24595,N_23817,N_23754);
and U24596 (N_24596,N_23758,N_23793);
xor U24597 (N_24597,N_23866,N_24286);
or U24598 (N_24598,N_23813,N_24243);
nand U24599 (N_24599,N_24250,N_23934);
or U24600 (N_24600,N_23927,N_24025);
xnor U24601 (N_24601,N_24217,N_24176);
nand U24602 (N_24602,N_23904,N_23880);
or U24603 (N_24603,N_23894,N_23846);
and U24604 (N_24604,N_24288,N_23803);
nor U24605 (N_24605,N_24266,N_23783);
nand U24606 (N_24606,N_24126,N_23978);
nor U24607 (N_24607,N_23809,N_24348);
and U24608 (N_24608,N_24347,N_23841);
nor U24609 (N_24609,N_24082,N_24002);
xnor U24610 (N_24610,N_24061,N_24162);
nand U24611 (N_24611,N_23859,N_23911);
nand U24612 (N_24612,N_23862,N_24107);
or U24613 (N_24613,N_23807,N_23814);
xnor U24614 (N_24614,N_24194,N_24187);
nor U24615 (N_24615,N_24041,N_24284);
or U24616 (N_24616,N_24049,N_23932);
xnor U24617 (N_24617,N_24353,N_23960);
nand U24618 (N_24618,N_24017,N_23839);
nor U24619 (N_24619,N_24106,N_24096);
nor U24620 (N_24620,N_23959,N_23929);
nand U24621 (N_24621,N_24210,N_24240);
or U24622 (N_24622,N_24218,N_24185);
or U24623 (N_24623,N_23891,N_23792);
nand U24624 (N_24624,N_23789,N_23977);
nor U24625 (N_24625,N_23890,N_23801);
xnor U24626 (N_24626,N_23774,N_24310);
xnor U24627 (N_24627,N_24260,N_24166);
or U24628 (N_24628,N_24221,N_24009);
and U24629 (N_24629,N_24206,N_24349);
xor U24630 (N_24630,N_24137,N_24131);
nor U24631 (N_24631,N_23884,N_23994);
nor U24632 (N_24632,N_24328,N_24228);
or U24633 (N_24633,N_24000,N_24364);
or U24634 (N_24634,N_23751,N_23889);
nand U24635 (N_24635,N_24088,N_23840);
and U24636 (N_24636,N_23883,N_24351);
nand U24637 (N_24637,N_23951,N_24230);
and U24638 (N_24638,N_23950,N_23805);
nand U24639 (N_24639,N_24358,N_24365);
and U24640 (N_24640,N_24119,N_24262);
nand U24641 (N_24641,N_24256,N_23987);
nor U24642 (N_24642,N_24071,N_24308);
nor U24643 (N_24643,N_23759,N_24261);
nor U24644 (N_24644,N_24094,N_24180);
nand U24645 (N_24645,N_23887,N_24200);
nand U24646 (N_24646,N_24158,N_23961);
and U24647 (N_24647,N_23892,N_24277);
or U24648 (N_24648,N_24178,N_24298);
or U24649 (N_24649,N_23769,N_23975);
nand U24650 (N_24650,N_24103,N_23812);
xor U24651 (N_24651,N_24203,N_23912);
xor U24652 (N_24652,N_24147,N_24189);
nand U24653 (N_24653,N_23853,N_24165);
xnor U24654 (N_24654,N_24214,N_24220);
nand U24655 (N_24655,N_23797,N_24145);
nand U24656 (N_24656,N_23775,N_24010);
or U24657 (N_24657,N_24095,N_23776);
nand U24658 (N_24658,N_24246,N_24090);
or U24659 (N_24659,N_24069,N_23869);
nor U24660 (N_24660,N_24135,N_23882);
and U24661 (N_24661,N_23885,N_24207);
and U24662 (N_24662,N_23771,N_24179);
or U24663 (N_24663,N_24316,N_23938);
nor U24664 (N_24664,N_23826,N_24023);
and U24665 (N_24665,N_24014,N_23808);
nor U24666 (N_24666,N_24092,N_23993);
nor U24667 (N_24667,N_23766,N_23825);
xor U24668 (N_24668,N_24028,N_24056);
nor U24669 (N_24669,N_24321,N_24015);
nor U24670 (N_24670,N_23983,N_23999);
nand U24671 (N_24671,N_23815,N_24184);
xnor U24672 (N_24672,N_24309,N_24159);
and U24673 (N_24673,N_23928,N_24311);
xor U24674 (N_24674,N_24335,N_24276);
or U24675 (N_24675,N_23897,N_24105);
nand U24676 (N_24676,N_24373,N_24342);
nand U24677 (N_24677,N_24340,N_24283);
and U24678 (N_24678,N_24153,N_23895);
nand U24679 (N_24679,N_24001,N_23905);
and U24680 (N_24680,N_24118,N_24251);
nor U24681 (N_24681,N_24232,N_24231);
and U24682 (N_24682,N_24154,N_23762);
xnor U24683 (N_24683,N_24065,N_23955);
and U24684 (N_24684,N_23764,N_24215);
nor U24685 (N_24685,N_24152,N_24297);
nand U24686 (N_24686,N_23970,N_23944);
nor U24687 (N_24687,N_24039,N_23958);
nor U24688 (N_24688,N_24336,N_24368);
nand U24689 (N_24689,N_23771,N_24048);
nor U24690 (N_24690,N_24021,N_24207);
nand U24691 (N_24691,N_23953,N_24066);
xor U24692 (N_24692,N_24109,N_23830);
and U24693 (N_24693,N_24193,N_23922);
and U24694 (N_24694,N_23827,N_23757);
nor U24695 (N_24695,N_24002,N_24313);
nand U24696 (N_24696,N_24077,N_24245);
or U24697 (N_24697,N_24174,N_24269);
nand U24698 (N_24698,N_24354,N_24051);
nand U24699 (N_24699,N_24045,N_23769);
nand U24700 (N_24700,N_24256,N_24153);
nand U24701 (N_24701,N_23901,N_24365);
and U24702 (N_24702,N_24008,N_24098);
and U24703 (N_24703,N_23845,N_23926);
nand U24704 (N_24704,N_23875,N_24191);
nand U24705 (N_24705,N_24113,N_23754);
xor U24706 (N_24706,N_24192,N_24164);
nand U24707 (N_24707,N_24154,N_24160);
nand U24708 (N_24708,N_24099,N_23911);
nand U24709 (N_24709,N_23756,N_23762);
and U24710 (N_24710,N_23991,N_24312);
nand U24711 (N_24711,N_24300,N_23771);
nor U24712 (N_24712,N_24002,N_23880);
nand U24713 (N_24713,N_23795,N_24157);
and U24714 (N_24714,N_23951,N_23797);
xor U24715 (N_24715,N_24121,N_24352);
nor U24716 (N_24716,N_24011,N_23778);
or U24717 (N_24717,N_23911,N_23993);
nand U24718 (N_24718,N_23776,N_23940);
nand U24719 (N_24719,N_24355,N_24198);
nor U24720 (N_24720,N_24338,N_23867);
or U24721 (N_24721,N_24329,N_24268);
and U24722 (N_24722,N_24027,N_24010);
nor U24723 (N_24723,N_24160,N_24291);
and U24724 (N_24724,N_23921,N_24107);
nor U24725 (N_24725,N_23960,N_24367);
nor U24726 (N_24726,N_24252,N_23876);
xor U24727 (N_24727,N_24128,N_23904);
or U24728 (N_24728,N_24085,N_23832);
xnor U24729 (N_24729,N_23916,N_23795);
xor U24730 (N_24730,N_24036,N_23900);
nand U24731 (N_24731,N_24159,N_24200);
xor U24732 (N_24732,N_24144,N_24343);
nor U24733 (N_24733,N_24347,N_24052);
nor U24734 (N_24734,N_23978,N_23941);
nor U24735 (N_24735,N_24080,N_24038);
xnor U24736 (N_24736,N_23852,N_23967);
or U24737 (N_24737,N_23805,N_23793);
nand U24738 (N_24738,N_24259,N_24305);
and U24739 (N_24739,N_24065,N_24359);
xor U24740 (N_24740,N_24002,N_24076);
xor U24741 (N_24741,N_24151,N_23773);
nor U24742 (N_24742,N_24309,N_23989);
xnor U24743 (N_24743,N_23993,N_23868);
or U24744 (N_24744,N_23917,N_23779);
and U24745 (N_24745,N_24140,N_24219);
nor U24746 (N_24746,N_23910,N_24247);
nor U24747 (N_24747,N_23795,N_24195);
xor U24748 (N_24748,N_23820,N_24049);
nand U24749 (N_24749,N_23813,N_24115);
or U24750 (N_24750,N_23986,N_24184);
nor U24751 (N_24751,N_24272,N_23772);
nand U24752 (N_24752,N_24147,N_24002);
nor U24753 (N_24753,N_24210,N_24047);
and U24754 (N_24754,N_23831,N_24122);
nand U24755 (N_24755,N_23894,N_24284);
and U24756 (N_24756,N_23954,N_23847);
nor U24757 (N_24757,N_24199,N_24281);
xor U24758 (N_24758,N_23835,N_23854);
and U24759 (N_24759,N_24160,N_24287);
nand U24760 (N_24760,N_24153,N_24004);
nand U24761 (N_24761,N_24274,N_24146);
or U24762 (N_24762,N_23974,N_23982);
and U24763 (N_24763,N_23888,N_24254);
nor U24764 (N_24764,N_23796,N_24184);
or U24765 (N_24765,N_23837,N_24237);
xor U24766 (N_24766,N_24011,N_23768);
nand U24767 (N_24767,N_23821,N_24195);
and U24768 (N_24768,N_23768,N_24083);
xnor U24769 (N_24769,N_24261,N_23958);
nor U24770 (N_24770,N_23826,N_24044);
nand U24771 (N_24771,N_23823,N_24001);
nand U24772 (N_24772,N_23996,N_24049);
nand U24773 (N_24773,N_23926,N_23914);
nand U24774 (N_24774,N_24009,N_23847);
and U24775 (N_24775,N_24300,N_24336);
and U24776 (N_24776,N_24268,N_23819);
xnor U24777 (N_24777,N_23875,N_24241);
or U24778 (N_24778,N_24218,N_23794);
nand U24779 (N_24779,N_23856,N_24016);
and U24780 (N_24780,N_24292,N_23806);
nand U24781 (N_24781,N_23813,N_23759);
xnor U24782 (N_24782,N_24329,N_23822);
nor U24783 (N_24783,N_24322,N_24095);
and U24784 (N_24784,N_24347,N_23801);
or U24785 (N_24785,N_24090,N_24272);
xor U24786 (N_24786,N_24296,N_24354);
or U24787 (N_24787,N_24010,N_24270);
and U24788 (N_24788,N_24255,N_24223);
or U24789 (N_24789,N_23989,N_23787);
xnor U24790 (N_24790,N_24138,N_24308);
nand U24791 (N_24791,N_23851,N_23758);
or U24792 (N_24792,N_24172,N_23773);
nand U24793 (N_24793,N_24202,N_24307);
or U24794 (N_24794,N_24250,N_23909);
nor U24795 (N_24795,N_24301,N_24336);
nand U24796 (N_24796,N_24158,N_23844);
xnor U24797 (N_24797,N_23794,N_23919);
nand U24798 (N_24798,N_24138,N_24258);
or U24799 (N_24799,N_24049,N_23792);
nand U24800 (N_24800,N_24027,N_23984);
xor U24801 (N_24801,N_23908,N_24252);
xnor U24802 (N_24802,N_23896,N_24141);
or U24803 (N_24803,N_24358,N_24333);
and U24804 (N_24804,N_24249,N_24303);
xor U24805 (N_24805,N_24072,N_23910);
xor U24806 (N_24806,N_24098,N_24365);
and U24807 (N_24807,N_24102,N_24229);
nor U24808 (N_24808,N_24167,N_23882);
nor U24809 (N_24809,N_24126,N_23778);
or U24810 (N_24810,N_23963,N_24325);
nor U24811 (N_24811,N_24017,N_24190);
nor U24812 (N_24812,N_24351,N_24247);
nand U24813 (N_24813,N_23878,N_23921);
nor U24814 (N_24814,N_24374,N_24294);
or U24815 (N_24815,N_24285,N_23924);
xor U24816 (N_24816,N_24097,N_24208);
and U24817 (N_24817,N_24037,N_23783);
nor U24818 (N_24818,N_23773,N_23874);
nor U24819 (N_24819,N_24148,N_24088);
nor U24820 (N_24820,N_23853,N_23880);
nand U24821 (N_24821,N_24223,N_23937);
xor U24822 (N_24822,N_23756,N_24144);
xnor U24823 (N_24823,N_23892,N_23947);
xor U24824 (N_24824,N_24079,N_24072);
nor U24825 (N_24825,N_23958,N_23918);
xnor U24826 (N_24826,N_24105,N_23807);
and U24827 (N_24827,N_23924,N_23912);
or U24828 (N_24828,N_24174,N_23899);
or U24829 (N_24829,N_24091,N_23874);
xor U24830 (N_24830,N_24146,N_23799);
or U24831 (N_24831,N_24351,N_23825);
or U24832 (N_24832,N_24104,N_24214);
nand U24833 (N_24833,N_23880,N_24254);
and U24834 (N_24834,N_24277,N_24160);
or U24835 (N_24835,N_24326,N_23849);
nand U24836 (N_24836,N_23840,N_23945);
nand U24837 (N_24837,N_24314,N_24080);
and U24838 (N_24838,N_23927,N_24269);
or U24839 (N_24839,N_23857,N_23812);
or U24840 (N_24840,N_24103,N_23782);
xnor U24841 (N_24841,N_24045,N_24157);
xnor U24842 (N_24842,N_24159,N_23973);
nor U24843 (N_24843,N_24136,N_24065);
nor U24844 (N_24844,N_24347,N_23985);
xnor U24845 (N_24845,N_23876,N_23896);
nor U24846 (N_24846,N_23809,N_24198);
nand U24847 (N_24847,N_24350,N_24256);
or U24848 (N_24848,N_24236,N_24030);
nor U24849 (N_24849,N_24098,N_23782);
xor U24850 (N_24850,N_24303,N_24205);
nand U24851 (N_24851,N_23839,N_24106);
nand U24852 (N_24852,N_24158,N_23875);
or U24853 (N_24853,N_23771,N_23866);
nand U24854 (N_24854,N_23845,N_24142);
nand U24855 (N_24855,N_24055,N_23775);
nor U24856 (N_24856,N_23888,N_24033);
nor U24857 (N_24857,N_24358,N_24364);
or U24858 (N_24858,N_24352,N_23828);
and U24859 (N_24859,N_24266,N_23885);
or U24860 (N_24860,N_23905,N_24118);
or U24861 (N_24861,N_24021,N_24255);
nor U24862 (N_24862,N_24254,N_24060);
nor U24863 (N_24863,N_23811,N_23781);
xnor U24864 (N_24864,N_23800,N_23947);
or U24865 (N_24865,N_23751,N_24172);
nand U24866 (N_24866,N_23814,N_24286);
and U24867 (N_24867,N_24276,N_23780);
xor U24868 (N_24868,N_24097,N_23824);
nand U24869 (N_24869,N_24248,N_24034);
xor U24870 (N_24870,N_24228,N_24311);
nand U24871 (N_24871,N_23985,N_24300);
xnor U24872 (N_24872,N_24176,N_24202);
or U24873 (N_24873,N_24275,N_23868);
nand U24874 (N_24874,N_24037,N_23971);
nand U24875 (N_24875,N_24087,N_23894);
nor U24876 (N_24876,N_23991,N_24107);
nand U24877 (N_24877,N_24109,N_24258);
or U24878 (N_24878,N_24357,N_23978);
nand U24879 (N_24879,N_23869,N_23970);
nand U24880 (N_24880,N_23885,N_23926);
nand U24881 (N_24881,N_24231,N_24307);
xnor U24882 (N_24882,N_23805,N_24163);
or U24883 (N_24883,N_23757,N_24307);
nor U24884 (N_24884,N_23864,N_24262);
nor U24885 (N_24885,N_23933,N_24041);
nand U24886 (N_24886,N_24217,N_24061);
nand U24887 (N_24887,N_23904,N_23944);
nor U24888 (N_24888,N_23753,N_24099);
or U24889 (N_24889,N_24370,N_23954);
xor U24890 (N_24890,N_24346,N_24098);
or U24891 (N_24891,N_24124,N_24036);
xnor U24892 (N_24892,N_24058,N_24073);
xor U24893 (N_24893,N_23766,N_24234);
or U24894 (N_24894,N_24081,N_24320);
or U24895 (N_24895,N_24241,N_24248);
xnor U24896 (N_24896,N_24310,N_24190);
nand U24897 (N_24897,N_24012,N_23853);
nor U24898 (N_24898,N_24031,N_23833);
nand U24899 (N_24899,N_24108,N_23867);
or U24900 (N_24900,N_24337,N_23915);
nand U24901 (N_24901,N_23902,N_23811);
and U24902 (N_24902,N_24111,N_23810);
and U24903 (N_24903,N_23782,N_24198);
nor U24904 (N_24904,N_24336,N_24260);
and U24905 (N_24905,N_23864,N_23752);
nor U24906 (N_24906,N_23837,N_23968);
xnor U24907 (N_24907,N_24274,N_23860);
xor U24908 (N_24908,N_24275,N_23888);
xnor U24909 (N_24909,N_24107,N_24091);
or U24910 (N_24910,N_24105,N_24075);
nand U24911 (N_24911,N_24137,N_24052);
nand U24912 (N_24912,N_24355,N_24109);
or U24913 (N_24913,N_24196,N_24000);
nand U24914 (N_24914,N_24043,N_24010);
nor U24915 (N_24915,N_24222,N_23862);
or U24916 (N_24916,N_23837,N_24010);
or U24917 (N_24917,N_24039,N_24353);
nor U24918 (N_24918,N_23914,N_23851);
nor U24919 (N_24919,N_24231,N_23933);
or U24920 (N_24920,N_24177,N_24360);
nand U24921 (N_24921,N_23919,N_24253);
nor U24922 (N_24922,N_24313,N_23809);
xnor U24923 (N_24923,N_24335,N_24146);
nand U24924 (N_24924,N_23810,N_23942);
or U24925 (N_24925,N_24083,N_24371);
xor U24926 (N_24926,N_23757,N_23756);
and U24927 (N_24927,N_24237,N_24341);
or U24928 (N_24928,N_24323,N_24194);
or U24929 (N_24929,N_24320,N_23829);
nor U24930 (N_24930,N_24281,N_23880);
and U24931 (N_24931,N_24116,N_24217);
or U24932 (N_24932,N_24246,N_24127);
xor U24933 (N_24933,N_24005,N_24050);
nor U24934 (N_24934,N_24097,N_24049);
nand U24935 (N_24935,N_23960,N_23901);
or U24936 (N_24936,N_23901,N_24204);
xnor U24937 (N_24937,N_24107,N_23847);
nand U24938 (N_24938,N_24211,N_23858);
and U24939 (N_24939,N_23941,N_24216);
nor U24940 (N_24940,N_23879,N_23988);
xor U24941 (N_24941,N_24282,N_23971);
or U24942 (N_24942,N_24054,N_23787);
and U24943 (N_24943,N_24182,N_23832);
xnor U24944 (N_24944,N_23944,N_24283);
nand U24945 (N_24945,N_24053,N_23918);
xnor U24946 (N_24946,N_24070,N_24048);
nor U24947 (N_24947,N_23769,N_24282);
xor U24948 (N_24948,N_24051,N_23991);
xnor U24949 (N_24949,N_24290,N_24365);
xor U24950 (N_24950,N_23816,N_24188);
or U24951 (N_24951,N_24303,N_24301);
nand U24952 (N_24952,N_24083,N_24129);
or U24953 (N_24953,N_23946,N_24165);
and U24954 (N_24954,N_23843,N_23879);
nand U24955 (N_24955,N_23844,N_24109);
xnor U24956 (N_24956,N_24028,N_24360);
and U24957 (N_24957,N_23891,N_24309);
xor U24958 (N_24958,N_23797,N_23956);
xor U24959 (N_24959,N_24194,N_24033);
or U24960 (N_24960,N_24167,N_24207);
nand U24961 (N_24961,N_24107,N_24098);
or U24962 (N_24962,N_23850,N_24164);
nand U24963 (N_24963,N_24171,N_24319);
and U24964 (N_24964,N_23860,N_23983);
or U24965 (N_24965,N_24061,N_24150);
nor U24966 (N_24966,N_23969,N_24268);
xnor U24967 (N_24967,N_24288,N_23824);
and U24968 (N_24968,N_24181,N_23820);
and U24969 (N_24969,N_24283,N_24127);
xor U24970 (N_24970,N_24166,N_24266);
nor U24971 (N_24971,N_24341,N_23849);
and U24972 (N_24972,N_24016,N_23806);
nand U24973 (N_24973,N_23977,N_24066);
or U24974 (N_24974,N_24295,N_24081);
xor U24975 (N_24975,N_24181,N_24231);
and U24976 (N_24976,N_24334,N_23890);
or U24977 (N_24977,N_24272,N_24125);
or U24978 (N_24978,N_23877,N_23980);
nand U24979 (N_24979,N_24189,N_23832);
nand U24980 (N_24980,N_23750,N_23978);
and U24981 (N_24981,N_23947,N_23790);
nand U24982 (N_24982,N_24115,N_23803);
xor U24983 (N_24983,N_24038,N_23826);
nor U24984 (N_24984,N_24320,N_23920);
nor U24985 (N_24985,N_24259,N_24014);
nor U24986 (N_24986,N_23967,N_24271);
or U24987 (N_24987,N_23754,N_24086);
and U24988 (N_24988,N_24086,N_23825);
nor U24989 (N_24989,N_23865,N_23825);
and U24990 (N_24990,N_24172,N_24003);
nor U24991 (N_24991,N_24035,N_24206);
nor U24992 (N_24992,N_24075,N_23789);
xnor U24993 (N_24993,N_23977,N_24059);
nand U24994 (N_24994,N_24003,N_24264);
xnor U24995 (N_24995,N_23785,N_24057);
or U24996 (N_24996,N_24247,N_24265);
or U24997 (N_24997,N_24292,N_24087);
and U24998 (N_24998,N_24181,N_24038);
and U24999 (N_24999,N_23808,N_24125);
or UO_0 (O_0,N_24608,N_24768);
and UO_1 (O_1,N_24431,N_24538);
nor UO_2 (O_2,N_24998,N_24535);
nor UO_3 (O_3,N_24919,N_24774);
xnor UO_4 (O_4,N_24408,N_24733);
xnor UO_5 (O_5,N_24427,N_24771);
xor UO_6 (O_6,N_24812,N_24454);
xor UO_7 (O_7,N_24776,N_24884);
nor UO_8 (O_8,N_24855,N_24601);
and UO_9 (O_9,N_24599,N_24539);
and UO_10 (O_10,N_24435,N_24870);
nand UO_11 (O_11,N_24527,N_24739);
nor UO_12 (O_12,N_24740,N_24916);
and UO_13 (O_13,N_24637,N_24517);
xnor UO_14 (O_14,N_24809,N_24693);
nand UO_15 (O_15,N_24876,N_24860);
nor UO_16 (O_16,N_24939,N_24629);
nand UO_17 (O_17,N_24568,N_24623);
and UO_18 (O_18,N_24666,N_24488);
nor UO_19 (O_19,N_24644,N_24668);
or UO_20 (O_20,N_24796,N_24694);
nor UO_21 (O_21,N_24839,N_24607);
nand UO_22 (O_22,N_24639,N_24907);
nand UO_23 (O_23,N_24953,N_24407);
and UO_24 (O_24,N_24600,N_24927);
nand UO_25 (O_25,N_24756,N_24626);
and UO_26 (O_26,N_24443,N_24890);
or UO_27 (O_27,N_24708,N_24522);
xnor UO_28 (O_28,N_24550,N_24924);
nor UO_29 (O_29,N_24388,N_24524);
xnor UO_30 (O_30,N_24753,N_24959);
and UO_31 (O_31,N_24417,N_24560);
xnor UO_32 (O_32,N_24494,N_24949);
xor UO_33 (O_33,N_24780,N_24791);
and UO_34 (O_34,N_24983,N_24605);
or UO_35 (O_35,N_24988,N_24707);
xnor UO_36 (O_36,N_24514,N_24409);
xor UO_37 (O_37,N_24686,N_24680);
nor UO_38 (O_38,N_24687,N_24399);
nand UO_39 (O_39,N_24596,N_24912);
nand UO_40 (O_40,N_24705,N_24458);
nand UO_41 (O_41,N_24935,N_24641);
xnor UO_42 (O_42,N_24845,N_24567);
and UO_43 (O_43,N_24647,N_24667);
nand UO_44 (O_44,N_24571,N_24944);
nor UO_45 (O_45,N_24795,N_24579);
xor UO_46 (O_46,N_24381,N_24671);
or UO_47 (O_47,N_24814,N_24398);
and UO_48 (O_48,N_24759,N_24730);
xnor UO_49 (O_49,N_24999,N_24893);
xor UO_50 (O_50,N_24700,N_24569);
and UO_51 (O_51,N_24670,N_24741);
and UO_52 (O_52,N_24932,N_24900);
and UO_53 (O_53,N_24824,N_24528);
nand UO_54 (O_54,N_24909,N_24719);
nor UO_55 (O_55,N_24718,N_24658);
nand UO_56 (O_56,N_24899,N_24383);
or UO_57 (O_57,N_24689,N_24546);
nor UO_58 (O_58,N_24624,N_24785);
xnor UO_59 (O_59,N_24688,N_24864);
nand UO_60 (O_60,N_24745,N_24572);
xor UO_61 (O_61,N_24473,N_24833);
nor UO_62 (O_62,N_24763,N_24564);
and UO_63 (O_63,N_24386,N_24464);
or UO_64 (O_64,N_24697,N_24404);
nor UO_65 (O_65,N_24575,N_24425);
xor UO_66 (O_66,N_24918,N_24760);
or UO_67 (O_67,N_24434,N_24789);
or UO_68 (O_68,N_24834,N_24875);
or UO_69 (O_69,N_24419,N_24881);
or UO_70 (O_70,N_24439,N_24946);
or UO_71 (O_71,N_24751,N_24610);
nor UO_72 (O_72,N_24818,N_24500);
or UO_73 (O_73,N_24905,N_24917);
nand UO_74 (O_74,N_24798,N_24611);
and UO_75 (O_75,N_24931,N_24561);
nand UO_76 (O_76,N_24423,N_24736);
nor UO_77 (O_77,N_24782,N_24574);
or UO_78 (O_78,N_24920,N_24835);
nand UO_79 (O_79,N_24861,N_24856);
xnor UO_80 (O_80,N_24971,N_24851);
and UO_81 (O_81,N_24429,N_24643);
or UO_82 (O_82,N_24551,N_24906);
nor UO_83 (O_83,N_24865,N_24677);
and UO_84 (O_84,N_24991,N_24886);
nand UO_85 (O_85,N_24980,N_24582);
xor UO_86 (O_86,N_24915,N_24992);
nor UO_87 (O_87,N_24754,N_24889);
or UO_88 (O_88,N_24468,N_24709);
xnor UO_89 (O_89,N_24485,N_24544);
and UO_90 (O_90,N_24808,N_24866);
nor UO_91 (O_91,N_24591,N_24595);
or UO_92 (O_92,N_24786,N_24747);
xor UO_93 (O_93,N_24987,N_24533);
and UO_94 (O_94,N_24593,N_24725);
and UO_95 (O_95,N_24836,N_24961);
nand UO_96 (O_96,N_24430,N_24462);
or UO_97 (O_97,N_24478,N_24586);
nand UO_98 (O_98,N_24547,N_24380);
xor UO_99 (O_99,N_24476,N_24631);
nor UO_100 (O_100,N_24698,N_24857);
or UO_101 (O_101,N_24681,N_24994);
or UO_102 (O_102,N_24772,N_24603);
or UO_103 (O_103,N_24606,N_24672);
xnor UO_104 (O_104,N_24728,N_24928);
and UO_105 (O_105,N_24902,N_24489);
xor UO_106 (O_106,N_24966,N_24649);
nor UO_107 (O_107,N_24438,N_24437);
or UO_108 (O_108,N_24685,N_24797);
nor UO_109 (O_109,N_24422,N_24512);
and UO_110 (O_110,N_24613,N_24981);
or UO_111 (O_111,N_24416,N_24376);
or UO_112 (O_112,N_24618,N_24804);
or UO_113 (O_113,N_24852,N_24752);
nor UO_114 (O_114,N_24682,N_24679);
xnor UO_115 (O_115,N_24993,N_24664);
and UO_116 (O_116,N_24841,N_24432);
nor UO_117 (O_117,N_24989,N_24807);
nor UO_118 (O_118,N_24502,N_24816);
nand UO_119 (O_119,N_24395,N_24982);
nand UO_120 (O_120,N_24499,N_24482);
nand UO_121 (O_121,N_24913,N_24453);
and UO_122 (O_122,N_24669,N_24825);
and UO_123 (O_123,N_24765,N_24545);
nor UO_124 (O_124,N_24878,N_24487);
nor UO_125 (O_125,N_24810,N_24457);
and UO_126 (O_126,N_24727,N_24492);
and UO_127 (O_127,N_24676,N_24471);
or UO_128 (O_128,N_24506,N_24630);
nand UO_129 (O_129,N_24832,N_24628);
nor UO_130 (O_130,N_24445,N_24387);
nor UO_131 (O_131,N_24632,N_24871);
or UO_132 (O_132,N_24862,N_24684);
xnor UO_133 (O_133,N_24849,N_24642);
and UO_134 (O_134,N_24475,N_24617);
nand UO_135 (O_135,N_24412,N_24384);
and UO_136 (O_136,N_24735,N_24691);
nand UO_137 (O_137,N_24926,N_24444);
and UO_138 (O_138,N_24844,N_24954);
and UO_139 (O_139,N_24778,N_24910);
xor UO_140 (O_140,N_24513,N_24703);
nand UO_141 (O_141,N_24405,N_24717);
and UO_142 (O_142,N_24699,N_24925);
xor UO_143 (O_143,N_24769,N_24732);
or UO_144 (O_144,N_24651,N_24377);
and UO_145 (O_145,N_24625,N_24616);
nand UO_146 (O_146,N_24466,N_24540);
and UO_147 (O_147,N_24830,N_24526);
and UO_148 (O_148,N_24938,N_24635);
and UO_149 (O_149,N_24465,N_24848);
and UO_150 (O_150,N_24652,N_24720);
and UO_151 (O_151,N_24716,N_24903);
nand UO_152 (O_152,N_24390,N_24933);
and UO_153 (O_153,N_24562,N_24577);
nand UO_154 (O_154,N_24737,N_24887);
or UO_155 (O_155,N_24621,N_24414);
or UO_156 (O_156,N_24588,N_24823);
xnor UO_157 (O_157,N_24790,N_24821);
and UO_158 (O_158,N_24721,N_24976);
nand UO_159 (O_159,N_24799,N_24755);
nor UO_160 (O_160,N_24880,N_24477);
xnor UO_161 (O_161,N_24518,N_24654);
or UO_162 (O_162,N_24587,N_24843);
nor UO_163 (O_163,N_24622,N_24516);
nand UO_164 (O_164,N_24748,N_24868);
nor UO_165 (O_165,N_24952,N_24418);
and UO_166 (O_166,N_24556,N_24660);
nand UO_167 (O_167,N_24634,N_24638);
xnor UO_168 (O_168,N_24777,N_24655);
nor UO_169 (O_169,N_24491,N_24396);
and UO_170 (O_170,N_24853,N_24389);
and UO_171 (O_171,N_24715,N_24873);
or UO_172 (O_172,N_24746,N_24558);
or UO_173 (O_173,N_24895,N_24766);
nor UO_174 (O_174,N_24744,N_24822);
xnor UO_175 (O_175,N_24509,N_24842);
nand UO_176 (O_176,N_24743,N_24484);
nand UO_177 (O_177,N_24662,N_24984);
xor UO_178 (O_178,N_24397,N_24609);
nor UO_179 (O_179,N_24483,N_24995);
xor UO_180 (O_180,N_24585,N_24554);
and UO_181 (O_181,N_24452,N_24879);
and UO_182 (O_182,N_24511,N_24440);
nand UO_183 (O_183,N_24702,N_24410);
nand UO_184 (O_184,N_24896,N_24403);
xor UO_185 (O_185,N_24520,N_24963);
nand UO_186 (O_186,N_24767,N_24723);
xor UO_187 (O_187,N_24433,N_24594);
and UO_188 (O_188,N_24461,N_24970);
and UO_189 (O_189,N_24507,N_24415);
or UO_190 (O_190,N_24529,N_24901);
nor UO_191 (O_191,N_24646,N_24555);
or UO_192 (O_192,N_24838,N_24820);
and UO_193 (O_193,N_24456,N_24469);
nor UO_194 (O_194,N_24542,N_24784);
xor UO_195 (O_195,N_24548,N_24451);
and UO_196 (O_196,N_24578,N_24867);
nor UO_197 (O_197,N_24503,N_24956);
xor UO_198 (O_198,N_24964,N_24570);
nand UO_199 (O_199,N_24770,N_24583);
xnor UO_200 (O_200,N_24428,N_24749);
or UO_201 (O_201,N_24937,N_24650);
nand UO_202 (O_202,N_24663,N_24627);
or UO_203 (O_203,N_24525,N_24576);
xnor UO_204 (O_204,N_24815,N_24612);
nand UO_205 (O_205,N_24584,N_24891);
or UO_206 (O_206,N_24773,N_24460);
nor UO_207 (O_207,N_24519,N_24534);
or UO_208 (O_208,N_24420,N_24758);
or UO_209 (O_209,N_24731,N_24455);
nand UO_210 (O_210,N_24921,N_24750);
or UO_211 (O_211,N_24496,N_24536);
xor UO_212 (O_212,N_24659,N_24883);
xnor UO_213 (O_213,N_24792,N_24467);
xor UO_214 (O_214,N_24950,N_24581);
or UO_215 (O_215,N_24775,N_24967);
and UO_216 (O_216,N_24490,N_24532);
or UO_217 (O_217,N_24801,N_24614);
or UO_218 (O_218,N_24972,N_24724);
or UO_219 (O_219,N_24831,N_24978);
or UO_220 (O_220,N_24897,N_24375);
nor UO_221 (O_221,N_24706,N_24783);
nand UO_222 (O_222,N_24923,N_24996);
xor UO_223 (O_223,N_24645,N_24779);
nor UO_224 (O_224,N_24947,N_24580);
xor UO_225 (O_225,N_24761,N_24592);
or UO_226 (O_226,N_24553,N_24828);
and UO_227 (O_227,N_24498,N_24882);
and UO_228 (O_228,N_24840,N_24442);
nand UO_229 (O_229,N_24975,N_24531);
nand UO_230 (O_230,N_24888,N_24690);
xor UO_231 (O_231,N_24382,N_24762);
and UO_232 (O_232,N_24379,N_24712);
nand UO_233 (O_233,N_24653,N_24448);
nor UO_234 (O_234,N_24885,N_24436);
or UO_235 (O_235,N_24413,N_24850);
nor UO_236 (O_236,N_24738,N_24965);
xnor UO_237 (O_237,N_24973,N_24378);
nor UO_238 (O_238,N_24406,N_24559);
nor UO_239 (O_239,N_24922,N_24537);
nand UO_240 (O_240,N_24819,N_24869);
nand UO_241 (O_241,N_24803,N_24657);
and UO_242 (O_242,N_24962,N_24446);
xor UO_243 (O_243,N_24904,N_24764);
nand UO_244 (O_244,N_24898,N_24892);
and UO_245 (O_245,N_24541,N_24805);
xor UO_246 (O_246,N_24549,N_24480);
nand UO_247 (O_247,N_24479,N_24497);
nor UO_248 (O_248,N_24450,N_24391);
or UO_249 (O_249,N_24800,N_24459);
nor UO_250 (O_250,N_24692,N_24573);
nand UO_251 (O_251,N_24486,N_24557);
nand UO_252 (O_252,N_24426,N_24504);
or UO_253 (O_253,N_24590,N_24675);
nor UO_254 (O_254,N_24523,N_24633);
nor UO_255 (O_255,N_24788,N_24794);
or UO_256 (O_256,N_24859,N_24392);
xnor UO_257 (O_257,N_24701,N_24463);
xor UO_258 (O_258,N_24874,N_24957);
nand UO_259 (O_259,N_24530,N_24521);
or UO_260 (O_260,N_24941,N_24793);
and UO_261 (O_261,N_24615,N_24449);
nand UO_262 (O_262,N_24472,N_24934);
nand UO_263 (O_263,N_24495,N_24936);
xnor UO_264 (O_264,N_24846,N_24908);
or UO_265 (O_265,N_24665,N_24474);
xor UO_266 (O_266,N_24447,N_24411);
or UO_267 (O_267,N_24863,N_24402);
nand UO_268 (O_268,N_24813,N_24604);
and UO_269 (O_269,N_24911,N_24722);
nand UO_270 (O_270,N_24385,N_24974);
or UO_271 (O_271,N_24620,N_24400);
nor UO_272 (O_272,N_24894,N_24713);
xnor UO_273 (O_273,N_24734,N_24552);
xor UO_274 (O_274,N_24837,N_24501);
and UO_275 (O_275,N_24781,N_24726);
and UO_276 (O_276,N_24589,N_24948);
or UO_277 (O_277,N_24640,N_24619);
and UO_278 (O_278,N_24424,N_24854);
xor UO_279 (O_279,N_24729,N_24817);
nor UO_280 (O_280,N_24811,N_24802);
or UO_281 (O_281,N_24543,N_24393);
xnor UO_282 (O_282,N_24979,N_24441);
nor UO_283 (O_283,N_24757,N_24711);
nand UO_284 (O_284,N_24597,N_24481);
nand UO_285 (O_285,N_24714,N_24636);
nand UO_286 (O_286,N_24598,N_24710);
xnor UO_287 (O_287,N_24508,N_24858);
xor UO_288 (O_288,N_24565,N_24942);
xor UO_289 (O_289,N_24997,N_24470);
or UO_290 (O_290,N_24704,N_24683);
nor UO_291 (O_291,N_24977,N_24958);
nor UO_292 (O_292,N_24505,N_24566);
nor UO_293 (O_293,N_24696,N_24787);
nand UO_294 (O_294,N_24656,N_24826);
nor UO_295 (O_295,N_24661,N_24968);
nand UO_296 (O_296,N_24929,N_24401);
or UO_297 (O_297,N_24674,N_24945);
nor UO_298 (O_298,N_24493,N_24648);
nor UO_299 (O_299,N_24510,N_24986);
nor UO_300 (O_300,N_24515,N_24742);
xor UO_301 (O_301,N_24872,N_24602);
nor UO_302 (O_302,N_24394,N_24421);
xnor UO_303 (O_303,N_24829,N_24673);
xnor UO_304 (O_304,N_24695,N_24678);
or UO_305 (O_305,N_24960,N_24969);
nand UO_306 (O_306,N_24990,N_24985);
nand UO_307 (O_307,N_24955,N_24827);
nand UO_308 (O_308,N_24930,N_24847);
and UO_309 (O_309,N_24951,N_24806);
nand UO_310 (O_310,N_24563,N_24914);
and UO_311 (O_311,N_24943,N_24940);
xor UO_312 (O_312,N_24877,N_24643);
or UO_313 (O_313,N_24585,N_24850);
or UO_314 (O_314,N_24473,N_24665);
nor UO_315 (O_315,N_24968,N_24732);
nand UO_316 (O_316,N_24872,N_24609);
xnor UO_317 (O_317,N_24556,N_24788);
xnor UO_318 (O_318,N_24897,N_24659);
or UO_319 (O_319,N_24511,N_24505);
nor UO_320 (O_320,N_24962,N_24476);
and UO_321 (O_321,N_24650,N_24666);
or UO_322 (O_322,N_24917,N_24882);
or UO_323 (O_323,N_24540,N_24730);
xnor UO_324 (O_324,N_24809,N_24587);
and UO_325 (O_325,N_24386,N_24944);
nor UO_326 (O_326,N_24749,N_24811);
nand UO_327 (O_327,N_24860,N_24990);
xor UO_328 (O_328,N_24379,N_24695);
or UO_329 (O_329,N_24419,N_24538);
and UO_330 (O_330,N_24585,N_24503);
or UO_331 (O_331,N_24448,N_24851);
nor UO_332 (O_332,N_24872,N_24519);
nor UO_333 (O_333,N_24929,N_24706);
or UO_334 (O_334,N_24432,N_24926);
xnor UO_335 (O_335,N_24878,N_24865);
nor UO_336 (O_336,N_24750,N_24556);
and UO_337 (O_337,N_24508,N_24847);
nand UO_338 (O_338,N_24806,N_24408);
or UO_339 (O_339,N_24920,N_24654);
or UO_340 (O_340,N_24881,N_24606);
nand UO_341 (O_341,N_24988,N_24987);
xnor UO_342 (O_342,N_24761,N_24404);
nor UO_343 (O_343,N_24989,N_24810);
or UO_344 (O_344,N_24743,N_24990);
or UO_345 (O_345,N_24938,N_24632);
and UO_346 (O_346,N_24725,N_24871);
and UO_347 (O_347,N_24859,N_24468);
nand UO_348 (O_348,N_24993,N_24957);
or UO_349 (O_349,N_24998,N_24414);
nand UO_350 (O_350,N_24504,N_24383);
and UO_351 (O_351,N_24691,N_24458);
nand UO_352 (O_352,N_24964,N_24985);
nor UO_353 (O_353,N_24898,N_24419);
nor UO_354 (O_354,N_24756,N_24777);
or UO_355 (O_355,N_24874,N_24726);
xor UO_356 (O_356,N_24617,N_24765);
nor UO_357 (O_357,N_24659,N_24418);
nand UO_358 (O_358,N_24461,N_24812);
nor UO_359 (O_359,N_24985,N_24836);
and UO_360 (O_360,N_24861,N_24477);
or UO_361 (O_361,N_24601,N_24517);
or UO_362 (O_362,N_24973,N_24497);
nand UO_363 (O_363,N_24816,N_24903);
and UO_364 (O_364,N_24984,N_24883);
or UO_365 (O_365,N_24711,N_24476);
nor UO_366 (O_366,N_24785,N_24747);
nand UO_367 (O_367,N_24476,N_24935);
or UO_368 (O_368,N_24747,N_24796);
xnor UO_369 (O_369,N_24887,N_24773);
and UO_370 (O_370,N_24720,N_24988);
and UO_371 (O_371,N_24875,N_24697);
nand UO_372 (O_372,N_24830,N_24397);
and UO_373 (O_373,N_24724,N_24765);
xnor UO_374 (O_374,N_24680,N_24919);
or UO_375 (O_375,N_24593,N_24978);
nand UO_376 (O_376,N_24930,N_24851);
nand UO_377 (O_377,N_24591,N_24622);
or UO_378 (O_378,N_24386,N_24465);
xor UO_379 (O_379,N_24735,N_24593);
xnor UO_380 (O_380,N_24650,N_24898);
nor UO_381 (O_381,N_24687,N_24652);
xor UO_382 (O_382,N_24539,N_24403);
xnor UO_383 (O_383,N_24422,N_24794);
xnor UO_384 (O_384,N_24593,N_24918);
xor UO_385 (O_385,N_24848,N_24886);
nor UO_386 (O_386,N_24752,N_24742);
nand UO_387 (O_387,N_24970,N_24451);
or UO_388 (O_388,N_24939,N_24562);
or UO_389 (O_389,N_24739,N_24705);
xor UO_390 (O_390,N_24713,N_24634);
nor UO_391 (O_391,N_24977,N_24626);
or UO_392 (O_392,N_24636,N_24663);
or UO_393 (O_393,N_24847,N_24496);
nand UO_394 (O_394,N_24681,N_24916);
xnor UO_395 (O_395,N_24612,N_24436);
and UO_396 (O_396,N_24674,N_24472);
xnor UO_397 (O_397,N_24704,N_24540);
nand UO_398 (O_398,N_24422,N_24559);
nand UO_399 (O_399,N_24446,N_24679);
nand UO_400 (O_400,N_24938,N_24977);
xor UO_401 (O_401,N_24649,N_24807);
and UO_402 (O_402,N_24442,N_24957);
nor UO_403 (O_403,N_24447,N_24535);
xor UO_404 (O_404,N_24438,N_24894);
or UO_405 (O_405,N_24910,N_24921);
nand UO_406 (O_406,N_24721,N_24462);
and UO_407 (O_407,N_24639,N_24710);
nor UO_408 (O_408,N_24412,N_24727);
or UO_409 (O_409,N_24875,N_24717);
and UO_410 (O_410,N_24978,N_24570);
and UO_411 (O_411,N_24562,N_24533);
and UO_412 (O_412,N_24702,N_24838);
nand UO_413 (O_413,N_24407,N_24810);
xor UO_414 (O_414,N_24678,N_24899);
xnor UO_415 (O_415,N_24524,N_24590);
or UO_416 (O_416,N_24456,N_24464);
xnor UO_417 (O_417,N_24857,N_24647);
or UO_418 (O_418,N_24762,N_24672);
nand UO_419 (O_419,N_24504,N_24847);
nor UO_420 (O_420,N_24568,N_24404);
or UO_421 (O_421,N_24564,N_24847);
xor UO_422 (O_422,N_24740,N_24599);
xnor UO_423 (O_423,N_24796,N_24571);
nor UO_424 (O_424,N_24384,N_24537);
xnor UO_425 (O_425,N_24859,N_24438);
nand UO_426 (O_426,N_24935,N_24961);
nor UO_427 (O_427,N_24508,N_24627);
or UO_428 (O_428,N_24584,N_24983);
or UO_429 (O_429,N_24577,N_24950);
or UO_430 (O_430,N_24647,N_24898);
nand UO_431 (O_431,N_24489,N_24404);
nand UO_432 (O_432,N_24708,N_24893);
and UO_433 (O_433,N_24510,N_24613);
or UO_434 (O_434,N_24826,N_24805);
and UO_435 (O_435,N_24739,N_24834);
nand UO_436 (O_436,N_24904,N_24892);
xnor UO_437 (O_437,N_24439,N_24795);
nand UO_438 (O_438,N_24928,N_24864);
nand UO_439 (O_439,N_24496,N_24939);
nand UO_440 (O_440,N_24787,N_24953);
nand UO_441 (O_441,N_24922,N_24376);
and UO_442 (O_442,N_24504,N_24496);
nor UO_443 (O_443,N_24707,N_24649);
nand UO_444 (O_444,N_24817,N_24836);
nor UO_445 (O_445,N_24892,N_24605);
nand UO_446 (O_446,N_24505,N_24805);
and UO_447 (O_447,N_24949,N_24574);
and UO_448 (O_448,N_24555,N_24759);
nand UO_449 (O_449,N_24746,N_24900);
or UO_450 (O_450,N_24777,N_24754);
nand UO_451 (O_451,N_24818,N_24780);
xnor UO_452 (O_452,N_24831,N_24602);
nand UO_453 (O_453,N_24588,N_24401);
xor UO_454 (O_454,N_24625,N_24802);
nand UO_455 (O_455,N_24834,N_24523);
and UO_456 (O_456,N_24989,N_24403);
nand UO_457 (O_457,N_24453,N_24534);
and UO_458 (O_458,N_24670,N_24613);
nand UO_459 (O_459,N_24699,N_24773);
nor UO_460 (O_460,N_24441,N_24657);
nor UO_461 (O_461,N_24899,N_24384);
and UO_462 (O_462,N_24674,N_24463);
xor UO_463 (O_463,N_24630,N_24939);
or UO_464 (O_464,N_24826,N_24871);
xnor UO_465 (O_465,N_24897,N_24794);
nand UO_466 (O_466,N_24697,N_24437);
and UO_467 (O_467,N_24880,N_24843);
nor UO_468 (O_468,N_24889,N_24865);
xnor UO_469 (O_469,N_24766,N_24531);
or UO_470 (O_470,N_24538,N_24894);
nor UO_471 (O_471,N_24436,N_24967);
or UO_472 (O_472,N_24687,N_24922);
xor UO_473 (O_473,N_24953,N_24405);
or UO_474 (O_474,N_24674,N_24800);
or UO_475 (O_475,N_24427,N_24663);
nor UO_476 (O_476,N_24482,N_24725);
or UO_477 (O_477,N_24841,N_24947);
and UO_478 (O_478,N_24693,N_24787);
nand UO_479 (O_479,N_24992,N_24491);
nor UO_480 (O_480,N_24802,N_24743);
xnor UO_481 (O_481,N_24559,N_24826);
or UO_482 (O_482,N_24834,N_24782);
and UO_483 (O_483,N_24482,N_24879);
nor UO_484 (O_484,N_24952,N_24548);
xnor UO_485 (O_485,N_24546,N_24854);
xor UO_486 (O_486,N_24755,N_24893);
nor UO_487 (O_487,N_24959,N_24990);
nor UO_488 (O_488,N_24392,N_24459);
and UO_489 (O_489,N_24590,N_24776);
nor UO_490 (O_490,N_24557,N_24769);
or UO_491 (O_491,N_24655,N_24567);
or UO_492 (O_492,N_24853,N_24914);
and UO_493 (O_493,N_24632,N_24515);
nor UO_494 (O_494,N_24916,N_24653);
and UO_495 (O_495,N_24704,N_24607);
nand UO_496 (O_496,N_24937,N_24655);
and UO_497 (O_497,N_24459,N_24999);
xnor UO_498 (O_498,N_24566,N_24533);
xnor UO_499 (O_499,N_24546,N_24658);
nand UO_500 (O_500,N_24500,N_24719);
or UO_501 (O_501,N_24466,N_24739);
xor UO_502 (O_502,N_24388,N_24681);
and UO_503 (O_503,N_24803,N_24939);
or UO_504 (O_504,N_24404,N_24668);
nand UO_505 (O_505,N_24583,N_24986);
xnor UO_506 (O_506,N_24864,N_24999);
and UO_507 (O_507,N_24875,N_24588);
nor UO_508 (O_508,N_24644,N_24741);
or UO_509 (O_509,N_24597,N_24720);
and UO_510 (O_510,N_24831,N_24848);
nand UO_511 (O_511,N_24578,N_24911);
or UO_512 (O_512,N_24687,N_24700);
xor UO_513 (O_513,N_24809,N_24756);
nor UO_514 (O_514,N_24513,N_24580);
and UO_515 (O_515,N_24423,N_24699);
and UO_516 (O_516,N_24427,N_24983);
and UO_517 (O_517,N_24507,N_24910);
or UO_518 (O_518,N_24503,N_24473);
or UO_519 (O_519,N_24558,N_24507);
nand UO_520 (O_520,N_24919,N_24681);
xor UO_521 (O_521,N_24387,N_24705);
xor UO_522 (O_522,N_24685,N_24647);
nor UO_523 (O_523,N_24499,N_24670);
or UO_524 (O_524,N_24523,N_24936);
nand UO_525 (O_525,N_24709,N_24877);
nand UO_526 (O_526,N_24502,N_24743);
xnor UO_527 (O_527,N_24610,N_24428);
xnor UO_528 (O_528,N_24780,N_24413);
nor UO_529 (O_529,N_24555,N_24929);
xor UO_530 (O_530,N_24389,N_24490);
nor UO_531 (O_531,N_24525,N_24865);
xor UO_532 (O_532,N_24741,N_24545);
nand UO_533 (O_533,N_24866,N_24892);
xnor UO_534 (O_534,N_24451,N_24648);
or UO_535 (O_535,N_24909,N_24998);
or UO_536 (O_536,N_24440,N_24673);
xnor UO_537 (O_537,N_24617,N_24932);
xor UO_538 (O_538,N_24717,N_24847);
or UO_539 (O_539,N_24657,N_24846);
nor UO_540 (O_540,N_24893,N_24926);
and UO_541 (O_541,N_24608,N_24505);
and UO_542 (O_542,N_24713,N_24969);
nand UO_543 (O_543,N_24727,N_24562);
and UO_544 (O_544,N_24412,N_24462);
nor UO_545 (O_545,N_24526,N_24494);
and UO_546 (O_546,N_24851,N_24584);
or UO_547 (O_547,N_24981,N_24514);
nor UO_548 (O_548,N_24482,N_24889);
or UO_549 (O_549,N_24644,N_24615);
and UO_550 (O_550,N_24854,N_24910);
or UO_551 (O_551,N_24693,N_24830);
nor UO_552 (O_552,N_24806,N_24520);
nand UO_553 (O_553,N_24877,N_24715);
or UO_554 (O_554,N_24750,N_24656);
or UO_555 (O_555,N_24521,N_24448);
or UO_556 (O_556,N_24841,N_24560);
nand UO_557 (O_557,N_24673,N_24504);
nor UO_558 (O_558,N_24431,N_24550);
nor UO_559 (O_559,N_24973,N_24622);
nand UO_560 (O_560,N_24783,N_24417);
or UO_561 (O_561,N_24838,N_24405);
and UO_562 (O_562,N_24565,N_24756);
nand UO_563 (O_563,N_24700,N_24616);
and UO_564 (O_564,N_24714,N_24590);
nor UO_565 (O_565,N_24809,N_24824);
or UO_566 (O_566,N_24417,N_24684);
and UO_567 (O_567,N_24732,N_24759);
nand UO_568 (O_568,N_24448,N_24429);
xnor UO_569 (O_569,N_24465,N_24629);
and UO_570 (O_570,N_24573,N_24553);
and UO_571 (O_571,N_24663,N_24378);
xor UO_572 (O_572,N_24764,N_24832);
or UO_573 (O_573,N_24612,N_24869);
xnor UO_574 (O_574,N_24906,N_24377);
nand UO_575 (O_575,N_24575,N_24970);
or UO_576 (O_576,N_24605,N_24588);
and UO_577 (O_577,N_24924,N_24662);
nor UO_578 (O_578,N_24877,N_24561);
and UO_579 (O_579,N_24463,N_24393);
nor UO_580 (O_580,N_24912,N_24744);
and UO_581 (O_581,N_24445,N_24620);
xnor UO_582 (O_582,N_24956,N_24731);
xnor UO_583 (O_583,N_24688,N_24971);
nor UO_584 (O_584,N_24462,N_24384);
and UO_585 (O_585,N_24774,N_24602);
nand UO_586 (O_586,N_24522,N_24840);
and UO_587 (O_587,N_24669,N_24515);
and UO_588 (O_588,N_24995,N_24969);
or UO_589 (O_589,N_24943,N_24577);
xor UO_590 (O_590,N_24788,N_24633);
xor UO_591 (O_591,N_24781,N_24796);
or UO_592 (O_592,N_24811,N_24584);
nor UO_593 (O_593,N_24571,N_24822);
or UO_594 (O_594,N_24547,N_24661);
or UO_595 (O_595,N_24605,N_24987);
nand UO_596 (O_596,N_24817,N_24605);
nand UO_597 (O_597,N_24498,N_24908);
and UO_598 (O_598,N_24881,N_24786);
xnor UO_599 (O_599,N_24941,N_24525);
nor UO_600 (O_600,N_24884,N_24783);
or UO_601 (O_601,N_24995,N_24884);
or UO_602 (O_602,N_24419,N_24862);
nand UO_603 (O_603,N_24941,N_24546);
and UO_604 (O_604,N_24809,N_24911);
nor UO_605 (O_605,N_24621,N_24830);
or UO_606 (O_606,N_24806,N_24792);
nor UO_607 (O_607,N_24980,N_24565);
nor UO_608 (O_608,N_24577,N_24677);
and UO_609 (O_609,N_24503,N_24533);
or UO_610 (O_610,N_24983,N_24539);
nand UO_611 (O_611,N_24380,N_24947);
and UO_612 (O_612,N_24852,N_24529);
and UO_613 (O_613,N_24541,N_24715);
nand UO_614 (O_614,N_24392,N_24890);
xor UO_615 (O_615,N_24954,N_24742);
and UO_616 (O_616,N_24559,N_24965);
or UO_617 (O_617,N_24670,N_24896);
or UO_618 (O_618,N_24477,N_24566);
nand UO_619 (O_619,N_24577,N_24482);
nand UO_620 (O_620,N_24771,N_24527);
nor UO_621 (O_621,N_24519,N_24905);
or UO_622 (O_622,N_24929,N_24538);
nor UO_623 (O_623,N_24991,N_24612);
and UO_624 (O_624,N_24853,N_24851);
nand UO_625 (O_625,N_24398,N_24450);
nor UO_626 (O_626,N_24871,N_24883);
xor UO_627 (O_627,N_24843,N_24584);
or UO_628 (O_628,N_24585,N_24805);
xor UO_629 (O_629,N_24402,N_24603);
xnor UO_630 (O_630,N_24724,N_24618);
xor UO_631 (O_631,N_24418,N_24469);
or UO_632 (O_632,N_24661,N_24862);
xor UO_633 (O_633,N_24489,N_24672);
nand UO_634 (O_634,N_24650,N_24445);
and UO_635 (O_635,N_24652,N_24757);
or UO_636 (O_636,N_24479,N_24971);
or UO_637 (O_637,N_24452,N_24909);
or UO_638 (O_638,N_24401,N_24465);
nand UO_639 (O_639,N_24710,N_24835);
and UO_640 (O_640,N_24957,N_24666);
and UO_641 (O_641,N_24437,N_24855);
nand UO_642 (O_642,N_24886,N_24441);
or UO_643 (O_643,N_24464,N_24419);
xnor UO_644 (O_644,N_24796,N_24861);
and UO_645 (O_645,N_24425,N_24914);
xnor UO_646 (O_646,N_24889,N_24864);
xor UO_647 (O_647,N_24574,N_24689);
and UO_648 (O_648,N_24831,N_24404);
and UO_649 (O_649,N_24761,N_24417);
xor UO_650 (O_650,N_24852,N_24758);
nand UO_651 (O_651,N_24657,N_24774);
nand UO_652 (O_652,N_24999,N_24404);
xnor UO_653 (O_653,N_24708,N_24408);
nor UO_654 (O_654,N_24904,N_24506);
and UO_655 (O_655,N_24841,N_24783);
nor UO_656 (O_656,N_24861,N_24534);
nand UO_657 (O_657,N_24571,N_24397);
or UO_658 (O_658,N_24792,N_24733);
or UO_659 (O_659,N_24426,N_24469);
xor UO_660 (O_660,N_24939,N_24403);
or UO_661 (O_661,N_24764,N_24396);
nor UO_662 (O_662,N_24832,N_24746);
and UO_663 (O_663,N_24993,N_24631);
xor UO_664 (O_664,N_24654,N_24501);
nor UO_665 (O_665,N_24542,N_24561);
or UO_666 (O_666,N_24580,N_24965);
or UO_667 (O_667,N_24545,N_24525);
xor UO_668 (O_668,N_24403,N_24729);
and UO_669 (O_669,N_24939,N_24525);
nor UO_670 (O_670,N_24700,N_24685);
xnor UO_671 (O_671,N_24816,N_24826);
nand UO_672 (O_672,N_24676,N_24731);
and UO_673 (O_673,N_24410,N_24878);
and UO_674 (O_674,N_24482,N_24692);
or UO_675 (O_675,N_24776,N_24710);
nand UO_676 (O_676,N_24648,N_24622);
and UO_677 (O_677,N_24383,N_24458);
or UO_678 (O_678,N_24970,N_24380);
and UO_679 (O_679,N_24964,N_24502);
nand UO_680 (O_680,N_24868,N_24640);
and UO_681 (O_681,N_24581,N_24426);
xnor UO_682 (O_682,N_24704,N_24864);
or UO_683 (O_683,N_24662,N_24779);
xor UO_684 (O_684,N_24903,N_24417);
or UO_685 (O_685,N_24983,N_24679);
nand UO_686 (O_686,N_24953,N_24615);
xor UO_687 (O_687,N_24852,N_24694);
and UO_688 (O_688,N_24535,N_24660);
or UO_689 (O_689,N_24988,N_24551);
nor UO_690 (O_690,N_24677,N_24544);
or UO_691 (O_691,N_24431,N_24514);
xor UO_692 (O_692,N_24592,N_24509);
nand UO_693 (O_693,N_24453,N_24460);
and UO_694 (O_694,N_24826,N_24726);
xnor UO_695 (O_695,N_24915,N_24890);
or UO_696 (O_696,N_24857,N_24498);
nand UO_697 (O_697,N_24837,N_24390);
or UO_698 (O_698,N_24882,N_24821);
nor UO_699 (O_699,N_24717,N_24896);
xnor UO_700 (O_700,N_24404,N_24475);
and UO_701 (O_701,N_24873,N_24401);
nor UO_702 (O_702,N_24554,N_24905);
nor UO_703 (O_703,N_24444,N_24717);
nand UO_704 (O_704,N_24894,N_24818);
nand UO_705 (O_705,N_24542,N_24425);
and UO_706 (O_706,N_24971,N_24425);
and UO_707 (O_707,N_24832,N_24740);
nor UO_708 (O_708,N_24612,N_24414);
nand UO_709 (O_709,N_24951,N_24521);
nor UO_710 (O_710,N_24706,N_24774);
nor UO_711 (O_711,N_24543,N_24929);
or UO_712 (O_712,N_24931,N_24816);
nor UO_713 (O_713,N_24433,N_24890);
and UO_714 (O_714,N_24554,N_24838);
xnor UO_715 (O_715,N_24622,N_24889);
nor UO_716 (O_716,N_24998,N_24994);
xor UO_717 (O_717,N_24876,N_24433);
or UO_718 (O_718,N_24879,N_24903);
and UO_719 (O_719,N_24951,N_24492);
nand UO_720 (O_720,N_24750,N_24700);
xnor UO_721 (O_721,N_24614,N_24832);
nor UO_722 (O_722,N_24423,N_24387);
and UO_723 (O_723,N_24750,N_24722);
or UO_724 (O_724,N_24409,N_24945);
nor UO_725 (O_725,N_24493,N_24387);
and UO_726 (O_726,N_24390,N_24508);
nand UO_727 (O_727,N_24396,N_24519);
nand UO_728 (O_728,N_24525,N_24698);
nand UO_729 (O_729,N_24800,N_24646);
nand UO_730 (O_730,N_24979,N_24415);
nand UO_731 (O_731,N_24676,N_24393);
xnor UO_732 (O_732,N_24589,N_24800);
xnor UO_733 (O_733,N_24896,N_24792);
nor UO_734 (O_734,N_24755,N_24833);
xnor UO_735 (O_735,N_24793,N_24788);
nor UO_736 (O_736,N_24414,N_24855);
xnor UO_737 (O_737,N_24827,N_24976);
xnor UO_738 (O_738,N_24752,N_24496);
or UO_739 (O_739,N_24426,N_24613);
nor UO_740 (O_740,N_24932,N_24675);
or UO_741 (O_741,N_24585,N_24943);
or UO_742 (O_742,N_24772,N_24642);
xnor UO_743 (O_743,N_24653,N_24902);
xnor UO_744 (O_744,N_24520,N_24937);
nor UO_745 (O_745,N_24897,N_24493);
xnor UO_746 (O_746,N_24800,N_24566);
xor UO_747 (O_747,N_24648,N_24867);
nand UO_748 (O_748,N_24426,N_24865);
and UO_749 (O_749,N_24709,N_24540);
or UO_750 (O_750,N_24588,N_24380);
xnor UO_751 (O_751,N_24647,N_24814);
and UO_752 (O_752,N_24538,N_24916);
and UO_753 (O_753,N_24456,N_24886);
nand UO_754 (O_754,N_24933,N_24908);
and UO_755 (O_755,N_24564,N_24693);
nand UO_756 (O_756,N_24482,N_24531);
xor UO_757 (O_757,N_24792,N_24862);
nor UO_758 (O_758,N_24657,N_24669);
nand UO_759 (O_759,N_24512,N_24399);
and UO_760 (O_760,N_24593,N_24446);
and UO_761 (O_761,N_24527,N_24523);
xor UO_762 (O_762,N_24807,N_24605);
or UO_763 (O_763,N_24692,N_24967);
and UO_764 (O_764,N_24640,N_24606);
xnor UO_765 (O_765,N_24887,N_24527);
or UO_766 (O_766,N_24493,N_24842);
nor UO_767 (O_767,N_24932,N_24727);
nor UO_768 (O_768,N_24780,N_24865);
or UO_769 (O_769,N_24555,N_24488);
and UO_770 (O_770,N_24891,N_24670);
nand UO_771 (O_771,N_24687,N_24857);
xnor UO_772 (O_772,N_24881,N_24439);
nand UO_773 (O_773,N_24634,N_24740);
or UO_774 (O_774,N_24817,N_24890);
or UO_775 (O_775,N_24770,N_24838);
nand UO_776 (O_776,N_24595,N_24934);
xnor UO_777 (O_777,N_24543,N_24520);
or UO_778 (O_778,N_24681,N_24611);
nor UO_779 (O_779,N_24990,N_24547);
nand UO_780 (O_780,N_24770,N_24482);
nor UO_781 (O_781,N_24433,N_24553);
xnor UO_782 (O_782,N_24727,N_24778);
or UO_783 (O_783,N_24567,N_24662);
xor UO_784 (O_784,N_24522,N_24687);
nand UO_785 (O_785,N_24996,N_24715);
xnor UO_786 (O_786,N_24507,N_24706);
xnor UO_787 (O_787,N_24502,N_24961);
nand UO_788 (O_788,N_24401,N_24720);
nor UO_789 (O_789,N_24967,N_24471);
nor UO_790 (O_790,N_24552,N_24777);
nor UO_791 (O_791,N_24926,N_24383);
nor UO_792 (O_792,N_24992,N_24575);
nand UO_793 (O_793,N_24819,N_24910);
nand UO_794 (O_794,N_24508,N_24427);
and UO_795 (O_795,N_24855,N_24656);
nand UO_796 (O_796,N_24731,N_24542);
xnor UO_797 (O_797,N_24503,N_24910);
nand UO_798 (O_798,N_24890,N_24399);
xnor UO_799 (O_799,N_24429,N_24642);
xor UO_800 (O_800,N_24911,N_24865);
nor UO_801 (O_801,N_24640,N_24502);
nand UO_802 (O_802,N_24787,N_24698);
and UO_803 (O_803,N_24758,N_24604);
nor UO_804 (O_804,N_24703,N_24573);
nand UO_805 (O_805,N_24956,N_24598);
nand UO_806 (O_806,N_24768,N_24911);
and UO_807 (O_807,N_24473,N_24587);
or UO_808 (O_808,N_24835,N_24752);
nor UO_809 (O_809,N_24785,N_24866);
nand UO_810 (O_810,N_24788,N_24701);
or UO_811 (O_811,N_24498,N_24873);
nor UO_812 (O_812,N_24643,N_24929);
xnor UO_813 (O_813,N_24693,N_24521);
or UO_814 (O_814,N_24450,N_24463);
xor UO_815 (O_815,N_24428,N_24476);
or UO_816 (O_816,N_24773,N_24997);
and UO_817 (O_817,N_24385,N_24516);
or UO_818 (O_818,N_24788,N_24985);
or UO_819 (O_819,N_24731,N_24628);
and UO_820 (O_820,N_24435,N_24845);
and UO_821 (O_821,N_24540,N_24916);
nand UO_822 (O_822,N_24966,N_24918);
nor UO_823 (O_823,N_24459,N_24942);
xnor UO_824 (O_824,N_24856,N_24797);
nand UO_825 (O_825,N_24903,N_24608);
nor UO_826 (O_826,N_24588,N_24630);
nor UO_827 (O_827,N_24528,N_24852);
and UO_828 (O_828,N_24494,N_24772);
nor UO_829 (O_829,N_24802,N_24383);
or UO_830 (O_830,N_24996,N_24601);
xor UO_831 (O_831,N_24952,N_24963);
and UO_832 (O_832,N_24972,N_24958);
or UO_833 (O_833,N_24464,N_24731);
and UO_834 (O_834,N_24757,N_24873);
xor UO_835 (O_835,N_24556,N_24698);
xnor UO_836 (O_836,N_24468,N_24478);
xor UO_837 (O_837,N_24812,N_24653);
nand UO_838 (O_838,N_24393,N_24816);
xnor UO_839 (O_839,N_24935,N_24926);
nor UO_840 (O_840,N_24910,N_24874);
nand UO_841 (O_841,N_24996,N_24963);
xnor UO_842 (O_842,N_24957,N_24556);
or UO_843 (O_843,N_24440,N_24631);
or UO_844 (O_844,N_24933,N_24913);
and UO_845 (O_845,N_24831,N_24671);
nand UO_846 (O_846,N_24593,N_24424);
nor UO_847 (O_847,N_24549,N_24968);
or UO_848 (O_848,N_24782,N_24993);
nor UO_849 (O_849,N_24848,N_24384);
nor UO_850 (O_850,N_24568,N_24461);
or UO_851 (O_851,N_24381,N_24811);
and UO_852 (O_852,N_24644,N_24777);
nor UO_853 (O_853,N_24847,N_24608);
xor UO_854 (O_854,N_24559,N_24589);
or UO_855 (O_855,N_24995,N_24415);
nor UO_856 (O_856,N_24781,N_24951);
nor UO_857 (O_857,N_24495,N_24397);
nor UO_858 (O_858,N_24651,N_24988);
and UO_859 (O_859,N_24497,N_24509);
or UO_860 (O_860,N_24958,N_24709);
nor UO_861 (O_861,N_24775,N_24972);
nor UO_862 (O_862,N_24432,N_24521);
xnor UO_863 (O_863,N_24830,N_24834);
or UO_864 (O_864,N_24430,N_24584);
or UO_865 (O_865,N_24744,N_24527);
xor UO_866 (O_866,N_24586,N_24579);
and UO_867 (O_867,N_24604,N_24714);
nor UO_868 (O_868,N_24935,N_24727);
nor UO_869 (O_869,N_24641,N_24690);
nor UO_870 (O_870,N_24795,N_24760);
nor UO_871 (O_871,N_24732,N_24934);
nand UO_872 (O_872,N_24622,N_24678);
and UO_873 (O_873,N_24411,N_24572);
or UO_874 (O_874,N_24752,N_24422);
xor UO_875 (O_875,N_24643,N_24792);
or UO_876 (O_876,N_24946,N_24852);
nor UO_877 (O_877,N_24904,N_24835);
nand UO_878 (O_878,N_24889,N_24599);
nor UO_879 (O_879,N_24438,N_24855);
and UO_880 (O_880,N_24650,N_24879);
and UO_881 (O_881,N_24530,N_24650);
xor UO_882 (O_882,N_24446,N_24643);
and UO_883 (O_883,N_24784,N_24773);
nor UO_884 (O_884,N_24993,N_24508);
nor UO_885 (O_885,N_24941,N_24433);
xnor UO_886 (O_886,N_24684,N_24561);
nand UO_887 (O_887,N_24859,N_24609);
nor UO_888 (O_888,N_24879,N_24421);
and UO_889 (O_889,N_24758,N_24995);
xnor UO_890 (O_890,N_24509,N_24833);
and UO_891 (O_891,N_24725,N_24375);
nand UO_892 (O_892,N_24745,N_24438);
xor UO_893 (O_893,N_24414,N_24662);
or UO_894 (O_894,N_24795,N_24567);
or UO_895 (O_895,N_24759,N_24910);
nor UO_896 (O_896,N_24477,N_24598);
nor UO_897 (O_897,N_24576,N_24743);
xnor UO_898 (O_898,N_24975,N_24568);
xor UO_899 (O_899,N_24993,N_24657);
or UO_900 (O_900,N_24795,N_24632);
nand UO_901 (O_901,N_24702,N_24753);
and UO_902 (O_902,N_24909,N_24424);
nand UO_903 (O_903,N_24380,N_24724);
xor UO_904 (O_904,N_24660,N_24411);
or UO_905 (O_905,N_24401,N_24413);
nor UO_906 (O_906,N_24721,N_24524);
nor UO_907 (O_907,N_24491,N_24459);
xnor UO_908 (O_908,N_24738,N_24422);
or UO_909 (O_909,N_24878,N_24634);
and UO_910 (O_910,N_24750,N_24789);
and UO_911 (O_911,N_24778,N_24978);
and UO_912 (O_912,N_24665,N_24553);
nand UO_913 (O_913,N_24991,N_24728);
and UO_914 (O_914,N_24746,N_24583);
or UO_915 (O_915,N_24759,N_24572);
and UO_916 (O_916,N_24628,N_24681);
xnor UO_917 (O_917,N_24385,N_24699);
xor UO_918 (O_918,N_24836,N_24705);
and UO_919 (O_919,N_24574,N_24765);
xnor UO_920 (O_920,N_24737,N_24603);
and UO_921 (O_921,N_24773,N_24855);
or UO_922 (O_922,N_24757,N_24816);
nor UO_923 (O_923,N_24991,N_24460);
or UO_924 (O_924,N_24624,N_24630);
xor UO_925 (O_925,N_24826,N_24451);
and UO_926 (O_926,N_24420,N_24889);
nor UO_927 (O_927,N_24895,N_24699);
or UO_928 (O_928,N_24516,N_24566);
xnor UO_929 (O_929,N_24833,N_24475);
nor UO_930 (O_930,N_24530,N_24777);
nor UO_931 (O_931,N_24872,N_24874);
and UO_932 (O_932,N_24478,N_24905);
nor UO_933 (O_933,N_24908,N_24871);
or UO_934 (O_934,N_24766,N_24896);
nor UO_935 (O_935,N_24792,N_24661);
or UO_936 (O_936,N_24863,N_24801);
nand UO_937 (O_937,N_24759,N_24633);
nor UO_938 (O_938,N_24482,N_24489);
nor UO_939 (O_939,N_24975,N_24786);
xor UO_940 (O_940,N_24947,N_24846);
nor UO_941 (O_941,N_24668,N_24476);
nor UO_942 (O_942,N_24543,N_24830);
and UO_943 (O_943,N_24529,N_24959);
xnor UO_944 (O_944,N_24495,N_24717);
or UO_945 (O_945,N_24484,N_24621);
nor UO_946 (O_946,N_24462,N_24518);
nor UO_947 (O_947,N_24987,N_24581);
or UO_948 (O_948,N_24522,N_24586);
xor UO_949 (O_949,N_24502,N_24957);
xor UO_950 (O_950,N_24776,N_24975);
and UO_951 (O_951,N_24926,N_24822);
or UO_952 (O_952,N_24688,N_24835);
nand UO_953 (O_953,N_24514,N_24921);
or UO_954 (O_954,N_24996,N_24917);
and UO_955 (O_955,N_24410,N_24957);
and UO_956 (O_956,N_24743,N_24758);
nor UO_957 (O_957,N_24519,N_24744);
nor UO_958 (O_958,N_24476,N_24709);
nor UO_959 (O_959,N_24918,N_24973);
and UO_960 (O_960,N_24704,N_24949);
xor UO_961 (O_961,N_24942,N_24787);
nor UO_962 (O_962,N_24627,N_24395);
xnor UO_963 (O_963,N_24933,N_24630);
nor UO_964 (O_964,N_24551,N_24912);
nor UO_965 (O_965,N_24550,N_24978);
nand UO_966 (O_966,N_24417,N_24654);
and UO_967 (O_967,N_24950,N_24683);
nor UO_968 (O_968,N_24568,N_24999);
nor UO_969 (O_969,N_24738,N_24402);
nor UO_970 (O_970,N_24893,N_24593);
nand UO_971 (O_971,N_24541,N_24597);
or UO_972 (O_972,N_24952,N_24664);
and UO_973 (O_973,N_24951,N_24467);
xor UO_974 (O_974,N_24745,N_24947);
nor UO_975 (O_975,N_24695,N_24674);
xor UO_976 (O_976,N_24722,N_24518);
or UO_977 (O_977,N_24432,N_24434);
and UO_978 (O_978,N_24884,N_24588);
or UO_979 (O_979,N_24453,N_24925);
nand UO_980 (O_980,N_24537,N_24525);
or UO_981 (O_981,N_24943,N_24544);
xnor UO_982 (O_982,N_24989,N_24932);
xor UO_983 (O_983,N_24842,N_24455);
or UO_984 (O_984,N_24475,N_24387);
xnor UO_985 (O_985,N_24392,N_24667);
nand UO_986 (O_986,N_24589,N_24484);
or UO_987 (O_987,N_24386,N_24810);
xor UO_988 (O_988,N_24679,N_24479);
nor UO_989 (O_989,N_24453,N_24808);
xnor UO_990 (O_990,N_24396,N_24824);
nand UO_991 (O_991,N_24896,N_24508);
nor UO_992 (O_992,N_24589,N_24729);
nand UO_993 (O_993,N_24761,N_24888);
nor UO_994 (O_994,N_24428,N_24592);
nor UO_995 (O_995,N_24736,N_24708);
nor UO_996 (O_996,N_24394,N_24599);
nand UO_997 (O_997,N_24896,N_24892);
nor UO_998 (O_998,N_24631,N_24873);
nand UO_999 (O_999,N_24748,N_24667);
nor UO_1000 (O_1000,N_24916,N_24697);
nand UO_1001 (O_1001,N_24895,N_24481);
nand UO_1002 (O_1002,N_24912,N_24544);
nand UO_1003 (O_1003,N_24533,N_24635);
nand UO_1004 (O_1004,N_24705,N_24512);
or UO_1005 (O_1005,N_24446,N_24481);
or UO_1006 (O_1006,N_24763,N_24732);
xnor UO_1007 (O_1007,N_24673,N_24415);
nor UO_1008 (O_1008,N_24730,N_24674);
nand UO_1009 (O_1009,N_24775,N_24452);
nand UO_1010 (O_1010,N_24897,N_24499);
or UO_1011 (O_1011,N_24560,N_24799);
nand UO_1012 (O_1012,N_24665,N_24391);
nor UO_1013 (O_1013,N_24909,N_24381);
nand UO_1014 (O_1014,N_24581,N_24509);
xnor UO_1015 (O_1015,N_24926,N_24806);
nand UO_1016 (O_1016,N_24941,N_24870);
xnor UO_1017 (O_1017,N_24634,N_24841);
nand UO_1018 (O_1018,N_24878,N_24768);
nand UO_1019 (O_1019,N_24648,N_24376);
nor UO_1020 (O_1020,N_24425,N_24970);
or UO_1021 (O_1021,N_24436,N_24497);
nand UO_1022 (O_1022,N_24707,N_24488);
nor UO_1023 (O_1023,N_24623,N_24774);
nand UO_1024 (O_1024,N_24690,N_24998);
xor UO_1025 (O_1025,N_24793,N_24817);
nand UO_1026 (O_1026,N_24649,N_24390);
or UO_1027 (O_1027,N_24511,N_24618);
xnor UO_1028 (O_1028,N_24960,N_24744);
nand UO_1029 (O_1029,N_24825,N_24737);
nand UO_1030 (O_1030,N_24787,N_24951);
nor UO_1031 (O_1031,N_24631,N_24395);
and UO_1032 (O_1032,N_24769,N_24660);
and UO_1033 (O_1033,N_24825,N_24635);
xor UO_1034 (O_1034,N_24922,N_24713);
xnor UO_1035 (O_1035,N_24521,N_24433);
nand UO_1036 (O_1036,N_24578,N_24559);
and UO_1037 (O_1037,N_24792,N_24776);
and UO_1038 (O_1038,N_24898,N_24913);
and UO_1039 (O_1039,N_24608,N_24824);
nor UO_1040 (O_1040,N_24954,N_24900);
xor UO_1041 (O_1041,N_24643,N_24927);
nand UO_1042 (O_1042,N_24616,N_24710);
or UO_1043 (O_1043,N_24885,N_24985);
or UO_1044 (O_1044,N_24826,N_24785);
nor UO_1045 (O_1045,N_24509,N_24907);
nand UO_1046 (O_1046,N_24559,N_24737);
nor UO_1047 (O_1047,N_24631,N_24966);
xor UO_1048 (O_1048,N_24531,N_24417);
or UO_1049 (O_1049,N_24936,N_24931);
nand UO_1050 (O_1050,N_24614,N_24680);
and UO_1051 (O_1051,N_24792,N_24866);
or UO_1052 (O_1052,N_24741,N_24582);
xor UO_1053 (O_1053,N_24457,N_24574);
nor UO_1054 (O_1054,N_24867,N_24566);
and UO_1055 (O_1055,N_24847,N_24413);
xor UO_1056 (O_1056,N_24506,N_24952);
and UO_1057 (O_1057,N_24549,N_24809);
or UO_1058 (O_1058,N_24806,N_24689);
and UO_1059 (O_1059,N_24738,N_24787);
nand UO_1060 (O_1060,N_24684,N_24571);
and UO_1061 (O_1061,N_24491,N_24378);
nand UO_1062 (O_1062,N_24484,N_24719);
xor UO_1063 (O_1063,N_24765,N_24967);
xor UO_1064 (O_1064,N_24401,N_24928);
or UO_1065 (O_1065,N_24473,N_24610);
xnor UO_1066 (O_1066,N_24589,N_24598);
and UO_1067 (O_1067,N_24867,N_24805);
nor UO_1068 (O_1068,N_24722,N_24640);
or UO_1069 (O_1069,N_24809,N_24602);
and UO_1070 (O_1070,N_24655,N_24865);
and UO_1071 (O_1071,N_24729,N_24489);
or UO_1072 (O_1072,N_24860,N_24792);
or UO_1073 (O_1073,N_24711,N_24671);
nand UO_1074 (O_1074,N_24385,N_24611);
or UO_1075 (O_1075,N_24542,N_24602);
or UO_1076 (O_1076,N_24934,N_24493);
nor UO_1077 (O_1077,N_24554,N_24695);
or UO_1078 (O_1078,N_24502,N_24530);
or UO_1079 (O_1079,N_24833,N_24959);
nor UO_1080 (O_1080,N_24915,N_24834);
xnor UO_1081 (O_1081,N_24924,N_24383);
nor UO_1082 (O_1082,N_24618,N_24377);
nand UO_1083 (O_1083,N_24543,N_24992);
nand UO_1084 (O_1084,N_24604,N_24910);
or UO_1085 (O_1085,N_24846,N_24821);
and UO_1086 (O_1086,N_24524,N_24441);
and UO_1087 (O_1087,N_24926,N_24686);
xnor UO_1088 (O_1088,N_24963,N_24726);
nor UO_1089 (O_1089,N_24608,N_24694);
nor UO_1090 (O_1090,N_24664,N_24997);
nor UO_1091 (O_1091,N_24515,N_24797);
or UO_1092 (O_1092,N_24952,N_24994);
or UO_1093 (O_1093,N_24605,N_24840);
and UO_1094 (O_1094,N_24646,N_24541);
xnor UO_1095 (O_1095,N_24790,N_24724);
nor UO_1096 (O_1096,N_24885,N_24605);
and UO_1097 (O_1097,N_24804,N_24837);
xor UO_1098 (O_1098,N_24510,N_24966);
nand UO_1099 (O_1099,N_24668,N_24575);
nand UO_1100 (O_1100,N_24589,N_24398);
or UO_1101 (O_1101,N_24987,N_24567);
xnor UO_1102 (O_1102,N_24907,N_24595);
and UO_1103 (O_1103,N_24433,N_24840);
and UO_1104 (O_1104,N_24712,N_24512);
nand UO_1105 (O_1105,N_24689,N_24460);
or UO_1106 (O_1106,N_24611,N_24748);
xnor UO_1107 (O_1107,N_24965,N_24519);
or UO_1108 (O_1108,N_24615,N_24965);
or UO_1109 (O_1109,N_24508,N_24422);
or UO_1110 (O_1110,N_24559,N_24438);
or UO_1111 (O_1111,N_24389,N_24631);
and UO_1112 (O_1112,N_24478,N_24548);
and UO_1113 (O_1113,N_24782,N_24446);
or UO_1114 (O_1114,N_24557,N_24671);
nor UO_1115 (O_1115,N_24560,N_24397);
or UO_1116 (O_1116,N_24739,N_24443);
xnor UO_1117 (O_1117,N_24400,N_24765);
and UO_1118 (O_1118,N_24592,N_24788);
nand UO_1119 (O_1119,N_24663,N_24999);
or UO_1120 (O_1120,N_24541,N_24516);
xor UO_1121 (O_1121,N_24855,N_24444);
nor UO_1122 (O_1122,N_24403,N_24507);
and UO_1123 (O_1123,N_24396,N_24789);
nor UO_1124 (O_1124,N_24862,N_24451);
and UO_1125 (O_1125,N_24861,N_24876);
and UO_1126 (O_1126,N_24432,N_24781);
nor UO_1127 (O_1127,N_24729,N_24865);
xor UO_1128 (O_1128,N_24678,N_24927);
xor UO_1129 (O_1129,N_24461,N_24508);
nand UO_1130 (O_1130,N_24793,N_24483);
and UO_1131 (O_1131,N_24477,N_24774);
or UO_1132 (O_1132,N_24419,N_24859);
xnor UO_1133 (O_1133,N_24389,N_24994);
nor UO_1134 (O_1134,N_24974,N_24682);
or UO_1135 (O_1135,N_24582,N_24748);
xnor UO_1136 (O_1136,N_24565,N_24921);
nor UO_1137 (O_1137,N_24439,N_24532);
nor UO_1138 (O_1138,N_24644,N_24658);
nor UO_1139 (O_1139,N_24732,N_24910);
nand UO_1140 (O_1140,N_24590,N_24731);
or UO_1141 (O_1141,N_24435,N_24814);
and UO_1142 (O_1142,N_24640,N_24981);
nor UO_1143 (O_1143,N_24551,N_24547);
and UO_1144 (O_1144,N_24611,N_24718);
nor UO_1145 (O_1145,N_24447,N_24797);
xnor UO_1146 (O_1146,N_24505,N_24900);
nand UO_1147 (O_1147,N_24831,N_24732);
or UO_1148 (O_1148,N_24649,N_24555);
or UO_1149 (O_1149,N_24851,N_24644);
or UO_1150 (O_1150,N_24527,N_24518);
nand UO_1151 (O_1151,N_24872,N_24911);
nor UO_1152 (O_1152,N_24401,N_24575);
or UO_1153 (O_1153,N_24668,N_24614);
nand UO_1154 (O_1154,N_24512,N_24788);
nor UO_1155 (O_1155,N_24771,N_24652);
nand UO_1156 (O_1156,N_24536,N_24624);
and UO_1157 (O_1157,N_24445,N_24773);
or UO_1158 (O_1158,N_24437,N_24699);
xor UO_1159 (O_1159,N_24864,N_24740);
and UO_1160 (O_1160,N_24471,N_24533);
or UO_1161 (O_1161,N_24531,N_24703);
xnor UO_1162 (O_1162,N_24711,N_24408);
xnor UO_1163 (O_1163,N_24693,N_24403);
and UO_1164 (O_1164,N_24546,N_24822);
nor UO_1165 (O_1165,N_24912,N_24716);
or UO_1166 (O_1166,N_24859,N_24997);
xnor UO_1167 (O_1167,N_24759,N_24743);
nand UO_1168 (O_1168,N_24757,N_24733);
nor UO_1169 (O_1169,N_24424,N_24883);
nand UO_1170 (O_1170,N_24433,N_24437);
and UO_1171 (O_1171,N_24997,N_24643);
and UO_1172 (O_1172,N_24585,N_24598);
nand UO_1173 (O_1173,N_24450,N_24889);
nor UO_1174 (O_1174,N_24878,N_24913);
xor UO_1175 (O_1175,N_24525,N_24740);
nand UO_1176 (O_1176,N_24481,N_24750);
nand UO_1177 (O_1177,N_24542,N_24638);
xnor UO_1178 (O_1178,N_24586,N_24837);
nand UO_1179 (O_1179,N_24389,N_24906);
or UO_1180 (O_1180,N_24563,N_24777);
or UO_1181 (O_1181,N_24422,N_24968);
or UO_1182 (O_1182,N_24767,N_24418);
nor UO_1183 (O_1183,N_24908,N_24492);
or UO_1184 (O_1184,N_24964,N_24596);
nand UO_1185 (O_1185,N_24975,N_24448);
nand UO_1186 (O_1186,N_24599,N_24847);
and UO_1187 (O_1187,N_24726,N_24588);
xor UO_1188 (O_1188,N_24399,N_24808);
nand UO_1189 (O_1189,N_24830,N_24984);
nor UO_1190 (O_1190,N_24408,N_24851);
xor UO_1191 (O_1191,N_24789,N_24390);
nor UO_1192 (O_1192,N_24804,N_24698);
and UO_1193 (O_1193,N_24835,N_24885);
nand UO_1194 (O_1194,N_24656,N_24949);
nor UO_1195 (O_1195,N_24792,N_24802);
nand UO_1196 (O_1196,N_24377,N_24652);
xor UO_1197 (O_1197,N_24445,N_24538);
or UO_1198 (O_1198,N_24657,N_24930);
nand UO_1199 (O_1199,N_24909,N_24664);
nand UO_1200 (O_1200,N_24899,N_24411);
xnor UO_1201 (O_1201,N_24914,N_24451);
xor UO_1202 (O_1202,N_24793,N_24706);
nand UO_1203 (O_1203,N_24798,N_24593);
or UO_1204 (O_1204,N_24657,N_24492);
and UO_1205 (O_1205,N_24852,N_24574);
nor UO_1206 (O_1206,N_24810,N_24648);
or UO_1207 (O_1207,N_24931,N_24967);
xnor UO_1208 (O_1208,N_24656,N_24753);
nor UO_1209 (O_1209,N_24622,N_24896);
or UO_1210 (O_1210,N_24521,N_24966);
nand UO_1211 (O_1211,N_24428,N_24542);
xnor UO_1212 (O_1212,N_24744,N_24835);
xnor UO_1213 (O_1213,N_24961,N_24400);
nand UO_1214 (O_1214,N_24911,N_24982);
nor UO_1215 (O_1215,N_24625,N_24543);
and UO_1216 (O_1216,N_24687,N_24701);
nor UO_1217 (O_1217,N_24892,N_24444);
or UO_1218 (O_1218,N_24384,N_24949);
nand UO_1219 (O_1219,N_24863,N_24448);
nand UO_1220 (O_1220,N_24791,N_24758);
or UO_1221 (O_1221,N_24442,N_24600);
and UO_1222 (O_1222,N_24378,N_24950);
xor UO_1223 (O_1223,N_24627,N_24972);
nand UO_1224 (O_1224,N_24469,N_24705);
and UO_1225 (O_1225,N_24514,N_24473);
nor UO_1226 (O_1226,N_24592,N_24664);
nor UO_1227 (O_1227,N_24971,N_24515);
or UO_1228 (O_1228,N_24987,N_24931);
xor UO_1229 (O_1229,N_24991,N_24858);
xnor UO_1230 (O_1230,N_24836,N_24783);
nor UO_1231 (O_1231,N_24643,N_24476);
or UO_1232 (O_1232,N_24765,N_24444);
and UO_1233 (O_1233,N_24953,N_24424);
nor UO_1234 (O_1234,N_24609,N_24597);
nor UO_1235 (O_1235,N_24850,N_24932);
or UO_1236 (O_1236,N_24628,N_24947);
or UO_1237 (O_1237,N_24522,N_24626);
nand UO_1238 (O_1238,N_24966,N_24532);
or UO_1239 (O_1239,N_24941,N_24748);
xor UO_1240 (O_1240,N_24862,N_24465);
xnor UO_1241 (O_1241,N_24591,N_24640);
nand UO_1242 (O_1242,N_24947,N_24983);
nor UO_1243 (O_1243,N_24650,N_24990);
nand UO_1244 (O_1244,N_24894,N_24776);
or UO_1245 (O_1245,N_24660,N_24768);
and UO_1246 (O_1246,N_24826,N_24725);
or UO_1247 (O_1247,N_24902,N_24813);
xnor UO_1248 (O_1248,N_24979,N_24835);
or UO_1249 (O_1249,N_24786,N_24413);
or UO_1250 (O_1250,N_24718,N_24408);
or UO_1251 (O_1251,N_24564,N_24708);
nor UO_1252 (O_1252,N_24966,N_24731);
nand UO_1253 (O_1253,N_24984,N_24877);
nor UO_1254 (O_1254,N_24795,N_24547);
or UO_1255 (O_1255,N_24406,N_24646);
nand UO_1256 (O_1256,N_24937,N_24494);
xnor UO_1257 (O_1257,N_24393,N_24597);
xnor UO_1258 (O_1258,N_24944,N_24778);
xor UO_1259 (O_1259,N_24863,N_24734);
and UO_1260 (O_1260,N_24749,N_24527);
or UO_1261 (O_1261,N_24913,N_24974);
nor UO_1262 (O_1262,N_24411,N_24754);
and UO_1263 (O_1263,N_24877,N_24610);
nand UO_1264 (O_1264,N_24465,N_24640);
nor UO_1265 (O_1265,N_24431,N_24596);
nor UO_1266 (O_1266,N_24634,N_24413);
xnor UO_1267 (O_1267,N_24733,N_24611);
and UO_1268 (O_1268,N_24864,N_24660);
xnor UO_1269 (O_1269,N_24983,N_24879);
or UO_1270 (O_1270,N_24895,N_24610);
nor UO_1271 (O_1271,N_24592,N_24873);
and UO_1272 (O_1272,N_24665,N_24623);
nand UO_1273 (O_1273,N_24552,N_24512);
or UO_1274 (O_1274,N_24599,N_24890);
and UO_1275 (O_1275,N_24629,N_24687);
nor UO_1276 (O_1276,N_24948,N_24500);
or UO_1277 (O_1277,N_24467,N_24883);
nor UO_1278 (O_1278,N_24716,N_24606);
or UO_1279 (O_1279,N_24567,N_24902);
nor UO_1280 (O_1280,N_24738,N_24993);
and UO_1281 (O_1281,N_24509,N_24673);
or UO_1282 (O_1282,N_24914,N_24771);
nand UO_1283 (O_1283,N_24397,N_24948);
nor UO_1284 (O_1284,N_24671,N_24649);
nor UO_1285 (O_1285,N_24553,N_24980);
and UO_1286 (O_1286,N_24876,N_24992);
nor UO_1287 (O_1287,N_24582,N_24733);
xor UO_1288 (O_1288,N_24760,N_24877);
nand UO_1289 (O_1289,N_24412,N_24936);
nor UO_1290 (O_1290,N_24759,N_24538);
nor UO_1291 (O_1291,N_24716,N_24413);
nor UO_1292 (O_1292,N_24378,N_24636);
nor UO_1293 (O_1293,N_24953,N_24735);
and UO_1294 (O_1294,N_24436,N_24564);
and UO_1295 (O_1295,N_24725,N_24620);
or UO_1296 (O_1296,N_24610,N_24772);
nor UO_1297 (O_1297,N_24691,N_24593);
nor UO_1298 (O_1298,N_24920,N_24778);
xor UO_1299 (O_1299,N_24595,N_24619);
or UO_1300 (O_1300,N_24710,N_24859);
xnor UO_1301 (O_1301,N_24993,N_24438);
and UO_1302 (O_1302,N_24939,N_24477);
or UO_1303 (O_1303,N_24552,N_24678);
xor UO_1304 (O_1304,N_24714,N_24848);
xor UO_1305 (O_1305,N_24465,N_24389);
nand UO_1306 (O_1306,N_24871,N_24683);
and UO_1307 (O_1307,N_24466,N_24756);
and UO_1308 (O_1308,N_24592,N_24998);
and UO_1309 (O_1309,N_24490,N_24675);
nand UO_1310 (O_1310,N_24682,N_24483);
xnor UO_1311 (O_1311,N_24508,N_24694);
or UO_1312 (O_1312,N_24678,N_24890);
nor UO_1313 (O_1313,N_24529,N_24911);
nand UO_1314 (O_1314,N_24946,N_24666);
nand UO_1315 (O_1315,N_24877,N_24423);
nand UO_1316 (O_1316,N_24440,N_24761);
nor UO_1317 (O_1317,N_24594,N_24463);
and UO_1318 (O_1318,N_24515,N_24785);
nor UO_1319 (O_1319,N_24378,N_24882);
and UO_1320 (O_1320,N_24617,N_24686);
nor UO_1321 (O_1321,N_24671,N_24706);
nand UO_1322 (O_1322,N_24957,N_24462);
xor UO_1323 (O_1323,N_24658,N_24465);
and UO_1324 (O_1324,N_24478,N_24805);
and UO_1325 (O_1325,N_24461,N_24802);
nand UO_1326 (O_1326,N_24705,N_24850);
or UO_1327 (O_1327,N_24634,N_24417);
nand UO_1328 (O_1328,N_24481,N_24671);
xnor UO_1329 (O_1329,N_24522,N_24766);
nand UO_1330 (O_1330,N_24870,N_24528);
nand UO_1331 (O_1331,N_24579,N_24566);
or UO_1332 (O_1332,N_24815,N_24693);
or UO_1333 (O_1333,N_24970,N_24626);
xnor UO_1334 (O_1334,N_24918,N_24410);
xor UO_1335 (O_1335,N_24906,N_24940);
xnor UO_1336 (O_1336,N_24627,N_24793);
and UO_1337 (O_1337,N_24822,N_24678);
nand UO_1338 (O_1338,N_24838,N_24903);
xnor UO_1339 (O_1339,N_24571,N_24594);
or UO_1340 (O_1340,N_24414,N_24597);
nor UO_1341 (O_1341,N_24961,N_24602);
nor UO_1342 (O_1342,N_24961,N_24685);
and UO_1343 (O_1343,N_24590,N_24591);
and UO_1344 (O_1344,N_24422,N_24471);
or UO_1345 (O_1345,N_24732,N_24542);
nor UO_1346 (O_1346,N_24665,N_24413);
nor UO_1347 (O_1347,N_24957,N_24949);
or UO_1348 (O_1348,N_24508,N_24452);
or UO_1349 (O_1349,N_24991,N_24906);
xnor UO_1350 (O_1350,N_24588,N_24500);
nor UO_1351 (O_1351,N_24741,N_24589);
xor UO_1352 (O_1352,N_24455,N_24609);
nand UO_1353 (O_1353,N_24722,N_24913);
nand UO_1354 (O_1354,N_24776,N_24636);
or UO_1355 (O_1355,N_24579,N_24398);
or UO_1356 (O_1356,N_24750,N_24624);
nor UO_1357 (O_1357,N_24870,N_24557);
or UO_1358 (O_1358,N_24648,N_24464);
or UO_1359 (O_1359,N_24514,N_24501);
nand UO_1360 (O_1360,N_24720,N_24563);
nor UO_1361 (O_1361,N_24997,N_24574);
and UO_1362 (O_1362,N_24890,N_24570);
and UO_1363 (O_1363,N_24545,N_24563);
and UO_1364 (O_1364,N_24858,N_24825);
nand UO_1365 (O_1365,N_24544,N_24513);
nor UO_1366 (O_1366,N_24515,N_24408);
nand UO_1367 (O_1367,N_24866,N_24649);
and UO_1368 (O_1368,N_24769,N_24832);
nand UO_1369 (O_1369,N_24984,N_24383);
nand UO_1370 (O_1370,N_24641,N_24915);
nor UO_1371 (O_1371,N_24576,N_24482);
and UO_1372 (O_1372,N_24689,N_24908);
xor UO_1373 (O_1373,N_24981,N_24453);
xnor UO_1374 (O_1374,N_24468,N_24980);
and UO_1375 (O_1375,N_24483,N_24447);
nor UO_1376 (O_1376,N_24630,N_24611);
or UO_1377 (O_1377,N_24405,N_24813);
nand UO_1378 (O_1378,N_24696,N_24711);
xnor UO_1379 (O_1379,N_24909,N_24783);
nand UO_1380 (O_1380,N_24634,N_24875);
xnor UO_1381 (O_1381,N_24699,N_24930);
xnor UO_1382 (O_1382,N_24673,N_24892);
xnor UO_1383 (O_1383,N_24844,N_24554);
or UO_1384 (O_1384,N_24959,N_24779);
and UO_1385 (O_1385,N_24433,N_24383);
nand UO_1386 (O_1386,N_24624,N_24375);
or UO_1387 (O_1387,N_24607,N_24899);
or UO_1388 (O_1388,N_24772,N_24568);
nor UO_1389 (O_1389,N_24783,N_24602);
and UO_1390 (O_1390,N_24813,N_24953);
xnor UO_1391 (O_1391,N_24532,N_24763);
xor UO_1392 (O_1392,N_24766,N_24876);
nor UO_1393 (O_1393,N_24850,N_24914);
nor UO_1394 (O_1394,N_24472,N_24460);
nor UO_1395 (O_1395,N_24913,N_24846);
nor UO_1396 (O_1396,N_24865,N_24810);
xor UO_1397 (O_1397,N_24519,N_24617);
nor UO_1398 (O_1398,N_24448,N_24824);
and UO_1399 (O_1399,N_24460,N_24912);
nand UO_1400 (O_1400,N_24865,N_24590);
nor UO_1401 (O_1401,N_24933,N_24820);
nand UO_1402 (O_1402,N_24977,N_24991);
xnor UO_1403 (O_1403,N_24451,N_24551);
or UO_1404 (O_1404,N_24476,N_24424);
and UO_1405 (O_1405,N_24883,N_24890);
and UO_1406 (O_1406,N_24825,N_24683);
or UO_1407 (O_1407,N_24570,N_24661);
nand UO_1408 (O_1408,N_24951,N_24591);
or UO_1409 (O_1409,N_24790,N_24533);
and UO_1410 (O_1410,N_24523,N_24733);
nand UO_1411 (O_1411,N_24634,N_24454);
xor UO_1412 (O_1412,N_24459,N_24947);
and UO_1413 (O_1413,N_24586,N_24708);
nand UO_1414 (O_1414,N_24784,N_24443);
nor UO_1415 (O_1415,N_24714,N_24436);
and UO_1416 (O_1416,N_24442,N_24806);
or UO_1417 (O_1417,N_24740,N_24840);
xor UO_1418 (O_1418,N_24976,N_24601);
or UO_1419 (O_1419,N_24531,N_24619);
and UO_1420 (O_1420,N_24399,N_24707);
nor UO_1421 (O_1421,N_24591,N_24537);
nand UO_1422 (O_1422,N_24874,N_24469);
or UO_1423 (O_1423,N_24462,N_24688);
and UO_1424 (O_1424,N_24942,N_24999);
or UO_1425 (O_1425,N_24882,N_24955);
xnor UO_1426 (O_1426,N_24512,N_24991);
and UO_1427 (O_1427,N_24968,N_24426);
nand UO_1428 (O_1428,N_24824,N_24578);
nor UO_1429 (O_1429,N_24729,N_24998);
nand UO_1430 (O_1430,N_24680,N_24873);
xor UO_1431 (O_1431,N_24402,N_24733);
nand UO_1432 (O_1432,N_24528,N_24846);
nor UO_1433 (O_1433,N_24980,N_24688);
xnor UO_1434 (O_1434,N_24620,N_24901);
nand UO_1435 (O_1435,N_24711,N_24959);
nor UO_1436 (O_1436,N_24950,N_24648);
and UO_1437 (O_1437,N_24678,N_24602);
xor UO_1438 (O_1438,N_24696,N_24447);
nand UO_1439 (O_1439,N_24729,N_24767);
nor UO_1440 (O_1440,N_24502,N_24949);
nand UO_1441 (O_1441,N_24428,N_24895);
nor UO_1442 (O_1442,N_24921,N_24939);
nand UO_1443 (O_1443,N_24730,N_24899);
nand UO_1444 (O_1444,N_24532,N_24955);
and UO_1445 (O_1445,N_24386,N_24927);
nand UO_1446 (O_1446,N_24649,N_24690);
nand UO_1447 (O_1447,N_24727,N_24888);
nand UO_1448 (O_1448,N_24763,N_24655);
xnor UO_1449 (O_1449,N_24779,N_24468);
or UO_1450 (O_1450,N_24523,N_24928);
nand UO_1451 (O_1451,N_24476,N_24941);
or UO_1452 (O_1452,N_24792,N_24442);
nor UO_1453 (O_1453,N_24999,N_24715);
and UO_1454 (O_1454,N_24690,N_24755);
nor UO_1455 (O_1455,N_24832,N_24828);
nand UO_1456 (O_1456,N_24759,N_24807);
nand UO_1457 (O_1457,N_24925,N_24818);
nor UO_1458 (O_1458,N_24907,N_24979);
nand UO_1459 (O_1459,N_24817,N_24978);
xor UO_1460 (O_1460,N_24837,N_24819);
and UO_1461 (O_1461,N_24461,N_24677);
xor UO_1462 (O_1462,N_24758,N_24506);
nor UO_1463 (O_1463,N_24824,N_24678);
xor UO_1464 (O_1464,N_24829,N_24449);
nor UO_1465 (O_1465,N_24910,N_24873);
xnor UO_1466 (O_1466,N_24419,N_24558);
nand UO_1467 (O_1467,N_24599,N_24466);
xnor UO_1468 (O_1468,N_24494,N_24953);
nand UO_1469 (O_1469,N_24677,N_24793);
xor UO_1470 (O_1470,N_24440,N_24525);
xor UO_1471 (O_1471,N_24744,N_24925);
nor UO_1472 (O_1472,N_24973,N_24767);
or UO_1473 (O_1473,N_24959,N_24412);
nand UO_1474 (O_1474,N_24530,N_24518);
nor UO_1475 (O_1475,N_24939,N_24967);
or UO_1476 (O_1476,N_24474,N_24901);
or UO_1477 (O_1477,N_24899,N_24468);
or UO_1478 (O_1478,N_24827,N_24731);
or UO_1479 (O_1479,N_24488,N_24379);
and UO_1480 (O_1480,N_24916,N_24950);
nor UO_1481 (O_1481,N_24798,N_24636);
and UO_1482 (O_1482,N_24733,N_24501);
nand UO_1483 (O_1483,N_24881,N_24983);
nand UO_1484 (O_1484,N_24533,N_24865);
xnor UO_1485 (O_1485,N_24669,N_24937);
or UO_1486 (O_1486,N_24502,N_24827);
nor UO_1487 (O_1487,N_24495,N_24497);
or UO_1488 (O_1488,N_24480,N_24551);
nor UO_1489 (O_1489,N_24880,N_24646);
nand UO_1490 (O_1490,N_24767,N_24903);
nand UO_1491 (O_1491,N_24828,N_24847);
xnor UO_1492 (O_1492,N_24632,N_24844);
and UO_1493 (O_1493,N_24821,N_24963);
nand UO_1494 (O_1494,N_24635,N_24586);
and UO_1495 (O_1495,N_24674,N_24527);
nand UO_1496 (O_1496,N_24567,N_24971);
xnor UO_1497 (O_1497,N_24884,N_24894);
nor UO_1498 (O_1498,N_24416,N_24465);
or UO_1499 (O_1499,N_24504,N_24899);
or UO_1500 (O_1500,N_24796,N_24661);
xnor UO_1501 (O_1501,N_24838,N_24872);
xnor UO_1502 (O_1502,N_24593,N_24563);
or UO_1503 (O_1503,N_24599,N_24462);
xnor UO_1504 (O_1504,N_24521,N_24942);
xnor UO_1505 (O_1505,N_24961,N_24485);
nand UO_1506 (O_1506,N_24616,N_24494);
nor UO_1507 (O_1507,N_24514,N_24524);
xor UO_1508 (O_1508,N_24730,N_24927);
nor UO_1509 (O_1509,N_24834,N_24380);
nor UO_1510 (O_1510,N_24427,N_24968);
and UO_1511 (O_1511,N_24534,N_24767);
xnor UO_1512 (O_1512,N_24824,N_24682);
and UO_1513 (O_1513,N_24774,N_24563);
nand UO_1514 (O_1514,N_24575,N_24618);
or UO_1515 (O_1515,N_24715,N_24630);
nor UO_1516 (O_1516,N_24878,N_24790);
nand UO_1517 (O_1517,N_24386,N_24614);
and UO_1518 (O_1518,N_24936,N_24614);
or UO_1519 (O_1519,N_24640,N_24841);
nor UO_1520 (O_1520,N_24649,N_24824);
and UO_1521 (O_1521,N_24782,N_24523);
nand UO_1522 (O_1522,N_24407,N_24845);
or UO_1523 (O_1523,N_24986,N_24747);
nand UO_1524 (O_1524,N_24944,N_24684);
xnor UO_1525 (O_1525,N_24950,N_24613);
xor UO_1526 (O_1526,N_24924,N_24861);
and UO_1527 (O_1527,N_24737,N_24891);
xor UO_1528 (O_1528,N_24579,N_24641);
nor UO_1529 (O_1529,N_24476,N_24467);
and UO_1530 (O_1530,N_24671,N_24625);
and UO_1531 (O_1531,N_24963,N_24571);
nor UO_1532 (O_1532,N_24431,N_24817);
nor UO_1533 (O_1533,N_24643,N_24435);
or UO_1534 (O_1534,N_24705,N_24962);
nor UO_1535 (O_1535,N_24741,N_24573);
or UO_1536 (O_1536,N_24694,N_24848);
or UO_1537 (O_1537,N_24653,N_24841);
xnor UO_1538 (O_1538,N_24942,N_24489);
nand UO_1539 (O_1539,N_24945,N_24658);
or UO_1540 (O_1540,N_24915,N_24817);
and UO_1541 (O_1541,N_24470,N_24918);
and UO_1542 (O_1542,N_24895,N_24739);
or UO_1543 (O_1543,N_24859,N_24595);
or UO_1544 (O_1544,N_24593,N_24666);
or UO_1545 (O_1545,N_24543,N_24672);
and UO_1546 (O_1546,N_24448,N_24475);
and UO_1547 (O_1547,N_24917,N_24723);
or UO_1548 (O_1548,N_24908,N_24835);
or UO_1549 (O_1549,N_24814,N_24884);
nor UO_1550 (O_1550,N_24599,N_24398);
and UO_1551 (O_1551,N_24681,N_24398);
nand UO_1552 (O_1552,N_24862,N_24942);
or UO_1553 (O_1553,N_24655,N_24629);
or UO_1554 (O_1554,N_24992,N_24430);
nand UO_1555 (O_1555,N_24807,N_24836);
xor UO_1556 (O_1556,N_24901,N_24615);
xnor UO_1557 (O_1557,N_24635,N_24704);
and UO_1558 (O_1558,N_24506,N_24470);
nor UO_1559 (O_1559,N_24719,N_24898);
nor UO_1560 (O_1560,N_24432,N_24897);
or UO_1561 (O_1561,N_24712,N_24444);
nand UO_1562 (O_1562,N_24862,N_24601);
nand UO_1563 (O_1563,N_24624,N_24673);
and UO_1564 (O_1564,N_24623,N_24884);
xor UO_1565 (O_1565,N_24447,N_24556);
nand UO_1566 (O_1566,N_24864,N_24623);
xor UO_1567 (O_1567,N_24753,N_24807);
nor UO_1568 (O_1568,N_24825,N_24781);
nor UO_1569 (O_1569,N_24862,N_24595);
nand UO_1570 (O_1570,N_24850,N_24936);
and UO_1571 (O_1571,N_24792,N_24530);
nand UO_1572 (O_1572,N_24648,N_24949);
nor UO_1573 (O_1573,N_24588,N_24747);
nor UO_1574 (O_1574,N_24398,N_24610);
or UO_1575 (O_1575,N_24872,N_24409);
nor UO_1576 (O_1576,N_24635,N_24775);
nor UO_1577 (O_1577,N_24890,N_24761);
or UO_1578 (O_1578,N_24609,N_24702);
nand UO_1579 (O_1579,N_24877,N_24987);
nand UO_1580 (O_1580,N_24527,N_24845);
xnor UO_1581 (O_1581,N_24976,N_24416);
and UO_1582 (O_1582,N_24818,N_24452);
or UO_1583 (O_1583,N_24562,N_24561);
nand UO_1584 (O_1584,N_24947,N_24854);
or UO_1585 (O_1585,N_24841,N_24681);
nor UO_1586 (O_1586,N_24526,N_24655);
xor UO_1587 (O_1587,N_24517,N_24524);
and UO_1588 (O_1588,N_24509,N_24405);
and UO_1589 (O_1589,N_24593,N_24776);
and UO_1590 (O_1590,N_24809,N_24556);
and UO_1591 (O_1591,N_24695,N_24947);
or UO_1592 (O_1592,N_24920,N_24934);
nand UO_1593 (O_1593,N_24935,N_24494);
nand UO_1594 (O_1594,N_24964,N_24983);
and UO_1595 (O_1595,N_24635,N_24949);
nand UO_1596 (O_1596,N_24641,N_24764);
and UO_1597 (O_1597,N_24429,N_24533);
nand UO_1598 (O_1598,N_24517,N_24839);
nand UO_1599 (O_1599,N_24555,N_24393);
nor UO_1600 (O_1600,N_24429,N_24811);
and UO_1601 (O_1601,N_24635,N_24539);
and UO_1602 (O_1602,N_24936,N_24668);
nor UO_1603 (O_1603,N_24626,N_24586);
nor UO_1604 (O_1604,N_24689,N_24445);
or UO_1605 (O_1605,N_24676,N_24534);
and UO_1606 (O_1606,N_24445,N_24904);
nand UO_1607 (O_1607,N_24726,N_24840);
nand UO_1608 (O_1608,N_24698,N_24734);
and UO_1609 (O_1609,N_24647,N_24765);
nor UO_1610 (O_1610,N_24815,N_24468);
xnor UO_1611 (O_1611,N_24448,N_24704);
xor UO_1612 (O_1612,N_24814,N_24541);
or UO_1613 (O_1613,N_24427,N_24792);
or UO_1614 (O_1614,N_24450,N_24532);
nor UO_1615 (O_1615,N_24766,N_24516);
nor UO_1616 (O_1616,N_24708,N_24544);
and UO_1617 (O_1617,N_24692,N_24869);
nor UO_1618 (O_1618,N_24601,N_24464);
nand UO_1619 (O_1619,N_24835,N_24616);
nor UO_1620 (O_1620,N_24659,N_24450);
and UO_1621 (O_1621,N_24587,N_24718);
or UO_1622 (O_1622,N_24406,N_24505);
nor UO_1623 (O_1623,N_24526,N_24424);
or UO_1624 (O_1624,N_24511,N_24609);
xor UO_1625 (O_1625,N_24969,N_24688);
xor UO_1626 (O_1626,N_24689,N_24511);
nand UO_1627 (O_1627,N_24901,N_24859);
and UO_1628 (O_1628,N_24772,N_24866);
and UO_1629 (O_1629,N_24440,N_24633);
nand UO_1630 (O_1630,N_24586,N_24662);
nor UO_1631 (O_1631,N_24408,N_24877);
xnor UO_1632 (O_1632,N_24422,N_24708);
xor UO_1633 (O_1633,N_24989,N_24573);
nand UO_1634 (O_1634,N_24861,N_24567);
nand UO_1635 (O_1635,N_24657,N_24840);
nor UO_1636 (O_1636,N_24488,N_24962);
and UO_1637 (O_1637,N_24909,N_24440);
nor UO_1638 (O_1638,N_24410,N_24934);
nand UO_1639 (O_1639,N_24397,N_24799);
or UO_1640 (O_1640,N_24519,N_24574);
or UO_1641 (O_1641,N_24855,N_24721);
xnor UO_1642 (O_1642,N_24894,N_24845);
nand UO_1643 (O_1643,N_24761,N_24475);
nor UO_1644 (O_1644,N_24836,N_24739);
xnor UO_1645 (O_1645,N_24673,N_24550);
nand UO_1646 (O_1646,N_24602,N_24853);
xnor UO_1647 (O_1647,N_24933,N_24604);
and UO_1648 (O_1648,N_24926,N_24525);
nor UO_1649 (O_1649,N_24565,N_24484);
xor UO_1650 (O_1650,N_24978,N_24919);
and UO_1651 (O_1651,N_24847,N_24730);
xor UO_1652 (O_1652,N_24708,N_24965);
or UO_1653 (O_1653,N_24475,N_24845);
and UO_1654 (O_1654,N_24543,N_24706);
nand UO_1655 (O_1655,N_24623,N_24702);
nand UO_1656 (O_1656,N_24550,N_24780);
xnor UO_1657 (O_1657,N_24741,N_24977);
and UO_1658 (O_1658,N_24792,N_24745);
or UO_1659 (O_1659,N_24649,N_24522);
nand UO_1660 (O_1660,N_24426,N_24388);
nand UO_1661 (O_1661,N_24605,N_24896);
nand UO_1662 (O_1662,N_24827,N_24745);
and UO_1663 (O_1663,N_24832,N_24847);
nor UO_1664 (O_1664,N_24986,N_24819);
or UO_1665 (O_1665,N_24515,N_24954);
nand UO_1666 (O_1666,N_24871,N_24894);
and UO_1667 (O_1667,N_24842,N_24515);
nand UO_1668 (O_1668,N_24993,N_24844);
and UO_1669 (O_1669,N_24421,N_24687);
and UO_1670 (O_1670,N_24690,N_24997);
xor UO_1671 (O_1671,N_24476,N_24388);
nor UO_1672 (O_1672,N_24731,N_24612);
nand UO_1673 (O_1673,N_24513,N_24656);
or UO_1674 (O_1674,N_24700,N_24432);
or UO_1675 (O_1675,N_24754,N_24848);
nand UO_1676 (O_1676,N_24690,N_24498);
and UO_1677 (O_1677,N_24907,N_24692);
or UO_1678 (O_1678,N_24771,N_24926);
xor UO_1679 (O_1679,N_24521,N_24837);
or UO_1680 (O_1680,N_24895,N_24983);
or UO_1681 (O_1681,N_24655,N_24942);
and UO_1682 (O_1682,N_24833,N_24770);
nor UO_1683 (O_1683,N_24564,N_24667);
or UO_1684 (O_1684,N_24692,N_24906);
or UO_1685 (O_1685,N_24869,N_24596);
nand UO_1686 (O_1686,N_24392,N_24942);
nor UO_1687 (O_1687,N_24419,N_24908);
and UO_1688 (O_1688,N_24845,N_24965);
and UO_1689 (O_1689,N_24681,N_24396);
or UO_1690 (O_1690,N_24444,N_24774);
and UO_1691 (O_1691,N_24899,N_24911);
and UO_1692 (O_1692,N_24444,N_24777);
nand UO_1693 (O_1693,N_24881,N_24533);
nor UO_1694 (O_1694,N_24403,N_24572);
xor UO_1695 (O_1695,N_24854,N_24684);
or UO_1696 (O_1696,N_24642,N_24822);
xor UO_1697 (O_1697,N_24575,N_24943);
or UO_1698 (O_1698,N_24750,N_24829);
nand UO_1699 (O_1699,N_24766,N_24378);
or UO_1700 (O_1700,N_24547,N_24922);
xor UO_1701 (O_1701,N_24957,N_24398);
nand UO_1702 (O_1702,N_24620,N_24630);
xnor UO_1703 (O_1703,N_24620,N_24908);
xnor UO_1704 (O_1704,N_24449,N_24872);
or UO_1705 (O_1705,N_24806,N_24910);
or UO_1706 (O_1706,N_24904,N_24751);
nor UO_1707 (O_1707,N_24961,N_24586);
nor UO_1708 (O_1708,N_24639,N_24411);
nand UO_1709 (O_1709,N_24605,N_24888);
nor UO_1710 (O_1710,N_24815,N_24983);
nand UO_1711 (O_1711,N_24825,N_24959);
xor UO_1712 (O_1712,N_24753,N_24490);
nor UO_1713 (O_1713,N_24530,N_24919);
nor UO_1714 (O_1714,N_24594,N_24443);
xnor UO_1715 (O_1715,N_24686,N_24595);
xnor UO_1716 (O_1716,N_24623,N_24465);
nor UO_1717 (O_1717,N_24529,N_24553);
xnor UO_1718 (O_1718,N_24560,N_24516);
or UO_1719 (O_1719,N_24426,N_24907);
nand UO_1720 (O_1720,N_24977,N_24928);
nor UO_1721 (O_1721,N_24917,N_24788);
nor UO_1722 (O_1722,N_24600,N_24812);
or UO_1723 (O_1723,N_24669,N_24576);
and UO_1724 (O_1724,N_24574,N_24794);
nand UO_1725 (O_1725,N_24671,N_24578);
nand UO_1726 (O_1726,N_24630,N_24997);
and UO_1727 (O_1727,N_24905,N_24999);
xor UO_1728 (O_1728,N_24548,N_24388);
nor UO_1729 (O_1729,N_24800,N_24926);
nor UO_1730 (O_1730,N_24855,N_24445);
nand UO_1731 (O_1731,N_24629,N_24679);
and UO_1732 (O_1732,N_24592,N_24539);
and UO_1733 (O_1733,N_24968,N_24424);
nand UO_1734 (O_1734,N_24409,N_24910);
nor UO_1735 (O_1735,N_24426,N_24465);
nand UO_1736 (O_1736,N_24509,N_24376);
xnor UO_1737 (O_1737,N_24395,N_24382);
and UO_1738 (O_1738,N_24700,N_24713);
xor UO_1739 (O_1739,N_24587,N_24980);
nor UO_1740 (O_1740,N_24566,N_24604);
and UO_1741 (O_1741,N_24585,N_24469);
nor UO_1742 (O_1742,N_24485,N_24522);
xor UO_1743 (O_1743,N_24486,N_24858);
xor UO_1744 (O_1744,N_24437,N_24822);
xnor UO_1745 (O_1745,N_24726,N_24692);
or UO_1746 (O_1746,N_24565,N_24586);
xor UO_1747 (O_1747,N_24638,N_24575);
or UO_1748 (O_1748,N_24599,N_24516);
nand UO_1749 (O_1749,N_24629,N_24993);
nand UO_1750 (O_1750,N_24477,N_24663);
nand UO_1751 (O_1751,N_24876,N_24487);
nand UO_1752 (O_1752,N_24462,N_24403);
nand UO_1753 (O_1753,N_24748,N_24871);
nand UO_1754 (O_1754,N_24599,N_24685);
nor UO_1755 (O_1755,N_24866,N_24441);
xor UO_1756 (O_1756,N_24861,N_24566);
nor UO_1757 (O_1757,N_24618,N_24576);
or UO_1758 (O_1758,N_24861,N_24824);
nor UO_1759 (O_1759,N_24460,N_24520);
or UO_1760 (O_1760,N_24686,N_24796);
and UO_1761 (O_1761,N_24756,N_24921);
nand UO_1762 (O_1762,N_24820,N_24939);
or UO_1763 (O_1763,N_24625,N_24880);
and UO_1764 (O_1764,N_24488,N_24413);
nor UO_1765 (O_1765,N_24695,N_24412);
nand UO_1766 (O_1766,N_24581,N_24801);
or UO_1767 (O_1767,N_24883,N_24457);
nor UO_1768 (O_1768,N_24947,N_24556);
xnor UO_1769 (O_1769,N_24595,N_24710);
or UO_1770 (O_1770,N_24434,N_24744);
xor UO_1771 (O_1771,N_24496,N_24822);
nor UO_1772 (O_1772,N_24846,N_24958);
nor UO_1773 (O_1773,N_24912,N_24562);
xnor UO_1774 (O_1774,N_24475,N_24417);
xnor UO_1775 (O_1775,N_24512,N_24521);
nand UO_1776 (O_1776,N_24469,N_24965);
xnor UO_1777 (O_1777,N_24725,N_24809);
and UO_1778 (O_1778,N_24729,N_24827);
nor UO_1779 (O_1779,N_24995,N_24890);
xnor UO_1780 (O_1780,N_24995,N_24610);
nand UO_1781 (O_1781,N_24654,N_24788);
xor UO_1782 (O_1782,N_24684,N_24526);
and UO_1783 (O_1783,N_24420,N_24933);
nand UO_1784 (O_1784,N_24460,N_24963);
and UO_1785 (O_1785,N_24935,N_24824);
xor UO_1786 (O_1786,N_24982,N_24747);
nand UO_1787 (O_1787,N_24477,N_24929);
nand UO_1788 (O_1788,N_24448,N_24962);
and UO_1789 (O_1789,N_24800,N_24509);
xor UO_1790 (O_1790,N_24710,N_24899);
xnor UO_1791 (O_1791,N_24792,N_24379);
nand UO_1792 (O_1792,N_24796,N_24837);
nor UO_1793 (O_1793,N_24547,N_24515);
or UO_1794 (O_1794,N_24939,N_24781);
nor UO_1795 (O_1795,N_24884,N_24980);
or UO_1796 (O_1796,N_24806,N_24583);
xor UO_1797 (O_1797,N_24388,N_24498);
and UO_1798 (O_1798,N_24422,N_24881);
and UO_1799 (O_1799,N_24685,N_24615);
or UO_1800 (O_1800,N_24567,N_24782);
nor UO_1801 (O_1801,N_24973,N_24648);
nand UO_1802 (O_1802,N_24627,N_24500);
and UO_1803 (O_1803,N_24821,N_24399);
nor UO_1804 (O_1804,N_24868,N_24957);
or UO_1805 (O_1805,N_24861,N_24544);
xor UO_1806 (O_1806,N_24685,N_24643);
and UO_1807 (O_1807,N_24556,N_24893);
xnor UO_1808 (O_1808,N_24496,N_24678);
xnor UO_1809 (O_1809,N_24632,N_24889);
nand UO_1810 (O_1810,N_24440,N_24865);
xor UO_1811 (O_1811,N_24517,N_24762);
nor UO_1812 (O_1812,N_24878,N_24398);
xor UO_1813 (O_1813,N_24684,N_24742);
nor UO_1814 (O_1814,N_24866,N_24588);
nor UO_1815 (O_1815,N_24712,N_24525);
nand UO_1816 (O_1816,N_24469,N_24402);
or UO_1817 (O_1817,N_24672,N_24376);
nand UO_1818 (O_1818,N_24450,N_24580);
xnor UO_1819 (O_1819,N_24868,N_24507);
nor UO_1820 (O_1820,N_24633,N_24460);
and UO_1821 (O_1821,N_24954,N_24445);
nand UO_1822 (O_1822,N_24797,N_24873);
or UO_1823 (O_1823,N_24605,N_24587);
nor UO_1824 (O_1824,N_24494,N_24698);
xnor UO_1825 (O_1825,N_24999,N_24487);
nand UO_1826 (O_1826,N_24840,N_24382);
or UO_1827 (O_1827,N_24761,N_24740);
xor UO_1828 (O_1828,N_24739,N_24375);
nor UO_1829 (O_1829,N_24925,N_24815);
or UO_1830 (O_1830,N_24963,N_24526);
nand UO_1831 (O_1831,N_24675,N_24627);
nor UO_1832 (O_1832,N_24798,N_24905);
xor UO_1833 (O_1833,N_24948,N_24648);
nor UO_1834 (O_1834,N_24512,N_24902);
nand UO_1835 (O_1835,N_24737,N_24959);
nand UO_1836 (O_1836,N_24960,N_24836);
or UO_1837 (O_1837,N_24478,N_24497);
xor UO_1838 (O_1838,N_24555,N_24750);
and UO_1839 (O_1839,N_24951,N_24703);
nor UO_1840 (O_1840,N_24413,N_24887);
nand UO_1841 (O_1841,N_24438,N_24666);
nor UO_1842 (O_1842,N_24867,N_24789);
or UO_1843 (O_1843,N_24744,N_24929);
xnor UO_1844 (O_1844,N_24953,N_24765);
and UO_1845 (O_1845,N_24827,N_24928);
or UO_1846 (O_1846,N_24622,N_24611);
and UO_1847 (O_1847,N_24922,N_24869);
nand UO_1848 (O_1848,N_24458,N_24868);
and UO_1849 (O_1849,N_24808,N_24479);
and UO_1850 (O_1850,N_24451,N_24846);
nor UO_1851 (O_1851,N_24418,N_24787);
and UO_1852 (O_1852,N_24770,N_24879);
xor UO_1853 (O_1853,N_24465,N_24856);
and UO_1854 (O_1854,N_24838,N_24945);
xnor UO_1855 (O_1855,N_24933,N_24714);
nand UO_1856 (O_1856,N_24393,N_24947);
nor UO_1857 (O_1857,N_24445,N_24432);
nor UO_1858 (O_1858,N_24540,N_24867);
nor UO_1859 (O_1859,N_24814,N_24601);
xnor UO_1860 (O_1860,N_24594,N_24761);
nor UO_1861 (O_1861,N_24618,N_24448);
or UO_1862 (O_1862,N_24772,N_24835);
and UO_1863 (O_1863,N_24825,N_24616);
nor UO_1864 (O_1864,N_24654,N_24697);
and UO_1865 (O_1865,N_24967,N_24520);
or UO_1866 (O_1866,N_24697,N_24703);
nand UO_1867 (O_1867,N_24508,N_24776);
nand UO_1868 (O_1868,N_24799,N_24509);
and UO_1869 (O_1869,N_24634,N_24867);
xnor UO_1870 (O_1870,N_24505,N_24884);
and UO_1871 (O_1871,N_24456,N_24538);
nand UO_1872 (O_1872,N_24964,N_24501);
or UO_1873 (O_1873,N_24947,N_24511);
xor UO_1874 (O_1874,N_24460,N_24747);
or UO_1875 (O_1875,N_24754,N_24869);
nor UO_1876 (O_1876,N_24864,N_24697);
nand UO_1877 (O_1877,N_24874,N_24577);
nor UO_1878 (O_1878,N_24805,N_24861);
nand UO_1879 (O_1879,N_24577,N_24990);
nand UO_1880 (O_1880,N_24737,N_24699);
nor UO_1881 (O_1881,N_24416,N_24581);
nand UO_1882 (O_1882,N_24532,N_24512);
xor UO_1883 (O_1883,N_24699,N_24890);
xnor UO_1884 (O_1884,N_24487,N_24491);
nand UO_1885 (O_1885,N_24563,N_24595);
nand UO_1886 (O_1886,N_24424,N_24402);
nor UO_1887 (O_1887,N_24638,N_24418);
xor UO_1888 (O_1888,N_24979,N_24817);
or UO_1889 (O_1889,N_24430,N_24896);
nor UO_1890 (O_1890,N_24850,N_24656);
xor UO_1891 (O_1891,N_24648,N_24551);
and UO_1892 (O_1892,N_24535,N_24496);
xor UO_1893 (O_1893,N_24576,N_24585);
nor UO_1894 (O_1894,N_24983,N_24399);
or UO_1895 (O_1895,N_24422,N_24876);
nand UO_1896 (O_1896,N_24910,N_24693);
xor UO_1897 (O_1897,N_24940,N_24418);
nor UO_1898 (O_1898,N_24728,N_24394);
and UO_1899 (O_1899,N_24787,N_24626);
and UO_1900 (O_1900,N_24883,N_24529);
and UO_1901 (O_1901,N_24998,N_24661);
and UO_1902 (O_1902,N_24511,N_24713);
or UO_1903 (O_1903,N_24951,N_24381);
and UO_1904 (O_1904,N_24456,N_24896);
and UO_1905 (O_1905,N_24925,N_24928);
or UO_1906 (O_1906,N_24945,N_24881);
nand UO_1907 (O_1907,N_24739,N_24817);
xnor UO_1908 (O_1908,N_24819,N_24419);
xnor UO_1909 (O_1909,N_24922,N_24502);
nor UO_1910 (O_1910,N_24856,N_24592);
nand UO_1911 (O_1911,N_24376,N_24906);
xor UO_1912 (O_1912,N_24509,N_24659);
or UO_1913 (O_1913,N_24909,N_24612);
xnor UO_1914 (O_1914,N_24675,N_24976);
or UO_1915 (O_1915,N_24620,N_24840);
nand UO_1916 (O_1916,N_24412,N_24773);
or UO_1917 (O_1917,N_24713,N_24749);
and UO_1918 (O_1918,N_24513,N_24906);
and UO_1919 (O_1919,N_24470,N_24760);
nor UO_1920 (O_1920,N_24603,N_24392);
nor UO_1921 (O_1921,N_24496,N_24658);
or UO_1922 (O_1922,N_24895,N_24691);
or UO_1923 (O_1923,N_24933,N_24460);
nand UO_1924 (O_1924,N_24380,N_24777);
nand UO_1925 (O_1925,N_24644,N_24763);
xor UO_1926 (O_1926,N_24501,N_24861);
and UO_1927 (O_1927,N_24864,N_24976);
nand UO_1928 (O_1928,N_24974,N_24479);
nand UO_1929 (O_1929,N_24787,N_24845);
and UO_1930 (O_1930,N_24941,N_24633);
and UO_1931 (O_1931,N_24990,N_24819);
xnor UO_1932 (O_1932,N_24494,N_24753);
nor UO_1933 (O_1933,N_24558,N_24881);
or UO_1934 (O_1934,N_24575,N_24991);
xnor UO_1935 (O_1935,N_24838,N_24647);
nand UO_1936 (O_1936,N_24946,N_24805);
or UO_1937 (O_1937,N_24817,N_24718);
or UO_1938 (O_1938,N_24807,N_24770);
xnor UO_1939 (O_1939,N_24497,N_24971);
and UO_1940 (O_1940,N_24713,N_24655);
or UO_1941 (O_1941,N_24835,N_24775);
nor UO_1942 (O_1942,N_24716,N_24633);
nand UO_1943 (O_1943,N_24719,N_24568);
or UO_1944 (O_1944,N_24740,N_24699);
and UO_1945 (O_1945,N_24905,N_24411);
and UO_1946 (O_1946,N_24703,N_24692);
nor UO_1947 (O_1947,N_24515,N_24802);
or UO_1948 (O_1948,N_24434,N_24385);
xnor UO_1949 (O_1949,N_24659,N_24607);
xor UO_1950 (O_1950,N_24624,N_24637);
xnor UO_1951 (O_1951,N_24936,N_24474);
and UO_1952 (O_1952,N_24463,N_24716);
or UO_1953 (O_1953,N_24732,N_24936);
or UO_1954 (O_1954,N_24496,N_24544);
nand UO_1955 (O_1955,N_24558,N_24671);
and UO_1956 (O_1956,N_24960,N_24714);
nor UO_1957 (O_1957,N_24732,N_24836);
xnor UO_1958 (O_1958,N_24379,N_24778);
or UO_1959 (O_1959,N_24440,N_24630);
nor UO_1960 (O_1960,N_24990,N_24517);
xnor UO_1961 (O_1961,N_24827,N_24934);
nor UO_1962 (O_1962,N_24921,N_24956);
xor UO_1963 (O_1963,N_24864,N_24516);
nand UO_1964 (O_1964,N_24903,N_24690);
or UO_1965 (O_1965,N_24502,N_24660);
or UO_1966 (O_1966,N_24997,N_24797);
nor UO_1967 (O_1967,N_24601,N_24927);
xor UO_1968 (O_1968,N_24887,N_24761);
or UO_1969 (O_1969,N_24623,N_24493);
or UO_1970 (O_1970,N_24662,N_24642);
and UO_1971 (O_1971,N_24788,N_24940);
nand UO_1972 (O_1972,N_24650,N_24690);
xnor UO_1973 (O_1973,N_24505,N_24421);
nand UO_1974 (O_1974,N_24493,N_24421);
xnor UO_1975 (O_1975,N_24706,N_24831);
nand UO_1976 (O_1976,N_24584,N_24574);
xor UO_1977 (O_1977,N_24817,N_24925);
nand UO_1978 (O_1978,N_24814,N_24894);
nand UO_1979 (O_1979,N_24905,N_24767);
or UO_1980 (O_1980,N_24993,N_24553);
nand UO_1981 (O_1981,N_24839,N_24832);
and UO_1982 (O_1982,N_24696,N_24859);
or UO_1983 (O_1983,N_24506,N_24973);
or UO_1984 (O_1984,N_24791,N_24434);
nand UO_1985 (O_1985,N_24554,N_24450);
xor UO_1986 (O_1986,N_24755,N_24689);
xor UO_1987 (O_1987,N_24518,N_24472);
and UO_1988 (O_1988,N_24907,N_24406);
nand UO_1989 (O_1989,N_24987,N_24787);
and UO_1990 (O_1990,N_24544,N_24992);
and UO_1991 (O_1991,N_24964,N_24489);
xnor UO_1992 (O_1992,N_24734,N_24405);
or UO_1993 (O_1993,N_24743,N_24457);
or UO_1994 (O_1994,N_24982,N_24898);
nor UO_1995 (O_1995,N_24378,N_24472);
or UO_1996 (O_1996,N_24882,N_24962);
or UO_1997 (O_1997,N_24545,N_24900);
xor UO_1998 (O_1998,N_24698,N_24691);
or UO_1999 (O_1999,N_24439,N_24700);
xnor UO_2000 (O_2000,N_24779,N_24550);
nor UO_2001 (O_2001,N_24673,N_24897);
xnor UO_2002 (O_2002,N_24486,N_24471);
and UO_2003 (O_2003,N_24493,N_24763);
or UO_2004 (O_2004,N_24747,N_24907);
xor UO_2005 (O_2005,N_24910,N_24465);
xnor UO_2006 (O_2006,N_24608,N_24379);
nor UO_2007 (O_2007,N_24813,N_24933);
nand UO_2008 (O_2008,N_24564,N_24549);
or UO_2009 (O_2009,N_24838,N_24464);
nand UO_2010 (O_2010,N_24420,N_24975);
nand UO_2011 (O_2011,N_24500,N_24999);
xor UO_2012 (O_2012,N_24702,N_24989);
or UO_2013 (O_2013,N_24807,N_24568);
nor UO_2014 (O_2014,N_24426,N_24857);
nor UO_2015 (O_2015,N_24923,N_24532);
nand UO_2016 (O_2016,N_24426,N_24805);
nand UO_2017 (O_2017,N_24936,N_24731);
and UO_2018 (O_2018,N_24975,N_24642);
or UO_2019 (O_2019,N_24681,N_24974);
or UO_2020 (O_2020,N_24480,N_24840);
nor UO_2021 (O_2021,N_24444,N_24672);
nor UO_2022 (O_2022,N_24699,N_24520);
and UO_2023 (O_2023,N_24768,N_24446);
xor UO_2024 (O_2024,N_24830,N_24600);
xor UO_2025 (O_2025,N_24951,N_24839);
or UO_2026 (O_2026,N_24884,N_24622);
nand UO_2027 (O_2027,N_24888,N_24978);
xor UO_2028 (O_2028,N_24855,N_24447);
or UO_2029 (O_2029,N_24621,N_24720);
and UO_2030 (O_2030,N_24661,N_24882);
nor UO_2031 (O_2031,N_24376,N_24839);
xnor UO_2032 (O_2032,N_24893,N_24502);
or UO_2033 (O_2033,N_24862,N_24703);
or UO_2034 (O_2034,N_24930,N_24666);
xor UO_2035 (O_2035,N_24897,N_24755);
or UO_2036 (O_2036,N_24693,N_24884);
and UO_2037 (O_2037,N_24483,N_24996);
and UO_2038 (O_2038,N_24471,N_24753);
nor UO_2039 (O_2039,N_24571,N_24552);
nor UO_2040 (O_2040,N_24865,N_24899);
or UO_2041 (O_2041,N_24834,N_24499);
nor UO_2042 (O_2042,N_24774,N_24565);
xnor UO_2043 (O_2043,N_24961,N_24661);
nor UO_2044 (O_2044,N_24984,N_24711);
or UO_2045 (O_2045,N_24589,N_24471);
xnor UO_2046 (O_2046,N_24742,N_24454);
and UO_2047 (O_2047,N_24698,N_24591);
and UO_2048 (O_2048,N_24997,N_24658);
nor UO_2049 (O_2049,N_24432,N_24430);
nor UO_2050 (O_2050,N_24839,N_24426);
xor UO_2051 (O_2051,N_24926,N_24823);
or UO_2052 (O_2052,N_24736,N_24383);
or UO_2053 (O_2053,N_24477,N_24829);
or UO_2054 (O_2054,N_24624,N_24821);
nor UO_2055 (O_2055,N_24711,N_24471);
nor UO_2056 (O_2056,N_24839,N_24963);
nand UO_2057 (O_2057,N_24631,N_24898);
nor UO_2058 (O_2058,N_24653,N_24539);
nor UO_2059 (O_2059,N_24925,N_24867);
nand UO_2060 (O_2060,N_24752,N_24939);
nor UO_2061 (O_2061,N_24522,N_24383);
or UO_2062 (O_2062,N_24941,N_24563);
nand UO_2063 (O_2063,N_24899,N_24721);
or UO_2064 (O_2064,N_24419,N_24850);
xnor UO_2065 (O_2065,N_24971,N_24568);
and UO_2066 (O_2066,N_24685,N_24563);
nor UO_2067 (O_2067,N_24536,N_24504);
or UO_2068 (O_2068,N_24425,N_24860);
or UO_2069 (O_2069,N_24920,N_24737);
and UO_2070 (O_2070,N_24800,N_24876);
or UO_2071 (O_2071,N_24856,N_24895);
or UO_2072 (O_2072,N_24388,N_24650);
and UO_2073 (O_2073,N_24641,N_24856);
or UO_2074 (O_2074,N_24406,N_24979);
or UO_2075 (O_2075,N_24715,N_24696);
or UO_2076 (O_2076,N_24444,N_24760);
xor UO_2077 (O_2077,N_24498,N_24636);
and UO_2078 (O_2078,N_24614,N_24850);
xor UO_2079 (O_2079,N_24564,N_24552);
nand UO_2080 (O_2080,N_24441,N_24701);
nor UO_2081 (O_2081,N_24543,N_24444);
nor UO_2082 (O_2082,N_24559,N_24985);
or UO_2083 (O_2083,N_24692,N_24824);
nor UO_2084 (O_2084,N_24796,N_24999);
nand UO_2085 (O_2085,N_24497,N_24629);
or UO_2086 (O_2086,N_24819,N_24662);
xor UO_2087 (O_2087,N_24670,N_24910);
and UO_2088 (O_2088,N_24570,N_24634);
xnor UO_2089 (O_2089,N_24848,N_24598);
or UO_2090 (O_2090,N_24953,N_24715);
nand UO_2091 (O_2091,N_24628,N_24412);
nor UO_2092 (O_2092,N_24547,N_24646);
nor UO_2093 (O_2093,N_24615,N_24704);
nand UO_2094 (O_2094,N_24951,N_24688);
nor UO_2095 (O_2095,N_24626,N_24917);
nor UO_2096 (O_2096,N_24798,N_24425);
xnor UO_2097 (O_2097,N_24877,N_24765);
xor UO_2098 (O_2098,N_24382,N_24636);
and UO_2099 (O_2099,N_24755,N_24734);
and UO_2100 (O_2100,N_24400,N_24608);
nand UO_2101 (O_2101,N_24822,N_24866);
and UO_2102 (O_2102,N_24485,N_24952);
nand UO_2103 (O_2103,N_24915,N_24605);
and UO_2104 (O_2104,N_24550,N_24819);
xnor UO_2105 (O_2105,N_24530,N_24950);
xor UO_2106 (O_2106,N_24628,N_24586);
nand UO_2107 (O_2107,N_24472,N_24946);
or UO_2108 (O_2108,N_24794,N_24937);
and UO_2109 (O_2109,N_24571,N_24778);
or UO_2110 (O_2110,N_24682,N_24700);
xor UO_2111 (O_2111,N_24496,N_24513);
xnor UO_2112 (O_2112,N_24863,N_24537);
or UO_2113 (O_2113,N_24417,N_24437);
or UO_2114 (O_2114,N_24816,N_24416);
nand UO_2115 (O_2115,N_24394,N_24905);
nand UO_2116 (O_2116,N_24725,N_24959);
and UO_2117 (O_2117,N_24952,N_24790);
nor UO_2118 (O_2118,N_24420,N_24450);
xor UO_2119 (O_2119,N_24396,N_24872);
and UO_2120 (O_2120,N_24710,N_24381);
or UO_2121 (O_2121,N_24580,N_24639);
xnor UO_2122 (O_2122,N_24500,N_24996);
or UO_2123 (O_2123,N_24606,N_24425);
xor UO_2124 (O_2124,N_24559,N_24537);
nand UO_2125 (O_2125,N_24661,N_24573);
nor UO_2126 (O_2126,N_24992,N_24535);
nor UO_2127 (O_2127,N_24437,N_24737);
and UO_2128 (O_2128,N_24672,N_24804);
nand UO_2129 (O_2129,N_24470,N_24653);
nand UO_2130 (O_2130,N_24519,N_24671);
xnor UO_2131 (O_2131,N_24503,N_24747);
nand UO_2132 (O_2132,N_24711,N_24944);
nand UO_2133 (O_2133,N_24506,N_24733);
nand UO_2134 (O_2134,N_24383,N_24761);
xnor UO_2135 (O_2135,N_24612,N_24706);
and UO_2136 (O_2136,N_24707,N_24962);
xnor UO_2137 (O_2137,N_24940,N_24438);
nand UO_2138 (O_2138,N_24394,N_24864);
nor UO_2139 (O_2139,N_24769,N_24643);
nor UO_2140 (O_2140,N_24450,N_24549);
xor UO_2141 (O_2141,N_24812,N_24782);
nor UO_2142 (O_2142,N_24673,N_24391);
xor UO_2143 (O_2143,N_24587,N_24742);
or UO_2144 (O_2144,N_24450,N_24941);
nor UO_2145 (O_2145,N_24464,N_24589);
nor UO_2146 (O_2146,N_24726,N_24888);
nand UO_2147 (O_2147,N_24975,N_24791);
nand UO_2148 (O_2148,N_24609,N_24487);
and UO_2149 (O_2149,N_24801,N_24791);
and UO_2150 (O_2150,N_24844,N_24818);
or UO_2151 (O_2151,N_24780,N_24676);
and UO_2152 (O_2152,N_24774,N_24526);
or UO_2153 (O_2153,N_24485,N_24461);
nand UO_2154 (O_2154,N_24706,N_24505);
nand UO_2155 (O_2155,N_24589,N_24719);
and UO_2156 (O_2156,N_24834,N_24548);
xnor UO_2157 (O_2157,N_24475,N_24494);
and UO_2158 (O_2158,N_24907,N_24571);
nand UO_2159 (O_2159,N_24952,N_24554);
nand UO_2160 (O_2160,N_24469,N_24823);
nand UO_2161 (O_2161,N_24548,N_24822);
nand UO_2162 (O_2162,N_24567,N_24564);
and UO_2163 (O_2163,N_24378,N_24470);
or UO_2164 (O_2164,N_24904,N_24566);
nor UO_2165 (O_2165,N_24387,N_24674);
or UO_2166 (O_2166,N_24800,N_24432);
and UO_2167 (O_2167,N_24815,N_24785);
xnor UO_2168 (O_2168,N_24438,N_24595);
and UO_2169 (O_2169,N_24947,N_24609);
or UO_2170 (O_2170,N_24425,N_24560);
nor UO_2171 (O_2171,N_24642,N_24727);
nand UO_2172 (O_2172,N_24596,N_24980);
nor UO_2173 (O_2173,N_24633,N_24703);
or UO_2174 (O_2174,N_24458,N_24986);
and UO_2175 (O_2175,N_24773,N_24728);
xor UO_2176 (O_2176,N_24525,N_24921);
and UO_2177 (O_2177,N_24929,N_24764);
or UO_2178 (O_2178,N_24735,N_24613);
nand UO_2179 (O_2179,N_24551,N_24687);
nand UO_2180 (O_2180,N_24966,N_24749);
or UO_2181 (O_2181,N_24454,N_24512);
nor UO_2182 (O_2182,N_24843,N_24704);
and UO_2183 (O_2183,N_24846,N_24593);
or UO_2184 (O_2184,N_24804,N_24520);
nor UO_2185 (O_2185,N_24678,N_24778);
and UO_2186 (O_2186,N_24732,N_24871);
and UO_2187 (O_2187,N_24774,N_24488);
or UO_2188 (O_2188,N_24426,N_24406);
nand UO_2189 (O_2189,N_24723,N_24701);
and UO_2190 (O_2190,N_24767,N_24983);
or UO_2191 (O_2191,N_24463,N_24587);
or UO_2192 (O_2192,N_24660,N_24470);
nor UO_2193 (O_2193,N_24652,N_24584);
or UO_2194 (O_2194,N_24970,N_24784);
nand UO_2195 (O_2195,N_24472,N_24842);
nor UO_2196 (O_2196,N_24752,N_24960);
nor UO_2197 (O_2197,N_24595,N_24572);
xnor UO_2198 (O_2198,N_24882,N_24443);
nor UO_2199 (O_2199,N_24619,N_24485);
or UO_2200 (O_2200,N_24787,N_24723);
and UO_2201 (O_2201,N_24717,N_24825);
nand UO_2202 (O_2202,N_24826,N_24597);
xor UO_2203 (O_2203,N_24582,N_24583);
and UO_2204 (O_2204,N_24436,N_24960);
xnor UO_2205 (O_2205,N_24982,N_24700);
or UO_2206 (O_2206,N_24556,N_24887);
and UO_2207 (O_2207,N_24466,N_24754);
or UO_2208 (O_2208,N_24472,N_24730);
xor UO_2209 (O_2209,N_24698,N_24658);
nor UO_2210 (O_2210,N_24530,N_24651);
xnor UO_2211 (O_2211,N_24873,N_24411);
and UO_2212 (O_2212,N_24500,N_24556);
or UO_2213 (O_2213,N_24952,N_24524);
nor UO_2214 (O_2214,N_24938,N_24901);
xor UO_2215 (O_2215,N_24714,N_24871);
or UO_2216 (O_2216,N_24891,N_24835);
nor UO_2217 (O_2217,N_24380,N_24553);
nor UO_2218 (O_2218,N_24653,N_24425);
or UO_2219 (O_2219,N_24533,N_24526);
or UO_2220 (O_2220,N_24781,N_24391);
xor UO_2221 (O_2221,N_24692,N_24700);
and UO_2222 (O_2222,N_24670,N_24822);
nand UO_2223 (O_2223,N_24819,N_24434);
nor UO_2224 (O_2224,N_24499,N_24970);
xor UO_2225 (O_2225,N_24569,N_24575);
or UO_2226 (O_2226,N_24902,N_24468);
nor UO_2227 (O_2227,N_24887,N_24927);
and UO_2228 (O_2228,N_24990,N_24970);
and UO_2229 (O_2229,N_24506,N_24624);
or UO_2230 (O_2230,N_24909,N_24676);
or UO_2231 (O_2231,N_24553,N_24752);
and UO_2232 (O_2232,N_24514,N_24624);
nor UO_2233 (O_2233,N_24816,N_24534);
xnor UO_2234 (O_2234,N_24614,N_24630);
xnor UO_2235 (O_2235,N_24633,N_24725);
nor UO_2236 (O_2236,N_24680,N_24788);
and UO_2237 (O_2237,N_24535,N_24887);
or UO_2238 (O_2238,N_24978,N_24451);
xnor UO_2239 (O_2239,N_24646,N_24806);
or UO_2240 (O_2240,N_24449,N_24881);
nand UO_2241 (O_2241,N_24564,N_24779);
or UO_2242 (O_2242,N_24469,N_24918);
xnor UO_2243 (O_2243,N_24941,N_24520);
or UO_2244 (O_2244,N_24538,N_24601);
or UO_2245 (O_2245,N_24480,N_24709);
or UO_2246 (O_2246,N_24627,N_24542);
nand UO_2247 (O_2247,N_24975,N_24556);
nor UO_2248 (O_2248,N_24836,N_24435);
nor UO_2249 (O_2249,N_24835,N_24667);
or UO_2250 (O_2250,N_24741,N_24560);
xnor UO_2251 (O_2251,N_24649,N_24612);
nand UO_2252 (O_2252,N_24519,N_24830);
and UO_2253 (O_2253,N_24700,N_24455);
nor UO_2254 (O_2254,N_24599,N_24992);
xnor UO_2255 (O_2255,N_24449,N_24526);
and UO_2256 (O_2256,N_24664,N_24822);
xor UO_2257 (O_2257,N_24655,N_24416);
and UO_2258 (O_2258,N_24627,N_24425);
nand UO_2259 (O_2259,N_24826,N_24934);
nor UO_2260 (O_2260,N_24696,N_24422);
and UO_2261 (O_2261,N_24693,N_24650);
xor UO_2262 (O_2262,N_24554,N_24375);
nand UO_2263 (O_2263,N_24945,N_24601);
nand UO_2264 (O_2264,N_24745,N_24931);
or UO_2265 (O_2265,N_24576,N_24766);
nor UO_2266 (O_2266,N_24532,N_24762);
xor UO_2267 (O_2267,N_24405,N_24627);
xor UO_2268 (O_2268,N_24448,N_24412);
or UO_2269 (O_2269,N_24757,N_24846);
or UO_2270 (O_2270,N_24837,N_24786);
xor UO_2271 (O_2271,N_24469,N_24629);
and UO_2272 (O_2272,N_24879,N_24985);
nor UO_2273 (O_2273,N_24743,N_24505);
and UO_2274 (O_2274,N_24787,N_24976);
and UO_2275 (O_2275,N_24752,N_24397);
xnor UO_2276 (O_2276,N_24466,N_24578);
nor UO_2277 (O_2277,N_24994,N_24956);
nor UO_2278 (O_2278,N_24927,N_24893);
nor UO_2279 (O_2279,N_24891,N_24704);
nor UO_2280 (O_2280,N_24455,N_24482);
xnor UO_2281 (O_2281,N_24656,N_24691);
nor UO_2282 (O_2282,N_24784,N_24930);
xnor UO_2283 (O_2283,N_24411,N_24638);
xnor UO_2284 (O_2284,N_24595,N_24695);
and UO_2285 (O_2285,N_24816,N_24376);
xor UO_2286 (O_2286,N_24781,N_24741);
and UO_2287 (O_2287,N_24872,N_24642);
nand UO_2288 (O_2288,N_24538,N_24440);
xnor UO_2289 (O_2289,N_24711,N_24752);
or UO_2290 (O_2290,N_24900,N_24394);
nor UO_2291 (O_2291,N_24380,N_24506);
nor UO_2292 (O_2292,N_24656,N_24737);
nor UO_2293 (O_2293,N_24967,N_24706);
xnor UO_2294 (O_2294,N_24863,N_24987);
nor UO_2295 (O_2295,N_24512,N_24899);
xnor UO_2296 (O_2296,N_24496,N_24751);
and UO_2297 (O_2297,N_24874,N_24622);
nor UO_2298 (O_2298,N_24885,N_24968);
or UO_2299 (O_2299,N_24606,N_24485);
nor UO_2300 (O_2300,N_24914,N_24380);
or UO_2301 (O_2301,N_24458,N_24490);
nand UO_2302 (O_2302,N_24828,N_24809);
xnor UO_2303 (O_2303,N_24606,N_24767);
nand UO_2304 (O_2304,N_24518,N_24478);
and UO_2305 (O_2305,N_24556,N_24655);
nand UO_2306 (O_2306,N_24612,N_24822);
and UO_2307 (O_2307,N_24894,N_24712);
and UO_2308 (O_2308,N_24456,N_24970);
or UO_2309 (O_2309,N_24967,N_24721);
or UO_2310 (O_2310,N_24750,N_24422);
and UO_2311 (O_2311,N_24700,N_24670);
xor UO_2312 (O_2312,N_24687,N_24966);
nor UO_2313 (O_2313,N_24406,N_24882);
nor UO_2314 (O_2314,N_24518,N_24640);
or UO_2315 (O_2315,N_24992,N_24642);
nand UO_2316 (O_2316,N_24890,N_24921);
nand UO_2317 (O_2317,N_24392,N_24708);
and UO_2318 (O_2318,N_24524,N_24784);
or UO_2319 (O_2319,N_24684,N_24478);
or UO_2320 (O_2320,N_24409,N_24984);
or UO_2321 (O_2321,N_24644,N_24907);
xor UO_2322 (O_2322,N_24746,N_24451);
nor UO_2323 (O_2323,N_24468,N_24833);
or UO_2324 (O_2324,N_24619,N_24797);
and UO_2325 (O_2325,N_24912,N_24778);
xnor UO_2326 (O_2326,N_24659,N_24621);
nor UO_2327 (O_2327,N_24943,N_24711);
or UO_2328 (O_2328,N_24475,N_24469);
and UO_2329 (O_2329,N_24492,N_24803);
nor UO_2330 (O_2330,N_24575,N_24988);
and UO_2331 (O_2331,N_24645,N_24727);
and UO_2332 (O_2332,N_24962,N_24985);
and UO_2333 (O_2333,N_24667,N_24860);
xnor UO_2334 (O_2334,N_24448,N_24741);
xnor UO_2335 (O_2335,N_24791,N_24864);
nor UO_2336 (O_2336,N_24924,N_24829);
nand UO_2337 (O_2337,N_24761,N_24680);
and UO_2338 (O_2338,N_24826,N_24700);
and UO_2339 (O_2339,N_24561,N_24535);
or UO_2340 (O_2340,N_24958,N_24463);
nor UO_2341 (O_2341,N_24633,N_24717);
xnor UO_2342 (O_2342,N_24486,N_24461);
and UO_2343 (O_2343,N_24939,N_24580);
xor UO_2344 (O_2344,N_24410,N_24406);
nand UO_2345 (O_2345,N_24707,N_24803);
and UO_2346 (O_2346,N_24878,N_24738);
nor UO_2347 (O_2347,N_24866,N_24736);
nand UO_2348 (O_2348,N_24645,N_24595);
or UO_2349 (O_2349,N_24641,N_24396);
xnor UO_2350 (O_2350,N_24417,N_24386);
or UO_2351 (O_2351,N_24935,N_24539);
and UO_2352 (O_2352,N_24823,N_24870);
or UO_2353 (O_2353,N_24940,N_24979);
or UO_2354 (O_2354,N_24965,N_24492);
and UO_2355 (O_2355,N_24814,N_24517);
nor UO_2356 (O_2356,N_24420,N_24537);
nand UO_2357 (O_2357,N_24901,N_24663);
xor UO_2358 (O_2358,N_24776,N_24413);
nand UO_2359 (O_2359,N_24708,N_24427);
nor UO_2360 (O_2360,N_24988,N_24716);
and UO_2361 (O_2361,N_24844,N_24860);
and UO_2362 (O_2362,N_24387,N_24419);
nand UO_2363 (O_2363,N_24434,N_24508);
nand UO_2364 (O_2364,N_24723,N_24449);
nand UO_2365 (O_2365,N_24859,N_24564);
nand UO_2366 (O_2366,N_24523,N_24524);
nor UO_2367 (O_2367,N_24637,N_24893);
xnor UO_2368 (O_2368,N_24933,N_24831);
nor UO_2369 (O_2369,N_24390,N_24757);
xnor UO_2370 (O_2370,N_24575,N_24829);
and UO_2371 (O_2371,N_24757,N_24501);
and UO_2372 (O_2372,N_24703,N_24660);
xor UO_2373 (O_2373,N_24558,N_24530);
nand UO_2374 (O_2374,N_24601,N_24780);
nand UO_2375 (O_2375,N_24666,N_24530);
nor UO_2376 (O_2376,N_24557,N_24550);
xor UO_2377 (O_2377,N_24464,N_24767);
xor UO_2378 (O_2378,N_24964,N_24850);
xnor UO_2379 (O_2379,N_24378,N_24874);
nand UO_2380 (O_2380,N_24846,N_24801);
xor UO_2381 (O_2381,N_24583,N_24827);
or UO_2382 (O_2382,N_24774,N_24445);
or UO_2383 (O_2383,N_24776,N_24486);
nand UO_2384 (O_2384,N_24949,N_24489);
nor UO_2385 (O_2385,N_24631,N_24388);
nand UO_2386 (O_2386,N_24847,N_24721);
nand UO_2387 (O_2387,N_24943,N_24459);
xor UO_2388 (O_2388,N_24862,N_24831);
or UO_2389 (O_2389,N_24429,N_24865);
nor UO_2390 (O_2390,N_24838,N_24390);
nor UO_2391 (O_2391,N_24857,N_24835);
nor UO_2392 (O_2392,N_24393,N_24834);
and UO_2393 (O_2393,N_24946,N_24583);
nand UO_2394 (O_2394,N_24493,N_24614);
nand UO_2395 (O_2395,N_24468,N_24509);
nor UO_2396 (O_2396,N_24839,N_24392);
and UO_2397 (O_2397,N_24549,N_24857);
and UO_2398 (O_2398,N_24626,N_24923);
nor UO_2399 (O_2399,N_24503,N_24810);
nor UO_2400 (O_2400,N_24982,N_24495);
nor UO_2401 (O_2401,N_24890,N_24690);
and UO_2402 (O_2402,N_24827,N_24442);
xnor UO_2403 (O_2403,N_24553,N_24610);
xor UO_2404 (O_2404,N_24898,N_24956);
or UO_2405 (O_2405,N_24886,N_24882);
and UO_2406 (O_2406,N_24415,N_24793);
nor UO_2407 (O_2407,N_24757,N_24653);
nand UO_2408 (O_2408,N_24649,N_24751);
and UO_2409 (O_2409,N_24705,N_24486);
xor UO_2410 (O_2410,N_24469,N_24718);
nand UO_2411 (O_2411,N_24922,N_24838);
and UO_2412 (O_2412,N_24536,N_24773);
xnor UO_2413 (O_2413,N_24731,N_24772);
xor UO_2414 (O_2414,N_24626,N_24690);
nor UO_2415 (O_2415,N_24896,N_24505);
nand UO_2416 (O_2416,N_24649,N_24666);
nor UO_2417 (O_2417,N_24432,N_24947);
nor UO_2418 (O_2418,N_24734,N_24967);
xnor UO_2419 (O_2419,N_24817,N_24578);
and UO_2420 (O_2420,N_24499,N_24966);
and UO_2421 (O_2421,N_24672,N_24497);
nor UO_2422 (O_2422,N_24778,N_24684);
xnor UO_2423 (O_2423,N_24530,N_24455);
xnor UO_2424 (O_2424,N_24548,N_24632);
nor UO_2425 (O_2425,N_24983,N_24993);
xnor UO_2426 (O_2426,N_24937,N_24502);
and UO_2427 (O_2427,N_24930,N_24700);
or UO_2428 (O_2428,N_24643,N_24767);
nor UO_2429 (O_2429,N_24668,N_24607);
nor UO_2430 (O_2430,N_24852,N_24659);
and UO_2431 (O_2431,N_24651,N_24750);
or UO_2432 (O_2432,N_24769,N_24542);
nor UO_2433 (O_2433,N_24514,N_24407);
nor UO_2434 (O_2434,N_24963,N_24898);
or UO_2435 (O_2435,N_24844,N_24469);
and UO_2436 (O_2436,N_24812,N_24586);
and UO_2437 (O_2437,N_24847,N_24986);
nand UO_2438 (O_2438,N_24992,N_24678);
nor UO_2439 (O_2439,N_24782,N_24912);
xnor UO_2440 (O_2440,N_24525,N_24977);
or UO_2441 (O_2441,N_24921,N_24955);
or UO_2442 (O_2442,N_24759,N_24376);
nand UO_2443 (O_2443,N_24478,N_24961);
xnor UO_2444 (O_2444,N_24767,N_24559);
or UO_2445 (O_2445,N_24483,N_24526);
xnor UO_2446 (O_2446,N_24913,N_24965);
nand UO_2447 (O_2447,N_24733,N_24799);
nand UO_2448 (O_2448,N_24929,N_24677);
xor UO_2449 (O_2449,N_24808,N_24701);
and UO_2450 (O_2450,N_24880,N_24747);
and UO_2451 (O_2451,N_24726,N_24987);
or UO_2452 (O_2452,N_24393,N_24785);
xnor UO_2453 (O_2453,N_24496,N_24543);
xnor UO_2454 (O_2454,N_24753,N_24796);
xnor UO_2455 (O_2455,N_24848,N_24605);
and UO_2456 (O_2456,N_24386,N_24615);
nor UO_2457 (O_2457,N_24691,N_24634);
nor UO_2458 (O_2458,N_24697,N_24836);
and UO_2459 (O_2459,N_24982,N_24469);
or UO_2460 (O_2460,N_24634,N_24822);
and UO_2461 (O_2461,N_24493,N_24773);
and UO_2462 (O_2462,N_24549,N_24879);
or UO_2463 (O_2463,N_24429,N_24549);
nor UO_2464 (O_2464,N_24485,N_24785);
or UO_2465 (O_2465,N_24800,N_24483);
or UO_2466 (O_2466,N_24693,N_24468);
nor UO_2467 (O_2467,N_24922,N_24736);
and UO_2468 (O_2468,N_24452,N_24592);
nand UO_2469 (O_2469,N_24376,N_24518);
nor UO_2470 (O_2470,N_24816,N_24774);
and UO_2471 (O_2471,N_24539,N_24441);
xor UO_2472 (O_2472,N_24898,N_24882);
or UO_2473 (O_2473,N_24746,N_24460);
nand UO_2474 (O_2474,N_24826,N_24497);
and UO_2475 (O_2475,N_24702,N_24498);
nor UO_2476 (O_2476,N_24475,N_24380);
xor UO_2477 (O_2477,N_24534,N_24780);
nand UO_2478 (O_2478,N_24603,N_24901);
xor UO_2479 (O_2479,N_24664,N_24827);
nor UO_2480 (O_2480,N_24680,N_24513);
nand UO_2481 (O_2481,N_24432,N_24750);
xnor UO_2482 (O_2482,N_24494,N_24891);
or UO_2483 (O_2483,N_24990,N_24652);
nor UO_2484 (O_2484,N_24501,N_24655);
nand UO_2485 (O_2485,N_24740,N_24456);
nand UO_2486 (O_2486,N_24887,N_24642);
and UO_2487 (O_2487,N_24574,N_24978);
xnor UO_2488 (O_2488,N_24400,N_24657);
xnor UO_2489 (O_2489,N_24770,N_24861);
or UO_2490 (O_2490,N_24850,N_24457);
xnor UO_2491 (O_2491,N_24874,N_24589);
and UO_2492 (O_2492,N_24851,N_24750);
nand UO_2493 (O_2493,N_24894,N_24512);
and UO_2494 (O_2494,N_24771,N_24387);
and UO_2495 (O_2495,N_24873,N_24945);
nor UO_2496 (O_2496,N_24393,N_24928);
nor UO_2497 (O_2497,N_24693,N_24873);
and UO_2498 (O_2498,N_24789,N_24985);
and UO_2499 (O_2499,N_24423,N_24603);
xnor UO_2500 (O_2500,N_24757,N_24717);
nand UO_2501 (O_2501,N_24449,N_24507);
nand UO_2502 (O_2502,N_24640,N_24870);
or UO_2503 (O_2503,N_24620,N_24935);
nand UO_2504 (O_2504,N_24561,N_24641);
xnor UO_2505 (O_2505,N_24721,N_24889);
nor UO_2506 (O_2506,N_24532,N_24563);
nor UO_2507 (O_2507,N_24538,N_24816);
nand UO_2508 (O_2508,N_24820,N_24743);
or UO_2509 (O_2509,N_24445,N_24976);
nand UO_2510 (O_2510,N_24779,N_24548);
xor UO_2511 (O_2511,N_24872,N_24703);
nand UO_2512 (O_2512,N_24965,N_24932);
nor UO_2513 (O_2513,N_24868,N_24597);
nand UO_2514 (O_2514,N_24558,N_24464);
xor UO_2515 (O_2515,N_24584,N_24645);
or UO_2516 (O_2516,N_24504,N_24692);
xor UO_2517 (O_2517,N_24772,N_24855);
and UO_2518 (O_2518,N_24863,N_24924);
or UO_2519 (O_2519,N_24437,N_24518);
and UO_2520 (O_2520,N_24467,N_24655);
nor UO_2521 (O_2521,N_24976,N_24707);
nor UO_2522 (O_2522,N_24419,N_24838);
or UO_2523 (O_2523,N_24720,N_24777);
or UO_2524 (O_2524,N_24538,N_24968);
nor UO_2525 (O_2525,N_24904,N_24826);
or UO_2526 (O_2526,N_24648,N_24687);
or UO_2527 (O_2527,N_24560,N_24993);
and UO_2528 (O_2528,N_24878,N_24719);
and UO_2529 (O_2529,N_24975,N_24675);
and UO_2530 (O_2530,N_24453,N_24444);
or UO_2531 (O_2531,N_24595,N_24558);
and UO_2532 (O_2532,N_24812,N_24856);
and UO_2533 (O_2533,N_24880,N_24721);
and UO_2534 (O_2534,N_24414,N_24377);
or UO_2535 (O_2535,N_24698,N_24509);
nor UO_2536 (O_2536,N_24653,N_24658);
and UO_2537 (O_2537,N_24719,N_24644);
xnor UO_2538 (O_2538,N_24881,N_24700);
and UO_2539 (O_2539,N_24855,N_24751);
nand UO_2540 (O_2540,N_24414,N_24713);
nand UO_2541 (O_2541,N_24388,N_24390);
nor UO_2542 (O_2542,N_24812,N_24650);
and UO_2543 (O_2543,N_24731,N_24702);
nand UO_2544 (O_2544,N_24936,N_24984);
nand UO_2545 (O_2545,N_24907,N_24393);
or UO_2546 (O_2546,N_24868,N_24554);
nand UO_2547 (O_2547,N_24706,N_24717);
and UO_2548 (O_2548,N_24667,N_24390);
xnor UO_2549 (O_2549,N_24522,N_24800);
and UO_2550 (O_2550,N_24456,N_24993);
and UO_2551 (O_2551,N_24832,N_24613);
and UO_2552 (O_2552,N_24749,N_24818);
nor UO_2553 (O_2553,N_24556,N_24627);
xnor UO_2554 (O_2554,N_24734,N_24472);
nor UO_2555 (O_2555,N_24860,N_24405);
xor UO_2556 (O_2556,N_24596,N_24583);
nand UO_2557 (O_2557,N_24506,N_24674);
nand UO_2558 (O_2558,N_24664,N_24666);
xor UO_2559 (O_2559,N_24489,N_24896);
and UO_2560 (O_2560,N_24961,N_24923);
xor UO_2561 (O_2561,N_24645,N_24897);
and UO_2562 (O_2562,N_24713,N_24508);
and UO_2563 (O_2563,N_24515,N_24789);
nor UO_2564 (O_2564,N_24795,N_24546);
nor UO_2565 (O_2565,N_24690,N_24671);
nand UO_2566 (O_2566,N_24766,N_24904);
or UO_2567 (O_2567,N_24475,N_24706);
nand UO_2568 (O_2568,N_24800,N_24397);
or UO_2569 (O_2569,N_24746,N_24609);
or UO_2570 (O_2570,N_24507,N_24902);
nand UO_2571 (O_2571,N_24981,N_24888);
or UO_2572 (O_2572,N_24995,N_24469);
and UO_2573 (O_2573,N_24433,N_24749);
xnor UO_2574 (O_2574,N_24592,N_24833);
xnor UO_2575 (O_2575,N_24647,N_24750);
nor UO_2576 (O_2576,N_24573,N_24683);
nor UO_2577 (O_2577,N_24670,N_24518);
or UO_2578 (O_2578,N_24872,N_24413);
xor UO_2579 (O_2579,N_24429,N_24729);
xor UO_2580 (O_2580,N_24857,N_24977);
and UO_2581 (O_2581,N_24875,N_24778);
xor UO_2582 (O_2582,N_24682,N_24746);
or UO_2583 (O_2583,N_24382,N_24724);
or UO_2584 (O_2584,N_24569,N_24725);
or UO_2585 (O_2585,N_24920,N_24427);
nand UO_2586 (O_2586,N_24794,N_24662);
nand UO_2587 (O_2587,N_24375,N_24642);
and UO_2588 (O_2588,N_24497,N_24520);
and UO_2589 (O_2589,N_24725,N_24545);
xor UO_2590 (O_2590,N_24828,N_24390);
or UO_2591 (O_2591,N_24973,N_24561);
and UO_2592 (O_2592,N_24724,N_24888);
xor UO_2593 (O_2593,N_24633,N_24399);
nand UO_2594 (O_2594,N_24593,N_24638);
xor UO_2595 (O_2595,N_24718,N_24830);
xnor UO_2596 (O_2596,N_24652,N_24626);
nor UO_2597 (O_2597,N_24704,N_24892);
nor UO_2598 (O_2598,N_24561,N_24922);
or UO_2599 (O_2599,N_24760,N_24609);
xor UO_2600 (O_2600,N_24548,N_24816);
or UO_2601 (O_2601,N_24697,N_24425);
xor UO_2602 (O_2602,N_24988,N_24849);
nor UO_2603 (O_2603,N_24801,N_24954);
or UO_2604 (O_2604,N_24969,N_24580);
xor UO_2605 (O_2605,N_24570,N_24377);
and UO_2606 (O_2606,N_24567,N_24515);
or UO_2607 (O_2607,N_24716,N_24421);
and UO_2608 (O_2608,N_24878,N_24562);
and UO_2609 (O_2609,N_24635,N_24816);
nor UO_2610 (O_2610,N_24991,N_24622);
xor UO_2611 (O_2611,N_24720,N_24998);
and UO_2612 (O_2612,N_24792,N_24628);
nor UO_2613 (O_2613,N_24412,N_24553);
and UO_2614 (O_2614,N_24543,N_24664);
or UO_2615 (O_2615,N_24391,N_24568);
xor UO_2616 (O_2616,N_24952,N_24875);
nand UO_2617 (O_2617,N_24872,N_24930);
and UO_2618 (O_2618,N_24583,N_24792);
nor UO_2619 (O_2619,N_24584,N_24849);
or UO_2620 (O_2620,N_24778,N_24791);
or UO_2621 (O_2621,N_24836,N_24991);
and UO_2622 (O_2622,N_24737,N_24627);
nor UO_2623 (O_2623,N_24538,N_24452);
nor UO_2624 (O_2624,N_24808,N_24501);
xor UO_2625 (O_2625,N_24628,N_24801);
and UO_2626 (O_2626,N_24828,N_24980);
nor UO_2627 (O_2627,N_24714,N_24623);
or UO_2628 (O_2628,N_24923,N_24479);
nor UO_2629 (O_2629,N_24513,N_24823);
nand UO_2630 (O_2630,N_24711,N_24870);
xnor UO_2631 (O_2631,N_24398,N_24807);
and UO_2632 (O_2632,N_24950,N_24970);
or UO_2633 (O_2633,N_24693,N_24519);
or UO_2634 (O_2634,N_24786,N_24773);
xnor UO_2635 (O_2635,N_24489,N_24518);
xnor UO_2636 (O_2636,N_24886,N_24945);
and UO_2637 (O_2637,N_24659,N_24753);
and UO_2638 (O_2638,N_24598,N_24648);
nor UO_2639 (O_2639,N_24921,N_24696);
nor UO_2640 (O_2640,N_24680,N_24859);
and UO_2641 (O_2641,N_24570,N_24895);
xor UO_2642 (O_2642,N_24535,N_24644);
and UO_2643 (O_2643,N_24901,N_24483);
nor UO_2644 (O_2644,N_24605,N_24633);
xor UO_2645 (O_2645,N_24843,N_24987);
or UO_2646 (O_2646,N_24649,N_24852);
and UO_2647 (O_2647,N_24532,N_24400);
and UO_2648 (O_2648,N_24648,N_24612);
nand UO_2649 (O_2649,N_24672,N_24924);
xnor UO_2650 (O_2650,N_24623,N_24782);
xor UO_2651 (O_2651,N_24655,N_24576);
or UO_2652 (O_2652,N_24631,N_24717);
and UO_2653 (O_2653,N_24876,N_24763);
nand UO_2654 (O_2654,N_24963,N_24447);
and UO_2655 (O_2655,N_24512,N_24942);
xnor UO_2656 (O_2656,N_24603,N_24984);
nor UO_2657 (O_2657,N_24424,N_24972);
xor UO_2658 (O_2658,N_24937,N_24489);
or UO_2659 (O_2659,N_24524,N_24936);
and UO_2660 (O_2660,N_24732,N_24937);
nor UO_2661 (O_2661,N_24631,N_24665);
and UO_2662 (O_2662,N_24667,N_24754);
nand UO_2663 (O_2663,N_24580,N_24849);
or UO_2664 (O_2664,N_24405,N_24631);
nand UO_2665 (O_2665,N_24582,N_24475);
nor UO_2666 (O_2666,N_24868,N_24569);
nand UO_2667 (O_2667,N_24744,N_24490);
and UO_2668 (O_2668,N_24873,N_24606);
xor UO_2669 (O_2669,N_24614,N_24753);
nand UO_2670 (O_2670,N_24565,N_24962);
xnor UO_2671 (O_2671,N_24719,N_24885);
nand UO_2672 (O_2672,N_24580,N_24475);
nor UO_2673 (O_2673,N_24645,N_24531);
or UO_2674 (O_2674,N_24939,N_24527);
or UO_2675 (O_2675,N_24776,N_24814);
or UO_2676 (O_2676,N_24977,N_24645);
nor UO_2677 (O_2677,N_24860,N_24641);
or UO_2678 (O_2678,N_24542,N_24900);
or UO_2679 (O_2679,N_24767,N_24472);
or UO_2680 (O_2680,N_24777,N_24749);
nor UO_2681 (O_2681,N_24404,N_24966);
and UO_2682 (O_2682,N_24440,N_24472);
nand UO_2683 (O_2683,N_24755,N_24477);
and UO_2684 (O_2684,N_24387,N_24611);
and UO_2685 (O_2685,N_24723,N_24630);
or UO_2686 (O_2686,N_24878,N_24995);
and UO_2687 (O_2687,N_24667,N_24921);
or UO_2688 (O_2688,N_24761,N_24811);
xor UO_2689 (O_2689,N_24459,N_24856);
and UO_2690 (O_2690,N_24818,N_24981);
nand UO_2691 (O_2691,N_24742,N_24605);
xnor UO_2692 (O_2692,N_24948,N_24434);
nand UO_2693 (O_2693,N_24906,N_24876);
or UO_2694 (O_2694,N_24799,N_24418);
nand UO_2695 (O_2695,N_24402,N_24382);
or UO_2696 (O_2696,N_24809,N_24390);
xnor UO_2697 (O_2697,N_24954,N_24513);
or UO_2698 (O_2698,N_24734,N_24525);
or UO_2699 (O_2699,N_24892,N_24573);
and UO_2700 (O_2700,N_24901,N_24948);
and UO_2701 (O_2701,N_24680,N_24457);
nand UO_2702 (O_2702,N_24934,N_24637);
nand UO_2703 (O_2703,N_24909,N_24522);
nor UO_2704 (O_2704,N_24591,N_24981);
xor UO_2705 (O_2705,N_24649,N_24483);
nand UO_2706 (O_2706,N_24563,N_24728);
nor UO_2707 (O_2707,N_24654,N_24610);
or UO_2708 (O_2708,N_24464,N_24810);
nor UO_2709 (O_2709,N_24683,N_24943);
and UO_2710 (O_2710,N_24725,N_24714);
and UO_2711 (O_2711,N_24599,N_24871);
xnor UO_2712 (O_2712,N_24795,N_24488);
nand UO_2713 (O_2713,N_24740,N_24737);
xor UO_2714 (O_2714,N_24719,N_24839);
xnor UO_2715 (O_2715,N_24405,N_24402);
and UO_2716 (O_2716,N_24456,N_24547);
nor UO_2717 (O_2717,N_24994,N_24509);
and UO_2718 (O_2718,N_24563,N_24375);
xor UO_2719 (O_2719,N_24789,N_24925);
nor UO_2720 (O_2720,N_24604,N_24527);
nor UO_2721 (O_2721,N_24666,N_24473);
xnor UO_2722 (O_2722,N_24409,N_24411);
nor UO_2723 (O_2723,N_24808,N_24407);
nor UO_2724 (O_2724,N_24865,N_24617);
nor UO_2725 (O_2725,N_24414,N_24401);
and UO_2726 (O_2726,N_24543,N_24914);
and UO_2727 (O_2727,N_24773,N_24771);
and UO_2728 (O_2728,N_24707,N_24668);
and UO_2729 (O_2729,N_24587,N_24554);
xor UO_2730 (O_2730,N_24505,N_24716);
nand UO_2731 (O_2731,N_24703,N_24671);
xnor UO_2732 (O_2732,N_24998,N_24794);
nand UO_2733 (O_2733,N_24578,N_24986);
and UO_2734 (O_2734,N_24710,N_24519);
or UO_2735 (O_2735,N_24714,N_24870);
xor UO_2736 (O_2736,N_24746,N_24918);
xor UO_2737 (O_2737,N_24712,N_24401);
and UO_2738 (O_2738,N_24688,N_24616);
or UO_2739 (O_2739,N_24942,N_24865);
nor UO_2740 (O_2740,N_24487,N_24794);
and UO_2741 (O_2741,N_24896,N_24440);
and UO_2742 (O_2742,N_24700,N_24470);
xnor UO_2743 (O_2743,N_24494,N_24607);
or UO_2744 (O_2744,N_24856,N_24849);
nor UO_2745 (O_2745,N_24971,N_24397);
and UO_2746 (O_2746,N_24644,N_24931);
xnor UO_2747 (O_2747,N_24866,N_24536);
nand UO_2748 (O_2748,N_24738,N_24732);
xor UO_2749 (O_2749,N_24450,N_24683);
or UO_2750 (O_2750,N_24380,N_24907);
nor UO_2751 (O_2751,N_24532,N_24842);
and UO_2752 (O_2752,N_24616,N_24552);
and UO_2753 (O_2753,N_24760,N_24633);
or UO_2754 (O_2754,N_24685,N_24865);
or UO_2755 (O_2755,N_24411,N_24642);
nand UO_2756 (O_2756,N_24913,N_24756);
xor UO_2757 (O_2757,N_24847,N_24754);
xor UO_2758 (O_2758,N_24526,N_24438);
nand UO_2759 (O_2759,N_24944,N_24929);
nor UO_2760 (O_2760,N_24534,N_24563);
or UO_2761 (O_2761,N_24726,N_24603);
xnor UO_2762 (O_2762,N_24426,N_24623);
nand UO_2763 (O_2763,N_24769,N_24549);
nand UO_2764 (O_2764,N_24754,N_24959);
nand UO_2765 (O_2765,N_24588,N_24467);
and UO_2766 (O_2766,N_24756,N_24464);
nor UO_2767 (O_2767,N_24860,N_24458);
and UO_2768 (O_2768,N_24865,N_24828);
nor UO_2769 (O_2769,N_24595,N_24507);
and UO_2770 (O_2770,N_24560,N_24538);
nand UO_2771 (O_2771,N_24998,N_24935);
xnor UO_2772 (O_2772,N_24516,N_24839);
or UO_2773 (O_2773,N_24970,N_24559);
or UO_2774 (O_2774,N_24580,N_24762);
xor UO_2775 (O_2775,N_24790,N_24433);
and UO_2776 (O_2776,N_24625,N_24587);
and UO_2777 (O_2777,N_24785,N_24501);
and UO_2778 (O_2778,N_24496,N_24931);
nor UO_2779 (O_2779,N_24435,N_24787);
nand UO_2780 (O_2780,N_24769,N_24567);
or UO_2781 (O_2781,N_24745,N_24509);
and UO_2782 (O_2782,N_24970,N_24925);
and UO_2783 (O_2783,N_24475,N_24511);
and UO_2784 (O_2784,N_24568,N_24988);
and UO_2785 (O_2785,N_24600,N_24823);
nand UO_2786 (O_2786,N_24452,N_24971);
nand UO_2787 (O_2787,N_24821,N_24504);
and UO_2788 (O_2788,N_24997,N_24855);
nand UO_2789 (O_2789,N_24502,N_24573);
xnor UO_2790 (O_2790,N_24524,N_24651);
nand UO_2791 (O_2791,N_24978,N_24663);
nand UO_2792 (O_2792,N_24677,N_24992);
nor UO_2793 (O_2793,N_24400,N_24503);
or UO_2794 (O_2794,N_24666,N_24849);
xnor UO_2795 (O_2795,N_24788,N_24902);
xnor UO_2796 (O_2796,N_24468,N_24936);
and UO_2797 (O_2797,N_24973,N_24696);
xor UO_2798 (O_2798,N_24717,N_24754);
nor UO_2799 (O_2799,N_24793,N_24858);
and UO_2800 (O_2800,N_24850,N_24747);
and UO_2801 (O_2801,N_24416,N_24564);
nor UO_2802 (O_2802,N_24505,N_24570);
and UO_2803 (O_2803,N_24707,N_24452);
nand UO_2804 (O_2804,N_24731,N_24859);
nand UO_2805 (O_2805,N_24515,N_24414);
nor UO_2806 (O_2806,N_24628,N_24639);
and UO_2807 (O_2807,N_24909,N_24375);
or UO_2808 (O_2808,N_24719,N_24929);
or UO_2809 (O_2809,N_24531,N_24777);
and UO_2810 (O_2810,N_24823,N_24884);
and UO_2811 (O_2811,N_24552,N_24473);
nand UO_2812 (O_2812,N_24869,N_24874);
or UO_2813 (O_2813,N_24967,N_24959);
or UO_2814 (O_2814,N_24942,N_24610);
nand UO_2815 (O_2815,N_24387,N_24918);
nand UO_2816 (O_2816,N_24534,N_24763);
nor UO_2817 (O_2817,N_24947,N_24966);
nand UO_2818 (O_2818,N_24897,N_24815);
or UO_2819 (O_2819,N_24897,N_24771);
and UO_2820 (O_2820,N_24557,N_24723);
nor UO_2821 (O_2821,N_24592,N_24989);
and UO_2822 (O_2822,N_24385,N_24455);
nand UO_2823 (O_2823,N_24577,N_24725);
or UO_2824 (O_2824,N_24507,N_24746);
nor UO_2825 (O_2825,N_24625,N_24835);
nand UO_2826 (O_2826,N_24438,N_24976);
xor UO_2827 (O_2827,N_24648,N_24415);
nand UO_2828 (O_2828,N_24804,N_24928);
nand UO_2829 (O_2829,N_24477,N_24460);
or UO_2830 (O_2830,N_24626,N_24681);
or UO_2831 (O_2831,N_24832,N_24409);
nor UO_2832 (O_2832,N_24779,N_24723);
nor UO_2833 (O_2833,N_24576,N_24578);
nand UO_2834 (O_2834,N_24965,N_24552);
and UO_2835 (O_2835,N_24433,N_24815);
xor UO_2836 (O_2836,N_24878,N_24563);
and UO_2837 (O_2837,N_24937,N_24793);
nor UO_2838 (O_2838,N_24912,N_24952);
and UO_2839 (O_2839,N_24676,N_24918);
xor UO_2840 (O_2840,N_24546,N_24376);
nor UO_2841 (O_2841,N_24455,N_24645);
xnor UO_2842 (O_2842,N_24413,N_24404);
nand UO_2843 (O_2843,N_24565,N_24685);
nand UO_2844 (O_2844,N_24586,N_24462);
xnor UO_2845 (O_2845,N_24920,N_24903);
nor UO_2846 (O_2846,N_24840,N_24860);
and UO_2847 (O_2847,N_24520,N_24743);
and UO_2848 (O_2848,N_24542,N_24879);
xor UO_2849 (O_2849,N_24415,N_24905);
nand UO_2850 (O_2850,N_24391,N_24955);
nor UO_2851 (O_2851,N_24755,N_24978);
or UO_2852 (O_2852,N_24396,N_24805);
xnor UO_2853 (O_2853,N_24403,N_24802);
or UO_2854 (O_2854,N_24695,N_24969);
and UO_2855 (O_2855,N_24460,N_24455);
xor UO_2856 (O_2856,N_24723,N_24726);
nor UO_2857 (O_2857,N_24422,N_24802);
xnor UO_2858 (O_2858,N_24834,N_24676);
xor UO_2859 (O_2859,N_24609,N_24720);
nor UO_2860 (O_2860,N_24521,N_24733);
and UO_2861 (O_2861,N_24710,N_24382);
and UO_2862 (O_2862,N_24789,N_24819);
and UO_2863 (O_2863,N_24441,N_24597);
and UO_2864 (O_2864,N_24680,N_24398);
and UO_2865 (O_2865,N_24959,N_24423);
or UO_2866 (O_2866,N_24772,N_24684);
and UO_2867 (O_2867,N_24657,N_24744);
and UO_2868 (O_2868,N_24586,N_24682);
or UO_2869 (O_2869,N_24526,N_24757);
nand UO_2870 (O_2870,N_24610,N_24860);
nor UO_2871 (O_2871,N_24422,N_24570);
or UO_2872 (O_2872,N_24447,N_24745);
nand UO_2873 (O_2873,N_24791,N_24677);
and UO_2874 (O_2874,N_24728,N_24622);
xnor UO_2875 (O_2875,N_24970,N_24571);
xor UO_2876 (O_2876,N_24821,N_24879);
nor UO_2877 (O_2877,N_24795,N_24712);
xnor UO_2878 (O_2878,N_24664,N_24631);
xor UO_2879 (O_2879,N_24463,N_24661);
xor UO_2880 (O_2880,N_24931,N_24732);
xnor UO_2881 (O_2881,N_24583,N_24468);
or UO_2882 (O_2882,N_24664,N_24891);
nor UO_2883 (O_2883,N_24762,N_24456);
and UO_2884 (O_2884,N_24577,N_24824);
xor UO_2885 (O_2885,N_24754,N_24735);
nand UO_2886 (O_2886,N_24484,N_24779);
and UO_2887 (O_2887,N_24503,N_24378);
nor UO_2888 (O_2888,N_24384,N_24770);
xnor UO_2889 (O_2889,N_24490,N_24672);
xor UO_2890 (O_2890,N_24401,N_24912);
or UO_2891 (O_2891,N_24385,N_24971);
nor UO_2892 (O_2892,N_24793,N_24669);
nand UO_2893 (O_2893,N_24489,N_24451);
nor UO_2894 (O_2894,N_24489,N_24812);
nor UO_2895 (O_2895,N_24592,N_24838);
nor UO_2896 (O_2896,N_24763,N_24779);
or UO_2897 (O_2897,N_24431,N_24773);
nand UO_2898 (O_2898,N_24760,N_24491);
nor UO_2899 (O_2899,N_24773,N_24886);
and UO_2900 (O_2900,N_24447,N_24684);
and UO_2901 (O_2901,N_24568,N_24764);
xnor UO_2902 (O_2902,N_24630,N_24730);
and UO_2903 (O_2903,N_24614,N_24944);
and UO_2904 (O_2904,N_24621,N_24909);
nand UO_2905 (O_2905,N_24666,N_24481);
or UO_2906 (O_2906,N_24628,N_24839);
and UO_2907 (O_2907,N_24919,N_24493);
and UO_2908 (O_2908,N_24893,N_24887);
or UO_2909 (O_2909,N_24905,N_24633);
xor UO_2910 (O_2910,N_24409,N_24550);
or UO_2911 (O_2911,N_24698,N_24774);
and UO_2912 (O_2912,N_24689,N_24666);
xnor UO_2913 (O_2913,N_24873,N_24978);
xor UO_2914 (O_2914,N_24695,N_24487);
nor UO_2915 (O_2915,N_24968,N_24559);
nor UO_2916 (O_2916,N_24506,N_24675);
nor UO_2917 (O_2917,N_24411,N_24901);
xnor UO_2918 (O_2918,N_24844,N_24995);
xnor UO_2919 (O_2919,N_24439,N_24432);
xor UO_2920 (O_2920,N_24571,N_24940);
and UO_2921 (O_2921,N_24888,N_24906);
nor UO_2922 (O_2922,N_24529,N_24636);
xnor UO_2923 (O_2923,N_24405,N_24964);
and UO_2924 (O_2924,N_24561,N_24974);
and UO_2925 (O_2925,N_24852,N_24967);
nand UO_2926 (O_2926,N_24398,N_24416);
nor UO_2927 (O_2927,N_24955,N_24954);
xnor UO_2928 (O_2928,N_24997,N_24396);
xnor UO_2929 (O_2929,N_24449,N_24795);
xor UO_2930 (O_2930,N_24451,N_24814);
nor UO_2931 (O_2931,N_24737,N_24520);
and UO_2932 (O_2932,N_24712,N_24758);
or UO_2933 (O_2933,N_24939,N_24473);
or UO_2934 (O_2934,N_24553,N_24926);
and UO_2935 (O_2935,N_24580,N_24466);
xnor UO_2936 (O_2936,N_24751,N_24508);
or UO_2937 (O_2937,N_24881,N_24694);
xor UO_2938 (O_2938,N_24791,N_24421);
or UO_2939 (O_2939,N_24580,N_24912);
nand UO_2940 (O_2940,N_24727,N_24700);
nor UO_2941 (O_2941,N_24774,N_24810);
nor UO_2942 (O_2942,N_24655,N_24522);
nor UO_2943 (O_2943,N_24585,N_24670);
xnor UO_2944 (O_2944,N_24530,N_24544);
xnor UO_2945 (O_2945,N_24817,N_24974);
xor UO_2946 (O_2946,N_24962,N_24634);
and UO_2947 (O_2947,N_24989,N_24730);
nor UO_2948 (O_2948,N_24401,N_24662);
and UO_2949 (O_2949,N_24715,N_24417);
nand UO_2950 (O_2950,N_24552,N_24578);
nand UO_2951 (O_2951,N_24655,N_24660);
or UO_2952 (O_2952,N_24942,N_24673);
and UO_2953 (O_2953,N_24685,N_24517);
xor UO_2954 (O_2954,N_24838,N_24842);
nor UO_2955 (O_2955,N_24708,N_24638);
and UO_2956 (O_2956,N_24796,N_24663);
and UO_2957 (O_2957,N_24733,N_24668);
xor UO_2958 (O_2958,N_24620,N_24948);
nor UO_2959 (O_2959,N_24971,N_24547);
xnor UO_2960 (O_2960,N_24754,N_24681);
nor UO_2961 (O_2961,N_24719,N_24454);
xor UO_2962 (O_2962,N_24391,N_24915);
nand UO_2963 (O_2963,N_24535,N_24634);
or UO_2964 (O_2964,N_24981,N_24723);
nand UO_2965 (O_2965,N_24669,N_24397);
and UO_2966 (O_2966,N_24900,N_24831);
and UO_2967 (O_2967,N_24963,N_24421);
or UO_2968 (O_2968,N_24851,N_24540);
nor UO_2969 (O_2969,N_24474,N_24768);
and UO_2970 (O_2970,N_24657,N_24416);
and UO_2971 (O_2971,N_24896,N_24679);
xnor UO_2972 (O_2972,N_24401,N_24378);
nor UO_2973 (O_2973,N_24690,N_24464);
nand UO_2974 (O_2974,N_24848,N_24796);
and UO_2975 (O_2975,N_24722,N_24936);
and UO_2976 (O_2976,N_24439,N_24603);
nand UO_2977 (O_2977,N_24422,N_24623);
nand UO_2978 (O_2978,N_24705,N_24696);
xnor UO_2979 (O_2979,N_24570,N_24989);
xnor UO_2980 (O_2980,N_24432,N_24913);
nor UO_2981 (O_2981,N_24538,N_24449);
or UO_2982 (O_2982,N_24981,N_24745);
xor UO_2983 (O_2983,N_24789,N_24796);
xor UO_2984 (O_2984,N_24544,N_24549);
nor UO_2985 (O_2985,N_24995,N_24444);
nor UO_2986 (O_2986,N_24455,N_24950);
and UO_2987 (O_2987,N_24756,N_24794);
and UO_2988 (O_2988,N_24692,N_24498);
nor UO_2989 (O_2989,N_24787,N_24663);
nor UO_2990 (O_2990,N_24624,N_24632);
nor UO_2991 (O_2991,N_24506,N_24734);
nand UO_2992 (O_2992,N_24375,N_24961);
or UO_2993 (O_2993,N_24783,N_24511);
nor UO_2994 (O_2994,N_24437,N_24769);
and UO_2995 (O_2995,N_24581,N_24478);
nand UO_2996 (O_2996,N_24947,N_24495);
and UO_2997 (O_2997,N_24698,N_24583);
nor UO_2998 (O_2998,N_24791,N_24980);
nand UO_2999 (O_2999,N_24791,N_24429);
endmodule