module basic_5000_50000_5000_100_levels_10xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999,N_30000,N_30001,N_30002,N_30003,N_30004,N_30005,N_30006,N_30007,N_30008,N_30009,N_30010,N_30011,N_30012,N_30013,N_30014,N_30015,N_30016,N_30017,N_30018,N_30019,N_30020,N_30021,N_30022,N_30023,N_30024,N_30025,N_30026,N_30027,N_30028,N_30029,N_30030,N_30031,N_30032,N_30033,N_30034,N_30035,N_30036,N_30037,N_30038,N_30039,N_30040,N_30041,N_30042,N_30043,N_30044,N_30045,N_30046,N_30047,N_30048,N_30049,N_30050,N_30051,N_30052,N_30053,N_30054,N_30055,N_30056,N_30057,N_30058,N_30059,N_30060,N_30061,N_30062,N_30063,N_30064,N_30065,N_30066,N_30067,N_30068,N_30069,N_30070,N_30071,N_30072,N_30073,N_30074,N_30075,N_30076,N_30077,N_30078,N_30079,N_30080,N_30081,N_30082,N_30083,N_30084,N_30085,N_30086,N_30087,N_30088,N_30089,N_30090,N_30091,N_30092,N_30093,N_30094,N_30095,N_30096,N_30097,N_30098,N_30099,N_30100,N_30101,N_30102,N_30103,N_30104,N_30105,N_30106,N_30107,N_30108,N_30109,N_30110,N_30111,N_30112,N_30113,N_30114,N_30115,N_30116,N_30117,N_30118,N_30119,N_30120,N_30121,N_30122,N_30123,N_30124,N_30125,N_30126,N_30127,N_30128,N_30129,N_30130,N_30131,N_30132,N_30133,N_30134,N_30135,N_30136,N_30137,N_30138,N_30139,N_30140,N_30141,N_30142,N_30143,N_30144,N_30145,N_30146,N_30147,N_30148,N_30149,N_30150,N_30151,N_30152,N_30153,N_30154,N_30155,N_30156,N_30157,N_30158,N_30159,N_30160,N_30161,N_30162,N_30163,N_30164,N_30165,N_30166,N_30167,N_30168,N_30169,N_30170,N_30171,N_30172,N_30173,N_30174,N_30175,N_30176,N_30177,N_30178,N_30179,N_30180,N_30181,N_30182,N_30183,N_30184,N_30185,N_30186,N_30187,N_30188,N_30189,N_30190,N_30191,N_30192,N_30193,N_30194,N_30195,N_30196,N_30197,N_30198,N_30199,N_30200,N_30201,N_30202,N_30203,N_30204,N_30205,N_30206,N_30207,N_30208,N_30209,N_30210,N_30211,N_30212,N_30213,N_30214,N_30215,N_30216,N_30217,N_30218,N_30219,N_30220,N_30221,N_30222,N_30223,N_30224,N_30225,N_30226,N_30227,N_30228,N_30229,N_30230,N_30231,N_30232,N_30233,N_30234,N_30235,N_30236,N_30237,N_30238,N_30239,N_30240,N_30241,N_30242,N_30243,N_30244,N_30245,N_30246,N_30247,N_30248,N_30249,N_30250,N_30251,N_30252,N_30253,N_30254,N_30255,N_30256,N_30257,N_30258,N_30259,N_30260,N_30261,N_30262,N_30263,N_30264,N_30265,N_30266,N_30267,N_30268,N_30269,N_30270,N_30271,N_30272,N_30273,N_30274,N_30275,N_30276,N_30277,N_30278,N_30279,N_30280,N_30281,N_30282,N_30283,N_30284,N_30285,N_30286,N_30287,N_30288,N_30289,N_30290,N_30291,N_30292,N_30293,N_30294,N_30295,N_30296,N_30297,N_30298,N_30299,N_30300,N_30301,N_30302,N_30303,N_30304,N_30305,N_30306,N_30307,N_30308,N_30309,N_30310,N_30311,N_30312,N_30313,N_30314,N_30315,N_30316,N_30317,N_30318,N_30319,N_30320,N_30321,N_30322,N_30323,N_30324,N_30325,N_30326,N_30327,N_30328,N_30329,N_30330,N_30331,N_30332,N_30333,N_30334,N_30335,N_30336,N_30337,N_30338,N_30339,N_30340,N_30341,N_30342,N_30343,N_30344,N_30345,N_30346,N_30347,N_30348,N_30349,N_30350,N_30351,N_30352,N_30353,N_30354,N_30355,N_30356,N_30357,N_30358,N_30359,N_30360,N_30361,N_30362,N_30363,N_30364,N_30365,N_30366,N_30367,N_30368,N_30369,N_30370,N_30371,N_30372,N_30373,N_30374,N_30375,N_30376,N_30377,N_30378,N_30379,N_30380,N_30381,N_30382,N_30383,N_30384,N_30385,N_30386,N_30387,N_30388,N_30389,N_30390,N_30391,N_30392,N_30393,N_30394,N_30395,N_30396,N_30397,N_30398,N_30399,N_30400,N_30401,N_30402,N_30403,N_30404,N_30405,N_30406,N_30407,N_30408,N_30409,N_30410,N_30411,N_30412,N_30413,N_30414,N_30415,N_30416,N_30417,N_30418,N_30419,N_30420,N_30421,N_30422,N_30423,N_30424,N_30425,N_30426,N_30427,N_30428,N_30429,N_30430,N_30431,N_30432,N_30433,N_30434,N_30435,N_30436,N_30437,N_30438,N_30439,N_30440,N_30441,N_30442,N_30443,N_30444,N_30445,N_30446,N_30447,N_30448,N_30449,N_30450,N_30451,N_30452,N_30453,N_30454,N_30455,N_30456,N_30457,N_30458,N_30459,N_30460,N_30461,N_30462,N_30463,N_30464,N_30465,N_30466,N_30467,N_30468,N_30469,N_30470,N_30471,N_30472,N_30473,N_30474,N_30475,N_30476,N_30477,N_30478,N_30479,N_30480,N_30481,N_30482,N_30483,N_30484,N_30485,N_30486,N_30487,N_30488,N_30489,N_30490,N_30491,N_30492,N_30493,N_30494,N_30495,N_30496,N_30497,N_30498,N_30499,N_30500,N_30501,N_30502,N_30503,N_30504,N_30505,N_30506,N_30507,N_30508,N_30509,N_30510,N_30511,N_30512,N_30513,N_30514,N_30515,N_30516,N_30517,N_30518,N_30519,N_30520,N_30521,N_30522,N_30523,N_30524,N_30525,N_30526,N_30527,N_30528,N_30529,N_30530,N_30531,N_30532,N_30533,N_30534,N_30535,N_30536,N_30537,N_30538,N_30539,N_30540,N_30541,N_30542,N_30543,N_30544,N_30545,N_30546,N_30547,N_30548,N_30549,N_30550,N_30551,N_30552,N_30553,N_30554,N_30555,N_30556,N_30557,N_30558,N_30559,N_30560,N_30561,N_30562,N_30563,N_30564,N_30565,N_30566,N_30567,N_30568,N_30569,N_30570,N_30571,N_30572,N_30573,N_30574,N_30575,N_30576,N_30577,N_30578,N_30579,N_30580,N_30581,N_30582,N_30583,N_30584,N_30585,N_30586,N_30587,N_30588,N_30589,N_30590,N_30591,N_30592,N_30593,N_30594,N_30595,N_30596,N_30597,N_30598,N_30599,N_30600,N_30601,N_30602,N_30603,N_30604,N_30605,N_30606,N_30607,N_30608,N_30609,N_30610,N_30611,N_30612,N_30613,N_30614,N_30615,N_30616,N_30617,N_30618,N_30619,N_30620,N_30621,N_30622,N_30623,N_30624,N_30625,N_30626,N_30627,N_30628,N_30629,N_30630,N_30631,N_30632,N_30633,N_30634,N_30635,N_30636,N_30637,N_30638,N_30639,N_30640,N_30641,N_30642,N_30643,N_30644,N_30645,N_30646,N_30647,N_30648,N_30649,N_30650,N_30651,N_30652,N_30653,N_30654,N_30655,N_30656,N_30657,N_30658,N_30659,N_30660,N_30661,N_30662,N_30663,N_30664,N_30665,N_30666,N_30667,N_30668,N_30669,N_30670,N_30671,N_30672,N_30673,N_30674,N_30675,N_30676,N_30677,N_30678,N_30679,N_30680,N_30681,N_30682,N_30683,N_30684,N_30685,N_30686,N_30687,N_30688,N_30689,N_30690,N_30691,N_30692,N_30693,N_30694,N_30695,N_30696,N_30697,N_30698,N_30699,N_30700,N_30701,N_30702,N_30703,N_30704,N_30705,N_30706,N_30707,N_30708,N_30709,N_30710,N_30711,N_30712,N_30713,N_30714,N_30715,N_30716,N_30717,N_30718,N_30719,N_30720,N_30721,N_30722,N_30723,N_30724,N_30725,N_30726,N_30727,N_30728,N_30729,N_30730,N_30731,N_30732,N_30733,N_30734,N_30735,N_30736,N_30737,N_30738,N_30739,N_30740,N_30741,N_30742,N_30743,N_30744,N_30745,N_30746,N_30747,N_30748,N_30749,N_30750,N_30751,N_30752,N_30753,N_30754,N_30755,N_30756,N_30757,N_30758,N_30759,N_30760,N_30761,N_30762,N_30763,N_30764,N_30765,N_30766,N_30767,N_30768,N_30769,N_30770,N_30771,N_30772,N_30773,N_30774,N_30775,N_30776,N_30777,N_30778,N_30779,N_30780,N_30781,N_30782,N_30783,N_30784,N_30785,N_30786,N_30787,N_30788,N_30789,N_30790,N_30791,N_30792,N_30793,N_30794,N_30795,N_30796,N_30797,N_30798,N_30799,N_30800,N_30801,N_30802,N_30803,N_30804,N_30805,N_30806,N_30807,N_30808,N_30809,N_30810,N_30811,N_30812,N_30813,N_30814,N_30815,N_30816,N_30817,N_30818,N_30819,N_30820,N_30821,N_30822,N_30823,N_30824,N_30825,N_30826,N_30827,N_30828,N_30829,N_30830,N_30831,N_30832,N_30833,N_30834,N_30835,N_30836,N_30837,N_30838,N_30839,N_30840,N_30841,N_30842,N_30843,N_30844,N_30845,N_30846,N_30847,N_30848,N_30849,N_30850,N_30851,N_30852,N_30853,N_30854,N_30855,N_30856,N_30857,N_30858,N_30859,N_30860,N_30861,N_30862,N_30863,N_30864,N_30865,N_30866,N_30867,N_30868,N_30869,N_30870,N_30871,N_30872,N_30873,N_30874,N_30875,N_30876,N_30877,N_30878,N_30879,N_30880,N_30881,N_30882,N_30883,N_30884,N_30885,N_30886,N_30887,N_30888,N_30889,N_30890,N_30891,N_30892,N_30893,N_30894,N_30895,N_30896,N_30897,N_30898,N_30899,N_30900,N_30901,N_30902,N_30903,N_30904,N_30905,N_30906,N_30907,N_30908,N_30909,N_30910,N_30911,N_30912,N_30913,N_30914,N_30915,N_30916,N_30917,N_30918,N_30919,N_30920,N_30921,N_30922,N_30923,N_30924,N_30925,N_30926,N_30927,N_30928,N_30929,N_30930,N_30931,N_30932,N_30933,N_30934,N_30935,N_30936,N_30937,N_30938,N_30939,N_30940,N_30941,N_30942,N_30943,N_30944,N_30945,N_30946,N_30947,N_30948,N_30949,N_30950,N_30951,N_30952,N_30953,N_30954,N_30955,N_30956,N_30957,N_30958,N_30959,N_30960,N_30961,N_30962,N_30963,N_30964,N_30965,N_30966,N_30967,N_30968,N_30969,N_30970,N_30971,N_30972,N_30973,N_30974,N_30975,N_30976,N_30977,N_30978,N_30979,N_30980,N_30981,N_30982,N_30983,N_30984,N_30985,N_30986,N_30987,N_30988,N_30989,N_30990,N_30991,N_30992,N_30993,N_30994,N_30995,N_30996,N_30997,N_30998,N_30999,N_31000,N_31001,N_31002,N_31003,N_31004,N_31005,N_31006,N_31007,N_31008,N_31009,N_31010,N_31011,N_31012,N_31013,N_31014,N_31015,N_31016,N_31017,N_31018,N_31019,N_31020,N_31021,N_31022,N_31023,N_31024,N_31025,N_31026,N_31027,N_31028,N_31029,N_31030,N_31031,N_31032,N_31033,N_31034,N_31035,N_31036,N_31037,N_31038,N_31039,N_31040,N_31041,N_31042,N_31043,N_31044,N_31045,N_31046,N_31047,N_31048,N_31049,N_31050,N_31051,N_31052,N_31053,N_31054,N_31055,N_31056,N_31057,N_31058,N_31059,N_31060,N_31061,N_31062,N_31063,N_31064,N_31065,N_31066,N_31067,N_31068,N_31069,N_31070,N_31071,N_31072,N_31073,N_31074,N_31075,N_31076,N_31077,N_31078,N_31079,N_31080,N_31081,N_31082,N_31083,N_31084,N_31085,N_31086,N_31087,N_31088,N_31089,N_31090,N_31091,N_31092,N_31093,N_31094,N_31095,N_31096,N_31097,N_31098,N_31099,N_31100,N_31101,N_31102,N_31103,N_31104,N_31105,N_31106,N_31107,N_31108,N_31109,N_31110,N_31111,N_31112,N_31113,N_31114,N_31115,N_31116,N_31117,N_31118,N_31119,N_31120,N_31121,N_31122,N_31123,N_31124,N_31125,N_31126,N_31127,N_31128,N_31129,N_31130,N_31131,N_31132,N_31133,N_31134,N_31135,N_31136,N_31137,N_31138,N_31139,N_31140,N_31141,N_31142,N_31143,N_31144,N_31145,N_31146,N_31147,N_31148,N_31149,N_31150,N_31151,N_31152,N_31153,N_31154,N_31155,N_31156,N_31157,N_31158,N_31159,N_31160,N_31161,N_31162,N_31163,N_31164,N_31165,N_31166,N_31167,N_31168,N_31169,N_31170,N_31171,N_31172,N_31173,N_31174,N_31175,N_31176,N_31177,N_31178,N_31179,N_31180,N_31181,N_31182,N_31183,N_31184,N_31185,N_31186,N_31187,N_31188,N_31189,N_31190,N_31191,N_31192,N_31193,N_31194,N_31195,N_31196,N_31197,N_31198,N_31199,N_31200,N_31201,N_31202,N_31203,N_31204,N_31205,N_31206,N_31207,N_31208,N_31209,N_31210,N_31211,N_31212,N_31213,N_31214,N_31215,N_31216,N_31217,N_31218,N_31219,N_31220,N_31221,N_31222,N_31223,N_31224,N_31225,N_31226,N_31227,N_31228,N_31229,N_31230,N_31231,N_31232,N_31233,N_31234,N_31235,N_31236,N_31237,N_31238,N_31239,N_31240,N_31241,N_31242,N_31243,N_31244,N_31245,N_31246,N_31247,N_31248,N_31249,N_31250,N_31251,N_31252,N_31253,N_31254,N_31255,N_31256,N_31257,N_31258,N_31259,N_31260,N_31261,N_31262,N_31263,N_31264,N_31265,N_31266,N_31267,N_31268,N_31269,N_31270,N_31271,N_31272,N_31273,N_31274,N_31275,N_31276,N_31277,N_31278,N_31279,N_31280,N_31281,N_31282,N_31283,N_31284,N_31285,N_31286,N_31287,N_31288,N_31289,N_31290,N_31291,N_31292,N_31293,N_31294,N_31295,N_31296,N_31297,N_31298,N_31299,N_31300,N_31301,N_31302,N_31303,N_31304,N_31305,N_31306,N_31307,N_31308,N_31309,N_31310,N_31311,N_31312,N_31313,N_31314,N_31315,N_31316,N_31317,N_31318,N_31319,N_31320,N_31321,N_31322,N_31323,N_31324,N_31325,N_31326,N_31327,N_31328,N_31329,N_31330,N_31331,N_31332,N_31333,N_31334,N_31335,N_31336,N_31337,N_31338,N_31339,N_31340,N_31341,N_31342,N_31343,N_31344,N_31345,N_31346,N_31347,N_31348,N_31349,N_31350,N_31351,N_31352,N_31353,N_31354,N_31355,N_31356,N_31357,N_31358,N_31359,N_31360,N_31361,N_31362,N_31363,N_31364,N_31365,N_31366,N_31367,N_31368,N_31369,N_31370,N_31371,N_31372,N_31373,N_31374,N_31375,N_31376,N_31377,N_31378,N_31379,N_31380,N_31381,N_31382,N_31383,N_31384,N_31385,N_31386,N_31387,N_31388,N_31389,N_31390,N_31391,N_31392,N_31393,N_31394,N_31395,N_31396,N_31397,N_31398,N_31399,N_31400,N_31401,N_31402,N_31403,N_31404,N_31405,N_31406,N_31407,N_31408,N_31409,N_31410,N_31411,N_31412,N_31413,N_31414,N_31415,N_31416,N_31417,N_31418,N_31419,N_31420,N_31421,N_31422,N_31423,N_31424,N_31425,N_31426,N_31427,N_31428,N_31429,N_31430,N_31431,N_31432,N_31433,N_31434,N_31435,N_31436,N_31437,N_31438,N_31439,N_31440,N_31441,N_31442,N_31443,N_31444,N_31445,N_31446,N_31447,N_31448,N_31449,N_31450,N_31451,N_31452,N_31453,N_31454,N_31455,N_31456,N_31457,N_31458,N_31459,N_31460,N_31461,N_31462,N_31463,N_31464,N_31465,N_31466,N_31467,N_31468,N_31469,N_31470,N_31471,N_31472,N_31473,N_31474,N_31475,N_31476,N_31477,N_31478,N_31479,N_31480,N_31481,N_31482,N_31483,N_31484,N_31485,N_31486,N_31487,N_31488,N_31489,N_31490,N_31491,N_31492,N_31493,N_31494,N_31495,N_31496,N_31497,N_31498,N_31499,N_31500,N_31501,N_31502,N_31503,N_31504,N_31505,N_31506,N_31507,N_31508,N_31509,N_31510,N_31511,N_31512,N_31513,N_31514,N_31515,N_31516,N_31517,N_31518,N_31519,N_31520,N_31521,N_31522,N_31523,N_31524,N_31525,N_31526,N_31527,N_31528,N_31529,N_31530,N_31531,N_31532,N_31533,N_31534,N_31535,N_31536,N_31537,N_31538,N_31539,N_31540,N_31541,N_31542,N_31543,N_31544,N_31545,N_31546,N_31547,N_31548,N_31549,N_31550,N_31551,N_31552,N_31553,N_31554,N_31555,N_31556,N_31557,N_31558,N_31559,N_31560,N_31561,N_31562,N_31563,N_31564,N_31565,N_31566,N_31567,N_31568,N_31569,N_31570,N_31571,N_31572,N_31573,N_31574,N_31575,N_31576,N_31577,N_31578,N_31579,N_31580,N_31581,N_31582,N_31583,N_31584,N_31585,N_31586,N_31587,N_31588,N_31589,N_31590,N_31591,N_31592,N_31593,N_31594,N_31595,N_31596,N_31597,N_31598,N_31599,N_31600,N_31601,N_31602,N_31603,N_31604,N_31605,N_31606,N_31607,N_31608,N_31609,N_31610,N_31611,N_31612,N_31613,N_31614,N_31615,N_31616,N_31617,N_31618,N_31619,N_31620,N_31621,N_31622,N_31623,N_31624,N_31625,N_31626,N_31627,N_31628,N_31629,N_31630,N_31631,N_31632,N_31633,N_31634,N_31635,N_31636,N_31637,N_31638,N_31639,N_31640,N_31641,N_31642,N_31643,N_31644,N_31645,N_31646,N_31647,N_31648,N_31649,N_31650,N_31651,N_31652,N_31653,N_31654,N_31655,N_31656,N_31657,N_31658,N_31659,N_31660,N_31661,N_31662,N_31663,N_31664,N_31665,N_31666,N_31667,N_31668,N_31669,N_31670,N_31671,N_31672,N_31673,N_31674,N_31675,N_31676,N_31677,N_31678,N_31679,N_31680,N_31681,N_31682,N_31683,N_31684,N_31685,N_31686,N_31687,N_31688,N_31689,N_31690,N_31691,N_31692,N_31693,N_31694,N_31695,N_31696,N_31697,N_31698,N_31699,N_31700,N_31701,N_31702,N_31703,N_31704,N_31705,N_31706,N_31707,N_31708,N_31709,N_31710,N_31711,N_31712,N_31713,N_31714,N_31715,N_31716,N_31717,N_31718,N_31719,N_31720,N_31721,N_31722,N_31723,N_31724,N_31725,N_31726,N_31727,N_31728,N_31729,N_31730,N_31731,N_31732,N_31733,N_31734,N_31735,N_31736,N_31737,N_31738,N_31739,N_31740,N_31741,N_31742,N_31743,N_31744,N_31745,N_31746,N_31747,N_31748,N_31749,N_31750,N_31751,N_31752,N_31753,N_31754,N_31755,N_31756,N_31757,N_31758,N_31759,N_31760,N_31761,N_31762,N_31763,N_31764,N_31765,N_31766,N_31767,N_31768,N_31769,N_31770,N_31771,N_31772,N_31773,N_31774,N_31775,N_31776,N_31777,N_31778,N_31779,N_31780,N_31781,N_31782,N_31783,N_31784,N_31785,N_31786,N_31787,N_31788,N_31789,N_31790,N_31791,N_31792,N_31793,N_31794,N_31795,N_31796,N_31797,N_31798,N_31799,N_31800,N_31801,N_31802,N_31803,N_31804,N_31805,N_31806,N_31807,N_31808,N_31809,N_31810,N_31811,N_31812,N_31813,N_31814,N_31815,N_31816,N_31817,N_31818,N_31819,N_31820,N_31821,N_31822,N_31823,N_31824,N_31825,N_31826,N_31827,N_31828,N_31829,N_31830,N_31831,N_31832,N_31833,N_31834,N_31835,N_31836,N_31837,N_31838,N_31839,N_31840,N_31841,N_31842,N_31843,N_31844,N_31845,N_31846,N_31847,N_31848,N_31849,N_31850,N_31851,N_31852,N_31853,N_31854,N_31855,N_31856,N_31857,N_31858,N_31859,N_31860,N_31861,N_31862,N_31863,N_31864,N_31865,N_31866,N_31867,N_31868,N_31869,N_31870,N_31871,N_31872,N_31873,N_31874,N_31875,N_31876,N_31877,N_31878,N_31879,N_31880,N_31881,N_31882,N_31883,N_31884,N_31885,N_31886,N_31887,N_31888,N_31889,N_31890,N_31891,N_31892,N_31893,N_31894,N_31895,N_31896,N_31897,N_31898,N_31899,N_31900,N_31901,N_31902,N_31903,N_31904,N_31905,N_31906,N_31907,N_31908,N_31909,N_31910,N_31911,N_31912,N_31913,N_31914,N_31915,N_31916,N_31917,N_31918,N_31919,N_31920,N_31921,N_31922,N_31923,N_31924,N_31925,N_31926,N_31927,N_31928,N_31929,N_31930,N_31931,N_31932,N_31933,N_31934,N_31935,N_31936,N_31937,N_31938,N_31939,N_31940,N_31941,N_31942,N_31943,N_31944,N_31945,N_31946,N_31947,N_31948,N_31949,N_31950,N_31951,N_31952,N_31953,N_31954,N_31955,N_31956,N_31957,N_31958,N_31959,N_31960,N_31961,N_31962,N_31963,N_31964,N_31965,N_31966,N_31967,N_31968,N_31969,N_31970,N_31971,N_31972,N_31973,N_31974,N_31975,N_31976,N_31977,N_31978,N_31979,N_31980,N_31981,N_31982,N_31983,N_31984,N_31985,N_31986,N_31987,N_31988,N_31989,N_31990,N_31991,N_31992,N_31993,N_31994,N_31995,N_31996,N_31997,N_31998,N_31999,N_32000,N_32001,N_32002,N_32003,N_32004,N_32005,N_32006,N_32007,N_32008,N_32009,N_32010,N_32011,N_32012,N_32013,N_32014,N_32015,N_32016,N_32017,N_32018,N_32019,N_32020,N_32021,N_32022,N_32023,N_32024,N_32025,N_32026,N_32027,N_32028,N_32029,N_32030,N_32031,N_32032,N_32033,N_32034,N_32035,N_32036,N_32037,N_32038,N_32039,N_32040,N_32041,N_32042,N_32043,N_32044,N_32045,N_32046,N_32047,N_32048,N_32049,N_32050,N_32051,N_32052,N_32053,N_32054,N_32055,N_32056,N_32057,N_32058,N_32059,N_32060,N_32061,N_32062,N_32063,N_32064,N_32065,N_32066,N_32067,N_32068,N_32069,N_32070,N_32071,N_32072,N_32073,N_32074,N_32075,N_32076,N_32077,N_32078,N_32079,N_32080,N_32081,N_32082,N_32083,N_32084,N_32085,N_32086,N_32087,N_32088,N_32089,N_32090,N_32091,N_32092,N_32093,N_32094,N_32095,N_32096,N_32097,N_32098,N_32099,N_32100,N_32101,N_32102,N_32103,N_32104,N_32105,N_32106,N_32107,N_32108,N_32109,N_32110,N_32111,N_32112,N_32113,N_32114,N_32115,N_32116,N_32117,N_32118,N_32119,N_32120,N_32121,N_32122,N_32123,N_32124,N_32125,N_32126,N_32127,N_32128,N_32129,N_32130,N_32131,N_32132,N_32133,N_32134,N_32135,N_32136,N_32137,N_32138,N_32139,N_32140,N_32141,N_32142,N_32143,N_32144,N_32145,N_32146,N_32147,N_32148,N_32149,N_32150,N_32151,N_32152,N_32153,N_32154,N_32155,N_32156,N_32157,N_32158,N_32159,N_32160,N_32161,N_32162,N_32163,N_32164,N_32165,N_32166,N_32167,N_32168,N_32169,N_32170,N_32171,N_32172,N_32173,N_32174,N_32175,N_32176,N_32177,N_32178,N_32179,N_32180,N_32181,N_32182,N_32183,N_32184,N_32185,N_32186,N_32187,N_32188,N_32189,N_32190,N_32191,N_32192,N_32193,N_32194,N_32195,N_32196,N_32197,N_32198,N_32199,N_32200,N_32201,N_32202,N_32203,N_32204,N_32205,N_32206,N_32207,N_32208,N_32209,N_32210,N_32211,N_32212,N_32213,N_32214,N_32215,N_32216,N_32217,N_32218,N_32219,N_32220,N_32221,N_32222,N_32223,N_32224,N_32225,N_32226,N_32227,N_32228,N_32229,N_32230,N_32231,N_32232,N_32233,N_32234,N_32235,N_32236,N_32237,N_32238,N_32239,N_32240,N_32241,N_32242,N_32243,N_32244,N_32245,N_32246,N_32247,N_32248,N_32249,N_32250,N_32251,N_32252,N_32253,N_32254,N_32255,N_32256,N_32257,N_32258,N_32259,N_32260,N_32261,N_32262,N_32263,N_32264,N_32265,N_32266,N_32267,N_32268,N_32269,N_32270,N_32271,N_32272,N_32273,N_32274,N_32275,N_32276,N_32277,N_32278,N_32279,N_32280,N_32281,N_32282,N_32283,N_32284,N_32285,N_32286,N_32287,N_32288,N_32289,N_32290,N_32291,N_32292,N_32293,N_32294,N_32295,N_32296,N_32297,N_32298,N_32299,N_32300,N_32301,N_32302,N_32303,N_32304,N_32305,N_32306,N_32307,N_32308,N_32309,N_32310,N_32311,N_32312,N_32313,N_32314,N_32315,N_32316,N_32317,N_32318,N_32319,N_32320,N_32321,N_32322,N_32323,N_32324,N_32325,N_32326,N_32327,N_32328,N_32329,N_32330,N_32331,N_32332,N_32333,N_32334,N_32335,N_32336,N_32337,N_32338,N_32339,N_32340,N_32341,N_32342,N_32343,N_32344,N_32345,N_32346,N_32347,N_32348,N_32349,N_32350,N_32351,N_32352,N_32353,N_32354,N_32355,N_32356,N_32357,N_32358,N_32359,N_32360,N_32361,N_32362,N_32363,N_32364,N_32365,N_32366,N_32367,N_32368,N_32369,N_32370,N_32371,N_32372,N_32373,N_32374,N_32375,N_32376,N_32377,N_32378,N_32379,N_32380,N_32381,N_32382,N_32383,N_32384,N_32385,N_32386,N_32387,N_32388,N_32389,N_32390,N_32391,N_32392,N_32393,N_32394,N_32395,N_32396,N_32397,N_32398,N_32399,N_32400,N_32401,N_32402,N_32403,N_32404,N_32405,N_32406,N_32407,N_32408,N_32409,N_32410,N_32411,N_32412,N_32413,N_32414,N_32415,N_32416,N_32417,N_32418,N_32419,N_32420,N_32421,N_32422,N_32423,N_32424,N_32425,N_32426,N_32427,N_32428,N_32429,N_32430,N_32431,N_32432,N_32433,N_32434,N_32435,N_32436,N_32437,N_32438,N_32439,N_32440,N_32441,N_32442,N_32443,N_32444,N_32445,N_32446,N_32447,N_32448,N_32449,N_32450,N_32451,N_32452,N_32453,N_32454,N_32455,N_32456,N_32457,N_32458,N_32459,N_32460,N_32461,N_32462,N_32463,N_32464,N_32465,N_32466,N_32467,N_32468,N_32469,N_32470,N_32471,N_32472,N_32473,N_32474,N_32475,N_32476,N_32477,N_32478,N_32479,N_32480,N_32481,N_32482,N_32483,N_32484,N_32485,N_32486,N_32487,N_32488,N_32489,N_32490,N_32491,N_32492,N_32493,N_32494,N_32495,N_32496,N_32497,N_32498,N_32499,N_32500,N_32501,N_32502,N_32503,N_32504,N_32505,N_32506,N_32507,N_32508,N_32509,N_32510,N_32511,N_32512,N_32513,N_32514,N_32515,N_32516,N_32517,N_32518,N_32519,N_32520,N_32521,N_32522,N_32523,N_32524,N_32525,N_32526,N_32527,N_32528,N_32529,N_32530,N_32531,N_32532,N_32533,N_32534,N_32535,N_32536,N_32537,N_32538,N_32539,N_32540,N_32541,N_32542,N_32543,N_32544,N_32545,N_32546,N_32547,N_32548,N_32549,N_32550,N_32551,N_32552,N_32553,N_32554,N_32555,N_32556,N_32557,N_32558,N_32559,N_32560,N_32561,N_32562,N_32563,N_32564,N_32565,N_32566,N_32567,N_32568,N_32569,N_32570,N_32571,N_32572,N_32573,N_32574,N_32575,N_32576,N_32577,N_32578,N_32579,N_32580,N_32581,N_32582,N_32583,N_32584,N_32585,N_32586,N_32587,N_32588,N_32589,N_32590,N_32591,N_32592,N_32593,N_32594,N_32595,N_32596,N_32597,N_32598,N_32599,N_32600,N_32601,N_32602,N_32603,N_32604,N_32605,N_32606,N_32607,N_32608,N_32609,N_32610,N_32611,N_32612,N_32613,N_32614,N_32615,N_32616,N_32617,N_32618,N_32619,N_32620,N_32621,N_32622,N_32623,N_32624,N_32625,N_32626,N_32627,N_32628,N_32629,N_32630,N_32631,N_32632,N_32633,N_32634,N_32635,N_32636,N_32637,N_32638,N_32639,N_32640,N_32641,N_32642,N_32643,N_32644,N_32645,N_32646,N_32647,N_32648,N_32649,N_32650,N_32651,N_32652,N_32653,N_32654,N_32655,N_32656,N_32657,N_32658,N_32659,N_32660,N_32661,N_32662,N_32663,N_32664,N_32665,N_32666,N_32667,N_32668,N_32669,N_32670,N_32671,N_32672,N_32673,N_32674,N_32675,N_32676,N_32677,N_32678,N_32679,N_32680,N_32681,N_32682,N_32683,N_32684,N_32685,N_32686,N_32687,N_32688,N_32689,N_32690,N_32691,N_32692,N_32693,N_32694,N_32695,N_32696,N_32697,N_32698,N_32699,N_32700,N_32701,N_32702,N_32703,N_32704,N_32705,N_32706,N_32707,N_32708,N_32709,N_32710,N_32711,N_32712,N_32713,N_32714,N_32715,N_32716,N_32717,N_32718,N_32719,N_32720,N_32721,N_32722,N_32723,N_32724,N_32725,N_32726,N_32727,N_32728,N_32729,N_32730,N_32731,N_32732,N_32733,N_32734,N_32735,N_32736,N_32737,N_32738,N_32739,N_32740,N_32741,N_32742,N_32743,N_32744,N_32745,N_32746,N_32747,N_32748,N_32749,N_32750,N_32751,N_32752,N_32753,N_32754,N_32755,N_32756,N_32757,N_32758,N_32759,N_32760,N_32761,N_32762,N_32763,N_32764,N_32765,N_32766,N_32767,N_32768,N_32769,N_32770,N_32771,N_32772,N_32773,N_32774,N_32775,N_32776,N_32777,N_32778,N_32779,N_32780,N_32781,N_32782,N_32783,N_32784,N_32785,N_32786,N_32787,N_32788,N_32789,N_32790,N_32791,N_32792,N_32793,N_32794,N_32795,N_32796,N_32797,N_32798,N_32799,N_32800,N_32801,N_32802,N_32803,N_32804,N_32805,N_32806,N_32807,N_32808,N_32809,N_32810,N_32811,N_32812,N_32813,N_32814,N_32815,N_32816,N_32817,N_32818,N_32819,N_32820,N_32821,N_32822,N_32823,N_32824,N_32825,N_32826,N_32827,N_32828,N_32829,N_32830,N_32831,N_32832,N_32833,N_32834,N_32835,N_32836,N_32837,N_32838,N_32839,N_32840,N_32841,N_32842,N_32843,N_32844,N_32845,N_32846,N_32847,N_32848,N_32849,N_32850,N_32851,N_32852,N_32853,N_32854,N_32855,N_32856,N_32857,N_32858,N_32859,N_32860,N_32861,N_32862,N_32863,N_32864,N_32865,N_32866,N_32867,N_32868,N_32869,N_32870,N_32871,N_32872,N_32873,N_32874,N_32875,N_32876,N_32877,N_32878,N_32879,N_32880,N_32881,N_32882,N_32883,N_32884,N_32885,N_32886,N_32887,N_32888,N_32889,N_32890,N_32891,N_32892,N_32893,N_32894,N_32895,N_32896,N_32897,N_32898,N_32899,N_32900,N_32901,N_32902,N_32903,N_32904,N_32905,N_32906,N_32907,N_32908,N_32909,N_32910,N_32911,N_32912,N_32913,N_32914,N_32915,N_32916,N_32917,N_32918,N_32919,N_32920,N_32921,N_32922,N_32923,N_32924,N_32925,N_32926,N_32927,N_32928,N_32929,N_32930,N_32931,N_32932,N_32933,N_32934,N_32935,N_32936,N_32937,N_32938,N_32939,N_32940,N_32941,N_32942,N_32943,N_32944,N_32945,N_32946,N_32947,N_32948,N_32949,N_32950,N_32951,N_32952,N_32953,N_32954,N_32955,N_32956,N_32957,N_32958,N_32959,N_32960,N_32961,N_32962,N_32963,N_32964,N_32965,N_32966,N_32967,N_32968,N_32969,N_32970,N_32971,N_32972,N_32973,N_32974,N_32975,N_32976,N_32977,N_32978,N_32979,N_32980,N_32981,N_32982,N_32983,N_32984,N_32985,N_32986,N_32987,N_32988,N_32989,N_32990,N_32991,N_32992,N_32993,N_32994,N_32995,N_32996,N_32997,N_32998,N_32999,N_33000,N_33001,N_33002,N_33003,N_33004,N_33005,N_33006,N_33007,N_33008,N_33009,N_33010,N_33011,N_33012,N_33013,N_33014,N_33015,N_33016,N_33017,N_33018,N_33019,N_33020,N_33021,N_33022,N_33023,N_33024,N_33025,N_33026,N_33027,N_33028,N_33029,N_33030,N_33031,N_33032,N_33033,N_33034,N_33035,N_33036,N_33037,N_33038,N_33039,N_33040,N_33041,N_33042,N_33043,N_33044,N_33045,N_33046,N_33047,N_33048,N_33049,N_33050,N_33051,N_33052,N_33053,N_33054,N_33055,N_33056,N_33057,N_33058,N_33059,N_33060,N_33061,N_33062,N_33063,N_33064,N_33065,N_33066,N_33067,N_33068,N_33069,N_33070,N_33071,N_33072,N_33073,N_33074,N_33075,N_33076,N_33077,N_33078,N_33079,N_33080,N_33081,N_33082,N_33083,N_33084,N_33085,N_33086,N_33087,N_33088,N_33089,N_33090,N_33091,N_33092,N_33093,N_33094,N_33095,N_33096,N_33097,N_33098,N_33099,N_33100,N_33101,N_33102,N_33103,N_33104,N_33105,N_33106,N_33107,N_33108,N_33109,N_33110,N_33111,N_33112,N_33113,N_33114,N_33115,N_33116,N_33117,N_33118,N_33119,N_33120,N_33121,N_33122,N_33123,N_33124,N_33125,N_33126,N_33127,N_33128,N_33129,N_33130,N_33131,N_33132,N_33133,N_33134,N_33135,N_33136,N_33137,N_33138,N_33139,N_33140,N_33141,N_33142,N_33143,N_33144,N_33145,N_33146,N_33147,N_33148,N_33149,N_33150,N_33151,N_33152,N_33153,N_33154,N_33155,N_33156,N_33157,N_33158,N_33159,N_33160,N_33161,N_33162,N_33163,N_33164,N_33165,N_33166,N_33167,N_33168,N_33169,N_33170,N_33171,N_33172,N_33173,N_33174,N_33175,N_33176,N_33177,N_33178,N_33179,N_33180,N_33181,N_33182,N_33183,N_33184,N_33185,N_33186,N_33187,N_33188,N_33189,N_33190,N_33191,N_33192,N_33193,N_33194,N_33195,N_33196,N_33197,N_33198,N_33199,N_33200,N_33201,N_33202,N_33203,N_33204,N_33205,N_33206,N_33207,N_33208,N_33209,N_33210,N_33211,N_33212,N_33213,N_33214,N_33215,N_33216,N_33217,N_33218,N_33219,N_33220,N_33221,N_33222,N_33223,N_33224,N_33225,N_33226,N_33227,N_33228,N_33229,N_33230,N_33231,N_33232,N_33233,N_33234,N_33235,N_33236,N_33237,N_33238,N_33239,N_33240,N_33241,N_33242,N_33243,N_33244,N_33245,N_33246,N_33247,N_33248,N_33249,N_33250,N_33251,N_33252,N_33253,N_33254,N_33255,N_33256,N_33257,N_33258,N_33259,N_33260,N_33261,N_33262,N_33263,N_33264,N_33265,N_33266,N_33267,N_33268,N_33269,N_33270,N_33271,N_33272,N_33273,N_33274,N_33275,N_33276,N_33277,N_33278,N_33279,N_33280,N_33281,N_33282,N_33283,N_33284,N_33285,N_33286,N_33287,N_33288,N_33289,N_33290,N_33291,N_33292,N_33293,N_33294,N_33295,N_33296,N_33297,N_33298,N_33299,N_33300,N_33301,N_33302,N_33303,N_33304,N_33305,N_33306,N_33307,N_33308,N_33309,N_33310,N_33311,N_33312,N_33313,N_33314,N_33315,N_33316,N_33317,N_33318,N_33319,N_33320,N_33321,N_33322,N_33323,N_33324,N_33325,N_33326,N_33327,N_33328,N_33329,N_33330,N_33331,N_33332,N_33333,N_33334,N_33335,N_33336,N_33337,N_33338,N_33339,N_33340,N_33341,N_33342,N_33343,N_33344,N_33345,N_33346,N_33347,N_33348,N_33349,N_33350,N_33351,N_33352,N_33353,N_33354,N_33355,N_33356,N_33357,N_33358,N_33359,N_33360,N_33361,N_33362,N_33363,N_33364,N_33365,N_33366,N_33367,N_33368,N_33369,N_33370,N_33371,N_33372,N_33373,N_33374,N_33375,N_33376,N_33377,N_33378,N_33379,N_33380,N_33381,N_33382,N_33383,N_33384,N_33385,N_33386,N_33387,N_33388,N_33389,N_33390,N_33391,N_33392,N_33393,N_33394,N_33395,N_33396,N_33397,N_33398,N_33399,N_33400,N_33401,N_33402,N_33403,N_33404,N_33405,N_33406,N_33407,N_33408,N_33409,N_33410,N_33411,N_33412,N_33413,N_33414,N_33415,N_33416,N_33417,N_33418,N_33419,N_33420,N_33421,N_33422,N_33423,N_33424,N_33425,N_33426,N_33427,N_33428,N_33429,N_33430,N_33431,N_33432,N_33433,N_33434,N_33435,N_33436,N_33437,N_33438,N_33439,N_33440,N_33441,N_33442,N_33443,N_33444,N_33445,N_33446,N_33447,N_33448,N_33449,N_33450,N_33451,N_33452,N_33453,N_33454,N_33455,N_33456,N_33457,N_33458,N_33459,N_33460,N_33461,N_33462,N_33463,N_33464,N_33465,N_33466,N_33467,N_33468,N_33469,N_33470,N_33471,N_33472,N_33473,N_33474,N_33475,N_33476,N_33477,N_33478,N_33479,N_33480,N_33481,N_33482,N_33483,N_33484,N_33485,N_33486,N_33487,N_33488,N_33489,N_33490,N_33491,N_33492,N_33493,N_33494,N_33495,N_33496,N_33497,N_33498,N_33499,N_33500,N_33501,N_33502,N_33503,N_33504,N_33505,N_33506,N_33507,N_33508,N_33509,N_33510,N_33511,N_33512,N_33513,N_33514,N_33515,N_33516,N_33517,N_33518,N_33519,N_33520,N_33521,N_33522,N_33523,N_33524,N_33525,N_33526,N_33527,N_33528,N_33529,N_33530,N_33531,N_33532,N_33533,N_33534,N_33535,N_33536,N_33537,N_33538,N_33539,N_33540,N_33541,N_33542,N_33543,N_33544,N_33545,N_33546,N_33547,N_33548,N_33549,N_33550,N_33551,N_33552,N_33553,N_33554,N_33555,N_33556,N_33557,N_33558,N_33559,N_33560,N_33561,N_33562,N_33563,N_33564,N_33565,N_33566,N_33567,N_33568,N_33569,N_33570,N_33571,N_33572,N_33573,N_33574,N_33575,N_33576,N_33577,N_33578,N_33579,N_33580,N_33581,N_33582,N_33583,N_33584,N_33585,N_33586,N_33587,N_33588,N_33589,N_33590,N_33591,N_33592,N_33593,N_33594,N_33595,N_33596,N_33597,N_33598,N_33599,N_33600,N_33601,N_33602,N_33603,N_33604,N_33605,N_33606,N_33607,N_33608,N_33609,N_33610,N_33611,N_33612,N_33613,N_33614,N_33615,N_33616,N_33617,N_33618,N_33619,N_33620,N_33621,N_33622,N_33623,N_33624,N_33625,N_33626,N_33627,N_33628,N_33629,N_33630,N_33631,N_33632,N_33633,N_33634,N_33635,N_33636,N_33637,N_33638,N_33639,N_33640,N_33641,N_33642,N_33643,N_33644,N_33645,N_33646,N_33647,N_33648,N_33649,N_33650,N_33651,N_33652,N_33653,N_33654,N_33655,N_33656,N_33657,N_33658,N_33659,N_33660,N_33661,N_33662,N_33663,N_33664,N_33665,N_33666,N_33667,N_33668,N_33669,N_33670,N_33671,N_33672,N_33673,N_33674,N_33675,N_33676,N_33677,N_33678,N_33679,N_33680,N_33681,N_33682,N_33683,N_33684,N_33685,N_33686,N_33687,N_33688,N_33689,N_33690,N_33691,N_33692,N_33693,N_33694,N_33695,N_33696,N_33697,N_33698,N_33699,N_33700,N_33701,N_33702,N_33703,N_33704,N_33705,N_33706,N_33707,N_33708,N_33709,N_33710,N_33711,N_33712,N_33713,N_33714,N_33715,N_33716,N_33717,N_33718,N_33719,N_33720,N_33721,N_33722,N_33723,N_33724,N_33725,N_33726,N_33727,N_33728,N_33729,N_33730,N_33731,N_33732,N_33733,N_33734,N_33735,N_33736,N_33737,N_33738,N_33739,N_33740,N_33741,N_33742,N_33743,N_33744,N_33745,N_33746,N_33747,N_33748,N_33749,N_33750,N_33751,N_33752,N_33753,N_33754,N_33755,N_33756,N_33757,N_33758,N_33759,N_33760,N_33761,N_33762,N_33763,N_33764,N_33765,N_33766,N_33767,N_33768,N_33769,N_33770,N_33771,N_33772,N_33773,N_33774,N_33775,N_33776,N_33777,N_33778,N_33779,N_33780,N_33781,N_33782,N_33783,N_33784,N_33785,N_33786,N_33787,N_33788,N_33789,N_33790,N_33791,N_33792,N_33793,N_33794,N_33795,N_33796,N_33797,N_33798,N_33799,N_33800,N_33801,N_33802,N_33803,N_33804,N_33805,N_33806,N_33807,N_33808,N_33809,N_33810,N_33811,N_33812,N_33813,N_33814,N_33815,N_33816,N_33817,N_33818,N_33819,N_33820,N_33821,N_33822,N_33823,N_33824,N_33825,N_33826,N_33827,N_33828,N_33829,N_33830,N_33831,N_33832,N_33833,N_33834,N_33835,N_33836,N_33837,N_33838,N_33839,N_33840,N_33841,N_33842,N_33843,N_33844,N_33845,N_33846,N_33847,N_33848,N_33849,N_33850,N_33851,N_33852,N_33853,N_33854,N_33855,N_33856,N_33857,N_33858,N_33859,N_33860,N_33861,N_33862,N_33863,N_33864,N_33865,N_33866,N_33867,N_33868,N_33869,N_33870,N_33871,N_33872,N_33873,N_33874,N_33875,N_33876,N_33877,N_33878,N_33879,N_33880,N_33881,N_33882,N_33883,N_33884,N_33885,N_33886,N_33887,N_33888,N_33889,N_33890,N_33891,N_33892,N_33893,N_33894,N_33895,N_33896,N_33897,N_33898,N_33899,N_33900,N_33901,N_33902,N_33903,N_33904,N_33905,N_33906,N_33907,N_33908,N_33909,N_33910,N_33911,N_33912,N_33913,N_33914,N_33915,N_33916,N_33917,N_33918,N_33919,N_33920,N_33921,N_33922,N_33923,N_33924,N_33925,N_33926,N_33927,N_33928,N_33929,N_33930,N_33931,N_33932,N_33933,N_33934,N_33935,N_33936,N_33937,N_33938,N_33939,N_33940,N_33941,N_33942,N_33943,N_33944,N_33945,N_33946,N_33947,N_33948,N_33949,N_33950,N_33951,N_33952,N_33953,N_33954,N_33955,N_33956,N_33957,N_33958,N_33959,N_33960,N_33961,N_33962,N_33963,N_33964,N_33965,N_33966,N_33967,N_33968,N_33969,N_33970,N_33971,N_33972,N_33973,N_33974,N_33975,N_33976,N_33977,N_33978,N_33979,N_33980,N_33981,N_33982,N_33983,N_33984,N_33985,N_33986,N_33987,N_33988,N_33989,N_33990,N_33991,N_33992,N_33993,N_33994,N_33995,N_33996,N_33997,N_33998,N_33999,N_34000,N_34001,N_34002,N_34003,N_34004,N_34005,N_34006,N_34007,N_34008,N_34009,N_34010,N_34011,N_34012,N_34013,N_34014,N_34015,N_34016,N_34017,N_34018,N_34019,N_34020,N_34021,N_34022,N_34023,N_34024,N_34025,N_34026,N_34027,N_34028,N_34029,N_34030,N_34031,N_34032,N_34033,N_34034,N_34035,N_34036,N_34037,N_34038,N_34039,N_34040,N_34041,N_34042,N_34043,N_34044,N_34045,N_34046,N_34047,N_34048,N_34049,N_34050,N_34051,N_34052,N_34053,N_34054,N_34055,N_34056,N_34057,N_34058,N_34059,N_34060,N_34061,N_34062,N_34063,N_34064,N_34065,N_34066,N_34067,N_34068,N_34069,N_34070,N_34071,N_34072,N_34073,N_34074,N_34075,N_34076,N_34077,N_34078,N_34079,N_34080,N_34081,N_34082,N_34083,N_34084,N_34085,N_34086,N_34087,N_34088,N_34089,N_34090,N_34091,N_34092,N_34093,N_34094,N_34095,N_34096,N_34097,N_34098,N_34099,N_34100,N_34101,N_34102,N_34103,N_34104,N_34105,N_34106,N_34107,N_34108,N_34109,N_34110,N_34111,N_34112,N_34113,N_34114,N_34115,N_34116,N_34117,N_34118,N_34119,N_34120,N_34121,N_34122,N_34123,N_34124,N_34125,N_34126,N_34127,N_34128,N_34129,N_34130,N_34131,N_34132,N_34133,N_34134,N_34135,N_34136,N_34137,N_34138,N_34139,N_34140,N_34141,N_34142,N_34143,N_34144,N_34145,N_34146,N_34147,N_34148,N_34149,N_34150,N_34151,N_34152,N_34153,N_34154,N_34155,N_34156,N_34157,N_34158,N_34159,N_34160,N_34161,N_34162,N_34163,N_34164,N_34165,N_34166,N_34167,N_34168,N_34169,N_34170,N_34171,N_34172,N_34173,N_34174,N_34175,N_34176,N_34177,N_34178,N_34179,N_34180,N_34181,N_34182,N_34183,N_34184,N_34185,N_34186,N_34187,N_34188,N_34189,N_34190,N_34191,N_34192,N_34193,N_34194,N_34195,N_34196,N_34197,N_34198,N_34199,N_34200,N_34201,N_34202,N_34203,N_34204,N_34205,N_34206,N_34207,N_34208,N_34209,N_34210,N_34211,N_34212,N_34213,N_34214,N_34215,N_34216,N_34217,N_34218,N_34219,N_34220,N_34221,N_34222,N_34223,N_34224,N_34225,N_34226,N_34227,N_34228,N_34229,N_34230,N_34231,N_34232,N_34233,N_34234,N_34235,N_34236,N_34237,N_34238,N_34239,N_34240,N_34241,N_34242,N_34243,N_34244,N_34245,N_34246,N_34247,N_34248,N_34249,N_34250,N_34251,N_34252,N_34253,N_34254,N_34255,N_34256,N_34257,N_34258,N_34259,N_34260,N_34261,N_34262,N_34263,N_34264,N_34265,N_34266,N_34267,N_34268,N_34269,N_34270,N_34271,N_34272,N_34273,N_34274,N_34275,N_34276,N_34277,N_34278,N_34279,N_34280,N_34281,N_34282,N_34283,N_34284,N_34285,N_34286,N_34287,N_34288,N_34289,N_34290,N_34291,N_34292,N_34293,N_34294,N_34295,N_34296,N_34297,N_34298,N_34299,N_34300,N_34301,N_34302,N_34303,N_34304,N_34305,N_34306,N_34307,N_34308,N_34309,N_34310,N_34311,N_34312,N_34313,N_34314,N_34315,N_34316,N_34317,N_34318,N_34319,N_34320,N_34321,N_34322,N_34323,N_34324,N_34325,N_34326,N_34327,N_34328,N_34329,N_34330,N_34331,N_34332,N_34333,N_34334,N_34335,N_34336,N_34337,N_34338,N_34339,N_34340,N_34341,N_34342,N_34343,N_34344,N_34345,N_34346,N_34347,N_34348,N_34349,N_34350,N_34351,N_34352,N_34353,N_34354,N_34355,N_34356,N_34357,N_34358,N_34359,N_34360,N_34361,N_34362,N_34363,N_34364,N_34365,N_34366,N_34367,N_34368,N_34369,N_34370,N_34371,N_34372,N_34373,N_34374,N_34375,N_34376,N_34377,N_34378,N_34379,N_34380,N_34381,N_34382,N_34383,N_34384,N_34385,N_34386,N_34387,N_34388,N_34389,N_34390,N_34391,N_34392,N_34393,N_34394,N_34395,N_34396,N_34397,N_34398,N_34399,N_34400,N_34401,N_34402,N_34403,N_34404,N_34405,N_34406,N_34407,N_34408,N_34409,N_34410,N_34411,N_34412,N_34413,N_34414,N_34415,N_34416,N_34417,N_34418,N_34419,N_34420,N_34421,N_34422,N_34423,N_34424,N_34425,N_34426,N_34427,N_34428,N_34429,N_34430,N_34431,N_34432,N_34433,N_34434,N_34435,N_34436,N_34437,N_34438,N_34439,N_34440,N_34441,N_34442,N_34443,N_34444,N_34445,N_34446,N_34447,N_34448,N_34449,N_34450,N_34451,N_34452,N_34453,N_34454,N_34455,N_34456,N_34457,N_34458,N_34459,N_34460,N_34461,N_34462,N_34463,N_34464,N_34465,N_34466,N_34467,N_34468,N_34469,N_34470,N_34471,N_34472,N_34473,N_34474,N_34475,N_34476,N_34477,N_34478,N_34479,N_34480,N_34481,N_34482,N_34483,N_34484,N_34485,N_34486,N_34487,N_34488,N_34489,N_34490,N_34491,N_34492,N_34493,N_34494,N_34495,N_34496,N_34497,N_34498,N_34499,N_34500,N_34501,N_34502,N_34503,N_34504,N_34505,N_34506,N_34507,N_34508,N_34509,N_34510,N_34511,N_34512,N_34513,N_34514,N_34515,N_34516,N_34517,N_34518,N_34519,N_34520,N_34521,N_34522,N_34523,N_34524,N_34525,N_34526,N_34527,N_34528,N_34529,N_34530,N_34531,N_34532,N_34533,N_34534,N_34535,N_34536,N_34537,N_34538,N_34539,N_34540,N_34541,N_34542,N_34543,N_34544,N_34545,N_34546,N_34547,N_34548,N_34549,N_34550,N_34551,N_34552,N_34553,N_34554,N_34555,N_34556,N_34557,N_34558,N_34559,N_34560,N_34561,N_34562,N_34563,N_34564,N_34565,N_34566,N_34567,N_34568,N_34569,N_34570,N_34571,N_34572,N_34573,N_34574,N_34575,N_34576,N_34577,N_34578,N_34579,N_34580,N_34581,N_34582,N_34583,N_34584,N_34585,N_34586,N_34587,N_34588,N_34589,N_34590,N_34591,N_34592,N_34593,N_34594,N_34595,N_34596,N_34597,N_34598,N_34599,N_34600,N_34601,N_34602,N_34603,N_34604,N_34605,N_34606,N_34607,N_34608,N_34609,N_34610,N_34611,N_34612,N_34613,N_34614,N_34615,N_34616,N_34617,N_34618,N_34619,N_34620,N_34621,N_34622,N_34623,N_34624,N_34625,N_34626,N_34627,N_34628,N_34629,N_34630,N_34631,N_34632,N_34633,N_34634,N_34635,N_34636,N_34637,N_34638,N_34639,N_34640,N_34641,N_34642,N_34643,N_34644,N_34645,N_34646,N_34647,N_34648,N_34649,N_34650,N_34651,N_34652,N_34653,N_34654,N_34655,N_34656,N_34657,N_34658,N_34659,N_34660,N_34661,N_34662,N_34663,N_34664,N_34665,N_34666,N_34667,N_34668,N_34669,N_34670,N_34671,N_34672,N_34673,N_34674,N_34675,N_34676,N_34677,N_34678,N_34679,N_34680,N_34681,N_34682,N_34683,N_34684,N_34685,N_34686,N_34687,N_34688,N_34689,N_34690,N_34691,N_34692,N_34693,N_34694,N_34695,N_34696,N_34697,N_34698,N_34699,N_34700,N_34701,N_34702,N_34703,N_34704,N_34705,N_34706,N_34707,N_34708,N_34709,N_34710,N_34711,N_34712,N_34713,N_34714,N_34715,N_34716,N_34717,N_34718,N_34719,N_34720,N_34721,N_34722,N_34723,N_34724,N_34725,N_34726,N_34727,N_34728,N_34729,N_34730,N_34731,N_34732,N_34733,N_34734,N_34735,N_34736,N_34737,N_34738,N_34739,N_34740,N_34741,N_34742,N_34743,N_34744,N_34745,N_34746,N_34747,N_34748,N_34749,N_34750,N_34751,N_34752,N_34753,N_34754,N_34755,N_34756,N_34757,N_34758,N_34759,N_34760,N_34761,N_34762,N_34763,N_34764,N_34765,N_34766,N_34767,N_34768,N_34769,N_34770,N_34771,N_34772,N_34773,N_34774,N_34775,N_34776,N_34777,N_34778,N_34779,N_34780,N_34781,N_34782,N_34783,N_34784,N_34785,N_34786,N_34787,N_34788,N_34789,N_34790,N_34791,N_34792,N_34793,N_34794,N_34795,N_34796,N_34797,N_34798,N_34799,N_34800,N_34801,N_34802,N_34803,N_34804,N_34805,N_34806,N_34807,N_34808,N_34809,N_34810,N_34811,N_34812,N_34813,N_34814,N_34815,N_34816,N_34817,N_34818,N_34819,N_34820,N_34821,N_34822,N_34823,N_34824,N_34825,N_34826,N_34827,N_34828,N_34829,N_34830,N_34831,N_34832,N_34833,N_34834,N_34835,N_34836,N_34837,N_34838,N_34839,N_34840,N_34841,N_34842,N_34843,N_34844,N_34845,N_34846,N_34847,N_34848,N_34849,N_34850,N_34851,N_34852,N_34853,N_34854,N_34855,N_34856,N_34857,N_34858,N_34859,N_34860,N_34861,N_34862,N_34863,N_34864,N_34865,N_34866,N_34867,N_34868,N_34869,N_34870,N_34871,N_34872,N_34873,N_34874,N_34875,N_34876,N_34877,N_34878,N_34879,N_34880,N_34881,N_34882,N_34883,N_34884,N_34885,N_34886,N_34887,N_34888,N_34889,N_34890,N_34891,N_34892,N_34893,N_34894,N_34895,N_34896,N_34897,N_34898,N_34899,N_34900,N_34901,N_34902,N_34903,N_34904,N_34905,N_34906,N_34907,N_34908,N_34909,N_34910,N_34911,N_34912,N_34913,N_34914,N_34915,N_34916,N_34917,N_34918,N_34919,N_34920,N_34921,N_34922,N_34923,N_34924,N_34925,N_34926,N_34927,N_34928,N_34929,N_34930,N_34931,N_34932,N_34933,N_34934,N_34935,N_34936,N_34937,N_34938,N_34939,N_34940,N_34941,N_34942,N_34943,N_34944,N_34945,N_34946,N_34947,N_34948,N_34949,N_34950,N_34951,N_34952,N_34953,N_34954,N_34955,N_34956,N_34957,N_34958,N_34959,N_34960,N_34961,N_34962,N_34963,N_34964,N_34965,N_34966,N_34967,N_34968,N_34969,N_34970,N_34971,N_34972,N_34973,N_34974,N_34975,N_34976,N_34977,N_34978,N_34979,N_34980,N_34981,N_34982,N_34983,N_34984,N_34985,N_34986,N_34987,N_34988,N_34989,N_34990,N_34991,N_34992,N_34993,N_34994,N_34995,N_34996,N_34997,N_34998,N_34999,N_35000,N_35001,N_35002,N_35003,N_35004,N_35005,N_35006,N_35007,N_35008,N_35009,N_35010,N_35011,N_35012,N_35013,N_35014,N_35015,N_35016,N_35017,N_35018,N_35019,N_35020,N_35021,N_35022,N_35023,N_35024,N_35025,N_35026,N_35027,N_35028,N_35029,N_35030,N_35031,N_35032,N_35033,N_35034,N_35035,N_35036,N_35037,N_35038,N_35039,N_35040,N_35041,N_35042,N_35043,N_35044,N_35045,N_35046,N_35047,N_35048,N_35049,N_35050,N_35051,N_35052,N_35053,N_35054,N_35055,N_35056,N_35057,N_35058,N_35059,N_35060,N_35061,N_35062,N_35063,N_35064,N_35065,N_35066,N_35067,N_35068,N_35069,N_35070,N_35071,N_35072,N_35073,N_35074,N_35075,N_35076,N_35077,N_35078,N_35079,N_35080,N_35081,N_35082,N_35083,N_35084,N_35085,N_35086,N_35087,N_35088,N_35089,N_35090,N_35091,N_35092,N_35093,N_35094,N_35095,N_35096,N_35097,N_35098,N_35099,N_35100,N_35101,N_35102,N_35103,N_35104,N_35105,N_35106,N_35107,N_35108,N_35109,N_35110,N_35111,N_35112,N_35113,N_35114,N_35115,N_35116,N_35117,N_35118,N_35119,N_35120,N_35121,N_35122,N_35123,N_35124,N_35125,N_35126,N_35127,N_35128,N_35129,N_35130,N_35131,N_35132,N_35133,N_35134,N_35135,N_35136,N_35137,N_35138,N_35139,N_35140,N_35141,N_35142,N_35143,N_35144,N_35145,N_35146,N_35147,N_35148,N_35149,N_35150,N_35151,N_35152,N_35153,N_35154,N_35155,N_35156,N_35157,N_35158,N_35159,N_35160,N_35161,N_35162,N_35163,N_35164,N_35165,N_35166,N_35167,N_35168,N_35169,N_35170,N_35171,N_35172,N_35173,N_35174,N_35175,N_35176,N_35177,N_35178,N_35179,N_35180,N_35181,N_35182,N_35183,N_35184,N_35185,N_35186,N_35187,N_35188,N_35189,N_35190,N_35191,N_35192,N_35193,N_35194,N_35195,N_35196,N_35197,N_35198,N_35199,N_35200,N_35201,N_35202,N_35203,N_35204,N_35205,N_35206,N_35207,N_35208,N_35209,N_35210,N_35211,N_35212,N_35213,N_35214,N_35215,N_35216,N_35217,N_35218,N_35219,N_35220,N_35221,N_35222,N_35223,N_35224,N_35225,N_35226,N_35227,N_35228,N_35229,N_35230,N_35231,N_35232,N_35233,N_35234,N_35235,N_35236,N_35237,N_35238,N_35239,N_35240,N_35241,N_35242,N_35243,N_35244,N_35245,N_35246,N_35247,N_35248,N_35249,N_35250,N_35251,N_35252,N_35253,N_35254,N_35255,N_35256,N_35257,N_35258,N_35259,N_35260,N_35261,N_35262,N_35263,N_35264,N_35265,N_35266,N_35267,N_35268,N_35269,N_35270,N_35271,N_35272,N_35273,N_35274,N_35275,N_35276,N_35277,N_35278,N_35279,N_35280,N_35281,N_35282,N_35283,N_35284,N_35285,N_35286,N_35287,N_35288,N_35289,N_35290,N_35291,N_35292,N_35293,N_35294,N_35295,N_35296,N_35297,N_35298,N_35299,N_35300,N_35301,N_35302,N_35303,N_35304,N_35305,N_35306,N_35307,N_35308,N_35309,N_35310,N_35311,N_35312,N_35313,N_35314,N_35315,N_35316,N_35317,N_35318,N_35319,N_35320,N_35321,N_35322,N_35323,N_35324,N_35325,N_35326,N_35327,N_35328,N_35329,N_35330,N_35331,N_35332,N_35333,N_35334,N_35335,N_35336,N_35337,N_35338,N_35339,N_35340,N_35341,N_35342,N_35343,N_35344,N_35345,N_35346,N_35347,N_35348,N_35349,N_35350,N_35351,N_35352,N_35353,N_35354,N_35355,N_35356,N_35357,N_35358,N_35359,N_35360,N_35361,N_35362,N_35363,N_35364,N_35365,N_35366,N_35367,N_35368,N_35369,N_35370,N_35371,N_35372,N_35373,N_35374,N_35375,N_35376,N_35377,N_35378,N_35379,N_35380,N_35381,N_35382,N_35383,N_35384,N_35385,N_35386,N_35387,N_35388,N_35389,N_35390,N_35391,N_35392,N_35393,N_35394,N_35395,N_35396,N_35397,N_35398,N_35399,N_35400,N_35401,N_35402,N_35403,N_35404,N_35405,N_35406,N_35407,N_35408,N_35409,N_35410,N_35411,N_35412,N_35413,N_35414,N_35415,N_35416,N_35417,N_35418,N_35419,N_35420,N_35421,N_35422,N_35423,N_35424,N_35425,N_35426,N_35427,N_35428,N_35429,N_35430,N_35431,N_35432,N_35433,N_35434,N_35435,N_35436,N_35437,N_35438,N_35439,N_35440,N_35441,N_35442,N_35443,N_35444,N_35445,N_35446,N_35447,N_35448,N_35449,N_35450,N_35451,N_35452,N_35453,N_35454,N_35455,N_35456,N_35457,N_35458,N_35459,N_35460,N_35461,N_35462,N_35463,N_35464,N_35465,N_35466,N_35467,N_35468,N_35469,N_35470,N_35471,N_35472,N_35473,N_35474,N_35475,N_35476,N_35477,N_35478,N_35479,N_35480,N_35481,N_35482,N_35483,N_35484,N_35485,N_35486,N_35487,N_35488,N_35489,N_35490,N_35491,N_35492,N_35493,N_35494,N_35495,N_35496,N_35497,N_35498,N_35499,N_35500,N_35501,N_35502,N_35503,N_35504,N_35505,N_35506,N_35507,N_35508,N_35509,N_35510,N_35511,N_35512,N_35513,N_35514,N_35515,N_35516,N_35517,N_35518,N_35519,N_35520,N_35521,N_35522,N_35523,N_35524,N_35525,N_35526,N_35527,N_35528,N_35529,N_35530,N_35531,N_35532,N_35533,N_35534,N_35535,N_35536,N_35537,N_35538,N_35539,N_35540,N_35541,N_35542,N_35543,N_35544,N_35545,N_35546,N_35547,N_35548,N_35549,N_35550,N_35551,N_35552,N_35553,N_35554,N_35555,N_35556,N_35557,N_35558,N_35559,N_35560,N_35561,N_35562,N_35563,N_35564,N_35565,N_35566,N_35567,N_35568,N_35569,N_35570,N_35571,N_35572,N_35573,N_35574,N_35575,N_35576,N_35577,N_35578,N_35579,N_35580,N_35581,N_35582,N_35583,N_35584,N_35585,N_35586,N_35587,N_35588,N_35589,N_35590,N_35591,N_35592,N_35593,N_35594,N_35595,N_35596,N_35597,N_35598,N_35599,N_35600,N_35601,N_35602,N_35603,N_35604,N_35605,N_35606,N_35607,N_35608,N_35609,N_35610,N_35611,N_35612,N_35613,N_35614,N_35615,N_35616,N_35617,N_35618,N_35619,N_35620,N_35621,N_35622,N_35623,N_35624,N_35625,N_35626,N_35627,N_35628,N_35629,N_35630,N_35631,N_35632,N_35633,N_35634,N_35635,N_35636,N_35637,N_35638,N_35639,N_35640,N_35641,N_35642,N_35643,N_35644,N_35645,N_35646,N_35647,N_35648,N_35649,N_35650,N_35651,N_35652,N_35653,N_35654,N_35655,N_35656,N_35657,N_35658,N_35659,N_35660,N_35661,N_35662,N_35663,N_35664,N_35665,N_35666,N_35667,N_35668,N_35669,N_35670,N_35671,N_35672,N_35673,N_35674,N_35675,N_35676,N_35677,N_35678,N_35679,N_35680,N_35681,N_35682,N_35683,N_35684,N_35685,N_35686,N_35687,N_35688,N_35689,N_35690,N_35691,N_35692,N_35693,N_35694,N_35695,N_35696,N_35697,N_35698,N_35699,N_35700,N_35701,N_35702,N_35703,N_35704,N_35705,N_35706,N_35707,N_35708,N_35709,N_35710,N_35711,N_35712,N_35713,N_35714,N_35715,N_35716,N_35717,N_35718,N_35719,N_35720,N_35721,N_35722,N_35723,N_35724,N_35725,N_35726,N_35727,N_35728,N_35729,N_35730,N_35731,N_35732,N_35733,N_35734,N_35735,N_35736,N_35737,N_35738,N_35739,N_35740,N_35741,N_35742,N_35743,N_35744,N_35745,N_35746,N_35747,N_35748,N_35749,N_35750,N_35751,N_35752,N_35753,N_35754,N_35755,N_35756,N_35757,N_35758,N_35759,N_35760,N_35761,N_35762,N_35763,N_35764,N_35765,N_35766,N_35767,N_35768,N_35769,N_35770,N_35771,N_35772,N_35773,N_35774,N_35775,N_35776,N_35777,N_35778,N_35779,N_35780,N_35781,N_35782,N_35783,N_35784,N_35785,N_35786,N_35787,N_35788,N_35789,N_35790,N_35791,N_35792,N_35793,N_35794,N_35795,N_35796,N_35797,N_35798,N_35799,N_35800,N_35801,N_35802,N_35803,N_35804,N_35805,N_35806,N_35807,N_35808,N_35809,N_35810,N_35811,N_35812,N_35813,N_35814,N_35815,N_35816,N_35817,N_35818,N_35819,N_35820,N_35821,N_35822,N_35823,N_35824,N_35825,N_35826,N_35827,N_35828,N_35829,N_35830,N_35831,N_35832,N_35833,N_35834,N_35835,N_35836,N_35837,N_35838,N_35839,N_35840,N_35841,N_35842,N_35843,N_35844,N_35845,N_35846,N_35847,N_35848,N_35849,N_35850,N_35851,N_35852,N_35853,N_35854,N_35855,N_35856,N_35857,N_35858,N_35859,N_35860,N_35861,N_35862,N_35863,N_35864,N_35865,N_35866,N_35867,N_35868,N_35869,N_35870,N_35871,N_35872,N_35873,N_35874,N_35875,N_35876,N_35877,N_35878,N_35879,N_35880,N_35881,N_35882,N_35883,N_35884,N_35885,N_35886,N_35887,N_35888,N_35889,N_35890,N_35891,N_35892,N_35893,N_35894,N_35895,N_35896,N_35897,N_35898,N_35899,N_35900,N_35901,N_35902,N_35903,N_35904,N_35905,N_35906,N_35907,N_35908,N_35909,N_35910,N_35911,N_35912,N_35913,N_35914,N_35915,N_35916,N_35917,N_35918,N_35919,N_35920,N_35921,N_35922,N_35923,N_35924,N_35925,N_35926,N_35927,N_35928,N_35929,N_35930,N_35931,N_35932,N_35933,N_35934,N_35935,N_35936,N_35937,N_35938,N_35939,N_35940,N_35941,N_35942,N_35943,N_35944,N_35945,N_35946,N_35947,N_35948,N_35949,N_35950,N_35951,N_35952,N_35953,N_35954,N_35955,N_35956,N_35957,N_35958,N_35959,N_35960,N_35961,N_35962,N_35963,N_35964,N_35965,N_35966,N_35967,N_35968,N_35969,N_35970,N_35971,N_35972,N_35973,N_35974,N_35975,N_35976,N_35977,N_35978,N_35979,N_35980,N_35981,N_35982,N_35983,N_35984,N_35985,N_35986,N_35987,N_35988,N_35989,N_35990,N_35991,N_35992,N_35993,N_35994,N_35995,N_35996,N_35997,N_35998,N_35999,N_36000,N_36001,N_36002,N_36003,N_36004,N_36005,N_36006,N_36007,N_36008,N_36009,N_36010,N_36011,N_36012,N_36013,N_36014,N_36015,N_36016,N_36017,N_36018,N_36019,N_36020,N_36021,N_36022,N_36023,N_36024,N_36025,N_36026,N_36027,N_36028,N_36029,N_36030,N_36031,N_36032,N_36033,N_36034,N_36035,N_36036,N_36037,N_36038,N_36039,N_36040,N_36041,N_36042,N_36043,N_36044,N_36045,N_36046,N_36047,N_36048,N_36049,N_36050,N_36051,N_36052,N_36053,N_36054,N_36055,N_36056,N_36057,N_36058,N_36059,N_36060,N_36061,N_36062,N_36063,N_36064,N_36065,N_36066,N_36067,N_36068,N_36069,N_36070,N_36071,N_36072,N_36073,N_36074,N_36075,N_36076,N_36077,N_36078,N_36079,N_36080,N_36081,N_36082,N_36083,N_36084,N_36085,N_36086,N_36087,N_36088,N_36089,N_36090,N_36091,N_36092,N_36093,N_36094,N_36095,N_36096,N_36097,N_36098,N_36099,N_36100,N_36101,N_36102,N_36103,N_36104,N_36105,N_36106,N_36107,N_36108,N_36109,N_36110,N_36111,N_36112,N_36113,N_36114,N_36115,N_36116,N_36117,N_36118,N_36119,N_36120,N_36121,N_36122,N_36123,N_36124,N_36125,N_36126,N_36127,N_36128,N_36129,N_36130,N_36131,N_36132,N_36133,N_36134,N_36135,N_36136,N_36137,N_36138,N_36139,N_36140,N_36141,N_36142,N_36143,N_36144,N_36145,N_36146,N_36147,N_36148,N_36149,N_36150,N_36151,N_36152,N_36153,N_36154,N_36155,N_36156,N_36157,N_36158,N_36159,N_36160,N_36161,N_36162,N_36163,N_36164,N_36165,N_36166,N_36167,N_36168,N_36169,N_36170,N_36171,N_36172,N_36173,N_36174,N_36175,N_36176,N_36177,N_36178,N_36179,N_36180,N_36181,N_36182,N_36183,N_36184,N_36185,N_36186,N_36187,N_36188,N_36189,N_36190,N_36191,N_36192,N_36193,N_36194,N_36195,N_36196,N_36197,N_36198,N_36199,N_36200,N_36201,N_36202,N_36203,N_36204,N_36205,N_36206,N_36207,N_36208,N_36209,N_36210,N_36211,N_36212,N_36213,N_36214,N_36215,N_36216,N_36217,N_36218,N_36219,N_36220,N_36221,N_36222,N_36223,N_36224,N_36225,N_36226,N_36227,N_36228,N_36229,N_36230,N_36231,N_36232,N_36233,N_36234,N_36235,N_36236,N_36237,N_36238,N_36239,N_36240,N_36241,N_36242,N_36243,N_36244,N_36245,N_36246,N_36247,N_36248,N_36249,N_36250,N_36251,N_36252,N_36253,N_36254,N_36255,N_36256,N_36257,N_36258,N_36259,N_36260,N_36261,N_36262,N_36263,N_36264,N_36265,N_36266,N_36267,N_36268,N_36269,N_36270,N_36271,N_36272,N_36273,N_36274,N_36275,N_36276,N_36277,N_36278,N_36279,N_36280,N_36281,N_36282,N_36283,N_36284,N_36285,N_36286,N_36287,N_36288,N_36289,N_36290,N_36291,N_36292,N_36293,N_36294,N_36295,N_36296,N_36297,N_36298,N_36299,N_36300,N_36301,N_36302,N_36303,N_36304,N_36305,N_36306,N_36307,N_36308,N_36309,N_36310,N_36311,N_36312,N_36313,N_36314,N_36315,N_36316,N_36317,N_36318,N_36319,N_36320,N_36321,N_36322,N_36323,N_36324,N_36325,N_36326,N_36327,N_36328,N_36329,N_36330,N_36331,N_36332,N_36333,N_36334,N_36335,N_36336,N_36337,N_36338,N_36339,N_36340,N_36341,N_36342,N_36343,N_36344,N_36345,N_36346,N_36347,N_36348,N_36349,N_36350,N_36351,N_36352,N_36353,N_36354,N_36355,N_36356,N_36357,N_36358,N_36359,N_36360,N_36361,N_36362,N_36363,N_36364,N_36365,N_36366,N_36367,N_36368,N_36369,N_36370,N_36371,N_36372,N_36373,N_36374,N_36375,N_36376,N_36377,N_36378,N_36379,N_36380,N_36381,N_36382,N_36383,N_36384,N_36385,N_36386,N_36387,N_36388,N_36389,N_36390,N_36391,N_36392,N_36393,N_36394,N_36395,N_36396,N_36397,N_36398,N_36399,N_36400,N_36401,N_36402,N_36403,N_36404,N_36405,N_36406,N_36407,N_36408,N_36409,N_36410,N_36411,N_36412,N_36413,N_36414,N_36415,N_36416,N_36417,N_36418,N_36419,N_36420,N_36421,N_36422,N_36423,N_36424,N_36425,N_36426,N_36427,N_36428,N_36429,N_36430,N_36431,N_36432,N_36433,N_36434,N_36435,N_36436,N_36437,N_36438,N_36439,N_36440,N_36441,N_36442,N_36443,N_36444,N_36445,N_36446,N_36447,N_36448,N_36449,N_36450,N_36451,N_36452,N_36453,N_36454,N_36455,N_36456,N_36457,N_36458,N_36459,N_36460,N_36461,N_36462,N_36463,N_36464,N_36465,N_36466,N_36467,N_36468,N_36469,N_36470,N_36471,N_36472,N_36473,N_36474,N_36475,N_36476,N_36477,N_36478,N_36479,N_36480,N_36481,N_36482,N_36483,N_36484,N_36485,N_36486,N_36487,N_36488,N_36489,N_36490,N_36491,N_36492,N_36493,N_36494,N_36495,N_36496,N_36497,N_36498,N_36499,N_36500,N_36501,N_36502,N_36503,N_36504,N_36505,N_36506,N_36507,N_36508,N_36509,N_36510,N_36511,N_36512,N_36513,N_36514,N_36515,N_36516,N_36517,N_36518,N_36519,N_36520,N_36521,N_36522,N_36523,N_36524,N_36525,N_36526,N_36527,N_36528,N_36529,N_36530,N_36531,N_36532,N_36533,N_36534,N_36535,N_36536,N_36537,N_36538,N_36539,N_36540,N_36541,N_36542,N_36543,N_36544,N_36545,N_36546,N_36547,N_36548,N_36549,N_36550,N_36551,N_36552,N_36553,N_36554,N_36555,N_36556,N_36557,N_36558,N_36559,N_36560,N_36561,N_36562,N_36563,N_36564,N_36565,N_36566,N_36567,N_36568,N_36569,N_36570,N_36571,N_36572,N_36573,N_36574,N_36575,N_36576,N_36577,N_36578,N_36579,N_36580,N_36581,N_36582,N_36583,N_36584,N_36585,N_36586,N_36587,N_36588,N_36589,N_36590,N_36591,N_36592,N_36593,N_36594,N_36595,N_36596,N_36597,N_36598,N_36599,N_36600,N_36601,N_36602,N_36603,N_36604,N_36605,N_36606,N_36607,N_36608,N_36609,N_36610,N_36611,N_36612,N_36613,N_36614,N_36615,N_36616,N_36617,N_36618,N_36619,N_36620,N_36621,N_36622,N_36623,N_36624,N_36625,N_36626,N_36627,N_36628,N_36629,N_36630,N_36631,N_36632,N_36633,N_36634,N_36635,N_36636,N_36637,N_36638,N_36639,N_36640,N_36641,N_36642,N_36643,N_36644,N_36645,N_36646,N_36647,N_36648,N_36649,N_36650,N_36651,N_36652,N_36653,N_36654,N_36655,N_36656,N_36657,N_36658,N_36659,N_36660,N_36661,N_36662,N_36663,N_36664,N_36665,N_36666,N_36667,N_36668,N_36669,N_36670,N_36671,N_36672,N_36673,N_36674,N_36675,N_36676,N_36677,N_36678,N_36679,N_36680,N_36681,N_36682,N_36683,N_36684,N_36685,N_36686,N_36687,N_36688,N_36689,N_36690,N_36691,N_36692,N_36693,N_36694,N_36695,N_36696,N_36697,N_36698,N_36699,N_36700,N_36701,N_36702,N_36703,N_36704,N_36705,N_36706,N_36707,N_36708,N_36709,N_36710,N_36711,N_36712,N_36713,N_36714,N_36715,N_36716,N_36717,N_36718,N_36719,N_36720,N_36721,N_36722,N_36723,N_36724,N_36725,N_36726,N_36727,N_36728,N_36729,N_36730,N_36731,N_36732,N_36733,N_36734,N_36735,N_36736,N_36737,N_36738,N_36739,N_36740,N_36741,N_36742,N_36743,N_36744,N_36745,N_36746,N_36747,N_36748,N_36749,N_36750,N_36751,N_36752,N_36753,N_36754,N_36755,N_36756,N_36757,N_36758,N_36759,N_36760,N_36761,N_36762,N_36763,N_36764,N_36765,N_36766,N_36767,N_36768,N_36769,N_36770,N_36771,N_36772,N_36773,N_36774,N_36775,N_36776,N_36777,N_36778,N_36779,N_36780,N_36781,N_36782,N_36783,N_36784,N_36785,N_36786,N_36787,N_36788,N_36789,N_36790,N_36791,N_36792,N_36793,N_36794,N_36795,N_36796,N_36797,N_36798,N_36799,N_36800,N_36801,N_36802,N_36803,N_36804,N_36805,N_36806,N_36807,N_36808,N_36809,N_36810,N_36811,N_36812,N_36813,N_36814,N_36815,N_36816,N_36817,N_36818,N_36819,N_36820,N_36821,N_36822,N_36823,N_36824,N_36825,N_36826,N_36827,N_36828,N_36829,N_36830,N_36831,N_36832,N_36833,N_36834,N_36835,N_36836,N_36837,N_36838,N_36839,N_36840,N_36841,N_36842,N_36843,N_36844,N_36845,N_36846,N_36847,N_36848,N_36849,N_36850,N_36851,N_36852,N_36853,N_36854,N_36855,N_36856,N_36857,N_36858,N_36859,N_36860,N_36861,N_36862,N_36863,N_36864,N_36865,N_36866,N_36867,N_36868,N_36869,N_36870,N_36871,N_36872,N_36873,N_36874,N_36875,N_36876,N_36877,N_36878,N_36879,N_36880,N_36881,N_36882,N_36883,N_36884,N_36885,N_36886,N_36887,N_36888,N_36889,N_36890,N_36891,N_36892,N_36893,N_36894,N_36895,N_36896,N_36897,N_36898,N_36899,N_36900,N_36901,N_36902,N_36903,N_36904,N_36905,N_36906,N_36907,N_36908,N_36909,N_36910,N_36911,N_36912,N_36913,N_36914,N_36915,N_36916,N_36917,N_36918,N_36919,N_36920,N_36921,N_36922,N_36923,N_36924,N_36925,N_36926,N_36927,N_36928,N_36929,N_36930,N_36931,N_36932,N_36933,N_36934,N_36935,N_36936,N_36937,N_36938,N_36939,N_36940,N_36941,N_36942,N_36943,N_36944,N_36945,N_36946,N_36947,N_36948,N_36949,N_36950,N_36951,N_36952,N_36953,N_36954,N_36955,N_36956,N_36957,N_36958,N_36959,N_36960,N_36961,N_36962,N_36963,N_36964,N_36965,N_36966,N_36967,N_36968,N_36969,N_36970,N_36971,N_36972,N_36973,N_36974,N_36975,N_36976,N_36977,N_36978,N_36979,N_36980,N_36981,N_36982,N_36983,N_36984,N_36985,N_36986,N_36987,N_36988,N_36989,N_36990,N_36991,N_36992,N_36993,N_36994,N_36995,N_36996,N_36997,N_36998,N_36999,N_37000,N_37001,N_37002,N_37003,N_37004,N_37005,N_37006,N_37007,N_37008,N_37009,N_37010,N_37011,N_37012,N_37013,N_37014,N_37015,N_37016,N_37017,N_37018,N_37019,N_37020,N_37021,N_37022,N_37023,N_37024,N_37025,N_37026,N_37027,N_37028,N_37029,N_37030,N_37031,N_37032,N_37033,N_37034,N_37035,N_37036,N_37037,N_37038,N_37039,N_37040,N_37041,N_37042,N_37043,N_37044,N_37045,N_37046,N_37047,N_37048,N_37049,N_37050,N_37051,N_37052,N_37053,N_37054,N_37055,N_37056,N_37057,N_37058,N_37059,N_37060,N_37061,N_37062,N_37063,N_37064,N_37065,N_37066,N_37067,N_37068,N_37069,N_37070,N_37071,N_37072,N_37073,N_37074,N_37075,N_37076,N_37077,N_37078,N_37079,N_37080,N_37081,N_37082,N_37083,N_37084,N_37085,N_37086,N_37087,N_37088,N_37089,N_37090,N_37091,N_37092,N_37093,N_37094,N_37095,N_37096,N_37097,N_37098,N_37099,N_37100,N_37101,N_37102,N_37103,N_37104,N_37105,N_37106,N_37107,N_37108,N_37109,N_37110,N_37111,N_37112,N_37113,N_37114,N_37115,N_37116,N_37117,N_37118,N_37119,N_37120,N_37121,N_37122,N_37123,N_37124,N_37125,N_37126,N_37127,N_37128,N_37129,N_37130,N_37131,N_37132,N_37133,N_37134,N_37135,N_37136,N_37137,N_37138,N_37139,N_37140,N_37141,N_37142,N_37143,N_37144,N_37145,N_37146,N_37147,N_37148,N_37149,N_37150,N_37151,N_37152,N_37153,N_37154,N_37155,N_37156,N_37157,N_37158,N_37159,N_37160,N_37161,N_37162,N_37163,N_37164,N_37165,N_37166,N_37167,N_37168,N_37169,N_37170,N_37171,N_37172,N_37173,N_37174,N_37175,N_37176,N_37177,N_37178,N_37179,N_37180,N_37181,N_37182,N_37183,N_37184,N_37185,N_37186,N_37187,N_37188,N_37189,N_37190,N_37191,N_37192,N_37193,N_37194,N_37195,N_37196,N_37197,N_37198,N_37199,N_37200,N_37201,N_37202,N_37203,N_37204,N_37205,N_37206,N_37207,N_37208,N_37209,N_37210,N_37211,N_37212,N_37213,N_37214,N_37215,N_37216,N_37217,N_37218,N_37219,N_37220,N_37221,N_37222,N_37223,N_37224,N_37225,N_37226,N_37227,N_37228,N_37229,N_37230,N_37231,N_37232,N_37233,N_37234,N_37235,N_37236,N_37237,N_37238,N_37239,N_37240,N_37241,N_37242,N_37243,N_37244,N_37245,N_37246,N_37247,N_37248,N_37249,N_37250,N_37251,N_37252,N_37253,N_37254,N_37255,N_37256,N_37257,N_37258,N_37259,N_37260,N_37261,N_37262,N_37263,N_37264,N_37265,N_37266,N_37267,N_37268,N_37269,N_37270,N_37271,N_37272,N_37273,N_37274,N_37275,N_37276,N_37277,N_37278,N_37279,N_37280,N_37281,N_37282,N_37283,N_37284,N_37285,N_37286,N_37287,N_37288,N_37289,N_37290,N_37291,N_37292,N_37293,N_37294,N_37295,N_37296,N_37297,N_37298,N_37299,N_37300,N_37301,N_37302,N_37303,N_37304,N_37305,N_37306,N_37307,N_37308,N_37309,N_37310,N_37311,N_37312,N_37313,N_37314,N_37315,N_37316,N_37317,N_37318,N_37319,N_37320,N_37321,N_37322,N_37323,N_37324,N_37325,N_37326,N_37327,N_37328,N_37329,N_37330,N_37331,N_37332,N_37333,N_37334,N_37335,N_37336,N_37337,N_37338,N_37339,N_37340,N_37341,N_37342,N_37343,N_37344,N_37345,N_37346,N_37347,N_37348,N_37349,N_37350,N_37351,N_37352,N_37353,N_37354,N_37355,N_37356,N_37357,N_37358,N_37359,N_37360,N_37361,N_37362,N_37363,N_37364,N_37365,N_37366,N_37367,N_37368,N_37369,N_37370,N_37371,N_37372,N_37373,N_37374,N_37375,N_37376,N_37377,N_37378,N_37379,N_37380,N_37381,N_37382,N_37383,N_37384,N_37385,N_37386,N_37387,N_37388,N_37389,N_37390,N_37391,N_37392,N_37393,N_37394,N_37395,N_37396,N_37397,N_37398,N_37399,N_37400,N_37401,N_37402,N_37403,N_37404,N_37405,N_37406,N_37407,N_37408,N_37409,N_37410,N_37411,N_37412,N_37413,N_37414,N_37415,N_37416,N_37417,N_37418,N_37419,N_37420,N_37421,N_37422,N_37423,N_37424,N_37425,N_37426,N_37427,N_37428,N_37429,N_37430,N_37431,N_37432,N_37433,N_37434,N_37435,N_37436,N_37437,N_37438,N_37439,N_37440,N_37441,N_37442,N_37443,N_37444,N_37445,N_37446,N_37447,N_37448,N_37449,N_37450,N_37451,N_37452,N_37453,N_37454,N_37455,N_37456,N_37457,N_37458,N_37459,N_37460,N_37461,N_37462,N_37463,N_37464,N_37465,N_37466,N_37467,N_37468,N_37469,N_37470,N_37471,N_37472,N_37473,N_37474,N_37475,N_37476,N_37477,N_37478,N_37479,N_37480,N_37481,N_37482,N_37483,N_37484,N_37485,N_37486,N_37487,N_37488,N_37489,N_37490,N_37491,N_37492,N_37493,N_37494,N_37495,N_37496,N_37497,N_37498,N_37499,N_37500,N_37501,N_37502,N_37503,N_37504,N_37505,N_37506,N_37507,N_37508,N_37509,N_37510,N_37511,N_37512,N_37513,N_37514,N_37515,N_37516,N_37517,N_37518,N_37519,N_37520,N_37521,N_37522,N_37523,N_37524,N_37525,N_37526,N_37527,N_37528,N_37529,N_37530,N_37531,N_37532,N_37533,N_37534,N_37535,N_37536,N_37537,N_37538,N_37539,N_37540,N_37541,N_37542,N_37543,N_37544,N_37545,N_37546,N_37547,N_37548,N_37549,N_37550,N_37551,N_37552,N_37553,N_37554,N_37555,N_37556,N_37557,N_37558,N_37559,N_37560,N_37561,N_37562,N_37563,N_37564,N_37565,N_37566,N_37567,N_37568,N_37569,N_37570,N_37571,N_37572,N_37573,N_37574,N_37575,N_37576,N_37577,N_37578,N_37579,N_37580,N_37581,N_37582,N_37583,N_37584,N_37585,N_37586,N_37587,N_37588,N_37589,N_37590,N_37591,N_37592,N_37593,N_37594,N_37595,N_37596,N_37597,N_37598,N_37599,N_37600,N_37601,N_37602,N_37603,N_37604,N_37605,N_37606,N_37607,N_37608,N_37609,N_37610,N_37611,N_37612,N_37613,N_37614,N_37615,N_37616,N_37617,N_37618,N_37619,N_37620,N_37621,N_37622,N_37623,N_37624,N_37625,N_37626,N_37627,N_37628,N_37629,N_37630,N_37631,N_37632,N_37633,N_37634,N_37635,N_37636,N_37637,N_37638,N_37639,N_37640,N_37641,N_37642,N_37643,N_37644,N_37645,N_37646,N_37647,N_37648,N_37649,N_37650,N_37651,N_37652,N_37653,N_37654,N_37655,N_37656,N_37657,N_37658,N_37659,N_37660,N_37661,N_37662,N_37663,N_37664,N_37665,N_37666,N_37667,N_37668,N_37669,N_37670,N_37671,N_37672,N_37673,N_37674,N_37675,N_37676,N_37677,N_37678,N_37679,N_37680,N_37681,N_37682,N_37683,N_37684,N_37685,N_37686,N_37687,N_37688,N_37689,N_37690,N_37691,N_37692,N_37693,N_37694,N_37695,N_37696,N_37697,N_37698,N_37699,N_37700,N_37701,N_37702,N_37703,N_37704,N_37705,N_37706,N_37707,N_37708,N_37709,N_37710,N_37711,N_37712,N_37713,N_37714,N_37715,N_37716,N_37717,N_37718,N_37719,N_37720,N_37721,N_37722,N_37723,N_37724,N_37725,N_37726,N_37727,N_37728,N_37729,N_37730,N_37731,N_37732,N_37733,N_37734,N_37735,N_37736,N_37737,N_37738,N_37739,N_37740,N_37741,N_37742,N_37743,N_37744,N_37745,N_37746,N_37747,N_37748,N_37749,N_37750,N_37751,N_37752,N_37753,N_37754,N_37755,N_37756,N_37757,N_37758,N_37759,N_37760,N_37761,N_37762,N_37763,N_37764,N_37765,N_37766,N_37767,N_37768,N_37769,N_37770,N_37771,N_37772,N_37773,N_37774,N_37775,N_37776,N_37777,N_37778,N_37779,N_37780,N_37781,N_37782,N_37783,N_37784,N_37785,N_37786,N_37787,N_37788,N_37789,N_37790,N_37791,N_37792,N_37793,N_37794,N_37795,N_37796,N_37797,N_37798,N_37799,N_37800,N_37801,N_37802,N_37803,N_37804,N_37805,N_37806,N_37807,N_37808,N_37809,N_37810,N_37811,N_37812,N_37813,N_37814,N_37815,N_37816,N_37817,N_37818,N_37819,N_37820,N_37821,N_37822,N_37823,N_37824,N_37825,N_37826,N_37827,N_37828,N_37829,N_37830,N_37831,N_37832,N_37833,N_37834,N_37835,N_37836,N_37837,N_37838,N_37839,N_37840,N_37841,N_37842,N_37843,N_37844,N_37845,N_37846,N_37847,N_37848,N_37849,N_37850,N_37851,N_37852,N_37853,N_37854,N_37855,N_37856,N_37857,N_37858,N_37859,N_37860,N_37861,N_37862,N_37863,N_37864,N_37865,N_37866,N_37867,N_37868,N_37869,N_37870,N_37871,N_37872,N_37873,N_37874,N_37875,N_37876,N_37877,N_37878,N_37879,N_37880,N_37881,N_37882,N_37883,N_37884,N_37885,N_37886,N_37887,N_37888,N_37889,N_37890,N_37891,N_37892,N_37893,N_37894,N_37895,N_37896,N_37897,N_37898,N_37899,N_37900,N_37901,N_37902,N_37903,N_37904,N_37905,N_37906,N_37907,N_37908,N_37909,N_37910,N_37911,N_37912,N_37913,N_37914,N_37915,N_37916,N_37917,N_37918,N_37919,N_37920,N_37921,N_37922,N_37923,N_37924,N_37925,N_37926,N_37927,N_37928,N_37929,N_37930,N_37931,N_37932,N_37933,N_37934,N_37935,N_37936,N_37937,N_37938,N_37939,N_37940,N_37941,N_37942,N_37943,N_37944,N_37945,N_37946,N_37947,N_37948,N_37949,N_37950,N_37951,N_37952,N_37953,N_37954,N_37955,N_37956,N_37957,N_37958,N_37959,N_37960,N_37961,N_37962,N_37963,N_37964,N_37965,N_37966,N_37967,N_37968,N_37969,N_37970,N_37971,N_37972,N_37973,N_37974,N_37975,N_37976,N_37977,N_37978,N_37979,N_37980,N_37981,N_37982,N_37983,N_37984,N_37985,N_37986,N_37987,N_37988,N_37989,N_37990,N_37991,N_37992,N_37993,N_37994,N_37995,N_37996,N_37997,N_37998,N_37999,N_38000,N_38001,N_38002,N_38003,N_38004,N_38005,N_38006,N_38007,N_38008,N_38009,N_38010,N_38011,N_38012,N_38013,N_38014,N_38015,N_38016,N_38017,N_38018,N_38019,N_38020,N_38021,N_38022,N_38023,N_38024,N_38025,N_38026,N_38027,N_38028,N_38029,N_38030,N_38031,N_38032,N_38033,N_38034,N_38035,N_38036,N_38037,N_38038,N_38039,N_38040,N_38041,N_38042,N_38043,N_38044,N_38045,N_38046,N_38047,N_38048,N_38049,N_38050,N_38051,N_38052,N_38053,N_38054,N_38055,N_38056,N_38057,N_38058,N_38059,N_38060,N_38061,N_38062,N_38063,N_38064,N_38065,N_38066,N_38067,N_38068,N_38069,N_38070,N_38071,N_38072,N_38073,N_38074,N_38075,N_38076,N_38077,N_38078,N_38079,N_38080,N_38081,N_38082,N_38083,N_38084,N_38085,N_38086,N_38087,N_38088,N_38089,N_38090,N_38091,N_38092,N_38093,N_38094,N_38095,N_38096,N_38097,N_38098,N_38099,N_38100,N_38101,N_38102,N_38103,N_38104,N_38105,N_38106,N_38107,N_38108,N_38109,N_38110,N_38111,N_38112,N_38113,N_38114,N_38115,N_38116,N_38117,N_38118,N_38119,N_38120,N_38121,N_38122,N_38123,N_38124,N_38125,N_38126,N_38127,N_38128,N_38129,N_38130,N_38131,N_38132,N_38133,N_38134,N_38135,N_38136,N_38137,N_38138,N_38139,N_38140,N_38141,N_38142,N_38143,N_38144,N_38145,N_38146,N_38147,N_38148,N_38149,N_38150,N_38151,N_38152,N_38153,N_38154,N_38155,N_38156,N_38157,N_38158,N_38159,N_38160,N_38161,N_38162,N_38163,N_38164,N_38165,N_38166,N_38167,N_38168,N_38169,N_38170,N_38171,N_38172,N_38173,N_38174,N_38175,N_38176,N_38177,N_38178,N_38179,N_38180,N_38181,N_38182,N_38183,N_38184,N_38185,N_38186,N_38187,N_38188,N_38189,N_38190,N_38191,N_38192,N_38193,N_38194,N_38195,N_38196,N_38197,N_38198,N_38199,N_38200,N_38201,N_38202,N_38203,N_38204,N_38205,N_38206,N_38207,N_38208,N_38209,N_38210,N_38211,N_38212,N_38213,N_38214,N_38215,N_38216,N_38217,N_38218,N_38219,N_38220,N_38221,N_38222,N_38223,N_38224,N_38225,N_38226,N_38227,N_38228,N_38229,N_38230,N_38231,N_38232,N_38233,N_38234,N_38235,N_38236,N_38237,N_38238,N_38239,N_38240,N_38241,N_38242,N_38243,N_38244,N_38245,N_38246,N_38247,N_38248,N_38249,N_38250,N_38251,N_38252,N_38253,N_38254,N_38255,N_38256,N_38257,N_38258,N_38259,N_38260,N_38261,N_38262,N_38263,N_38264,N_38265,N_38266,N_38267,N_38268,N_38269,N_38270,N_38271,N_38272,N_38273,N_38274,N_38275,N_38276,N_38277,N_38278,N_38279,N_38280,N_38281,N_38282,N_38283,N_38284,N_38285,N_38286,N_38287,N_38288,N_38289,N_38290,N_38291,N_38292,N_38293,N_38294,N_38295,N_38296,N_38297,N_38298,N_38299,N_38300,N_38301,N_38302,N_38303,N_38304,N_38305,N_38306,N_38307,N_38308,N_38309,N_38310,N_38311,N_38312,N_38313,N_38314,N_38315,N_38316,N_38317,N_38318,N_38319,N_38320,N_38321,N_38322,N_38323,N_38324,N_38325,N_38326,N_38327,N_38328,N_38329,N_38330,N_38331,N_38332,N_38333,N_38334,N_38335,N_38336,N_38337,N_38338,N_38339,N_38340,N_38341,N_38342,N_38343,N_38344,N_38345,N_38346,N_38347,N_38348,N_38349,N_38350,N_38351,N_38352,N_38353,N_38354,N_38355,N_38356,N_38357,N_38358,N_38359,N_38360,N_38361,N_38362,N_38363,N_38364,N_38365,N_38366,N_38367,N_38368,N_38369,N_38370,N_38371,N_38372,N_38373,N_38374,N_38375,N_38376,N_38377,N_38378,N_38379,N_38380,N_38381,N_38382,N_38383,N_38384,N_38385,N_38386,N_38387,N_38388,N_38389,N_38390,N_38391,N_38392,N_38393,N_38394,N_38395,N_38396,N_38397,N_38398,N_38399,N_38400,N_38401,N_38402,N_38403,N_38404,N_38405,N_38406,N_38407,N_38408,N_38409,N_38410,N_38411,N_38412,N_38413,N_38414,N_38415,N_38416,N_38417,N_38418,N_38419,N_38420,N_38421,N_38422,N_38423,N_38424,N_38425,N_38426,N_38427,N_38428,N_38429,N_38430,N_38431,N_38432,N_38433,N_38434,N_38435,N_38436,N_38437,N_38438,N_38439,N_38440,N_38441,N_38442,N_38443,N_38444,N_38445,N_38446,N_38447,N_38448,N_38449,N_38450,N_38451,N_38452,N_38453,N_38454,N_38455,N_38456,N_38457,N_38458,N_38459,N_38460,N_38461,N_38462,N_38463,N_38464,N_38465,N_38466,N_38467,N_38468,N_38469,N_38470,N_38471,N_38472,N_38473,N_38474,N_38475,N_38476,N_38477,N_38478,N_38479,N_38480,N_38481,N_38482,N_38483,N_38484,N_38485,N_38486,N_38487,N_38488,N_38489,N_38490,N_38491,N_38492,N_38493,N_38494,N_38495,N_38496,N_38497,N_38498,N_38499,N_38500,N_38501,N_38502,N_38503,N_38504,N_38505,N_38506,N_38507,N_38508,N_38509,N_38510,N_38511,N_38512,N_38513,N_38514,N_38515,N_38516,N_38517,N_38518,N_38519,N_38520,N_38521,N_38522,N_38523,N_38524,N_38525,N_38526,N_38527,N_38528,N_38529,N_38530,N_38531,N_38532,N_38533,N_38534,N_38535,N_38536,N_38537,N_38538,N_38539,N_38540,N_38541,N_38542,N_38543,N_38544,N_38545,N_38546,N_38547,N_38548,N_38549,N_38550,N_38551,N_38552,N_38553,N_38554,N_38555,N_38556,N_38557,N_38558,N_38559,N_38560,N_38561,N_38562,N_38563,N_38564,N_38565,N_38566,N_38567,N_38568,N_38569,N_38570,N_38571,N_38572,N_38573,N_38574,N_38575,N_38576,N_38577,N_38578,N_38579,N_38580,N_38581,N_38582,N_38583,N_38584,N_38585,N_38586,N_38587,N_38588,N_38589,N_38590,N_38591,N_38592,N_38593,N_38594,N_38595,N_38596,N_38597,N_38598,N_38599,N_38600,N_38601,N_38602,N_38603,N_38604,N_38605,N_38606,N_38607,N_38608,N_38609,N_38610,N_38611,N_38612,N_38613,N_38614,N_38615,N_38616,N_38617,N_38618,N_38619,N_38620,N_38621,N_38622,N_38623,N_38624,N_38625,N_38626,N_38627,N_38628,N_38629,N_38630,N_38631,N_38632,N_38633,N_38634,N_38635,N_38636,N_38637,N_38638,N_38639,N_38640,N_38641,N_38642,N_38643,N_38644,N_38645,N_38646,N_38647,N_38648,N_38649,N_38650,N_38651,N_38652,N_38653,N_38654,N_38655,N_38656,N_38657,N_38658,N_38659,N_38660,N_38661,N_38662,N_38663,N_38664,N_38665,N_38666,N_38667,N_38668,N_38669,N_38670,N_38671,N_38672,N_38673,N_38674,N_38675,N_38676,N_38677,N_38678,N_38679,N_38680,N_38681,N_38682,N_38683,N_38684,N_38685,N_38686,N_38687,N_38688,N_38689,N_38690,N_38691,N_38692,N_38693,N_38694,N_38695,N_38696,N_38697,N_38698,N_38699,N_38700,N_38701,N_38702,N_38703,N_38704,N_38705,N_38706,N_38707,N_38708,N_38709,N_38710,N_38711,N_38712,N_38713,N_38714,N_38715,N_38716,N_38717,N_38718,N_38719,N_38720,N_38721,N_38722,N_38723,N_38724,N_38725,N_38726,N_38727,N_38728,N_38729,N_38730,N_38731,N_38732,N_38733,N_38734,N_38735,N_38736,N_38737,N_38738,N_38739,N_38740,N_38741,N_38742,N_38743,N_38744,N_38745,N_38746,N_38747,N_38748,N_38749,N_38750,N_38751,N_38752,N_38753,N_38754,N_38755,N_38756,N_38757,N_38758,N_38759,N_38760,N_38761,N_38762,N_38763,N_38764,N_38765,N_38766,N_38767,N_38768,N_38769,N_38770,N_38771,N_38772,N_38773,N_38774,N_38775,N_38776,N_38777,N_38778,N_38779,N_38780,N_38781,N_38782,N_38783,N_38784,N_38785,N_38786,N_38787,N_38788,N_38789,N_38790,N_38791,N_38792,N_38793,N_38794,N_38795,N_38796,N_38797,N_38798,N_38799,N_38800,N_38801,N_38802,N_38803,N_38804,N_38805,N_38806,N_38807,N_38808,N_38809,N_38810,N_38811,N_38812,N_38813,N_38814,N_38815,N_38816,N_38817,N_38818,N_38819,N_38820,N_38821,N_38822,N_38823,N_38824,N_38825,N_38826,N_38827,N_38828,N_38829,N_38830,N_38831,N_38832,N_38833,N_38834,N_38835,N_38836,N_38837,N_38838,N_38839,N_38840,N_38841,N_38842,N_38843,N_38844,N_38845,N_38846,N_38847,N_38848,N_38849,N_38850,N_38851,N_38852,N_38853,N_38854,N_38855,N_38856,N_38857,N_38858,N_38859,N_38860,N_38861,N_38862,N_38863,N_38864,N_38865,N_38866,N_38867,N_38868,N_38869,N_38870,N_38871,N_38872,N_38873,N_38874,N_38875,N_38876,N_38877,N_38878,N_38879,N_38880,N_38881,N_38882,N_38883,N_38884,N_38885,N_38886,N_38887,N_38888,N_38889,N_38890,N_38891,N_38892,N_38893,N_38894,N_38895,N_38896,N_38897,N_38898,N_38899,N_38900,N_38901,N_38902,N_38903,N_38904,N_38905,N_38906,N_38907,N_38908,N_38909,N_38910,N_38911,N_38912,N_38913,N_38914,N_38915,N_38916,N_38917,N_38918,N_38919,N_38920,N_38921,N_38922,N_38923,N_38924,N_38925,N_38926,N_38927,N_38928,N_38929,N_38930,N_38931,N_38932,N_38933,N_38934,N_38935,N_38936,N_38937,N_38938,N_38939,N_38940,N_38941,N_38942,N_38943,N_38944,N_38945,N_38946,N_38947,N_38948,N_38949,N_38950,N_38951,N_38952,N_38953,N_38954,N_38955,N_38956,N_38957,N_38958,N_38959,N_38960,N_38961,N_38962,N_38963,N_38964,N_38965,N_38966,N_38967,N_38968,N_38969,N_38970,N_38971,N_38972,N_38973,N_38974,N_38975,N_38976,N_38977,N_38978,N_38979,N_38980,N_38981,N_38982,N_38983,N_38984,N_38985,N_38986,N_38987,N_38988,N_38989,N_38990,N_38991,N_38992,N_38993,N_38994,N_38995,N_38996,N_38997,N_38998,N_38999,N_39000,N_39001,N_39002,N_39003,N_39004,N_39005,N_39006,N_39007,N_39008,N_39009,N_39010,N_39011,N_39012,N_39013,N_39014,N_39015,N_39016,N_39017,N_39018,N_39019,N_39020,N_39021,N_39022,N_39023,N_39024,N_39025,N_39026,N_39027,N_39028,N_39029,N_39030,N_39031,N_39032,N_39033,N_39034,N_39035,N_39036,N_39037,N_39038,N_39039,N_39040,N_39041,N_39042,N_39043,N_39044,N_39045,N_39046,N_39047,N_39048,N_39049,N_39050,N_39051,N_39052,N_39053,N_39054,N_39055,N_39056,N_39057,N_39058,N_39059,N_39060,N_39061,N_39062,N_39063,N_39064,N_39065,N_39066,N_39067,N_39068,N_39069,N_39070,N_39071,N_39072,N_39073,N_39074,N_39075,N_39076,N_39077,N_39078,N_39079,N_39080,N_39081,N_39082,N_39083,N_39084,N_39085,N_39086,N_39087,N_39088,N_39089,N_39090,N_39091,N_39092,N_39093,N_39094,N_39095,N_39096,N_39097,N_39098,N_39099,N_39100,N_39101,N_39102,N_39103,N_39104,N_39105,N_39106,N_39107,N_39108,N_39109,N_39110,N_39111,N_39112,N_39113,N_39114,N_39115,N_39116,N_39117,N_39118,N_39119,N_39120,N_39121,N_39122,N_39123,N_39124,N_39125,N_39126,N_39127,N_39128,N_39129,N_39130,N_39131,N_39132,N_39133,N_39134,N_39135,N_39136,N_39137,N_39138,N_39139,N_39140,N_39141,N_39142,N_39143,N_39144,N_39145,N_39146,N_39147,N_39148,N_39149,N_39150,N_39151,N_39152,N_39153,N_39154,N_39155,N_39156,N_39157,N_39158,N_39159,N_39160,N_39161,N_39162,N_39163,N_39164,N_39165,N_39166,N_39167,N_39168,N_39169,N_39170,N_39171,N_39172,N_39173,N_39174,N_39175,N_39176,N_39177,N_39178,N_39179,N_39180,N_39181,N_39182,N_39183,N_39184,N_39185,N_39186,N_39187,N_39188,N_39189,N_39190,N_39191,N_39192,N_39193,N_39194,N_39195,N_39196,N_39197,N_39198,N_39199,N_39200,N_39201,N_39202,N_39203,N_39204,N_39205,N_39206,N_39207,N_39208,N_39209,N_39210,N_39211,N_39212,N_39213,N_39214,N_39215,N_39216,N_39217,N_39218,N_39219,N_39220,N_39221,N_39222,N_39223,N_39224,N_39225,N_39226,N_39227,N_39228,N_39229,N_39230,N_39231,N_39232,N_39233,N_39234,N_39235,N_39236,N_39237,N_39238,N_39239,N_39240,N_39241,N_39242,N_39243,N_39244,N_39245,N_39246,N_39247,N_39248,N_39249,N_39250,N_39251,N_39252,N_39253,N_39254,N_39255,N_39256,N_39257,N_39258,N_39259,N_39260,N_39261,N_39262,N_39263,N_39264,N_39265,N_39266,N_39267,N_39268,N_39269,N_39270,N_39271,N_39272,N_39273,N_39274,N_39275,N_39276,N_39277,N_39278,N_39279,N_39280,N_39281,N_39282,N_39283,N_39284,N_39285,N_39286,N_39287,N_39288,N_39289,N_39290,N_39291,N_39292,N_39293,N_39294,N_39295,N_39296,N_39297,N_39298,N_39299,N_39300,N_39301,N_39302,N_39303,N_39304,N_39305,N_39306,N_39307,N_39308,N_39309,N_39310,N_39311,N_39312,N_39313,N_39314,N_39315,N_39316,N_39317,N_39318,N_39319,N_39320,N_39321,N_39322,N_39323,N_39324,N_39325,N_39326,N_39327,N_39328,N_39329,N_39330,N_39331,N_39332,N_39333,N_39334,N_39335,N_39336,N_39337,N_39338,N_39339,N_39340,N_39341,N_39342,N_39343,N_39344,N_39345,N_39346,N_39347,N_39348,N_39349,N_39350,N_39351,N_39352,N_39353,N_39354,N_39355,N_39356,N_39357,N_39358,N_39359,N_39360,N_39361,N_39362,N_39363,N_39364,N_39365,N_39366,N_39367,N_39368,N_39369,N_39370,N_39371,N_39372,N_39373,N_39374,N_39375,N_39376,N_39377,N_39378,N_39379,N_39380,N_39381,N_39382,N_39383,N_39384,N_39385,N_39386,N_39387,N_39388,N_39389,N_39390,N_39391,N_39392,N_39393,N_39394,N_39395,N_39396,N_39397,N_39398,N_39399,N_39400,N_39401,N_39402,N_39403,N_39404,N_39405,N_39406,N_39407,N_39408,N_39409,N_39410,N_39411,N_39412,N_39413,N_39414,N_39415,N_39416,N_39417,N_39418,N_39419,N_39420,N_39421,N_39422,N_39423,N_39424,N_39425,N_39426,N_39427,N_39428,N_39429,N_39430,N_39431,N_39432,N_39433,N_39434,N_39435,N_39436,N_39437,N_39438,N_39439,N_39440,N_39441,N_39442,N_39443,N_39444,N_39445,N_39446,N_39447,N_39448,N_39449,N_39450,N_39451,N_39452,N_39453,N_39454,N_39455,N_39456,N_39457,N_39458,N_39459,N_39460,N_39461,N_39462,N_39463,N_39464,N_39465,N_39466,N_39467,N_39468,N_39469,N_39470,N_39471,N_39472,N_39473,N_39474,N_39475,N_39476,N_39477,N_39478,N_39479,N_39480,N_39481,N_39482,N_39483,N_39484,N_39485,N_39486,N_39487,N_39488,N_39489,N_39490,N_39491,N_39492,N_39493,N_39494,N_39495,N_39496,N_39497,N_39498,N_39499,N_39500,N_39501,N_39502,N_39503,N_39504,N_39505,N_39506,N_39507,N_39508,N_39509,N_39510,N_39511,N_39512,N_39513,N_39514,N_39515,N_39516,N_39517,N_39518,N_39519,N_39520,N_39521,N_39522,N_39523,N_39524,N_39525,N_39526,N_39527,N_39528,N_39529,N_39530,N_39531,N_39532,N_39533,N_39534,N_39535,N_39536,N_39537,N_39538,N_39539,N_39540,N_39541,N_39542,N_39543,N_39544,N_39545,N_39546,N_39547,N_39548,N_39549,N_39550,N_39551,N_39552,N_39553,N_39554,N_39555,N_39556,N_39557,N_39558,N_39559,N_39560,N_39561,N_39562,N_39563,N_39564,N_39565,N_39566,N_39567,N_39568,N_39569,N_39570,N_39571,N_39572,N_39573,N_39574,N_39575,N_39576,N_39577,N_39578,N_39579,N_39580,N_39581,N_39582,N_39583,N_39584,N_39585,N_39586,N_39587,N_39588,N_39589,N_39590,N_39591,N_39592,N_39593,N_39594,N_39595,N_39596,N_39597,N_39598,N_39599,N_39600,N_39601,N_39602,N_39603,N_39604,N_39605,N_39606,N_39607,N_39608,N_39609,N_39610,N_39611,N_39612,N_39613,N_39614,N_39615,N_39616,N_39617,N_39618,N_39619,N_39620,N_39621,N_39622,N_39623,N_39624,N_39625,N_39626,N_39627,N_39628,N_39629,N_39630,N_39631,N_39632,N_39633,N_39634,N_39635,N_39636,N_39637,N_39638,N_39639,N_39640,N_39641,N_39642,N_39643,N_39644,N_39645,N_39646,N_39647,N_39648,N_39649,N_39650,N_39651,N_39652,N_39653,N_39654,N_39655,N_39656,N_39657,N_39658,N_39659,N_39660,N_39661,N_39662,N_39663,N_39664,N_39665,N_39666,N_39667,N_39668,N_39669,N_39670,N_39671,N_39672,N_39673,N_39674,N_39675,N_39676,N_39677,N_39678,N_39679,N_39680,N_39681,N_39682,N_39683,N_39684,N_39685,N_39686,N_39687,N_39688,N_39689,N_39690,N_39691,N_39692,N_39693,N_39694,N_39695,N_39696,N_39697,N_39698,N_39699,N_39700,N_39701,N_39702,N_39703,N_39704,N_39705,N_39706,N_39707,N_39708,N_39709,N_39710,N_39711,N_39712,N_39713,N_39714,N_39715,N_39716,N_39717,N_39718,N_39719,N_39720,N_39721,N_39722,N_39723,N_39724,N_39725,N_39726,N_39727,N_39728,N_39729,N_39730,N_39731,N_39732,N_39733,N_39734,N_39735,N_39736,N_39737,N_39738,N_39739,N_39740,N_39741,N_39742,N_39743,N_39744,N_39745,N_39746,N_39747,N_39748,N_39749,N_39750,N_39751,N_39752,N_39753,N_39754,N_39755,N_39756,N_39757,N_39758,N_39759,N_39760,N_39761,N_39762,N_39763,N_39764,N_39765,N_39766,N_39767,N_39768,N_39769,N_39770,N_39771,N_39772,N_39773,N_39774,N_39775,N_39776,N_39777,N_39778,N_39779,N_39780,N_39781,N_39782,N_39783,N_39784,N_39785,N_39786,N_39787,N_39788,N_39789,N_39790,N_39791,N_39792,N_39793,N_39794,N_39795,N_39796,N_39797,N_39798,N_39799,N_39800,N_39801,N_39802,N_39803,N_39804,N_39805,N_39806,N_39807,N_39808,N_39809,N_39810,N_39811,N_39812,N_39813,N_39814,N_39815,N_39816,N_39817,N_39818,N_39819,N_39820,N_39821,N_39822,N_39823,N_39824,N_39825,N_39826,N_39827,N_39828,N_39829,N_39830,N_39831,N_39832,N_39833,N_39834,N_39835,N_39836,N_39837,N_39838,N_39839,N_39840,N_39841,N_39842,N_39843,N_39844,N_39845,N_39846,N_39847,N_39848,N_39849,N_39850,N_39851,N_39852,N_39853,N_39854,N_39855,N_39856,N_39857,N_39858,N_39859,N_39860,N_39861,N_39862,N_39863,N_39864,N_39865,N_39866,N_39867,N_39868,N_39869,N_39870,N_39871,N_39872,N_39873,N_39874,N_39875,N_39876,N_39877,N_39878,N_39879,N_39880,N_39881,N_39882,N_39883,N_39884,N_39885,N_39886,N_39887,N_39888,N_39889,N_39890,N_39891,N_39892,N_39893,N_39894,N_39895,N_39896,N_39897,N_39898,N_39899,N_39900,N_39901,N_39902,N_39903,N_39904,N_39905,N_39906,N_39907,N_39908,N_39909,N_39910,N_39911,N_39912,N_39913,N_39914,N_39915,N_39916,N_39917,N_39918,N_39919,N_39920,N_39921,N_39922,N_39923,N_39924,N_39925,N_39926,N_39927,N_39928,N_39929,N_39930,N_39931,N_39932,N_39933,N_39934,N_39935,N_39936,N_39937,N_39938,N_39939,N_39940,N_39941,N_39942,N_39943,N_39944,N_39945,N_39946,N_39947,N_39948,N_39949,N_39950,N_39951,N_39952,N_39953,N_39954,N_39955,N_39956,N_39957,N_39958,N_39959,N_39960,N_39961,N_39962,N_39963,N_39964,N_39965,N_39966,N_39967,N_39968,N_39969,N_39970,N_39971,N_39972,N_39973,N_39974,N_39975,N_39976,N_39977,N_39978,N_39979,N_39980,N_39981,N_39982,N_39983,N_39984,N_39985,N_39986,N_39987,N_39988,N_39989,N_39990,N_39991,N_39992,N_39993,N_39994,N_39995,N_39996,N_39997,N_39998,N_39999,N_40000,N_40001,N_40002,N_40003,N_40004,N_40005,N_40006,N_40007,N_40008,N_40009,N_40010,N_40011,N_40012,N_40013,N_40014,N_40015,N_40016,N_40017,N_40018,N_40019,N_40020,N_40021,N_40022,N_40023,N_40024,N_40025,N_40026,N_40027,N_40028,N_40029,N_40030,N_40031,N_40032,N_40033,N_40034,N_40035,N_40036,N_40037,N_40038,N_40039,N_40040,N_40041,N_40042,N_40043,N_40044,N_40045,N_40046,N_40047,N_40048,N_40049,N_40050,N_40051,N_40052,N_40053,N_40054,N_40055,N_40056,N_40057,N_40058,N_40059,N_40060,N_40061,N_40062,N_40063,N_40064,N_40065,N_40066,N_40067,N_40068,N_40069,N_40070,N_40071,N_40072,N_40073,N_40074,N_40075,N_40076,N_40077,N_40078,N_40079,N_40080,N_40081,N_40082,N_40083,N_40084,N_40085,N_40086,N_40087,N_40088,N_40089,N_40090,N_40091,N_40092,N_40093,N_40094,N_40095,N_40096,N_40097,N_40098,N_40099,N_40100,N_40101,N_40102,N_40103,N_40104,N_40105,N_40106,N_40107,N_40108,N_40109,N_40110,N_40111,N_40112,N_40113,N_40114,N_40115,N_40116,N_40117,N_40118,N_40119,N_40120,N_40121,N_40122,N_40123,N_40124,N_40125,N_40126,N_40127,N_40128,N_40129,N_40130,N_40131,N_40132,N_40133,N_40134,N_40135,N_40136,N_40137,N_40138,N_40139,N_40140,N_40141,N_40142,N_40143,N_40144,N_40145,N_40146,N_40147,N_40148,N_40149,N_40150,N_40151,N_40152,N_40153,N_40154,N_40155,N_40156,N_40157,N_40158,N_40159,N_40160,N_40161,N_40162,N_40163,N_40164,N_40165,N_40166,N_40167,N_40168,N_40169,N_40170,N_40171,N_40172,N_40173,N_40174,N_40175,N_40176,N_40177,N_40178,N_40179,N_40180,N_40181,N_40182,N_40183,N_40184,N_40185,N_40186,N_40187,N_40188,N_40189,N_40190,N_40191,N_40192,N_40193,N_40194,N_40195,N_40196,N_40197,N_40198,N_40199,N_40200,N_40201,N_40202,N_40203,N_40204,N_40205,N_40206,N_40207,N_40208,N_40209,N_40210,N_40211,N_40212,N_40213,N_40214,N_40215,N_40216,N_40217,N_40218,N_40219,N_40220,N_40221,N_40222,N_40223,N_40224,N_40225,N_40226,N_40227,N_40228,N_40229,N_40230,N_40231,N_40232,N_40233,N_40234,N_40235,N_40236,N_40237,N_40238,N_40239,N_40240,N_40241,N_40242,N_40243,N_40244,N_40245,N_40246,N_40247,N_40248,N_40249,N_40250,N_40251,N_40252,N_40253,N_40254,N_40255,N_40256,N_40257,N_40258,N_40259,N_40260,N_40261,N_40262,N_40263,N_40264,N_40265,N_40266,N_40267,N_40268,N_40269,N_40270,N_40271,N_40272,N_40273,N_40274,N_40275,N_40276,N_40277,N_40278,N_40279,N_40280,N_40281,N_40282,N_40283,N_40284,N_40285,N_40286,N_40287,N_40288,N_40289,N_40290,N_40291,N_40292,N_40293,N_40294,N_40295,N_40296,N_40297,N_40298,N_40299,N_40300,N_40301,N_40302,N_40303,N_40304,N_40305,N_40306,N_40307,N_40308,N_40309,N_40310,N_40311,N_40312,N_40313,N_40314,N_40315,N_40316,N_40317,N_40318,N_40319,N_40320,N_40321,N_40322,N_40323,N_40324,N_40325,N_40326,N_40327,N_40328,N_40329,N_40330,N_40331,N_40332,N_40333,N_40334,N_40335,N_40336,N_40337,N_40338,N_40339,N_40340,N_40341,N_40342,N_40343,N_40344,N_40345,N_40346,N_40347,N_40348,N_40349,N_40350,N_40351,N_40352,N_40353,N_40354,N_40355,N_40356,N_40357,N_40358,N_40359,N_40360,N_40361,N_40362,N_40363,N_40364,N_40365,N_40366,N_40367,N_40368,N_40369,N_40370,N_40371,N_40372,N_40373,N_40374,N_40375,N_40376,N_40377,N_40378,N_40379,N_40380,N_40381,N_40382,N_40383,N_40384,N_40385,N_40386,N_40387,N_40388,N_40389,N_40390,N_40391,N_40392,N_40393,N_40394,N_40395,N_40396,N_40397,N_40398,N_40399,N_40400,N_40401,N_40402,N_40403,N_40404,N_40405,N_40406,N_40407,N_40408,N_40409,N_40410,N_40411,N_40412,N_40413,N_40414,N_40415,N_40416,N_40417,N_40418,N_40419,N_40420,N_40421,N_40422,N_40423,N_40424,N_40425,N_40426,N_40427,N_40428,N_40429,N_40430,N_40431,N_40432,N_40433,N_40434,N_40435,N_40436,N_40437,N_40438,N_40439,N_40440,N_40441,N_40442,N_40443,N_40444,N_40445,N_40446,N_40447,N_40448,N_40449,N_40450,N_40451,N_40452,N_40453,N_40454,N_40455,N_40456,N_40457,N_40458,N_40459,N_40460,N_40461,N_40462,N_40463,N_40464,N_40465,N_40466,N_40467,N_40468,N_40469,N_40470,N_40471,N_40472,N_40473,N_40474,N_40475,N_40476,N_40477,N_40478,N_40479,N_40480,N_40481,N_40482,N_40483,N_40484,N_40485,N_40486,N_40487,N_40488,N_40489,N_40490,N_40491,N_40492,N_40493,N_40494,N_40495,N_40496,N_40497,N_40498,N_40499,N_40500,N_40501,N_40502,N_40503,N_40504,N_40505,N_40506,N_40507,N_40508,N_40509,N_40510,N_40511,N_40512,N_40513,N_40514,N_40515,N_40516,N_40517,N_40518,N_40519,N_40520,N_40521,N_40522,N_40523,N_40524,N_40525,N_40526,N_40527,N_40528,N_40529,N_40530,N_40531,N_40532,N_40533,N_40534,N_40535,N_40536,N_40537,N_40538,N_40539,N_40540,N_40541,N_40542,N_40543,N_40544,N_40545,N_40546,N_40547,N_40548,N_40549,N_40550,N_40551,N_40552,N_40553,N_40554,N_40555,N_40556,N_40557,N_40558,N_40559,N_40560,N_40561,N_40562,N_40563,N_40564,N_40565,N_40566,N_40567,N_40568,N_40569,N_40570,N_40571,N_40572,N_40573,N_40574,N_40575,N_40576,N_40577,N_40578,N_40579,N_40580,N_40581,N_40582,N_40583,N_40584,N_40585,N_40586,N_40587,N_40588,N_40589,N_40590,N_40591,N_40592,N_40593,N_40594,N_40595,N_40596,N_40597,N_40598,N_40599,N_40600,N_40601,N_40602,N_40603,N_40604,N_40605,N_40606,N_40607,N_40608,N_40609,N_40610,N_40611,N_40612,N_40613,N_40614,N_40615,N_40616,N_40617,N_40618,N_40619,N_40620,N_40621,N_40622,N_40623,N_40624,N_40625,N_40626,N_40627,N_40628,N_40629,N_40630,N_40631,N_40632,N_40633,N_40634,N_40635,N_40636,N_40637,N_40638,N_40639,N_40640,N_40641,N_40642,N_40643,N_40644,N_40645,N_40646,N_40647,N_40648,N_40649,N_40650,N_40651,N_40652,N_40653,N_40654,N_40655,N_40656,N_40657,N_40658,N_40659,N_40660,N_40661,N_40662,N_40663,N_40664,N_40665,N_40666,N_40667,N_40668,N_40669,N_40670,N_40671,N_40672,N_40673,N_40674,N_40675,N_40676,N_40677,N_40678,N_40679,N_40680,N_40681,N_40682,N_40683,N_40684,N_40685,N_40686,N_40687,N_40688,N_40689,N_40690,N_40691,N_40692,N_40693,N_40694,N_40695,N_40696,N_40697,N_40698,N_40699,N_40700,N_40701,N_40702,N_40703,N_40704,N_40705,N_40706,N_40707,N_40708,N_40709,N_40710,N_40711,N_40712,N_40713,N_40714,N_40715,N_40716,N_40717,N_40718,N_40719,N_40720,N_40721,N_40722,N_40723,N_40724,N_40725,N_40726,N_40727,N_40728,N_40729,N_40730,N_40731,N_40732,N_40733,N_40734,N_40735,N_40736,N_40737,N_40738,N_40739,N_40740,N_40741,N_40742,N_40743,N_40744,N_40745,N_40746,N_40747,N_40748,N_40749,N_40750,N_40751,N_40752,N_40753,N_40754,N_40755,N_40756,N_40757,N_40758,N_40759,N_40760,N_40761,N_40762,N_40763,N_40764,N_40765,N_40766,N_40767,N_40768,N_40769,N_40770,N_40771,N_40772,N_40773,N_40774,N_40775,N_40776,N_40777,N_40778,N_40779,N_40780,N_40781,N_40782,N_40783,N_40784,N_40785,N_40786,N_40787,N_40788,N_40789,N_40790,N_40791,N_40792,N_40793,N_40794,N_40795,N_40796,N_40797,N_40798,N_40799,N_40800,N_40801,N_40802,N_40803,N_40804,N_40805,N_40806,N_40807,N_40808,N_40809,N_40810,N_40811,N_40812,N_40813,N_40814,N_40815,N_40816,N_40817,N_40818,N_40819,N_40820,N_40821,N_40822,N_40823,N_40824,N_40825,N_40826,N_40827,N_40828,N_40829,N_40830,N_40831,N_40832,N_40833,N_40834,N_40835,N_40836,N_40837,N_40838,N_40839,N_40840,N_40841,N_40842,N_40843,N_40844,N_40845,N_40846,N_40847,N_40848,N_40849,N_40850,N_40851,N_40852,N_40853,N_40854,N_40855,N_40856,N_40857,N_40858,N_40859,N_40860,N_40861,N_40862,N_40863,N_40864,N_40865,N_40866,N_40867,N_40868,N_40869,N_40870,N_40871,N_40872,N_40873,N_40874,N_40875,N_40876,N_40877,N_40878,N_40879,N_40880,N_40881,N_40882,N_40883,N_40884,N_40885,N_40886,N_40887,N_40888,N_40889,N_40890,N_40891,N_40892,N_40893,N_40894,N_40895,N_40896,N_40897,N_40898,N_40899,N_40900,N_40901,N_40902,N_40903,N_40904,N_40905,N_40906,N_40907,N_40908,N_40909,N_40910,N_40911,N_40912,N_40913,N_40914,N_40915,N_40916,N_40917,N_40918,N_40919,N_40920,N_40921,N_40922,N_40923,N_40924,N_40925,N_40926,N_40927,N_40928,N_40929,N_40930,N_40931,N_40932,N_40933,N_40934,N_40935,N_40936,N_40937,N_40938,N_40939,N_40940,N_40941,N_40942,N_40943,N_40944,N_40945,N_40946,N_40947,N_40948,N_40949,N_40950,N_40951,N_40952,N_40953,N_40954,N_40955,N_40956,N_40957,N_40958,N_40959,N_40960,N_40961,N_40962,N_40963,N_40964,N_40965,N_40966,N_40967,N_40968,N_40969,N_40970,N_40971,N_40972,N_40973,N_40974,N_40975,N_40976,N_40977,N_40978,N_40979,N_40980,N_40981,N_40982,N_40983,N_40984,N_40985,N_40986,N_40987,N_40988,N_40989,N_40990,N_40991,N_40992,N_40993,N_40994,N_40995,N_40996,N_40997,N_40998,N_40999,N_41000,N_41001,N_41002,N_41003,N_41004,N_41005,N_41006,N_41007,N_41008,N_41009,N_41010,N_41011,N_41012,N_41013,N_41014,N_41015,N_41016,N_41017,N_41018,N_41019,N_41020,N_41021,N_41022,N_41023,N_41024,N_41025,N_41026,N_41027,N_41028,N_41029,N_41030,N_41031,N_41032,N_41033,N_41034,N_41035,N_41036,N_41037,N_41038,N_41039,N_41040,N_41041,N_41042,N_41043,N_41044,N_41045,N_41046,N_41047,N_41048,N_41049,N_41050,N_41051,N_41052,N_41053,N_41054,N_41055,N_41056,N_41057,N_41058,N_41059,N_41060,N_41061,N_41062,N_41063,N_41064,N_41065,N_41066,N_41067,N_41068,N_41069,N_41070,N_41071,N_41072,N_41073,N_41074,N_41075,N_41076,N_41077,N_41078,N_41079,N_41080,N_41081,N_41082,N_41083,N_41084,N_41085,N_41086,N_41087,N_41088,N_41089,N_41090,N_41091,N_41092,N_41093,N_41094,N_41095,N_41096,N_41097,N_41098,N_41099,N_41100,N_41101,N_41102,N_41103,N_41104,N_41105,N_41106,N_41107,N_41108,N_41109,N_41110,N_41111,N_41112,N_41113,N_41114,N_41115,N_41116,N_41117,N_41118,N_41119,N_41120,N_41121,N_41122,N_41123,N_41124,N_41125,N_41126,N_41127,N_41128,N_41129,N_41130,N_41131,N_41132,N_41133,N_41134,N_41135,N_41136,N_41137,N_41138,N_41139,N_41140,N_41141,N_41142,N_41143,N_41144,N_41145,N_41146,N_41147,N_41148,N_41149,N_41150,N_41151,N_41152,N_41153,N_41154,N_41155,N_41156,N_41157,N_41158,N_41159,N_41160,N_41161,N_41162,N_41163,N_41164,N_41165,N_41166,N_41167,N_41168,N_41169,N_41170,N_41171,N_41172,N_41173,N_41174,N_41175,N_41176,N_41177,N_41178,N_41179,N_41180,N_41181,N_41182,N_41183,N_41184,N_41185,N_41186,N_41187,N_41188,N_41189,N_41190,N_41191,N_41192,N_41193,N_41194,N_41195,N_41196,N_41197,N_41198,N_41199,N_41200,N_41201,N_41202,N_41203,N_41204,N_41205,N_41206,N_41207,N_41208,N_41209,N_41210,N_41211,N_41212,N_41213,N_41214,N_41215,N_41216,N_41217,N_41218,N_41219,N_41220,N_41221,N_41222,N_41223,N_41224,N_41225,N_41226,N_41227,N_41228,N_41229,N_41230,N_41231,N_41232,N_41233,N_41234,N_41235,N_41236,N_41237,N_41238,N_41239,N_41240,N_41241,N_41242,N_41243,N_41244,N_41245,N_41246,N_41247,N_41248,N_41249,N_41250,N_41251,N_41252,N_41253,N_41254,N_41255,N_41256,N_41257,N_41258,N_41259,N_41260,N_41261,N_41262,N_41263,N_41264,N_41265,N_41266,N_41267,N_41268,N_41269,N_41270,N_41271,N_41272,N_41273,N_41274,N_41275,N_41276,N_41277,N_41278,N_41279,N_41280,N_41281,N_41282,N_41283,N_41284,N_41285,N_41286,N_41287,N_41288,N_41289,N_41290,N_41291,N_41292,N_41293,N_41294,N_41295,N_41296,N_41297,N_41298,N_41299,N_41300,N_41301,N_41302,N_41303,N_41304,N_41305,N_41306,N_41307,N_41308,N_41309,N_41310,N_41311,N_41312,N_41313,N_41314,N_41315,N_41316,N_41317,N_41318,N_41319,N_41320,N_41321,N_41322,N_41323,N_41324,N_41325,N_41326,N_41327,N_41328,N_41329,N_41330,N_41331,N_41332,N_41333,N_41334,N_41335,N_41336,N_41337,N_41338,N_41339,N_41340,N_41341,N_41342,N_41343,N_41344,N_41345,N_41346,N_41347,N_41348,N_41349,N_41350,N_41351,N_41352,N_41353,N_41354,N_41355,N_41356,N_41357,N_41358,N_41359,N_41360,N_41361,N_41362,N_41363,N_41364,N_41365,N_41366,N_41367,N_41368,N_41369,N_41370,N_41371,N_41372,N_41373,N_41374,N_41375,N_41376,N_41377,N_41378,N_41379,N_41380,N_41381,N_41382,N_41383,N_41384,N_41385,N_41386,N_41387,N_41388,N_41389,N_41390,N_41391,N_41392,N_41393,N_41394,N_41395,N_41396,N_41397,N_41398,N_41399,N_41400,N_41401,N_41402,N_41403,N_41404,N_41405,N_41406,N_41407,N_41408,N_41409,N_41410,N_41411,N_41412,N_41413,N_41414,N_41415,N_41416,N_41417,N_41418,N_41419,N_41420,N_41421,N_41422,N_41423,N_41424,N_41425,N_41426,N_41427,N_41428,N_41429,N_41430,N_41431,N_41432,N_41433,N_41434,N_41435,N_41436,N_41437,N_41438,N_41439,N_41440,N_41441,N_41442,N_41443,N_41444,N_41445,N_41446,N_41447,N_41448,N_41449,N_41450,N_41451,N_41452,N_41453,N_41454,N_41455,N_41456,N_41457,N_41458,N_41459,N_41460,N_41461,N_41462,N_41463,N_41464,N_41465,N_41466,N_41467,N_41468,N_41469,N_41470,N_41471,N_41472,N_41473,N_41474,N_41475,N_41476,N_41477,N_41478,N_41479,N_41480,N_41481,N_41482,N_41483,N_41484,N_41485,N_41486,N_41487,N_41488,N_41489,N_41490,N_41491,N_41492,N_41493,N_41494,N_41495,N_41496,N_41497,N_41498,N_41499,N_41500,N_41501,N_41502,N_41503,N_41504,N_41505,N_41506,N_41507,N_41508,N_41509,N_41510,N_41511,N_41512,N_41513,N_41514,N_41515,N_41516,N_41517,N_41518,N_41519,N_41520,N_41521,N_41522,N_41523,N_41524,N_41525,N_41526,N_41527,N_41528,N_41529,N_41530,N_41531,N_41532,N_41533,N_41534,N_41535,N_41536,N_41537,N_41538,N_41539,N_41540,N_41541,N_41542,N_41543,N_41544,N_41545,N_41546,N_41547,N_41548,N_41549,N_41550,N_41551,N_41552,N_41553,N_41554,N_41555,N_41556,N_41557,N_41558,N_41559,N_41560,N_41561,N_41562,N_41563,N_41564,N_41565,N_41566,N_41567,N_41568,N_41569,N_41570,N_41571,N_41572,N_41573,N_41574,N_41575,N_41576,N_41577,N_41578,N_41579,N_41580,N_41581,N_41582,N_41583,N_41584,N_41585,N_41586,N_41587,N_41588,N_41589,N_41590,N_41591,N_41592,N_41593,N_41594,N_41595,N_41596,N_41597,N_41598,N_41599,N_41600,N_41601,N_41602,N_41603,N_41604,N_41605,N_41606,N_41607,N_41608,N_41609,N_41610,N_41611,N_41612,N_41613,N_41614,N_41615,N_41616,N_41617,N_41618,N_41619,N_41620,N_41621,N_41622,N_41623,N_41624,N_41625,N_41626,N_41627,N_41628,N_41629,N_41630,N_41631,N_41632,N_41633,N_41634,N_41635,N_41636,N_41637,N_41638,N_41639,N_41640,N_41641,N_41642,N_41643,N_41644,N_41645,N_41646,N_41647,N_41648,N_41649,N_41650,N_41651,N_41652,N_41653,N_41654,N_41655,N_41656,N_41657,N_41658,N_41659,N_41660,N_41661,N_41662,N_41663,N_41664,N_41665,N_41666,N_41667,N_41668,N_41669,N_41670,N_41671,N_41672,N_41673,N_41674,N_41675,N_41676,N_41677,N_41678,N_41679,N_41680,N_41681,N_41682,N_41683,N_41684,N_41685,N_41686,N_41687,N_41688,N_41689,N_41690,N_41691,N_41692,N_41693,N_41694,N_41695,N_41696,N_41697,N_41698,N_41699,N_41700,N_41701,N_41702,N_41703,N_41704,N_41705,N_41706,N_41707,N_41708,N_41709,N_41710,N_41711,N_41712,N_41713,N_41714,N_41715,N_41716,N_41717,N_41718,N_41719,N_41720,N_41721,N_41722,N_41723,N_41724,N_41725,N_41726,N_41727,N_41728,N_41729,N_41730,N_41731,N_41732,N_41733,N_41734,N_41735,N_41736,N_41737,N_41738,N_41739,N_41740,N_41741,N_41742,N_41743,N_41744,N_41745,N_41746,N_41747,N_41748,N_41749,N_41750,N_41751,N_41752,N_41753,N_41754,N_41755,N_41756,N_41757,N_41758,N_41759,N_41760,N_41761,N_41762,N_41763,N_41764,N_41765,N_41766,N_41767,N_41768,N_41769,N_41770,N_41771,N_41772,N_41773,N_41774,N_41775,N_41776,N_41777,N_41778,N_41779,N_41780,N_41781,N_41782,N_41783,N_41784,N_41785,N_41786,N_41787,N_41788,N_41789,N_41790,N_41791,N_41792,N_41793,N_41794,N_41795,N_41796,N_41797,N_41798,N_41799,N_41800,N_41801,N_41802,N_41803,N_41804,N_41805,N_41806,N_41807,N_41808,N_41809,N_41810,N_41811,N_41812,N_41813,N_41814,N_41815,N_41816,N_41817,N_41818,N_41819,N_41820,N_41821,N_41822,N_41823,N_41824,N_41825,N_41826,N_41827,N_41828,N_41829,N_41830,N_41831,N_41832,N_41833,N_41834,N_41835,N_41836,N_41837,N_41838,N_41839,N_41840,N_41841,N_41842,N_41843,N_41844,N_41845,N_41846,N_41847,N_41848,N_41849,N_41850,N_41851,N_41852,N_41853,N_41854,N_41855,N_41856,N_41857,N_41858,N_41859,N_41860,N_41861,N_41862,N_41863,N_41864,N_41865,N_41866,N_41867,N_41868,N_41869,N_41870,N_41871,N_41872,N_41873,N_41874,N_41875,N_41876,N_41877,N_41878,N_41879,N_41880,N_41881,N_41882,N_41883,N_41884,N_41885,N_41886,N_41887,N_41888,N_41889,N_41890,N_41891,N_41892,N_41893,N_41894,N_41895,N_41896,N_41897,N_41898,N_41899,N_41900,N_41901,N_41902,N_41903,N_41904,N_41905,N_41906,N_41907,N_41908,N_41909,N_41910,N_41911,N_41912,N_41913,N_41914,N_41915,N_41916,N_41917,N_41918,N_41919,N_41920,N_41921,N_41922,N_41923,N_41924,N_41925,N_41926,N_41927,N_41928,N_41929,N_41930,N_41931,N_41932,N_41933,N_41934,N_41935,N_41936,N_41937,N_41938,N_41939,N_41940,N_41941,N_41942,N_41943,N_41944,N_41945,N_41946,N_41947,N_41948,N_41949,N_41950,N_41951,N_41952,N_41953,N_41954,N_41955,N_41956,N_41957,N_41958,N_41959,N_41960,N_41961,N_41962,N_41963,N_41964,N_41965,N_41966,N_41967,N_41968,N_41969,N_41970,N_41971,N_41972,N_41973,N_41974,N_41975,N_41976,N_41977,N_41978,N_41979,N_41980,N_41981,N_41982,N_41983,N_41984,N_41985,N_41986,N_41987,N_41988,N_41989,N_41990,N_41991,N_41992,N_41993,N_41994,N_41995,N_41996,N_41997,N_41998,N_41999,N_42000,N_42001,N_42002,N_42003,N_42004,N_42005,N_42006,N_42007,N_42008,N_42009,N_42010,N_42011,N_42012,N_42013,N_42014,N_42015,N_42016,N_42017,N_42018,N_42019,N_42020,N_42021,N_42022,N_42023,N_42024,N_42025,N_42026,N_42027,N_42028,N_42029,N_42030,N_42031,N_42032,N_42033,N_42034,N_42035,N_42036,N_42037,N_42038,N_42039,N_42040,N_42041,N_42042,N_42043,N_42044,N_42045,N_42046,N_42047,N_42048,N_42049,N_42050,N_42051,N_42052,N_42053,N_42054,N_42055,N_42056,N_42057,N_42058,N_42059,N_42060,N_42061,N_42062,N_42063,N_42064,N_42065,N_42066,N_42067,N_42068,N_42069,N_42070,N_42071,N_42072,N_42073,N_42074,N_42075,N_42076,N_42077,N_42078,N_42079,N_42080,N_42081,N_42082,N_42083,N_42084,N_42085,N_42086,N_42087,N_42088,N_42089,N_42090,N_42091,N_42092,N_42093,N_42094,N_42095,N_42096,N_42097,N_42098,N_42099,N_42100,N_42101,N_42102,N_42103,N_42104,N_42105,N_42106,N_42107,N_42108,N_42109,N_42110,N_42111,N_42112,N_42113,N_42114,N_42115,N_42116,N_42117,N_42118,N_42119,N_42120,N_42121,N_42122,N_42123,N_42124,N_42125,N_42126,N_42127,N_42128,N_42129,N_42130,N_42131,N_42132,N_42133,N_42134,N_42135,N_42136,N_42137,N_42138,N_42139,N_42140,N_42141,N_42142,N_42143,N_42144,N_42145,N_42146,N_42147,N_42148,N_42149,N_42150,N_42151,N_42152,N_42153,N_42154,N_42155,N_42156,N_42157,N_42158,N_42159,N_42160,N_42161,N_42162,N_42163,N_42164,N_42165,N_42166,N_42167,N_42168,N_42169,N_42170,N_42171,N_42172,N_42173,N_42174,N_42175,N_42176,N_42177,N_42178,N_42179,N_42180,N_42181,N_42182,N_42183,N_42184,N_42185,N_42186,N_42187,N_42188,N_42189,N_42190,N_42191,N_42192,N_42193,N_42194,N_42195,N_42196,N_42197,N_42198,N_42199,N_42200,N_42201,N_42202,N_42203,N_42204,N_42205,N_42206,N_42207,N_42208,N_42209,N_42210,N_42211,N_42212,N_42213,N_42214,N_42215,N_42216,N_42217,N_42218,N_42219,N_42220,N_42221,N_42222,N_42223,N_42224,N_42225,N_42226,N_42227,N_42228,N_42229,N_42230,N_42231,N_42232,N_42233,N_42234,N_42235,N_42236,N_42237,N_42238,N_42239,N_42240,N_42241,N_42242,N_42243,N_42244,N_42245,N_42246,N_42247,N_42248,N_42249,N_42250,N_42251,N_42252,N_42253,N_42254,N_42255,N_42256,N_42257,N_42258,N_42259,N_42260,N_42261,N_42262,N_42263,N_42264,N_42265,N_42266,N_42267,N_42268,N_42269,N_42270,N_42271,N_42272,N_42273,N_42274,N_42275,N_42276,N_42277,N_42278,N_42279,N_42280,N_42281,N_42282,N_42283,N_42284,N_42285,N_42286,N_42287,N_42288,N_42289,N_42290,N_42291,N_42292,N_42293,N_42294,N_42295,N_42296,N_42297,N_42298,N_42299,N_42300,N_42301,N_42302,N_42303,N_42304,N_42305,N_42306,N_42307,N_42308,N_42309,N_42310,N_42311,N_42312,N_42313,N_42314,N_42315,N_42316,N_42317,N_42318,N_42319,N_42320,N_42321,N_42322,N_42323,N_42324,N_42325,N_42326,N_42327,N_42328,N_42329,N_42330,N_42331,N_42332,N_42333,N_42334,N_42335,N_42336,N_42337,N_42338,N_42339,N_42340,N_42341,N_42342,N_42343,N_42344,N_42345,N_42346,N_42347,N_42348,N_42349,N_42350,N_42351,N_42352,N_42353,N_42354,N_42355,N_42356,N_42357,N_42358,N_42359,N_42360,N_42361,N_42362,N_42363,N_42364,N_42365,N_42366,N_42367,N_42368,N_42369,N_42370,N_42371,N_42372,N_42373,N_42374,N_42375,N_42376,N_42377,N_42378,N_42379,N_42380,N_42381,N_42382,N_42383,N_42384,N_42385,N_42386,N_42387,N_42388,N_42389,N_42390,N_42391,N_42392,N_42393,N_42394,N_42395,N_42396,N_42397,N_42398,N_42399,N_42400,N_42401,N_42402,N_42403,N_42404,N_42405,N_42406,N_42407,N_42408,N_42409,N_42410,N_42411,N_42412,N_42413,N_42414,N_42415,N_42416,N_42417,N_42418,N_42419,N_42420,N_42421,N_42422,N_42423,N_42424,N_42425,N_42426,N_42427,N_42428,N_42429,N_42430,N_42431,N_42432,N_42433,N_42434,N_42435,N_42436,N_42437,N_42438,N_42439,N_42440,N_42441,N_42442,N_42443,N_42444,N_42445,N_42446,N_42447,N_42448,N_42449,N_42450,N_42451,N_42452,N_42453,N_42454,N_42455,N_42456,N_42457,N_42458,N_42459,N_42460,N_42461,N_42462,N_42463,N_42464,N_42465,N_42466,N_42467,N_42468,N_42469,N_42470,N_42471,N_42472,N_42473,N_42474,N_42475,N_42476,N_42477,N_42478,N_42479,N_42480,N_42481,N_42482,N_42483,N_42484,N_42485,N_42486,N_42487,N_42488,N_42489,N_42490,N_42491,N_42492,N_42493,N_42494,N_42495,N_42496,N_42497,N_42498,N_42499,N_42500,N_42501,N_42502,N_42503,N_42504,N_42505,N_42506,N_42507,N_42508,N_42509,N_42510,N_42511,N_42512,N_42513,N_42514,N_42515,N_42516,N_42517,N_42518,N_42519,N_42520,N_42521,N_42522,N_42523,N_42524,N_42525,N_42526,N_42527,N_42528,N_42529,N_42530,N_42531,N_42532,N_42533,N_42534,N_42535,N_42536,N_42537,N_42538,N_42539,N_42540,N_42541,N_42542,N_42543,N_42544,N_42545,N_42546,N_42547,N_42548,N_42549,N_42550,N_42551,N_42552,N_42553,N_42554,N_42555,N_42556,N_42557,N_42558,N_42559,N_42560,N_42561,N_42562,N_42563,N_42564,N_42565,N_42566,N_42567,N_42568,N_42569,N_42570,N_42571,N_42572,N_42573,N_42574,N_42575,N_42576,N_42577,N_42578,N_42579,N_42580,N_42581,N_42582,N_42583,N_42584,N_42585,N_42586,N_42587,N_42588,N_42589,N_42590,N_42591,N_42592,N_42593,N_42594,N_42595,N_42596,N_42597,N_42598,N_42599,N_42600,N_42601,N_42602,N_42603,N_42604,N_42605,N_42606,N_42607,N_42608,N_42609,N_42610,N_42611,N_42612,N_42613,N_42614,N_42615,N_42616,N_42617,N_42618,N_42619,N_42620,N_42621,N_42622,N_42623,N_42624,N_42625,N_42626,N_42627,N_42628,N_42629,N_42630,N_42631,N_42632,N_42633,N_42634,N_42635,N_42636,N_42637,N_42638,N_42639,N_42640,N_42641,N_42642,N_42643,N_42644,N_42645,N_42646,N_42647,N_42648,N_42649,N_42650,N_42651,N_42652,N_42653,N_42654,N_42655,N_42656,N_42657,N_42658,N_42659,N_42660,N_42661,N_42662,N_42663,N_42664,N_42665,N_42666,N_42667,N_42668,N_42669,N_42670,N_42671,N_42672,N_42673,N_42674,N_42675,N_42676,N_42677,N_42678,N_42679,N_42680,N_42681,N_42682,N_42683,N_42684,N_42685,N_42686,N_42687,N_42688,N_42689,N_42690,N_42691,N_42692,N_42693,N_42694,N_42695,N_42696,N_42697,N_42698,N_42699,N_42700,N_42701,N_42702,N_42703,N_42704,N_42705,N_42706,N_42707,N_42708,N_42709,N_42710,N_42711,N_42712,N_42713,N_42714,N_42715,N_42716,N_42717,N_42718,N_42719,N_42720,N_42721,N_42722,N_42723,N_42724,N_42725,N_42726,N_42727,N_42728,N_42729,N_42730,N_42731,N_42732,N_42733,N_42734,N_42735,N_42736,N_42737,N_42738,N_42739,N_42740,N_42741,N_42742,N_42743,N_42744,N_42745,N_42746,N_42747,N_42748,N_42749,N_42750,N_42751,N_42752,N_42753,N_42754,N_42755,N_42756,N_42757,N_42758,N_42759,N_42760,N_42761,N_42762,N_42763,N_42764,N_42765,N_42766,N_42767,N_42768,N_42769,N_42770,N_42771,N_42772,N_42773,N_42774,N_42775,N_42776,N_42777,N_42778,N_42779,N_42780,N_42781,N_42782,N_42783,N_42784,N_42785,N_42786,N_42787,N_42788,N_42789,N_42790,N_42791,N_42792,N_42793,N_42794,N_42795,N_42796,N_42797,N_42798,N_42799,N_42800,N_42801,N_42802,N_42803,N_42804,N_42805,N_42806,N_42807,N_42808,N_42809,N_42810,N_42811,N_42812,N_42813,N_42814,N_42815,N_42816,N_42817,N_42818,N_42819,N_42820,N_42821,N_42822,N_42823,N_42824,N_42825,N_42826,N_42827,N_42828,N_42829,N_42830,N_42831,N_42832,N_42833,N_42834,N_42835,N_42836,N_42837,N_42838,N_42839,N_42840,N_42841,N_42842,N_42843,N_42844,N_42845,N_42846,N_42847,N_42848,N_42849,N_42850,N_42851,N_42852,N_42853,N_42854,N_42855,N_42856,N_42857,N_42858,N_42859,N_42860,N_42861,N_42862,N_42863,N_42864,N_42865,N_42866,N_42867,N_42868,N_42869,N_42870,N_42871,N_42872,N_42873,N_42874,N_42875,N_42876,N_42877,N_42878,N_42879,N_42880,N_42881,N_42882,N_42883,N_42884,N_42885,N_42886,N_42887,N_42888,N_42889,N_42890,N_42891,N_42892,N_42893,N_42894,N_42895,N_42896,N_42897,N_42898,N_42899,N_42900,N_42901,N_42902,N_42903,N_42904,N_42905,N_42906,N_42907,N_42908,N_42909,N_42910,N_42911,N_42912,N_42913,N_42914,N_42915,N_42916,N_42917,N_42918,N_42919,N_42920,N_42921,N_42922,N_42923,N_42924,N_42925,N_42926,N_42927,N_42928,N_42929,N_42930,N_42931,N_42932,N_42933,N_42934,N_42935,N_42936,N_42937,N_42938,N_42939,N_42940,N_42941,N_42942,N_42943,N_42944,N_42945,N_42946,N_42947,N_42948,N_42949,N_42950,N_42951,N_42952,N_42953,N_42954,N_42955,N_42956,N_42957,N_42958,N_42959,N_42960,N_42961,N_42962,N_42963,N_42964,N_42965,N_42966,N_42967,N_42968,N_42969,N_42970,N_42971,N_42972,N_42973,N_42974,N_42975,N_42976,N_42977,N_42978,N_42979,N_42980,N_42981,N_42982,N_42983,N_42984,N_42985,N_42986,N_42987,N_42988,N_42989,N_42990,N_42991,N_42992,N_42993,N_42994,N_42995,N_42996,N_42997,N_42998,N_42999,N_43000,N_43001,N_43002,N_43003,N_43004,N_43005,N_43006,N_43007,N_43008,N_43009,N_43010,N_43011,N_43012,N_43013,N_43014,N_43015,N_43016,N_43017,N_43018,N_43019,N_43020,N_43021,N_43022,N_43023,N_43024,N_43025,N_43026,N_43027,N_43028,N_43029,N_43030,N_43031,N_43032,N_43033,N_43034,N_43035,N_43036,N_43037,N_43038,N_43039,N_43040,N_43041,N_43042,N_43043,N_43044,N_43045,N_43046,N_43047,N_43048,N_43049,N_43050,N_43051,N_43052,N_43053,N_43054,N_43055,N_43056,N_43057,N_43058,N_43059,N_43060,N_43061,N_43062,N_43063,N_43064,N_43065,N_43066,N_43067,N_43068,N_43069,N_43070,N_43071,N_43072,N_43073,N_43074,N_43075,N_43076,N_43077,N_43078,N_43079,N_43080,N_43081,N_43082,N_43083,N_43084,N_43085,N_43086,N_43087,N_43088,N_43089,N_43090,N_43091,N_43092,N_43093,N_43094,N_43095,N_43096,N_43097,N_43098,N_43099,N_43100,N_43101,N_43102,N_43103,N_43104,N_43105,N_43106,N_43107,N_43108,N_43109,N_43110,N_43111,N_43112,N_43113,N_43114,N_43115,N_43116,N_43117,N_43118,N_43119,N_43120,N_43121,N_43122,N_43123,N_43124,N_43125,N_43126,N_43127,N_43128,N_43129,N_43130,N_43131,N_43132,N_43133,N_43134,N_43135,N_43136,N_43137,N_43138,N_43139,N_43140,N_43141,N_43142,N_43143,N_43144,N_43145,N_43146,N_43147,N_43148,N_43149,N_43150,N_43151,N_43152,N_43153,N_43154,N_43155,N_43156,N_43157,N_43158,N_43159,N_43160,N_43161,N_43162,N_43163,N_43164,N_43165,N_43166,N_43167,N_43168,N_43169,N_43170,N_43171,N_43172,N_43173,N_43174,N_43175,N_43176,N_43177,N_43178,N_43179,N_43180,N_43181,N_43182,N_43183,N_43184,N_43185,N_43186,N_43187,N_43188,N_43189,N_43190,N_43191,N_43192,N_43193,N_43194,N_43195,N_43196,N_43197,N_43198,N_43199,N_43200,N_43201,N_43202,N_43203,N_43204,N_43205,N_43206,N_43207,N_43208,N_43209,N_43210,N_43211,N_43212,N_43213,N_43214,N_43215,N_43216,N_43217,N_43218,N_43219,N_43220,N_43221,N_43222,N_43223,N_43224,N_43225,N_43226,N_43227,N_43228,N_43229,N_43230,N_43231,N_43232,N_43233,N_43234,N_43235,N_43236,N_43237,N_43238,N_43239,N_43240,N_43241,N_43242,N_43243,N_43244,N_43245,N_43246,N_43247,N_43248,N_43249,N_43250,N_43251,N_43252,N_43253,N_43254,N_43255,N_43256,N_43257,N_43258,N_43259,N_43260,N_43261,N_43262,N_43263,N_43264,N_43265,N_43266,N_43267,N_43268,N_43269,N_43270,N_43271,N_43272,N_43273,N_43274,N_43275,N_43276,N_43277,N_43278,N_43279,N_43280,N_43281,N_43282,N_43283,N_43284,N_43285,N_43286,N_43287,N_43288,N_43289,N_43290,N_43291,N_43292,N_43293,N_43294,N_43295,N_43296,N_43297,N_43298,N_43299,N_43300,N_43301,N_43302,N_43303,N_43304,N_43305,N_43306,N_43307,N_43308,N_43309,N_43310,N_43311,N_43312,N_43313,N_43314,N_43315,N_43316,N_43317,N_43318,N_43319,N_43320,N_43321,N_43322,N_43323,N_43324,N_43325,N_43326,N_43327,N_43328,N_43329,N_43330,N_43331,N_43332,N_43333,N_43334,N_43335,N_43336,N_43337,N_43338,N_43339,N_43340,N_43341,N_43342,N_43343,N_43344,N_43345,N_43346,N_43347,N_43348,N_43349,N_43350,N_43351,N_43352,N_43353,N_43354,N_43355,N_43356,N_43357,N_43358,N_43359,N_43360,N_43361,N_43362,N_43363,N_43364,N_43365,N_43366,N_43367,N_43368,N_43369,N_43370,N_43371,N_43372,N_43373,N_43374,N_43375,N_43376,N_43377,N_43378,N_43379,N_43380,N_43381,N_43382,N_43383,N_43384,N_43385,N_43386,N_43387,N_43388,N_43389,N_43390,N_43391,N_43392,N_43393,N_43394,N_43395,N_43396,N_43397,N_43398,N_43399,N_43400,N_43401,N_43402,N_43403,N_43404,N_43405,N_43406,N_43407,N_43408,N_43409,N_43410,N_43411,N_43412,N_43413,N_43414,N_43415,N_43416,N_43417,N_43418,N_43419,N_43420,N_43421,N_43422,N_43423,N_43424,N_43425,N_43426,N_43427,N_43428,N_43429,N_43430,N_43431,N_43432,N_43433,N_43434,N_43435,N_43436,N_43437,N_43438,N_43439,N_43440,N_43441,N_43442,N_43443,N_43444,N_43445,N_43446,N_43447,N_43448,N_43449,N_43450,N_43451,N_43452,N_43453,N_43454,N_43455,N_43456,N_43457,N_43458,N_43459,N_43460,N_43461,N_43462,N_43463,N_43464,N_43465,N_43466,N_43467,N_43468,N_43469,N_43470,N_43471,N_43472,N_43473,N_43474,N_43475,N_43476,N_43477,N_43478,N_43479,N_43480,N_43481,N_43482,N_43483,N_43484,N_43485,N_43486,N_43487,N_43488,N_43489,N_43490,N_43491,N_43492,N_43493,N_43494,N_43495,N_43496,N_43497,N_43498,N_43499,N_43500,N_43501,N_43502,N_43503,N_43504,N_43505,N_43506,N_43507,N_43508,N_43509,N_43510,N_43511,N_43512,N_43513,N_43514,N_43515,N_43516,N_43517,N_43518,N_43519,N_43520,N_43521,N_43522,N_43523,N_43524,N_43525,N_43526,N_43527,N_43528,N_43529,N_43530,N_43531,N_43532,N_43533,N_43534,N_43535,N_43536,N_43537,N_43538,N_43539,N_43540,N_43541,N_43542,N_43543,N_43544,N_43545,N_43546,N_43547,N_43548,N_43549,N_43550,N_43551,N_43552,N_43553,N_43554,N_43555,N_43556,N_43557,N_43558,N_43559,N_43560,N_43561,N_43562,N_43563,N_43564,N_43565,N_43566,N_43567,N_43568,N_43569,N_43570,N_43571,N_43572,N_43573,N_43574,N_43575,N_43576,N_43577,N_43578,N_43579,N_43580,N_43581,N_43582,N_43583,N_43584,N_43585,N_43586,N_43587,N_43588,N_43589,N_43590,N_43591,N_43592,N_43593,N_43594,N_43595,N_43596,N_43597,N_43598,N_43599,N_43600,N_43601,N_43602,N_43603,N_43604,N_43605,N_43606,N_43607,N_43608,N_43609,N_43610,N_43611,N_43612,N_43613,N_43614,N_43615,N_43616,N_43617,N_43618,N_43619,N_43620,N_43621,N_43622,N_43623,N_43624,N_43625,N_43626,N_43627,N_43628,N_43629,N_43630,N_43631,N_43632,N_43633,N_43634,N_43635,N_43636,N_43637,N_43638,N_43639,N_43640,N_43641,N_43642,N_43643,N_43644,N_43645,N_43646,N_43647,N_43648,N_43649,N_43650,N_43651,N_43652,N_43653,N_43654,N_43655,N_43656,N_43657,N_43658,N_43659,N_43660,N_43661,N_43662,N_43663,N_43664,N_43665,N_43666,N_43667,N_43668,N_43669,N_43670,N_43671,N_43672,N_43673,N_43674,N_43675,N_43676,N_43677,N_43678,N_43679,N_43680,N_43681,N_43682,N_43683,N_43684,N_43685,N_43686,N_43687,N_43688,N_43689,N_43690,N_43691,N_43692,N_43693,N_43694,N_43695,N_43696,N_43697,N_43698,N_43699,N_43700,N_43701,N_43702,N_43703,N_43704,N_43705,N_43706,N_43707,N_43708,N_43709,N_43710,N_43711,N_43712,N_43713,N_43714,N_43715,N_43716,N_43717,N_43718,N_43719,N_43720,N_43721,N_43722,N_43723,N_43724,N_43725,N_43726,N_43727,N_43728,N_43729,N_43730,N_43731,N_43732,N_43733,N_43734,N_43735,N_43736,N_43737,N_43738,N_43739,N_43740,N_43741,N_43742,N_43743,N_43744,N_43745,N_43746,N_43747,N_43748,N_43749,N_43750,N_43751,N_43752,N_43753,N_43754,N_43755,N_43756,N_43757,N_43758,N_43759,N_43760,N_43761,N_43762,N_43763,N_43764,N_43765,N_43766,N_43767,N_43768,N_43769,N_43770,N_43771,N_43772,N_43773,N_43774,N_43775,N_43776,N_43777,N_43778,N_43779,N_43780,N_43781,N_43782,N_43783,N_43784,N_43785,N_43786,N_43787,N_43788,N_43789,N_43790,N_43791,N_43792,N_43793,N_43794,N_43795,N_43796,N_43797,N_43798,N_43799,N_43800,N_43801,N_43802,N_43803,N_43804,N_43805,N_43806,N_43807,N_43808,N_43809,N_43810,N_43811,N_43812,N_43813,N_43814,N_43815,N_43816,N_43817,N_43818,N_43819,N_43820,N_43821,N_43822,N_43823,N_43824,N_43825,N_43826,N_43827,N_43828,N_43829,N_43830,N_43831,N_43832,N_43833,N_43834,N_43835,N_43836,N_43837,N_43838,N_43839,N_43840,N_43841,N_43842,N_43843,N_43844,N_43845,N_43846,N_43847,N_43848,N_43849,N_43850,N_43851,N_43852,N_43853,N_43854,N_43855,N_43856,N_43857,N_43858,N_43859,N_43860,N_43861,N_43862,N_43863,N_43864,N_43865,N_43866,N_43867,N_43868,N_43869,N_43870,N_43871,N_43872,N_43873,N_43874,N_43875,N_43876,N_43877,N_43878,N_43879,N_43880,N_43881,N_43882,N_43883,N_43884,N_43885,N_43886,N_43887,N_43888,N_43889,N_43890,N_43891,N_43892,N_43893,N_43894,N_43895,N_43896,N_43897,N_43898,N_43899,N_43900,N_43901,N_43902,N_43903,N_43904,N_43905,N_43906,N_43907,N_43908,N_43909,N_43910,N_43911,N_43912,N_43913,N_43914,N_43915,N_43916,N_43917,N_43918,N_43919,N_43920,N_43921,N_43922,N_43923,N_43924,N_43925,N_43926,N_43927,N_43928,N_43929,N_43930,N_43931,N_43932,N_43933,N_43934,N_43935,N_43936,N_43937,N_43938,N_43939,N_43940,N_43941,N_43942,N_43943,N_43944,N_43945,N_43946,N_43947,N_43948,N_43949,N_43950,N_43951,N_43952,N_43953,N_43954,N_43955,N_43956,N_43957,N_43958,N_43959,N_43960,N_43961,N_43962,N_43963,N_43964,N_43965,N_43966,N_43967,N_43968,N_43969,N_43970,N_43971,N_43972,N_43973,N_43974,N_43975,N_43976,N_43977,N_43978,N_43979,N_43980,N_43981,N_43982,N_43983,N_43984,N_43985,N_43986,N_43987,N_43988,N_43989,N_43990,N_43991,N_43992,N_43993,N_43994,N_43995,N_43996,N_43997,N_43998,N_43999,N_44000,N_44001,N_44002,N_44003,N_44004,N_44005,N_44006,N_44007,N_44008,N_44009,N_44010,N_44011,N_44012,N_44013,N_44014,N_44015,N_44016,N_44017,N_44018,N_44019,N_44020,N_44021,N_44022,N_44023,N_44024,N_44025,N_44026,N_44027,N_44028,N_44029,N_44030,N_44031,N_44032,N_44033,N_44034,N_44035,N_44036,N_44037,N_44038,N_44039,N_44040,N_44041,N_44042,N_44043,N_44044,N_44045,N_44046,N_44047,N_44048,N_44049,N_44050,N_44051,N_44052,N_44053,N_44054,N_44055,N_44056,N_44057,N_44058,N_44059,N_44060,N_44061,N_44062,N_44063,N_44064,N_44065,N_44066,N_44067,N_44068,N_44069,N_44070,N_44071,N_44072,N_44073,N_44074,N_44075,N_44076,N_44077,N_44078,N_44079,N_44080,N_44081,N_44082,N_44083,N_44084,N_44085,N_44086,N_44087,N_44088,N_44089,N_44090,N_44091,N_44092,N_44093,N_44094,N_44095,N_44096,N_44097,N_44098,N_44099,N_44100,N_44101,N_44102,N_44103,N_44104,N_44105,N_44106,N_44107,N_44108,N_44109,N_44110,N_44111,N_44112,N_44113,N_44114,N_44115,N_44116,N_44117,N_44118,N_44119,N_44120,N_44121,N_44122,N_44123,N_44124,N_44125,N_44126,N_44127,N_44128,N_44129,N_44130,N_44131,N_44132,N_44133,N_44134,N_44135,N_44136,N_44137,N_44138,N_44139,N_44140,N_44141,N_44142,N_44143,N_44144,N_44145,N_44146,N_44147,N_44148,N_44149,N_44150,N_44151,N_44152,N_44153,N_44154,N_44155,N_44156,N_44157,N_44158,N_44159,N_44160,N_44161,N_44162,N_44163,N_44164,N_44165,N_44166,N_44167,N_44168,N_44169,N_44170,N_44171,N_44172,N_44173,N_44174,N_44175,N_44176,N_44177,N_44178,N_44179,N_44180,N_44181,N_44182,N_44183,N_44184,N_44185,N_44186,N_44187,N_44188,N_44189,N_44190,N_44191,N_44192,N_44193,N_44194,N_44195,N_44196,N_44197,N_44198,N_44199,N_44200,N_44201,N_44202,N_44203,N_44204,N_44205,N_44206,N_44207,N_44208,N_44209,N_44210,N_44211,N_44212,N_44213,N_44214,N_44215,N_44216,N_44217,N_44218,N_44219,N_44220,N_44221,N_44222,N_44223,N_44224,N_44225,N_44226,N_44227,N_44228,N_44229,N_44230,N_44231,N_44232,N_44233,N_44234,N_44235,N_44236,N_44237,N_44238,N_44239,N_44240,N_44241,N_44242,N_44243,N_44244,N_44245,N_44246,N_44247,N_44248,N_44249,N_44250,N_44251,N_44252,N_44253,N_44254,N_44255,N_44256,N_44257,N_44258,N_44259,N_44260,N_44261,N_44262,N_44263,N_44264,N_44265,N_44266,N_44267,N_44268,N_44269,N_44270,N_44271,N_44272,N_44273,N_44274,N_44275,N_44276,N_44277,N_44278,N_44279,N_44280,N_44281,N_44282,N_44283,N_44284,N_44285,N_44286,N_44287,N_44288,N_44289,N_44290,N_44291,N_44292,N_44293,N_44294,N_44295,N_44296,N_44297,N_44298,N_44299,N_44300,N_44301,N_44302,N_44303,N_44304,N_44305,N_44306,N_44307,N_44308,N_44309,N_44310,N_44311,N_44312,N_44313,N_44314,N_44315,N_44316,N_44317,N_44318,N_44319,N_44320,N_44321,N_44322,N_44323,N_44324,N_44325,N_44326,N_44327,N_44328,N_44329,N_44330,N_44331,N_44332,N_44333,N_44334,N_44335,N_44336,N_44337,N_44338,N_44339,N_44340,N_44341,N_44342,N_44343,N_44344,N_44345,N_44346,N_44347,N_44348,N_44349,N_44350,N_44351,N_44352,N_44353,N_44354,N_44355,N_44356,N_44357,N_44358,N_44359,N_44360,N_44361,N_44362,N_44363,N_44364,N_44365,N_44366,N_44367,N_44368,N_44369,N_44370,N_44371,N_44372,N_44373,N_44374,N_44375,N_44376,N_44377,N_44378,N_44379,N_44380,N_44381,N_44382,N_44383,N_44384,N_44385,N_44386,N_44387,N_44388,N_44389,N_44390,N_44391,N_44392,N_44393,N_44394,N_44395,N_44396,N_44397,N_44398,N_44399,N_44400,N_44401,N_44402,N_44403,N_44404,N_44405,N_44406,N_44407,N_44408,N_44409,N_44410,N_44411,N_44412,N_44413,N_44414,N_44415,N_44416,N_44417,N_44418,N_44419,N_44420,N_44421,N_44422,N_44423,N_44424,N_44425,N_44426,N_44427,N_44428,N_44429,N_44430,N_44431,N_44432,N_44433,N_44434,N_44435,N_44436,N_44437,N_44438,N_44439,N_44440,N_44441,N_44442,N_44443,N_44444,N_44445,N_44446,N_44447,N_44448,N_44449,N_44450,N_44451,N_44452,N_44453,N_44454,N_44455,N_44456,N_44457,N_44458,N_44459,N_44460,N_44461,N_44462,N_44463,N_44464,N_44465,N_44466,N_44467,N_44468,N_44469,N_44470,N_44471,N_44472,N_44473,N_44474,N_44475,N_44476,N_44477,N_44478,N_44479,N_44480,N_44481,N_44482,N_44483,N_44484,N_44485,N_44486,N_44487,N_44488,N_44489,N_44490,N_44491,N_44492,N_44493,N_44494,N_44495,N_44496,N_44497,N_44498,N_44499,N_44500,N_44501,N_44502,N_44503,N_44504,N_44505,N_44506,N_44507,N_44508,N_44509,N_44510,N_44511,N_44512,N_44513,N_44514,N_44515,N_44516,N_44517,N_44518,N_44519,N_44520,N_44521,N_44522,N_44523,N_44524,N_44525,N_44526,N_44527,N_44528,N_44529,N_44530,N_44531,N_44532,N_44533,N_44534,N_44535,N_44536,N_44537,N_44538,N_44539,N_44540,N_44541,N_44542,N_44543,N_44544,N_44545,N_44546,N_44547,N_44548,N_44549,N_44550,N_44551,N_44552,N_44553,N_44554,N_44555,N_44556,N_44557,N_44558,N_44559,N_44560,N_44561,N_44562,N_44563,N_44564,N_44565,N_44566,N_44567,N_44568,N_44569,N_44570,N_44571,N_44572,N_44573,N_44574,N_44575,N_44576,N_44577,N_44578,N_44579,N_44580,N_44581,N_44582,N_44583,N_44584,N_44585,N_44586,N_44587,N_44588,N_44589,N_44590,N_44591,N_44592,N_44593,N_44594,N_44595,N_44596,N_44597,N_44598,N_44599,N_44600,N_44601,N_44602,N_44603,N_44604,N_44605,N_44606,N_44607,N_44608,N_44609,N_44610,N_44611,N_44612,N_44613,N_44614,N_44615,N_44616,N_44617,N_44618,N_44619,N_44620,N_44621,N_44622,N_44623,N_44624,N_44625,N_44626,N_44627,N_44628,N_44629,N_44630,N_44631,N_44632,N_44633,N_44634,N_44635,N_44636,N_44637,N_44638,N_44639,N_44640,N_44641,N_44642,N_44643,N_44644,N_44645,N_44646,N_44647,N_44648,N_44649,N_44650,N_44651,N_44652,N_44653,N_44654,N_44655,N_44656,N_44657,N_44658,N_44659,N_44660,N_44661,N_44662,N_44663,N_44664,N_44665,N_44666,N_44667,N_44668,N_44669,N_44670,N_44671,N_44672,N_44673,N_44674,N_44675,N_44676,N_44677,N_44678,N_44679,N_44680,N_44681,N_44682,N_44683,N_44684,N_44685,N_44686,N_44687,N_44688,N_44689,N_44690,N_44691,N_44692,N_44693,N_44694,N_44695,N_44696,N_44697,N_44698,N_44699,N_44700,N_44701,N_44702,N_44703,N_44704,N_44705,N_44706,N_44707,N_44708,N_44709,N_44710,N_44711,N_44712,N_44713,N_44714,N_44715,N_44716,N_44717,N_44718,N_44719,N_44720,N_44721,N_44722,N_44723,N_44724,N_44725,N_44726,N_44727,N_44728,N_44729,N_44730,N_44731,N_44732,N_44733,N_44734,N_44735,N_44736,N_44737,N_44738,N_44739,N_44740,N_44741,N_44742,N_44743,N_44744,N_44745,N_44746,N_44747,N_44748,N_44749,N_44750,N_44751,N_44752,N_44753,N_44754,N_44755,N_44756,N_44757,N_44758,N_44759,N_44760,N_44761,N_44762,N_44763,N_44764,N_44765,N_44766,N_44767,N_44768,N_44769,N_44770,N_44771,N_44772,N_44773,N_44774,N_44775,N_44776,N_44777,N_44778,N_44779,N_44780,N_44781,N_44782,N_44783,N_44784,N_44785,N_44786,N_44787,N_44788,N_44789,N_44790,N_44791,N_44792,N_44793,N_44794,N_44795,N_44796,N_44797,N_44798,N_44799,N_44800,N_44801,N_44802,N_44803,N_44804,N_44805,N_44806,N_44807,N_44808,N_44809,N_44810,N_44811,N_44812,N_44813,N_44814,N_44815,N_44816,N_44817,N_44818,N_44819,N_44820,N_44821,N_44822,N_44823,N_44824,N_44825,N_44826,N_44827,N_44828,N_44829,N_44830,N_44831,N_44832,N_44833,N_44834,N_44835,N_44836,N_44837,N_44838,N_44839,N_44840,N_44841,N_44842,N_44843,N_44844,N_44845,N_44846,N_44847,N_44848,N_44849,N_44850,N_44851,N_44852,N_44853,N_44854,N_44855,N_44856,N_44857,N_44858,N_44859,N_44860,N_44861,N_44862,N_44863,N_44864,N_44865,N_44866,N_44867,N_44868,N_44869,N_44870,N_44871,N_44872,N_44873,N_44874,N_44875,N_44876,N_44877,N_44878,N_44879,N_44880,N_44881,N_44882,N_44883,N_44884,N_44885,N_44886,N_44887,N_44888,N_44889,N_44890,N_44891,N_44892,N_44893,N_44894,N_44895,N_44896,N_44897,N_44898,N_44899,N_44900,N_44901,N_44902,N_44903,N_44904,N_44905,N_44906,N_44907,N_44908,N_44909,N_44910,N_44911,N_44912,N_44913,N_44914,N_44915,N_44916,N_44917,N_44918,N_44919,N_44920,N_44921,N_44922,N_44923,N_44924,N_44925,N_44926,N_44927,N_44928,N_44929,N_44930,N_44931,N_44932,N_44933,N_44934,N_44935,N_44936,N_44937,N_44938,N_44939,N_44940,N_44941,N_44942,N_44943,N_44944,N_44945,N_44946,N_44947,N_44948,N_44949,N_44950,N_44951,N_44952,N_44953,N_44954,N_44955,N_44956,N_44957,N_44958,N_44959,N_44960,N_44961,N_44962,N_44963,N_44964,N_44965,N_44966,N_44967,N_44968,N_44969,N_44970,N_44971,N_44972,N_44973,N_44974,N_44975,N_44976,N_44977,N_44978,N_44979,N_44980,N_44981,N_44982,N_44983,N_44984,N_44985,N_44986,N_44987,N_44988,N_44989,N_44990,N_44991,N_44992,N_44993,N_44994,N_44995,N_44996,N_44997,N_44998,N_44999,N_45000,N_45001,N_45002,N_45003,N_45004,N_45005,N_45006,N_45007,N_45008,N_45009,N_45010,N_45011,N_45012,N_45013,N_45014,N_45015,N_45016,N_45017,N_45018,N_45019,N_45020,N_45021,N_45022,N_45023,N_45024,N_45025,N_45026,N_45027,N_45028,N_45029,N_45030,N_45031,N_45032,N_45033,N_45034,N_45035,N_45036,N_45037,N_45038,N_45039,N_45040,N_45041,N_45042,N_45043,N_45044,N_45045,N_45046,N_45047,N_45048,N_45049,N_45050,N_45051,N_45052,N_45053,N_45054,N_45055,N_45056,N_45057,N_45058,N_45059,N_45060,N_45061,N_45062,N_45063,N_45064,N_45065,N_45066,N_45067,N_45068,N_45069,N_45070,N_45071,N_45072,N_45073,N_45074,N_45075,N_45076,N_45077,N_45078,N_45079,N_45080,N_45081,N_45082,N_45083,N_45084,N_45085,N_45086,N_45087,N_45088,N_45089,N_45090,N_45091,N_45092,N_45093,N_45094,N_45095,N_45096,N_45097,N_45098,N_45099,N_45100,N_45101,N_45102,N_45103,N_45104,N_45105,N_45106,N_45107,N_45108,N_45109,N_45110,N_45111,N_45112,N_45113,N_45114,N_45115,N_45116,N_45117,N_45118,N_45119,N_45120,N_45121,N_45122,N_45123,N_45124,N_45125,N_45126,N_45127,N_45128,N_45129,N_45130,N_45131,N_45132,N_45133,N_45134,N_45135,N_45136,N_45137,N_45138,N_45139,N_45140,N_45141,N_45142,N_45143,N_45144,N_45145,N_45146,N_45147,N_45148,N_45149,N_45150,N_45151,N_45152,N_45153,N_45154,N_45155,N_45156,N_45157,N_45158,N_45159,N_45160,N_45161,N_45162,N_45163,N_45164,N_45165,N_45166,N_45167,N_45168,N_45169,N_45170,N_45171,N_45172,N_45173,N_45174,N_45175,N_45176,N_45177,N_45178,N_45179,N_45180,N_45181,N_45182,N_45183,N_45184,N_45185,N_45186,N_45187,N_45188,N_45189,N_45190,N_45191,N_45192,N_45193,N_45194,N_45195,N_45196,N_45197,N_45198,N_45199,N_45200,N_45201,N_45202,N_45203,N_45204,N_45205,N_45206,N_45207,N_45208,N_45209,N_45210,N_45211,N_45212,N_45213,N_45214,N_45215,N_45216,N_45217,N_45218,N_45219,N_45220,N_45221,N_45222,N_45223,N_45224,N_45225,N_45226,N_45227,N_45228,N_45229,N_45230,N_45231,N_45232,N_45233,N_45234,N_45235,N_45236,N_45237,N_45238,N_45239,N_45240,N_45241,N_45242,N_45243,N_45244,N_45245,N_45246,N_45247,N_45248,N_45249,N_45250,N_45251,N_45252,N_45253,N_45254,N_45255,N_45256,N_45257,N_45258,N_45259,N_45260,N_45261,N_45262,N_45263,N_45264,N_45265,N_45266,N_45267,N_45268,N_45269,N_45270,N_45271,N_45272,N_45273,N_45274,N_45275,N_45276,N_45277,N_45278,N_45279,N_45280,N_45281,N_45282,N_45283,N_45284,N_45285,N_45286,N_45287,N_45288,N_45289,N_45290,N_45291,N_45292,N_45293,N_45294,N_45295,N_45296,N_45297,N_45298,N_45299,N_45300,N_45301,N_45302,N_45303,N_45304,N_45305,N_45306,N_45307,N_45308,N_45309,N_45310,N_45311,N_45312,N_45313,N_45314,N_45315,N_45316,N_45317,N_45318,N_45319,N_45320,N_45321,N_45322,N_45323,N_45324,N_45325,N_45326,N_45327,N_45328,N_45329,N_45330,N_45331,N_45332,N_45333,N_45334,N_45335,N_45336,N_45337,N_45338,N_45339,N_45340,N_45341,N_45342,N_45343,N_45344,N_45345,N_45346,N_45347,N_45348,N_45349,N_45350,N_45351,N_45352,N_45353,N_45354,N_45355,N_45356,N_45357,N_45358,N_45359,N_45360,N_45361,N_45362,N_45363,N_45364,N_45365,N_45366,N_45367,N_45368,N_45369,N_45370,N_45371,N_45372,N_45373,N_45374,N_45375,N_45376,N_45377,N_45378,N_45379,N_45380,N_45381,N_45382,N_45383,N_45384,N_45385,N_45386,N_45387,N_45388,N_45389,N_45390,N_45391,N_45392,N_45393,N_45394,N_45395,N_45396,N_45397,N_45398,N_45399,N_45400,N_45401,N_45402,N_45403,N_45404,N_45405,N_45406,N_45407,N_45408,N_45409,N_45410,N_45411,N_45412,N_45413,N_45414,N_45415,N_45416,N_45417,N_45418,N_45419,N_45420,N_45421,N_45422,N_45423,N_45424,N_45425,N_45426,N_45427,N_45428,N_45429,N_45430,N_45431,N_45432,N_45433,N_45434,N_45435,N_45436,N_45437,N_45438,N_45439,N_45440,N_45441,N_45442,N_45443,N_45444,N_45445,N_45446,N_45447,N_45448,N_45449,N_45450,N_45451,N_45452,N_45453,N_45454,N_45455,N_45456,N_45457,N_45458,N_45459,N_45460,N_45461,N_45462,N_45463,N_45464,N_45465,N_45466,N_45467,N_45468,N_45469,N_45470,N_45471,N_45472,N_45473,N_45474,N_45475,N_45476,N_45477,N_45478,N_45479,N_45480,N_45481,N_45482,N_45483,N_45484,N_45485,N_45486,N_45487,N_45488,N_45489,N_45490,N_45491,N_45492,N_45493,N_45494,N_45495,N_45496,N_45497,N_45498,N_45499,N_45500,N_45501,N_45502,N_45503,N_45504,N_45505,N_45506,N_45507,N_45508,N_45509,N_45510,N_45511,N_45512,N_45513,N_45514,N_45515,N_45516,N_45517,N_45518,N_45519,N_45520,N_45521,N_45522,N_45523,N_45524,N_45525,N_45526,N_45527,N_45528,N_45529,N_45530,N_45531,N_45532,N_45533,N_45534,N_45535,N_45536,N_45537,N_45538,N_45539,N_45540,N_45541,N_45542,N_45543,N_45544,N_45545,N_45546,N_45547,N_45548,N_45549,N_45550,N_45551,N_45552,N_45553,N_45554,N_45555,N_45556,N_45557,N_45558,N_45559,N_45560,N_45561,N_45562,N_45563,N_45564,N_45565,N_45566,N_45567,N_45568,N_45569,N_45570,N_45571,N_45572,N_45573,N_45574,N_45575,N_45576,N_45577,N_45578,N_45579,N_45580,N_45581,N_45582,N_45583,N_45584,N_45585,N_45586,N_45587,N_45588,N_45589,N_45590,N_45591,N_45592,N_45593,N_45594,N_45595,N_45596,N_45597,N_45598,N_45599,N_45600,N_45601,N_45602,N_45603,N_45604,N_45605,N_45606,N_45607,N_45608,N_45609,N_45610,N_45611,N_45612,N_45613,N_45614,N_45615,N_45616,N_45617,N_45618,N_45619,N_45620,N_45621,N_45622,N_45623,N_45624,N_45625,N_45626,N_45627,N_45628,N_45629,N_45630,N_45631,N_45632,N_45633,N_45634,N_45635,N_45636,N_45637,N_45638,N_45639,N_45640,N_45641,N_45642,N_45643,N_45644,N_45645,N_45646,N_45647,N_45648,N_45649,N_45650,N_45651,N_45652,N_45653,N_45654,N_45655,N_45656,N_45657,N_45658,N_45659,N_45660,N_45661,N_45662,N_45663,N_45664,N_45665,N_45666,N_45667,N_45668,N_45669,N_45670,N_45671,N_45672,N_45673,N_45674,N_45675,N_45676,N_45677,N_45678,N_45679,N_45680,N_45681,N_45682,N_45683,N_45684,N_45685,N_45686,N_45687,N_45688,N_45689,N_45690,N_45691,N_45692,N_45693,N_45694,N_45695,N_45696,N_45697,N_45698,N_45699,N_45700,N_45701,N_45702,N_45703,N_45704,N_45705,N_45706,N_45707,N_45708,N_45709,N_45710,N_45711,N_45712,N_45713,N_45714,N_45715,N_45716,N_45717,N_45718,N_45719,N_45720,N_45721,N_45722,N_45723,N_45724,N_45725,N_45726,N_45727,N_45728,N_45729,N_45730,N_45731,N_45732,N_45733,N_45734,N_45735,N_45736,N_45737,N_45738,N_45739,N_45740,N_45741,N_45742,N_45743,N_45744,N_45745,N_45746,N_45747,N_45748,N_45749,N_45750,N_45751,N_45752,N_45753,N_45754,N_45755,N_45756,N_45757,N_45758,N_45759,N_45760,N_45761,N_45762,N_45763,N_45764,N_45765,N_45766,N_45767,N_45768,N_45769,N_45770,N_45771,N_45772,N_45773,N_45774,N_45775,N_45776,N_45777,N_45778,N_45779,N_45780,N_45781,N_45782,N_45783,N_45784,N_45785,N_45786,N_45787,N_45788,N_45789,N_45790,N_45791,N_45792,N_45793,N_45794,N_45795,N_45796,N_45797,N_45798,N_45799,N_45800,N_45801,N_45802,N_45803,N_45804,N_45805,N_45806,N_45807,N_45808,N_45809,N_45810,N_45811,N_45812,N_45813,N_45814,N_45815,N_45816,N_45817,N_45818,N_45819,N_45820,N_45821,N_45822,N_45823,N_45824,N_45825,N_45826,N_45827,N_45828,N_45829,N_45830,N_45831,N_45832,N_45833,N_45834,N_45835,N_45836,N_45837,N_45838,N_45839,N_45840,N_45841,N_45842,N_45843,N_45844,N_45845,N_45846,N_45847,N_45848,N_45849,N_45850,N_45851,N_45852,N_45853,N_45854,N_45855,N_45856,N_45857,N_45858,N_45859,N_45860,N_45861,N_45862,N_45863,N_45864,N_45865,N_45866,N_45867,N_45868,N_45869,N_45870,N_45871,N_45872,N_45873,N_45874,N_45875,N_45876,N_45877,N_45878,N_45879,N_45880,N_45881,N_45882,N_45883,N_45884,N_45885,N_45886,N_45887,N_45888,N_45889,N_45890,N_45891,N_45892,N_45893,N_45894,N_45895,N_45896,N_45897,N_45898,N_45899,N_45900,N_45901,N_45902,N_45903,N_45904,N_45905,N_45906,N_45907,N_45908,N_45909,N_45910,N_45911,N_45912,N_45913,N_45914,N_45915,N_45916,N_45917,N_45918,N_45919,N_45920,N_45921,N_45922,N_45923,N_45924,N_45925,N_45926,N_45927,N_45928,N_45929,N_45930,N_45931,N_45932,N_45933,N_45934,N_45935,N_45936,N_45937,N_45938,N_45939,N_45940,N_45941,N_45942,N_45943,N_45944,N_45945,N_45946,N_45947,N_45948,N_45949,N_45950,N_45951,N_45952,N_45953,N_45954,N_45955,N_45956,N_45957,N_45958,N_45959,N_45960,N_45961,N_45962,N_45963,N_45964,N_45965,N_45966,N_45967,N_45968,N_45969,N_45970,N_45971,N_45972,N_45973,N_45974,N_45975,N_45976,N_45977,N_45978,N_45979,N_45980,N_45981,N_45982,N_45983,N_45984,N_45985,N_45986,N_45987,N_45988,N_45989,N_45990,N_45991,N_45992,N_45993,N_45994,N_45995,N_45996,N_45997,N_45998,N_45999,N_46000,N_46001,N_46002,N_46003,N_46004,N_46005,N_46006,N_46007,N_46008,N_46009,N_46010,N_46011,N_46012,N_46013,N_46014,N_46015,N_46016,N_46017,N_46018,N_46019,N_46020,N_46021,N_46022,N_46023,N_46024,N_46025,N_46026,N_46027,N_46028,N_46029,N_46030,N_46031,N_46032,N_46033,N_46034,N_46035,N_46036,N_46037,N_46038,N_46039,N_46040,N_46041,N_46042,N_46043,N_46044,N_46045,N_46046,N_46047,N_46048,N_46049,N_46050,N_46051,N_46052,N_46053,N_46054,N_46055,N_46056,N_46057,N_46058,N_46059,N_46060,N_46061,N_46062,N_46063,N_46064,N_46065,N_46066,N_46067,N_46068,N_46069,N_46070,N_46071,N_46072,N_46073,N_46074,N_46075,N_46076,N_46077,N_46078,N_46079,N_46080,N_46081,N_46082,N_46083,N_46084,N_46085,N_46086,N_46087,N_46088,N_46089,N_46090,N_46091,N_46092,N_46093,N_46094,N_46095,N_46096,N_46097,N_46098,N_46099,N_46100,N_46101,N_46102,N_46103,N_46104,N_46105,N_46106,N_46107,N_46108,N_46109,N_46110,N_46111,N_46112,N_46113,N_46114,N_46115,N_46116,N_46117,N_46118,N_46119,N_46120,N_46121,N_46122,N_46123,N_46124,N_46125,N_46126,N_46127,N_46128,N_46129,N_46130,N_46131,N_46132,N_46133,N_46134,N_46135,N_46136,N_46137,N_46138,N_46139,N_46140,N_46141,N_46142,N_46143,N_46144,N_46145,N_46146,N_46147,N_46148,N_46149,N_46150,N_46151,N_46152,N_46153,N_46154,N_46155,N_46156,N_46157,N_46158,N_46159,N_46160,N_46161,N_46162,N_46163,N_46164,N_46165,N_46166,N_46167,N_46168,N_46169,N_46170,N_46171,N_46172,N_46173,N_46174,N_46175,N_46176,N_46177,N_46178,N_46179,N_46180,N_46181,N_46182,N_46183,N_46184,N_46185,N_46186,N_46187,N_46188,N_46189,N_46190,N_46191,N_46192,N_46193,N_46194,N_46195,N_46196,N_46197,N_46198,N_46199,N_46200,N_46201,N_46202,N_46203,N_46204,N_46205,N_46206,N_46207,N_46208,N_46209,N_46210,N_46211,N_46212,N_46213,N_46214,N_46215,N_46216,N_46217,N_46218,N_46219,N_46220,N_46221,N_46222,N_46223,N_46224,N_46225,N_46226,N_46227,N_46228,N_46229,N_46230,N_46231,N_46232,N_46233,N_46234,N_46235,N_46236,N_46237,N_46238,N_46239,N_46240,N_46241,N_46242,N_46243,N_46244,N_46245,N_46246,N_46247,N_46248,N_46249,N_46250,N_46251,N_46252,N_46253,N_46254,N_46255,N_46256,N_46257,N_46258,N_46259,N_46260,N_46261,N_46262,N_46263,N_46264,N_46265,N_46266,N_46267,N_46268,N_46269,N_46270,N_46271,N_46272,N_46273,N_46274,N_46275,N_46276,N_46277,N_46278,N_46279,N_46280,N_46281,N_46282,N_46283,N_46284,N_46285,N_46286,N_46287,N_46288,N_46289,N_46290,N_46291,N_46292,N_46293,N_46294,N_46295,N_46296,N_46297,N_46298,N_46299,N_46300,N_46301,N_46302,N_46303,N_46304,N_46305,N_46306,N_46307,N_46308,N_46309,N_46310,N_46311,N_46312,N_46313,N_46314,N_46315,N_46316,N_46317,N_46318,N_46319,N_46320,N_46321,N_46322,N_46323,N_46324,N_46325,N_46326,N_46327,N_46328,N_46329,N_46330,N_46331,N_46332,N_46333,N_46334,N_46335,N_46336,N_46337,N_46338,N_46339,N_46340,N_46341,N_46342,N_46343,N_46344,N_46345,N_46346,N_46347,N_46348,N_46349,N_46350,N_46351,N_46352,N_46353,N_46354,N_46355,N_46356,N_46357,N_46358,N_46359,N_46360,N_46361,N_46362,N_46363,N_46364,N_46365,N_46366,N_46367,N_46368,N_46369,N_46370,N_46371,N_46372,N_46373,N_46374,N_46375,N_46376,N_46377,N_46378,N_46379,N_46380,N_46381,N_46382,N_46383,N_46384,N_46385,N_46386,N_46387,N_46388,N_46389,N_46390,N_46391,N_46392,N_46393,N_46394,N_46395,N_46396,N_46397,N_46398,N_46399,N_46400,N_46401,N_46402,N_46403,N_46404,N_46405,N_46406,N_46407,N_46408,N_46409,N_46410,N_46411,N_46412,N_46413,N_46414,N_46415,N_46416,N_46417,N_46418,N_46419,N_46420,N_46421,N_46422,N_46423,N_46424,N_46425,N_46426,N_46427,N_46428,N_46429,N_46430,N_46431,N_46432,N_46433,N_46434,N_46435,N_46436,N_46437,N_46438,N_46439,N_46440,N_46441,N_46442,N_46443,N_46444,N_46445,N_46446,N_46447,N_46448,N_46449,N_46450,N_46451,N_46452,N_46453,N_46454,N_46455,N_46456,N_46457,N_46458,N_46459,N_46460,N_46461,N_46462,N_46463,N_46464,N_46465,N_46466,N_46467,N_46468,N_46469,N_46470,N_46471,N_46472,N_46473,N_46474,N_46475,N_46476,N_46477,N_46478,N_46479,N_46480,N_46481,N_46482,N_46483,N_46484,N_46485,N_46486,N_46487,N_46488,N_46489,N_46490,N_46491,N_46492,N_46493,N_46494,N_46495,N_46496,N_46497,N_46498,N_46499,N_46500,N_46501,N_46502,N_46503,N_46504,N_46505,N_46506,N_46507,N_46508,N_46509,N_46510,N_46511,N_46512,N_46513,N_46514,N_46515,N_46516,N_46517,N_46518,N_46519,N_46520,N_46521,N_46522,N_46523,N_46524,N_46525,N_46526,N_46527,N_46528,N_46529,N_46530,N_46531,N_46532,N_46533,N_46534,N_46535,N_46536,N_46537,N_46538,N_46539,N_46540,N_46541,N_46542,N_46543,N_46544,N_46545,N_46546,N_46547,N_46548,N_46549,N_46550,N_46551,N_46552,N_46553,N_46554,N_46555,N_46556,N_46557,N_46558,N_46559,N_46560,N_46561,N_46562,N_46563,N_46564,N_46565,N_46566,N_46567,N_46568,N_46569,N_46570,N_46571,N_46572,N_46573,N_46574,N_46575,N_46576,N_46577,N_46578,N_46579,N_46580,N_46581,N_46582,N_46583,N_46584,N_46585,N_46586,N_46587,N_46588,N_46589,N_46590,N_46591,N_46592,N_46593,N_46594,N_46595,N_46596,N_46597,N_46598,N_46599,N_46600,N_46601,N_46602,N_46603,N_46604,N_46605,N_46606,N_46607,N_46608,N_46609,N_46610,N_46611,N_46612,N_46613,N_46614,N_46615,N_46616,N_46617,N_46618,N_46619,N_46620,N_46621,N_46622,N_46623,N_46624,N_46625,N_46626,N_46627,N_46628,N_46629,N_46630,N_46631,N_46632,N_46633,N_46634,N_46635,N_46636,N_46637,N_46638,N_46639,N_46640,N_46641,N_46642,N_46643,N_46644,N_46645,N_46646,N_46647,N_46648,N_46649,N_46650,N_46651,N_46652,N_46653,N_46654,N_46655,N_46656,N_46657,N_46658,N_46659,N_46660,N_46661,N_46662,N_46663,N_46664,N_46665,N_46666,N_46667,N_46668,N_46669,N_46670,N_46671,N_46672,N_46673,N_46674,N_46675,N_46676,N_46677,N_46678,N_46679,N_46680,N_46681,N_46682,N_46683,N_46684,N_46685,N_46686,N_46687,N_46688,N_46689,N_46690,N_46691,N_46692,N_46693,N_46694,N_46695,N_46696,N_46697,N_46698,N_46699,N_46700,N_46701,N_46702,N_46703,N_46704,N_46705,N_46706,N_46707,N_46708,N_46709,N_46710,N_46711,N_46712,N_46713,N_46714,N_46715,N_46716,N_46717,N_46718,N_46719,N_46720,N_46721,N_46722,N_46723,N_46724,N_46725,N_46726,N_46727,N_46728,N_46729,N_46730,N_46731,N_46732,N_46733,N_46734,N_46735,N_46736,N_46737,N_46738,N_46739,N_46740,N_46741,N_46742,N_46743,N_46744,N_46745,N_46746,N_46747,N_46748,N_46749,N_46750,N_46751,N_46752,N_46753,N_46754,N_46755,N_46756,N_46757,N_46758,N_46759,N_46760,N_46761,N_46762,N_46763,N_46764,N_46765,N_46766,N_46767,N_46768,N_46769,N_46770,N_46771,N_46772,N_46773,N_46774,N_46775,N_46776,N_46777,N_46778,N_46779,N_46780,N_46781,N_46782,N_46783,N_46784,N_46785,N_46786,N_46787,N_46788,N_46789,N_46790,N_46791,N_46792,N_46793,N_46794,N_46795,N_46796,N_46797,N_46798,N_46799,N_46800,N_46801,N_46802,N_46803,N_46804,N_46805,N_46806,N_46807,N_46808,N_46809,N_46810,N_46811,N_46812,N_46813,N_46814,N_46815,N_46816,N_46817,N_46818,N_46819,N_46820,N_46821,N_46822,N_46823,N_46824,N_46825,N_46826,N_46827,N_46828,N_46829,N_46830,N_46831,N_46832,N_46833,N_46834,N_46835,N_46836,N_46837,N_46838,N_46839,N_46840,N_46841,N_46842,N_46843,N_46844,N_46845,N_46846,N_46847,N_46848,N_46849,N_46850,N_46851,N_46852,N_46853,N_46854,N_46855,N_46856,N_46857,N_46858,N_46859,N_46860,N_46861,N_46862,N_46863,N_46864,N_46865,N_46866,N_46867,N_46868,N_46869,N_46870,N_46871,N_46872,N_46873,N_46874,N_46875,N_46876,N_46877,N_46878,N_46879,N_46880,N_46881,N_46882,N_46883,N_46884,N_46885,N_46886,N_46887,N_46888,N_46889,N_46890,N_46891,N_46892,N_46893,N_46894,N_46895,N_46896,N_46897,N_46898,N_46899,N_46900,N_46901,N_46902,N_46903,N_46904,N_46905,N_46906,N_46907,N_46908,N_46909,N_46910,N_46911,N_46912,N_46913,N_46914,N_46915,N_46916,N_46917,N_46918,N_46919,N_46920,N_46921,N_46922,N_46923,N_46924,N_46925,N_46926,N_46927,N_46928,N_46929,N_46930,N_46931,N_46932,N_46933,N_46934,N_46935,N_46936,N_46937,N_46938,N_46939,N_46940,N_46941,N_46942,N_46943,N_46944,N_46945,N_46946,N_46947,N_46948,N_46949,N_46950,N_46951,N_46952,N_46953,N_46954,N_46955,N_46956,N_46957,N_46958,N_46959,N_46960,N_46961,N_46962,N_46963,N_46964,N_46965,N_46966,N_46967,N_46968,N_46969,N_46970,N_46971,N_46972,N_46973,N_46974,N_46975,N_46976,N_46977,N_46978,N_46979,N_46980,N_46981,N_46982,N_46983,N_46984,N_46985,N_46986,N_46987,N_46988,N_46989,N_46990,N_46991,N_46992,N_46993,N_46994,N_46995,N_46996,N_46997,N_46998,N_46999,N_47000,N_47001,N_47002,N_47003,N_47004,N_47005,N_47006,N_47007,N_47008,N_47009,N_47010,N_47011,N_47012,N_47013,N_47014,N_47015,N_47016,N_47017,N_47018,N_47019,N_47020,N_47021,N_47022,N_47023,N_47024,N_47025,N_47026,N_47027,N_47028,N_47029,N_47030,N_47031,N_47032,N_47033,N_47034,N_47035,N_47036,N_47037,N_47038,N_47039,N_47040,N_47041,N_47042,N_47043,N_47044,N_47045,N_47046,N_47047,N_47048,N_47049,N_47050,N_47051,N_47052,N_47053,N_47054,N_47055,N_47056,N_47057,N_47058,N_47059,N_47060,N_47061,N_47062,N_47063,N_47064,N_47065,N_47066,N_47067,N_47068,N_47069,N_47070,N_47071,N_47072,N_47073,N_47074,N_47075,N_47076,N_47077,N_47078,N_47079,N_47080,N_47081,N_47082,N_47083,N_47084,N_47085,N_47086,N_47087,N_47088,N_47089,N_47090,N_47091,N_47092,N_47093,N_47094,N_47095,N_47096,N_47097,N_47098,N_47099,N_47100,N_47101,N_47102,N_47103,N_47104,N_47105,N_47106,N_47107,N_47108,N_47109,N_47110,N_47111,N_47112,N_47113,N_47114,N_47115,N_47116,N_47117,N_47118,N_47119,N_47120,N_47121,N_47122,N_47123,N_47124,N_47125,N_47126,N_47127,N_47128,N_47129,N_47130,N_47131,N_47132,N_47133,N_47134,N_47135,N_47136,N_47137,N_47138,N_47139,N_47140,N_47141,N_47142,N_47143,N_47144,N_47145,N_47146,N_47147,N_47148,N_47149,N_47150,N_47151,N_47152,N_47153,N_47154,N_47155,N_47156,N_47157,N_47158,N_47159,N_47160,N_47161,N_47162,N_47163,N_47164,N_47165,N_47166,N_47167,N_47168,N_47169,N_47170,N_47171,N_47172,N_47173,N_47174,N_47175,N_47176,N_47177,N_47178,N_47179,N_47180,N_47181,N_47182,N_47183,N_47184,N_47185,N_47186,N_47187,N_47188,N_47189,N_47190,N_47191,N_47192,N_47193,N_47194,N_47195,N_47196,N_47197,N_47198,N_47199,N_47200,N_47201,N_47202,N_47203,N_47204,N_47205,N_47206,N_47207,N_47208,N_47209,N_47210,N_47211,N_47212,N_47213,N_47214,N_47215,N_47216,N_47217,N_47218,N_47219,N_47220,N_47221,N_47222,N_47223,N_47224,N_47225,N_47226,N_47227,N_47228,N_47229,N_47230,N_47231,N_47232,N_47233,N_47234,N_47235,N_47236,N_47237,N_47238,N_47239,N_47240,N_47241,N_47242,N_47243,N_47244,N_47245,N_47246,N_47247,N_47248,N_47249,N_47250,N_47251,N_47252,N_47253,N_47254,N_47255,N_47256,N_47257,N_47258,N_47259,N_47260,N_47261,N_47262,N_47263,N_47264,N_47265,N_47266,N_47267,N_47268,N_47269,N_47270,N_47271,N_47272,N_47273,N_47274,N_47275,N_47276,N_47277,N_47278,N_47279,N_47280,N_47281,N_47282,N_47283,N_47284,N_47285,N_47286,N_47287,N_47288,N_47289,N_47290,N_47291,N_47292,N_47293,N_47294,N_47295,N_47296,N_47297,N_47298,N_47299,N_47300,N_47301,N_47302,N_47303,N_47304,N_47305,N_47306,N_47307,N_47308,N_47309,N_47310,N_47311,N_47312,N_47313,N_47314,N_47315,N_47316,N_47317,N_47318,N_47319,N_47320,N_47321,N_47322,N_47323,N_47324,N_47325,N_47326,N_47327,N_47328,N_47329,N_47330,N_47331,N_47332,N_47333,N_47334,N_47335,N_47336,N_47337,N_47338,N_47339,N_47340,N_47341,N_47342,N_47343,N_47344,N_47345,N_47346,N_47347,N_47348,N_47349,N_47350,N_47351,N_47352,N_47353,N_47354,N_47355,N_47356,N_47357,N_47358,N_47359,N_47360,N_47361,N_47362,N_47363,N_47364,N_47365,N_47366,N_47367,N_47368,N_47369,N_47370,N_47371,N_47372,N_47373,N_47374,N_47375,N_47376,N_47377,N_47378,N_47379,N_47380,N_47381,N_47382,N_47383,N_47384,N_47385,N_47386,N_47387,N_47388,N_47389,N_47390,N_47391,N_47392,N_47393,N_47394,N_47395,N_47396,N_47397,N_47398,N_47399,N_47400,N_47401,N_47402,N_47403,N_47404,N_47405,N_47406,N_47407,N_47408,N_47409,N_47410,N_47411,N_47412,N_47413,N_47414,N_47415,N_47416,N_47417,N_47418,N_47419,N_47420,N_47421,N_47422,N_47423,N_47424,N_47425,N_47426,N_47427,N_47428,N_47429,N_47430,N_47431,N_47432,N_47433,N_47434,N_47435,N_47436,N_47437,N_47438,N_47439,N_47440,N_47441,N_47442,N_47443,N_47444,N_47445,N_47446,N_47447,N_47448,N_47449,N_47450,N_47451,N_47452,N_47453,N_47454,N_47455,N_47456,N_47457,N_47458,N_47459,N_47460,N_47461,N_47462,N_47463,N_47464,N_47465,N_47466,N_47467,N_47468,N_47469,N_47470,N_47471,N_47472,N_47473,N_47474,N_47475,N_47476,N_47477,N_47478,N_47479,N_47480,N_47481,N_47482,N_47483,N_47484,N_47485,N_47486,N_47487,N_47488,N_47489,N_47490,N_47491,N_47492,N_47493,N_47494,N_47495,N_47496,N_47497,N_47498,N_47499,N_47500,N_47501,N_47502,N_47503,N_47504,N_47505,N_47506,N_47507,N_47508,N_47509,N_47510,N_47511,N_47512,N_47513,N_47514,N_47515,N_47516,N_47517,N_47518,N_47519,N_47520,N_47521,N_47522,N_47523,N_47524,N_47525,N_47526,N_47527,N_47528,N_47529,N_47530,N_47531,N_47532,N_47533,N_47534,N_47535,N_47536,N_47537,N_47538,N_47539,N_47540,N_47541,N_47542,N_47543,N_47544,N_47545,N_47546,N_47547,N_47548,N_47549,N_47550,N_47551,N_47552,N_47553,N_47554,N_47555,N_47556,N_47557,N_47558,N_47559,N_47560,N_47561,N_47562,N_47563,N_47564,N_47565,N_47566,N_47567,N_47568,N_47569,N_47570,N_47571,N_47572,N_47573,N_47574,N_47575,N_47576,N_47577,N_47578,N_47579,N_47580,N_47581,N_47582,N_47583,N_47584,N_47585,N_47586,N_47587,N_47588,N_47589,N_47590,N_47591,N_47592,N_47593,N_47594,N_47595,N_47596,N_47597,N_47598,N_47599,N_47600,N_47601,N_47602,N_47603,N_47604,N_47605,N_47606,N_47607,N_47608,N_47609,N_47610,N_47611,N_47612,N_47613,N_47614,N_47615,N_47616,N_47617,N_47618,N_47619,N_47620,N_47621,N_47622,N_47623,N_47624,N_47625,N_47626,N_47627,N_47628,N_47629,N_47630,N_47631,N_47632,N_47633,N_47634,N_47635,N_47636,N_47637,N_47638,N_47639,N_47640,N_47641,N_47642,N_47643,N_47644,N_47645,N_47646,N_47647,N_47648,N_47649,N_47650,N_47651,N_47652,N_47653,N_47654,N_47655,N_47656,N_47657,N_47658,N_47659,N_47660,N_47661,N_47662,N_47663,N_47664,N_47665,N_47666,N_47667,N_47668,N_47669,N_47670,N_47671,N_47672,N_47673,N_47674,N_47675,N_47676,N_47677,N_47678,N_47679,N_47680,N_47681,N_47682,N_47683,N_47684,N_47685,N_47686,N_47687,N_47688,N_47689,N_47690,N_47691,N_47692,N_47693,N_47694,N_47695,N_47696,N_47697,N_47698,N_47699,N_47700,N_47701,N_47702,N_47703,N_47704,N_47705,N_47706,N_47707,N_47708,N_47709,N_47710,N_47711,N_47712,N_47713,N_47714,N_47715,N_47716,N_47717,N_47718,N_47719,N_47720,N_47721,N_47722,N_47723,N_47724,N_47725,N_47726,N_47727,N_47728,N_47729,N_47730,N_47731,N_47732,N_47733,N_47734,N_47735,N_47736,N_47737,N_47738,N_47739,N_47740,N_47741,N_47742,N_47743,N_47744,N_47745,N_47746,N_47747,N_47748,N_47749,N_47750,N_47751,N_47752,N_47753,N_47754,N_47755,N_47756,N_47757,N_47758,N_47759,N_47760,N_47761,N_47762,N_47763,N_47764,N_47765,N_47766,N_47767,N_47768,N_47769,N_47770,N_47771,N_47772,N_47773,N_47774,N_47775,N_47776,N_47777,N_47778,N_47779,N_47780,N_47781,N_47782,N_47783,N_47784,N_47785,N_47786,N_47787,N_47788,N_47789,N_47790,N_47791,N_47792,N_47793,N_47794,N_47795,N_47796,N_47797,N_47798,N_47799,N_47800,N_47801,N_47802,N_47803,N_47804,N_47805,N_47806,N_47807,N_47808,N_47809,N_47810,N_47811,N_47812,N_47813,N_47814,N_47815,N_47816,N_47817,N_47818,N_47819,N_47820,N_47821,N_47822,N_47823,N_47824,N_47825,N_47826,N_47827,N_47828,N_47829,N_47830,N_47831,N_47832,N_47833,N_47834,N_47835,N_47836,N_47837,N_47838,N_47839,N_47840,N_47841,N_47842,N_47843,N_47844,N_47845,N_47846,N_47847,N_47848,N_47849,N_47850,N_47851,N_47852,N_47853,N_47854,N_47855,N_47856,N_47857,N_47858,N_47859,N_47860,N_47861,N_47862,N_47863,N_47864,N_47865,N_47866,N_47867,N_47868,N_47869,N_47870,N_47871,N_47872,N_47873,N_47874,N_47875,N_47876,N_47877,N_47878,N_47879,N_47880,N_47881,N_47882,N_47883,N_47884,N_47885,N_47886,N_47887,N_47888,N_47889,N_47890,N_47891,N_47892,N_47893,N_47894,N_47895,N_47896,N_47897,N_47898,N_47899,N_47900,N_47901,N_47902,N_47903,N_47904,N_47905,N_47906,N_47907,N_47908,N_47909,N_47910,N_47911,N_47912,N_47913,N_47914,N_47915,N_47916,N_47917,N_47918,N_47919,N_47920,N_47921,N_47922,N_47923,N_47924,N_47925,N_47926,N_47927,N_47928,N_47929,N_47930,N_47931,N_47932,N_47933,N_47934,N_47935,N_47936,N_47937,N_47938,N_47939,N_47940,N_47941,N_47942,N_47943,N_47944,N_47945,N_47946,N_47947,N_47948,N_47949,N_47950,N_47951,N_47952,N_47953,N_47954,N_47955,N_47956,N_47957,N_47958,N_47959,N_47960,N_47961,N_47962,N_47963,N_47964,N_47965,N_47966,N_47967,N_47968,N_47969,N_47970,N_47971,N_47972,N_47973,N_47974,N_47975,N_47976,N_47977,N_47978,N_47979,N_47980,N_47981,N_47982,N_47983,N_47984,N_47985,N_47986,N_47987,N_47988,N_47989,N_47990,N_47991,N_47992,N_47993,N_47994,N_47995,N_47996,N_47997,N_47998,N_47999,N_48000,N_48001,N_48002,N_48003,N_48004,N_48005,N_48006,N_48007,N_48008,N_48009,N_48010,N_48011,N_48012,N_48013,N_48014,N_48015,N_48016,N_48017,N_48018,N_48019,N_48020,N_48021,N_48022,N_48023,N_48024,N_48025,N_48026,N_48027,N_48028,N_48029,N_48030,N_48031,N_48032,N_48033,N_48034,N_48035,N_48036,N_48037,N_48038,N_48039,N_48040,N_48041,N_48042,N_48043,N_48044,N_48045,N_48046,N_48047,N_48048,N_48049,N_48050,N_48051,N_48052,N_48053,N_48054,N_48055,N_48056,N_48057,N_48058,N_48059,N_48060,N_48061,N_48062,N_48063,N_48064,N_48065,N_48066,N_48067,N_48068,N_48069,N_48070,N_48071,N_48072,N_48073,N_48074,N_48075,N_48076,N_48077,N_48078,N_48079,N_48080,N_48081,N_48082,N_48083,N_48084,N_48085,N_48086,N_48087,N_48088,N_48089,N_48090,N_48091,N_48092,N_48093,N_48094,N_48095,N_48096,N_48097,N_48098,N_48099,N_48100,N_48101,N_48102,N_48103,N_48104,N_48105,N_48106,N_48107,N_48108,N_48109,N_48110,N_48111,N_48112,N_48113,N_48114,N_48115,N_48116,N_48117,N_48118,N_48119,N_48120,N_48121,N_48122,N_48123,N_48124,N_48125,N_48126,N_48127,N_48128,N_48129,N_48130,N_48131,N_48132,N_48133,N_48134,N_48135,N_48136,N_48137,N_48138,N_48139,N_48140,N_48141,N_48142,N_48143,N_48144,N_48145,N_48146,N_48147,N_48148,N_48149,N_48150,N_48151,N_48152,N_48153,N_48154,N_48155,N_48156,N_48157,N_48158,N_48159,N_48160,N_48161,N_48162,N_48163,N_48164,N_48165,N_48166,N_48167,N_48168,N_48169,N_48170,N_48171,N_48172,N_48173,N_48174,N_48175,N_48176,N_48177,N_48178,N_48179,N_48180,N_48181,N_48182,N_48183,N_48184,N_48185,N_48186,N_48187,N_48188,N_48189,N_48190,N_48191,N_48192,N_48193,N_48194,N_48195,N_48196,N_48197,N_48198,N_48199,N_48200,N_48201,N_48202,N_48203,N_48204,N_48205,N_48206,N_48207,N_48208,N_48209,N_48210,N_48211,N_48212,N_48213,N_48214,N_48215,N_48216,N_48217,N_48218,N_48219,N_48220,N_48221,N_48222,N_48223,N_48224,N_48225,N_48226,N_48227,N_48228,N_48229,N_48230,N_48231,N_48232,N_48233,N_48234,N_48235,N_48236,N_48237,N_48238,N_48239,N_48240,N_48241,N_48242,N_48243,N_48244,N_48245,N_48246,N_48247,N_48248,N_48249,N_48250,N_48251,N_48252,N_48253,N_48254,N_48255,N_48256,N_48257,N_48258,N_48259,N_48260,N_48261,N_48262,N_48263,N_48264,N_48265,N_48266,N_48267,N_48268,N_48269,N_48270,N_48271,N_48272,N_48273,N_48274,N_48275,N_48276,N_48277,N_48278,N_48279,N_48280,N_48281,N_48282,N_48283,N_48284,N_48285,N_48286,N_48287,N_48288,N_48289,N_48290,N_48291,N_48292,N_48293,N_48294,N_48295,N_48296,N_48297,N_48298,N_48299,N_48300,N_48301,N_48302,N_48303,N_48304,N_48305,N_48306,N_48307,N_48308,N_48309,N_48310,N_48311,N_48312,N_48313,N_48314,N_48315,N_48316,N_48317,N_48318,N_48319,N_48320,N_48321,N_48322,N_48323,N_48324,N_48325,N_48326,N_48327,N_48328,N_48329,N_48330,N_48331,N_48332,N_48333,N_48334,N_48335,N_48336,N_48337,N_48338,N_48339,N_48340,N_48341,N_48342,N_48343,N_48344,N_48345,N_48346,N_48347,N_48348,N_48349,N_48350,N_48351,N_48352,N_48353,N_48354,N_48355,N_48356,N_48357,N_48358,N_48359,N_48360,N_48361,N_48362,N_48363,N_48364,N_48365,N_48366,N_48367,N_48368,N_48369,N_48370,N_48371,N_48372,N_48373,N_48374,N_48375,N_48376,N_48377,N_48378,N_48379,N_48380,N_48381,N_48382,N_48383,N_48384,N_48385,N_48386,N_48387,N_48388,N_48389,N_48390,N_48391,N_48392,N_48393,N_48394,N_48395,N_48396,N_48397,N_48398,N_48399,N_48400,N_48401,N_48402,N_48403,N_48404,N_48405,N_48406,N_48407,N_48408,N_48409,N_48410,N_48411,N_48412,N_48413,N_48414,N_48415,N_48416,N_48417,N_48418,N_48419,N_48420,N_48421,N_48422,N_48423,N_48424,N_48425,N_48426,N_48427,N_48428,N_48429,N_48430,N_48431,N_48432,N_48433,N_48434,N_48435,N_48436,N_48437,N_48438,N_48439,N_48440,N_48441,N_48442,N_48443,N_48444,N_48445,N_48446,N_48447,N_48448,N_48449,N_48450,N_48451,N_48452,N_48453,N_48454,N_48455,N_48456,N_48457,N_48458,N_48459,N_48460,N_48461,N_48462,N_48463,N_48464,N_48465,N_48466,N_48467,N_48468,N_48469,N_48470,N_48471,N_48472,N_48473,N_48474,N_48475,N_48476,N_48477,N_48478,N_48479,N_48480,N_48481,N_48482,N_48483,N_48484,N_48485,N_48486,N_48487,N_48488,N_48489,N_48490,N_48491,N_48492,N_48493,N_48494,N_48495,N_48496,N_48497,N_48498,N_48499,N_48500,N_48501,N_48502,N_48503,N_48504,N_48505,N_48506,N_48507,N_48508,N_48509,N_48510,N_48511,N_48512,N_48513,N_48514,N_48515,N_48516,N_48517,N_48518,N_48519,N_48520,N_48521,N_48522,N_48523,N_48524,N_48525,N_48526,N_48527,N_48528,N_48529,N_48530,N_48531,N_48532,N_48533,N_48534,N_48535,N_48536,N_48537,N_48538,N_48539,N_48540,N_48541,N_48542,N_48543,N_48544,N_48545,N_48546,N_48547,N_48548,N_48549,N_48550,N_48551,N_48552,N_48553,N_48554,N_48555,N_48556,N_48557,N_48558,N_48559,N_48560,N_48561,N_48562,N_48563,N_48564,N_48565,N_48566,N_48567,N_48568,N_48569,N_48570,N_48571,N_48572,N_48573,N_48574,N_48575,N_48576,N_48577,N_48578,N_48579,N_48580,N_48581,N_48582,N_48583,N_48584,N_48585,N_48586,N_48587,N_48588,N_48589,N_48590,N_48591,N_48592,N_48593,N_48594,N_48595,N_48596,N_48597,N_48598,N_48599,N_48600,N_48601,N_48602,N_48603,N_48604,N_48605,N_48606,N_48607,N_48608,N_48609,N_48610,N_48611,N_48612,N_48613,N_48614,N_48615,N_48616,N_48617,N_48618,N_48619,N_48620,N_48621,N_48622,N_48623,N_48624,N_48625,N_48626,N_48627,N_48628,N_48629,N_48630,N_48631,N_48632,N_48633,N_48634,N_48635,N_48636,N_48637,N_48638,N_48639,N_48640,N_48641,N_48642,N_48643,N_48644,N_48645,N_48646,N_48647,N_48648,N_48649,N_48650,N_48651,N_48652,N_48653,N_48654,N_48655,N_48656,N_48657,N_48658,N_48659,N_48660,N_48661,N_48662,N_48663,N_48664,N_48665,N_48666,N_48667,N_48668,N_48669,N_48670,N_48671,N_48672,N_48673,N_48674,N_48675,N_48676,N_48677,N_48678,N_48679,N_48680,N_48681,N_48682,N_48683,N_48684,N_48685,N_48686,N_48687,N_48688,N_48689,N_48690,N_48691,N_48692,N_48693,N_48694,N_48695,N_48696,N_48697,N_48698,N_48699,N_48700,N_48701,N_48702,N_48703,N_48704,N_48705,N_48706,N_48707,N_48708,N_48709,N_48710,N_48711,N_48712,N_48713,N_48714,N_48715,N_48716,N_48717,N_48718,N_48719,N_48720,N_48721,N_48722,N_48723,N_48724,N_48725,N_48726,N_48727,N_48728,N_48729,N_48730,N_48731,N_48732,N_48733,N_48734,N_48735,N_48736,N_48737,N_48738,N_48739,N_48740,N_48741,N_48742,N_48743,N_48744,N_48745,N_48746,N_48747,N_48748,N_48749,N_48750,N_48751,N_48752,N_48753,N_48754,N_48755,N_48756,N_48757,N_48758,N_48759,N_48760,N_48761,N_48762,N_48763,N_48764,N_48765,N_48766,N_48767,N_48768,N_48769,N_48770,N_48771,N_48772,N_48773,N_48774,N_48775,N_48776,N_48777,N_48778,N_48779,N_48780,N_48781,N_48782,N_48783,N_48784,N_48785,N_48786,N_48787,N_48788,N_48789,N_48790,N_48791,N_48792,N_48793,N_48794,N_48795,N_48796,N_48797,N_48798,N_48799,N_48800,N_48801,N_48802,N_48803,N_48804,N_48805,N_48806,N_48807,N_48808,N_48809,N_48810,N_48811,N_48812,N_48813,N_48814,N_48815,N_48816,N_48817,N_48818,N_48819,N_48820,N_48821,N_48822,N_48823,N_48824,N_48825,N_48826,N_48827,N_48828,N_48829,N_48830,N_48831,N_48832,N_48833,N_48834,N_48835,N_48836,N_48837,N_48838,N_48839,N_48840,N_48841,N_48842,N_48843,N_48844,N_48845,N_48846,N_48847,N_48848,N_48849,N_48850,N_48851,N_48852,N_48853,N_48854,N_48855,N_48856,N_48857,N_48858,N_48859,N_48860,N_48861,N_48862,N_48863,N_48864,N_48865,N_48866,N_48867,N_48868,N_48869,N_48870,N_48871,N_48872,N_48873,N_48874,N_48875,N_48876,N_48877,N_48878,N_48879,N_48880,N_48881,N_48882,N_48883,N_48884,N_48885,N_48886,N_48887,N_48888,N_48889,N_48890,N_48891,N_48892,N_48893,N_48894,N_48895,N_48896,N_48897,N_48898,N_48899,N_48900,N_48901,N_48902,N_48903,N_48904,N_48905,N_48906,N_48907,N_48908,N_48909,N_48910,N_48911,N_48912,N_48913,N_48914,N_48915,N_48916,N_48917,N_48918,N_48919,N_48920,N_48921,N_48922,N_48923,N_48924,N_48925,N_48926,N_48927,N_48928,N_48929,N_48930,N_48931,N_48932,N_48933,N_48934,N_48935,N_48936,N_48937,N_48938,N_48939,N_48940,N_48941,N_48942,N_48943,N_48944,N_48945,N_48946,N_48947,N_48948,N_48949,N_48950,N_48951,N_48952,N_48953,N_48954,N_48955,N_48956,N_48957,N_48958,N_48959,N_48960,N_48961,N_48962,N_48963,N_48964,N_48965,N_48966,N_48967,N_48968,N_48969,N_48970,N_48971,N_48972,N_48973,N_48974,N_48975,N_48976,N_48977,N_48978,N_48979,N_48980,N_48981,N_48982,N_48983,N_48984,N_48985,N_48986,N_48987,N_48988,N_48989,N_48990,N_48991,N_48992,N_48993,N_48994,N_48995,N_48996,N_48997,N_48998,N_48999,N_49000,N_49001,N_49002,N_49003,N_49004,N_49005,N_49006,N_49007,N_49008,N_49009,N_49010,N_49011,N_49012,N_49013,N_49014,N_49015,N_49016,N_49017,N_49018,N_49019,N_49020,N_49021,N_49022,N_49023,N_49024,N_49025,N_49026,N_49027,N_49028,N_49029,N_49030,N_49031,N_49032,N_49033,N_49034,N_49035,N_49036,N_49037,N_49038,N_49039,N_49040,N_49041,N_49042,N_49043,N_49044,N_49045,N_49046,N_49047,N_49048,N_49049,N_49050,N_49051,N_49052,N_49053,N_49054,N_49055,N_49056,N_49057,N_49058,N_49059,N_49060,N_49061,N_49062,N_49063,N_49064,N_49065,N_49066,N_49067,N_49068,N_49069,N_49070,N_49071,N_49072,N_49073,N_49074,N_49075,N_49076,N_49077,N_49078,N_49079,N_49080,N_49081,N_49082,N_49083,N_49084,N_49085,N_49086,N_49087,N_49088,N_49089,N_49090,N_49091,N_49092,N_49093,N_49094,N_49095,N_49096,N_49097,N_49098,N_49099,N_49100,N_49101,N_49102,N_49103,N_49104,N_49105,N_49106,N_49107,N_49108,N_49109,N_49110,N_49111,N_49112,N_49113,N_49114,N_49115,N_49116,N_49117,N_49118,N_49119,N_49120,N_49121,N_49122,N_49123,N_49124,N_49125,N_49126,N_49127,N_49128,N_49129,N_49130,N_49131,N_49132,N_49133,N_49134,N_49135,N_49136,N_49137,N_49138,N_49139,N_49140,N_49141,N_49142,N_49143,N_49144,N_49145,N_49146,N_49147,N_49148,N_49149,N_49150,N_49151,N_49152,N_49153,N_49154,N_49155,N_49156,N_49157,N_49158,N_49159,N_49160,N_49161,N_49162,N_49163,N_49164,N_49165,N_49166,N_49167,N_49168,N_49169,N_49170,N_49171,N_49172,N_49173,N_49174,N_49175,N_49176,N_49177,N_49178,N_49179,N_49180,N_49181,N_49182,N_49183,N_49184,N_49185,N_49186,N_49187,N_49188,N_49189,N_49190,N_49191,N_49192,N_49193,N_49194,N_49195,N_49196,N_49197,N_49198,N_49199,N_49200,N_49201,N_49202,N_49203,N_49204,N_49205,N_49206,N_49207,N_49208,N_49209,N_49210,N_49211,N_49212,N_49213,N_49214,N_49215,N_49216,N_49217,N_49218,N_49219,N_49220,N_49221,N_49222,N_49223,N_49224,N_49225,N_49226,N_49227,N_49228,N_49229,N_49230,N_49231,N_49232,N_49233,N_49234,N_49235,N_49236,N_49237,N_49238,N_49239,N_49240,N_49241,N_49242,N_49243,N_49244,N_49245,N_49246,N_49247,N_49248,N_49249,N_49250,N_49251,N_49252,N_49253,N_49254,N_49255,N_49256,N_49257,N_49258,N_49259,N_49260,N_49261,N_49262,N_49263,N_49264,N_49265,N_49266,N_49267,N_49268,N_49269,N_49270,N_49271,N_49272,N_49273,N_49274,N_49275,N_49276,N_49277,N_49278,N_49279,N_49280,N_49281,N_49282,N_49283,N_49284,N_49285,N_49286,N_49287,N_49288,N_49289,N_49290,N_49291,N_49292,N_49293,N_49294,N_49295,N_49296,N_49297,N_49298,N_49299,N_49300,N_49301,N_49302,N_49303,N_49304,N_49305,N_49306,N_49307,N_49308,N_49309,N_49310,N_49311,N_49312,N_49313,N_49314,N_49315,N_49316,N_49317,N_49318,N_49319,N_49320,N_49321,N_49322,N_49323,N_49324,N_49325,N_49326,N_49327,N_49328,N_49329,N_49330,N_49331,N_49332,N_49333,N_49334,N_49335,N_49336,N_49337,N_49338,N_49339,N_49340,N_49341,N_49342,N_49343,N_49344,N_49345,N_49346,N_49347,N_49348,N_49349,N_49350,N_49351,N_49352,N_49353,N_49354,N_49355,N_49356,N_49357,N_49358,N_49359,N_49360,N_49361,N_49362,N_49363,N_49364,N_49365,N_49366,N_49367,N_49368,N_49369,N_49370,N_49371,N_49372,N_49373,N_49374,N_49375,N_49376,N_49377,N_49378,N_49379,N_49380,N_49381,N_49382,N_49383,N_49384,N_49385,N_49386,N_49387,N_49388,N_49389,N_49390,N_49391,N_49392,N_49393,N_49394,N_49395,N_49396,N_49397,N_49398,N_49399,N_49400,N_49401,N_49402,N_49403,N_49404,N_49405,N_49406,N_49407,N_49408,N_49409,N_49410,N_49411,N_49412,N_49413,N_49414,N_49415,N_49416,N_49417,N_49418,N_49419,N_49420,N_49421,N_49422,N_49423,N_49424,N_49425,N_49426,N_49427,N_49428,N_49429,N_49430,N_49431,N_49432,N_49433,N_49434,N_49435,N_49436,N_49437,N_49438,N_49439,N_49440,N_49441,N_49442,N_49443,N_49444,N_49445,N_49446,N_49447,N_49448,N_49449,N_49450,N_49451,N_49452,N_49453,N_49454,N_49455,N_49456,N_49457,N_49458,N_49459,N_49460,N_49461,N_49462,N_49463,N_49464,N_49465,N_49466,N_49467,N_49468,N_49469,N_49470,N_49471,N_49472,N_49473,N_49474,N_49475,N_49476,N_49477,N_49478,N_49479,N_49480,N_49481,N_49482,N_49483,N_49484,N_49485,N_49486,N_49487,N_49488,N_49489,N_49490,N_49491,N_49492,N_49493,N_49494,N_49495,N_49496,N_49497,N_49498,N_49499,N_49500,N_49501,N_49502,N_49503,N_49504,N_49505,N_49506,N_49507,N_49508,N_49509,N_49510,N_49511,N_49512,N_49513,N_49514,N_49515,N_49516,N_49517,N_49518,N_49519,N_49520,N_49521,N_49522,N_49523,N_49524,N_49525,N_49526,N_49527,N_49528,N_49529,N_49530,N_49531,N_49532,N_49533,N_49534,N_49535,N_49536,N_49537,N_49538,N_49539,N_49540,N_49541,N_49542,N_49543,N_49544,N_49545,N_49546,N_49547,N_49548,N_49549,N_49550,N_49551,N_49552,N_49553,N_49554,N_49555,N_49556,N_49557,N_49558,N_49559,N_49560,N_49561,N_49562,N_49563,N_49564,N_49565,N_49566,N_49567,N_49568,N_49569,N_49570,N_49571,N_49572,N_49573,N_49574,N_49575,N_49576,N_49577,N_49578,N_49579,N_49580,N_49581,N_49582,N_49583,N_49584,N_49585,N_49586,N_49587,N_49588,N_49589,N_49590,N_49591,N_49592,N_49593,N_49594,N_49595,N_49596,N_49597,N_49598,N_49599,N_49600,N_49601,N_49602,N_49603,N_49604,N_49605,N_49606,N_49607,N_49608,N_49609,N_49610,N_49611,N_49612,N_49613,N_49614,N_49615,N_49616,N_49617,N_49618,N_49619,N_49620,N_49621,N_49622,N_49623,N_49624,N_49625,N_49626,N_49627,N_49628,N_49629,N_49630,N_49631,N_49632,N_49633,N_49634,N_49635,N_49636,N_49637,N_49638,N_49639,N_49640,N_49641,N_49642,N_49643,N_49644,N_49645,N_49646,N_49647,N_49648,N_49649,N_49650,N_49651,N_49652,N_49653,N_49654,N_49655,N_49656,N_49657,N_49658,N_49659,N_49660,N_49661,N_49662,N_49663,N_49664,N_49665,N_49666,N_49667,N_49668,N_49669,N_49670,N_49671,N_49672,N_49673,N_49674,N_49675,N_49676,N_49677,N_49678,N_49679,N_49680,N_49681,N_49682,N_49683,N_49684,N_49685,N_49686,N_49687,N_49688,N_49689,N_49690,N_49691,N_49692,N_49693,N_49694,N_49695,N_49696,N_49697,N_49698,N_49699,N_49700,N_49701,N_49702,N_49703,N_49704,N_49705,N_49706,N_49707,N_49708,N_49709,N_49710,N_49711,N_49712,N_49713,N_49714,N_49715,N_49716,N_49717,N_49718,N_49719,N_49720,N_49721,N_49722,N_49723,N_49724,N_49725,N_49726,N_49727,N_49728,N_49729,N_49730,N_49731,N_49732,N_49733,N_49734,N_49735,N_49736,N_49737,N_49738,N_49739,N_49740,N_49741,N_49742,N_49743,N_49744,N_49745,N_49746,N_49747,N_49748,N_49749,N_49750,N_49751,N_49752,N_49753,N_49754,N_49755,N_49756,N_49757,N_49758,N_49759,N_49760,N_49761,N_49762,N_49763,N_49764,N_49765,N_49766,N_49767,N_49768,N_49769,N_49770,N_49771,N_49772,N_49773,N_49774,N_49775,N_49776,N_49777,N_49778,N_49779,N_49780,N_49781,N_49782,N_49783,N_49784,N_49785,N_49786,N_49787,N_49788,N_49789,N_49790,N_49791,N_49792,N_49793,N_49794,N_49795,N_49796,N_49797,N_49798,N_49799,N_49800,N_49801,N_49802,N_49803,N_49804,N_49805,N_49806,N_49807,N_49808,N_49809,N_49810,N_49811,N_49812,N_49813,N_49814,N_49815,N_49816,N_49817,N_49818,N_49819,N_49820,N_49821,N_49822,N_49823,N_49824,N_49825,N_49826,N_49827,N_49828,N_49829,N_49830,N_49831,N_49832,N_49833,N_49834,N_49835,N_49836,N_49837,N_49838,N_49839,N_49840,N_49841,N_49842,N_49843,N_49844,N_49845,N_49846,N_49847,N_49848,N_49849,N_49850,N_49851,N_49852,N_49853,N_49854,N_49855,N_49856,N_49857,N_49858,N_49859,N_49860,N_49861,N_49862,N_49863,N_49864,N_49865,N_49866,N_49867,N_49868,N_49869,N_49870,N_49871,N_49872,N_49873,N_49874,N_49875,N_49876,N_49877,N_49878,N_49879,N_49880,N_49881,N_49882,N_49883,N_49884,N_49885,N_49886,N_49887,N_49888,N_49889,N_49890,N_49891,N_49892,N_49893,N_49894,N_49895,N_49896,N_49897,N_49898,N_49899,N_49900,N_49901,N_49902,N_49903,N_49904,N_49905,N_49906,N_49907,N_49908,N_49909,N_49910,N_49911,N_49912,N_49913,N_49914,N_49915,N_49916,N_49917,N_49918,N_49919,N_49920,N_49921,N_49922,N_49923,N_49924,N_49925,N_49926,N_49927,N_49928,N_49929,N_49930,N_49931,N_49932,N_49933,N_49934,N_49935,N_49936,N_49937,N_49938,N_49939,N_49940,N_49941,N_49942,N_49943,N_49944,N_49945,N_49946,N_49947,N_49948,N_49949,N_49950,N_49951,N_49952,N_49953,N_49954,N_49955,N_49956,N_49957,N_49958,N_49959,N_49960,N_49961,N_49962,N_49963,N_49964,N_49965,N_49966,N_49967,N_49968,N_49969,N_49970,N_49971,N_49972,N_49973,N_49974,N_49975,N_49976,N_49977,N_49978,N_49979,N_49980,N_49981,N_49982,N_49983,N_49984,N_49985,N_49986,N_49987,N_49988,N_49989,N_49990,N_49991,N_49992,N_49993,N_49994,N_49995,N_49996,N_49997,N_49998,N_49999;
nand U0 (N_0,In_2206,In_4446);
xnor U1 (N_1,In_3642,In_3148);
nor U2 (N_2,In_1850,In_4717);
xor U3 (N_3,In_3923,In_4287);
nor U4 (N_4,In_2318,In_171);
nor U5 (N_5,In_4360,In_2483);
nand U6 (N_6,In_2857,In_2234);
and U7 (N_7,In_2145,In_1594);
or U8 (N_8,In_1158,In_2360);
nand U9 (N_9,In_3918,In_1958);
and U10 (N_10,In_3111,In_1191);
nand U11 (N_11,In_670,In_1146);
nand U12 (N_12,In_4310,In_3429);
nand U13 (N_13,In_663,In_1034);
and U14 (N_14,In_3000,In_4846);
nor U15 (N_15,In_70,In_458);
or U16 (N_16,In_2773,In_3309);
xor U17 (N_17,In_937,In_4740);
or U18 (N_18,In_2062,In_2501);
nand U19 (N_19,In_3407,In_1996);
and U20 (N_20,In_4133,In_3088);
or U21 (N_21,In_2278,In_2979);
nor U22 (N_22,In_3020,In_3871);
xor U23 (N_23,In_929,In_2306);
nand U24 (N_24,In_1095,In_688);
and U25 (N_25,In_1873,In_4732);
nor U26 (N_26,In_1061,In_2027);
nor U27 (N_27,In_2737,In_1316);
nor U28 (N_28,In_3784,In_4006);
nor U29 (N_29,In_133,In_1428);
and U30 (N_30,In_3463,In_1438);
and U31 (N_31,In_38,In_3953);
nor U32 (N_32,In_418,In_488);
nand U33 (N_33,In_3455,In_4612);
xnor U34 (N_34,In_3692,In_2976);
nand U35 (N_35,In_2601,In_1832);
or U36 (N_36,In_507,In_4866);
nand U37 (N_37,In_4134,In_4794);
nand U38 (N_38,In_4649,In_2210);
and U39 (N_39,In_2741,In_991);
nand U40 (N_40,In_1202,In_2943);
nor U41 (N_41,In_1214,In_4149);
xor U42 (N_42,In_4034,In_4731);
or U43 (N_43,In_2526,In_344);
and U44 (N_44,In_4874,In_260);
nor U45 (N_45,In_1371,In_255);
nand U46 (N_46,In_650,In_2980);
nor U47 (N_47,In_269,In_1354);
xor U48 (N_48,In_3457,In_1197);
nand U49 (N_49,In_1041,In_4154);
and U50 (N_50,In_642,In_4291);
and U51 (N_51,In_652,In_559);
nand U52 (N_52,In_747,In_4011);
or U53 (N_53,In_4334,In_1263);
or U54 (N_54,In_3855,In_4945);
nor U55 (N_55,In_662,In_1646);
xor U56 (N_56,In_74,In_4630);
xnor U57 (N_57,In_1939,In_184);
nor U58 (N_58,In_2950,In_1471);
nand U59 (N_59,In_2612,In_2585);
xnor U60 (N_60,In_1603,In_3936);
or U61 (N_61,In_1261,In_2772);
and U62 (N_62,In_4242,In_3329);
nand U63 (N_63,In_4458,In_1600);
nand U64 (N_64,In_4581,In_432);
and U65 (N_65,In_1487,In_811);
nand U66 (N_66,In_2494,In_53);
or U67 (N_67,In_3717,In_2322);
nor U68 (N_68,In_2411,In_2299);
nand U69 (N_69,In_1147,In_3114);
or U70 (N_70,In_3859,In_414);
nor U71 (N_71,In_3829,In_4986);
and U72 (N_72,In_2012,In_1784);
nor U73 (N_73,In_1301,In_2005);
nor U74 (N_74,In_2706,In_4471);
and U75 (N_75,In_1200,In_1307);
xnor U76 (N_76,In_590,In_3914);
nand U77 (N_77,In_157,In_4275);
or U78 (N_78,In_1442,In_1888);
and U79 (N_79,In_208,In_1419);
xnor U80 (N_80,In_2888,In_1489);
and U81 (N_81,In_1120,In_3048);
or U82 (N_82,In_1390,In_1836);
and U83 (N_83,In_2044,In_2783);
or U84 (N_84,In_3769,In_50);
xnor U85 (N_85,In_1479,In_1139);
and U86 (N_86,In_1008,In_1765);
and U87 (N_87,In_3804,In_2242);
nand U88 (N_88,In_3704,In_3690);
nor U89 (N_89,In_3683,In_4604);
or U90 (N_90,In_1098,In_4748);
and U91 (N_91,In_4441,In_3549);
and U92 (N_92,In_3198,In_4135);
or U93 (N_93,In_1551,In_4737);
or U94 (N_94,In_1967,In_1851);
nor U95 (N_95,In_837,In_323);
nor U96 (N_96,In_3567,In_2918);
or U97 (N_97,In_1258,In_2766);
nand U98 (N_98,In_1607,In_2368);
nor U99 (N_99,In_2220,In_3856);
nand U100 (N_100,In_2836,In_483);
xor U101 (N_101,In_3946,In_3343);
nor U102 (N_102,In_617,In_3112);
or U103 (N_103,In_4033,In_3365);
nand U104 (N_104,In_4433,In_4518);
xnor U105 (N_105,In_4286,In_1955);
nor U106 (N_106,In_3587,In_2059);
nor U107 (N_107,In_1229,In_3781);
nand U108 (N_108,In_164,In_4515);
nor U109 (N_109,In_2257,In_235);
and U110 (N_110,In_3864,In_4907);
and U111 (N_111,In_3865,In_637);
and U112 (N_112,In_3065,In_1367);
nor U113 (N_113,In_2952,In_3540);
xor U114 (N_114,In_4372,In_217);
nand U115 (N_115,In_1156,In_425);
xnor U116 (N_116,In_586,In_553);
or U117 (N_117,In_1020,In_2125);
xnor U118 (N_118,In_211,In_1647);
or U119 (N_119,In_3500,In_3612);
nor U120 (N_120,In_4123,In_4597);
xnor U121 (N_121,In_4009,In_2431);
and U122 (N_122,In_4750,In_3009);
and U123 (N_123,In_1122,In_2513);
or U124 (N_124,In_1302,In_3279);
and U125 (N_125,In_4652,In_897);
and U126 (N_126,In_3284,In_1802);
xnor U127 (N_127,In_1266,In_601);
xnor U128 (N_128,In_3830,In_1491);
and U129 (N_129,In_2058,In_2009);
nor U130 (N_130,In_1854,In_1525);
xor U131 (N_131,In_1773,In_979);
or U132 (N_132,In_2093,In_2759);
or U133 (N_133,In_4055,In_2003);
nand U134 (N_134,In_1231,In_3051);
nor U135 (N_135,In_1051,In_3396);
nand U136 (N_136,In_876,In_1159);
and U137 (N_137,In_2630,In_2860);
or U138 (N_138,In_1568,In_2427);
nand U139 (N_139,In_3815,In_915);
nand U140 (N_140,In_4582,In_1633);
or U141 (N_141,In_1726,In_819);
xnor U142 (N_142,In_1698,In_4200);
nand U143 (N_143,In_555,In_2111);
xnor U144 (N_144,In_1276,In_3214);
nand U145 (N_145,In_1183,In_1865);
or U146 (N_146,In_306,In_2907);
and U147 (N_147,In_2912,In_756);
or U148 (N_148,In_1547,In_4529);
nor U149 (N_149,In_3025,In_225);
or U150 (N_150,In_2792,In_4340);
and U151 (N_151,In_4807,In_1452);
xnor U152 (N_152,In_404,In_3403);
nand U153 (N_153,In_2345,In_4467);
xor U154 (N_154,In_4840,In_236);
and U155 (N_155,In_4451,In_2280);
nor U156 (N_156,In_1971,In_1256);
nand U157 (N_157,In_2964,In_3398);
nor U158 (N_158,In_4682,In_3057);
and U159 (N_159,In_630,In_316);
and U160 (N_160,In_1553,In_2130);
xnor U161 (N_161,In_441,In_4184);
xor U162 (N_162,In_2960,In_3139);
or U163 (N_163,In_2618,In_3966);
nor U164 (N_164,In_4815,In_4627);
and U165 (N_165,In_4653,In_4051);
and U166 (N_166,In_603,In_1816);
xor U167 (N_167,In_4657,In_4912);
and U168 (N_168,In_1524,In_277);
nor U169 (N_169,In_407,In_3318);
or U170 (N_170,In_4931,In_2372);
xor U171 (N_171,In_3597,In_176);
nor U172 (N_172,In_697,In_4877);
xor U173 (N_173,In_1017,In_1086);
or U174 (N_174,In_147,In_4332);
nand U175 (N_175,In_2935,In_227);
xnor U176 (N_176,In_291,In_4338);
xor U177 (N_177,In_93,In_1897);
or U178 (N_178,In_1255,In_2340);
or U179 (N_179,In_651,In_1578);
or U180 (N_180,In_2064,In_3723);
or U181 (N_181,In_3054,In_2507);
nor U182 (N_182,In_3615,In_885);
or U183 (N_183,In_421,In_3509);
and U184 (N_184,In_1507,In_2356);
xor U185 (N_185,In_2073,In_1523);
and U186 (N_186,In_268,In_1096);
and U187 (N_187,In_2538,In_354);
nand U188 (N_188,In_2853,In_1601);
nand U189 (N_189,In_1722,In_3640);
nor U190 (N_190,In_3473,In_3027);
nand U191 (N_191,In_3110,In_2877);
nand U192 (N_192,In_2108,In_1709);
nor U193 (N_193,In_992,In_4554);
nand U194 (N_194,In_3577,In_1628);
and U195 (N_195,In_2388,In_3145);
nand U196 (N_196,In_658,In_710);
nor U197 (N_197,In_1678,In_139);
nor U198 (N_198,In_1269,In_3444);
xnor U199 (N_199,In_2515,In_1430);
nand U200 (N_200,In_1552,In_3967);
xnor U201 (N_201,In_2365,In_1397);
xor U202 (N_202,In_1410,In_4754);
nor U203 (N_203,In_537,In_195);
nand U204 (N_204,In_3226,In_4647);
nor U205 (N_205,In_1683,In_455);
or U206 (N_206,In_2803,In_2495);
nor U207 (N_207,In_3311,In_365);
and U208 (N_208,In_3093,In_2545);
or U209 (N_209,In_3312,In_1192);
nor U210 (N_210,In_1282,In_3419);
xor U211 (N_211,In_2939,In_2705);
or U212 (N_212,In_411,In_2995);
or U213 (N_213,In_1198,In_4884);
and U214 (N_214,In_3087,In_4867);
xnor U215 (N_215,In_1223,In_3903);
nor U216 (N_216,In_813,In_3228);
nand U217 (N_217,In_2413,In_817);
nor U218 (N_218,In_2508,In_4054);
and U219 (N_219,In_3132,In_2861);
and U220 (N_220,In_620,In_3122);
and U221 (N_221,In_2711,In_2488);
or U222 (N_222,In_4041,In_1129);
nand U223 (N_223,In_2250,In_4428);
nand U224 (N_224,In_3432,In_4082);
nor U225 (N_225,In_47,In_3123);
or U226 (N_226,In_3080,In_341);
and U227 (N_227,In_242,In_3031);
nor U228 (N_228,In_3512,In_2347);
or U229 (N_229,In_1405,In_3584);
nand U230 (N_230,In_1974,In_1981);
or U231 (N_231,In_1799,In_2219);
nor U232 (N_232,In_2164,In_3861);
nand U233 (N_233,In_494,In_1277);
xor U234 (N_234,In_922,In_1614);
nor U235 (N_235,In_3131,In_3958);
and U236 (N_236,In_2118,In_2821);
xor U237 (N_237,In_1372,In_482);
xnor U238 (N_238,In_4537,In_4295);
nor U239 (N_239,In_606,In_3655);
nor U240 (N_240,In_2900,In_4519);
or U241 (N_241,In_1447,In_207);
nor U242 (N_242,In_281,In_3975);
xnor U243 (N_243,In_2933,In_4421);
or U244 (N_244,In_2983,In_4013);
nand U245 (N_245,In_1808,In_849);
nor U246 (N_246,In_4882,In_4853);
nand U247 (N_247,In_4959,In_3824);
nand U248 (N_248,In_2307,In_4021);
nand U249 (N_249,In_1220,In_3092);
nand U250 (N_250,In_1777,In_2049);
nand U251 (N_251,In_2668,In_4371);
or U252 (N_252,In_3108,In_2337);
and U253 (N_253,In_4778,In_2634);
xor U254 (N_254,In_704,In_2167);
nor U255 (N_255,In_2449,In_4313);
and U256 (N_256,In_4916,In_2566);
and U257 (N_257,In_493,In_874);
nand U258 (N_258,In_3186,In_3603);
nand U259 (N_259,In_2778,In_4160);
and U260 (N_260,In_3167,In_554);
nor U261 (N_261,In_1875,In_1323);
and U262 (N_262,In_2509,In_2977);
nor U263 (N_263,In_761,In_2894);
nor U264 (N_264,In_955,In_4536);
nand U265 (N_265,In_3870,In_4068);
nand U266 (N_266,In_1572,In_2863);
xnor U267 (N_267,In_615,In_135);
or U268 (N_268,In_1844,In_4486);
xnor U269 (N_269,In_4927,In_2727);
nand U270 (N_270,In_449,In_906);
or U271 (N_271,In_869,In_2987);
nand U272 (N_272,In_2826,In_2609);
nand U273 (N_273,In_327,In_1494);
or U274 (N_274,In_1920,In_2400);
and U275 (N_275,In_2619,In_2958);
xnor U276 (N_276,In_2382,In_179);
or U277 (N_277,In_3077,In_3336);
nor U278 (N_278,In_836,In_4150);
xnor U279 (N_279,In_917,In_290);
nor U280 (N_280,In_2945,In_2922);
or U281 (N_281,In_2066,In_2555);
and U282 (N_282,In_818,In_3443);
nor U283 (N_283,In_4684,In_1977);
and U284 (N_284,In_72,In_4022);
xnor U285 (N_285,In_2040,In_4863);
xor U286 (N_286,In_4662,In_2847);
or U287 (N_287,In_787,In_2442);
nor U288 (N_288,In_1260,In_4665);
and U289 (N_289,In_1758,In_1480);
and U290 (N_290,In_1846,In_4449);
and U291 (N_291,In_863,In_1610);
nand U292 (N_292,In_1927,In_2166);
xnor U293 (N_293,In_599,In_3873);
nand U294 (N_294,In_1993,In_4012);
xnor U295 (N_295,In_3394,In_3227);
or U296 (N_296,In_1420,In_3686);
or U297 (N_297,In_4583,In_1);
nor U298 (N_298,In_4819,In_959);
nand U299 (N_299,In_2386,In_4880);
and U300 (N_300,In_4786,In_1895);
or U301 (N_301,In_3204,In_3565);
and U302 (N_302,In_1132,In_4125);
nor U303 (N_303,In_873,In_1576);
and U304 (N_304,In_248,In_275);
xnor U305 (N_305,In_575,In_1626);
xor U306 (N_306,In_4557,In_487);
and U307 (N_307,In_1924,In_2190);
nor U308 (N_308,In_1217,In_2001);
and U309 (N_309,In_3192,In_1407);
nor U310 (N_310,In_4052,In_409);
or U311 (N_311,In_3633,In_4909);
and U312 (N_312,In_3260,In_3733);
xnor U313 (N_313,In_1885,In_760);
xor U314 (N_314,In_1327,In_3722);
nor U315 (N_315,In_3384,In_2461);
nand U316 (N_316,In_1393,In_3575);
and U317 (N_317,In_4553,In_2419);
xor U318 (N_318,In_947,In_4197);
xnor U319 (N_319,In_2045,In_1794);
xor U320 (N_320,In_739,In_3180);
xor U321 (N_321,In_990,In_2240);
nand U322 (N_322,In_717,In_2672);
xor U323 (N_323,In_4110,In_4997);
xor U324 (N_324,In_1554,In_1415);
and U325 (N_325,In_3168,In_2812);
xnor U326 (N_326,In_1731,In_3928);
xor U327 (N_327,In_726,In_4069);
nand U328 (N_328,In_2834,In_2344);
nor U329 (N_329,In_750,In_3357);
nand U330 (N_330,In_2680,In_4514);
xnor U331 (N_331,In_4812,In_3818);
xor U332 (N_332,In_4100,In_191);
nor U333 (N_333,In_3304,In_1374);
nor U334 (N_334,In_4131,In_2641);
xnor U335 (N_335,In_2645,In_4668);
nand U336 (N_336,In_2039,In_3295);
or U337 (N_337,In_2712,In_3202);
xnor U338 (N_338,In_1224,In_933);
xnor U339 (N_339,In_2774,In_4018);
and U340 (N_340,In_2915,In_1081);
and U341 (N_341,In_2055,In_2750);
nor U342 (N_342,In_4132,In_4233);
and U343 (N_343,In_1210,In_2937);
and U344 (N_344,In_1821,In_2971);
or U345 (N_345,In_4396,In_517);
or U346 (N_346,In_2004,In_3361);
xor U347 (N_347,In_1619,In_2006);
or U348 (N_348,In_764,In_3619);
nand U349 (N_349,In_2200,In_1026);
and U350 (N_350,In_2588,In_4602);
xnor U351 (N_351,In_4829,In_2867);
and U352 (N_352,In_4715,In_4593);
nand U353 (N_353,In_4698,In_1272);
nor U354 (N_354,In_4353,In_2137);
nor U355 (N_355,In_4228,In_4106);
xor U356 (N_356,In_4580,In_439);
xnor U357 (N_357,In_1687,In_4254);
or U358 (N_358,In_1597,In_1617);
nand U359 (N_359,In_2898,In_2684);
xnor U360 (N_360,In_3935,In_3024);
and U361 (N_361,In_1054,In_3511);
xnor U362 (N_362,In_3454,In_1715);
nor U363 (N_363,In_0,In_2238);
nor U364 (N_364,In_294,In_4071);
nand U365 (N_365,In_3833,In_1331);
and U366 (N_366,In_4605,In_2830);
nor U367 (N_367,In_311,In_3594);
or U368 (N_368,In_3089,In_745);
nand U369 (N_369,In_349,In_3327);
or U370 (N_370,In_2000,In_2729);
xor U371 (N_371,In_351,In_340);
xnor U372 (N_372,In_998,In_1696);
and U373 (N_373,In_2571,In_4445);
and U374 (N_374,In_1216,In_4845);
and U375 (N_375,In_461,In_1842);
nor U376 (N_376,In_4574,In_1182);
xnor U377 (N_377,In_2338,In_3947);
nand U378 (N_378,In_1475,In_4457);
xnor U379 (N_379,In_3694,In_4492);
and U380 (N_380,In_1596,In_373);
xnor U381 (N_381,In_4642,In_4891);
nand U382 (N_382,In_4911,In_206);
nand U383 (N_383,In_2472,In_3210);
or U384 (N_384,In_656,In_4356);
xor U385 (N_385,In_4152,In_2549);
xor U386 (N_386,In_4464,In_6);
or U387 (N_387,In_3240,In_4683);
xor U388 (N_388,In_4048,In_4671);
nor U389 (N_389,In_4424,In_3300);
nand U390 (N_390,In_1297,In_623);
nand U391 (N_391,In_1298,In_390);
xnor U392 (N_392,In_3090,In_1421);
nand U393 (N_393,In_1150,In_3413);
nor U394 (N_394,In_4820,In_3750);
nand U395 (N_395,In_941,In_1733);
xnor U396 (N_396,In_1819,In_1792);
nor U397 (N_397,In_989,In_1115);
xnor U398 (N_398,In_3430,In_3339);
nor U399 (N_399,In_1291,In_4147);
nand U400 (N_400,In_28,In_3047);
or U401 (N_401,In_1716,In_3360);
nand U402 (N_402,In_2463,In_4221);
and U403 (N_403,In_2196,In_2734);
nor U404 (N_404,In_2581,In_2870);
xnor U405 (N_405,In_3941,In_4024);
nand U406 (N_406,In_3620,In_1212);
and U407 (N_407,In_4250,In_3098);
xor U408 (N_408,In_2473,In_244);
xor U409 (N_409,In_2321,In_4251);
or U410 (N_410,In_4118,In_4249);
nor U411 (N_411,In_154,In_4643);
nand U412 (N_412,In_346,In_752);
nand U413 (N_413,In_3472,In_1933);
and U414 (N_414,In_1768,In_829);
and U415 (N_415,In_3171,In_2956);
nor U416 (N_416,In_4323,In_2379);
xor U417 (N_417,In_3673,In_2046);
nand U418 (N_418,In_2273,In_4259);
nand U419 (N_419,In_1416,In_1798);
nand U420 (N_420,In_584,In_1353);
and U421 (N_421,In_2702,In_4072);
and U422 (N_422,In_2673,In_2291);
xnor U423 (N_423,In_4383,In_2113);
xnor U424 (N_424,In_2840,In_2047);
or U425 (N_425,In_4103,In_2896);
xnor U426 (N_426,In_4699,In_2035);
and U427 (N_427,In_4512,In_3458);
and U428 (N_428,In_2380,In_2228);
nor U429 (N_429,In_1840,In_3126);
and U430 (N_430,In_3943,In_3726);
nand U431 (N_431,In_1395,In_249);
and U432 (N_432,In_2363,In_1848);
and U433 (N_433,In_4425,In_1668);
nor U434 (N_434,In_1339,In_705);
nor U435 (N_435,In_1860,In_1676);
or U436 (N_436,In_3654,In_4470);
and U437 (N_437,In_2532,In_3405);
or U438 (N_438,In_4212,In_51);
xor U439 (N_439,In_3544,In_3041);
nand U440 (N_440,In_4640,In_2224);
xnor U441 (N_441,In_2985,In_3516);
xnor U442 (N_442,In_1903,In_423);
and U443 (N_443,In_846,In_803);
nand U444 (N_444,In_2008,In_3113);
xor U445 (N_445,In_3306,In_4533);
or U446 (N_446,In_4994,In_4592);
nand U447 (N_447,In_3973,In_3996);
and U448 (N_448,In_1942,In_4155);
nand U449 (N_449,In_3397,In_3682);
and U450 (N_450,In_3857,In_1398);
xor U451 (N_451,In_2676,In_3888);
or U452 (N_452,In_151,In_796);
nand U453 (N_453,In_324,In_4830);
nor U454 (N_454,In_516,In_1930);
xnor U455 (N_455,In_3959,In_1082);
and U456 (N_456,In_4609,In_2133);
and U457 (N_457,In_4292,In_4113);
or U458 (N_458,In_800,In_1899);
or U459 (N_459,In_1664,In_1692);
and U460 (N_460,In_3158,In_3066);
or U461 (N_461,In_773,In_3847);
xor U462 (N_462,In_1677,In_1786);
nor U463 (N_463,In_1448,In_547);
nand U464 (N_464,In_1399,In_1097);
nand U465 (N_465,In_3207,In_3939);
or U466 (N_466,In_1278,In_823);
xor U467 (N_467,In_1176,In_2270);
and U468 (N_468,In_1136,In_3596);
nor U469 (N_469,In_742,In_4573);
nor U470 (N_470,In_4713,In_678);
nor U471 (N_471,In_3431,In_875);
nand U472 (N_472,In_610,In_4141);
or U473 (N_473,In_2042,In_375);
nor U474 (N_474,In_169,In_1028);
or U475 (N_475,In_196,In_2085);
or U476 (N_476,In_1834,In_489);
xnor U477 (N_477,In_76,In_138);
xnor U478 (N_478,In_2586,In_443);
and U479 (N_479,In_3745,In_1235);
or U480 (N_480,In_2409,In_2893);
nor U481 (N_481,In_1810,In_1591);
and U482 (N_482,In_2289,In_3749);
nand U483 (N_483,In_446,In_1824);
nand U484 (N_484,In_4809,In_3890);
nand U485 (N_485,In_4306,In_4925);
nor U486 (N_486,In_1239,In_15);
nor U487 (N_487,In_1247,In_2496);
and U488 (N_488,In_4238,In_531);
or U489 (N_489,In_473,In_4870);
nand U490 (N_490,In_2050,In_301);
or U491 (N_491,In_2267,In_2715);
xor U492 (N_492,In_2086,In_4146);
and U493 (N_493,In_769,In_2546);
nand U494 (N_494,In_2784,In_746);
xor U495 (N_495,In_4472,In_2747);
nand U496 (N_496,In_3561,In_3412);
xor U497 (N_497,In_2686,In_1121);
nand U498 (N_498,In_3743,In_3618);
nor U499 (N_499,In_768,In_320);
and U500 (N_500,In_1392,In_4172);
and U501 (N_501,N_46,In_4491);
nand U502 (N_502,In_2389,In_490);
and U503 (N_503,In_1157,In_4333);
or U504 (N_504,In_776,In_2357);
nand U505 (N_505,In_3359,In_2597);
or U506 (N_506,In_1329,In_4823);
nor U507 (N_507,N_100,In_556);
xnor U508 (N_508,In_1651,In_730);
xor U509 (N_509,In_629,In_4667);
nand U510 (N_510,In_3524,In_850);
nand U511 (N_511,In_4269,In_210);
xor U512 (N_512,In_2478,In_3545);
and U513 (N_513,In_3484,In_827);
nand U514 (N_514,In_4465,In_4431);
nor U515 (N_515,N_324,In_3799);
or U516 (N_516,In_2858,In_4168);
xor U517 (N_517,In_307,N_397);
and U518 (N_518,In_1826,In_3060);
xnor U519 (N_519,In_4596,In_2126);
or U520 (N_520,In_3528,In_3466);
nand U521 (N_521,In_999,N_112);
xnor U522 (N_522,In_880,In_4896);
and U523 (N_523,In_1883,In_2189);
or U524 (N_524,In_3572,In_2757);
or U525 (N_525,In_2829,In_2755);
xor U526 (N_526,In_644,In_2685);
xnor U527 (N_527,In_4436,In_595);
nand U528 (N_528,In_3156,In_382);
nor U529 (N_529,N_258,N_419);
or U530 (N_530,N_388,In_1859);
and U531 (N_531,In_2819,In_2623);
and U532 (N_532,In_2390,N_72);
or U533 (N_533,In_3628,In_2470);
nor U534 (N_534,In_3526,In_4375);
nand U535 (N_535,In_4215,In_3201);
nor U536 (N_536,In_2724,N_235);
nand U537 (N_537,N_311,N_134);
or U538 (N_538,In_3119,In_4349);
nor U539 (N_539,In_3518,In_2611);
and U540 (N_540,In_1847,In_3033);
xor U541 (N_541,In_3345,In_1673);
and U542 (N_542,In_1771,In_3677);
or U543 (N_543,In_3366,In_3464);
and U544 (N_544,In_2060,In_2453);
xor U545 (N_545,In_1749,In_4374);
nand U546 (N_546,In_3950,N_318);
nor U547 (N_547,In_4037,In_4852);
xnor U548 (N_548,In_2481,In_1338);
and U549 (N_549,In_121,In_2855);
nand U550 (N_550,In_358,In_1881);
or U551 (N_551,In_284,In_1712);
nor U552 (N_552,In_1403,In_3424);
nand U553 (N_553,In_3601,In_1118);
nor U554 (N_554,In_4361,N_273);
xor U555 (N_555,In_4237,N_474);
xnor U556 (N_556,In_4834,In_1040);
or U557 (N_557,In_2997,In_2521);
nand U558 (N_558,In_1242,N_67);
xnor U559 (N_559,In_4127,In_1584);
xor U560 (N_560,In_1569,In_218);
and U561 (N_561,In_1230,In_1478);
nand U562 (N_562,In_4305,In_743);
nand U563 (N_563,In_4173,In_3332);
or U564 (N_564,N_269,In_1005);
nor U565 (N_565,N_454,In_977);
nor U566 (N_566,In_3208,In_4634);
or U567 (N_567,In_95,In_3338);
xnor U568 (N_568,In_216,In_4452);
nor U569 (N_569,In_4569,In_4183);
and U570 (N_570,In_2231,In_1906);
nand U571 (N_571,In_1295,In_638);
xor U572 (N_572,In_611,In_660);
nand U573 (N_573,In_3016,In_3627);
xor U574 (N_574,In_986,In_312);
or U575 (N_575,In_701,In_1624);
xnor U576 (N_576,In_2010,In_4454);
or U577 (N_577,In_1439,In_1076);
nor U578 (N_578,In_2092,In_1679);
or U579 (N_579,In_1623,In_3288);
or U580 (N_580,In_3417,In_3991);
or U581 (N_581,In_1658,In_2805);
nor U582 (N_582,In_1805,In_3449);
xnor U583 (N_583,N_262,In_1706);
nor U584 (N_584,In_4507,N_74);
nand U585 (N_585,In_3255,In_1886);
xor U586 (N_586,N_38,N_481);
xor U587 (N_587,In_2341,In_4921);
xor U588 (N_588,N_449,In_2930);
nand U589 (N_589,N_244,In_2214);
and U590 (N_590,In_48,In_2667);
xor U591 (N_591,In_1953,In_4772);
xnor U592 (N_592,In_2769,In_1417);
xnor U593 (N_593,N_33,In_4900);
and U594 (N_594,In_1219,In_3287);
xnor U595 (N_595,N_445,N_93);
xnor U596 (N_596,In_799,In_3906);
xor U597 (N_597,In_566,In_2107);
or U598 (N_598,In_1383,In_145);
nand U599 (N_599,In_1112,In_408);
and U600 (N_600,In_4303,In_1822);
xor U601 (N_601,In_1917,In_1249);
or U602 (N_602,In_2296,In_2293);
and U603 (N_603,In_3889,In_1669);
and U604 (N_604,In_3795,In_3703);
and U605 (N_605,In_2403,In_2054);
nand U606 (N_606,In_3957,In_3532);
nor U607 (N_607,In_2799,In_1288);
nand U608 (N_608,In_713,In_385);
and U609 (N_609,In_627,In_526);
nor U610 (N_610,N_149,In_3043);
xnor U611 (N_611,In_3141,In_3154);
or U612 (N_612,In_3301,In_4014);
nor U613 (N_613,In_1342,In_3130);
or U614 (N_614,In_3945,In_864);
or U615 (N_615,In_1545,In_3868);
xnor U616 (N_616,In_4746,In_3489);
xor U617 (N_617,In_3370,In_3036);
and U618 (N_618,In_946,In_4535);
or U619 (N_619,In_1621,In_1501);
or U620 (N_620,In_1270,N_391);
and U621 (N_621,In_3334,In_58);
or U622 (N_622,In_2831,N_225);
xor U623 (N_623,In_3556,N_107);
nand U624 (N_624,In_1779,In_4130);
nor U625 (N_625,In_2816,In_3965);
xnor U626 (N_626,In_3028,In_2034);
nor U627 (N_627,In_4500,In_2777);
nor U628 (N_628,In_924,In_4965);
xor U629 (N_629,In_4969,In_2942);
xor U630 (N_630,In_4148,In_1688);
and U631 (N_631,In_731,In_4261);
nor U632 (N_632,In_4932,In_833);
and U633 (N_633,In_2543,In_4129);
nor U634 (N_634,In_4979,In_238);
or U635 (N_635,In_2193,N_349);
or U636 (N_636,N_166,In_2802);
nor U637 (N_637,In_4387,In_4047);
nand U638 (N_638,In_241,In_4347);
nand U639 (N_639,In_3460,In_1563);
nor U640 (N_640,In_1546,In_3143);
and U641 (N_641,In_485,In_4416);
or U642 (N_642,In_1063,In_4290);
or U643 (N_643,In_1376,In_347);
nand U644 (N_644,In_2638,N_286);
nand U645 (N_645,In_2175,In_4545);
xnor U646 (N_646,In_362,In_2304);
xnor U647 (N_647,In_699,In_3529);
and U648 (N_648,In_2259,In_4119);
or U649 (N_649,In_65,In_3003);
or U650 (N_650,In_4502,In_3035);
or U651 (N_651,In_3513,In_2701);
or U652 (N_652,In_1473,In_2725);
nand U653 (N_653,N_461,In_1032);
xor U654 (N_654,In_465,In_1818);
xnor U655 (N_655,In_1530,In_1740);
and U656 (N_656,In_545,In_370);
and U657 (N_657,In_4547,In_1556);
nand U658 (N_658,In_797,N_360);
xor U659 (N_659,In_278,In_3492);
xnor U660 (N_660,In_1893,In_549);
nand U661 (N_661,In_3705,In_198);
nor U662 (N_662,In_4708,In_1533);
nor U663 (N_663,In_1711,N_317);
and U664 (N_664,In_1887,In_3978);
or U665 (N_665,In_4996,In_3802);
and U666 (N_666,In_1037,N_69);
or U667 (N_667,In_4504,In_264);
nor U668 (N_668,In_4030,In_4940);
and U669 (N_669,In_4289,In_1155);
nand U670 (N_670,In_2332,In_3969);
nor U671 (N_671,In_4548,In_4962);
xnor U672 (N_672,In_4190,N_338);
nor U673 (N_673,In_3095,In_2535);
nand U674 (N_674,N_144,N_48);
and U675 (N_675,N_22,In_3034);
nand U676 (N_676,In_2462,In_1205);
xor U677 (N_677,In_2810,In_2838);
nor U678 (N_678,In_2517,In_724);
xnor U679 (N_679,In_22,In_3068);
or U680 (N_680,In_910,In_2726);
nor U681 (N_681,In_1046,In_180);
nor U682 (N_682,N_230,In_1666);
nor U683 (N_683,In_4344,N_190);
nand U684 (N_684,In_1222,In_616);
xnor U685 (N_685,In_3465,In_194);
and U686 (N_686,In_31,In_2536);
xnor U687 (N_687,In_529,In_2244);
nand U688 (N_688,In_2459,In_2872);
and U689 (N_689,In_2433,In_1055);
or U690 (N_690,In_129,In_2529);
xnor U691 (N_691,In_4894,In_1286);
and U692 (N_692,In_1434,In_3951);
and U693 (N_693,In_4097,In_3650);
nor U694 (N_694,In_4495,In_2974);
nor U695 (N_695,In_463,N_217);
nor U696 (N_696,N_373,In_2608);
or U697 (N_697,In_3563,N_276);
nand U698 (N_698,In_1170,In_1066);
nand U699 (N_699,In_4263,In_4493);
nand U700 (N_700,N_293,In_3013);
and U701 (N_701,In_142,In_2984);
nand U702 (N_702,In_2681,In_3931);
xnor U703 (N_703,In_3747,N_95);
nor U704 (N_704,N_196,In_3976);
and U705 (N_705,In_3600,In_4817);
xnor U706 (N_706,In_1234,In_4542);
xnor U707 (N_707,In_1163,In_3985);
and U708 (N_708,In_605,In_1188);
nor U709 (N_709,In_4769,N_362);
nand U710 (N_710,In_4074,In_150);
nor U711 (N_711,In_2664,In_4384);
or U712 (N_712,In_794,In_3919);
nor U713 (N_713,In_1583,In_3867);
or U714 (N_714,In_4297,In_4111);
or U715 (N_715,In_73,In_3152);
or U716 (N_716,In_4283,In_4838);
xnor U717 (N_717,In_363,In_3566);
nand U718 (N_718,In_994,In_433);
nand U719 (N_719,In_520,In_3026);
and U720 (N_720,In_3354,In_3586);
nor U721 (N_721,In_583,In_4217);
xor U722 (N_722,In_4762,In_3685);
nor U723 (N_723,In_1328,N_188);
nor U724 (N_724,In_305,In_1500);
nor U725 (N_725,In_4453,In_4423);
xnor U726 (N_726,In_3581,In_3712);
xnor U727 (N_727,In_4329,In_2312);
and U728 (N_728,In_4721,N_36);
nand U729 (N_729,In_124,N_4);
nor U730 (N_730,In_3663,In_3199);
xor U731 (N_731,In_2941,In_4905);
xor U732 (N_732,In_4831,In_3831);
or U733 (N_733,In_997,In_1761);
nor U734 (N_734,In_2541,In_4232);
and U735 (N_735,In_1631,In_2225);
xnor U736 (N_736,In_3753,In_3725);
xor U737 (N_737,In_2573,In_3948);
or U738 (N_738,In_203,In_1265);
or U739 (N_739,In_3254,N_426);
nor U740 (N_740,In_3713,In_4610);
nor U741 (N_741,In_4555,In_1208);
and U742 (N_742,In_2670,In_1634);
nor U743 (N_743,In_2839,In_1693);
xor U744 (N_744,In_4067,In_3508);
xor U745 (N_745,In_1078,In_4419);
nand U746 (N_746,In_2947,In_466);
nand U747 (N_747,In_2110,N_363);
and U748 (N_748,In_2222,N_227);
xnor U749 (N_749,N_249,In_1294);
nand U750 (N_750,In_1152,In_1817);
or U751 (N_751,In_3693,In_3569);
nor U752 (N_752,N_471,N_212);
nor U753 (N_753,In_1187,In_4801);
xor U754 (N_754,In_3876,In_1868);
xor U755 (N_755,In_2173,In_4955);
xor U756 (N_756,In_4968,In_4505);
xor U757 (N_757,In_1045,In_966);
nor U758 (N_758,In_2731,N_404);
xor U759 (N_759,In_1029,In_3729);
nor U760 (N_760,In_292,In_263);
xor U761 (N_761,N_270,In_1598);
and U762 (N_762,In_49,In_4177);
xnor U763 (N_763,In_4296,In_1505);
or U764 (N_764,N_18,In_1769);
xnor U765 (N_765,In_3698,In_4524);
nand U766 (N_766,In_3793,In_1253);
and U767 (N_767,N_468,In_3219);
nor U768 (N_768,In_1861,In_1548);
nor U769 (N_769,In_3900,In_4784);
xnor U770 (N_770,In_187,In_355);
nor U771 (N_771,In_2767,In_1511);
or U772 (N_772,In_3913,In_1093);
nor U773 (N_773,In_3271,In_2444);
xor U774 (N_774,In_4355,N_400);
xor U775 (N_775,In_3758,In_4083);
and U776 (N_776,In_1522,In_534);
and U777 (N_777,In_230,N_442);
xnor U778 (N_778,In_2075,In_808);
xor U779 (N_779,In_1788,In_4007);
nand U780 (N_780,In_1474,In_4753);
and U781 (N_781,In_4543,In_896);
and U782 (N_782,In_1935,In_2435);
xnor U783 (N_783,In_3149,In_1657);
nor U784 (N_784,In_4140,In_1517);
nand U785 (N_785,In_1827,N_403);
xor U786 (N_786,In_4725,In_3992);
nor U787 (N_787,In_4633,In_3368);
or U788 (N_788,In_3911,In_286);
xor U789 (N_789,In_2275,In_3651);
and U790 (N_790,In_708,In_4564);
nand U791 (N_791,In_3780,In_2656);
nor U792 (N_792,In_1510,In_2445);
nor U793 (N_793,In_1549,In_3428);
nand U794 (N_794,In_2825,In_1469);
nand U795 (N_795,In_3721,In_1320);
or U796 (N_796,In_2785,In_4923);
or U797 (N_797,In_1322,In_4015);
or U798 (N_798,In_4770,In_4941);
nor U799 (N_799,In_550,In_1825);
or U800 (N_800,In_396,In_4676);
and U801 (N_801,In_3296,N_302);
nand U802 (N_802,In_2690,In_3351);
or U803 (N_803,In_2642,In_4760);
xor U804 (N_804,In_1453,In_2161);
xnor U805 (N_805,In_3183,In_4622);
nor U806 (N_806,N_353,N_272);
or U807 (N_807,N_171,In_3647);
nor U808 (N_808,In_2547,In_3006);
or U809 (N_809,In_1684,In_3588);
nand U810 (N_810,In_1318,In_4330);
or U811 (N_811,In_18,In_2598);
nand U812 (N_812,N_265,In_672);
or U813 (N_813,In_4225,In_877);
xor U814 (N_814,In_1701,In_2868);
nand U815 (N_815,In_3944,In_3017);
or U816 (N_816,In_444,In_2334);
xnor U817 (N_817,In_237,N_389);
nor U818 (N_818,In_4503,In_4785);
and U819 (N_819,In_3987,In_329);
or U820 (N_820,In_3872,In_2636);
or U821 (N_821,In_934,In_464);
nor U822 (N_822,In_4243,In_4977);
xnor U823 (N_823,In_1739,In_591);
nand U824 (N_824,In_2120,In_457);
nor U825 (N_825,In_1084,In_1720);
xnor U826 (N_826,In_3744,In_14);
and U827 (N_827,In_4585,In_3427);
xor U828 (N_828,In_3225,N_469);
and U829 (N_829,In_852,In_2313);
nand U830 (N_830,In_4394,In_2071);
nand U831 (N_831,In_2248,N_147);
and U832 (N_832,In_1841,In_4181);
nand U833 (N_833,In_1815,In_4116);
xnor U834 (N_834,In_3246,In_4039);
or U835 (N_835,In_4187,In_4624);
or U836 (N_836,In_3882,In_4205);
xnor U837 (N_837,In_2089,In_231);
nand U838 (N_838,In_2697,In_2973);
nand U839 (N_839,In_4366,In_4641);
nand U840 (N_840,N_24,In_3536);
or U841 (N_841,In_3999,In_578);
or U842 (N_842,In_4170,In_4090);
or U843 (N_843,In_265,In_2644);
and U844 (N_844,In_2421,In_3420);
nor U845 (N_845,N_122,In_1332);
xor U846 (N_846,In_3467,In_4796);
or U847 (N_847,In_2707,N_495);
nand U848 (N_848,In_3238,In_4318);
xnor U849 (N_849,In_767,N_384);
and U850 (N_850,In_1542,In_4953);
nor U851 (N_851,In_551,In_3699);
xor U852 (N_852,In_4860,In_3515);
nand U853 (N_853,In_4903,In_4065);
nand U854 (N_854,In_2768,In_3589);
or U855 (N_855,In_2522,In_522);
and U856 (N_856,In_1512,In_502);
xor U857 (N_857,In_4917,In_1637);
or U858 (N_858,In_4218,In_1340);
nand U859 (N_859,In_4586,In_10);
nand U860 (N_860,N_145,In_4010);
nand U861 (N_861,In_3261,In_3280);
nor U862 (N_862,In_2245,N_352);
or U863 (N_863,In_4989,In_352);
or U864 (N_864,In_618,In_2070);
and U865 (N_865,In_4144,In_2735);
nand U866 (N_866,In_2438,In_851);
nand U867 (N_867,In_1360,In_3496);
xor U868 (N_868,In_749,N_115);
nand U869 (N_869,In_3008,In_3738);
and U870 (N_870,N_300,In_3748);
nor U871 (N_871,In_394,In_4397);
xor U872 (N_872,In_4326,In_4744);
xnor U873 (N_873,N_152,In_1655);
nor U874 (N_874,In_3325,In_1465);
and U875 (N_875,N_176,In_4966);
nand U876 (N_876,In_883,In_4673);
or U877 (N_877,In_3099,In_3814);
and U878 (N_878,In_77,In_82);
and U879 (N_879,In_830,In_3337);
nand U880 (N_880,In_2286,In_2391);
or U881 (N_881,In_3477,In_378);
nor U882 (N_882,N_448,In_921);
nand U883 (N_883,In_1285,In_2511);
nand U884 (N_884,In_1648,In_2370);
and U885 (N_885,In_1990,In_1386);
nor U886 (N_886,In_3754,In_2703);
and U887 (N_887,In_2780,In_3211);
nor U888 (N_888,In_4828,In_598);
nand U889 (N_889,In_2910,In_4724);
xor U890 (N_890,In_4992,In_943);
and U891 (N_891,In_4922,In_4983);
nand U892 (N_892,In_1661,In_1141);
xnor U893 (N_893,In_1632,In_92);
nand U894 (N_894,In_3574,In_3475);
nor U895 (N_895,In_1206,In_3984);
nand U896 (N_896,In_2119,N_260);
nor U897 (N_897,In_4407,In_3531);
nand U898 (N_898,In_2213,In_4985);
nor U899 (N_899,In_114,In_3399);
and U900 (N_900,In_1049,N_224);
or U901 (N_901,In_2663,In_832);
or U902 (N_902,N_344,In_3811);
or U903 (N_903,In_1388,In_4246);
xor U904 (N_904,N_44,N_2);
nand U905 (N_905,N_370,In_4764);
xnor U906 (N_906,In_1314,In_3789);
nor U907 (N_907,In_1864,In_969);
xor U908 (N_908,In_4273,N_98);
or U909 (N_909,N_140,In_1986);
nand U910 (N_910,In_3638,In_3487);
and U911 (N_911,In_1615,In_2800);
or U912 (N_912,In_2714,In_3562);
xor U913 (N_913,In_714,In_2704);
xor U914 (N_914,In_3030,In_3840);
and U915 (N_915,In_2843,In_1377);
nor U916 (N_916,In_1562,In_734);
or U917 (N_917,In_4053,In_3249);
xor U918 (N_918,In_4352,In_319);
and U919 (N_919,In_3495,N_51);
nor U920 (N_920,In_313,N_173);
nor U921 (N_921,In_1088,In_1418);
nor U922 (N_922,In_3004,In_1128);
xor U923 (N_923,In_2405,In_4060);
and U924 (N_924,In_256,In_3055);
or U925 (N_925,In_4063,In_4961);
nand U926 (N_926,N_256,In_3082);
xnor U927 (N_927,In_480,In_4489);
xnor U928 (N_928,N_472,In_4114);
nand U929 (N_929,In_2660,In_3897);
or U930 (N_930,In_3352,In_2294);
nor U931 (N_931,In_2355,In_4049);
or U932 (N_932,In_4162,In_1884);
xor U933 (N_933,In_2455,In_2415);
and U934 (N_934,In_2096,In_1236);
nand U935 (N_935,In_2474,In_1570);
and U936 (N_936,In_1605,In_140);
and U937 (N_937,In_2394,In_1267);
nor U938 (N_938,In_1889,In_3502);
nor U939 (N_939,In_3174,In_2978);
xor U940 (N_940,In_4936,In_552);
or U941 (N_941,In_2441,In_3373);
nor U942 (N_942,In_4697,In_2874);
or U943 (N_943,N_17,In_3303);
nand U944 (N_944,N_58,In_3348);
nor U945 (N_945,In_2765,In_3385);
xor U946 (N_946,In_589,In_4368);
nor U947 (N_947,In_2466,In_1918);
and U948 (N_948,In_3349,In_2019);
xor U949 (N_949,In_2954,In_4678);
xor U950 (N_950,In_612,In_3172);
nand U951 (N_951,In_4002,N_444);
xnor U952 (N_952,In_1459,In_952);
nor U953 (N_953,N_63,N_335);
or U954 (N_954,N_329,In_403);
or U955 (N_955,In_3474,In_646);
and U956 (N_956,In_1014,In_2723);
or U957 (N_957,In_2317,In_2677);
xnor U958 (N_958,In_2559,In_3740);
or U959 (N_959,In_4001,In_1496);
xnor U960 (N_960,In_2795,In_858);
xor U961 (N_961,N_39,In_2208);
or U962 (N_962,N_108,In_4319);
xor U963 (N_963,In_532,In_1988);
and U964 (N_964,In_3493,In_1516);
xnor U965 (N_965,In_4851,In_1718);
xnor U966 (N_966,In_1999,In_4498);
xor U967 (N_967,In_4913,In_86);
or U968 (N_968,In_3353,N_83);
xor U969 (N_969,In_26,N_455);
xor U970 (N_970,In_2621,N_0);
nand U971 (N_971,In_4781,In_4659);
and U972 (N_972,In_3267,In_930);
xnor U973 (N_973,In_4525,In_2077);
nor U974 (N_974,N_345,In_4193);
nand U975 (N_975,N_390,In_4398);
nor U976 (N_976,In_628,In_3825);
xor U977 (N_977,N_385,In_406);
nand U978 (N_978,In_2600,In_1109);
and U979 (N_979,In_1482,In_1738);
nor U980 (N_980,In_366,In_492);
or U981 (N_981,In_2106,In_2940);
xor U982 (N_982,In_2653,In_1675);
or U983 (N_983,In_1599,In_2187);
xnor U984 (N_984,In_1401,In_1774);
nor U985 (N_985,In_1912,In_1901);
and U986 (N_986,In_2216,In_951);
nand U987 (N_987,N_197,In_4156);
or U988 (N_988,In_2457,N_240);
nand U989 (N_989,In_4145,In_2505);
xor U990 (N_990,In_219,In_4689);
nand U991 (N_991,In_2763,N_143);
nor U992 (N_992,In_2142,In_4635);
nor U993 (N_993,In_755,In_4924);
or U994 (N_994,In_1303,In_3422);
xnor U995 (N_995,In_3711,In_1535);
nand U996 (N_996,In_4918,In_2846);
nand U997 (N_997,In_1364,In_4681);
nor U998 (N_998,N_132,In_753);
xnor U999 (N_999,N_223,In_3101);
and U1000 (N_1000,In_4755,In_1201);
or U1001 (N_1001,In_4229,In_356);
nor U1002 (N_1002,In_859,N_208);
xor U1003 (N_1003,In_3012,In_4484);
and U1004 (N_1004,In_450,In_1268);
and U1005 (N_1005,In_3848,In_2651);
nor U1006 (N_1006,In_926,N_733);
nor U1007 (N_1007,In_2625,In_2336);
nor U1008 (N_1008,N_975,In_4971);
nor U1009 (N_1009,In_1504,In_2258);
nand U1010 (N_1010,In_2364,In_2820);
and U1011 (N_1011,In_2396,In_1373);
nand U1012 (N_1012,In_4849,N_572);
xnor U1013 (N_1013,In_4915,In_436);
or U1014 (N_1014,In_2078,In_1160);
nand U1015 (N_1015,In_931,N_123);
and U1016 (N_1016,In_2639,In_2822);
and U1017 (N_1017,In_3218,In_3018);
nand U1018 (N_1018,In_1400,In_233);
and U1019 (N_1019,N_264,In_166);
and U1020 (N_1020,In_1567,In_4531);
or U1021 (N_1021,N_53,N_763);
xor U1022 (N_1022,In_2450,In_3741);
nand U1023 (N_1023,In_4862,In_1056);
nand U1024 (N_1024,N_927,In_1352);
or U1025 (N_1025,In_4095,In_98);
nand U1026 (N_1026,In_633,In_1379);
and U1027 (N_1027,N_999,In_434);
and U1028 (N_1028,In_252,In_119);
nor U1029 (N_1029,In_3269,In_1311);
or U1030 (N_1030,In_770,N_906);
or U1031 (N_1031,In_2565,In_1464);
and U1032 (N_1032,In_1685,In_3137);
or U1033 (N_1033,N_587,In_4253);
nand U1034 (N_1034,In_4220,In_1426);
nand U1035 (N_1035,In_2352,In_308);
nand U1036 (N_1036,In_2856,N_738);
nand U1037 (N_1037,In_3525,In_3039);
and U1038 (N_1038,In_3448,In_3081);
nand U1039 (N_1039,In_1934,In_2832);
or U1040 (N_1040,In_1994,In_4782);
and U1041 (N_1041,N_50,In_3850);
xor U1042 (N_1042,In_1870,In_2742);
nand U1043 (N_1043,In_1645,In_4739);
and U1044 (N_1044,In_42,In_4795);
or U1045 (N_1045,In_3878,In_888);
xor U1046 (N_1046,In_1780,N_887);
xor U1047 (N_1047,N_770,In_3406);
or U1048 (N_1048,In_872,N_599);
xor U1049 (N_1049,In_3237,In_3342);
or U1050 (N_1050,In_105,In_2132);
xor U1051 (N_1051,In_4705,In_4165);
or U1052 (N_1052,In_1089,In_3494);
nor U1053 (N_1053,N_483,In_3049);
nand U1054 (N_1054,In_2349,In_1488);
and U1055 (N_1055,In_4901,In_2782);
and U1056 (N_1056,In_1173,N_592);
nand U1057 (N_1057,In_90,In_1345);
or U1058 (N_1058,In_1245,In_1103);
nand U1059 (N_1059,In_3389,In_3164);
and U1060 (N_1060,In_2290,In_326);
and U1061 (N_1061,In_985,In_4223);
xnor U1062 (N_1062,N_159,In_2276);
xor U1063 (N_1063,In_3229,In_3050);
nor U1064 (N_1064,N_901,N_429);
and U1065 (N_1065,In_1010,In_4272);
or U1066 (N_1066,N_82,In_1812);
nand U1067 (N_1067,In_4879,In_4696);
nor U1068 (N_1068,In_2593,In_2996);
and U1069 (N_1069,In_866,In_2594);
xor U1070 (N_1070,In_2962,In_4245);
nand U1071 (N_1071,In_2342,In_1306);
nor U1072 (N_1072,In_727,In_683);
xnor U1073 (N_1073,In_845,N_456);
or U1074 (N_1074,In_4710,In_904);
and U1075 (N_1075,In_3297,N_307);
and U1076 (N_1076,In_4209,In_4672);
or U1077 (N_1077,In_2076,N_245);
and U1078 (N_1078,N_868,In_1347);
and U1079 (N_1079,In_1110,In_523);
and U1080 (N_1080,In_691,In_37);
nor U1081 (N_1081,In_1030,In_2695);
nand U1082 (N_1082,In_1957,In_4422);
and U1083 (N_1083,N_976,In_1804);
xnor U1084 (N_1084,In_1050,In_3021);
xnor U1085 (N_1085,In_2968,In_3922);
nor U1086 (N_1086,In_3203,In_1938);
nor U1087 (N_1087,In_1035,In_3274);
xnor U1088 (N_1088,In_4089,N_40);
nor U1089 (N_1089,In_2011,In_3185);
nand U1090 (N_1090,In_4307,N_586);
and U1091 (N_1091,In_1140,In_2574);
nor U1092 (N_1092,In_1620,N_303);
xor U1093 (N_1093,N_674,In_4546);
nand U1094 (N_1094,In_804,In_1370);
and U1095 (N_1095,In_3307,In_2764);
and U1096 (N_1096,In_213,N_170);
and U1097 (N_1097,N_951,N_1);
xnor U1098 (N_1098,N_747,In_735);
and U1099 (N_1099,N_325,N_984);
or U1100 (N_1100,N_517,In_4481);
xor U1101 (N_1101,In_1734,N_237);
nand U1102 (N_1102,In_2051,In_4316);
nand U1103 (N_1103,In_160,In_2146);
and U1104 (N_1104,In_667,In_1514);
xnor U1105 (N_1105,N_973,N_343);
nand U1106 (N_1106,In_1196,In_2330);
and U1107 (N_1107,N_96,N_155);
xor U1108 (N_1108,N_486,In_1166);
and U1109 (N_1109,In_4718,N_814);
nor U1110 (N_1110,In_4391,In_2875);
nand U1111 (N_1111,N_940,N_626);
xor U1112 (N_1112,N_470,In_780);
nand U1113 (N_1113,In_2432,N_116);
nand U1114 (N_1114,N_891,In_3425);
nor U1115 (N_1115,N_160,In_3893);
nand U1116 (N_1116,In_2889,N_588);
nor U1117 (N_1117,In_4380,In_2647);
or U1118 (N_1118,In_4878,In_2253);
xnor U1119 (N_1119,In_1012,In_405);
or U1120 (N_1120,In_3904,N_179);
nand U1121 (N_1121,In_4709,In_2969);
xnor U1122 (N_1122,In_3634,In_2953);
nand U1123 (N_1123,In_920,In_3952);
nand U1124 (N_1124,N_997,In_1843);
nor U1125 (N_1125,In_1335,In_2603);
xor U1126 (N_1126,In_2627,N_742);
xor U1127 (N_1127,In_3541,In_197);
nor U1128 (N_1128,In_1589,In_3925);
or U1129 (N_1129,In_322,In_254);
nor U1130 (N_1130,In_212,In_1114);
xor U1131 (N_1131,N_547,In_2662);
and U1132 (N_1132,In_2243,In_2849);
or U1133 (N_1133,In_3480,In_143);
or U1134 (N_1134,In_2972,In_4248);
or U1135 (N_1135,In_2249,N_769);
nand U1136 (N_1136,N_417,In_1165);
or U1137 (N_1137,N_501,In_1437);
nor U1138 (N_1138,In_1604,In_512);
nand U1139 (N_1139,In_1275,N_500);
nor U1140 (N_1140,In_3233,In_2654);
or U1141 (N_1141,N_573,In_81);
or U1142 (N_1142,In_215,In_2553);
xnor U1143 (N_1143,In_3653,N_818);
and U1144 (N_1144,In_521,In_2626);
nor U1145 (N_1145,N_735,In_2602);
and U1146 (N_1146,In_1048,In_2624);
nor U1147 (N_1147,In_4179,In_1389);
or U1148 (N_1148,In_4325,In_1300);
nor U1149 (N_1149,N_760,In_4902);
and U1150 (N_1150,In_2414,In_1343);
and U1151 (N_1151,In_1867,N_575);
xor U1152 (N_1152,N_219,N_142);
nor U1153 (N_1153,In_3933,In_901);
nor U1154 (N_1154,In_3503,N_582);
and U1155 (N_1155,In_1811,In_2739);
nor U1156 (N_1156,In_3375,N_675);
or U1157 (N_1157,In_4459,In_2961);
xor U1158 (N_1158,In_1039,In_706);
xnor U1159 (N_1159,In_3102,In_369);
nand U1160 (N_1160,In_4405,In_940);
or U1161 (N_1161,In_3220,In_1564);
or U1162 (N_1162,In_2315,In_170);
or U1163 (N_1163,In_4666,N_866);
nor U1164 (N_1164,In_223,In_2970);
or U1165 (N_1165,In_2580,N_630);
and U1166 (N_1166,In_295,In_1060);
nor U1167 (N_1167,In_4651,In_604);
nor U1168 (N_1168,In_177,In_2679);
or U1169 (N_1169,N_889,In_2994);
and U1170 (N_1170,N_700,In_524);
or U1171 (N_1171,In_4331,N_539);
and U1172 (N_1172,In_2850,N_741);
nor U1173 (N_1173,In_1915,In_1697);
xor U1174 (N_1174,N_114,In_4342);
and U1175 (N_1175,In_120,In_3837);
or U1176 (N_1176,In_2484,In_4277);
or U1177 (N_1177,In_1111,In_4378);
nand U1178 (N_1178,N_734,N_55);
xnor U1179 (N_1179,In_2254,In_200);
xnor U1180 (N_1180,In_2957,N_974);
xnor U1181 (N_1181,In_427,In_2416);
xor U1182 (N_1182,In_3905,N_649);
nand U1183 (N_1183,In_1581,N_576);
xnor U1184 (N_1184,In_3990,In_2615);
nor U1185 (N_1185,In_448,In_4399);
xor U1186 (N_1186,In_3507,In_4700);
xor U1187 (N_1187,N_151,In_2115);
and U1188 (N_1188,In_417,In_4008);
or U1189 (N_1189,N_433,In_2353);
xor U1190 (N_1190,N_832,N_202);
xor U1191 (N_1191,In_3330,In_892);
nand U1192 (N_1192,N_989,In_4285);
xor U1193 (N_1193,In_1254,In_4881);
nor U1194 (N_1194,N_136,In_1172);
nand U1195 (N_1195,In_2437,In_3823);
xor U1196 (N_1196,N_291,In_4534);
nor U1197 (N_1197,In_825,N_650);
or U1198 (N_1198,In_3648,In_1194);
and U1199 (N_1199,In_2103,In_2669);
xnor U1200 (N_1200,In_3418,In_4523);
or U1201 (N_1201,In_4898,In_4268);
xor U1202 (N_1202,In_1641,In_3989);
nor U1203 (N_1203,N_858,In_4958);
nand U1204 (N_1204,In_3129,N_137);
xnor U1205 (N_1205,In_2762,In_4702);
xnor U1206 (N_1206,In_2744,In_3205);
nand U1207 (N_1207,In_1296,In_3550);
nand U1208 (N_1208,In_3762,In_4541);
nand U1209 (N_1209,In_2447,In_2884);
nor U1210 (N_1210,N_460,In_1913);
nand U1211 (N_1211,In_4045,N_175);
and U1212 (N_1212,N_169,In_855);
or U1213 (N_1213,In_3986,In_1909);
nor U1214 (N_1214,N_666,In_1998);
nand U1215 (N_1215,In_422,In_1727);
xnor U1216 (N_1216,In_1271,In_3560);
nand U1217 (N_1217,N_347,In_3212);
nand U1218 (N_1218,In_2,In_2564);
nor U1219 (N_1219,In_3666,N_736);
nor U1220 (N_1220,In_2719,In_2885);
xor U1221 (N_1221,In_172,N_790);
and U1222 (N_1222,In_4645,In_3052);
or U1223 (N_1223,In_3636,In_4964);
xnor U1224 (N_1224,In_1751,In_3875);
and U1225 (N_1225,In_1719,In_2828);
xor U1226 (N_1226,In_2114,In_626);
xor U1227 (N_1227,In_67,In_3401);
nor U1228 (N_1228,In_2256,N_242);
or U1229 (N_1229,In_1928,In_3727);
xor U1230 (N_1230,N_7,N_65);
nor U1231 (N_1231,In_4972,In_798);
and U1232 (N_1232,In_460,In_2124);
nor U1233 (N_1233,In_106,In_389);
or U1234 (N_1234,In_958,In_1280);
or U1235 (N_1235,N_439,In_887);
or U1236 (N_1236,In_865,In_3841);
nor U1237 (N_1237,In_107,N_795);
or U1238 (N_1238,In_1476,N_523);
nand U1239 (N_1239,N_157,In_2016);
nand U1240 (N_1240,In_2141,N_552);
nand U1241 (N_1241,In_274,In_3235);
or U1242 (N_1242,In_826,N_604);
nand U1243 (N_1243,In_546,In_3294);
nand U1244 (N_1244,In_4230,In_3323);
xor U1245 (N_1245,In_536,N_101);
or U1246 (N_1246,N_606,In_3390);
xnor U1247 (N_1247,In_4571,N_691);
and U1248 (N_1248,In_3146,N_758);
nand U1249 (N_1249,N_9,In_508);
or U1250 (N_1250,In_4720,In_1361);
nor U1251 (N_1251,N_715,In_4204);
or U1252 (N_1252,In_3346,In_687);
nor U1253 (N_1253,N_844,In_2746);
xor U1254 (N_1254,N_530,In_173);
nor U1255 (N_1255,In_881,In_3979);
nand U1256 (N_1256,In_964,In_1717);
and U1257 (N_1257,N_898,In_3971);
and U1258 (N_1258,In_4701,N_764);
and U1259 (N_1259,N_948,In_2468);
xnor U1260 (N_1260,In_1425,N_996);
and U1261 (N_1261,In_4670,In_805);
nand U1262 (N_1262,In_2139,In_1644);
and U1263 (N_1263,In_4496,N_550);
or U1264 (N_1264,In_1073,In_1609);
or U1265 (N_1265,In_3144,In_2905);
nand U1266 (N_1266,In_4889,In_3236);
nand U1267 (N_1267,In_1879,N_861);
nor U1268 (N_1268,In_1033,N_210);
nor U1269 (N_1269,In_2177,In_4362);
or U1270 (N_1270,N_644,N_31);
xnor U1271 (N_1271,N_900,In_2392);
or U1272 (N_1272,In_4339,In_148);
and U1273 (N_1273,In_1778,In_2297);
or U1274 (N_1274,In_1925,In_1264);
xnor U1275 (N_1275,N_903,In_4429);
or U1276 (N_1276,N_49,In_4084);
nand U1277 (N_1277,N_396,In_1659);
xnor U1278 (N_1278,In_186,In_3716);
or U1279 (N_1279,In_2512,In_3103);
nand U1280 (N_1280,In_3708,In_4777);
nor U1281 (N_1281,In_296,In_4026);
or U1282 (N_1282,In_1813,In_3812);
and U1283 (N_1283,In_1094,N_634);
xnor U1284 (N_1284,N_379,N_865);
xnor U1285 (N_1285,In_3213,In_1950);
and U1286 (N_1286,In_91,N_757);
nand U1287 (N_1287,In_2425,In_55);
nand U1288 (N_1288,In_3954,In_185);
nand U1289 (N_1289,In_2144,In_4175);
and U1290 (N_1290,In_4417,N_938);
xnor U1291 (N_1291,N_277,In_1506);
nor U1292 (N_1292,In_4843,In_29);
and U1293 (N_1293,In_3506,In_4163);
xnor U1294 (N_1294,In_3641,In_4094);
and U1295 (N_1295,N_520,In_2482);
xnor U1296 (N_1296,In_4793,In_2351);
xor U1297 (N_1297,N_684,In_3446);
nor U1298 (N_1298,In_1062,In_2485);
or U1299 (N_1299,In_2186,In_3604);
nand U1300 (N_1300,In_3283,N_499);
nand U1301 (N_1301,In_3488,In_199);
nand U1302 (N_1302,In_3378,In_3340);
nand U1303 (N_1303,In_2866,In_1767);
nand U1304 (N_1304,In_1814,N_703);
nand U1305 (N_1305,In_4939,In_2026);
nor U1306 (N_1306,In_3902,In_835);
xnor U1307 (N_1307,In_671,In_2383);
xnor U1308 (N_1308,In_518,N_506);
nor U1309 (N_1309,In_3476,In_2657);
xnor U1310 (N_1310,N_886,N_829);
xor U1311 (N_1311,N_233,In_45);
xor U1312 (N_1312,In_856,In_4260);
or U1313 (N_1313,In_4365,In_505);
and U1314 (N_1314,In_4637,In_1869);
nor U1315 (N_1315,N_936,N_518);
and U1316 (N_1316,N_986,In_822);
nor U1317 (N_1317,In_1571,In_3230);
nand U1318 (N_1318,In_4549,In_3746);
or U1319 (N_1319,N_924,In_3423);
or U1320 (N_1320,N_354,N_730);
and U1321 (N_1321,In_3834,N_62);
and U1322 (N_1322,In_4078,In_167);
or U1323 (N_1323,In_175,In_3632);
nand U1324 (N_1324,In_4745,In_1672);
nand U1325 (N_1325,In_3456,In_1613);
nor U1326 (N_1326,In_118,In_20);
nor U1327 (N_1327,In_4798,N_556);
and U1328 (N_1328,In_3022,N_118);
nand U1329 (N_1329,In_1877,In_3846);
or U1330 (N_1330,In_1211,In_3216);
nand U1331 (N_1331,In_66,In_3469);
and U1332 (N_1332,In_4899,In_3960);
nand U1333 (N_1333,In_3790,In_653);
nor U1334 (N_1334,In_3613,In_938);
xnor U1335 (N_1335,N_238,N_200);
xnor U1336 (N_1336,In_2153,N_513);
or U1337 (N_1337,In_944,In_4926);
or U1338 (N_1338,N_358,In_3827);
nand U1339 (N_1339,In_2959,In_2184);
nor U1340 (N_1340,In_562,In_1989);
nor U1341 (N_1341,N_441,In_2990);
xor U1342 (N_1342,In_3165,N_670);
xor U1343 (N_1343,In_3116,In_3061);
xnor U1344 (N_1344,In_364,In_1135);
nor U1345 (N_1345,N_488,In_3912);
and U1346 (N_1346,N_813,N_902);
and U1347 (N_1347,In_2815,In_3313);
or U1348 (N_1348,N_564,In_3910);
nand U1349 (N_1349,In_331,In_23);
and U1350 (N_1350,In_3701,N_218);
and U1351 (N_1351,N_121,In_3435);
nor U1352 (N_1352,In_2903,In_3363);
xor U1353 (N_1353,In_2923,In_3191);
and U1354 (N_1354,In_533,In_2020);
xor U1355 (N_1355,In_1611,In_1625);
nand U1356 (N_1356,In_1274,In_1443);
xor U1357 (N_1357,In_987,In_3367);
nor U1358 (N_1358,N_125,N_553);
or U1359 (N_1359,N_708,In_4773);
nor U1360 (N_1360,In_1574,In_1590);
xnor U1361 (N_1361,N_150,In_3854);
nor U1362 (N_1362,In_4842,In_3672);
or U1363 (N_1363,In_871,In_4343);
xnor U1364 (N_1364,N_321,In_608);
and U1365 (N_1365,In_1167,In_1031);
nor U1366 (N_1366,In_1783,In_2587);
and U1367 (N_1367,In_2199,In_1852);
nand U1368 (N_1368,In_3724,In_3688);
nand U1369 (N_1369,In_3079,In_4943);
xnor U1370 (N_1370,In_4595,N_612);
nand U1371 (N_1371,In_4791,In_4722);
xnor U1372 (N_1372,In_467,In_1126);
or U1373 (N_1373,In_3842,In_2456);
xor U1374 (N_1374,In_2084,N_12);
and U1375 (N_1375,In_1987,In_2057);
nand U1376 (N_1376,In_2015,In_1789);
or U1377 (N_1377,In_1273,N_645);
and U1378 (N_1378,In_2013,N_357);
or U1379 (N_1379,In_4774,In_2048);
xnor U1380 (N_1380,In_4461,In_894);
or U1381 (N_1381,In_234,In_4482);
nand U1382 (N_1382,In_12,In_1575);
xnor U1383 (N_1383,In_1287,N_752);
and U1384 (N_1384,In_1127,N_802);
or U1385 (N_1385,In_4763,In_3625);
xnor U1386 (N_1386,In_3898,N_937);
nor U1387 (N_1387,In_2924,In_348);
and U1388 (N_1388,In_779,In_1785);
nand U1389 (N_1389,In_4077,In_4897);
nor U1390 (N_1390,In_619,In_2104);
or U1391 (N_1391,In_1947,In_936);
nor U1392 (N_1392,N_751,In_4138);
xor U1393 (N_1393,In_3256,N_540);
and U1394 (N_1394,In_2659,In_4675);
and U1395 (N_1395,In_46,In_3921);
xor U1396 (N_1396,In_4761,In_1193);
and U1397 (N_1397,N_731,In_3819);
and U1398 (N_1398,In_2476,In_1334);
or U1399 (N_1399,In_4735,In_914);
xor U1400 (N_1400,In_1946,In_2925);
and U1401 (N_1401,In_2233,In_342);
nor U1402 (N_1402,In_2033,In_3932);
xnor U1403 (N_1403,In_1209,In_4513);
xor U1404 (N_1404,In_3874,In_479);
and U1405 (N_1405,N_480,In_659);
or U1406 (N_1406,In_128,In_1123);
xor U1407 (N_1407,N_549,In_2149);
and U1408 (N_1408,In_2572,In_675);
and U1409 (N_1409,In_183,N_744);
and U1410 (N_1410,In_844,In_1940);
nand U1411 (N_1411,In_4468,In_398);
xor U1412 (N_1412,In_353,In_569);
nand U1413 (N_1413,In_821,N_640);
xor U1414 (N_1414,In_4759,In_1384);
nor U1415 (N_1415,In_1959,In_2281);
or U1416 (N_1416,N_451,In_649);
nand U1417 (N_1417,In_87,In_3756);
nor U1418 (N_1418,In_2728,In_2756);
xor U1419 (N_1419,In_4320,In_1363);
nand U1420 (N_1420,N_935,In_4835);
and U1421 (N_1421,In_3438,In_751);
and U1422 (N_1422,In_3644,In_3072);
nand U1423 (N_1423,In_2174,In_4598);
nor U1424 (N_1424,In_371,In_4201);
nand U1425 (N_1425,N_103,N_771);
xnor U1426 (N_1426,N_987,In_32);
or U1427 (N_1427,N_524,In_3687);
xnor U1428 (N_1428,N_611,In_1142);
nor U1429 (N_1429,N_412,N_828);
nand U1430 (N_1430,In_945,In_4389);
or U1431 (N_1431,In_2643,In_108);
and U1432 (N_1432,In_2592,In_572);
and U1433 (N_1433,In_3335,In_737);
nor U1434 (N_1434,In_1932,In_4216);
or U1435 (N_1435,In_841,N_653);
and U1436 (N_1436,In_1820,In_3785);
nor U1437 (N_1437,N_206,In_3980);
nor U1438 (N_1438,N_655,N_187);
nor U1439 (N_1439,In_3646,In_3775);
nand U1440 (N_1440,N_346,In_2558);
nand U1441 (N_1441,N_287,In_462);
nor U1442 (N_1442,In_3534,In_1493);
or U1443 (N_1443,N_128,In_468);
and U1444 (N_1444,In_4516,In_2302);
xnor U1445 (N_1445,N_879,In_4488);
and U1446 (N_1446,N_877,In_309);
xnor U1447 (N_1447,In_3533,In_4151);
nand U1448 (N_1448,In_1406,In_2191);
and U1449 (N_1449,In_4247,In_3362);
nor U1450 (N_1450,In_2053,In_579);
xor U1451 (N_1451,In_3270,In_2617);
xor U1452 (N_1452,In_1629,In_4208);
nand U1453 (N_1453,N_310,In_376);
or U1454 (N_1454,In_1466,In_563);
xor U1455 (N_1455,In_3656,In_1460);
xor U1456 (N_1456,In_4414,In_4040);
or U1457 (N_1457,In_2018,In_1538);
nor U1458 (N_1458,N_339,In_2030);
or U1459 (N_1459,In_3252,In_4613);
or U1460 (N_1460,In_4115,In_205);
or U1461 (N_1461,In_2326,In_2237);
or U1462 (N_1462,In_3277,In_967);
and U1463 (N_1463,In_4,In_878);
nor U1464 (N_1464,In_4528,In_3771);
nor U1465 (N_1465,In_962,In_807);
xnor U1466 (N_1466,In_415,N_654);
xnor U1467 (N_1467,In_3161,In_4563);
nor U1468 (N_1468,N_192,In_1508);
nand U1469 (N_1469,N_94,N_850);
nor U1470 (N_1470,In_4847,In_1527);
or U1471 (N_1471,In_4444,In_4615);
xnor U1472 (N_1472,In_4057,N_398);
or U1473 (N_1473,In_318,In_3883);
or U1474 (N_1474,In_2616,In_4410);
xor U1475 (N_1475,In_942,In_4854);
or U1476 (N_1476,In_4227,N_11);
or U1477 (N_1477,In_136,In_3331);
xor U1478 (N_1478,In_3442,N_526);
xor U1479 (N_1479,N_477,In_2477);
or U1480 (N_1480,N_904,In_648);
xnor U1481 (N_1481,In_2448,In_1184);
nor U1482 (N_1482,N_41,N_165);
or U1483 (N_1483,In_2790,In_2099);
nand U1484 (N_1484,In_4679,In_360);
xnor U1485 (N_1485,In_4706,N_80);
xor U1486 (N_1486,In_3019,In_3962);
xor U1487 (N_1487,N_706,In_2993);
or U1488 (N_1488,In_332,In_3657);
nor U1489 (N_1489,In_4346,In_445);
xnor U1490 (N_1490,N_234,In_729);
xnor U1491 (N_1491,In_775,In_2770);
nand U1492 (N_1492,In_1830,In_4736);
xnor U1493 (N_1493,In_3843,In_4358);
or U1494 (N_1494,N_693,In_3231);
nor U1495 (N_1495,N_542,In_4101);
nand U1496 (N_1496,In_1451,In_2032);
xor U1497 (N_1497,In_3381,In_1057);
or U1498 (N_1498,N_418,In_786);
nor U1499 (N_1499,In_367,N_135);
and U1500 (N_1500,In_3559,In_3319);
nand U1501 (N_1501,In_4357,N_280);
nand U1502 (N_1502,In_2279,N_1229);
and U1503 (N_1503,N_807,In_3552);
or U1504 (N_1504,In_791,N_1161);
or U1505 (N_1505,In_3383,In_3153);
nand U1506 (N_1506,N_1250,N_1387);
and U1507 (N_1507,In_2211,In_2451);
nand U1508 (N_1508,In_2467,In_4532);
nand U1509 (N_1509,N_985,In_1874);
and U1510 (N_1510,In_1833,In_1662);
nand U1511 (N_1511,In_2154,N_334);
xor U1512 (N_1512,In_3285,In_7);
or U1513 (N_1513,N_977,In_1532);
nor U1514 (N_1514,In_4590,N_559);
or U1515 (N_1515,N_849,N_1272);
nand U1516 (N_1516,N_304,In_614);
or U1517 (N_1517,N_297,In_1682);
or U1518 (N_1518,In_4239,In_1905);
nor U1519 (N_1519,In_1309,In_1304);
nand U1520 (N_1520,In_2486,In_4483);
nand U1521 (N_1521,N_1047,In_2917);
xor U1522 (N_1522,In_1561,In_2693);
nand U1523 (N_1523,In_1762,In_4426);
nor U1524 (N_1524,In_2577,In_2882);
and U1525 (N_1525,In_3779,In_4105);
nand U1526 (N_1526,In_3862,N_162);
and U1527 (N_1527,In_1161,In_4712);
and U1528 (N_1528,In_4046,In_3259);
nor U1529 (N_1529,In_165,N_1193);
nor U1530 (N_1530,In_4463,In_202);
or U1531 (N_1531,In_4271,N_327);
or U1532 (N_1532,In_1558,N_1071);
nor U1533 (N_1533,In_3253,In_4411);
nor U1534 (N_1534,In_1910,In_2381);
nand U1535 (N_1535,In_3570,In_3736);
nand U1536 (N_1536,In_402,N_1473);
or U1537 (N_1537,In_4241,In_1346);
and U1538 (N_1538,In_1725,In_2156);
nand U1539 (N_1539,N_207,In_782);
and U1540 (N_1540,N_1255,N_1237);
nand U1541 (N_1541,In_2479,In_4810);
nand U1542 (N_1542,N_658,N_1344);
or U1543 (N_1543,In_3482,In_302);
and U1544 (N_1544,N_966,N_837);
and U1545 (N_1545,In_3468,In_2989);
nor U1546 (N_1546,In_2948,N_1391);
nand U1547 (N_1547,N_378,In_3372);
xor U1548 (N_1548,N_830,In_3731);
nor U1549 (N_1549,N_646,N_37);
and U1550 (N_1550,N_1445,In_1293);
nand U1551 (N_1551,N_1115,In_950);
and U1552 (N_1552,In_1023,N_478);
nand U1553 (N_1553,In_4050,N_797);
or U1554 (N_1554,In_1336,In_4509);
nor U1555 (N_1555,N_1267,In_2183);
or U1556 (N_1556,In_4797,N_620);
xor U1557 (N_1557,In_2880,In_2285);
and U1558 (N_1558,In_4822,In_3530);
and U1559 (N_1559,In_4914,N_1066);
and U1560 (N_1560,In_2215,In_3832);
or U1561 (N_1561,N_1227,N_1368);
and U1562 (N_1562,N_410,N_279);
nand U1563 (N_1563,In_1992,In_4169);
or U1564 (N_1564,In_4359,N_367);
and U1565 (N_1565,In_1179,N_704);
or U1566 (N_1566,N_68,In_953);
nor U1567 (N_1567,In_2371,In_3059);
nand U1568 (N_1568,N_1280,In_4478);
nor U1569 (N_1569,N_1221,In_1228);
and U1570 (N_1570,In_251,In_3808);
xnor U1571 (N_1571,In_3504,In_609);
xnor U1572 (N_1572,In_1858,In_3510);
nand U1573 (N_1573,N_919,In_3937);
nor U1574 (N_1574,In_1431,In_280);
xor U1575 (N_1575,In_2236,In_3879);
nand U1576 (N_1576,N_774,In_4729);
nor U1577 (N_1577,In_684,N_846);
nor U1578 (N_1578,In_4158,N_1011);
or U1579 (N_1579,In_336,In_1963);
or U1580 (N_1580,In_1743,N_21);
and U1581 (N_1581,In_3767,N_1435);
or U1582 (N_1582,In_1462,In_1776);
or U1583 (N_1583,In_2890,In_4300);
nor U1584 (N_1584,In_240,In_397);
or U1585 (N_1585,N_1150,N_504);
and U1586 (N_1586,In_1707,In_3881);
xnor U1587 (N_1587,In_2635,In_4404);
or U1588 (N_1588,In_975,In_2936);
xnor U1589 (N_1589,In_1124,In_4363);
and U1590 (N_1590,In_3155,N_182);
xor U1591 (N_1591,In_381,In_2823);
nand U1592 (N_1592,N_1033,In_2387);
nor U1593 (N_1593,In_1800,In_2740);
xnor U1594 (N_1594,N_912,N_1114);
nand U1595 (N_1595,In_4747,In_3316);
nor U1596 (N_1596,In_4161,In_4723);
nor U1597 (N_1597,N_1048,In_3010);
and U1598 (N_1598,N_298,In_4032);
and U1599 (N_1599,In_2373,In_4086);
nand U1600 (N_1600,In_1423,In_3232);
nor U1601 (N_1601,In_2428,In_2551);
nor U1602 (N_1602,N_1409,In_1705);
nand U1603 (N_1603,N_57,In_2169);
or U1604 (N_1604,In_1616,In_2926);
nand U1605 (N_1605,N_372,In_3884);
or U1606 (N_1606,In_4443,N_146);
nor U1607 (N_1607,In_4742,N_928);
nor U1608 (N_1608,N_1080,N_1025);
or U1609 (N_1609,N_1256,N_177);
xor U1610 (N_1610,In_3909,N_724);
or U1611 (N_1611,In_2929,In_2377);
xor U1612 (N_1612,In_2949,N_1246);
nor U1613 (N_1613,In_1555,N_972);
and U1614 (N_1614,N_671,N_386);
and U1615 (N_1615,In_703,N_1101);
or U1616 (N_1616,In_2397,In_1724);
nand U1617 (N_1617,In_1667,In_984);
nand U1618 (N_1618,In_4000,In_2399);
or U1619 (N_1619,In_828,In_1965);
xnor U1620 (N_1620,In_1486,In_1015);
xor U1621 (N_1621,N_1451,N_880);
nand U1622 (N_1622,In_995,In_3321);
nand U1623 (N_1623,In_2556,N_1417);
or U1624 (N_1624,In_4107,In_2135);
xor U1625 (N_1625,In_3645,N_787);
xor U1626 (N_1626,In_1979,N_595);
and U1627 (N_1627,In_1823,In_16);
xnor U1628 (N_1628,In_2152,In_3757);
nor U1629 (N_1629,N_609,In_4226);
nand U1630 (N_1630,In_4309,N_1337);
nand U1631 (N_1631,In_673,N_1226);
nand U1632 (N_1632,In_3461,In_1723);
and U1633 (N_1633,In_2292,In_1310);
and U1634 (N_1634,N_1053,In_4195);
xnor U1635 (N_1635,In_840,N_1373);
and U1636 (N_1636,N_1298,In_1937);
nand U1637 (N_1637,In_4873,In_3542);
xnor U1638 (N_1638,N_1320,N_594);
nand U1639 (N_1639,In_338,N_1336);
nand U1640 (N_1640,In_1246,In_1252);
or U1641 (N_1641,In_3374,In_1240);
and U1642 (N_1642,In_2640,In_3981);
or U1643 (N_1643,In_2140,In_4180);
or U1644 (N_1644,In_1748,N_833);
nor U1645 (N_1645,In_2171,In_4669);
nand U1646 (N_1646,In_335,In_700);
and U1647 (N_1647,In_3416,In_3742);
nand U1648 (N_1648,In_698,N_864);
nand U1649 (N_1649,In_4073,In_3478);
xor U1650 (N_1650,N_16,In_625);
xor U1651 (N_1651,N_1077,In_4198);
nor U1652 (N_1652,In_1404,In_2787);
or U1653 (N_1653,In_3067,In_3675);
xor U1654 (N_1654,In_2319,N_856);
and U1655 (N_1655,In_2283,In_3617);
nand U1656 (N_1656,In_1499,In_2303);
and U1657 (N_1657,N_183,N_1326);
xnor U1658 (N_1658,In_2718,In_631);
and U1659 (N_1659,N_1313,In_1052);
or U1660 (N_1660,N_382,In_132);
or U1661 (N_1661,In_3266,N_638);
xnor U1662 (N_1662,In_916,In_2401);
and U1663 (N_1663,N_1200,In_2404);
xor U1664 (N_1664,In_2359,In_2348);
or U1665 (N_1665,In_3763,N_1089);
nand U1666 (N_1666,In_3822,In_80);
xnor U1667 (N_1667,N_248,N_854);
xor U1668 (N_1668,N_1384,N_482);
and U1669 (N_1669,In_168,In_596);
nor U1670 (N_1670,In_968,N_1009);
or U1671 (N_1671,N_1109,In_3624);
nor U1672 (N_1672,In_4112,In_1892);
nor U1673 (N_1673,In_899,N_401);
and U1674 (N_1674,N_78,N_158);
nand U1675 (N_1675,N_1263,In_3669);
or U1676 (N_1676,N_863,N_193);
and U1677 (N_1677,N_810,In_2827);
nand U1678 (N_1678,In_839,In_1042);
nor U1679 (N_1679,In_3483,In_1756);
and U1680 (N_1680,N_1305,N_1359);
or U1681 (N_1681,N_1211,In_3681);
and U1682 (N_1682,N_616,In_1498);
and U1683 (N_1683,In_560,N_720);
xor U1684 (N_1684,N_952,N_834);
nand U1685 (N_1685,In_2658,In_2674);
or U1686 (N_1686,In_4606,In_2582);
or U1687 (N_1687,In_2065,In_4646);
or U1688 (N_1688,N_794,In_2560);
or U1689 (N_1689,In_4816,In_1606);
nand U1690 (N_1690,N_463,In_3011);
nor U1691 (N_1691,N_178,In_4887);
nand U1692 (N_1692,N_1152,In_174);
and U1693 (N_1693,N_1324,In_3451);
or U1694 (N_1694,In_4644,In_4321);
or U1695 (N_1695,In_1138,In_654);
nor U1696 (N_1696,In_4058,N_399);
nand U1697 (N_1697,In_1580,In_2265);
nand U1698 (N_1698,In_3821,In_4108);
and U1699 (N_1699,In_4206,N_1428);
nor U1700 (N_1700,In_2876,N_631);
xor U1701 (N_1701,In_4079,N_800);
or U1702 (N_1702,N_1355,N_1470);
and U1703 (N_1703,In_4813,In_4768);
and U1704 (N_1704,In_1513,In_4076);
nand U1705 (N_1705,N_1455,In_2090);
or U1706 (N_1706,N_278,In_1068);
or U1707 (N_1707,N_436,N_130);
nor U1708 (N_1708,N_1151,In_1699);
nor U1709 (N_1709,In_3684,In_2869);
nor U1710 (N_1710,N_1153,N_316);
nor U1711 (N_1711,N_1319,In_870);
and U1712 (N_1712,In_495,In_777);
nand U1713 (N_1713,N_1195,N_543);
xnor U1714 (N_1714,N_855,N_811);
nor U1715 (N_1715,In_388,In_971);
or U1716 (N_1716,In_3298,In_4995);
nand U1717 (N_1717,In_723,In_3289);
nand U1718 (N_1718,In_209,In_784);
nor U1719 (N_1719,In_3993,In_2251);
and U1720 (N_1720,In_491,In_2328);
nor U1721 (N_1721,In_221,In_2902);
and U1722 (N_1722,In_3115,N_1129);
or U1723 (N_1723,In_1923,N_1423);
and U1724 (N_1724,In_2088,In_1502);
nor U1725 (N_1725,N_1341,In_4935);
nor U1726 (N_1726,In_1125,In_1801);
nor U1727 (N_1727,N_1058,In_3142);
and U1728 (N_1728,In_1117,In_4556);
nor U1729 (N_1729,In_2963,In_1195);
and U1730 (N_1730,In_239,In_4415);
xor U1731 (N_1731,In_40,N_1310);
nor U1732 (N_1732,In_2944,N_605);
and U1733 (N_1733,In_1856,N_1042);
nor U1734 (N_1734,N_371,In_2675);
nand U1735 (N_1735,N_292,N_32);
and U1736 (N_1736,In_1145,In_41);
nor U1737 (N_1737,In_1350,In_2375);
or U1738 (N_1738,In_1454,In_1226);
nor U1739 (N_1739,N_961,In_2837);
nand U1740 (N_1740,In_101,N_1163);
nor U1741 (N_1741,In_1612,In_3195);
nand U1742 (N_1742,In_3133,N_1145);
nand U1743 (N_1743,N_1349,In_4530);
or U1744 (N_1744,N_1427,N_447);
nand U1745 (N_1745,In_702,In_3927);
nor U1746 (N_1746,In_1772,N_1443);
or U1747 (N_1747,N_838,In_1663);
nand U1748 (N_1748,N_1148,In_4629);
or U1749 (N_1749,In_540,N_555);
nand U1750 (N_1750,In_1759,In_4981);
or U1751 (N_1751,N_1438,N_873);
and U1752 (N_1752,In_2176,In_3809);
nand U1753 (N_1753,N_743,In_2534);
and U1754 (N_1754,In_1174,In_1449);
nor U1755 (N_1755,In_4951,In_4987);
xor U1756 (N_1756,N_1421,In_4381);
nor U1757 (N_1757,In_3614,In_1793);
or U1758 (N_1758,In_2992,In_1075);
xor U1759 (N_1759,In_3520,In_1244);
xor U1760 (N_1760,In_1457,In_4749);
nand U1761 (N_1761,N_598,In_2842);
and U1762 (N_1762,In_2417,In_3224);
or U1763 (N_1763,In_1003,N_1060);
or U1764 (N_1764,N_561,N_337);
nor U1765 (N_1765,In_4990,In_1650);
and U1766 (N_1766,In_3554,N_920);
xnor U1767 (N_1767,N_1155,In_4734);
xor U1768 (N_1768,N_374,N_1454);
and U1769 (N_1769,In_3268,In_1670);
nand U1770 (N_1770,N_842,N_516);
nor U1771 (N_1771,In_4322,In_4837);
and U1772 (N_1772,N_534,N_1179);
nor U1773 (N_1773,N_1466,N_804);
nor U1774 (N_1774,In_4023,In_1638);
xnor U1775 (N_1775,In_1964,In_2550);
nor U1776 (N_1776,N_683,In_1162);
and U1777 (N_1777,N_1192,N_950);
nand U1778 (N_1778,In_4185,In_3977);
and U1779 (N_1779,In_1190,N_35);
nor U1780 (N_1780,In_2480,N_185);
xnor U1781 (N_1781,In_1803,In_3083);
or U1782 (N_1782,In_78,N_895);
nand U1783 (N_1783,In_4603,In_2080);
or U1784 (N_1784,N_1199,In_530);
nand U1785 (N_1785,N_435,In_4475);
nand U1786 (N_1786,In_3801,In_1674);
nand U1787 (N_1787,N_1307,In_4858);
or U1788 (N_1788,In_2570,In_4438);
nand U1789 (N_1789,N_319,In_902);
nand U1790 (N_1790,In_71,N_945);
nor U1791 (N_1791,In_2094,In_712);
xnor U1792 (N_1792,In_1872,In_321);
or U1793 (N_1793,N_579,In_297);
nand U1794 (N_1794,In_2916,In_1791);
xnor U1795 (N_1795,In_2203,N_320);
nor U1796 (N_1796,In_4650,N_593);
nor U1797 (N_1797,In_1151,In_1587);
or U1798 (N_1798,N_1219,In_4274);
and U1799 (N_1799,In_3546,In_2865);
xor U1800 (N_1800,In_2041,In_4460);
or U1801 (N_1801,In_1248,In_1890);
xnor U1802 (N_1802,In_2696,N_514);
nand U1803 (N_1803,In_3187,In_4298);
nand U1804 (N_1804,In_925,N_881);
nor U1805 (N_1805,N_1488,In_3553);
and U1806 (N_1806,In_1143,In_1721);
nand U1807 (N_1807,In_1595,In_2246);
and U1808 (N_1808,In_24,In_44);
nor U1809 (N_1809,In_3002,In_500);
nor U1810 (N_1810,N_1224,In_4080);
nand U1811 (N_1811,In_657,N_963);
and U1812 (N_1812,In_3094,In_3755);
nor U1813 (N_1813,In_3194,N_577);
xnor U1814 (N_1814,In_1871,In_276);
nand U1815 (N_1815,N_1007,N_970);
nand U1816 (N_1816,N_1383,N_648);
and U1817 (N_1817,N_885,In_4733);
nand U1818 (N_1818,N_1029,N_251);
nand U1819 (N_1819,In_2305,In_2721);
or U1820 (N_1820,In_5,N_527);
xnor U1821 (N_1821,In_1907,In_3151);
nand U1822 (N_1822,In_3800,In_2491);
xnor U1823 (N_1823,N_1225,In_247);
or U1824 (N_1824,In_983,N_1490);
nor U1825 (N_1825,In_1070,In_558);
nand U1826 (N_1826,In_1185,N_259);
nand U1827 (N_1827,N_624,N_580);
or U1828 (N_1828,N_536,In_1241);
or U1829 (N_1829,In_2758,N_458);
and U1830 (N_1830,N_1019,In_4980);
xor U1831 (N_1831,In_4572,N_753);
and U1832 (N_1832,N_168,In_903);
or U1833 (N_1833,N_727,In_2087);
nor U1834 (N_1834,In_3659,In_2722);
and U1835 (N_1835,N_1311,In_686);
and U1836 (N_1836,In_4256,N_1103);
xor U1837 (N_1837,In_300,N_1094);
nand U1838 (N_1838,In_4207,In_905);
or U1839 (N_1839,In_2282,In_860);
nor U1840 (N_1840,In_2443,In_4790);
and U1841 (N_1841,N_629,In_2179);
xor U1842 (N_1842,In_3395,In_287);
nand U1843 (N_1843,N_773,N_1169);
xnor U1844 (N_1844,In_3471,In_1737);
nand U1845 (N_1845,N_1330,In_4685);
nor U1846 (N_1846,N_377,N_105);
nor U1847 (N_1847,N_943,In_3393);
or U1848 (N_1848,N_1485,In_4210);
and U1849 (N_1849,N_1457,In_155);
nand U1850 (N_1850,N_1260,In_4929);
nor U1851 (N_1851,In_325,In_4403);
or U1852 (N_1852,In_3606,In_3680);
and U1853 (N_1853,N_1201,In_2314);
nor U1854 (N_1854,In_178,In_2788);
xor U1855 (N_1855,N_30,N_211);
xnor U1856 (N_1856,In_3315,In_1308);
and U1857 (N_1857,In_3118,N_1301);
xnor U1858 (N_1858,In_4868,In_1622);
and U1859 (N_1859,N_1400,In_1321);
and U1860 (N_1860,N_139,In_741);
nor U1861 (N_1861,In_1863,N_673);
or U1862 (N_1862,In_2192,In_456);
xor U1863 (N_1863,N_1141,In_978);
nor U1864 (N_1864,N_1189,In_1006);
nand U1865 (N_1865,N_1117,In_3209);
nand U1866 (N_1866,In_593,N_1068);
xor U1867 (N_1867,In_3995,In_3085);
nand U1868 (N_1868,In_2497,N_475);
and U1869 (N_1869,In_3302,In_3894);
xor U1870 (N_1870,N_1035,In_1995);
and U1871 (N_1871,In_372,N_1134);
or U1872 (N_1872,In_976,In_1543);
nor U1873 (N_1873,In_2561,In_4789);
and U1874 (N_1874,N_92,In_2682);
nand U1875 (N_1875,In_2873,In_3265);
nor U1876 (N_1876,N_405,N_1499);
nor U1877 (N_1877,In_33,In_568);
or U1878 (N_1878,In_1259,In_4194);
nor U1879 (N_1879,In_4974,N_1001);
xor U1880 (N_1880,N_333,In_2514);
nor U1881 (N_1881,In_4388,N_1149);
xor U1882 (N_1882,In_4395,In_430);
nand U1883 (N_1883,In_4821,In_117);
or U1884 (N_1884,In_3942,In_3182);
nand U1885 (N_1885,In_2891,N_1247);
nand U1886 (N_1886,In_2683,N_968);
and U1887 (N_1887,In_3734,N_425);
xor U1888 (N_1888,In_4814,In_3696);
xor U1889 (N_1889,In_2614,N_1107);
or U1890 (N_1890,In_2988,N_947);
nor U1891 (N_1891,In_918,In_3044);
and U1892 (N_1892,N_380,N_1165);
nand U1893 (N_1893,In_3714,In_1557);
nand U1894 (N_1894,In_4539,N_1140);
and U1895 (N_1895,N_1044,In_472);
nor U1896 (N_1896,In_152,In_3695);
xnor U1897 (N_1897,In_4508,In_3844);
or U1898 (N_1898,In_2037,In_4447);
nand U1899 (N_1899,N_843,In_2052);
nand U1900 (N_1900,In_2014,In_1540);
xor U1901 (N_1901,In_868,In_3630);
or U1902 (N_1902,In_1976,N_584);
or U1903 (N_1903,In_2458,In_1358);
nand U1904 (N_1904,In_498,N_301);
nand U1905 (N_1905,N_485,In_3437);
nor U1906 (N_1906,In_3853,In_204);
nand U1907 (N_1907,In_2752,N_1054);
nor U1908 (N_1908,N_652,N_239);
nand U1909 (N_1909,In_3106,In_647);
xor U1910 (N_1910,In_4947,In_2123);
nand U1911 (N_1911,N_1098,In_3940);
and U1912 (N_1912,In_201,In_4824);
nand U1913 (N_1913,In_3075,In_774);
or U1914 (N_1914,In_954,N_1174);
nor U1915 (N_1915,N_466,N_1350);
xor U1916 (N_1916,N_1171,N_510);
nor U1917 (N_1917,In_3599,In_442);
nor U1918 (N_1918,N_1446,N_1100);
nor U1919 (N_1919,In_3652,In_4663);
and U1920 (N_1920,In_4920,In_4281);
nor U1921 (N_1921,N_331,N_1498);
nand U1922 (N_1922,In_2794,In_1602);
nor U1923 (N_1923,N_1397,N_284);
nor U1924 (N_1924,In_565,In_3798);
nor U1925 (N_1925,N_979,In_1741);
nand U1926 (N_1926,In_4196,In_3730);
xor U1927 (N_1927,N_836,In_27);
and U1928 (N_1928,In_4166,N_205);
xnor U1929 (N_1929,In_4540,In_2986);
and U1930 (N_1930,In_61,In_4991);
or U1931 (N_1931,In_2398,In_1985);
nand U1932 (N_1932,In_506,In_3273);
xnor U1933 (N_1933,In_3983,In_4787);
xor U1934 (N_1934,N_781,In_1016);
and U1935 (N_1935,N_827,N_847);
xnor U1936 (N_1936,N_782,In_477);
and U1937 (N_1937,In_253,In_3621);
nor U1938 (N_1938,In_3970,N_745);
nand U1939 (N_1939,N_1031,In_783);
or U1940 (N_1940,In_2796,In_592);
or U1941 (N_1941,N_110,In_693);
or U1942 (N_1942,N_268,N_988);
nand U1943 (N_1943,In_748,In_965);
nand U1944 (N_1944,In_1579,In_3040);
xnor U1945 (N_1945,In_1232,In_4799);
and U1946 (N_1946,N_956,N_326);
and U1947 (N_1947,N_725,In_1153);
and U1948 (N_1948,In_2730,N_1388);
and U1949 (N_1949,In_2017,In_4904);
nor U1950 (N_1950,In_3796,In_1969);
or U1951 (N_1951,In_2150,N_420);
nand U1952 (N_1952,In_4999,N_1477);
and U1953 (N_1953,In_1243,N_1469);
and U1954 (N_1954,In_1133,N_60);
xor U1955 (N_1955,In_842,In_1412);
nor U1956 (N_1956,N_1131,N_1461);
nor U1957 (N_1957,N_440,N_473);
and U1958 (N_1958,In_2808,N_1002);
nand U1959 (N_1959,N_583,In_270);
and U1960 (N_1960,In_258,N_263);
xor U1961 (N_1961,In_1047,N_799);
nand U1962 (N_1962,In_163,In_3440);
nand U1963 (N_1963,In_2028,In_721);
xnor U1964 (N_1964,N_1018,In_2753);
nor U1965 (N_1965,In_110,In_3777);
xor U1966 (N_1966,In_3774,In_4872);
xor U1967 (N_1967,In_4956,In_542);
xnor U1968 (N_1968,In_4485,In_4584);
xor U1969 (N_1969,In_2366,In_636);
nor U1970 (N_1970,N_27,In_383);
or U1971 (N_1971,In_1326,N_672);
nand U1972 (N_1972,In_820,In_1021);
nand U1973 (N_1973,In_1101,In_2862);
nor U1974 (N_1974,N_1363,In_2528);
and U1975 (N_1975,In_600,In_1831);
and U1976 (N_1976,In_4088,In_4806);
nor U1977 (N_1977,In_1461,In_3895);
or U1978 (N_1978,In_1215,In_181);
nand U1979 (N_1979,In_4128,In_3491);
nor U1980 (N_1980,In_1168,In_4510);
or U1981 (N_1981,In_824,N_1406);
xor U1982 (N_1982,N_1196,In_594);
nor U1983 (N_1983,N_479,In_669);
and U1984 (N_1984,In_4143,In_339);
nor U1985 (N_1985,In_4164,In_4301);
or U1986 (N_1986,N_1372,N_133);
nand U1987 (N_1987,In_2709,In_2568);
xnor U1988 (N_1988,N_1218,N_309);
xnor U1989 (N_1989,In_334,In_2194);
and U1990 (N_1990,N_1143,In_1137);
nor U1991 (N_1991,N_25,N_1178);
nor U1992 (N_1992,In_3189,In_1521);
or U1993 (N_1993,In_1991,In_1978);
and U1994 (N_1994,In_2298,In_144);
and U1995 (N_1995,N_1070,In_4235);
or U1996 (N_1996,N_127,In_4124);
nor U1997 (N_1997,In_1218,In_1531);
or U1998 (N_1998,In_3058,N_1234);
xor U1999 (N_1999,In_1085,In_350);
and U2000 (N_2000,N_1212,N_1828);
and U2001 (N_2001,N_1644,N_1204);
nor U2002 (N_2002,In_3892,N_627);
and U2003 (N_2003,N_1444,In_2074);
and U2004 (N_2004,In_4559,N_969);
nor U2005 (N_2005,In_2999,N_1905);
xnor U2006 (N_2006,N_980,In_838);
and U2007 (N_2007,N_1713,In_3835);
nand U2008 (N_2008,N_1886,In_1891);
nand U2009 (N_2009,In_890,N_1594);
nor U2010 (N_2010,In_232,In_3527);
xor U2011 (N_2011,In_4780,In_1708);
nor U2012 (N_2012,In_1427,N_1616);
and U2013 (N_2013,In_3333,In_4203);
nand U2014 (N_2014,N_1422,In_809);
nor U2015 (N_2015,In_3974,N_1971);
and U2016 (N_2016,N_1198,In_2965);
xor U2017 (N_2017,In_1391,In_3376);
and U2018 (N_2018,In_4406,N_1957);
or U2019 (N_2019,In_3163,N_1291);
nor U2020 (N_2020,N_1617,In_1108);
nand U2021 (N_2021,In_1735,In_3415);
nor U2022 (N_2022,N_1663,N_1015);
xor U2023 (N_2023,In_2260,In_2781);
and U2024 (N_2024,In_3521,N_1899);
nand U2025 (N_2025,In_4213,In_2650);
and U2026 (N_2026,N_1425,N_1823);
nand U2027 (N_2027,In_3768,N_1282);
nor U2028 (N_2028,N_1529,In_3907);
xor U2029 (N_2029,N_1630,In_692);
or U2030 (N_2030,N_1038,N_1814);
or U2031 (N_2031,N_1640,In_2316);
or U2032 (N_2032,In_4758,N_1442);
and U2033 (N_2033,In_1837,In_182);
nand U2034 (N_2034,In_2938,In_3193);
nand U2035 (N_2035,In_3159,In_1660);
and U2036 (N_2036,In_3263,In_3250);
xnor U2037 (N_2037,In_2232,In_2418);
or U2038 (N_2038,In_2354,N_1792);
xor U2039 (N_2039,In_1186,N_131);
or U2040 (N_2040,N_680,N_777);
or U2041 (N_2041,N_1973,In_3776);
xnor U2042 (N_2042,In_11,N_1603);
nand U2043 (N_2043,In_85,N_897);
xor U2044 (N_2044,In_1537,N_1075);
xor U2045 (N_2045,N_1673,In_3702);
nor U2046 (N_2046,N_431,N_289);
nor U2047 (N_2047,In_4893,N_1340);
or U2048 (N_2048,In_109,In_2901);
nand U2049 (N_2049,In_2732,N_299);
and U2050 (N_2050,N_1577,In_3062);
or U2051 (N_2051,In_3441,N_1206);
nand U2052 (N_2052,N_1168,N_647);
xor U2053 (N_2053,In_3105,N_1133);
or U2054 (N_2054,In_3547,N_659);
xor U2055 (N_2055,In_2036,N_1785);
nor U2056 (N_2056,N_637,In_3450);
nor U2057 (N_2057,N_1286,N_1184);
or U2058 (N_2058,In_2446,N_1412);
nand U2059 (N_2059,In_1853,N_1289);
nor U2060 (N_2060,N_1612,N_1586);
and U2061 (N_2061,In_100,In_3097);
xor U2062 (N_2062,N_718,In_1013);
xor U2063 (N_2063,In_1528,In_279);
or U2064 (N_2064,In_1695,N_870);
or U2065 (N_2065,N_1587,In_3005);
xor U2066 (N_2066,N_1562,In_3127);
and U2067 (N_2067,In_2395,In_97);
and U2068 (N_2068,In_4139,In_4591);
or U2069 (N_2069,In_1189,In_1495);
nand U2070 (N_2070,N_1284,In_2909);
xor U2071 (N_2071,In_3305,In_386);
and U2072 (N_2072,In_571,In_4199);
and U2073 (N_2073,In_3759,In_2362);
nor U2074 (N_2074,N_965,In_299);
nand U2075 (N_2075,In_993,N_340);
xor U2076 (N_2076,In_1385,N_1241);
nor U2077 (N_2077,N_1393,In_1729);
xor U2078 (N_2078,N_20,N_1596);
and U2079 (N_2079,In_3286,N_1657);
and U2080 (N_2080,In_2661,In_4930);
nor U2081 (N_2081,N_163,In_3071);
nand U2082 (N_2082,N_1074,N_521);
and U2083 (N_2083,N_1652,N_1123);
nor U2084 (N_2084,In_2471,In_793);
xor U2085 (N_2085,In_343,In_2218);
and U2086 (N_2086,N_894,In_1880);
nand U2087 (N_2087,N_1979,N_737);
nand U2088 (N_2088,In_1492,In_3787);
xnor U2089 (N_2089,N_465,In_3197);
xnor U2090 (N_2090,N_1530,In_2227);
nand U2091 (N_2091,In_4126,In_4656);
nor U2092 (N_2092,N_1118,In_645);
nor U2093 (N_2093,N_1618,N_1811);
nor U2094 (N_2094,In_1763,N_1687);
xnor U2095 (N_2095,In_3791,In_2178);
xor U2096 (N_2096,N_1420,In_981);
nor U2097 (N_2097,N_6,In_3938);
nor U2098 (N_2098,N_1097,N_1874);
nand U2099 (N_2099,In_39,N_1087);
xor U2100 (N_2100,N_709,N_359);
or U2101 (N_2101,N_1669,In_4876);
xnor U2102 (N_2102,In_156,In_2165);
and U2103 (N_2103,In_624,N_1795);
nand U2104 (N_2104,N_1448,In_1091);
nor U2105 (N_2105,N_1726,In_1027);
xor U2106 (N_2106,In_2188,N_1760);
xor U2107 (N_2107,N_1126,In_2465);
nor U2108 (N_2108,N_1916,N_1911);
and U2109 (N_2109,N_1995,In_1387);
or U2110 (N_2110,N_1659,N_453);
xnor U2111 (N_2111,N_778,In_3064);
nand U2112 (N_2112,In_3869,In_1067);
or U2113 (N_2113,N_1877,In_1424);
xnor U2114 (N_2114,In_2883,N_571);
or U2115 (N_2115,N_1733,N_1798);
nor U2116 (N_2116,N_1782,In_3117);
nor U2117 (N_2117,In_3045,In_2841);
xor U2118 (N_2118,In_2920,N_1385);
and U2119 (N_2119,In_1324,In_1973);
xor U2120 (N_2120,In_4618,In_4589);
or U2121 (N_2121,N_911,In_3689);
nor U2122 (N_2122,In_4511,In_982);
nand U2123 (N_2123,In_4182,In_2454);
nand U2124 (N_2124,In_1896,N_1935);
xor U2125 (N_2125,In_226,In_1857);
xor U2126 (N_2126,N_1239,In_766);
and U2127 (N_2127,N_1034,In_3806);
nor U2128 (N_2128,N_1922,In_2424);
nand U2129 (N_2129,In_867,In_1806);
nor U2130 (N_2130,In_778,In_2255);
nand U2131 (N_2131,In_4988,In_4430);
and U2132 (N_2132,N_1944,N_1032);
xor U2133 (N_2133,In_1106,In_1882);
nor U2134 (N_2134,In_548,N_1364);
nand U2135 (N_2135,In_2881,In_3720);
or U2136 (N_2136,N_1315,In_1952);
nand U2137 (N_2137,N_283,In_1653);
nand U2138 (N_2138,N_1285,N_1749);
or U2139 (N_2139,N_489,N_1519);
or U2140 (N_2140,In_2063,In_1703);
or U2141 (N_2141,In_357,In_3576);
xnor U2142 (N_2142,In_831,In_3453);
and U2143 (N_2143,In_4284,N_1050);
and U2144 (N_2144,N_1549,In_1351);
and U2145 (N_2145,N_1411,In_1966);
nand U2146 (N_2146,N_220,N_1615);
or U2147 (N_2147,N_525,In_588);
and U2148 (N_2148,In_2932,N_546);
xor U2149 (N_2149,In_438,In_4240);
nand U2150 (N_2150,In_1058,In_2589);
nand U2151 (N_2151,In_4222,N_1667);
xnor U2152 (N_2152,N_1346,In_4757);
xnor U2153 (N_2153,In_4219,In_4687);
and U2154 (N_2154,In_4655,In_1038);
xnor U2155 (N_2155,N_1261,N_1860);
xnor U2156 (N_2156,In_961,In_3439);
nand U2157 (N_2157,In_3391,N_1022);
and U2158 (N_2158,In_4056,In_3175);
nor U2159 (N_2159,In_1809,In_4264);
nand U2160 (N_2160,In_3836,N_617);
or U2161 (N_2161,In_4019,In_3788);
nand U2162 (N_2162,In_814,N_1841);
or U2163 (N_2163,N_1614,In_3535);
nand U2164 (N_2164,In_2300,N_1505);
and U2165 (N_2165,N_126,In_401);
xor U2166 (N_2166,N_755,N_1410);
or U2167 (N_2167,In_4257,N_1972);
xor U2168 (N_2168,In_587,In_935);
nor U2169 (N_2169,In_1074,N_1538);
nand U2170 (N_2170,In_1690,N_502);
nand U2171 (N_2171,In_288,In_1378);
xnor U2172 (N_2172,In_725,In_243);
nand U2173 (N_2173,N_1173,In_639);
xnor U2174 (N_2174,N_762,N_1819);
nor U2175 (N_2175,In_3029,N_1496);
nand U2176 (N_2176,In_3592,In_4214);
xnor U2177 (N_2177,In_4280,In_2576);
nor U2178 (N_2178,N_1249,In_3053);
or U2179 (N_2179,N_1278,In_4400);
and U2180 (N_2180,In_4719,In_1181);
nor U2181 (N_2181,In_2708,In_111);
xnor U2182 (N_2182,In_1315,N_1605);
or U2183 (N_2183,N_408,In_3485);
and U2184 (N_2184,In_1251,N_1637);
or U2185 (N_2185,N_761,In_4522);
and U2186 (N_2186,In_2666,In_3387);
nand U2187 (N_2187,N_1106,In_4029);
xor U2188 (N_2188,N_1479,In_3551);
or U2189 (N_2189,In_3408,N_702);
nand U2190 (N_2190,N_164,In_3505);
xor U2191 (N_2191,In_744,In_2143);
or U2192 (N_2192,In_3037,In_2393);
and U2193 (N_2193,N_1102,In_834);
and U2194 (N_2194,N_1744,In_3783);
and U2195 (N_2195,In_2700,In_4910);
or U2196 (N_2196,In_2067,In_1916);
or U2197 (N_2197,In_3414,N_1697);
nand U2198 (N_2198,N_1848,In_4538);
and U2199 (N_2199,In_2738,In_1408);
xor U2200 (N_2200,N_84,N_1240);
or U2201 (N_2201,In_304,In_2420);
nand U2202 (N_2202,In_539,N_1205);
nand U2203 (N_2203,In_4327,N_1789);
nand U2204 (N_2204,In_431,In_3188);
or U2205 (N_2205,N_1046,In_3091);
nand U2206 (N_2206,In_1134,In_3886);
and U2207 (N_2207,In_1083,In_2308);
nor U2208 (N_2208,In_1262,N_551);
nand U2209 (N_2209,N_416,In_2043);
nand U2210 (N_2210,In_1237,N_285);
or U2211 (N_2211,In_854,In_932);
or U2212 (N_2212,N_172,In_4270);
nand U2213 (N_2213,In_1079,In_581);
nand U2214 (N_2214,N_1306,In_3400);
or U2215 (N_2215,N_1521,N_1774);
nor U2216 (N_2216,In_893,N_841);
xor U2217 (N_2217,In_453,In_4418);
or U2218 (N_2218,N_1607,N_1660);
xnor U2219 (N_2219,N_1960,N_1559);
nor U2220 (N_2220,In_4474,N_759);
and U2221 (N_2221,N_618,N_1925);
nand U2222 (N_2222,N_971,N_1868);
or U2223 (N_2223,N_1555,In_3988);
and U2224 (N_2224,In_3138,In_3462);
and U2225 (N_2225,N_1907,N_622);
xor U2226 (N_2226,N_1674,N_1917);
nor U2227 (N_2227,N_1331,In_503);
xor U2228 (N_2228,N_1459,N_1820);
and U2229 (N_2229,In_1948,N_1724);
nor U2230 (N_2230,In_3514,In_4850);
or U2231 (N_2231,In_1072,In_4480);
nor U2232 (N_2232,N_625,In_2148);
and U2233 (N_2233,N_1497,In_980);
and U2234 (N_2234,N_381,N_1950);
xnor U2235 (N_2235,In_2262,In_4616);
nand U2236 (N_2236,In_1754,In_3147);
or U2237 (N_2237,N_1191,N_567);
nand U2238 (N_2238,N_1745,In_3109);
xor U2239 (N_2239,In_3605,In_909);
nand U2240 (N_2240,N_1366,In_2596);
nand U2241 (N_2241,N_1378,In_2530);
or U2242 (N_2242,N_129,N_52);
and U2243 (N_2243,N_1808,N_1354);
or U2244 (N_2244,N_1535,N_1863);
nor U2245 (N_2245,N_1804,N_1351);
nor U2246 (N_2246,In_2083,In_4661);
xor U2247 (N_2247,N_689,N_1158);
nor U2248 (N_2248,N_1684,In_3371);
nand U2249 (N_2249,In_695,N_871);
or U2250 (N_2250,N_1997,N_1990);
or U2251 (N_2251,N_892,N_1550);
and U2252 (N_2252,N_1052,N_198);
nand U2253 (N_2253,In_2068,In_511);
and U2254 (N_2254,In_3863,In_3697);
nor U2255 (N_2255,In_1747,In_3411);
and U2256 (N_2256,In_3322,N_1276);
and U2257 (N_2257,In_484,N_1419);
nand U2258 (N_2258,In_4826,N_56);
nand U2259 (N_2259,N_124,In_4064);
and U2260 (N_2260,In_4892,In_4188);
nor U2261 (N_2261,N_1881,N_423);
xor U2262 (N_2262,In_3447,N_722);
xor U2263 (N_2263,N_1861,In_2207);
nand U2264 (N_2264,In_1997,N_1871);
nor U2265 (N_2265,In_919,In_4276);
nand U2266 (N_2266,N_1921,In_4288);
nand U2267 (N_2267,N_1472,In_525);
xor U2268 (N_2268,In_1984,N_1898);
nor U2269 (N_2269,N_1902,In_4427);
nor U2270 (N_2270,In_1007,In_4626);
or U2271 (N_2271,N_1539,N_1028);
xnor U2272 (N_2272,In_3032,In_4693);
nand U2273 (N_2273,N_1269,In_4315);
or U2274 (N_2274,N_1494,In_1100);
or U2275 (N_2275,In_4186,In_63);
nor U2276 (N_2276,N_1680,N_1611);
xor U2277 (N_2277,N_1253,N_1965);
or U2278 (N_2278,N_1735,In_1702);
xor U2279 (N_2279,In_3190,In_3078);
nand U2280 (N_2280,In_891,N_1124);
or U2281 (N_2281,N_1283,In_4282);
xor U2282 (N_2282,In_635,In_3);
nand U2283 (N_2283,In_1225,N_1413);
xor U2284 (N_2284,In_715,N_1401);
xnor U2285 (N_2285,N_1867,In_585);
and U2286 (N_2286,In_4385,N_77);
and U2287 (N_2287,N_917,In_2430);
nand U2288 (N_2288,N_1251,In_2197);
nor U2289 (N_2289,N_1274,In_4576);
nor U2290 (N_2290,In_3409,In_4442);
xnor U2291 (N_2291,In_1975,In_2061);
or U2292 (N_2292,N_189,N_1099);
nor U2293 (N_2293,In_1337,In_429);
or U2294 (N_2294,N_643,N_332);
xor U2295 (N_2295,In_736,In_4092);
or U2296 (N_2296,In_2263,In_960);
and U2297 (N_2297,In_3104,N_754);
or U2298 (N_2298,In_4704,N_690);
or U2299 (N_2299,N_1092,N_167);
or U2300 (N_2300,N_1748,N_1138);
nor U2301 (N_2301,N_411,In_3667);
xor U2302 (N_2302,N_28,In_848);
nand U2303 (N_2303,N_1458,In_1382);
and U2304 (N_2304,In_2429,In_4841);
or U2305 (N_2305,In_4727,N_1999);
nand U2306 (N_2306,In_718,In_4544);
xnor U2307 (N_2307,N_1216,In_3963);
nor U2308 (N_2308,In_2367,N_1197);
and U2309 (N_2309,In_1355,In_1839);
nand U2310 (N_2310,In_1941,In_666);
and U2311 (N_2311,In_3579,In_597);
nand U2312 (N_2312,In_4350,In_3276);
or U2313 (N_2313,N_1758,In_4957);
or U2314 (N_2314,In_1330,N_1547);
or U2315 (N_2315,In_1643,N_628);
or U2316 (N_2316,N_1962,In_137);
nand U2317 (N_2317,In_1529,N_1433);
nand U2318 (N_2318,In_2710,N_1527);
xnor U2319 (N_2319,In_3660,In_576);
and U2320 (N_2320,In_1526,N_1716);
and U2321 (N_2321,N_1981,N_229);
nor U2322 (N_2322,N_982,N_1554);
and U2323 (N_2323,In_1943,In_2817);
xnor U2324 (N_2324,In_345,In_387);
nor U2325 (N_2325,N_1369,In_454);
nor U2326 (N_2326,In_2928,N_1938);
nor U2327 (N_2327,In_2628,N_484);
or U2328 (N_2328,In_2021,In_4832);
or U2329 (N_2329,In_3877,In_1149);
nor U2330 (N_2330,In_4839,In_1642);
and U2331 (N_2331,In_2160,In_567);
nor U2332 (N_2332,In_3299,In_4628);
nand U2333 (N_2333,In_2116,In_3282);
nand U2334 (N_2334,In_4386,In_3074);
or U2335 (N_2335,In_246,N_1086);
nor U2336 (N_2336,In_4379,N_663);
and U2337 (N_2337,N_1910,In_4122);
or U2338 (N_2338,N_1055,In_4066);
nand U2339 (N_2339,N_636,In_400);
nand U2340 (N_2340,In_2464,In_513);
nand U2341 (N_2341,In_1503,In_3813);
or U2342 (N_2342,In_3166,In_2982);
nor U2343 (N_2343,In_2072,In_3222);
nor U2344 (N_2344,In_3314,In_3196);
nor U2345 (N_2345,N_1091,In_4864);
nand U2346 (N_2346,N_1418,In_3324);
nand U2347 (N_2347,N_1185,In_882);
nor U2348 (N_2348,In_4751,In_4570);
or U2349 (N_2349,In_2252,In_1746);
nand U2350 (N_2350,In_17,In_3805);
and U2351 (N_2351,In_1559,In_1422);
nand U2352 (N_2352,N_1599,In_2274);
or U2353 (N_2353,N_1453,In_3452);
or U2354 (N_2354,In_682,In_3272);
and U2355 (N_2355,In_3585,N_1984);
and U2356 (N_2356,In_2631,N_1348);
nor U2357 (N_2357,N_1486,In_4059);
xor U2358 (N_2358,In_4527,N_1180);
nand U2359 (N_2359,In_69,In_4861);
and U2360 (N_2360,N_1837,N_1290);
or U2361 (N_2361,N_1356,N_42);
or U2362 (N_2362,N_1509,In_1931);
nand U2363 (N_2363,N_796,In_4434);
nand U2364 (N_2364,In_4348,N_1753);
or U2365 (N_2365,In_266,N_1629);
nand U2366 (N_2366,N_222,N_748);
and U2367 (N_2367,N_548,N_1426);
nand U2368 (N_2368,N_76,In_4691);
or U2369 (N_2369,N_281,In_2655);
or U2370 (N_2370,N_1686,N_740);
xor U2371 (N_2371,N_1913,N_707);
nor U2372 (N_2372,In_515,N_1665);
or U2373 (N_2373,In_3665,In_2975);
nor U2374 (N_2374,In_3181,In_2760);
xnor U2375 (N_2375,In_1694,N_282);
nor U2376 (N_2376,In_3470,N_1259);
nand U2377 (N_2377,N_1772,In_4621);
and U2378 (N_2378,N_1016,In_4707);
nor U2379 (N_2379,N_99,In_3637);
nor U2380 (N_2380,In_3956,In_4805);
xor U2381 (N_2381,N_1642,In_622);
and U2382 (N_2382,N_1790,In_2605);
nor U2383 (N_2383,In_3707,In_1618);
and U2384 (N_2384,In_4087,N_944);
or U2385 (N_2385,In_3643,In_3706);
and U2386 (N_2386,In_3994,N_1878);
nand U2387 (N_2387,N_1403,N_494);
nor U2388 (N_2388,In_3239,N_1974);
or U2389 (N_2389,N_942,N_967);
or U2390 (N_2390,In_4401,N_955);
nand U2391 (N_2391,In_4648,In_149);
xor U2392 (N_2392,In_1257,In_4888);
nor U2393 (N_2393,N_1480,In_738);
nand U2394 (N_2394,N_1010,In_2374);
nand U2395 (N_2395,N_430,In_4623);
and U2396 (N_2396,In_4171,In_1689);
nor U2397 (N_2397,N_1362,In_3803);
and U2398 (N_2398,N_875,In_2172);
xnor U2399 (N_2399,In_3810,In_2637);
nand U2400 (N_2400,In_4714,In_4075);
xor U2401 (N_2401,In_3498,N_1851);
or U2402 (N_2402,N_1928,N_1856);
nor U2403 (N_2403,N_662,N_934);
and U2404 (N_2404,In_4136,N_569);
and U2405 (N_2405,In_1753,In_1178);
or U2406 (N_2406,N_1623,N_214);
or U2407 (N_2407,In_99,In_141);
nand U2408 (N_2408,N_1656,In_1541);
nor U2409 (N_2409,In_4954,In_3674);
xor U2410 (N_2410,N_566,In_285);
nand U2411 (N_2411,In_720,N_1706);
or U2412 (N_2412,In_158,N_1424);
and U2413 (N_2413,In_2775,In_3096);
xor U2414 (N_2414,N_1793,In_1835);
or U2415 (N_2415,N_1013,N_1845);
nand U2416 (N_2416,In_2105,In_2272);
xor U2417 (N_2417,In_3838,In_3241);
nor U2418 (N_2418,N_1711,N_296);
nor U2419 (N_2419,In_3001,N_1317);
and U2420 (N_2420,N_1342,In_3782);
nand U2421 (N_2421,In_4550,N_1915);
and U2422 (N_2422,In_641,In_857);
nand U2423 (N_2423,In_3244,In_368);
xnor U2424 (N_2424,In_4933,N_1210);
xor U2425 (N_2425,In_3916,In_420);
nor U2426 (N_2426,N_528,N_1523);
nor U2427 (N_2427,N_1815,N_817);
xnor U2428 (N_2428,N_323,N_1604);
or U2429 (N_2429,In_2533,In_4265);
nand U2430 (N_2430,N_1941,In_271);
or U2431 (N_2431,N_845,In_2069);
nand U2432 (N_2432,In_939,In_3828);
nor U2433 (N_2433,N_1689,In_361);
and U2434 (N_2434,In_3816,In_1982);
nand U2435 (N_2435,In_2818,N_1736);
or U2436 (N_2436,N_1737,N_816);
and U2437 (N_2437,In_4439,In_3678);
xor U2438 (N_2438,N_1456,In_189);
nand U2439 (N_2439,N_79,N_656);
xnor U2440 (N_2440,In_2327,N_1670);
nand U2441 (N_2441,N_1039,In_2506);
or U2442 (N_2442,N_141,In_3851);
and U2443 (N_2443,In_3056,N_1405);
nand U2444 (N_2444,N_138,In_2904);
nor U2445 (N_2445,N_247,In_3086);
nor U2446 (N_2446,In_84,N_228);
or U2447 (N_2447,In_2813,N_1727);
and U2448 (N_2448,In_3899,N_364);
or U2449 (N_2449,In_504,N_1112);
or U2450 (N_2450,In_25,In_3281);
nor U2451 (N_2451,In_4908,N_1365);
xnor U2452 (N_2452,In_1090,N_1213);
xnor U2453 (N_2453,In_392,N_1606);
or U2454 (N_2454,N_993,In_1520);
or U2455 (N_2455,In_4501,N_1183);
or U2456 (N_2456,In_2748,In_2230);
nand U2457 (N_2457,In_471,In_4803);
and U2458 (N_2458,In_122,In_3786);
or U2459 (N_2459,In_1279,In_3543);
nand U2460 (N_2460,N_815,N_1432);
nand U2461 (N_2461,In_3662,In_2699);
and U2462 (N_2462,In_4614,In_2913);
and U2463 (N_2463,In_4836,N_288);
or U2464 (N_2464,In_4808,N_1989);
nor U2465 (N_2465,N_1352,In_2023);
and U2466 (N_2466,In_898,N_255);
and U2467 (N_2467,In_2871,In_3206);
nor U2468 (N_2468,In_4369,In_4561);
xnor U2469 (N_2469,In_2261,In_2407);
or U2470 (N_2470,In_2412,In_419);
nand U2471 (N_2471,In_2544,In_728);
and U2472 (N_2472,N_915,In_3718);
and U2473 (N_2473,In_3732,N_635);
xor U2474 (N_2474,In_96,In_2271);
or U2475 (N_2475,In_4895,N_1090);
xnor U2476 (N_2476,In_2851,N_1396);
xor U2477 (N_2477,N_601,N_1452);
and U2478 (N_2478,In_4278,N_1762);
or U2479 (N_2479,In_544,In_3728);
nand U2480 (N_2480,N_1954,In_2346);
and U2481 (N_2481,N_120,In_2689);
and U2482 (N_2482,N_1177,In_3766);
nor U2483 (N_2483,N_1436,In_1755);
and U2484 (N_2484,N_676,In_1064);
nand U2485 (N_2485,N_174,N_221);
and U2486 (N_2486,N_1951,In_4081);
or U2487 (N_2487,In_4202,N_1967);
or U2488 (N_2488,In_2927,N_633);
or U2489 (N_2489,In_4476,N_888);
or U2490 (N_2490,N_711,N_728);
xor U2491 (N_2491,In_3901,In_497);
nand U2492 (N_2492,In_4857,In_3436);
and U2493 (N_2493,N_1572,N_43);
xnor U2494 (N_2494,N_805,N_1631);
xnor U2495 (N_2495,In_2269,In_475);
or U2496 (N_2496,N_793,N_1347);
nand U2497 (N_2497,In_4611,In_3328);
xnor U2498 (N_2498,In_2887,In_963);
nand U2499 (N_2499,N_1575,In_4490);
or U2500 (N_2500,N_2188,In_3015);
xor U2501 (N_2501,In_4102,N_1244);
nand U2502 (N_2502,N_1756,N_498);
nand U2503 (N_2503,In_328,N_1721);
xor U2504 (N_2504,N_1932,In_1732);
xnor U2505 (N_2505,N_2236,N_1649);
or U2506 (N_2506,N_1818,In_315);
or U2507 (N_2507,N_687,N_1740);
or U2508 (N_2508,In_4244,N_1020);
and U2509 (N_2509,N_70,In_1949);
or U2510 (N_2510,N_2058,In_1484);
xnor U2511 (N_2511,In_1766,N_2292);
nand U2512 (N_2512,N_45,N_1514);
nor U2513 (N_2513,In_54,N_250);
xnor U2514 (N_2514,In_3610,N_1846);
or U2515 (N_2515,In_4975,In_3555);
xnor U2516 (N_2516,In_1911,In_957);
nand U2517 (N_2517,N_2177,In_4189);
xor U2518 (N_2518,N_34,N_2126);
nand U2519 (N_2519,N_1076,In_428);
or U2520 (N_2520,In_3773,In_2239);
and U2521 (N_2521,In_4328,In_2440);
xor U2522 (N_2522,N_1993,In_1866);
xor U2523 (N_2523,N_1621,N_1407);
xnor U2524 (N_2524,N_104,N_848);
or U2525 (N_2525,In_3765,In_19);
nand U2526 (N_2526,N_1390,N_2189);
and U2527 (N_2527,N_1855,N_2433);
or U2528 (N_2528,N_1838,N_1172);
xnor U2529 (N_2529,N_2065,N_464);
xor U2530 (N_2530,N_2335,In_3649);
nand U2531 (N_2531,N_2305,N_2293);
nor U2532 (N_2532,N_54,In_4440);
nor U2533 (N_2533,In_2489,In_795);
nand U2534 (N_2534,N_511,N_823);
xnor U2535 (N_2535,N_1705,In_2811);
or U2536 (N_2536,N_801,N_2088);
nand U2537 (N_2537,N_1111,N_1489);
nor U2538 (N_2538,N_632,N_1732);
xnor U2539 (N_2539,N_2456,In_2385);
xor U2540 (N_2540,N_1645,N_2493);
or U2541 (N_2541,N_529,N_2480);
or U2542 (N_2542,In_272,In_395);
and U2543 (N_2543,N_2406,In_4304);
and U2544 (N_2544,N_1694,In_1284);
or U2545 (N_2545,N_1595,In_501);
xnor U2546 (N_2546,In_3709,N_2331);
xor U2547 (N_2547,N_1677,In_4575);
nand U2548 (N_2548,N_1160,N_615);
and U2549 (N_2549,N_2294,N_1113);
nand U2550 (N_2550,In_2499,In_2854);
and U2551 (N_2551,N_701,In_996);
or U2552 (N_2552,N_241,In_1440);
or U2553 (N_2553,N_788,N_1926);
nor U2554 (N_2554,In_4526,In_655);
and U2555 (N_2555,N_958,N_1940);
or U2556 (N_2556,N_2124,N_1541);
nor U2557 (N_2557,In_134,N_2322);
nand U2558 (N_2558,N_2439,N_2073);
nor U2559 (N_2559,In_4494,In_3839);
nor U2560 (N_2560,In_2914,In_2733);
nand U2561 (N_2561,N_2400,N_1968);
xor U2562 (N_2562,In_543,In_4382);
and U2563 (N_2563,N_685,In_2895);
nand U2564 (N_2564,N_2499,N_2415);
nor U2565 (N_2565,In_21,N_608);
and U2566 (N_2566,N_1501,In_4042);
nand U2567 (N_2567,N_1788,In_3317);
xor U2568 (N_2568,N_1872,N_2375);
nand U2569 (N_2569,N_2410,In_3358);
nor U2570 (N_2570,In_527,N_2068);
nor U2571 (N_2571,N_749,In_2717);
nand U2572 (N_2572,In_2519,In_451);
nand U2573 (N_2573,In_4266,N_939);
nand U2574 (N_2574,N_2061,N_941);
or U2575 (N_2575,In_2886,In_3764);
nor U2576 (N_2576,In_3658,N_1801);
and U2577 (N_2577,N_767,In_1744);
or U2578 (N_2578,In_2002,In_1381);
or U2579 (N_2579,N_1471,N_2216);
nand U2580 (N_2580,N_1842,N_2053);
or U2581 (N_2581,N_803,N_2184);
nor U2582 (N_2582,N_949,N_1966);
and U2583 (N_2583,N_1975,In_3611);
nand U2584 (N_2584,N_1879,N_2369);
nor U2585 (N_2585,N_1650,N_2143);
nand U2586 (N_2586,In_1919,In_3184);
xor U2587 (N_2587,In_1483,N_1651);
nor U2588 (N_2588,N_1429,In_469);
and U2589 (N_2589,In_1681,In_3014);
nor U2590 (N_2590,In_1458,N_1853);
nand U2591 (N_2591,In_3858,In_886);
nor U2592 (N_2592,N_1892,In_4390);
nand U2593 (N_2593,N_1394,In_3924);
nand U2594 (N_2594,N_2027,In_4159);
xnor U2595 (N_2595,N_723,N_2266);
nor U2596 (N_2596,In_3150,In_514);
xor U2597 (N_2597,N_1232,In_1380);
or U2598 (N_2598,N_1122,In_2264);
nor U2599 (N_2599,N_496,N_1067);
nand U2600 (N_2600,N_2172,In_193);
nand U2601 (N_2601,In_3668,In_528);
and U2602 (N_2602,N_667,N_2078);
nor U2603 (N_2603,In_3136,N_878);
or U2604 (N_2604,N_1608,In_4262);
nand U2605 (N_2605,N_1803,N_2149);
nor U2606 (N_2606,N_696,N_1081);
and U2607 (N_2607,In_2079,N_2116);
and U2608 (N_2608,In_412,N_712);
or U2609 (N_2609,In_4311,N_1585);
xnor U2610 (N_2610,N_14,N_697);
nand U2611 (N_2611,In_2688,In_188);
or U2612 (N_2612,In_3930,N_1398);
and U2613 (N_2613,In_2716,N_1794);
or U2614 (N_2614,N_424,N_2226);
nor U2615 (N_2615,N_1715,N_2133);
or U2616 (N_2616,N_2214,In_1341);
or U2617 (N_2617,N_1482,N_2145);
or U2618 (N_2618,N_1909,N_1265);
and U2619 (N_2619,N_375,N_1491);
nand U2620 (N_2620,In_1787,In_519);
nor U2621 (N_2621,N_1021,N_729);
nand U2622 (N_2622,In_3700,N_1208);
nand U2623 (N_2623,N_2477,N_1203);
or U2624 (N_2624,In_4377,In_1113);
or U2625 (N_2625,N_2045,N_2208);
nor U2626 (N_2626,N_983,N_2316);
or U2627 (N_2627,N_1701,In_4811);
nor U2628 (N_2628,In_4766,N_992);
and U2629 (N_2629,N_2302,N_1752);
or U2630 (N_2630,In_162,In_3291);
xnor U2631 (N_2631,In_948,N_1088);
nor U2632 (N_2632,N_1381,In_1845);
and U2633 (N_2633,N_2330,In_4934);
and U2634 (N_2634,In_3679,In_2804);
xnor U2635 (N_2635,N_1299,N_2037);
nor U2636 (N_2636,In_1539,N_204);
nand U2637 (N_2637,N_2368,In_1855);
nand U2638 (N_2638,In_2579,N_1775);
xnor U2639 (N_2639,N_1061,N_2039);
nand U2640 (N_2640,N_2253,N_2026);
nand U2641 (N_2641,In_2648,N_2082);
or U2642 (N_2642,In_2038,In_4984);
nor U2643 (N_2643,In_1630,In_1534);
nand U2644 (N_2644,In_2022,N_1293);
nor U2645 (N_2645,N_681,In_3275);
or U2646 (N_2646,In_2955,N_119);
and U2647 (N_2647,N_2141,In_3582);
xor U2648 (N_2648,N_2256,N_2171);
xnor U2649 (N_2649,In_3245,In_3866);
and U2650 (N_2650,In_3344,N_2270);
xnor U2651 (N_2651,N_1105,N_2281);
nor U2652 (N_2652,In_2966,N_2234);
and U2653 (N_2653,N_2144,In_3479);
or U2654 (N_2654,N_2176,N_2190);
and U2655 (N_2655,N_2212,In_3257);
xor U2656 (N_2656,In_4976,N_954);
xnor U2657 (N_2657,In_2422,N_2121);
nand U2658 (N_2658,In_1429,In_2369);
and U2659 (N_2659,N_541,In_3402);
and U2660 (N_2660,N_1182,N_2066);
xor U2661 (N_2661,In_1468,In_788);
and U2662 (N_2662,In_317,N_2217);
or U2663 (N_2663,In_2320,In_1790);
nand U2664 (N_2664,N_1449,N_2285);
nand U2665 (N_2665,N_1463,In_4928);
nor U2666 (N_2666,In_4680,In_3797);
xnor U2667 (N_2667,In_2845,In_1233);
or U2668 (N_2668,In_4883,In_190);
or U2669 (N_2669,In_949,In_3497);
nand U2670 (N_2670,In_75,In_4677);
or U2671 (N_2671,N_1063,In_2736);
and U2672 (N_2672,In_3121,In_1983);
nor U2673 (N_2673,N_1887,N_899);
and U2674 (N_2674,N_2057,N_2060);
or U2675 (N_2675,In_4044,N_682);
nand U2676 (N_2676,In_722,N_1565);
or U2677 (N_2677,N_1478,In_574);
nor U2678 (N_2678,N_23,N_2008);
nand U2679 (N_2679,N_1441,In_1970);
and U2680 (N_2680,In_192,N_623);
nor U2681 (N_2681,N_2470,N_1664);
or U2682 (N_2682,N_602,In_2157);
or U2683 (N_2683,N_2489,N_1593);
or U2684 (N_2684,N_1648,N_2003);
nand U2685 (N_2685,In_3608,N_1750);
nor U2686 (N_2686,N_1655,N_1884);
or U2687 (N_2687,N_2150,N_565);
and U2688 (N_2688,In_3069,In_1365);
nor U2689 (N_2689,In_478,In_1333);
and U2690 (N_2690,In_4587,N_2185);
nand U2691 (N_2691,In_3073,N_1207);
nor U2692 (N_2692,N_2136,N_2367);
or U2693 (N_2693,N_669,In_1102);
and U2694 (N_2694,N_209,N_1512);
and U2695 (N_2695,In_1394,In_3278);
or U2696 (N_2696,N_1231,In_541);
nand U2697 (N_2697,In_1577,In_1962);
nand U2698 (N_2698,N_1929,N_2249);
or U2699 (N_2699,In_685,In_677);
xor U2700 (N_2700,In_4568,In_1691);
nor U2701 (N_2701,In_4477,In_4003);
or U2702 (N_2702,In_293,N_1408);
nand U2703 (N_2703,N_1827,N_2040);
xor U2704 (N_2704,N_532,N_2430);
xnor U2705 (N_2705,N_1440,N_710);
or U2706 (N_2706,N_1187,N_2411);
or U2707 (N_2707,In_102,N_1776);
or U2708 (N_2708,N_2206,In_2288);
nor U2709 (N_2709,In_4402,N_1710);
or U2710 (N_2710,N_1228,In_4600);
nand U2711 (N_2711,N_2173,N_66);
or U2712 (N_2712,In_3490,N_2312);
or U2713 (N_2713,N_1729,In_1446);
and U2714 (N_2714,N_2224,N_853);
nor U2715 (N_2715,In_2151,N_2319);
nand U2716 (N_2716,In_4314,N_2409);
nor U2717 (N_2717,N_1996,N_2052);
or U2718 (N_2718,N_2260,N_2055);
nand U2719 (N_2719,N_1992,N_1882);
nor U2720 (N_2720,In_1470,In_2713);
nor U2721 (N_2721,N_201,N_252);
and U2722 (N_2722,In_4567,N_2444);
xnor U2723 (N_2723,In_4825,N_421);
nand U2724 (N_2724,N_2106,In_4594);
nand U2725 (N_2725,N_1988,In_4875);
nand U2726 (N_2726,In_229,N_1186);
xnor U2727 (N_2727,N_910,In_2584);
and U2728 (N_2728,In_970,In_2776);
xor U2729 (N_2729,In_632,In_913);
nor U2730 (N_2730,N_117,N_1634);
nor U2731 (N_2731,In_1795,N_2381);
nor U2732 (N_2732,N_8,N_1132);
or U2733 (N_2733,In_2678,N_2455);
nand U2734 (N_2734,In_4312,N_1245);
xnor U2735 (N_2735,N_2397,N_859);
xnor U2736 (N_2736,In_1686,N_2424);
xor U2737 (N_2737,In_4142,In_3481);
xor U2738 (N_2738,N_1865,N_1885);
nand U2739 (N_2739,In_4191,In_4487);
xor U2740 (N_2740,N_2278,N_2084);
nand U2741 (N_2741,N_457,N_2228);
xor U2742 (N_2742,N_1275,In_564);
or U2743 (N_2743,In_1036,N_2183);
xnor U2744 (N_2744,N_1468,In_424);
nor U2745 (N_2745,In_410,In_3293);
and U2746 (N_2746,In_104,N_661);
and U2747 (N_2747,N_1564,In_674);
nand U2748 (N_2748,N_1376,N_1936);
nor U2749 (N_2749,In_1375,N_2342);
and U2750 (N_2750,N_195,N_916);
nor U2751 (N_2751,In_4499,In_496);
and U2752 (N_2752,In_3157,In_2646);
nor U2753 (N_2753,N_2488,N_1730);
and U2754 (N_2754,In_2807,N_772);
xor U2755 (N_2755,In_283,In_4692);
nor U2756 (N_2756,N_1517,N_226);
or U2757 (N_2757,In_3251,In_391);
nor U2758 (N_2758,N_341,In_607);
xor U2759 (N_2759,In_2155,N_2394);
nor U2760 (N_2760,N_2021,N_2401);
xor U2761 (N_2761,In_1944,N_1238);
and U2762 (N_2762,N_694,N_2324);
nand U2763 (N_2763,N_1335,N_1377);
and U2764 (N_2764,N_1653,N_1937);
nand U2765 (N_2765,N_2459,In_1961);
and U2766 (N_2766,In_538,N_161);
nor U2767 (N_2767,N_2491,In_4588);
xnor U2768 (N_2768,In_4607,In_1704);
or U2769 (N_2769,In_2620,In_4016);
nor U2770 (N_2770,In_4948,N_271);
nor U2771 (N_2771,N_1327,N_2180);
or U2772 (N_2772,In_4031,N_557);
or U2773 (N_2773,N_1288,N_505);
and U2774 (N_2774,N_295,In_3955);
or U2775 (N_2775,N_2123,N_2336);
and U2776 (N_2776,In_2510,In_4608);
or U2777 (N_2777,In_4993,In_4871);
or U2778 (N_2778,In_3778,In_4730);
nor U2779 (N_2779,N_71,N_862);
nor U2780 (N_2780,In_3023,N_1835);
xnor U2781 (N_2781,N_1942,In_1455);
nor U2782 (N_2782,In_912,N_2469);
or U2783 (N_2783,N_2317,In_573);
and U2784 (N_2784,N_642,N_2359);
nor U2785 (N_2785,N_191,In_3602);
nand U2786 (N_2786,N_1522,N_1434);
nor U2787 (N_2787,In_4738,In_3173);
and U2788 (N_2788,N_1939,In_4520);
xnor U2789 (N_2789,N_1844,In_4783);
nand U2790 (N_2790,N_106,N_2135);
nor U2791 (N_2791,In_1445,In_1071);
nand U2792 (N_2792,In_812,In_509);
nand U2793 (N_2793,N_1934,In_3715);
xnor U2794 (N_2794,In_4558,N_1300);
xnor U2795 (N_2795,In_2575,N_2452);
nand U2796 (N_2796,N_1248,N_1830);
and U2797 (N_2797,N_5,In_2557);
nand U2798 (N_2798,In_3070,In_3710);
or U2799 (N_2799,In_2610,N_2209);
nand U2800 (N_2800,N_1069,In_1585);
nand U2801 (N_2801,N_2428,In_1898);
and U2802 (N_2802,N_1906,N_869);
nand U2803 (N_2803,In_127,In_2934);
or U2804 (N_2804,N_2178,In_3308);
and U2805 (N_2805,In_4620,In_2031);
xnor U2806 (N_2806,In_3248,N_2479);
nor U2807 (N_2807,In_802,N_2181);
and U2808 (N_2808,In_1593,In_2502);
nand U2809 (N_2809,In_4455,N_113);
or U2810 (N_2810,In_3234,In_440);
nand U2811 (N_2811,In_4690,In_1636);
and U2812 (N_2812,In_4364,N_2403);
xor U2813 (N_2813,In_3258,N_1281);
nor U2814 (N_2814,N_213,N_2320);
or U2815 (N_2815,N_2283,In_2247);
and U2816 (N_2816,N_884,In_224);
or U2817 (N_2817,N_1154,N_2240);
or U2818 (N_2818,In_2527,In_2097);
or U2819 (N_2819,In_861,In_447);
and U2820 (N_2820,In_621,In_2848);
and U2821 (N_2821,N_721,In_289);
xor U2822 (N_2822,N_97,In_3794);
and U2823 (N_2823,In_2204,N_253);
or U2824 (N_2824,In_4978,In_2743);
nor U2825 (N_2825,N_2227,N_2207);
xor U2826 (N_2826,In_1515,N_1912);
xnor U2827 (N_2827,N_2458,N_1590);
and U2828 (N_2828,In_3595,In_3845);
nor U2829 (N_2829,In_3735,N_432);
nand U2830 (N_2830,In_3290,In_4062);
nand U2831 (N_2831,In_3751,In_4027);
xnor U2832 (N_2832,N_1703,N_824);
xnor U2833 (N_2833,N_1323,N_2352);
and U2834 (N_2834,N_1375,In_3076);
and U2835 (N_2835,In_2201,N_422);
and U2836 (N_2836,In_2163,In_2343);
nand U2837 (N_2837,N_821,In_1807);
and U2838 (N_2838,In_4566,N_2000);
nor U2839 (N_2839,N_2273,N_1734);
and U2840 (N_2840,N_2257,N_1610);
nand U2841 (N_2841,In_4765,In_3170);
and U2842 (N_2842,N_2417,In_3326);
nor U2843 (N_2843,N_1946,N_1639);
nand U2844 (N_2844,In_1313,N_2169);
and U2845 (N_2845,In_2779,N_607);
and U2846 (N_2846,N_562,N_826);
nand U2847 (N_2847,In_3341,In_2325);
or U2848 (N_2848,In_62,N_2453);
xor U2849 (N_2849,N_2310,In_2562);
nor U2850 (N_2850,N_962,N_1854);
nand U2851 (N_2851,N_313,N_243);
nor U2852 (N_2852,In_57,N_2402);
or U2853 (N_2853,In_2295,In_2434);
xnor U2854 (N_2854,In_3564,In_4855);
xnor U2855 (N_2855,In_1207,In_2604);
nand U2856 (N_2856,N_1742,N_2481);
nand U2857 (N_2857,N_348,N_450);
and U2858 (N_2858,N_1005,In_4392);
and U2859 (N_2859,In_113,N_369);
and U2860 (N_2860,In_3631,N_308);
nand U2861 (N_2861,N_1699,In_3616);
nand U2862 (N_2862,In_2101,N_1328);
xor U2863 (N_2863,N_2490,In_3379);
nor U2864 (N_2864,N_990,N_2168);
nand U2865 (N_2865,In_1770,In_3739);
nor U2866 (N_2866,In_1144,N_2354);
nor U2867 (N_2867,In_2136,N_1130);
or U2868 (N_2868,N_2005,N_1104);
and U2869 (N_2869,In_4448,In_1357);
and U2870 (N_2870,In_4688,In_2946);
xnor U2871 (N_2871,In_4432,N_812);
xor U2872 (N_2872,In_1728,In_1586);
nand U2873 (N_2873,In_64,In_2629);
xnor U2874 (N_2874,N_1613,In_2525);
and U2875 (N_2875,N_621,N_2496);
or U2876 (N_2876,In_3571,N_1704);
xnor U2877 (N_2877,N_2419,N_487);
nand U2878 (N_2878,N_1316,In_2991);
and U2879 (N_2879,In_3517,N_2364);
xnor U2880 (N_2880,N_2395,N_1557);
xor U2881 (N_2881,N_231,N_2081);
xor U2882 (N_2882,In_2180,N_1708);
xor U2883 (N_2883,N_585,N_29);
xor U2884 (N_2884,N_1164,N_806);
or U2885 (N_2885,In_4632,In_3364);
or U2886 (N_2886,N_1869,N_1542);
nor U2887 (N_2887,N_2159,In_4450);
nand U2888 (N_2888,In_2751,In_2358);
nor U2889 (N_2889,In_4756,N_1622);
and U2890 (N_2890,In_1972,N_2011);
and U2891 (N_2891,In_2503,N_1714);
xor U2892 (N_2892,N_2473,In_4192);
and U2893 (N_2893,In_2323,In_2754);
nand U2894 (N_2894,N_1142,N_1382);
and U2895 (N_2895,N_1592,In_3964);
or U2896 (N_2896,N_2271,N_1215);
nand U2897 (N_2897,In_337,N_1548);
nand U2898 (N_2898,N_1404,N_13);
xnor U2899 (N_2899,N_610,In_2217);
nor U2900 (N_2900,N_1551,N_203);
nor U2901 (N_2901,N_312,In_1000);
and U2902 (N_2902,N_413,In_3523);
nand U2903 (N_2903,N_2229,In_2198);
nor U2904 (N_2904,In_1736,N_1709);
nand U2905 (N_2905,N_1889,In_3459);
nor U2906 (N_2906,N_1252,N_274);
nand U2907 (N_2907,N_515,N_1812);
nand U2908 (N_2908,N_2476,In_3310);
nor U2909 (N_2909,N_1620,In_679);
nand U2910 (N_2910,In_3982,In_3063);
xor U2911 (N_2911,In_2967,N_1857);
nand U2912 (N_2912,N_2357,N_995);
nor U2913 (N_2913,In_1904,N_2391);
or U2914 (N_2914,N_2265,N_2163);
nand U2915 (N_2915,N_350,N_808);
nor U2916 (N_2916,In_4351,N_2353);
or U2917 (N_2917,N_2118,N_1543);
or U2918 (N_2918,N_1135,N_1475);
nor U2919 (N_2919,N_254,In_3623);
nand U2920 (N_2920,N_839,N_2376);
nor U2921 (N_2921,In_1204,In_222);
and U2922 (N_2922,N_2105,In_4020);
nor U2923 (N_2923,In_4636,In_146);
and U2924 (N_2924,In_3264,N_1643);
and U2925 (N_2925,N_1904,In_52);
nand U2926 (N_2926,In_1878,N_1144);
xor U2927 (N_2927,In_3499,In_1656);
nor U2928 (N_2928,In_2452,In_2408);
nor U2929 (N_2929,In_643,In_2892);
nand U2930 (N_2930,N_581,N_1718);
nor U2931 (N_2931,N_1556,In_785);
nor U2932 (N_2932,N_1712,N_2162);
nor U2933 (N_2933,N_315,N_1374);
xnor U2934 (N_2934,N_1994,In_4982);
and U2935 (N_2935,In_709,N_660);
xor U2936 (N_2936,N_1725,In_535);
or U2937 (N_2937,In_1250,In_88);
or U2938 (N_2938,In_314,N_957);
and U2939 (N_2939,In_1764,N_2497);
xor U2940 (N_2940,N_558,N_2160);
or U2941 (N_2941,N_2007,In_2998);
nand U2942 (N_2942,N_768,In_1171);
nand U2943 (N_2943,In_1509,N_2321);
xor U2944 (N_2944,N_1769,In_2102);
nor U2945 (N_2945,N_2076,N_2102);
nor U2946 (N_2946,In_3972,N_2225);
nor U2947 (N_2947,N_2464,N_427);
and U2948 (N_2948,In_36,N_2363);
or U2949 (N_2949,N_2018,In_2652);
nand U2950 (N_2950,In_4337,N_1450);
nor U2951 (N_2951,N_2498,N_657);
and U2952 (N_2952,N_1264,N_507);
xor U2953 (N_2953,N_1901,In_2852);
or U2954 (N_2954,N_1271,In_2516);
nor U2955 (N_2955,In_30,N_393);
nor U2956 (N_2956,N_2298,In_2761);
nand U2957 (N_2957,In_613,N_394);
xnor U2958 (N_2958,N_1110,N_1439);
xor U2959 (N_2959,N_1502,N_2386);
nand U2960 (N_2960,N_2091,N_1588);
nand U2961 (N_2961,In_1640,N_2431);
and U2962 (N_2962,In_2212,In_4800);
xnor U2963 (N_2963,N_443,N_2250);
nand U2964 (N_2964,In_4617,In_4109);
and U2965 (N_2965,N_2445,N_194);
nor U2966 (N_2966,In_2595,In_561);
nor U2967 (N_2967,In_1485,In_2540);
xnor U2968 (N_2968,N_64,N_1707);
and U2969 (N_2969,N_1602,N_86);
and U2970 (N_2970,N_2243,In_435);
nor U2971 (N_2971,In_680,N_1516);
nor U2972 (N_2972,In_1077,In_416);
or U2973 (N_2973,N_2156,In_4367);
and U2974 (N_2974,In_927,In_1518);
and U2975 (N_2975,N_1043,N_336);
or U2976 (N_2976,N_90,N_570);
nor U2977 (N_2977,In_1359,N_1826);
xor U2978 (N_2978,N_2194,N_1116);
nor U2979 (N_2979,In_1828,N_2117);
nand U2980 (N_2980,In_2266,N_2289);
or U2981 (N_2981,N_1392,In_707);
or U2982 (N_2982,N_2245,N_1194);
or U2983 (N_2983,N_1849,In_1221);
nor U2984 (N_2984,N_1127,N_1220);
nand U2985 (N_2985,N_181,N_199);
and U2986 (N_2986,N_792,N_2384);
or U2987 (N_2987,In_1956,N_1589);
or U2988 (N_2988,In_4224,In_374);
and U2989 (N_2989,N_1520,In_2523);
xnor U2990 (N_2990,In_4792,N_1574);
xnor U2991 (N_2991,N_438,In_557);
nand U2992 (N_2992,N_2344,N_1956);
xnor U2993 (N_2993,N_2340,N_2108);
and U2994 (N_2994,N_688,N_2179);
and U2995 (N_2995,N_409,N_2019);
and U2996 (N_2996,In_2518,N_2235);
nand U2997 (N_2997,N_923,In_1180);
nor U2998 (N_2998,In_4938,In_2745);
or U2999 (N_2999,N_2094,In_1635);
xnor U3000 (N_3000,In_3915,N_2507);
or U3001 (N_3001,In_3388,In_577);
and U3002 (N_3002,N_2529,N_2770);
or U3003 (N_3003,In_2128,In_4479);
or U3004 (N_3004,N_1692,In_4788);
nand U3005 (N_3005,N_2592,In_4578);
nand U3006 (N_3006,In_393,N_2855);
and U3007 (N_3007,In_2081,In_3607);
and U3008 (N_3008,N_603,N_402);
nor U3009 (N_3009,N_2709,N_1379);
xnor U3010 (N_3010,In_1550,N_1361);
nor U3011 (N_3011,N_2380,N_1279);
nand U3012 (N_3012,N_2775,N_2727);
xnor U3013 (N_3013,N_2441,N_2943);
nor U3014 (N_3014,N_368,N_2296);
and U3015 (N_3015,N_257,N_921);
xnor U3016 (N_3016,N_493,N_3);
and U3017 (N_3017,N_1078,In_1299);
nand U3018 (N_3018,N_2815,N_1465);
nand U3019 (N_3019,In_4025,N_2902);
xor U3020 (N_3020,In_3849,N_2790);
or U3021 (N_3021,N_2789,In_923);
nand U3022 (N_3022,In_4324,N_2511);
xnor U3023 (N_3023,N_1786,N_365);
nor U3024 (N_3024,N_2203,In_3519);
nor U3025 (N_3025,N_2286,In_665);
and U3026 (N_3026,In_1025,N_1147);
nor U3027 (N_3027,N_2760,N_1467);
nor U3028 (N_3028,In_3622,N_154);
and U3029 (N_3029,N_1528,N_2443);
nor U3030 (N_3030,In_2029,N_508);
nand U3031 (N_3031,N_2939,N_2128);
and U3032 (N_3032,In_3355,In_2209);
and U3033 (N_3033,N_1137,N_2640);
nand U3034 (N_3034,N_2593,N_2350);
or U3035 (N_3035,N_2609,N_2515);
and U3036 (N_3036,N_2110,N_2619);
and U3037 (N_3037,N_2842,N_1233);
nor U3038 (N_3038,N_2523,N_2337);
or U3039 (N_3039,N_2304,N_1510);
and U3040 (N_3040,N_2528,In_4167);
nor U3041 (N_3041,N_1552,N_1720);
xor U3042 (N_3042,N_1876,In_2056);
nor U3043 (N_3043,N_2941,In_2687);
nor U3044 (N_3044,N_2835,In_1368);
and U3045 (N_3045,N_1791,In_843);
or U3046 (N_3046,N_2744,N_2556);
or U3047 (N_3047,In_3217,N_2997);
and U3048 (N_3048,In_1894,N_2862);
nor U3049 (N_3049,N_2877,In_771);
nor U3050 (N_3050,N_2538,N_361);
or U3051 (N_3051,N_2001,N_2536);
nor U3052 (N_3052,N_2699,N_775);
nand U3053 (N_3053,In_4258,N_2998);
nor U3054 (N_3054,N_2090,In_1921);
nor U3055 (N_3055,N_2086,In_4104);
or U3056 (N_3056,In_1797,N_1977);
or U3057 (N_3057,N_2526,N_2072);
nor U3058 (N_3058,N_2780,In_4654);
nor U3059 (N_3059,N_1500,N_2089);
nor U3060 (N_3060,In_1175,N_1870);
or U3061 (N_3061,In_2771,N_2891);
nand U3062 (N_3062,In_1105,N_1963);
xor U3063 (N_3063,N_2962,N_699);
or U3064 (N_3064,N_1544,N_2944);
xor U3065 (N_3065,N_1806,In_245);
or U3066 (N_3066,N_1821,In_2806);
nand U3067 (N_3067,In_3609,In_2552);
nand U3068 (N_3068,N_2355,N_2233);
or U3069 (N_3069,N_1008,N_780);
or U3070 (N_3070,In_4775,N_2648);
and U3071 (N_3071,N_2134,N_2697);
or U3072 (N_3072,N_2462,N_2516);
nor U3073 (N_3073,N_2127,N_2740);
nand U3074 (N_3074,N_1333,In_303);
and U3075 (N_3075,N_2890,N_1430);
nor U3076 (N_3076,N_1983,In_1024);
and U3077 (N_3077,In_228,In_380);
xor U3078 (N_3078,N_2732,In_1004);
or U3079 (N_3079,N_1257,N_1026);
xnor U3080 (N_3080,N_73,N_1638);
xnor U3081 (N_3081,N_2010,In_4293);
and U3082 (N_3082,In_4952,N_2696);
nand U3083 (N_3083,N_713,In_2112);
nand U3084 (N_3084,N_2042,In_83);
nor U3085 (N_3085,N_2119,In_1876);
or U3086 (N_3086,N_1998,N_2611);
or U3087 (N_3087,In_399,N_2280);
xor U3088 (N_3088,In_1104,N_1223);
or U3089 (N_3089,N_857,N_964);
xor U3090 (N_3090,N_2158,N_2936);
nand U3091 (N_3091,In_1001,In_4153);
nand U3092 (N_3092,In_4035,In_740);
nand U3093 (N_3093,N_215,N_2182);
nand U3094 (N_3094,In_4373,In_1710);
nand U3095 (N_3095,N_714,In_2091);
xnor U3096 (N_3096,N_2687,In_1954);
or U3097 (N_3097,N_2765,N_820);
and U3098 (N_3098,In_3917,N_1072);
nor U3099 (N_3099,N_2773,N_2070);
nand U3100 (N_3100,N_1781,N_2518);
xor U3101 (N_3101,In_4716,In_792);
or U3102 (N_3102,N_1474,N_2098);
and U3103 (N_3103,N_2432,N_2492);
or U3104 (N_3104,N_305,N_1802);
nor U3105 (N_3105,In_298,N_2661);
or U3106 (N_3106,N_1139,N_2259);
nor U3107 (N_3107,N_1695,N_959);
or U3108 (N_3108,N_1460,N_2851);
xor U3109 (N_3109,N_698,In_1796);
and U3110 (N_3110,N_2097,N_2041);
xor U3111 (N_3111,N_2202,N_2993);
nor U3112 (N_3112,N_1796,N_2313);
or U3113 (N_3113,N_2530,In_3664);
nand U3114 (N_3114,N_1987,N_2724);
nor U3115 (N_3115,In_261,N_2418);
and U3116 (N_3116,In_2524,N_2122);
nand U3117 (N_3117,N_2734,N_2562);
and U3118 (N_3118,In_2793,In_3135);
xnor U3119 (N_3119,N_1778,In_2613);
nand U3120 (N_3120,In_1444,N_2781);
nor U3121 (N_3121,N_1702,N_2650);
xor U3122 (N_3122,In_4664,In_801);
nor U3123 (N_3123,N_1312,In_2537);
and U3124 (N_3124,In_2844,N_831);
or U3125 (N_3125,N_2218,N_2554);
xor U3126 (N_3126,N_852,N_1546);
nor U3127 (N_3127,N_2980,In_2284);
xor U3128 (N_3128,N_2950,N_2920);
xnor U3129 (N_3129,In_2007,N_2940);
xnor U3130 (N_3130,N_491,N_2139);
xnor U3131 (N_3131,N_2351,In_1087);
and U3132 (N_3132,In_130,In_757);
and U3133 (N_3133,N_2617,N_2038);
nor U3134 (N_3134,N_1167,In_1900);
and U3135 (N_3135,In_3434,N_1832);
xnor U3136 (N_3136,In_1402,N_2864);
nand U3137 (N_3137,N_2193,N_2146);
xnor U3138 (N_3138,In_2814,N_2755);
and U3139 (N_3139,In_2554,N_2804);
or U3140 (N_3140,N_668,N_1262);
nand U3141 (N_3141,N_1339,In_580);
nor U3142 (N_3142,In_4695,In_1752);
nand U3143 (N_3143,N_732,In_2162);
xor U3144 (N_3144,In_259,N_490);
and U3145 (N_3145,N_2654,In_772);
xor U3146 (N_3146,In_4255,In_2671);
nor U3147 (N_3147,In_1344,N_2385);
nand U3148 (N_3148,N_2546,N_2754);
nor U3149 (N_3149,N_2738,In_4944);
nor U3150 (N_3150,N_1626,N_2646);
nor U3151 (N_3151,N_2628,N_2390);
nor U3152 (N_3152,N_876,In_3262);
nor U3153 (N_3153,In_459,N_2627);
or U3154 (N_3154,N_2783,N_2131);
xor U3155 (N_3155,N_2875,N_2818);
nand U3156 (N_3156,N_2147,N_522);
nand U3157 (N_3157,N_2111,In_1490);
and U3158 (N_3158,In_2578,In_2931);
xnor U3159 (N_3159,N_1978,N_2140);
or U3160 (N_3160,N_2288,N_1675);
xnor U3161 (N_3161,N_2502,N_2942);
and U3162 (N_3162,N_2692,In_1608);
and U3163 (N_3163,N_2210,N_563);
or U3164 (N_3164,In_4579,N_1121);
nand U3165 (N_3165,N_2618,N_1676);
and U3166 (N_3166,N_2840,N_2196);
nand U3167 (N_3167,In_1319,N_2635);
and U3168 (N_3168,In_4551,N_2797);
or U3169 (N_3169,In_2786,In_9);
and U3170 (N_3170,N_2984,N_1809);
nand U3171 (N_3171,In_1566,In_3243);
nor U3172 (N_3172,N_2239,N_1969);
nand U3173 (N_3173,In_4117,N_236);
and U3174 (N_3174,In_2691,N_750);
nor U3175 (N_3175,N_867,In_384);
nand U3176 (N_3176,N_2398,In_2824);
or U3177 (N_3177,N_2085,N_2374);
nand U3178 (N_3178,N_1671,N_2413);
and U3179 (N_3179,In_4435,N_2537);
xor U3180 (N_3180,N_930,N_2487);
xor U3181 (N_3181,N_437,N_1591);
nor U3182 (N_3182,In_4967,N_366);
nor U3183 (N_3183,N_1345,N_1880);
xor U3184 (N_3184,N_2805,In_1914);
nand U3185 (N_3185,N_2129,N_1897);
and U3186 (N_3186,N_1258,N_1023);
nor U3187 (N_3187,N_545,N_2888);
nor U3188 (N_3188,N_1230,N_2563);
xor U3189 (N_3189,N_1093,N_1582);
nor U3190 (N_3190,In_1760,N_1537);
nand U3191 (N_3191,In_4963,In_3380);
xnor U3192 (N_3192,N_392,N_2557);
and U3193 (N_3193,In_911,N_1386);
and U3194 (N_3194,N_2884,In_1413);
or U3195 (N_3195,In_758,In_2539);
nand U3196 (N_3196,N_2577,N_1672);
nand U3197 (N_3197,In_2221,N_75);
nor U3198 (N_3198,N_1481,N_2971);
and U3199 (N_3199,N_1636,N_2358);
or U3200 (N_3200,N_1560,N_2894);
nand U3201 (N_3201,N_290,N_2230);
and U3202 (N_3202,N_2155,N_1570);
and U3203 (N_3203,In_3792,In_4703);
and U3204 (N_3204,N_2307,In_1582);
or U3205 (N_3205,N_2356,N_1325);
or U3206 (N_3206,N_2615,N_2876);
and U3207 (N_3207,N_1900,N_2112);
or U3208 (N_3208,N_1578,N_929);
nor U3209 (N_3209,N_1524,In_816);
nor U3210 (N_3210,N_2975,In_2487);
or U3211 (N_3211,N_578,N_2747);
nand U3212 (N_3212,N_2077,In_3737);
nor U3213 (N_3213,In_3880,In_3961);
and U3214 (N_3214,N_2689,In_470);
nor U3215 (N_3215,N_2248,N_2796);
or U3216 (N_3216,N_2130,N_2982);
and U3217 (N_3217,N_2581,In_2301);
nand U3218 (N_3218,In_94,N_2625);
and U3219 (N_3219,N_2623,N_882);
and U3220 (N_3220,In_3176,N_2263);
xnor U3221 (N_3221,N_1014,In_3038);
xor U3222 (N_3222,N_2631,In_4070);
and U3223 (N_3223,In_1312,N_2680);
or U3224 (N_3224,N_2585,N_2904);
or U3225 (N_3225,N_2028,In_4267);
nor U3226 (N_3226,N_739,In_689);
nand U3227 (N_3227,N_2669,In_2548);
or U3228 (N_3228,N_415,N_2752);
or U3229 (N_3229,N_2691,N_1757);
or U3230 (N_3230,In_1750,In_1467);
nand U3231 (N_3231,In_2095,N_1743);
or U3232 (N_3232,N_2211,In_79);
nor U3233 (N_3233,In_3433,In_4625);
nand U3234 (N_3234,In_815,N_2421);
and U3235 (N_3235,N_109,N_651);
nor U3236 (N_3236,N_1095,N_1862);
nor U3237 (N_3237,N_1679,N_2315);
xnor U3238 (N_3238,In_2310,N_2768);
xnor U3239 (N_3239,N_2004,N_2996);
or U3240 (N_3240,In_4694,In_4752);
and U3241 (N_3241,N_2478,N_2838);
or U3242 (N_3242,N_2705,N_2301);
nand U3243 (N_3243,N_1970,N_1329);
xnor U3244 (N_3244,In_640,N_2025);
or U3245 (N_3245,In_4848,N_2764);
and U3246 (N_3246,N_2987,N_2774);
and U3247 (N_3247,N_2914,N_2449);
nor U3248 (N_3248,In_2134,N_2567);
and U3249 (N_3249,N_2079,N_1576);
or U3250 (N_3250,In_2329,N_994);
nor U3251 (N_3251,In_1018,N_2013);
nor U3252 (N_3252,In_4619,N_2870);
nand U3253 (N_3253,N_2104,N_2454);
and U3254 (N_3254,In_4506,N_1321);
or U3255 (N_3255,N_2372,In_1059);
or U3256 (N_3256,In_2859,In_1154);
nor U3257 (N_3257,N_2595,In_4231);
and U3258 (N_3258,N_2924,N_2779);
or U3259 (N_3259,N_896,In_1119);
xor U3260 (N_3260,N_1037,N_1062);
nand U3261 (N_3261,N_2938,N_2960);
or U3262 (N_3262,N_2204,In_1148);
xnor U3263 (N_3263,In_4601,N_2148);
or U3264 (N_3264,N_913,In_2147);
and U3265 (N_3265,In_2520,N_1017);
or U3266 (N_3266,N_2300,In_4252);
or U3267 (N_3267,N_2659,N_2915);
and U3268 (N_3268,N_1027,In_2168);
nor U3269 (N_3269,N_2677,N_2165);
and U3270 (N_3270,In_3223,In_4599);
nor U3271 (N_3271,In_2897,N_2437);
nand U3272 (N_3272,N_2152,N_2685);
nor U3273 (N_3273,N_2571,N_1266);
nand U3274 (N_3274,N_544,In_3770);
xnor U3275 (N_3275,N_2872,N_2534);
xnor U3276 (N_3276,In_1281,N_2334);
and U3277 (N_3277,N_1759,In_125);
nor U3278 (N_3278,N_2954,N_1571);
nand U3279 (N_3279,N_2101,N_2032);
and U3280 (N_3280,In_2864,In_1463);
or U3281 (N_3281,In_1926,In_2127);
and U3282 (N_3282,N_2782,N_2868);
and U3283 (N_3283,N_1813,N_1635);
and U3284 (N_3284,N_2632,In_4420);
nand U3285 (N_3285,N_2535,In_4631);
xnor U3286 (N_3286,In_220,N_1690);
nor U3287 (N_3287,N_2978,In_103);
nor U3288 (N_3288,N_2525,In_2835);
and U3289 (N_3289,In_4085,In_2268);
nor U3290 (N_3290,N_1728,N_2881);
nor U3291 (N_3291,In_4176,N_2909);
xnor U3292 (N_3292,N_2174,N_1598);
and U3293 (N_3293,N_1181,In_161);
and U3294 (N_3294,N_2096,In_3578);
and U3295 (N_3295,In_3807,In_879);
or U3296 (N_3296,In_676,In_1238);
xor U3297 (N_3297,In_2082,N_2231);
and U3298 (N_3298,In_3539,In_4462);
nand U3299 (N_3299,N_1209,N_1064);
and U3300 (N_3300,N_1783,N_2853);
or U3301 (N_3301,N_1961,N_2125);
xor U3302 (N_3302,N_2800,N_2036);
and U3303 (N_3303,In_2131,N_2850);
nand U3304 (N_3304,N_2652,In_474);
nor U3305 (N_3305,N_1722,N_87);
nand U3306 (N_3306,N_1930,N_835);
or U3307 (N_3307,N_2532,In_2809);
nand U3308 (N_3308,In_3120,In_4728);
nor U3309 (N_3309,N_2629,In_2632);
nor U3310 (N_3310,N_1051,N_1314);
nand U3311 (N_3311,N_1834,In_1652);
nor U3312 (N_3312,N_2861,In_2109);
nor U3313 (N_3313,N_1318,In_3752);
xor U3314 (N_3314,N_2063,N_2863);
nand U3315 (N_3315,N_2603,In_974);
nor U3316 (N_3316,N_2034,N_2509);
and U3317 (N_3317,N_1609,N_1894);
or U3318 (N_3318,In_2402,N_2605);
and U3319 (N_3319,N_2521,In_1349);
or U3320 (N_3320,N_2860,N_2869);
and U3321 (N_3321,In_214,N_2252);
or U3322 (N_3322,In_4638,N_2533);
nand U3323 (N_3323,N_2670,N_2604);
and U3324 (N_3324,N_261,In_2410);
and U3325 (N_3325,N_2587,N_2291);
xnor U3326 (N_3326,N_2396,N_2761);
nand U3327 (N_3327,In_3369,In_4473);
xor U3328 (N_3328,N_1000,N_2934);
xor U3329 (N_3329,N_1096,In_681);
xor U3330 (N_3330,N_2120,In_4093);
xnor U3331 (N_3331,N_2241,N_2720);
nand U3332 (N_3332,N_695,N_88);
and U3333 (N_3333,N_2429,N_2539);
and U3334 (N_3334,N_1297,N_2959);
nor U3335 (N_3335,N_2423,In_4409);
nor U3336 (N_3336,In_4802,N_2594);
and U3337 (N_3337,N_2326,In_3920);
xor U3338 (N_3338,In_1730,N_1380);
xor U3339 (N_3339,N_1668,N_2048);
nand U3340 (N_3340,N_756,N_1654);
nor U3341 (N_3341,N_2472,N_2834);
or U3342 (N_3342,In_2492,N_1235);
nor U3343 (N_3343,N_2484,N_2757);
nand U3344 (N_3344,In_956,N_2540);
xnor U3345 (N_3345,In_1022,In_1305);
or U3346 (N_3346,N_1119,N_246);
or U3347 (N_3347,N_2610,N_1156);
nor U3348 (N_3348,In_1164,In_2335);
or U3349 (N_3349,N_746,N_2795);
or U3350 (N_3350,In_3817,In_889);
or U3351 (N_3351,In_754,N_1030);
nor U3352 (N_3352,N_908,N_2848);
xor U3353 (N_3353,N_1825,In_3949);
nor U3354 (N_3354,In_3760,In_4906);
xor U3355 (N_3355,In_1450,N_2588);
and U3356 (N_3356,N_2682,N_2383);
xnor U3357 (N_3357,In_4211,N_2899);
or U3358 (N_3358,In_2241,N_2932);
nand U3359 (N_3359,In_3761,N_314);
or U3360 (N_3360,In_4779,In_4036);
xor U3361 (N_3361,N_184,N_1784);
xor U3362 (N_3362,N_1641,N_932);
nor U3363 (N_3363,N_2989,In_2791);
xnor U3364 (N_3364,In_570,In_3392);
nor U3365 (N_3365,N_574,N_2961);
nand U3366 (N_3366,N_1918,N_538);
xor U3367 (N_3367,N_2733,N_922);
nor U3368 (N_3368,In_413,N_1964);
nor U3369 (N_3369,N_1919,N_2658);
and U3370 (N_3370,In_973,N_2831);
nor U3371 (N_3371,N_2044,In_1536);
or U3372 (N_3372,In_1369,In_2531);
nor U3373 (N_3373,In_2439,N_2282);
or U3374 (N_3374,N_2043,In_2878);
or U3375 (N_3375,N_2816,In_68);
and U3376 (N_3376,N_2921,In_4061);
nand U3377 (N_3377,In_3580,N_1254);
nor U3378 (N_3378,In_1107,N_2660);
and U3379 (N_3379,In_3178,In_4844);
or U3380 (N_3380,In_3860,In_2423);
nor U3381 (N_3381,N_2849,In_762);
or U3382 (N_3382,N_1492,N_2722);
xnor U3383 (N_3383,In_790,N_1627);
nand U3384 (N_3384,N_462,N_925);
nor U3385 (N_3385,N_2712,N_2050);
nand U3386 (N_3386,N_2776,N_2333);
nand U3387 (N_3387,In_2309,In_131);
xor U3388 (N_3388,N_1146,N_2657);
nor U3389 (N_3389,N_1003,In_2493);
nand U3390 (N_3390,N_2295,N_2318);
or U3391 (N_3391,In_153,In_3426);
nand U3392 (N_3392,N_2678,In_4711);
xor U3393 (N_3393,N_1816,In_476);
nor U3394 (N_3394,In_1960,In_3100);
xnor U3395 (N_3395,In_3639,N_1875);
nand U3396 (N_3396,In_2490,In_4234);
nand U3397 (N_3397,N_851,N_2846);
and U3398 (N_3398,N_2711,In_159);
nor U3399 (N_3399,N_1082,In_4294);
or U3400 (N_3400,N_2284,N_2064);
nor U3401 (N_3401,N_2569,In_3320);
nand U3402 (N_3402,In_3377,In_3042);
and U3403 (N_3403,In_56,N_2446);
or U3404 (N_3404,In_1356,N_2514);
and U3405 (N_3405,N_2836,N_822);
or U3406 (N_3406,In_1116,N_2949);
nor U3407 (N_3407,N_2475,N_692);
or U3408 (N_3408,N_2893,N_2485);
and U3409 (N_3409,N_791,In_765);
xnor U3410 (N_3410,N_2597,N_2708);
nand U3411 (N_3411,N_2823,N_2109);
or U3412 (N_3412,In_895,N_2845);
xnor U3413 (N_3413,N_597,N_2666);
or U3414 (N_3414,N_2438,N_1719);
and U3415 (N_3415,In_4120,N_2739);
and U3416 (N_3416,In_1203,In_2202);
nand U3417 (N_3417,N_2325,In_847);
or U3418 (N_3418,In_4236,In_884);
or U3419 (N_3419,N_1360,In_1862);
and U3420 (N_3420,In_4827,N_2328);
nand U3421 (N_3421,N_2197,In_2797);
nand U3422 (N_3422,N_395,N_2327);
nand U3423 (N_3423,N_1569,N_1852);
nand U3424 (N_3424,N_2655,N_840);
nor U3425 (N_3425,In_1213,In_4950);
nand U3426 (N_3426,In_4497,N_2675);
and U3427 (N_3427,In_2460,N_1302);
xnor U3428 (N_3428,In_3661,In_4741);
nor U3429 (N_3429,N_789,N_2999);
or U3430 (N_3430,In_250,N_1309);
nand U3431 (N_3431,N_2866,In_3626);
nor U3432 (N_3432,N_560,N_2827);
nand U3433 (N_3433,N_2388,N_1980);
xor U3434 (N_3434,N_1831,In_4674);
and U3435 (N_3435,N_907,N_2933);
xnor U3436 (N_3436,N_1170,N_2926);
and U3437 (N_3437,In_781,In_4174);
nor U3438 (N_3438,In_4376,N_2972);
nand U3439 (N_3439,N_2841,In_3826);
nor U3440 (N_3440,N_1402,N_2387);
nor U3441 (N_3441,In_3557,In_1456);
nor U3442 (N_3442,N_1503,N_2012);
nand U3443 (N_3443,In_668,In_3598);
nand U3444 (N_3444,In_262,N_2642);
and U3445 (N_3445,N_2138,N_2447);
nand U3446 (N_3446,N_2794,N_2728);
nor U3447 (N_3447,N_2544,In_1714);
xnor U3448 (N_3448,N_2974,N_2157);
and U3449 (N_3449,N_1079,In_2121);
and U3450 (N_3450,N_2683,N_2602);
or U3451 (N_3451,N_2222,In_2159);
nand U3452 (N_3452,N_591,In_3772);
nand U3453 (N_3453,N_2742,N_1948);
nand U3454 (N_3454,N_914,N_2969);
or U3455 (N_3455,N_2991,N_1024);
nand U3456 (N_3456,In_3558,N_785);
xor U3457 (N_3457,N_2192,N_1924);
xnor U3458 (N_3458,N_2663,N_1415);
xnor U3459 (N_3459,N_2854,In_3676);
and U3460 (N_3460,In_3386,In_2350);
or U3461 (N_3461,N_825,N_2913);
or U3462 (N_3462,N_328,In_3179);
nor U3463 (N_3463,N_2772,N_1065);
and U3464 (N_3464,N_1661,N_1859);
or U3465 (N_3465,N_1303,N_330);
nor U3466 (N_3466,In_3934,N_2584);
or U3467 (N_3467,In_359,N_2956);
nand U3468 (N_3468,N_1159,In_3169);
nor U3469 (N_3469,N_2268,In_2583);
and U3470 (N_3470,N_1770,N_2220);
nor U3471 (N_3471,N_2448,N_1073);
nand U3472 (N_3472,N_1949,In_4408);
or U3473 (N_3473,N_2508,N_2483);
xor U3474 (N_3474,In_2426,In_1639);
or U3475 (N_3475,In_3671,N_2132);
or U3476 (N_3476,N_89,N_2730);
nor U3477 (N_3477,In_2182,N_2731);
nor U3478 (N_3478,N_266,N_2935);
or U3479 (N_3479,N_2929,N_2748);
nor U3480 (N_3480,N_2880,N_1525);
or U3481 (N_3481,In_1130,N_2948);
and U3482 (N_3482,N_2501,N_1822);
xnor U3483 (N_3483,N_1864,N_2763);
and U3484 (N_3484,In_1781,N_798);
nor U3485 (N_3485,N_2267,N_568);
and U3486 (N_3486,In_4970,N_2373);
xnor U3487 (N_3487,N_2531,N_960);
nor U3488 (N_3488,N_2814,N_1296);
or U3489 (N_3489,N_59,N_2598);
nor U3490 (N_3490,N_766,N_2957);
xnor U3491 (N_3491,N_459,N_1691);
or U3492 (N_3492,N_2404,N_2006);
and U3493 (N_3493,In_3347,N_1108);
nor U3494 (N_3494,In_1169,In_908);
or U3495 (N_3495,N_1399,N_1343);
and U3496 (N_3496,N_2074,In_4949);
and U3497 (N_3497,In_3356,In_4776);
xnor U3498 (N_3498,N_1891,N_2599);
xor U3499 (N_3499,N_860,N_2681);
xor U3500 (N_3500,In_499,N_1829);
or U3501 (N_3501,N_1747,N_1367);
nand U3502 (N_3502,N_1584,N_1270);
nand U3503 (N_3503,N_2737,N_2054);
nand U3504 (N_3504,N_883,In_582);
or U3505 (N_3505,N_2261,In_4517);
nand U3506 (N_3506,N_1493,In_4804);
nor U3507 (N_3507,In_3635,In_1951);
xor U3508 (N_3508,N_1761,N_3440);
or U3509 (N_3509,N_2644,N_1991);
nand U3510 (N_3510,N_2596,N_3094);
nand U3511 (N_3511,N_2830,N_890);
nor U3512 (N_3512,In_3140,N_3067);
xor U3513 (N_3513,N_1414,N_3395);
or U3514 (N_3514,N_2901,N_3010);
xor U3515 (N_3515,N_3371,N_2067);
or U3516 (N_3516,N_428,N_2741);
or U3517 (N_3517,N_3294,N_2897);
nand U3518 (N_3518,N_2633,N_2551);
or U3519 (N_3519,N_946,N_2784);
xnor U3520 (N_3520,N_3258,N_2486);
nor U3521 (N_3521,N_3069,N_3063);
xnor U3522 (N_3522,N_2254,N_3488);
and U3523 (N_3523,In_116,N_3231);
and U3524 (N_3524,N_1765,N_2549);
xor U3525 (N_3525,N_2339,N_2015);
and U3526 (N_3526,N_2608,In_716);
xor U3527 (N_3527,In_1902,N_3206);
nor U3528 (N_3528,In_4833,N_1755);
nand U3529 (N_3529,In_3125,N_3448);
nand U3530 (N_3530,N_3381,N_2371);
nand U3531 (N_3531,N_2865,N_2702);
or U3532 (N_3532,N_3159,N_1056);
nand U3533 (N_3533,N_3278,N_3077);
or U3534 (N_3534,N_1682,In_1592);
nand U3535 (N_3535,N_3450,N_2907);
and U3536 (N_3536,In_1588,In_377);
and U3537 (N_3537,N_3302,N_3459);
and U3538 (N_3538,N_1873,N_3148);
nand U3539 (N_3539,In_3501,In_2542);
xnor U3540 (N_3540,N_2912,In_4317);
or U3541 (N_3541,N_2323,N_434);
or U3542 (N_3542,In_4818,N_2858);
xnor U3543 (N_3543,N_2719,N_2308);
or U3544 (N_3544,N_3075,N_3243);
and U3545 (N_3545,N_1515,N_2698);
nor U3546 (N_3546,N_3122,N_3079);
or U3547 (N_3547,N_2785,In_2361);
nand U3548 (N_3548,N_1295,N_2435);
nand U3549 (N_3549,In_1700,N_2262);
or U3550 (N_3550,In_3007,In_3968);
or U3551 (N_3551,N_2638,In_2384);
or U3552 (N_3552,N_819,N_1799);
xor U3553 (N_3553,N_3308,In_1936);
and U3554 (N_3554,N_641,N_3241);
nand U3555 (N_3555,N_2826,In_2498);
or U3556 (N_3556,N_2887,N_1836);
nor U3557 (N_3557,N_406,N_2885);
nand U3558 (N_3558,N_3420,N_1495);
xor U3559 (N_3559,N_3337,N_2710);
xor U3560 (N_3560,N_2992,N_3324);
nand U3561 (N_3561,N_1580,In_4469);
xor U3562 (N_3562,In_3200,N_2911);
nand U3563 (N_3563,N_998,In_972);
and U3564 (N_3564,N_2612,N_3499);
nand U3565 (N_3565,N_2758,N_3326);
nand U3566 (N_3566,N_3037,N_893);
nor U3567 (N_3567,In_4946,N_3312);
nand U3568 (N_3568,N_3264,N_3249);
and U3569 (N_3569,N_3123,N_1006);
nor U3570 (N_3570,N_2442,N_3051);
nor U3571 (N_3571,N_2009,In_4521);
and U3572 (N_3572,N_26,N_2736);
nand U3573 (N_3573,N_1561,N_3307);
and U3574 (N_3574,N_3284,N_1843);
xnor U3575 (N_3575,N_3048,N_2095);
nand U3576 (N_3576,N_1824,N_2922);
and U3577 (N_3577,N_2201,In_13);
and U3578 (N_3578,N_232,N_2504);
nor U3579 (N_3579,N_2931,In_1829);
nand U3580 (N_3580,N_2346,N_3286);
or U3581 (N_3581,N_2798,N_1004);
or U3582 (N_3582,In_3128,N_1955);
or U3583 (N_3583,N_3199,N_3054);
and U3584 (N_3584,N_294,N_3328);
or U3585 (N_3585,N_1507,N_3246);
nor U3586 (N_3586,N_3460,In_1929);
nand U3587 (N_3587,N_2647,N_2771);
or U3588 (N_3588,N_1012,N_1532);
nor U3589 (N_3589,N_3389,N_3049);
or U3590 (N_3590,N_3065,In_4299);
nor U3591 (N_3591,In_3691,N_1294);
nor U3592 (N_3592,N_1681,N_2813);
and U3593 (N_3593,N_3113,N_2543);
nor U3594 (N_3594,N_3379,N_1533);
xor U3595 (N_3595,N_3301,N_1357);
and U3596 (N_3596,N_3432,N_3026);
or U3597 (N_3597,N_717,N_111);
xnor U3598 (N_3598,N_3194,N_2806);
and U3599 (N_3599,N_3036,In_4960);
and U3600 (N_3600,N_3425,In_2911);
nor U3601 (N_3601,N_1431,N_2867);
xor U3602 (N_3602,N_2020,N_2667);
nand U3603 (N_3603,N_3263,N_2303);
xnor U3604 (N_3604,N_3314,N_3035);
nand U3605 (N_3605,N_1847,N_1986);
xnor U3606 (N_3606,N_2451,In_1908);
and U3607 (N_3607,N_497,N_2142);
xnor U3608 (N_3608,N_3491,In_1441);
or U3609 (N_3609,N_3416,In_2622);
nor U3610 (N_3610,In_330,N_3422);
and U3611 (N_3611,N_2164,In_1317);
xnor U3612 (N_3612,N_3350,In_4771);
nand U3613 (N_3613,N_3485,N_1888);
nor U3614 (N_3614,N_2947,N_2634);
xor U3615 (N_3615,N_3449,N_2973);
xnor U3616 (N_3616,N_991,N_2777);
nor U3617 (N_3617,N_3158,N_3368);
or U3618 (N_3618,N_3078,N_3162);
nor U3619 (N_3619,N_509,N_2994);
nor U3620 (N_3620,N_2791,N_3393);
or U3621 (N_3621,N_3346,In_3820);
xor U3622 (N_3622,N_3124,N_3180);
nand U3623 (N_3623,N_2620,N_2264);
nand U3624 (N_3624,N_2839,N_3207);
nor U3625 (N_3625,N_2637,N_3423);
and U3626 (N_3626,N_2033,N_3087);
or U3627 (N_3627,N_2056,In_4743);
nor U3628 (N_3628,N_267,N_3320);
and U3629 (N_3629,N_2345,N_3155);
nor U3630 (N_3630,N_3106,N_905);
nand U3631 (N_3631,In_4412,N_3409);
or U3632 (N_3632,N_874,N_503);
xnor U3633 (N_3633,N_1619,N_2970);
and U3634 (N_3634,N_2186,N_3315);
nor U3635 (N_3635,N_2087,N_3340);
nand U3636 (N_3636,N_2983,N_2154);
xor U3637 (N_3637,N_1563,N_2945);
xnor U3638 (N_3638,N_3082,N_2365);
xor U3639 (N_3639,In_60,In_4345);
nor U3640 (N_3640,N_2238,N_2246);
nand U3641 (N_3641,N_3330,In_1325);
or U3642 (N_3642,N_3404,N_3099);
or U3643 (N_3643,N_2272,N_619);
xor U3644 (N_3644,N_3351,N_3479);
or U3645 (N_3645,In_1838,N_3474);
and U3646 (N_3646,In_1396,N_3107);
or U3647 (N_3647,N_3372,N_2906);
nor U3648 (N_3648,N_3038,In_2951);
xnor U3649 (N_3649,N_664,N_953);
xnor U3650 (N_3650,N_2953,In_3107);
xnor U3651 (N_3651,N_3455,In_3537);
xor U3652 (N_3652,In_4466,N_2693);
xnor U3653 (N_3653,N_3300,N_3221);
or U3654 (N_3654,In_4565,N_3325);
or U3655 (N_3655,N_1308,N_3215);
nand U3656 (N_3656,N_2700,N_1040);
nand U3657 (N_3657,N_3208,N_1723);
xor U3658 (N_3658,N_2471,N_2671);
or U3659 (N_3659,N_1157,In_3926);
xor U3660 (N_3660,N_3084,N_639);
xor U3661 (N_3661,N_3354,N_2161);
and U3662 (N_3662,In_1362,N_3327);
and U3663 (N_3663,N_2908,N_3253);
or U3664 (N_3664,N_2347,N_1646);
xnor U3665 (N_3665,N_2986,N_2889);
nor U3666 (N_3666,N_1771,N_47);
nand U3667 (N_3667,N_3282,N_3390);
or U3668 (N_3668,In_3247,In_1477);
and U3669 (N_3669,N_3471,N_2290);
and U3670 (N_3670,N_2769,N_2586);
nor U3671 (N_3671,N_3001,In_1177);
or U3672 (N_3672,N_3085,N_2083);
or U3673 (N_3673,In_1627,In_2798);
xnor U3674 (N_3674,N_2495,In_2277);
xor U3675 (N_3675,N_2701,N_1839);
and U3676 (N_3676,N_554,N_2219);
or U3677 (N_3677,In_2436,N_1188);
or U3678 (N_3678,N_3000,N_1658);
nand U3679 (N_3679,N_3187,N_3104);
xor U3680 (N_3680,In_2567,N_3118);
nor U3681 (N_3681,N_2242,N_3233);
xor U3682 (N_3682,In_3670,N_2688);
xnor U3683 (N_3683,N_3341,N_3358);
or U3684 (N_3684,In_3177,N_3374);
and U3685 (N_3685,N_614,N_2279);
and U3686 (N_3686,In_2692,N_2622);
and U3687 (N_3687,N_3186,In_1292);
or U3688 (N_3688,N_2461,N_3152);
nand U3689 (N_3689,N_1292,In_2606);
and U3690 (N_3690,N_3343,In_2921);
and U3691 (N_3691,N_2590,In_2138);
nand U3692 (N_3692,In_4157,N_1120);
or U3693 (N_3693,N_3071,N_2799);
nand U3694 (N_3694,N_3133,In_3162);
nor U3695 (N_3695,In_1671,N_2047);
xnor U3696 (N_3696,N_3273,N_3114);
and U3697 (N_3697,In_1009,N_1531);
and U3698 (N_3698,N_3019,N_2579);
or U3699 (N_3699,In_1968,In_126);
xor U3700 (N_3700,N_3109,N_3127);
nand U3701 (N_3701,N_1085,In_1745);
or U3702 (N_3702,N_2046,N_3018);
nand U3703 (N_3703,N_2749,N_3046);
or U3704 (N_3704,N_3008,In_928);
nand U3705 (N_3705,N_2882,N_2927);
nand U3706 (N_3706,N_1959,N_414);
and U3707 (N_3707,N_2847,N_2564);
nor U3708 (N_3708,N_3059,N_3034);
and U3709 (N_3709,N_3201,N_3211);
or U3710 (N_3710,N_1447,N_2937);
or U3711 (N_3711,N_3213,N_2434);
and U3712 (N_3712,N_3212,In_3852);
and U3713 (N_3713,In_3885,N_3387);
nor U3714 (N_3714,In_2229,N_3295);
xor U3715 (N_3715,N_3424,N_2099);
xor U3716 (N_3716,N_1914,N_1624);
nand U3717 (N_3717,N_2237,N_3403);
or U3718 (N_3718,In_2158,N_2787);
xnor U3719 (N_3719,N_2030,In_486);
xnor U3720 (N_3720,N_1176,In_1654);
xnor U3721 (N_3721,N_3120,N_3369);
nor U3722 (N_3722,N_2420,In_1472);
nor U3723 (N_3723,N_2482,In_862);
nor U3724 (N_3724,N_2524,N_1583);
or U3725 (N_3725,N_2717,N_2759);
and U3726 (N_3726,In_2665,N_3384);
nand U3727 (N_3727,N_1573,N_2706);
nand U3728 (N_3728,N_2002,N_2407);
nand U3729 (N_3729,N_783,N_1850);
and U3730 (N_3730,N_2656,N_3470);
and U3731 (N_3731,N_3198,N_2824);
nand U3732 (N_3732,N_1083,N_2059);
or U3733 (N_3733,N_677,In_1519);
nand U3734 (N_3734,In_1649,N_3003);
and U3735 (N_3735,In_1775,N_2723);
xor U3736 (N_3736,N_3050,N_678);
nand U3737 (N_3737,In_112,In_900);
and U3738 (N_3738,In_4099,N_3197);
and U3739 (N_3739,N_3149,In_3929);
nand U3740 (N_3740,In_694,N_2910);
nor U3741 (N_3741,N_3394,In_2475);
nor U3742 (N_3742,N_2191,N_3032);
xor U3743 (N_3743,N_2726,N_2463);
or U3744 (N_3744,N_2750,In_3887);
or U3745 (N_3745,N_1698,N_3115);
xor U3746 (N_3746,N_3406,N_2107);
and U3747 (N_3747,N_2844,N_3280);
xor U3748 (N_3748,In_4767,N_2223);
and U3749 (N_3749,N_3150,N_3184);
or U3750 (N_3750,N_2255,N_1242);
xnor U3751 (N_3751,N_2967,N_2565);
nand U3752 (N_3752,In_1680,In_3350);
or U3753 (N_3753,In_2607,N_2566);
or U3754 (N_3754,N_2399,N_3042);
and U3755 (N_3755,N_3434,N_2069);
nand U3756 (N_3756,N_1908,In_733);
nand U3757 (N_3757,N_3380,N_1534);
xnor U3758 (N_3758,N_2093,N_1476);
xor U3759 (N_3759,N_719,N_1927);
xnor U3760 (N_3760,N_3495,N_2545);
nor U3761 (N_3761,N_1217,N_2965);
or U3762 (N_3762,N_2274,In_810);
or U3763 (N_3763,N_2519,In_732);
xnor U3764 (N_3764,N_1536,N_2995);
and U3765 (N_3765,N_3247,In_1560);
and U3766 (N_3766,N_1045,N_1768);
and U3767 (N_3767,In_853,N_2247);
or U3768 (N_3768,N_3012,N_2195);
xor U3769 (N_3769,N_2500,N_1764);
and U3770 (N_3770,N_2166,N_3494);
or U3771 (N_3771,In_1782,N_2153);
or U3772 (N_3772,N_2721,N_2892);
or U3773 (N_3773,In_1290,N_2976);
nand U3774 (N_3774,N_467,In_3891);
nor U3775 (N_3775,N_2051,N_3259);
nor U3776 (N_3776,N_3086,N_1763);
or U3777 (N_3777,In_452,N_1805);
or U3778 (N_3778,N_3375,N_2762);
xnor U3779 (N_3779,N_3081,In_282);
or U3780 (N_3780,N_1136,N_3292);
and U3781 (N_3781,N_102,N_1581);
and U3782 (N_3782,N_2450,N_2793);
or U3783 (N_3783,N_2925,N_148);
or U3784 (N_3784,N_2338,N_3335);
or U3785 (N_3785,N_2560,N_2951);
nor U3786 (N_3786,N_2664,N_3347);
xnor U3787 (N_3787,N_3256,N_376);
nand U3788 (N_3788,N_3009,N_407);
nor U3789 (N_3789,N_2833,N_1696);
or U3790 (N_3790,In_2226,In_4886);
and U3791 (N_3791,N_2460,In_4335);
xor U3792 (N_3792,In_661,N_15);
nand U3793 (N_3793,N_1840,In_1665);
nor U3794 (N_3794,N_3168,N_3296);
nand U3795 (N_3795,N_383,N_3285);
or U3796 (N_3796,N_3480,N_3417);
and U3797 (N_3797,N_3428,N_2766);
or U3798 (N_3798,N_3245,In_1019);
nand U3799 (N_3799,N_2024,N_3193);
nand U3800 (N_3800,N_2883,N_3021);
and U3801 (N_3801,In_2749,N_3016);
xnor U3802 (N_3802,N_1817,In_2098);
nand U3803 (N_3803,N_3402,N_3452);
or U3804 (N_3804,In_2504,N_2314);
or U3805 (N_3805,N_2979,N_2258);
or U3806 (N_3806,N_3287,N_3265);
nand U3807 (N_3807,N_153,In_4562);
xor U3808 (N_3808,N_3056,N_2810);
and U3809 (N_3809,In_789,N_2269);
or U3810 (N_3810,In_1573,In_4919);
nor U3811 (N_3811,N_2520,N_1633);
and U3812 (N_3812,N_3465,N_3200);
nor U3813 (N_3813,N_3323,In_1044);
and U3814 (N_3814,N_3454,N_2468);
or U3815 (N_3815,N_3092,N_3289);
nor U3816 (N_3816,N_931,N_3142);
and U3817 (N_3817,N_3293,N_3329);
or U3818 (N_3818,N_2704,In_123);
and U3819 (N_3819,N_3005,N_275);
or U3820 (N_3820,N_3370,N_2100);
xor U3821 (N_3821,N_3283,N_3476);
and U3822 (N_3822,In_2117,N_2553);
nor U3823 (N_3823,N_3468,N_726);
xnor U3824 (N_3824,N_1545,N_3041);
nor U3825 (N_3825,N_3209,N_3111);
or U3826 (N_3826,N_2825,N_1511);
xnor U3827 (N_3827,N_1601,N_537);
xor U3828 (N_3828,In_4413,In_310);
and U3829 (N_3829,In_3593,In_1757);
or U3830 (N_3830,N_2811,N_3397);
nor U3831 (N_3831,N_3110,N_3281);
nand U3832 (N_3832,N_2718,N_2600);
nand U3833 (N_3833,N_1797,N_2311);
nand U3834 (N_3834,N_2729,N_3177);
nor U3835 (N_3835,N_2382,N_3291);
nor U3836 (N_3836,N_2606,N_2803);
xor U3837 (N_3837,N_3456,N_3316);
nand U3838 (N_3838,N_3429,N_2167);
nor U3839 (N_3839,N_1685,N_3181);
xnor U3840 (N_3840,In_696,N_2198);
or U3841 (N_3841,N_1693,N_3458);
or U3842 (N_3842,N_3108,N_1700);
nor U3843 (N_3843,N_3267,N_2022);
nand U3844 (N_3844,In_379,N_3382);
nand U3845 (N_3845,N_1976,In_634);
xor U3846 (N_3846,N_3436,N_3386);
or U3847 (N_3847,N_2175,N_1662);
nand U3848 (N_3848,In_1544,N_3064);
and U3849 (N_3849,N_3131,N_2977);
and U3850 (N_3850,N_2964,In_3568);
or U3851 (N_3851,N_2832,In_763);
and U3852 (N_3852,N_1773,N_2422);
xor U3853 (N_3853,N_3288,In_3719);
xnor U3854 (N_3854,In_1849,N_3310);
nor U3855 (N_3855,In_2287,N_2297);
and U3856 (N_3856,N_3144,In_4341);
or U3857 (N_3857,N_3451,N_1746);
xnor U3858 (N_3858,In_3896,N_3091);
nand U3859 (N_3859,N_3160,N_3344);
xnor U3860 (N_3860,N_2651,N_3385);
and U3861 (N_3861,N_3029,N_3473);
or U3862 (N_3862,In_1289,N_3205);
xor U3863 (N_3863,N_1332,N_2668);
nor U3864 (N_3864,In_273,In_3292);
and U3865 (N_3865,N_2905,N_3189);
xnor U3866 (N_3866,In_1565,N_3222);
xnor U3867 (N_3867,In_907,N_1666);
or U3868 (N_3868,In_1043,In_3404);
nand U3869 (N_3869,In_1080,N_2653);
nand U3870 (N_3870,In_3410,N_3236);
nor U3871 (N_3871,N_3317,N_3490);
or U3872 (N_3872,N_1688,N_1437);
nor U3873 (N_3873,N_3225,In_4017);
and U3874 (N_3874,N_3153,N_3028);
nor U3875 (N_3875,In_257,N_2576);
nor U3876 (N_3876,N_3146,N_1125);
nor U3877 (N_3877,N_1304,N_2414);
or U3878 (N_3878,In_4393,N_2426);
xnor U3879 (N_3879,N_1858,N_765);
nor U3880 (N_3880,N_3363,N_1958);
and U3881 (N_3881,In_1348,N_786);
xor U3882 (N_3882,N_3360,N_3483);
nand U3883 (N_3883,In_1131,In_2024);
nor U3884 (N_3884,N_3255,In_1432);
nor U3885 (N_3885,In_437,N_2092);
xor U3886 (N_3886,N_533,N_2788);
xnor U3887 (N_3887,N_3044,N_2299);
nor U3888 (N_3888,N_2856,In_1065);
or U3889 (N_3889,N_2828,In_426);
xor U3890 (N_3890,N_2114,N_3006);
xnor U3891 (N_3891,N_926,N_3413);
or U3892 (N_3892,N_1416,N_3164);
nand U3893 (N_3893,N_2955,N_2548);
or U3894 (N_3894,N_3447,N_1866);
or U3895 (N_3895,N_2580,N_2745);
and U3896 (N_3896,In_2698,N_1506);
nor U3897 (N_3897,N_3224,N_3342);
nand U3898 (N_3898,N_2467,N_2200);
nand U3899 (N_3899,N_3421,N_3105);
nor U3900 (N_3900,In_4998,N_3234);
nor U3901 (N_3901,N_3481,N_1358);
or U3902 (N_3902,In_2649,N_2466);
nor U3903 (N_3903,In_3548,N_3126);
nand U3904 (N_3904,In_1002,N_3377);
xnor U3905 (N_3905,In_3134,In_4639);
nor U3906 (N_3906,N_2919,N_2205);
xor U3907 (N_3907,N_1214,N_2221);
xor U3908 (N_3908,N_1807,In_1011);
or U3909 (N_3909,In_4121,N_3173);
nand U3910 (N_3910,N_1890,N_2822);
nor U3911 (N_3911,N_3128,In_4577);
nor U3912 (N_3912,In_2633,N_2626);
and U3913 (N_3913,N_1683,N_1462);
or U3914 (N_3914,N_2348,In_2569);
and U3915 (N_3915,In_2789,In_1481);
nor U3916 (N_3916,In_4091,N_3392);
or U3917 (N_3917,N_2809,N_1945);
nand U3918 (N_3918,N_1731,N_3176);
xnor U3919 (N_3919,N_1464,In_2223);
nor U3920 (N_3920,In_1092,N_2694);
and U3921 (N_3921,N_3446,N_3378);
and U3922 (N_3922,N_492,In_4279);
or U3923 (N_3923,N_2812,N_1049);
or U3924 (N_3924,N_3414,N_387);
nor U3925 (N_3925,N_3174,N_2614);
or U3926 (N_3926,N_2690,N_3229);
and U3927 (N_3927,N_2049,N_3100);
or U3928 (N_3928,N_2503,N_1084);
xor U3929 (N_3929,N_3356,N_2023);
nor U3930 (N_3930,N_2213,N_3102);
and U3931 (N_3931,N_779,N_2244);
or U3932 (N_3932,N_3055,N_2792);
nand U3933 (N_3933,N_3017,In_2195);
nor U3934 (N_3934,N_1166,N_3306);
xor U3935 (N_3935,N_3066,N_2306);
and U3936 (N_3936,N_3388,N_2820);
nor U3937 (N_3937,N_1059,In_4658);
xnor U3938 (N_3938,N_2817,N_10);
nor U3939 (N_3939,In_2469,N_3298);
nand U3940 (N_3940,N_1338,N_2583);
or U3941 (N_3941,N_3401,N_3031);
or U3942 (N_3942,N_3033,N_1893);
nand U3943 (N_3943,In_2563,N_2591);
nor U3944 (N_3944,N_2930,In_2324);
nand U3945 (N_3945,N_2918,N_3154);
nand U3946 (N_3946,N_3175,N_1513);
xnor U3947 (N_3947,N_3134,N_2645);
or U3948 (N_3948,N_3223,N_2952);
nor U3949 (N_3949,N_1568,In_3591);
nor U3950 (N_3950,In_4038,N_3254);
or U3951 (N_3951,N_3463,N_1566);
nor U3952 (N_3952,N_2703,N_2541);
and U3953 (N_3953,N_2405,N_3353);
nor U3954 (N_3954,N_1738,N_2071);
and U3955 (N_3955,In_2906,N_3216);
nor U3956 (N_3956,N_3430,N_1766);
or U3957 (N_3957,N_3166,In_2235);
or U3958 (N_3958,N_2199,In_2331);
nand U3959 (N_3959,N_2859,N_3191);
or U3960 (N_3960,N_2341,N_2558);
xnor U3961 (N_3961,N_81,In_115);
or U3962 (N_3962,N_1389,In_1435);
nor U3963 (N_3963,N_809,N_2016);
xnor U3964 (N_3964,N_1779,N_1484);
nand U3965 (N_3965,N_2649,In_3997);
nand U3966 (N_3966,N_356,N_1751);
nor U3967 (N_3967,N_3014,N_3352);
nand U3968 (N_3968,N_2389,N_1487);
or U3969 (N_3969,N_535,N_1353);
nand U3970 (N_3970,N_2276,N_3489);
nor U3971 (N_3971,N_2630,N_2695);
nand U3972 (N_3972,N_3015,N_3274);
nand U3973 (N_3973,N_1273,N_2601);
nand U3974 (N_3974,In_4005,N_3269);
and U3975 (N_3975,N_3023,In_1742);
or U3976 (N_3976,N_216,In_3242);
nand U3977 (N_3977,N_3367,In_2981);
nand U3978 (N_3978,N_3203,N_3047);
xor U3979 (N_3979,N_2017,N_3096);
xor U3980 (N_3980,N_3266,In_4178);
nand U3981 (N_3981,N_3147,N_3411);
xnor U3982 (N_3982,N_3355,N_3348);
nor U3983 (N_3983,N_3024,N_3469);
or U3984 (N_3984,In_1283,N_2725);
xor U3985 (N_3985,In_2376,N_2552);
xor U3986 (N_3986,N_2735,N_3275);
xnor U3987 (N_3987,N_2756,N_3410);
nor U3988 (N_3988,In_2406,N_2575);
nor U3989 (N_3989,N_3376,In_3583);
nand U3990 (N_3990,N_1628,N_3362);
or U3991 (N_3991,N_3299,N_2895);
xnor U3992 (N_3992,N_512,N_3262);
and U3993 (N_3993,N_2636,N_2578);
nor U3994 (N_3994,N_3244,N_3196);
and U3995 (N_3995,N_3361,N_2819);
nor U3996 (N_3996,N_2510,N_3486);
nand U3997 (N_3997,N_3027,N_1777);
nand U3998 (N_3998,N_2275,N_3313);
nand U3999 (N_3999,N_3169,N_3138);
nand U4000 (N_4000,N_3536,N_590);
nand U4001 (N_4001,In_2694,N_3725);
nor U4002 (N_4002,N_3741,N_3606);
and U4003 (N_4003,N_1370,In_3538);
xor U4004 (N_4004,N_1558,N_3778);
nand U4005 (N_4005,N_2589,In_481);
xor U4006 (N_4006,N_716,In_43);
xnor U4007 (N_4007,N_2251,N_3880);
or U4008 (N_4008,N_2370,N_3513);
and U4009 (N_4009,N_2582,N_3912);
or U4010 (N_4010,N_3866,N_2436);
and U4011 (N_4011,N_3807,N_2896);
or U4012 (N_4012,In_690,N_2527);
or U4013 (N_4013,N_3603,N_3250);
nor U4014 (N_4014,N_3461,In_4973);
xnor U4015 (N_4015,N_1483,N_2802);
or U4016 (N_4016,N_2917,In_1945);
and U4017 (N_4017,N_2474,N_3228);
nor U4018 (N_4018,N_3934,N_3730);
xnor U4019 (N_4019,N_3586,N_3841);
or U4020 (N_4020,N_2641,N_3692);
nand U4021 (N_4021,In_2879,N_3568);
xor U4022 (N_4022,N_3982,N_2494);
xnor U4023 (N_4023,In_4096,N_3659);
xor U4024 (N_4024,N_3562,N_3678);
nor U4025 (N_4025,N_1985,N_2287);
or U4026 (N_4026,In_35,N_3530);
nor U4027 (N_4027,N_3204,N_1943);
and U4028 (N_4028,N_3673,N_3622);
and U4029 (N_4029,N_3574,N_3101);
and U4030 (N_4030,N_3573,N_3837);
nor U4031 (N_4031,N_2343,In_8);
nand U4032 (N_4032,N_3710,N_3339);
nor U4033 (N_4033,N_3412,N_1678);
or U4034 (N_4034,N_3058,N_3878);
or U4035 (N_4035,N_3702,N_1508);
nand U4036 (N_4036,N_3969,N_3801);
nor U4037 (N_4037,N_1567,N_3439);
and U4038 (N_4038,N_3501,N_1947);
or U4039 (N_4039,N_2232,In_1099);
nand U4040 (N_4040,N_3167,N_3804);
xor U4041 (N_4041,N_3681,N_3235);
nor U4042 (N_4042,N_3475,N_3698);
and U4043 (N_4043,N_3525,N_2713);
nor U4044 (N_4044,In_4890,In_3084);
and U4045 (N_4045,N_3917,N_3090);
and U4046 (N_4046,N_3727,N_2412);
nand U4047 (N_4047,N_3514,N_3179);
nand U4048 (N_4048,N_3701,In_2181);
nand U4049 (N_4049,N_3947,N_3610);
nand U4050 (N_4050,N_1982,N_686);
nor U4051 (N_4051,N_3680,N_3214);
xor U4052 (N_4052,In_719,N_3443);
and U4053 (N_4053,N_3493,N_3578);
nand U4054 (N_4054,N_180,In_988);
and U4055 (N_4055,N_3635,N_3013);
nor U4056 (N_4056,N_3997,N_3759);
nand U4057 (N_4057,N_3498,N_3823);
xor U4058 (N_4058,N_1287,N_3004);
and U4059 (N_4059,N_3140,In_3215);
or U4060 (N_4060,N_3336,N_3157);
xor U4061 (N_4061,N_3545,N_3931);
nand U4062 (N_4062,N_3137,N_3400);
xnor U4063 (N_4063,N_3894,N_3643);
nand U4064 (N_4064,In_2720,N_3760);
nand U4065 (N_4065,N_3068,N_3074);
xor U4066 (N_4066,N_3775,N_1057);
xnor U4067 (N_4067,N_3967,N_3549);
nand U4068 (N_4068,N_3986,In_664);
xnor U4069 (N_4069,N_3851,N_3672);
xor U4070 (N_4070,N_3195,N_3773);
nand U4071 (N_4071,N_3093,N_2377);
nand U4072 (N_4072,N_3852,N_3887);
xnor U4073 (N_4073,In_2129,N_3910);
xor U4074 (N_4074,N_3943,N_2505);
xor U4075 (N_4075,N_3901,N_3509);
nor U4076 (N_4076,In_3124,N_2031);
and U4077 (N_4077,N_3136,In_4859);
or U4078 (N_4078,N_446,N_3828);
nand U4079 (N_4079,N_1277,N_3478);
and U4080 (N_4080,N_3708,N_3752);
and U4081 (N_4081,In_4869,N_3579);
nor U4082 (N_4082,N_3699,N_918);
xnor U4083 (N_4083,N_3952,N_3407);
and U4084 (N_4084,N_3713,N_3057);
nand U4085 (N_4085,In_2185,N_3666);
xor U4086 (N_4086,N_3620,N_1625);
xnor U4087 (N_4087,N_3563,N_3500);
and U4088 (N_4088,N_3898,N_776);
nor U4089 (N_4089,N_3572,N_3891);
and U4090 (N_4090,N_3884,N_3251);
nor U4091 (N_4091,N_3913,N_3125);
xor U4092 (N_4092,N_596,N_2555);
xnor U4093 (N_4093,N_3944,N_3897);
or U4094 (N_4094,N_2115,N_3634);
xnor U4095 (N_4095,N_3627,N_3321);
and U4096 (N_4096,N_3865,N_3960);
xnor U4097 (N_4097,N_3663,N_3818);
xnor U4098 (N_4098,N_3918,In_3522);
and U4099 (N_4099,N_3805,N_3889);
or U4100 (N_4100,N_3905,N_1923);
or U4101 (N_4101,In_2100,N_2676);
nand U4102 (N_4102,N_2607,In_3421);
or U4103 (N_4103,N_3405,N_3747);
nand U4104 (N_4104,N_3808,N_3846);
nor U4105 (N_4105,In_4942,N_3743);
nand U4106 (N_4106,N_3540,N_3772);
or U4107 (N_4107,N_3958,N_2035);
nor U4108 (N_4108,N_2465,N_2679);
xnor U4109 (N_4109,N_3650,N_3873);
and U4110 (N_4110,In_3445,N_3881);
nor U4111 (N_4111,N_3976,N_3613);
xor U4112 (N_4112,N_2898,N_3726);
or U4113 (N_4113,N_1162,N_3571);
xor U4114 (N_4114,N_3872,N_3970);
and U4115 (N_4115,N_3819,N_3532);
nor U4116 (N_4116,N_3145,N_3399);
and U4117 (N_4117,N_3529,N_3860);
and U4118 (N_4118,N_3700,N_3116);
xor U4119 (N_4119,N_3585,N_3319);
xnor U4120 (N_4120,N_3826,N_3564);
xor U4121 (N_4121,N_3629,N_3297);
xor U4122 (N_4122,N_3861,In_1414);
nor U4123 (N_4123,N_3924,N_1717);
or U4124 (N_4124,N_3318,N_2753);
and U4125 (N_4125,N_3641,N_2871);
or U4126 (N_4126,N_3900,N_3276);
nand U4127 (N_4127,N_2559,N_2080);
and U4128 (N_4128,N_3217,N_2506);
or U4129 (N_4129,In_2378,N_186);
nor U4130 (N_4130,N_3950,N_3492);
nor U4131 (N_4131,N_1810,N_3636);
nor U4132 (N_4132,N_3978,N_3907);
and U4133 (N_4133,N_1268,In_4043);
and U4134 (N_4134,N_3906,In_4302);
and U4135 (N_4135,N_3533,N_1800);
and U4136 (N_4136,N_2393,N_3761);
nor U4137 (N_4137,N_3914,N_3979);
xnor U4138 (N_4138,N_3121,N_3868);
nor U4139 (N_4139,N_3656,N_1632);
or U4140 (N_4140,N_3239,N_2821);
nor U4141 (N_4141,N_3512,N_3467);
nor U4142 (N_4142,N_3756,N_3604);
or U4143 (N_4143,N_3838,N_2873);
and U4144 (N_4144,N_3558,N_2075);
nor U4145 (N_4145,N_3528,N_3011);
nor U4146 (N_4146,N_3926,N_3795);
xor U4147 (N_4147,In_4308,N_2440);
nor U4148 (N_4148,N_3771,N_3770);
nand U4149 (N_4149,N_3190,N_3553);
xnor U4150 (N_4150,N_3602,N_3002);
or U4151 (N_4151,N_3630,N_3832);
or U4152 (N_4152,N_2829,N_3991);
and U4153 (N_4153,N_3734,N_3728);
or U4154 (N_4154,N_3915,N_3764);
nor U4155 (N_4155,N_3848,N_3651);
or U4156 (N_4156,N_3511,N_1036);
and U4157 (N_4157,N_2542,N_3431);
nand U4158 (N_4158,N_3592,N_3981);
nor U4159 (N_4159,N_3129,In_2025);
or U4160 (N_4160,N_2928,N_3694);
or U4161 (N_4161,N_3597,N_61);
nand U4162 (N_4162,N_3909,N_3060);
nor U4163 (N_4163,N_2574,N_679);
xnor U4164 (N_4164,In_4560,N_3793);
xor U4165 (N_4165,N_3497,N_3835);
nand U4166 (N_4166,N_3565,N_3645);
nor U4167 (N_4167,N_3802,N_3677);
or U4168 (N_4168,N_3812,N_2743);
xor U4169 (N_4169,N_3715,N_3218);
nand U4170 (N_4170,N_3272,N_3437);
nor U4171 (N_4171,N_3980,N_3594);
xnor U4172 (N_4172,N_3631,N_3987);
nor U4173 (N_4173,In_4004,N_3615);
or U4174 (N_4174,N_3591,N_2837);
nand U4175 (N_4175,N_2674,N_3863);
and U4176 (N_4176,N_3797,N_3248);
nand U4177 (N_4177,N_3345,N_2686);
nor U4178 (N_4178,N_3665,N_2408);
and U4179 (N_4179,In_1199,N_3847);
nor U4180 (N_4180,N_519,N_19);
and U4181 (N_4181,N_3570,N_3908);
nand U4182 (N_4182,N_2746,N_3977);
xor U4183 (N_4183,N_3445,N_3238);
nand U4184 (N_4184,N_3453,In_2801);
nor U4185 (N_4185,N_3151,N_3830);
and U4186 (N_4186,N_3030,N_3040);
or U4187 (N_4187,N_3739,In_1069);
and U4188 (N_4188,N_3538,N_3202);
and U4189 (N_4189,N_3911,N_1128);
or U4190 (N_4190,N_3813,N_3457);
nand U4191 (N_4191,In_4856,N_3724);
nor U4192 (N_4192,N_3920,N_3607);
nand U4193 (N_4193,N_2170,N_3053);
xnor U4194 (N_4194,N_3616,N_3955);
or U4195 (N_4195,N_3675,N_933);
xnor U4196 (N_4196,In_2205,N_3810);
nand U4197 (N_4197,N_3933,In_3590);
or U4198 (N_4198,N_3751,N_3798);
or U4199 (N_4199,N_3141,N_1597);
nand U4200 (N_4200,N_981,In_602);
and U4201 (N_4201,N_3964,N_1787);
or U4202 (N_4202,N_2513,N_3855);
and U4203 (N_4203,N_3716,In_4098);
and U4204 (N_4204,N_3596,N_3945);
nand U4205 (N_4205,N_3043,N_3686);
or U4206 (N_4206,N_3829,N_3780);
or U4207 (N_4207,N_1041,N_3062);
nor U4208 (N_4208,N_3112,N_3858);
nor U4209 (N_4209,In_3573,N_3261);
nor U4210 (N_4210,In_3160,N_1236);
and U4211 (N_4211,N_3738,N_2843);
nor U4212 (N_4212,N_3357,N_3279);
and U4213 (N_4213,N_3640,N_3589);
nand U4214 (N_4214,N_3322,N_3618);
nor U4215 (N_4215,In_2919,N_3583);
and U4216 (N_4216,N_3661,N_2379);
nand U4217 (N_4217,N_3117,N_3587);
or U4218 (N_4218,N_3839,N_2643);
and U4219 (N_4219,N_3814,N_3623);
xor U4220 (N_4220,N_1540,In_1053);
and U4221 (N_4221,In_267,N_1920);
xor U4222 (N_4222,N_2624,N_3824);
nor U4223 (N_4223,In_1922,N_2425);
and U4224 (N_4224,N_3521,N_1334);
or U4225 (N_4225,N_1579,N_3506);
or U4226 (N_4226,N_665,N_3693);
and U4227 (N_4227,N_1600,N_2751);
and U4228 (N_4228,N_3626,N_3840);
xnor U4229 (N_4229,N_3925,N_3025);
and U4230 (N_4230,N_3546,N_3888);
xor U4231 (N_4231,N_531,N_3704);
and U4232 (N_4232,N_3598,N_3785);
nor U4233 (N_4233,N_2416,N_3435);
nand U4234 (N_4234,N_3608,N_2715);
xor U4235 (N_4235,N_3720,N_3849);
nor U4236 (N_4236,N_3737,N_3842);
xnor U4237 (N_4237,N_3577,N_3242);
and U4238 (N_4238,N_3783,N_3582);
xor U4239 (N_4239,N_3268,N_3938);
nand U4240 (N_4240,N_3083,N_3895);
xnor U4241 (N_4241,N_2808,In_3998);
nand U4242 (N_4242,N_1371,N_3763);
and U4243 (N_4243,N_2517,N_1243);
nor U4244 (N_4244,N_3237,N_1202);
and U4245 (N_4245,N_3526,N_3088);
nor U4246 (N_4246,N_3754,N_3648);
and U4247 (N_4247,N_2946,In_3908);
nand U4248 (N_4248,N_3338,N_3729);
and U4249 (N_4249,N_3182,N_3788);
and U4250 (N_4250,N_3975,N_3717);
and U4251 (N_4251,N_3796,N_3966);
or U4252 (N_4252,N_2277,N_3718);
nor U4253 (N_4253,N_3444,N_3803);
or U4254 (N_4254,In_2833,N_1518);
xor U4255 (N_4255,N_2062,N_3935);
nand U4256 (N_4256,N_3647,N_2916);
or U4257 (N_4257,In_1497,N_3921);
or U4258 (N_4258,N_3867,N_3876);
nand U4259 (N_4259,N_3171,N_3484);
or U4260 (N_4260,N_3581,N_3080);
xor U4261 (N_4261,N_3304,N_3580);
or U4262 (N_4262,N_2639,N_3990);
nand U4263 (N_4263,N_3968,N_3426);
nand U4264 (N_4264,N_1190,N_3667);
nor U4265 (N_4265,N_2786,N_3566);
nor U4266 (N_4266,N_784,N_3595);
nor U4267 (N_4267,N_3714,N_589);
nor U4268 (N_4268,N_1222,N_3954);
xnor U4269 (N_4269,N_342,In_2590);
xor U4270 (N_4270,N_2547,N_3309);
xor U4271 (N_4271,N_3786,N_3172);
or U4272 (N_4272,N_3505,N_613);
or U4273 (N_4273,In_1433,N_3719);
nor U4274 (N_4274,N_3588,N_3210);
and U4275 (N_4275,In_4370,N_909);
nor U4276 (N_4276,N_3707,In_2333);
and U4277 (N_4277,N_2137,N_3709);
and U4278 (N_4278,N_3649,N_3520);
and U4279 (N_4279,N_3517,N_3736);
or U4280 (N_4280,N_3790,N_3518);
nor U4281 (N_4281,N_2857,N_3653);
nor U4282 (N_4282,N_3541,N_3612);
nor U4283 (N_4283,In_4354,In_2599);
xor U4284 (N_4284,N_2309,N_3932);
nand U4285 (N_4285,N_3559,N_3857);
nor U4286 (N_4286,N_3922,N_3877);
nand U4287 (N_4287,N_2662,N_705);
xnor U4288 (N_4288,N_3682,N_3904);
nor U4289 (N_4289,N_3961,N_3687);
nand U4290 (N_4290,N_2672,N_3644);
xnor U4291 (N_4291,N_3496,N_3836);
xnor U4292 (N_4292,N_3519,N_3902);
nand U4293 (N_4293,N_2392,N_156);
or U4294 (N_4294,N_3948,N_2613);
nand U4295 (N_4295,N_3311,N_2966);
nor U4296 (N_4296,N_1833,N_2349);
nand U4297 (N_4297,N_3537,N_3590);
or U4298 (N_4298,N_3834,N_3984);
and U4299 (N_4299,N_3072,N_3703);
nor U4300 (N_4300,N_3601,N_3776);
nor U4301 (N_4301,N_3742,N_2573);
and U4302 (N_4302,N_3799,In_1366);
nand U4303 (N_4303,N_3879,N_3373);
and U4304 (N_4304,N_3784,N_1780);
or U4305 (N_4305,In_759,N_3816);
nor U4306 (N_4306,N_3482,N_2801);
nand U4307 (N_4307,N_3531,N_2113);
nor U4308 (N_4308,In_4552,N_3185);
and U4309 (N_4309,N_3192,N_1741);
or U4310 (N_4310,N_3535,N_1903);
or U4311 (N_4311,N_3706,N_3561);
xnor U4312 (N_4312,N_2522,N_2550);
xnor U4313 (N_4313,N_3972,In_2908);
xnor U4314 (N_4314,N_3923,N_3504);
and U4315 (N_4315,N_3551,N_3232);
nand U4316 (N_4316,N_2778,N_2561);
nor U4317 (N_4317,N_3765,N_3614);
xor U4318 (N_4318,N_3662,N_3359);
xor U4319 (N_4319,N_3441,N_3119);
xnor U4320 (N_4320,N_306,N_2673);
or U4321 (N_4321,N_3170,N_3766);
xor U4322 (N_4322,N_3749,N_3625);
nor U4323 (N_4323,N_3953,N_3696);
nand U4324 (N_4324,N_3774,N_3230);
or U4325 (N_4325,N_3864,N_3523);
or U4326 (N_4326,N_3815,N_3098);
nand U4327 (N_4327,N_2886,N_3745);
xnor U4328 (N_4328,N_3856,N_3748);
or U4329 (N_4329,N_3593,N_3637);
nor U4330 (N_4330,N_3227,N_351);
and U4331 (N_4331,N_1739,In_711);
or U4332 (N_4332,In_333,N_3557);
nor U4333 (N_4333,N_3721,N_3507);
and U4334 (N_4334,In_4137,N_3022);
nand U4335 (N_4335,N_3165,N_3963);
nand U4336 (N_4336,In_4336,N_2958);
and U4337 (N_4337,N_2512,N_3632);
xnor U4338 (N_4338,N_2707,N_2714);
or U4339 (N_4339,N_3472,N_3477);
and U4340 (N_4340,N_3899,In_1227);
or U4341 (N_4341,N_2903,In_4456);
and U4342 (N_4342,N_1395,N_3464);
and U4343 (N_4343,N_2716,N_3854);
xnor U4344 (N_4344,N_2014,N_2362);
or U4345 (N_4345,N_2366,In_1436);
and U4346 (N_4346,N_3791,N_3903);
or U4347 (N_4347,N_3624,N_3219);
or U4348 (N_4348,In_3046,N_3039);
or U4349 (N_4349,In_4437,N_2923);
or U4350 (N_4350,N_3845,N_3886);
or U4351 (N_4351,N_3705,N_2427);
or U4352 (N_4352,N_3668,N_3466);
or U4353 (N_4353,N_3527,N_3271);
nor U4354 (N_4354,N_3391,N_3366);
nor U4355 (N_4355,N_2767,N_3995);
nor U4356 (N_4356,N_3697,N_3132);
or U4357 (N_4357,N_3781,N_3733);
nand U4358 (N_4358,N_3052,N_1526);
or U4359 (N_4359,N_3691,N_3188);
and U4360 (N_4360,N_3642,N_3735);
and U4361 (N_4361,N_3660,N_476);
nor U4362 (N_4362,N_3787,N_3103);
nand U4363 (N_4363,N_3503,N_3020);
and U4364 (N_4364,N_3290,N_3685);
and U4365 (N_4365,N_3516,In_2122);
and U4366 (N_4366,N_3270,N_3850);
xor U4367 (N_4367,In_2170,N_3962);
xnor U4368 (N_4368,N_3821,N_3628);
and U4369 (N_4369,In_4726,N_3916);
or U4370 (N_4370,N_2621,N_3746);
xor U4371 (N_4371,N_3927,N_3928);
and U4372 (N_4372,In_2311,In_4028);
nor U4373 (N_4373,N_3408,N_2988);
and U4374 (N_4374,N_3669,N_3575);
nand U4375 (N_4375,N_3638,N_3674);
nand U4376 (N_4376,N_1553,N_3779);
xnor U4377 (N_4377,N_3621,N_2215);
xor U4378 (N_4378,N_3542,N_3833);
xnor U4379 (N_4379,N_3946,N_3139);
or U4380 (N_4380,N_3869,N_1933);
nor U4381 (N_4381,N_3089,N_3547);
or U4382 (N_4382,N_3679,N_2457);
or U4383 (N_4383,N_2981,N_3722);
and U4384 (N_4384,N_1952,N_3862);
xor U4385 (N_4385,N_3843,N_2103);
or U4386 (N_4386,N_3870,N_3794);
and U4387 (N_4387,N_3883,In_4937);
and U4388 (N_4388,In_2899,N_3871);
nor U4389 (N_4389,N_3045,N_3951);
xnor U4390 (N_4390,N_3240,N_3655);
or U4391 (N_4391,N_3156,In_1411);
or U4392 (N_4392,N_3731,N_3939);
or U4393 (N_4393,N_3252,N_3893);
nor U4394 (N_4394,N_2360,N_2684);
nand U4395 (N_4395,N_3664,In_3221);
or U4396 (N_4396,N_3959,N_2572);
nor U4397 (N_4397,N_3522,N_1754);
or U4398 (N_4398,N_85,N_872);
or U4399 (N_4399,N_3755,In_4660);
and U4400 (N_4400,N_3515,N_3487);
and U4401 (N_4401,N_1647,N_3875);
xnor U4402 (N_4402,N_3070,N_2570);
nor U4403 (N_4403,N_3508,N_3600);
nand U4404 (N_4404,N_3768,N_452);
nor U4405 (N_4405,N_2568,N_3983);
or U4406 (N_4406,N_3609,N_3061);
nand U4407 (N_4407,N_3949,N_3757);
nand U4408 (N_4408,N_3993,N_3646);
nand U4409 (N_4409,N_1895,N_3740);
and U4410 (N_4410,N_3332,N_3989);
or U4411 (N_4411,N_3605,N_3539);
and U4412 (N_4412,N_1504,N_2963);
or U4413 (N_4413,N_3859,N_3789);
and U4414 (N_4414,N_3817,N_1767);
and U4415 (N_4415,N_1883,N_3383);
or U4416 (N_4416,N_3633,In_2339);
and U4417 (N_4417,N_3994,N_3974);
nand U4418 (N_4418,N_3534,N_3130);
xor U4419 (N_4419,N_3695,N_3885);
xnor U4420 (N_4420,N_2852,N_3548);
nand U4421 (N_4421,N_3226,N_3364);
or U4422 (N_4422,N_3800,N_355);
or U4423 (N_4423,In_510,N_2151);
nand U4424 (N_4424,N_3712,N_3723);
or U4425 (N_4425,N_3163,N_3688);
or U4426 (N_4426,N_3576,N_3135);
nor U4427 (N_4427,N_3965,N_3333);
or U4428 (N_4428,N_3097,N_3971);
nand U4429 (N_4429,N_3882,N_3654);
xor U4430 (N_4430,N_3822,N_3844);
and U4431 (N_4431,N_1322,N_3684);
xnor U4432 (N_4432,N_3811,N_3973);
nand U4433 (N_4433,N_3892,N_1896);
xnor U4434 (N_4434,N_3556,N_3820);
nor U4435 (N_4435,N_3178,N_3940);
or U4436 (N_4436,In_59,N_3260);
nand U4437 (N_4437,N_3992,N_322);
nor U4438 (N_4438,N_978,N_3919);
nor U4439 (N_4439,N_3942,N_3396);
or U4440 (N_4440,N_3831,N_3985);
or U4441 (N_4441,N_2900,N_3349);
nand U4442 (N_4442,N_3183,N_3670);
nor U4443 (N_4443,N_3552,N_3220);
nor U4444 (N_4444,N_3936,N_2029);
or U4445 (N_4445,N_3657,N_3676);
and U4446 (N_4446,N_3777,N_3365);
nand U4447 (N_4447,N_2985,N_3331);
xnor U4448 (N_4448,N_3143,In_1409);
nand U4449 (N_4449,N_3711,N_3433);
or U4450 (N_4450,N_3782,N_3442);
nand U4451 (N_4451,N_2378,In_4686);
and U4452 (N_4452,N_3438,N_3874);
nand U4453 (N_4453,N_3415,N_3427);
nand U4454 (N_4454,N_3095,N_3753);
xor U4455 (N_4455,N_3550,N_600);
or U4456 (N_4456,N_3809,N_3825);
nand U4457 (N_4457,N_2361,N_3257);
xor U4458 (N_4458,N_2878,N_3567);
xor U4459 (N_4459,N_2665,N_3758);
and U4460 (N_4460,N_2329,N_3584);
nand U4461 (N_4461,N_3689,N_91);
nor U4462 (N_4462,N_3806,N_3956);
or U4463 (N_4463,N_3652,N_3510);
nand U4464 (N_4464,In_2591,In_3382);
nor U4465 (N_4465,In_34,N_3076);
xnor U4466 (N_4466,In_3486,N_3619);
or U4467 (N_4467,N_3569,N_2332);
or U4468 (N_4468,N_3599,N_3305);
or U4469 (N_4469,N_2968,N_3683);
or U4470 (N_4470,N_3658,N_3303);
nor U4471 (N_4471,N_3937,N_2187);
and U4472 (N_4472,N_1175,N_3890);
nand U4473 (N_4473,N_3073,N_3462);
nor U4474 (N_4474,In_1713,N_3896);
or U4475 (N_4475,N_2807,In_4885);
nor U4476 (N_4476,In_4865,N_3502);
xnor U4477 (N_4477,N_3617,N_3161);
or U4478 (N_4478,N_3769,N_3999);
or U4479 (N_4479,N_3007,N_3767);
nor U4480 (N_4480,N_3418,N_3277);
xnor U4481 (N_4481,N_3853,N_3690);
or U4482 (N_4482,N_3792,N_3543);
and U4483 (N_4483,N_3639,N_3827);
nand U4484 (N_4484,N_3998,N_3671);
or U4485 (N_4485,N_3929,N_3554);
xnor U4486 (N_4486,N_3334,N_3941);
or U4487 (N_4487,N_3762,N_3560);
xor U4488 (N_4488,N_3524,N_3611);
or U4489 (N_4489,In_3629,N_3750);
xor U4490 (N_4490,N_3930,N_2874);
or U4491 (N_4491,In_89,N_1931);
or U4492 (N_4492,N_3419,N_3544);
xnor U4493 (N_4493,N_3732,N_3744);
nor U4494 (N_4494,N_2879,N_3398);
nand U4495 (N_4495,N_3996,N_3555);
and U4496 (N_4496,N_3957,N_2616);
nand U4497 (N_4497,In_806,N_3988);
nand U4498 (N_4498,In_2500,N_1953);
or U4499 (N_4499,N_2990,In_1980);
nor U4500 (N_4500,N_4355,N_4231);
and U4501 (N_4501,N_4146,N_4173);
nor U4502 (N_4502,N_4049,N_4382);
or U4503 (N_4503,N_4140,N_4130);
or U4504 (N_4504,N_4292,N_4278);
xnor U4505 (N_4505,N_4251,N_4096);
xnor U4506 (N_4506,N_4000,N_4415);
nand U4507 (N_4507,N_4077,N_4439);
and U4508 (N_4508,N_4236,N_4396);
and U4509 (N_4509,N_4070,N_4466);
nand U4510 (N_4510,N_4248,N_4308);
and U4511 (N_4511,N_4034,N_4001);
and U4512 (N_4512,N_4452,N_4455);
or U4513 (N_4513,N_4004,N_4088);
nor U4514 (N_4514,N_4095,N_4499);
and U4515 (N_4515,N_4158,N_4317);
and U4516 (N_4516,N_4230,N_4057);
and U4517 (N_4517,N_4240,N_4329);
or U4518 (N_4518,N_4435,N_4356);
and U4519 (N_4519,N_4293,N_4234);
nand U4520 (N_4520,N_4348,N_4351);
xor U4521 (N_4521,N_4281,N_4301);
xnor U4522 (N_4522,N_4303,N_4300);
nor U4523 (N_4523,N_4109,N_4128);
xnor U4524 (N_4524,N_4144,N_4309);
or U4525 (N_4525,N_4440,N_4461);
and U4526 (N_4526,N_4105,N_4083);
nand U4527 (N_4527,N_4196,N_4101);
or U4528 (N_4528,N_4016,N_4357);
and U4529 (N_4529,N_4274,N_4084);
or U4530 (N_4530,N_4311,N_4444);
nand U4531 (N_4531,N_4022,N_4218);
nand U4532 (N_4532,N_4275,N_4165);
nor U4533 (N_4533,N_4098,N_4395);
nand U4534 (N_4534,N_4390,N_4202);
nor U4535 (N_4535,N_4087,N_4185);
or U4536 (N_4536,N_4430,N_4488);
or U4537 (N_4537,N_4447,N_4495);
nor U4538 (N_4538,N_4229,N_4262);
or U4539 (N_4539,N_4244,N_4002);
or U4540 (N_4540,N_4371,N_4012);
xnor U4541 (N_4541,N_4204,N_4368);
nor U4542 (N_4542,N_4143,N_4413);
nor U4543 (N_4543,N_4014,N_4325);
xnor U4544 (N_4544,N_4107,N_4183);
xor U4545 (N_4545,N_4349,N_4178);
xnor U4546 (N_4546,N_4347,N_4268);
nand U4547 (N_4547,N_4380,N_4160);
nand U4548 (N_4548,N_4375,N_4186);
xnor U4549 (N_4549,N_4184,N_4449);
and U4550 (N_4550,N_4392,N_4033);
and U4551 (N_4551,N_4485,N_4362);
and U4552 (N_4552,N_4135,N_4386);
xnor U4553 (N_4553,N_4214,N_4136);
nand U4554 (N_4554,N_4132,N_4172);
xnor U4555 (N_4555,N_4483,N_4490);
nand U4556 (N_4556,N_4320,N_4156);
and U4557 (N_4557,N_4476,N_4441);
nor U4558 (N_4558,N_4005,N_4114);
nand U4559 (N_4559,N_4420,N_4209);
xnor U4560 (N_4560,N_4494,N_4113);
or U4561 (N_4561,N_4225,N_4052);
xnor U4562 (N_4562,N_4051,N_4175);
and U4563 (N_4563,N_4223,N_4482);
nand U4564 (N_4564,N_4010,N_4062);
xnor U4565 (N_4565,N_4474,N_4217);
xor U4566 (N_4566,N_4145,N_4161);
and U4567 (N_4567,N_4418,N_4063);
and U4568 (N_4568,N_4133,N_4221);
nor U4569 (N_4569,N_4024,N_4264);
nand U4570 (N_4570,N_4450,N_4360);
nor U4571 (N_4571,N_4287,N_4411);
or U4572 (N_4572,N_4469,N_4359);
xor U4573 (N_4573,N_4270,N_4467);
and U4574 (N_4574,N_4048,N_4043);
nand U4575 (N_4575,N_4028,N_4445);
xnor U4576 (N_4576,N_4066,N_4417);
nor U4577 (N_4577,N_4112,N_4255);
xor U4578 (N_4578,N_4489,N_4389);
nor U4579 (N_4579,N_4331,N_4198);
nand U4580 (N_4580,N_4330,N_4342);
or U4581 (N_4581,N_4354,N_4405);
xor U4582 (N_4582,N_4493,N_4438);
nor U4583 (N_4583,N_4092,N_4341);
or U4584 (N_4584,N_4394,N_4176);
nor U4585 (N_4585,N_4369,N_4378);
nor U4586 (N_4586,N_4100,N_4310);
or U4587 (N_4587,N_4307,N_4167);
and U4588 (N_4588,N_4477,N_4023);
and U4589 (N_4589,N_4451,N_4208);
and U4590 (N_4590,N_4212,N_4094);
and U4591 (N_4591,N_4080,N_4276);
xor U4592 (N_4592,N_4280,N_4150);
nand U4593 (N_4593,N_4302,N_4038);
xnor U4594 (N_4594,N_4139,N_4243);
nor U4595 (N_4595,N_4025,N_4383);
or U4596 (N_4596,N_4104,N_4261);
xor U4597 (N_4597,N_4267,N_4199);
xnor U4598 (N_4598,N_4027,N_4367);
xnor U4599 (N_4599,N_4037,N_4409);
or U4600 (N_4600,N_4400,N_4106);
or U4601 (N_4601,N_4434,N_4045);
xnor U4602 (N_4602,N_4194,N_4102);
nand U4603 (N_4603,N_4170,N_4412);
xnor U4604 (N_4604,N_4259,N_4319);
or U4605 (N_4605,N_4366,N_4465);
xnor U4606 (N_4606,N_4304,N_4350);
xor U4607 (N_4607,N_4031,N_4436);
xor U4608 (N_4608,N_4110,N_4487);
nor U4609 (N_4609,N_4463,N_4074);
or U4610 (N_4610,N_4296,N_4117);
and U4611 (N_4611,N_4235,N_4174);
or U4612 (N_4612,N_4055,N_4182);
xnor U4613 (N_4613,N_4123,N_4336);
or U4614 (N_4614,N_4437,N_4254);
or U4615 (N_4615,N_4213,N_4408);
nor U4616 (N_4616,N_4338,N_4426);
nand U4617 (N_4617,N_4076,N_4059);
and U4618 (N_4618,N_4053,N_4364);
nor U4619 (N_4619,N_4042,N_4006);
nand U4620 (N_4620,N_4191,N_4265);
xnor U4621 (N_4621,N_4376,N_4335);
nand U4622 (N_4622,N_4228,N_4155);
nor U4623 (N_4623,N_4298,N_4171);
or U4624 (N_4624,N_4353,N_4361);
nand U4625 (N_4625,N_4036,N_4305);
nand U4626 (N_4626,N_4423,N_4456);
and U4627 (N_4627,N_4233,N_4099);
nor U4628 (N_4628,N_4397,N_4385);
nand U4629 (N_4629,N_4011,N_4147);
and U4630 (N_4630,N_4428,N_4203);
nand U4631 (N_4631,N_4166,N_4344);
nor U4632 (N_4632,N_4232,N_4021);
and U4633 (N_4633,N_4370,N_4097);
nor U4634 (N_4634,N_4306,N_4442);
or U4635 (N_4635,N_4443,N_4374);
nor U4636 (N_4636,N_4239,N_4398);
nand U4637 (N_4637,N_4219,N_4237);
nor U4638 (N_4638,N_4480,N_4065);
and U4639 (N_4639,N_4425,N_4497);
xnor U4640 (N_4640,N_4041,N_4082);
nor U4641 (N_4641,N_4315,N_4326);
nand U4642 (N_4642,N_4157,N_4283);
and U4643 (N_4643,N_4189,N_4111);
or U4644 (N_4644,N_4127,N_4468);
nor U4645 (N_4645,N_4269,N_4013);
nor U4646 (N_4646,N_4072,N_4168);
xnor U4647 (N_4647,N_4210,N_4471);
or U4648 (N_4648,N_4035,N_4419);
and U4649 (N_4649,N_4365,N_4312);
and U4650 (N_4650,N_4009,N_4256);
xor U4651 (N_4651,N_4294,N_4498);
xor U4652 (N_4652,N_4429,N_4388);
nor U4653 (N_4653,N_4472,N_4192);
and U4654 (N_4654,N_4093,N_4299);
xor U4655 (N_4655,N_4484,N_4081);
and U4656 (N_4656,N_4163,N_4020);
nor U4657 (N_4657,N_4180,N_4491);
or U4658 (N_4658,N_4138,N_4462);
nor U4659 (N_4659,N_4148,N_4121);
and U4660 (N_4660,N_4401,N_4324);
or U4661 (N_4661,N_4431,N_4116);
and U4662 (N_4662,N_4416,N_4432);
nand U4663 (N_4663,N_4071,N_4164);
xnor U4664 (N_4664,N_4029,N_4181);
nand U4665 (N_4665,N_4205,N_4075);
nor U4666 (N_4666,N_4289,N_4047);
or U4667 (N_4667,N_4050,N_4263);
nand U4668 (N_4668,N_4407,N_4448);
nor U4669 (N_4669,N_4177,N_4060);
nand U4670 (N_4670,N_4067,N_4241);
xor U4671 (N_4671,N_4187,N_4424);
or U4672 (N_4672,N_4279,N_4115);
or U4673 (N_4673,N_4124,N_4188);
and U4674 (N_4674,N_4478,N_4297);
and U4675 (N_4675,N_4141,N_4242);
and U4676 (N_4676,N_4046,N_4152);
and U4677 (N_4677,N_4222,N_4085);
and U4678 (N_4678,N_4019,N_4126);
nor U4679 (N_4679,N_4272,N_4260);
or U4680 (N_4680,N_4220,N_4340);
nand U4681 (N_4681,N_4108,N_4216);
nand U4682 (N_4682,N_4149,N_4040);
or U4683 (N_4683,N_4201,N_4404);
nand U4684 (N_4684,N_4288,N_4227);
or U4685 (N_4685,N_4266,N_4313);
or U4686 (N_4686,N_4457,N_4142);
and U4687 (N_4687,N_4026,N_4381);
xnor U4688 (N_4688,N_4334,N_4427);
or U4689 (N_4689,N_4496,N_4403);
nor U4690 (N_4690,N_4197,N_4323);
and U4691 (N_4691,N_4337,N_4103);
nor U4692 (N_4692,N_4079,N_4179);
nor U4693 (N_4693,N_4018,N_4257);
or U4694 (N_4694,N_4134,N_4078);
or U4695 (N_4695,N_4492,N_4193);
nor U4696 (N_4696,N_4460,N_4414);
xnor U4697 (N_4697,N_4479,N_4154);
nor U4698 (N_4698,N_4089,N_4162);
and U4699 (N_4699,N_4481,N_4246);
nand U4700 (N_4700,N_4131,N_4007);
nor U4701 (N_4701,N_4250,N_4091);
nor U4702 (N_4702,N_4318,N_4332);
nand U4703 (N_4703,N_4295,N_4486);
xor U4704 (N_4704,N_4433,N_4327);
xnor U4705 (N_4705,N_4195,N_4137);
and U4706 (N_4706,N_4410,N_4273);
or U4707 (N_4707,N_4316,N_4151);
nor U4708 (N_4708,N_4238,N_4122);
and U4709 (N_4709,N_4008,N_4384);
nand U4710 (N_4710,N_4387,N_4379);
or U4711 (N_4711,N_4215,N_4169);
xor U4712 (N_4712,N_4352,N_4343);
and U4713 (N_4713,N_4258,N_4190);
nand U4714 (N_4714,N_4271,N_4345);
nand U4715 (N_4715,N_4321,N_4284);
nand U4716 (N_4716,N_4090,N_4086);
xnor U4717 (N_4717,N_4453,N_4030);
and U4718 (N_4718,N_4118,N_4039);
nor U4719 (N_4719,N_4373,N_4333);
or U4720 (N_4720,N_4458,N_4363);
or U4721 (N_4721,N_4346,N_4286);
and U4722 (N_4722,N_4358,N_4282);
nand U4723 (N_4723,N_4393,N_4056);
nand U4724 (N_4724,N_4245,N_4399);
or U4725 (N_4725,N_4470,N_4224);
and U4726 (N_4726,N_4119,N_4206);
nor U4727 (N_4727,N_4247,N_4054);
nand U4728 (N_4728,N_4068,N_4249);
xnor U4729 (N_4729,N_4129,N_4153);
or U4730 (N_4730,N_4475,N_4015);
or U4731 (N_4731,N_4125,N_4322);
and U4732 (N_4732,N_4120,N_4459);
nor U4733 (N_4733,N_4290,N_4391);
and U4734 (N_4734,N_4226,N_4314);
xnor U4735 (N_4735,N_4044,N_4207);
nor U4736 (N_4736,N_4372,N_4339);
nand U4737 (N_4737,N_4446,N_4058);
or U4738 (N_4738,N_4422,N_4211);
and U4739 (N_4739,N_4377,N_4253);
nand U4740 (N_4740,N_4402,N_4454);
and U4741 (N_4741,N_4285,N_4032);
and U4742 (N_4742,N_4328,N_4003);
or U4743 (N_4743,N_4159,N_4473);
nand U4744 (N_4744,N_4421,N_4073);
xor U4745 (N_4745,N_4291,N_4252);
nand U4746 (N_4746,N_4406,N_4200);
nor U4747 (N_4747,N_4017,N_4069);
and U4748 (N_4748,N_4061,N_4064);
and U4749 (N_4749,N_4277,N_4464);
or U4750 (N_4750,N_4387,N_4183);
nand U4751 (N_4751,N_4234,N_4452);
and U4752 (N_4752,N_4136,N_4147);
nand U4753 (N_4753,N_4181,N_4457);
xnor U4754 (N_4754,N_4477,N_4268);
nand U4755 (N_4755,N_4143,N_4103);
xnor U4756 (N_4756,N_4295,N_4332);
nor U4757 (N_4757,N_4429,N_4325);
xor U4758 (N_4758,N_4334,N_4401);
and U4759 (N_4759,N_4000,N_4293);
and U4760 (N_4760,N_4041,N_4179);
nor U4761 (N_4761,N_4357,N_4301);
or U4762 (N_4762,N_4307,N_4255);
nand U4763 (N_4763,N_4423,N_4218);
nand U4764 (N_4764,N_4461,N_4218);
or U4765 (N_4765,N_4199,N_4495);
nor U4766 (N_4766,N_4420,N_4078);
nor U4767 (N_4767,N_4326,N_4043);
and U4768 (N_4768,N_4184,N_4332);
and U4769 (N_4769,N_4129,N_4096);
or U4770 (N_4770,N_4072,N_4408);
and U4771 (N_4771,N_4446,N_4303);
xor U4772 (N_4772,N_4435,N_4013);
or U4773 (N_4773,N_4352,N_4353);
xor U4774 (N_4774,N_4419,N_4370);
and U4775 (N_4775,N_4455,N_4157);
and U4776 (N_4776,N_4038,N_4254);
and U4777 (N_4777,N_4338,N_4441);
nor U4778 (N_4778,N_4486,N_4355);
nor U4779 (N_4779,N_4471,N_4085);
nand U4780 (N_4780,N_4329,N_4048);
nand U4781 (N_4781,N_4479,N_4280);
and U4782 (N_4782,N_4429,N_4370);
and U4783 (N_4783,N_4244,N_4476);
xor U4784 (N_4784,N_4003,N_4445);
or U4785 (N_4785,N_4337,N_4307);
nand U4786 (N_4786,N_4003,N_4433);
nor U4787 (N_4787,N_4084,N_4153);
and U4788 (N_4788,N_4329,N_4146);
nor U4789 (N_4789,N_4032,N_4147);
xnor U4790 (N_4790,N_4084,N_4444);
xnor U4791 (N_4791,N_4293,N_4009);
xnor U4792 (N_4792,N_4086,N_4103);
or U4793 (N_4793,N_4499,N_4305);
or U4794 (N_4794,N_4080,N_4327);
nand U4795 (N_4795,N_4043,N_4437);
nand U4796 (N_4796,N_4008,N_4245);
nor U4797 (N_4797,N_4173,N_4298);
or U4798 (N_4798,N_4419,N_4039);
and U4799 (N_4799,N_4289,N_4074);
xnor U4800 (N_4800,N_4190,N_4202);
or U4801 (N_4801,N_4040,N_4135);
nand U4802 (N_4802,N_4255,N_4319);
and U4803 (N_4803,N_4347,N_4458);
nand U4804 (N_4804,N_4001,N_4259);
and U4805 (N_4805,N_4165,N_4250);
xnor U4806 (N_4806,N_4192,N_4009);
and U4807 (N_4807,N_4124,N_4223);
nand U4808 (N_4808,N_4169,N_4402);
or U4809 (N_4809,N_4410,N_4029);
nand U4810 (N_4810,N_4162,N_4462);
and U4811 (N_4811,N_4135,N_4100);
and U4812 (N_4812,N_4373,N_4449);
or U4813 (N_4813,N_4000,N_4385);
nor U4814 (N_4814,N_4022,N_4255);
nand U4815 (N_4815,N_4385,N_4178);
nand U4816 (N_4816,N_4328,N_4267);
xnor U4817 (N_4817,N_4251,N_4209);
or U4818 (N_4818,N_4050,N_4000);
xnor U4819 (N_4819,N_4408,N_4059);
and U4820 (N_4820,N_4055,N_4038);
xor U4821 (N_4821,N_4015,N_4322);
xor U4822 (N_4822,N_4156,N_4474);
xnor U4823 (N_4823,N_4121,N_4286);
or U4824 (N_4824,N_4169,N_4475);
or U4825 (N_4825,N_4005,N_4199);
xor U4826 (N_4826,N_4417,N_4324);
nand U4827 (N_4827,N_4454,N_4446);
nor U4828 (N_4828,N_4244,N_4246);
and U4829 (N_4829,N_4061,N_4274);
and U4830 (N_4830,N_4486,N_4285);
and U4831 (N_4831,N_4412,N_4384);
nand U4832 (N_4832,N_4379,N_4292);
and U4833 (N_4833,N_4202,N_4463);
and U4834 (N_4834,N_4411,N_4470);
or U4835 (N_4835,N_4103,N_4034);
xnor U4836 (N_4836,N_4326,N_4169);
or U4837 (N_4837,N_4110,N_4305);
and U4838 (N_4838,N_4052,N_4315);
nand U4839 (N_4839,N_4124,N_4299);
or U4840 (N_4840,N_4237,N_4313);
nand U4841 (N_4841,N_4261,N_4200);
nor U4842 (N_4842,N_4398,N_4309);
nor U4843 (N_4843,N_4013,N_4477);
xor U4844 (N_4844,N_4006,N_4382);
and U4845 (N_4845,N_4072,N_4415);
and U4846 (N_4846,N_4087,N_4041);
and U4847 (N_4847,N_4179,N_4131);
nor U4848 (N_4848,N_4203,N_4232);
xnor U4849 (N_4849,N_4453,N_4447);
nor U4850 (N_4850,N_4460,N_4254);
nand U4851 (N_4851,N_4187,N_4284);
nor U4852 (N_4852,N_4311,N_4194);
or U4853 (N_4853,N_4161,N_4286);
and U4854 (N_4854,N_4160,N_4114);
and U4855 (N_4855,N_4452,N_4174);
and U4856 (N_4856,N_4275,N_4193);
nand U4857 (N_4857,N_4103,N_4033);
nor U4858 (N_4858,N_4233,N_4199);
nor U4859 (N_4859,N_4120,N_4069);
or U4860 (N_4860,N_4299,N_4083);
or U4861 (N_4861,N_4277,N_4123);
and U4862 (N_4862,N_4165,N_4480);
or U4863 (N_4863,N_4348,N_4189);
and U4864 (N_4864,N_4231,N_4488);
and U4865 (N_4865,N_4340,N_4219);
and U4866 (N_4866,N_4030,N_4184);
or U4867 (N_4867,N_4492,N_4050);
or U4868 (N_4868,N_4280,N_4214);
and U4869 (N_4869,N_4129,N_4289);
or U4870 (N_4870,N_4327,N_4243);
nor U4871 (N_4871,N_4405,N_4389);
and U4872 (N_4872,N_4464,N_4146);
nand U4873 (N_4873,N_4106,N_4139);
and U4874 (N_4874,N_4077,N_4323);
xnor U4875 (N_4875,N_4354,N_4045);
nand U4876 (N_4876,N_4423,N_4412);
xor U4877 (N_4877,N_4337,N_4114);
or U4878 (N_4878,N_4410,N_4452);
nand U4879 (N_4879,N_4078,N_4486);
nor U4880 (N_4880,N_4127,N_4084);
xnor U4881 (N_4881,N_4117,N_4002);
nor U4882 (N_4882,N_4177,N_4220);
and U4883 (N_4883,N_4224,N_4079);
nand U4884 (N_4884,N_4126,N_4266);
nand U4885 (N_4885,N_4256,N_4261);
nor U4886 (N_4886,N_4184,N_4200);
xnor U4887 (N_4887,N_4383,N_4167);
nand U4888 (N_4888,N_4427,N_4441);
and U4889 (N_4889,N_4003,N_4289);
nand U4890 (N_4890,N_4471,N_4176);
nand U4891 (N_4891,N_4133,N_4322);
xor U4892 (N_4892,N_4154,N_4183);
nand U4893 (N_4893,N_4465,N_4263);
nand U4894 (N_4894,N_4133,N_4188);
xnor U4895 (N_4895,N_4356,N_4041);
and U4896 (N_4896,N_4403,N_4239);
nor U4897 (N_4897,N_4366,N_4499);
and U4898 (N_4898,N_4387,N_4369);
and U4899 (N_4899,N_4025,N_4330);
nor U4900 (N_4900,N_4036,N_4406);
nand U4901 (N_4901,N_4023,N_4240);
and U4902 (N_4902,N_4152,N_4388);
nand U4903 (N_4903,N_4395,N_4431);
or U4904 (N_4904,N_4194,N_4408);
and U4905 (N_4905,N_4122,N_4153);
nand U4906 (N_4906,N_4142,N_4118);
and U4907 (N_4907,N_4484,N_4417);
and U4908 (N_4908,N_4479,N_4157);
or U4909 (N_4909,N_4312,N_4264);
or U4910 (N_4910,N_4005,N_4034);
nand U4911 (N_4911,N_4100,N_4032);
nand U4912 (N_4912,N_4241,N_4063);
and U4913 (N_4913,N_4468,N_4359);
xor U4914 (N_4914,N_4135,N_4185);
nand U4915 (N_4915,N_4197,N_4403);
and U4916 (N_4916,N_4126,N_4223);
nand U4917 (N_4917,N_4019,N_4321);
xor U4918 (N_4918,N_4196,N_4461);
or U4919 (N_4919,N_4345,N_4259);
and U4920 (N_4920,N_4357,N_4265);
and U4921 (N_4921,N_4247,N_4366);
xnor U4922 (N_4922,N_4076,N_4088);
nor U4923 (N_4923,N_4281,N_4231);
or U4924 (N_4924,N_4460,N_4488);
nor U4925 (N_4925,N_4397,N_4218);
nor U4926 (N_4926,N_4047,N_4422);
nand U4927 (N_4927,N_4427,N_4347);
and U4928 (N_4928,N_4345,N_4184);
or U4929 (N_4929,N_4352,N_4335);
or U4930 (N_4930,N_4332,N_4400);
and U4931 (N_4931,N_4438,N_4265);
and U4932 (N_4932,N_4128,N_4011);
and U4933 (N_4933,N_4307,N_4037);
xnor U4934 (N_4934,N_4272,N_4487);
and U4935 (N_4935,N_4343,N_4482);
nand U4936 (N_4936,N_4474,N_4171);
or U4937 (N_4937,N_4427,N_4326);
nand U4938 (N_4938,N_4070,N_4136);
nor U4939 (N_4939,N_4147,N_4018);
or U4940 (N_4940,N_4008,N_4227);
and U4941 (N_4941,N_4305,N_4227);
nand U4942 (N_4942,N_4138,N_4400);
and U4943 (N_4943,N_4444,N_4392);
xnor U4944 (N_4944,N_4274,N_4123);
xnor U4945 (N_4945,N_4182,N_4072);
or U4946 (N_4946,N_4282,N_4453);
nand U4947 (N_4947,N_4035,N_4131);
nor U4948 (N_4948,N_4267,N_4182);
xnor U4949 (N_4949,N_4224,N_4149);
or U4950 (N_4950,N_4131,N_4458);
nor U4951 (N_4951,N_4309,N_4027);
or U4952 (N_4952,N_4094,N_4130);
and U4953 (N_4953,N_4084,N_4314);
and U4954 (N_4954,N_4301,N_4344);
xor U4955 (N_4955,N_4391,N_4490);
nand U4956 (N_4956,N_4415,N_4195);
nand U4957 (N_4957,N_4268,N_4376);
nand U4958 (N_4958,N_4357,N_4146);
and U4959 (N_4959,N_4017,N_4133);
and U4960 (N_4960,N_4393,N_4430);
nor U4961 (N_4961,N_4221,N_4140);
nand U4962 (N_4962,N_4230,N_4045);
nand U4963 (N_4963,N_4112,N_4012);
nor U4964 (N_4964,N_4350,N_4302);
nand U4965 (N_4965,N_4327,N_4118);
or U4966 (N_4966,N_4338,N_4180);
nor U4967 (N_4967,N_4147,N_4092);
xor U4968 (N_4968,N_4075,N_4412);
nand U4969 (N_4969,N_4199,N_4463);
xnor U4970 (N_4970,N_4447,N_4352);
nor U4971 (N_4971,N_4137,N_4225);
xor U4972 (N_4972,N_4320,N_4035);
nand U4973 (N_4973,N_4360,N_4371);
nor U4974 (N_4974,N_4455,N_4426);
and U4975 (N_4975,N_4023,N_4403);
and U4976 (N_4976,N_4220,N_4178);
or U4977 (N_4977,N_4061,N_4469);
xor U4978 (N_4978,N_4196,N_4091);
nand U4979 (N_4979,N_4241,N_4385);
and U4980 (N_4980,N_4300,N_4271);
or U4981 (N_4981,N_4134,N_4434);
nor U4982 (N_4982,N_4325,N_4240);
or U4983 (N_4983,N_4402,N_4475);
nand U4984 (N_4984,N_4296,N_4429);
nand U4985 (N_4985,N_4478,N_4471);
nand U4986 (N_4986,N_4399,N_4118);
nor U4987 (N_4987,N_4432,N_4206);
xnor U4988 (N_4988,N_4359,N_4128);
or U4989 (N_4989,N_4294,N_4086);
nand U4990 (N_4990,N_4319,N_4155);
or U4991 (N_4991,N_4389,N_4249);
and U4992 (N_4992,N_4484,N_4063);
nand U4993 (N_4993,N_4098,N_4277);
nor U4994 (N_4994,N_4373,N_4196);
and U4995 (N_4995,N_4191,N_4226);
and U4996 (N_4996,N_4190,N_4252);
nor U4997 (N_4997,N_4452,N_4040);
nand U4998 (N_4998,N_4114,N_4120);
xnor U4999 (N_4999,N_4263,N_4106);
nor U5000 (N_5000,N_4708,N_4871);
nand U5001 (N_5001,N_4998,N_4875);
nand U5002 (N_5002,N_4901,N_4851);
nor U5003 (N_5003,N_4528,N_4833);
nand U5004 (N_5004,N_4870,N_4687);
or U5005 (N_5005,N_4644,N_4521);
nand U5006 (N_5006,N_4817,N_4936);
nor U5007 (N_5007,N_4795,N_4966);
xnor U5008 (N_5008,N_4918,N_4762);
nand U5009 (N_5009,N_4682,N_4945);
or U5010 (N_5010,N_4948,N_4745);
nand U5011 (N_5011,N_4533,N_4712);
nor U5012 (N_5012,N_4897,N_4661);
nor U5013 (N_5013,N_4520,N_4699);
or U5014 (N_5014,N_4578,N_4916);
and U5015 (N_5015,N_4738,N_4880);
or U5016 (N_5016,N_4927,N_4911);
nand U5017 (N_5017,N_4696,N_4786);
or U5018 (N_5018,N_4859,N_4991);
and U5019 (N_5019,N_4548,N_4526);
and U5020 (N_5020,N_4685,N_4693);
and U5021 (N_5021,N_4804,N_4669);
and U5022 (N_5022,N_4743,N_4524);
nor U5023 (N_5023,N_4912,N_4813);
xor U5024 (N_5024,N_4536,N_4710);
xnor U5025 (N_5025,N_4836,N_4519);
nand U5026 (N_5026,N_4860,N_4941);
and U5027 (N_5027,N_4826,N_4718);
xnor U5028 (N_5028,N_4955,N_4959);
nor U5029 (N_5029,N_4976,N_4765);
nor U5030 (N_5030,N_4660,N_4512);
and U5031 (N_5031,N_4575,N_4891);
and U5032 (N_5032,N_4540,N_4585);
xnor U5033 (N_5033,N_4717,N_4613);
nor U5034 (N_5034,N_4665,N_4729);
and U5035 (N_5035,N_4815,N_4734);
and U5036 (N_5036,N_4985,N_4968);
nor U5037 (N_5037,N_4632,N_4970);
xor U5038 (N_5038,N_4603,N_4705);
or U5039 (N_5039,N_4652,N_4720);
nand U5040 (N_5040,N_4760,N_4997);
or U5041 (N_5041,N_4781,N_4510);
nor U5042 (N_5042,N_4986,N_4645);
nand U5043 (N_5043,N_4648,N_4910);
or U5044 (N_5044,N_4576,N_4647);
xor U5045 (N_5045,N_4843,N_4742);
nor U5046 (N_5046,N_4516,N_4971);
nor U5047 (N_5047,N_4772,N_4549);
nand U5048 (N_5048,N_4925,N_4964);
and U5049 (N_5049,N_4572,N_4597);
nor U5050 (N_5050,N_4675,N_4819);
nand U5051 (N_5051,N_4539,N_4563);
nand U5052 (N_5052,N_4898,N_4704);
nor U5053 (N_5053,N_4820,N_4562);
nand U5054 (N_5054,N_4967,N_4621);
xnor U5055 (N_5055,N_4957,N_4917);
nor U5056 (N_5056,N_4601,N_4878);
nand U5057 (N_5057,N_4668,N_4796);
nand U5058 (N_5058,N_4513,N_4502);
or U5059 (N_5059,N_4748,N_4777);
and U5060 (N_5060,N_4972,N_4617);
and U5061 (N_5061,N_4564,N_4611);
nor U5062 (N_5062,N_4546,N_4756);
nor U5063 (N_5063,N_4733,N_4679);
or U5064 (N_5064,N_4994,N_4628);
or U5065 (N_5065,N_4749,N_4853);
and U5066 (N_5066,N_4622,N_4571);
and U5067 (N_5067,N_4906,N_4580);
xor U5068 (N_5068,N_4943,N_4773);
or U5069 (N_5069,N_4690,N_4792);
nor U5070 (N_5070,N_4633,N_4584);
or U5071 (N_5071,N_4863,N_4755);
and U5072 (N_5072,N_4747,N_4653);
and U5073 (N_5073,N_4716,N_4514);
and U5074 (N_5074,N_4594,N_4893);
nor U5075 (N_5075,N_4861,N_4629);
xor U5076 (N_5076,N_4583,N_4662);
nand U5077 (N_5077,N_4636,N_4511);
and U5078 (N_5078,N_4935,N_4907);
nand U5079 (N_5079,N_4686,N_4832);
nor U5080 (N_5080,N_4958,N_4737);
and U5081 (N_5081,N_4806,N_4530);
or U5082 (N_5082,N_4922,N_4780);
xnor U5083 (N_5083,N_4680,N_4504);
nor U5084 (N_5084,N_4518,N_4915);
xor U5085 (N_5085,N_4625,N_4586);
and U5086 (N_5086,N_4827,N_4894);
xnor U5087 (N_5087,N_4837,N_4515);
or U5088 (N_5088,N_4552,N_4570);
nand U5089 (N_5089,N_4558,N_4574);
or U5090 (N_5090,N_4608,N_4609);
nand U5091 (N_5091,N_4766,N_4788);
nand U5092 (N_5092,N_4544,N_4759);
or U5093 (N_5093,N_4973,N_4924);
and U5094 (N_5094,N_4944,N_4803);
and U5095 (N_5095,N_4757,N_4569);
nand U5096 (N_5096,N_4637,N_4650);
xnor U5097 (N_5097,N_4542,N_4744);
nand U5098 (N_5098,N_4855,N_4933);
nand U5099 (N_5099,N_4844,N_4754);
and U5100 (N_5100,N_4579,N_4509);
nand U5101 (N_5101,N_4534,N_4869);
and U5102 (N_5102,N_4726,N_4954);
or U5103 (N_5103,N_4960,N_4663);
or U5104 (N_5104,N_4550,N_4776);
and U5105 (N_5105,N_4876,N_4920);
or U5106 (N_5106,N_4599,N_4684);
nor U5107 (N_5107,N_4874,N_4545);
nand U5108 (N_5108,N_4522,N_4980);
nor U5109 (N_5109,N_4787,N_4649);
nand U5110 (N_5110,N_4565,N_4646);
xor U5111 (N_5111,N_4501,N_4969);
nand U5112 (N_5112,N_4989,N_4721);
and U5113 (N_5113,N_4557,N_4677);
nor U5114 (N_5114,N_4556,N_4824);
nand U5115 (N_5115,N_4990,N_4658);
nor U5116 (N_5116,N_4840,N_4672);
nand U5117 (N_5117,N_4779,N_4821);
xnor U5118 (N_5118,N_4950,N_4707);
or U5119 (N_5119,N_4854,N_4688);
or U5120 (N_5120,N_4949,N_4541);
and U5121 (N_5121,N_4651,N_4730);
and U5122 (N_5122,N_4926,N_4600);
and U5123 (N_5123,N_4790,N_4838);
xor U5124 (N_5124,N_4931,N_4961);
or U5125 (N_5125,N_4940,N_4816);
nor U5126 (N_5126,N_4602,N_4805);
and U5127 (N_5127,N_4883,N_4914);
xor U5128 (N_5128,N_4885,N_4929);
xor U5129 (N_5129,N_4753,N_4532);
nand U5130 (N_5130,N_4605,N_4877);
and U5131 (N_5131,N_4698,N_4610);
or U5132 (N_5132,N_4593,N_4939);
xor U5133 (N_5133,N_4866,N_4631);
xnor U5134 (N_5134,N_4951,N_4567);
nand U5135 (N_5135,N_4828,N_4769);
nand U5136 (N_5136,N_4626,N_4896);
nor U5137 (N_5137,N_4607,N_4835);
and U5138 (N_5138,N_4823,N_4538);
xnor U5139 (N_5139,N_4992,N_4864);
xnor U5140 (N_5140,N_4616,N_4592);
or U5141 (N_5141,N_4624,N_4659);
or U5142 (N_5142,N_4751,N_4825);
xnor U5143 (N_5143,N_4879,N_4736);
and U5144 (N_5144,N_4887,N_4785);
and U5145 (N_5145,N_4767,N_4867);
nor U5146 (N_5146,N_4890,N_4500);
or U5147 (N_5147,N_4674,N_4666);
xnor U5148 (N_5148,N_4523,N_4770);
or U5149 (N_5149,N_4689,N_4553);
nor U5150 (N_5150,N_4664,N_4681);
xnor U5151 (N_5151,N_4711,N_4995);
nand U5152 (N_5152,N_4850,N_4993);
nor U5153 (N_5153,N_4678,N_4793);
and U5154 (N_5154,N_4507,N_4642);
or U5155 (N_5155,N_4531,N_4547);
and U5156 (N_5156,N_4761,N_4620);
or U5157 (N_5157,N_4899,N_4517);
xor U5158 (N_5158,N_4789,N_4892);
or U5159 (N_5159,N_4978,N_4627);
or U5160 (N_5160,N_4981,N_4846);
nand U5161 (N_5161,N_4845,N_4728);
nand U5162 (N_5162,N_4731,N_4640);
nand U5163 (N_5163,N_4799,N_4857);
or U5164 (N_5164,N_4551,N_4529);
xnor U5165 (N_5165,N_4582,N_4695);
nor U5166 (N_5166,N_4655,N_4947);
and U5167 (N_5167,N_4831,N_4975);
nand U5168 (N_5168,N_4938,N_4559);
or U5169 (N_5169,N_4700,N_4612);
and U5170 (N_5170,N_4618,N_4987);
nand U5171 (N_5171,N_4566,N_4984);
nor U5172 (N_5172,N_4604,N_4800);
nor U5173 (N_5173,N_4982,N_4709);
nand U5174 (N_5174,N_4818,N_4715);
nor U5175 (N_5175,N_4872,N_4886);
xnor U5176 (N_5176,N_4849,N_4527);
and U5177 (N_5177,N_4508,N_4812);
nor U5178 (N_5178,N_4525,N_4810);
xnor U5179 (N_5179,N_4930,N_4937);
xor U5180 (N_5180,N_4724,N_4921);
or U5181 (N_5181,N_4581,N_4573);
nand U5182 (N_5182,N_4641,N_4903);
or U5183 (N_5183,N_4758,N_4746);
xnor U5184 (N_5184,N_4862,N_4798);
nor U5185 (N_5185,N_4829,N_4671);
xor U5186 (N_5186,N_4895,N_4676);
and U5187 (N_5187,N_4928,N_4657);
xor U5188 (N_5188,N_4701,N_4889);
nor U5189 (N_5189,N_4596,N_4555);
xor U5190 (N_5190,N_4673,N_4847);
nand U5191 (N_5191,N_4983,N_4577);
xor U5192 (N_5192,N_4900,N_4590);
nor U5193 (N_5193,N_4725,N_4830);
and U5194 (N_5194,N_4852,N_4839);
nor U5195 (N_5195,N_4784,N_4909);
nand U5196 (N_5196,N_4735,N_4768);
and U5197 (N_5197,N_4667,N_4763);
and U5198 (N_5198,N_4723,N_4750);
nor U5199 (N_5199,N_4764,N_4808);
nand U5200 (N_5200,N_4953,N_4741);
or U5201 (N_5201,N_4811,N_4619);
or U5202 (N_5202,N_4719,N_4554);
xor U5203 (N_5203,N_4999,N_4630);
nand U5204 (N_5204,N_4979,N_4834);
nor U5205 (N_5205,N_4739,N_4797);
and U5206 (N_5206,N_4974,N_4904);
nand U5207 (N_5207,N_4882,N_4683);
nor U5208 (N_5208,N_4595,N_4606);
and U5209 (N_5209,N_4656,N_4848);
nor U5210 (N_5210,N_4615,N_4740);
xor U5211 (N_5211,N_4561,N_4752);
xnor U5212 (N_5212,N_4856,N_4560);
xnor U5213 (N_5213,N_4694,N_4635);
and U5214 (N_5214,N_4868,N_4775);
or U5215 (N_5215,N_4822,N_4952);
and U5216 (N_5216,N_4670,N_4703);
and U5217 (N_5217,N_4774,N_4919);
xor U5218 (N_5218,N_4691,N_4842);
nor U5219 (N_5219,N_4732,N_4702);
nor U5220 (N_5220,N_4801,N_4807);
and U5221 (N_5221,N_4962,N_4722);
and U5222 (N_5222,N_4506,N_4598);
and U5223 (N_5223,N_4923,N_4873);
nor U5224 (N_5224,N_4503,N_4913);
xnor U5225 (N_5225,N_4639,N_4587);
xnor U5226 (N_5226,N_4505,N_4946);
nand U5227 (N_5227,N_4932,N_4908);
nand U5228 (N_5228,N_4589,N_4543);
or U5229 (N_5229,N_4942,N_4634);
nor U5230 (N_5230,N_4888,N_4714);
nor U5231 (N_5231,N_4614,N_4697);
nor U5232 (N_5232,N_4588,N_4841);
nor U5233 (N_5233,N_4881,N_4623);
nand U5234 (N_5234,N_4643,N_4865);
nor U5235 (N_5235,N_4783,N_4568);
and U5236 (N_5236,N_4791,N_4727);
nand U5237 (N_5237,N_4713,N_4934);
or U5238 (N_5238,N_4809,N_4794);
xnor U5239 (N_5239,N_4905,N_4858);
xnor U5240 (N_5240,N_4771,N_4537);
nand U5241 (N_5241,N_4884,N_4988);
and U5242 (N_5242,N_4591,N_4814);
xor U5243 (N_5243,N_4654,N_4778);
nand U5244 (N_5244,N_4902,N_4963);
nor U5245 (N_5245,N_4638,N_4535);
or U5246 (N_5246,N_4977,N_4692);
and U5247 (N_5247,N_4965,N_4706);
xnor U5248 (N_5248,N_4996,N_4782);
and U5249 (N_5249,N_4802,N_4956);
and U5250 (N_5250,N_4911,N_4972);
nor U5251 (N_5251,N_4832,N_4661);
nand U5252 (N_5252,N_4776,N_4908);
nand U5253 (N_5253,N_4890,N_4549);
nand U5254 (N_5254,N_4821,N_4537);
xor U5255 (N_5255,N_4858,N_4586);
nand U5256 (N_5256,N_4951,N_4502);
xor U5257 (N_5257,N_4638,N_4846);
xor U5258 (N_5258,N_4666,N_4760);
xor U5259 (N_5259,N_4933,N_4866);
nor U5260 (N_5260,N_4745,N_4552);
xor U5261 (N_5261,N_4599,N_4899);
and U5262 (N_5262,N_4797,N_4790);
nor U5263 (N_5263,N_4650,N_4535);
or U5264 (N_5264,N_4927,N_4747);
nand U5265 (N_5265,N_4822,N_4597);
or U5266 (N_5266,N_4757,N_4517);
nand U5267 (N_5267,N_4784,N_4718);
xnor U5268 (N_5268,N_4789,N_4611);
and U5269 (N_5269,N_4987,N_4686);
xnor U5270 (N_5270,N_4786,N_4651);
xor U5271 (N_5271,N_4831,N_4742);
nor U5272 (N_5272,N_4887,N_4587);
nor U5273 (N_5273,N_4823,N_4835);
or U5274 (N_5274,N_4758,N_4876);
or U5275 (N_5275,N_4794,N_4709);
nor U5276 (N_5276,N_4597,N_4979);
or U5277 (N_5277,N_4836,N_4611);
or U5278 (N_5278,N_4787,N_4770);
and U5279 (N_5279,N_4532,N_4932);
nor U5280 (N_5280,N_4740,N_4570);
nand U5281 (N_5281,N_4962,N_4557);
xor U5282 (N_5282,N_4934,N_4682);
nand U5283 (N_5283,N_4566,N_4729);
or U5284 (N_5284,N_4594,N_4661);
nand U5285 (N_5285,N_4941,N_4504);
nand U5286 (N_5286,N_4800,N_4825);
xor U5287 (N_5287,N_4738,N_4896);
nor U5288 (N_5288,N_4666,N_4724);
xnor U5289 (N_5289,N_4638,N_4863);
and U5290 (N_5290,N_4965,N_4902);
nand U5291 (N_5291,N_4842,N_4626);
xnor U5292 (N_5292,N_4852,N_4729);
xnor U5293 (N_5293,N_4976,N_4806);
nand U5294 (N_5294,N_4741,N_4598);
and U5295 (N_5295,N_4514,N_4776);
nand U5296 (N_5296,N_4821,N_4923);
nand U5297 (N_5297,N_4981,N_4639);
xor U5298 (N_5298,N_4777,N_4728);
nand U5299 (N_5299,N_4618,N_4963);
or U5300 (N_5300,N_4986,N_4501);
and U5301 (N_5301,N_4580,N_4554);
xnor U5302 (N_5302,N_4941,N_4789);
and U5303 (N_5303,N_4523,N_4521);
nor U5304 (N_5304,N_4803,N_4521);
or U5305 (N_5305,N_4583,N_4504);
nor U5306 (N_5306,N_4903,N_4517);
xnor U5307 (N_5307,N_4600,N_4997);
nand U5308 (N_5308,N_4970,N_4576);
xnor U5309 (N_5309,N_4895,N_4528);
nor U5310 (N_5310,N_4820,N_4838);
nor U5311 (N_5311,N_4956,N_4707);
or U5312 (N_5312,N_4703,N_4961);
xor U5313 (N_5313,N_4821,N_4669);
nor U5314 (N_5314,N_4925,N_4907);
xnor U5315 (N_5315,N_4862,N_4522);
nor U5316 (N_5316,N_4943,N_4992);
nand U5317 (N_5317,N_4955,N_4692);
nor U5318 (N_5318,N_4734,N_4765);
nor U5319 (N_5319,N_4674,N_4916);
and U5320 (N_5320,N_4987,N_4683);
nand U5321 (N_5321,N_4620,N_4665);
and U5322 (N_5322,N_4994,N_4737);
nor U5323 (N_5323,N_4787,N_4589);
nand U5324 (N_5324,N_4605,N_4803);
nor U5325 (N_5325,N_4917,N_4552);
xor U5326 (N_5326,N_4593,N_4774);
and U5327 (N_5327,N_4702,N_4799);
xor U5328 (N_5328,N_4831,N_4825);
or U5329 (N_5329,N_4984,N_4657);
nand U5330 (N_5330,N_4881,N_4625);
and U5331 (N_5331,N_4539,N_4699);
and U5332 (N_5332,N_4674,N_4855);
and U5333 (N_5333,N_4609,N_4649);
nand U5334 (N_5334,N_4751,N_4708);
nand U5335 (N_5335,N_4847,N_4540);
nor U5336 (N_5336,N_4538,N_4747);
xor U5337 (N_5337,N_4871,N_4612);
xor U5338 (N_5338,N_4621,N_4702);
or U5339 (N_5339,N_4506,N_4669);
nand U5340 (N_5340,N_4810,N_4942);
or U5341 (N_5341,N_4754,N_4968);
nand U5342 (N_5342,N_4575,N_4643);
xor U5343 (N_5343,N_4867,N_4784);
nand U5344 (N_5344,N_4519,N_4643);
and U5345 (N_5345,N_4628,N_4998);
nor U5346 (N_5346,N_4663,N_4696);
or U5347 (N_5347,N_4600,N_4901);
nand U5348 (N_5348,N_4818,N_4886);
or U5349 (N_5349,N_4947,N_4589);
or U5350 (N_5350,N_4767,N_4798);
nor U5351 (N_5351,N_4723,N_4825);
nor U5352 (N_5352,N_4756,N_4731);
xnor U5353 (N_5353,N_4629,N_4814);
and U5354 (N_5354,N_4665,N_4899);
nor U5355 (N_5355,N_4644,N_4524);
or U5356 (N_5356,N_4997,N_4692);
nand U5357 (N_5357,N_4737,N_4721);
nor U5358 (N_5358,N_4883,N_4668);
nor U5359 (N_5359,N_4637,N_4543);
xor U5360 (N_5360,N_4677,N_4660);
nor U5361 (N_5361,N_4807,N_4957);
nand U5362 (N_5362,N_4787,N_4857);
and U5363 (N_5363,N_4743,N_4770);
nor U5364 (N_5364,N_4739,N_4644);
nand U5365 (N_5365,N_4839,N_4540);
or U5366 (N_5366,N_4616,N_4998);
nand U5367 (N_5367,N_4558,N_4620);
or U5368 (N_5368,N_4534,N_4968);
nand U5369 (N_5369,N_4831,N_4711);
and U5370 (N_5370,N_4697,N_4897);
and U5371 (N_5371,N_4826,N_4798);
or U5372 (N_5372,N_4786,N_4797);
or U5373 (N_5373,N_4720,N_4875);
or U5374 (N_5374,N_4612,N_4827);
and U5375 (N_5375,N_4599,N_4800);
nor U5376 (N_5376,N_4501,N_4620);
xor U5377 (N_5377,N_4983,N_4608);
and U5378 (N_5378,N_4579,N_4670);
nor U5379 (N_5379,N_4745,N_4572);
xor U5380 (N_5380,N_4586,N_4724);
nor U5381 (N_5381,N_4883,N_4695);
nand U5382 (N_5382,N_4811,N_4977);
and U5383 (N_5383,N_4546,N_4750);
nor U5384 (N_5384,N_4827,N_4591);
nand U5385 (N_5385,N_4574,N_4701);
or U5386 (N_5386,N_4683,N_4687);
nor U5387 (N_5387,N_4946,N_4762);
nor U5388 (N_5388,N_4591,N_4982);
or U5389 (N_5389,N_4701,N_4692);
and U5390 (N_5390,N_4819,N_4562);
nor U5391 (N_5391,N_4717,N_4639);
or U5392 (N_5392,N_4652,N_4849);
xor U5393 (N_5393,N_4889,N_4770);
or U5394 (N_5394,N_4684,N_4573);
and U5395 (N_5395,N_4858,N_4800);
nand U5396 (N_5396,N_4804,N_4617);
and U5397 (N_5397,N_4577,N_4736);
xor U5398 (N_5398,N_4884,N_4632);
nand U5399 (N_5399,N_4860,N_4831);
or U5400 (N_5400,N_4556,N_4683);
and U5401 (N_5401,N_4643,N_4876);
xnor U5402 (N_5402,N_4652,N_4952);
or U5403 (N_5403,N_4540,N_4970);
nand U5404 (N_5404,N_4946,N_4770);
or U5405 (N_5405,N_4615,N_4677);
xor U5406 (N_5406,N_4744,N_4806);
xor U5407 (N_5407,N_4803,N_4527);
or U5408 (N_5408,N_4631,N_4929);
and U5409 (N_5409,N_4895,N_4906);
xor U5410 (N_5410,N_4581,N_4531);
or U5411 (N_5411,N_4500,N_4654);
nor U5412 (N_5412,N_4570,N_4988);
or U5413 (N_5413,N_4646,N_4692);
xor U5414 (N_5414,N_4964,N_4637);
xor U5415 (N_5415,N_4986,N_4897);
or U5416 (N_5416,N_4851,N_4731);
nand U5417 (N_5417,N_4953,N_4682);
and U5418 (N_5418,N_4537,N_4647);
nand U5419 (N_5419,N_4533,N_4970);
nand U5420 (N_5420,N_4794,N_4917);
and U5421 (N_5421,N_4662,N_4922);
and U5422 (N_5422,N_4994,N_4970);
or U5423 (N_5423,N_4538,N_4999);
nand U5424 (N_5424,N_4815,N_4867);
nor U5425 (N_5425,N_4722,N_4828);
nand U5426 (N_5426,N_4973,N_4894);
nand U5427 (N_5427,N_4729,N_4563);
nor U5428 (N_5428,N_4747,N_4552);
and U5429 (N_5429,N_4768,N_4566);
and U5430 (N_5430,N_4691,N_4659);
nand U5431 (N_5431,N_4835,N_4914);
nand U5432 (N_5432,N_4958,N_4662);
xnor U5433 (N_5433,N_4689,N_4633);
nand U5434 (N_5434,N_4966,N_4927);
or U5435 (N_5435,N_4764,N_4986);
nor U5436 (N_5436,N_4626,N_4793);
xor U5437 (N_5437,N_4546,N_4825);
nand U5438 (N_5438,N_4874,N_4608);
xnor U5439 (N_5439,N_4514,N_4724);
and U5440 (N_5440,N_4938,N_4684);
and U5441 (N_5441,N_4575,N_4794);
or U5442 (N_5442,N_4882,N_4629);
nor U5443 (N_5443,N_4562,N_4584);
and U5444 (N_5444,N_4918,N_4856);
and U5445 (N_5445,N_4848,N_4938);
xnor U5446 (N_5446,N_4585,N_4706);
nand U5447 (N_5447,N_4835,N_4514);
nand U5448 (N_5448,N_4684,N_4786);
or U5449 (N_5449,N_4644,N_4987);
nor U5450 (N_5450,N_4785,N_4868);
nor U5451 (N_5451,N_4803,N_4763);
or U5452 (N_5452,N_4665,N_4543);
or U5453 (N_5453,N_4858,N_4693);
and U5454 (N_5454,N_4848,N_4593);
nor U5455 (N_5455,N_4884,N_4883);
xor U5456 (N_5456,N_4576,N_4691);
and U5457 (N_5457,N_4815,N_4915);
nor U5458 (N_5458,N_4871,N_4649);
nor U5459 (N_5459,N_4820,N_4551);
nand U5460 (N_5460,N_4672,N_4523);
nand U5461 (N_5461,N_4559,N_4696);
or U5462 (N_5462,N_4548,N_4817);
nand U5463 (N_5463,N_4871,N_4753);
nand U5464 (N_5464,N_4512,N_4750);
nor U5465 (N_5465,N_4585,N_4718);
and U5466 (N_5466,N_4768,N_4745);
or U5467 (N_5467,N_4732,N_4617);
xor U5468 (N_5468,N_4718,N_4612);
and U5469 (N_5469,N_4952,N_4638);
xnor U5470 (N_5470,N_4529,N_4653);
and U5471 (N_5471,N_4805,N_4789);
nor U5472 (N_5472,N_4696,N_4922);
and U5473 (N_5473,N_4868,N_4720);
xor U5474 (N_5474,N_4564,N_4805);
or U5475 (N_5475,N_4967,N_4673);
and U5476 (N_5476,N_4909,N_4792);
xnor U5477 (N_5477,N_4574,N_4835);
or U5478 (N_5478,N_4680,N_4929);
nand U5479 (N_5479,N_4735,N_4821);
nor U5480 (N_5480,N_4623,N_4961);
or U5481 (N_5481,N_4881,N_4794);
nand U5482 (N_5482,N_4561,N_4582);
nand U5483 (N_5483,N_4665,N_4761);
or U5484 (N_5484,N_4750,N_4638);
xnor U5485 (N_5485,N_4995,N_4620);
xor U5486 (N_5486,N_4682,N_4781);
and U5487 (N_5487,N_4719,N_4672);
or U5488 (N_5488,N_4562,N_4629);
xnor U5489 (N_5489,N_4741,N_4900);
or U5490 (N_5490,N_4502,N_4735);
and U5491 (N_5491,N_4965,N_4745);
nand U5492 (N_5492,N_4895,N_4871);
nor U5493 (N_5493,N_4682,N_4803);
and U5494 (N_5494,N_4681,N_4538);
and U5495 (N_5495,N_4786,N_4725);
xor U5496 (N_5496,N_4506,N_4618);
or U5497 (N_5497,N_4698,N_4893);
nor U5498 (N_5498,N_4605,N_4599);
nor U5499 (N_5499,N_4780,N_4744);
xnor U5500 (N_5500,N_5156,N_5430);
nand U5501 (N_5501,N_5149,N_5075);
nor U5502 (N_5502,N_5268,N_5161);
or U5503 (N_5503,N_5215,N_5187);
nor U5504 (N_5504,N_5303,N_5236);
nand U5505 (N_5505,N_5457,N_5346);
or U5506 (N_5506,N_5017,N_5091);
or U5507 (N_5507,N_5221,N_5154);
nor U5508 (N_5508,N_5269,N_5064);
nand U5509 (N_5509,N_5033,N_5189);
or U5510 (N_5510,N_5420,N_5447);
or U5511 (N_5511,N_5116,N_5280);
nor U5512 (N_5512,N_5047,N_5314);
nor U5513 (N_5513,N_5065,N_5066);
nand U5514 (N_5514,N_5068,N_5060);
nor U5515 (N_5515,N_5050,N_5436);
xor U5516 (N_5516,N_5455,N_5308);
nand U5517 (N_5517,N_5467,N_5493);
and U5518 (N_5518,N_5492,N_5421);
and U5519 (N_5519,N_5078,N_5416);
or U5520 (N_5520,N_5106,N_5213);
and U5521 (N_5521,N_5177,N_5401);
nor U5522 (N_5522,N_5301,N_5443);
xor U5523 (N_5523,N_5082,N_5342);
nor U5524 (N_5524,N_5333,N_5316);
xnor U5525 (N_5525,N_5118,N_5331);
xnor U5526 (N_5526,N_5003,N_5124);
nand U5527 (N_5527,N_5466,N_5260);
xor U5528 (N_5528,N_5037,N_5107);
and U5529 (N_5529,N_5405,N_5144);
or U5530 (N_5530,N_5191,N_5016);
xnor U5531 (N_5531,N_5497,N_5427);
and U5532 (N_5532,N_5136,N_5234);
nor U5533 (N_5533,N_5160,N_5379);
nor U5534 (N_5534,N_5406,N_5120);
xnor U5535 (N_5535,N_5245,N_5356);
or U5536 (N_5536,N_5272,N_5336);
nand U5537 (N_5537,N_5434,N_5079);
and U5538 (N_5538,N_5031,N_5418);
xor U5539 (N_5539,N_5393,N_5454);
nand U5540 (N_5540,N_5203,N_5139);
nand U5541 (N_5541,N_5178,N_5055);
nand U5542 (N_5542,N_5230,N_5367);
nand U5543 (N_5543,N_5086,N_5038);
and U5544 (N_5544,N_5369,N_5036);
and U5545 (N_5545,N_5372,N_5053);
and U5546 (N_5546,N_5171,N_5122);
xor U5547 (N_5547,N_5473,N_5061);
nor U5548 (N_5548,N_5469,N_5209);
or U5549 (N_5549,N_5253,N_5435);
nor U5550 (N_5550,N_5130,N_5085);
xnor U5551 (N_5551,N_5432,N_5476);
nor U5552 (N_5552,N_5001,N_5229);
or U5553 (N_5553,N_5121,N_5226);
nand U5554 (N_5554,N_5417,N_5362);
or U5555 (N_5555,N_5153,N_5207);
or U5556 (N_5556,N_5373,N_5010);
nor U5557 (N_5557,N_5448,N_5378);
and U5558 (N_5558,N_5340,N_5045);
xnor U5559 (N_5559,N_5477,N_5408);
nand U5560 (N_5560,N_5415,N_5096);
nand U5561 (N_5561,N_5168,N_5030);
nor U5562 (N_5562,N_5487,N_5232);
xnor U5563 (N_5563,N_5310,N_5483);
xor U5564 (N_5564,N_5433,N_5142);
nand U5565 (N_5565,N_5345,N_5444);
xnor U5566 (N_5566,N_5228,N_5163);
and U5567 (N_5567,N_5298,N_5489);
xnor U5568 (N_5568,N_5081,N_5238);
xnor U5569 (N_5569,N_5088,N_5145);
nand U5570 (N_5570,N_5000,N_5276);
or U5571 (N_5571,N_5446,N_5468);
nand U5572 (N_5572,N_5488,N_5227);
xor U5573 (N_5573,N_5004,N_5292);
nand U5574 (N_5574,N_5322,N_5470);
nor U5575 (N_5575,N_5248,N_5319);
nand U5576 (N_5576,N_5257,N_5196);
and U5577 (N_5577,N_5256,N_5026);
or U5578 (N_5578,N_5425,N_5201);
nand U5579 (N_5579,N_5471,N_5093);
nand U5580 (N_5580,N_5135,N_5043);
xor U5581 (N_5581,N_5158,N_5296);
nor U5582 (N_5582,N_5354,N_5185);
xnor U5583 (N_5583,N_5219,N_5323);
xor U5584 (N_5584,N_5294,N_5042);
and U5585 (N_5585,N_5208,N_5205);
nor U5586 (N_5586,N_5181,N_5325);
nand U5587 (N_5587,N_5353,N_5199);
nor U5588 (N_5588,N_5162,N_5383);
and U5589 (N_5589,N_5242,N_5478);
nand U5590 (N_5590,N_5251,N_5214);
nand U5591 (N_5591,N_5289,N_5022);
xnor U5592 (N_5592,N_5307,N_5452);
nand U5593 (N_5593,N_5374,N_5442);
nor U5594 (N_5594,N_5380,N_5009);
xnor U5595 (N_5595,N_5456,N_5264);
nand U5596 (N_5596,N_5271,N_5391);
or U5597 (N_5597,N_5411,N_5239);
and U5598 (N_5598,N_5140,N_5029);
xor U5599 (N_5599,N_5388,N_5148);
or U5600 (N_5600,N_5258,N_5089);
nand U5601 (N_5601,N_5463,N_5222);
or U5602 (N_5602,N_5225,N_5499);
xnor U5603 (N_5603,N_5460,N_5044);
or U5604 (N_5604,N_5198,N_5327);
nand U5605 (N_5605,N_5376,N_5461);
nor U5606 (N_5606,N_5324,N_5375);
xor U5607 (N_5607,N_5063,N_5167);
or U5608 (N_5608,N_5397,N_5250);
and U5609 (N_5609,N_5368,N_5328);
or U5610 (N_5610,N_5414,N_5223);
and U5611 (N_5611,N_5220,N_5287);
xnor U5612 (N_5612,N_5123,N_5173);
nor U5613 (N_5613,N_5057,N_5180);
or U5614 (N_5614,N_5073,N_5265);
xor U5615 (N_5615,N_5424,N_5283);
xnor U5616 (N_5616,N_5194,N_5495);
nor U5617 (N_5617,N_5361,N_5494);
xnor U5618 (N_5618,N_5051,N_5034);
nor U5619 (N_5619,N_5103,N_5138);
or U5620 (N_5620,N_5335,N_5218);
and U5621 (N_5621,N_5024,N_5170);
and U5622 (N_5622,N_5182,N_5498);
nand U5623 (N_5623,N_5392,N_5472);
xor U5624 (N_5624,N_5491,N_5312);
nor U5625 (N_5625,N_5146,N_5217);
and U5626 (N_5626,N_5246,N_5326);
nor U5627 (N_5627,N_5098,N_5113);
or U5628 (N_5628,N_5126,N_5077);
or U5629 (N_5629,N_5211,N_5249);
or U5630 (N_5630,N_5147,N_5422);
nand U5631 (N_5631,N_5451,N_5216);
nor U5632 (N_5632,N_5008,N_5100);
xor U5633 (N_5633,N_5290,N_5370);
or U5634 (N_5634,N_5315,N_5385);
xnor U5635 (N_5635,N_5465,N_5450);
nand U5636 (N_5636,N_5054,N_5302);
and U5637 (N_5637,N_5150,N_5202);
or U5638 (N_5638,N_5412,N_5143);
xnor U5639 (N_5639,N_5020,N_5363);
nor U5640 (N_5640,N_5394,N_5224);
nand U5641 (N_5641,N_5067,N_5243);
nand U5642 (N_5642,N_5058,N_5350);
xor U5643 (N_5643,N_5459,N_5400);
or U5644 (N_5644,N_5359,N_5090);
or U5645 (N_5645,N_5083,N_5048);
nand U5646 (N_5646,N_5304,N_5396);
and U5647 (N_5647,N_5266,N_5481);
nor U5648 (N_5648,N_5399,N_5186);
nand U5649 (N_5649,N_5413,N_5329);
xnor U5650 (N_5650,N_5440,N_5395);
and U5651 (N_5651,N_5006,N_5099);
nor U5652 (N_5652,N_5259,N_5423);
nor U5653 (N_5653,N_5458,N_5231);
and U5654 (N_5654,N_5384,N_5371);
or U5655 (N_5655,N_5095,N_5108);
nor U5656 (N_5656,N_5041,N_5437);
and U5657 (N_5657,N_5119,N_5129);
xnor U5658 (N_5658,N_5313,N_5348);
xor U5659 (N_5659,N_5255,N_5190);
or U5660 (N_5660,N_5012,N_5358);
and U5661 (N_5661,N_5152,N_5351);
or U5662 (N_5662,N_5131,N_5134);
xor U5663 (N_5663,N_5141,N_5453);
nand U5664 (N_5664,N_5431,N_5309);
and U5665 (N_5665,N_5021,N_5349);
nor U5666 (N_5666,N_5254,N_5339);
nor U5667 (N_5667,N_5115,N_5111);
nor U5668 (N_5668,N_5052,N_5027);
nor U5669 (N_5669,N_5321,N_5407);
xor U5670 (N_5670,N_5005,N_5267);
nor U5671 (N_5671,N_5352,N_5252);
nand U5672 (N_5672,N_5341,N_5014);
or U5673 (N_5673,N_5398,N_5019);
or U5674 (N_5674,N_5200,N_5428);
and U5675 (N_5675,N_5278,N_5485);
xor U5676 (N_5676,N_5300,N_5032);
or U5677 (N_5677,N_5076,N_5480);
nor U5678 (N_5678,N_5332,N_5059);
nor U5679 (N_5679,N_5184,N_5305);
and U5680 (N_5680,N_5285,N_5484);
nor U5681 (N_5681,N_5377,N_5273);
or U5682 (N_5682,N_5013,N_5311);
nand U5683 (N_5683,N_5334,N_5365);
nand U5684 (N_5684,N_5474,N_5175);
nor U5685 (N_5685,N_5475,N_5237);
or U5686 (N_5686,N_5482,N_5344);
nor U5687 (N_5687,N_5125,N_5409);
or U5688 (N_5688,N_5132,N_5049);
or U5689 (N_5689,N_5410,N_5306);
nand U5690 (N_5690,N_5261,N_5382);
nor U5691 (N_5691,N_5188,N_5288);
and U5692 (N_5692,N_5101,N_5159);
and U5693 (N_5693,N_5381,N_5429);
nand U5694 (N_5694,N_5110,N_5404);
nor U5695 (N_5695,N_5011,N_5133);
or U5696 (N_5696,N_5072,N_5212);
nand U5697 (N_5697,N_5233,N_5439);
xor U5698 (N_5698,N_5172,N_5317);
or U5699 (N_5699,N_5069,N_5281);
and U5700 (N_5700,N_5357,N_5389);
xor U5701 (N_5701,N_5299,N_5240);
or U5702 (N_5702,N_5007,N_5002);
xor U5703 (N_5703,N_5056,N_5270);
nand U5704 (N_5704,N_5241,N_5137);
xor U5705 (N_5705,N_5235,N_5204);
nand U5706 (N_5706,N_5169,N_5114);
nor U5707 (N_5707,N_5070,N_5355);
and U5708 (N_5708,N_5360,N_5155);
nor U5709 (N_5709,N_5151,N_5028);
nand U5710 (N_5710,N_5274,N_5176);
nand U5711 (N_5711,N_5210,N_5174);
xor U5712 (N_5712,N_5275,N_5479);
nand U5713 (N_5713,N_5486,N_5286);
nor U5714 (N_5714,N_5337,N_5157);
nand U5715 (N_5715,N_5282,N_5295);
nand U5716 (N_5716,N_5318,N_5426);
or U5717 (N_5717,N_5263,N_5183);
nand U5718 (N_5718,N_5039,N_5297);
or U5719 (N_5719,N_5015,N_5364);
nor U5720 (N_5720,N_5035,N_5330);
xor U5721 (N_5721,N_5347,N_5195);
nand U5722 (N_5722,N_5366,N_5496);
or U5723 (N_5723,N_5441,N_5128);
or U5724 (N_5724,N_5291,N_5206);
or U5725 (N_5725,N_5102,N_5192);
xnor U5726 (N_5726,N_5390,N_5386);
and U5727 (N_5727,N_5046,N_5462);
nand U5728 (N_5728,N_5464,N_5071);
or U5729 (N_5729,N_5025,N_5293);
nand U5730 (N_5730,N_5445,N_5279);
nand U5731 (N_5731,N_5097,N_5438);
xnor U5732 (N_5732,N_5164,N_5165);
or U5733 (N_5733,N_5094,N_5244);
xnor U5734 (N_5734,N_5084,N_5104);
or U5735 (N_5735,N_5419,N_5018);
and U5736 (N_5736,N_5490,N_5109);
xnor U5737 (N_5737,N_5284,N_5320);
and U5738 (N_5738,N_5023,N_5449);
xnor U5739 (N_5739,N_5105,N_5117);
nand U5740 (N_5740,N_5197,N_5087);
or U5741 (N_5741,N_5179,N_5402);
xnor U5742 (N_5742,N_5166,N_5040);
or U5743 (N_5743,N_5343,N_5277);
xnor U5744 (N_5744,N_5074,N_5262);
or U5745 (N_5745,N_5338,N_5062);
nor U5746 (N_5746,N_5127,N_5080);
xor U5747 (N_5747,N_5112,N_5092);
xnor U5748 (N_5748,N_5403,N_5193);
nor U5749 (N_5749,N_5387,N_5247);
and U5750 (N_5750,N_5005,N_5450);
xnor U5751 (N_5751,N_5416,N_5072);
xor U5752 (N_5752,N_5230,N_5227);
and U5753 (N_5753,N_5321,N_5360);
and U5754 (N_5754,N_5442,N_5449);
or U5755 (N_5755,N_5420,N_5364);
nand U5756 (N_5756,N_5423,N_5454);
or U5757 (N_5757,N_5253,N_5251);
or U5758 (N_5758,N_5041,N_5010);
nor U5759 (N_5759,N_5030,N_5132);
xor U5760 (N_5760,N_5407,N_5164);
nor U5761 (N_5761,N_5132,N_5118);
or U5762 (N_5762,N_5279,N_5299);
xnor U5763 (N_5763,N_5047,N_5268);
xor U5764 (N_5764,N_5477,N_5140);
xnor U5765 (N_5765,N_5285,N_5493);
nor U5766 (N_5766,N_5494,N_5278);
or U5767 (N_5767,N_5255,N_5101);
xnor U5768 (N_5768,N_5174,N_5320);
and U5769 (N_5769,N_5316,N_5359);
or U5770 (N_5770,N_5121,N_5450);
nor U5771 (N_5771,N_5456,N_5418);
and U5772 (N_5772,N_5177,N_5481);
xnor U5773 (N_5773,N_5118,N_5176);
nor U5774 (N_5774,N_5264,N_5180);
or U5775 (N_5775,N_5039,N_5354);
and U5776 (N_5776,N_5036,N_5198);
xor U5777 (N_5777,N_5457,N_5496);
nand U5778 (N_5778,N_5154,N_5452);
or U5779 (N_5779,N_5314,N_5090);
nor U5780 (N_5780,N_5149,N_5351);
or U5781 (N_5781,N_5339,N_5032);
xnor U5782 (N_5782,N_5360,N_5033);
nand U5783 (N_5783,N_5216,N_5411);
nand U5784 (N_5784,N_5048,N_5080);
nand U5785 (N_5785,N_5431,N_5189);
nor U5786 (N_5786,N_5179,N_5238);
or U5787 (N_5787,N_5214,N_5292);
nor U5788 (N_5788,N_5408,N_5006);
or U5789 (N_5789,N_5433,N_5419);
xnor U5790 (N_5790,N_5121,N_5088);
or U5791 (N_5791,N_5183,N_5294);
nand U5792 (N_5792,N_5039,N_5362);
xnor U5793 (N_5793,N_5277,N_5444);
nand U5794 (N_5794,N_5250,N_5011);
xor U5795 (N_5795,N_5358,N_5194);
nor U5796 (N_5796,N_5370,N_5492);
xnor U5797 (N_5797,N_5311,N_5393);
xor U5798 (N_5798,N_5215,N_5343);
nand U5799 (N_5799,N_5224,N_5144);
and U5800 (N_5800,N_5380,N_5142);
xor U5801 (N_5801,N_5090,N_5489);
and U5802 (N_5802,N_5052,N_5116);
xor U5803 (N_5803,N_5304,N_5336);
nor U5804 (N_5804,N_5140,N_5055);
and U5805 (N_5805,N_5092,N_5035);
nand U5806 (N_5806,N_5080,N_5457);
xnor U5807 (N_5807,N_5262,N_5203);
and U5808 (N_5808,N_5164,N_5495);
or U5809 (N_5809,N_5050,N_5329);
nor U5810 (N_5810,N_5101,N_5413);
nand U5811 (N_5811,N_5211,N_5159);
or U5812 (N_5812,N_5444,N_5034);
or U5813 (N_5813,N_5467,N_5450);
or U5814 (N_5814,N_5336,N_5300);
nand U5815 (N_5815,N_5440,N_5284);
xnor U5816 (N_5816,N_5141,N_5354);
nand U5817 (N_5817,N_5194,N_5477);
xor U5818 (N_5818,N_5220,N_5139);
nor U5819 (N_5819,N_5239,N_5011);
and U5820 (N_5820,N_5369,N_5200);
nor U5821 (N_5821,N_5129,N_5211);
nor U5822 (N_5822,N_5124,N_5048);
nand U5823 (N_5823,N_5323,N_5032);
or U5824 (N_5824,N_5374,N_5294);
nand U5825 (N_5825,N_5212,N_5382);
xor U5826 (N_5826,N_5188,N_5147);
and U5827 (N_5827,N_5145,N_5282);
nand U5828 (N_5828,N_5050,N_5176);
nand U5829 (N_5829,N_5398,N_5284);
nand U5830 (N_5830,N_5185,N_5153);
nand U5831 (N_5831,N_5012,N_5407);
xnor U5832 (N_5832,N_5071,N_5066);
or U5833 (N_5833,N_5446,N_5389);
and U5834 (N_5834,N_5462,N_5027);
nor U5835 (N_5835,N_5476,N_5023);
xor U5836 (N_5836,N_5179,N_5246);
and U5837 (N_5837,N_5397,N_5292);
and U5838 (N_5838,N_5427,N_5073);
and U5839 (N_5839,N_5237,N_5318);
xor U5840 (N_5840,N_5102,N_5053);
nor U5841 (N_5841,N_5375,N_5069);
and U5842 (N_5842,N_5457,N_5466);
nor U5843 (N_5843,N_5242,N_5446);
xor U5844 (N_5844,N_5110,N_5133);
nand U5845 (N_5845,N_5228,N_5012);
or U5846 (N_5846,N_5250,N_5142);
or U5847 (N_5847,N_5368,N_5188);
nor U5848 (N_5848,N_5433,N_5222);
nand U5849 (N_5849,N_5300,N_5127);
nor U5850 (N_5850,N_5046,N_5197);
and U5851 (N_5851,N_5141,N_5346);
nor U5852 (N_5852,N_5449,N_5453);
nor U5853 (N_5853,N_5416,N_5081);
or U5854 (N_5854,N_5346,N_5171);
nor U5855 (N_5855,N_5141,N_5045);
xnor U5856 (N_5856,N_5122,N_5424);
nand U5857 (N_5857,N_5089,N_5339);
nand U5858 (N_5858,N_5325,N_5037);
or U5859 (N_5859,N_5409,N_5149);
xor U5860 (N_5860,N_5072,N_5310);
nand U5861 (N_5861,N_5482,N_5330);
xor U5862 (N_5862,N_5181,N_5205);
and U5863 (N_5863,N_5020,N_5270);
or U5864 (N_5864,N_5221,N_5151);
or U5865 (N_5865,N_5304,N_5387);
xnor U5866 (N_5866,N_5287,N_5088);
nor U5867 (N_5867,N_5152,N_5303);
xor U5868 (N_5868,N_5301,N_5017);
xnor U5869 (N_5869,N_5098,N_5392);
xnor U5870 (N_5870,N_5417,N_5300);
nor U5871 (N_5871,N_5195,N_5431);
xor U5872 (N_5872,N_5317,N_5249);
and U5873 (N_5873,N_5210,N_5467);
or U5874 (N_5874,N_5393,N_5342);
or U5875 (N_5875,N_5358,N_5091);
nand U5876 (N_5876,N_5348,N_5436);
nand U5877 (N_5877,N_5331,N_5087);
xnor U5878 (N_5878,N_5496,N_5432);
nor U5879 (N_5879,N_5181,N_5140);
xor U5880 (N_5880,N_5185,N_5044);
xor U5881 (N_5881,N_5252,N_5350);
xor U5882 (N_5882,N_5366,N_5004);
or U5883 (N_5883,N_5395,N_5071);
or U5884 (N_5884,N_5197,N_5054);
nand U5885 (N_5885,N_5036,N_5056);
and U5886 (N_5886,N_5467,N_5455);
and U5887 (N_5887,N_5202,N_5357);
nand U5888 (N_5888,N_5141,N_5131);
or U5889 (N_5889,N_5079,N_5243);
or U5890 (N_5890,N_5382,N_5333);
nand U5891 (N_5891,N_5143,N_5107);
nor U5892 (N_5892,N_5429,N_5335);
xnor U5893 (N_5893,N_5003,N_5069);
xnor U5894 (N_5894,N_5199,N_5154);
and U5895 (N_5895,N_5332,N_5202);
xnor U5896 (N_5896,N_5421,N_5184);
xor U5897 (N_5897,N_5124,N_5411);
or U5898 (N_5898,N_5080,N_5155);
xor U5899 (N_5899,N_5070,N_5169);
nand U5900 (N_5900,N_5450,N_5383);
and U5901 (N_5901,N_5301,N_5132);
nand U5902 (N_5902,N_5270,N_5050);
nor U5903 (N_5903,N_5272,N_5191);
and U5904 (N_5904,N_5079,N_5051);
nor U5905 (N_5905,N_5309,N_5229);
nor U5906 (N_5906,N_5165,N_5365);
nor U5907 (N_5907,N_5211,N_5313);
nor U5908 (N_5908,N_5281,N_5153);
nor U5909 (N_5909,N_5421,N_5354);
nand U5910 (N_5910,N_5456,N_5244);
and U5911 (N_5911,N_5132,N_5355);
nor U5912 (N_5912,N_5246,N_5117);
xnor U5913 (N_5913,N_5060,N_5100);
nor U5914 (N_5914,N_5252,N_5078);
nor U5915 (N_5915,N_5131,N_5002);
and U5916 (N_5916,N_5431,N_5300);
nand U5917 (N_5917,N_5326,N_5382);
nand U5918 (N_5918,N_5331,N_5236);
nand U5919 (N_5919,N_5329,N_5042);
or U5920 (N_5920,N_5346,N_5422);
nor U5921 (N_5921,N_5194,N_5008);
nand U5922 (N_5922,N_5132,N_5468);
and U5923 (N_5923,N_5074,N_5024);
xor U5924 (N_5924,N_5076,N_5088);
nor U5925 (N_5925,N_5463,N_5045);
nand U5926 (N_5926,N_5016,N_5489);
or U5927 (N_5927,N_5271,N_5017);
and U5928 (N_5928,N_5345,N_5382);
nand U5929 (N_5929,N_5237,N_5093);
or U5930 (N_5930,N_5208,N_5474);
nor U5931 (N_5931,N_5360,N_5490);
or U5932 (N_5932,N_5276,N_5153);
nand U5933 (N_5933,N_5123,N_5169);
nand U5934 (N_5934,N_5347,N_5408);
xnor U5935 (N_5935,N_5123,N_5029);
or U5936 (N_5936,N_5105,N_5409);
nor U5937 (N_5937,N_5460,N_5170);
nand U5938 (N_5938,N_5256,N_5001);
or U5939 (N_5939,N_5214,N_5135);
nand U5940 (N_5940,N_5143,N_5484);
and U5941 (N_5941,N_5003,N_5129);
xor U5942 (N_5942,N_5211,N_5311);
and U5943 (N_5943,N_5001,N_5032);
or U5944 (N_5944,N_5000,N_5233);
and U5945 (N_5945,N_5335,N_5316);
or U5946 (N_5946,N_5253,N_5371);
nor U5947 (N_5947,N_5069,N_5193);
nor U5948 (N_5948,N_5254,N_5464);
nor U5949 (N_5949,N_5011,N_5432);
and U5950 (N_5950,N_5385,N_5495);
or U5951 (N_5951,N_5207,N_5174);
and U5952 (N_5952,N_5016,N_5450);
nor U5953 (N_5953,N_5243,N_5004);
or U5954 (N_5954,N_5205,N_5452);
xor U5955 (N_5955,N_5214,N_5150);
xnor U5956 (N_5956,N_5328,N_5380);
nand U5957 (N_5957,N_5022,N_5031);
and U5958 (N_5958,N_5200,N_5144);
nand U5959 (N_5959,N_5493,N_5408);
nand U5960 (N_5960,N_5152,N_5325);
nand U5961 (N_5961,N_5101,N_5188);
nor U5962 (N_5962,N_5301,N_5243);
or U5963 (N_5963,N_5056,N_5188);
nand U5964 (N_5964,N_5482,N_5396);
nand U5965 (N_5965,N_5190,N_5331);
and U5966 (N_5966,N_5132,N_5367);
nand U5967 (N_5967,N_5335,N_5492);
xnor U5968 (N_5968,N_5449,N_5437);
nor U5969 (N_5969,N_5055,N_5037);
nand U5970 (N_5970,N_5149,N_5293);
nor U5971 (N_5971,N_5132,N_5128);
nor U5972 (N_5972,N_5461,N_5067);
nand U5973 (N_5973,N_5270,N_5097);
or U5974 (N_5974,N_5168,N_5413);
or U5975 (N_5975,N_5495,N_5147);
nor U5976 (N_5976,N_5310,N_5028);
nor U5977 (N_5977,N_5229,N_5061);
or U5978 (N_5978,N_5154,N_5092);
nor U5979 (N_5979,N_5151,N_5466);
or U5980 (N_5980,N_5170,N_5347);
nor U5981 (N_5981,N_5211,N_5341);
nor U5982 (N_5982,N_5164,N_5034);
or U5983 (N_5983,N_5381,N_5495);
or U5984 (N_5984,N_5422,N_5463);
and U5985 (N_5985,N_5267,N_5024);
and U5986 (N_5986,N_5118,N_5163);
nor U5987 (N_5987,N_5272,N_5212);
and U5988 (N_5988,N_5294,N_5168);
nand U5989 (N_5989,N_5179,N_5064);
xor U5990 (N_5990,N_5340,N_5429);
or U5991 (N_5991,N_5169,N_5087);
nand U5992 (N_5992,N_5385,N_5256);
nand U5993 (N_5993,N_5315,N_5432);
nand U5994 (N_5994,N_5089,N_5314);
nand U5995 (N_5995,N_5181,N_5232);
and U5996 (N_5996,N_5297,N_5288);
nand U5997 (N_5997,N_5270,N_5111);
or U5998 (N_5998,N_5358,N_5212);
nor U5999 (N_5999,N_5272,N_5401);
nand U6000 (N_6000,N_5865,N_5537);
nand U6001 (N_6001,N_5760,N_5837);
or U6002 (N_6002,N_5626,N_5606);
nand U6003 (N_6003,N_5696,N_5776);
xnor U6004 (N_6004,N_5857,N_5659);
nand U6005 (N_6005,N_5732,N_5563);
nand U6006 (N_6006,N_5541,N_5831);
or U6007 (N_6007,N_5940,N_5918);
and U6008 (N_6008,N_5785,N_5858);
and U6009 (N_6009,N_5889,N_5731);
or U6010 (N_6010,N_5583,N_5624);
xnor U6011 (N_6011,N_5892,N_5882);
nor U6012 (N_6012,N_5597,N_5799);
nand U6013 (N_6013,N_5744,N_5933);
and U6014 (N_6014,N_5978,N_5794);
or U6015 (N_6015,N_5902,N_5920);
nor U6016 (N_6016,N_5868,N_5993);
and U6017 (N_6017,N_5756,N_5554);
xor U6018 (N_6018,N_5701,N_5680);
or U6019 (N_6019,N_5848,N_5658);
nor U6020 (N_6020,N_5518,N_5965);
nor U6021 (N_6021,N_5772,N_5915);
and U6022 (N_6022,N_5833,N_5854);
and U6023 (N_6023,N_5517,N_5611);
or U6024 (N_6024,N_5675,N_5710);
xor U6025 (N_6025,N_5651,N_5951);
xnor U6026 (N_6026,N_5793,N_5938);
nor U6027 (N_6027,N_5571,N_5847);
or U6028 (N_6028,N_5888,N_5755);
nor U6029 (N_6029,N_5620,N_5769);
and U6030 (N_6030,N_5643,N_5797);
xnor U6031 (N_6031,N_5973,N_5500);
nor U6032 (N_6032,N_5861,N_5851);
nor U6033 (N_6033,N_5578,N_5780);
and U6034 (N_6034,N_5788,N_5979);
or U6035 (N_6035,N_5766,N_5535);
or U6036 (N_6036,N_5530,N_5691);
nand U6037 (N_6037,N_5507,N_5525);
or U6038 (N_6038,N_5588,N_5768);
and U6039 (N_6039,N_5976,N_5536);
xor U6040 (N_6040,N_5655,N_5670);
nand U6041 (N_6041,N_5947,N_5543);
and U6042 (N_6042,N_5593,N_5502);
nor U6043 (N_6043,N_5879,N_5757);
and U6044 (N_6044,N_5953,N_5985);
xnor U6045 (N_6045,N_5549,N_5773);
or U6046 (N_6046,N_5844,N_5817);
nor U6047 (N_6047,N_5689,N_5742);
nor U6048 (N_6048,N_5908,N_5615);
xor U6049 (N_6049,N_5955,N_5722);
xor U6050 (N_6050,N_5919,N_5647);
nand U6051 (N_6051,N_5505,N_5635);
nor U6052 (N_6052,N_5820,N_5846);
xnor U6053 (N_6053,N_5666,N_5907);
nand U6054 (N_6054,N_5891,N_5787);
or U6055 (N_6055,N_5555,N_5547);
xnor U6056 (N_6056,N_5561,N_5763);
and U6057 (N_6057,N_5790,N_5661);
xnor U6058 (N_6058,N_5568,N_5786);
and U6059 (N_6059,N_5754,N_5894);
and U6060 (N_6060,N_5683,N_5913);
and U6061 (N_6061,N_5596,N_5967);
and U6062 (N_6062,N_5531,N_5640);
or U6063 (N_6063,N_5717,N_5909);
and U6064 (N_6064,N_5912,N_5688);
nor U6065 (N_6065,N_5660,N_5840);
and U6066 (N_6066,N_5641,N_5823);
nor U6067 (N_6067,N_5897,N_5692);
nand U6068 (N_6068,N_5726,N_5644);
xor U6069 (N_6069,N_5649,N_5816);
and U6070 (N_6070,N_5671,N_5822);
xnor U6071 (N_6071,N_5628,N_5927);
nor U6072 (N_6072,N_5564,N_5825);
and U6073 (N_6073,N_5770,N_5910);
or U6074 (N_6074,N_5950,N_5715);
nor U6075 (N_6075,N_5608,N_5896);
nor U6076 (N_6076,N_5903,N_5806);
and U6077 (N_6077,N_5952,N_5815);
nor U6078 (N_6078,N_5610,N_5805);
nor U6079 (N_6079,N_5570,N_5634);
and U6080 (N_6080,N_5874,N_5709);
and U6081 (N_6081,N_5599,N_5632);
and U6082 (N_6082,N_5562,N_5703);
xor U6083 (N_6083,N_5998,N_5512);
and U6084 (N_6084,N_5591,N_5665);
nor U6085 (N_6085,N_5827,N_5975);
or U6086 (N_6086,N_5576,N_5546);
or U6087 (N_6087,N_5859,N_5949);
xor U6088 (N_6088,N_5522,N_5695);
xnor U6089 (N_6089,N_5601,N_5807);
and U6090 (N_6090,N_5727,N_5533);
nand U6091 (N_6091,N_5600,N_5566);
nor U6092 (N_6092,N_5690,N_5914);
or U6093 (N_6093,N_5829,N_5542);
xor U6094 (N_6094,N_5867,N_5828);
nor U6095 (N_6095,N_5612,N_5946);
nand U6096 (N_6096,N_5934,N_5989);
nor U6097 (N_6097,N_5916,N_5728);
and U6098 (N_6098,N_5771,N_5852);
nand U6099 (N_6099,N_5883,N_5923);
nor U6100 (N_6100,N_5981,N_5849);
and U6101 (N_6101,N_5876,N_5761);
nor U6102 (N_6102,N_5996,N_5906);
or U6103 (N_6103,N_5712,N_5924);
xnor U6104 (N_6104,N_5669,N_5759);
nand U6105 (N_6105,N_5551,N_5745);
nand U6106 (N_6106,N_5977,N_5871);
xnor U6107 (N_6107,N_5552,N_5521);
nand U6108 (N_6108,N_5528,N_5872);
nor U6109 (N_6109,N_5835,N_5839);
and U6110 (N_6110,N_5887,N_5884);
xnor U6111 (N_6111,N_5804,N_5824);
xnor U6112 (N_6112,N_5639,N_5704);
and U6113 (N_6113,N_5990,N_5932);
and U6114 (N_6114,N_5589,N_5516);
or U6115 (N_6115,N_5523,N_5988);
or U6116 (N_6116,N_5750,N_5974);
nor U6117 (N_6117,N_5743,N_5557);
and U6118 (N_6118,N_5706,N_5506);
and U6119 (N_6119,N_5654,N_5698);
xor U6120 (N_6120,N_5791,N_5767);
xnor U6121 (N_6121,N_5926,N_5880);
nor U6122 (N_6122,N_5713,N_5936);
nand U6123 (N_6123,N_5784,N_5866);
and U6124 (N_6124,N_5685,N_5718);
xnor U6125 (N_6125,N_5735,N_5961);
nand U6126 (N_6126,N_5774,N_5656);
xnor U6127 (N_6127,N_5603,N_5834);
nand U6128 (N_6128,N_5734,N_5573);
nand U6129 (N_6129,N_5982,N_5818);
xor U6130 (N_6130,N_5513,N_5987);
or U6131 (N_6131,N_5682,N_5559);
nand U6132 (N_6132,N_5813,N_5808);
or U6133 (N_6133,N_5963,N_5992);
and U6134 (N_6134,N_5623,N_5648);
and U6135 (N_6135,N_5838,N_5602);
and U6136 (N_6136,N_5752,N_5592);
or U6137 (N_6137,N_5687,N_5870);
nand U6138 (N_6138,N_5618,N_5779);
xor U6139 (N_6139,N_5605,N_5520);
or U6140 (N_6140,N_5796,N_5504);
nor U6141 (N_6141,N_5629,N_5637);
and U6142 (N_6142,N_5925,N_5901);
and U6143 (N_6143,N_5937,N_5650);
nand U6144 (N_6144,N_5556,N_5764);
or U6145 (N_6145,N_5613,N_5590);
nor U6146 (N_6146,N_5809,N_5677);
xnor U6147 (N_6147,N_5850,N_5594);
and U6148 (N_6148,N_5877,N_5777);
and U6149 (N_6149,N_5792,N_5811);
nand U6150 (N_6150,N_5935,N_5730);
nor U6151 (N_6151,N_5748,N_5911);
and U6152 (N_6152,N_5739,N_5524);
nand U6153 (N_6153,N_5509,N_5970);
or U6154 (N_6154,N_5994,N_5842);
and U6155 (N_6155,N_5821,N_5720);
nand U6156 (N_6156,N_5803,N_5881);
nand U6157 (N_6157,N_5636,N_5968);
xor U6158 (N_6158,N_5587,N_5515);
nand U6159 (N_6159,N_5630,N_5997);
nor U6160 (N_6160,N_5853,N_5569);
and U6161 (N_6161,N_5954,N_5939);
nor U6162 (N_6162,N_5686,N_5674);
or U6163 (N_6163,N_5598,N_5751);
and U6164 (N_6164,N_5890,N_5789);
and U6165 (N_6165,N_5856,N_5733);
and U6166 (N_6166,N_5798,N_5595);
nor U6167 (N_6167,N_5575,N_5527);
nand U6168 (N_6168,N_5638,N_5740);
xor U6169 (N_6169,N_5960,N_5943);
xnor U6170 (N_6170,N_5653,N_5714);
xnor U6171 (N_6171,N_5614,N_5969);
nor U6172 (N_6172,N_5544,N_5539);
and U6173 (N_6173,N_5681,N_5986);
nand U6174 (N_6174,N_5526,N_5810);
nor U6175 (N_6175,N_5607,N_5944);
nor U6176 (N_6176,N_5921,N_5999);
or U6177 (N_6177,N_5869,N_5905);
or U6178 (N_6178,N_5622,N_5765);
nor U6179 (N_6179,N_5893,N_5972);
nand U6180 (N_6180,N_5991,N_5529);
nor U6181 (N_6181,N_5633,N_5514);
xnor U6182 (N_6182,N_5721,N_5645);
nor U6183 (N_6183,N_5948,N_5737);
and U6184 (N_6184,N_5673,N_5708);
or U6185 (N_6185,N_5627,N_5716);
nand U6186 (N_6186,N_5758,N_5705);
and U6187 (N_6187,N_5885,N_5625);
nand U6188 (N_6188,N_5707,N_5738);
nand U6189 (N_6189,N_5663,N_5971);
nor U6190 (N_6190,N_5503,N_5560);
and U6191 (N_6191,N_5832,N_5642);
and U6192 (N_6192,N_5995,N_5668);
and U6193 (N_6193,N_5841,N_5711);
or U6194 (N_6194,N_5580,N_5574);
xnor U6195 (N_6195,N_5778,N_5814);
or U6196 (N_6196,N_5558,N_5510);
xor U6197 (N_6197,N_5862,N_5577);
or U6198 (N_6198,N_5945,N_5966);
nor U6199 (N_6199,N_5782,N_5878);
or U6200 (N_6200,N_5609,N_5679);
and U6201 (N_6201,N_5619,N_5678);
nand U6202 (N_6202,N_5697,N_5781);
nand U6203 (N_6203,N_5917,N_5900);
nand U6204 (N_6204,N_5929,N_5724);
nor U6205 (N_6205,N_5579,N_5723);
and U6206 (N_6206,N_5875,N_5959);
nand U6207 (N_6207,N_5550,N_5672);
nand U6208 (N_6208,N_5631,N_5753);
or U6209 (N_6209,N_5581,N_5962);
and U6210 (N_6210,N_5958,N_5741);
xor U6211 (N_6211,N_5930,N_5617);
xor U6212 (N_6212,N_5899,N_5729);
or U6213 (N_6213,N_5747,N_5775);
xor U6214 (N_6214,N_5886,N_5942);
xor U6215 (N_6215,N_5662,N_5702);
and U6216 (N_6216,N_5928,N_5795);
or U6217 (N_6217,N_5957,N_5548);
xnor U6218 (N_6218,N_5836,N_5826);
nand U6219 (N_6219,N_5983,N_5898);
xnor U6220 (N_6220,N_5984,N_5621);
or U6221 (N_6221,N_5553,N_5855);
nand U6222 (N_6222,N_5699,N_5664);
and U6223 (N_6223,N_5783,N_5922);
and U6224 (N_6224,N_5538,N_5586);
nor U6225 (N_6225,N_5904,N_5956);
and U6226 (N_6226,N_5843,N_5830);
and U6227 (N_6227,N_5746,N_5565);
nor U6228 (N_6228,N_5657,N_5511);
and U6229 (N_6229,N_5860,N_5532);
nor U6230 (N_6230,N_5693,N_5684);
and U6231 (N_6231,N_5895,N_5694);
nand U6232 (N_6232,N_5676,N_5519);
and U6233 (N_6233,N_5508,N_5545);
and U6234 (N_6234,N_5941,N_5801);
xnor U6235 (N_6235,N_5845,N_5700);
nand U6236 (N_6236,N_5652,N_5819);
nand U6237 (N_6237,N_5567,N_5873);
nand U6238 (N_6238,N_5719,N_5980);
nand U6239 (N_6239,N_5572,N_5736);
and U6240 (N_6240,N_5616,N_5964);
or U6241 (N_6241,N_5584,N_5800);
xnor U6242 (N_6242,N_5812,N_5534);
and U6243 (N_6243,N_5582,N_5667);
and U6244 (N_6244,N_5540,N_5604);
xor U6245 (N_6245,N_5863,N_5762);
nand U6246 (N_6246,N_5931,N_5864);
xnor U6247 (N_6247,N_5749,N_5501);
and U6248 (N_6248,N_5802,N_5646);
xor U6249 (N_6249,N_5725,N_5585);
and U6250 (N_6250,N_5542,N_5942);
and U6251 (N_6251,N_5719,N_5517);
xnor U6252 (N_6252,N_5566,N_5730);
or U6253 (N_6253,N_5723,N_5978);
nor U6254 (N_6254,N_5996,N_5649);
or U6255 (N_6255,N_5596,N_5758);
or U6256 (N_6256,N_5852,N_5603);
xnor U6257 (N_6257,N_5985,N_5536);
xor U6258 (N_6258,N_5565,N_5834);
xnor U6259 (N_6259,N_5659,N_5554);
and U6260 (N_6260,N_5524,N_5995);
nor U6261 (N_6261,N_5569,N_5555);
or U6262 (N_6262,N_5721,N_5816);
and U6263 (N_6263,N_5898,N_5924);
or U6264 (N_6264,N_5803,N_5938);
or U6265 (N_6265,N_5698,N_5686);
or U6266 (N_6266,N_5873,N_5578);
nor U6267 (N_6267,N_5509,N_5819);
and U6268 (N_6268,N_5682,N_5989);
xnor U6269 (N_6269,N_5753,N_5658);
nor U6270 (N_6270,N_5703,N_5509);
nand U6271 (N_6271,N_5728,N_5921);
xor U6272 (N_6272,N_5652,N_5992);
xnor U6273 (N_6273,N_5786,N_5798);
or U6274 (N_6274,N_5579,N_5742);
or U6275 (N_6275,N_5742,N_5622);
or U6276 (N_6276,N_5793,N_5565);
xnor U6277 (N_6277,N_5722,N_5609);
or U6278 (N_6278,N_5915,N_5590);
and U6279 (N_6279,N_5820,N_5986);
and U6280 (N_6280,N_5763,N_5707);
nand U6281 (N_6281,N_5791,N_5795);
nor U6282 (N_6282,N_5961,N_5837);
or U6283 (N_6283,N_5948,N_5630);
nand U6284 (N_6284,N_5880,N_5624);
nor U6285 (N_6285,N_5525,N_5501);
nand U6286 (N_6286,N_5664,N_5921);
nor U6287 (N_6287,N_5849,N_5620);
and U6288 (N_6288,N_5741,N_5833);
xor U6289 (N_6289,N_5973,N_5798);
or U6290 (N_6290,N_5730,N_5588);
or U6291 (N_6291,N_5533,N_5958);
xnor U6292 (N_6292,N_5656,N_5857);
nor U6293 (N_6293,N_5877,N_5900);
or U6294 (N_6294,N_5603,N_5689);
nor U6295 (N_6295,N_5737,N_5833);
or U6296 (N_6296,N_5656,N_5590);
or U6297 (N_6297,N_5522,N_5553);
xor U6298 (N_6298,N_5766,N_5608);
or U6299 (N_6299,N_5675,N_5731);
and U6300 (N_6300,N_5772,N_5563);
nor U6301 (N_6301,N_5883,N_5899);
and U6302 (N_6302,N_5524,N_5961);
xor U6303 (N_6303,N_5980,N_5972);
and U6304 (N_6304,N_5613,N_5945);
xor U6305 (N_6305,N_5636,N_5689);
nand U6306 (N_6306,N_5535,N_5606);
nor U6307 (N_6307,N_5527,N_5917);
nand U6308 (N_6308,N_5915,N_5871);
nand U6309 (N_6309,N_5720,N_5722);
xor U6310 (N_6310,N_5855,N_5951);
nand U6311 (N_6311,N_5787,N_5952);
and U6312 (N_6312,N_5733,N_5909);
and U6313 (N_6313,N_5942,N_5806);
or U6314 (N_6314,N_5947,N_5569);
or U6315 (N_6315,N_5502,N_5637);
nand U6316 (N_6316,N_5633,N_5750);
nand U6317 (N_6317,N_5831,N_5723);
or U6318 (N_6318,N_5992,N_5524);
or U6319 (N_6319,N_5603,N_5782);
or U6320 (N_6320,N_5733,N_5718);
nor U6321 (N_6321,N_5613,N_5650);
nor U6322 (N_6322,N_5996,N_5654);
and U6323 (N_6323,N_5679,N_5594);
xor U6324 (N_6324,N_5875,N_5775);
xor U6325 (N_6325,N_5687,N_5888);
nand U6326 (N_6326,N_5856,N_5593);
nor U6327 (N_6327,N_5746,N_5617);
or U6328 (N_6328,N_5557,N_5902);
and U6329 (N_6329,N_5994,N_5790);
and U6330 (N_6330,N_5740,N_5811);
nand U6331 (N_6331,N_5775,N_5776);
and U6332 (N_6332,N_5997,N_5635);
nand U6333 (N_6333,N_5503,N_5952);
xnor U6334 (N_6334,N_5900,N_5723);
nor U6335 (N_6335,N_5742,N_5915);
nor U6336 (N_6336,N_5683,N_5741);
xor U6337 (N_6337,N_5766,N_5553);
and U6338 (N_6338,N_5652,N_5760);
and U6339 (N_6339,N_5574,N_5997);
xor U6340 (N_6340,N_5889,N_5810);
and U6341 (N_6341,N_5878,N_5717);
or U6342 (N_6342,N_5954,N_5716);
and U6343 (N_6343,N_5621,N_5561);
or U6344 (N_6344,N_5623,N_5747);
and U6345 (N_6345,N_5531,N_5870);
or U6346 (N_6346,N_5525,N_5547);
or U6347 (N_6347,N_5596,N_5512);
nor U6348 (N_6348,N_5853,N_5992);
nand U6349 (N_6349,N_5611,N_5913);
nor U6350 (N_6350,N_5912,N_5566);
or U6351 (N_6351,N_5766,N_5821);
nand U6352 (N_6352,N_5698,N_5988);
xnor U6353 (N_6353,N_5728,N_5878);
and U6354 (N_6354,N_5703,N_5800);
nor U6355 (N_6355,N_5876,N_5517);
nor U6356 (N_6356,N_5572,N_5554);
nand U6357 (N_6357,N_5654,N_5724);
xnor U6358 (N_6358,N_5981,N_5883);
nand U6359 (N_6359,N_5769,N_5692);
nor U6360 (N_6360,N_5519,N_5893);
and U6361 (N_6361,N_5840,N_5696);
or U6362 (N_6362,N_5882,N_5648);
xor U6363 (N_6363,N_5853,N_5843);
nand U6364 (N_6364,N_5803,N_5971);
and U6365 (N_6365,N_5629,N_5686);
nor U6366 (N_6366,N_5903,N_5559);
nor U6367 (N_6367,N_5707,N_5820);
nor U6368 (N_6368,N_5694,N_5585);
xnor U6369 (N_6369,N_5553,N_5690);
or U6370 (N_6370,N_5837,N_5829);
nand U6371 (N_6371,N_5613,N_5660);
nor U6372 (N_6372,N_5673,N_5617);
nand U6373 (N_6373,N_5902,N_5664);
nand U6374 (N_6374,N_5713,N_5881);
or U6375 (N_6375,N_5615,N_5533);
or U6376 (N_6376,N_5568,N_5628);
and U6377 (N_6377,N_5987,N_5665);
and U6378 (N_6378,N_5657,N_5675);
or U6379 (N_6379,N_5929,N_5885);
and U6380 (N_6380,N_5653,N_5617);
and U6381 (N_6381,N_5528,N_5759);
nor U6382 (N_6382,N_5519,N_5960);
nor U6383 (N_6383,N_5805,N_5869);
or U6384 (N_6384,N_5506,N_5660);
and U6385 (N_6385,N_5838,N_5633);
and U6386 (N_6386,N_5535,N_5734);
nor U6387 (N_6387,N_5542,N_5926);
nor U6388 (N_6388,N_5617,N_5607);
nand U6389 (N_6389,N_5980,N_5589);
nor U6390 (N_6390,N_5965,N_5813);
xor U6391 (N_6391,N_5644,N_5895);
and U6392 (N_6392,N_5847,N_5784);
nand U6393 (N_6393,N_5506,N_5826);
or U6394 (N_6394,N_5939,N_5644);
xor U6395 (N_6395,N_5907,N_5935);
xor U6396 (N_6396,N_5523,N_5754);
xor U6397 (N_6397,N_5814,N_5703);
xnor U6398 (N_6398,N_5857,N_5985);
nand U6399 (N_6399,N_5812,N_5777);
xor U6400 (N_6400,N_5596,N_5964);
nor U6401 (N_6401,N_5504,N_5784);
or U6402 (N_6402,N_5889,N_5686);
or U6403 (N_6403,N_5625,N_5640);
xor U6404 (N_6404,N_5677,N_5958);
xnor U6405 (N_6405,N_5811,N_5563);
or U6406 (N_6406,N_5680,N_5681);
nor U6407 (N_6407,N_5614,N_5774);
nor U6408 (N_6408,N_5959,N_5894);
and U6409 (N_6409,N_5732,N_5977);
nor U6410 (N_6410,N_5524,N_5867);
and U6411 (N_6411,N_5658,N_5939);
nor U6412 (N_6412,N_5996,N_5616);
nor U6413 (N_6413,N_5905,N_5806);
and U6414 (N_6414,N_5887,N_5761);
nand U6415 (N_6415,N_5668,N_5513);
xnor U6416 (N_6416,N_5951,N_5825);
or U6417 (N_6417,N_5923,N_5537);
nor U6418 (N_6418,N_5629,N_5982);
nand U6419 (N_6419,N_5811,N_5538);
or U6420 (N_6420,N_5824,N_5742);
nand U6421 (N_6421,N_5970,N_5782);
xor U6422 (N_6422,N_5635,N_5873);
nand U6423 (N_6423,N_5959,N_5759);
nor U6424 (N_6424,N_5529,N_5844);
nand U6425 (N_6425,N_5704,N_5894);
or U6426 (N_6426,N_5732,N_5520);
nor U6427 (N_6427,N_5632,N_5967);
nor U6428 (N_6428,N_5846,N_5502);
nand U6429 (N_6429,N_5573,N_5535);
nor U6430 (N_6430,N_5568,N_5838);
nand U6431 (N_6431,N_5907,N_5858);
and U6432 (N_6432,N_5515,N_5829);
nand U6433 (N_6433,N_5891,N_5734);
or U6434 (N_6434,N_5792,N_5667);
or U6435 (N_6435,N_5996,N_5870);
nand U6436 (N_6436,N_5896,N_5824);
nand U6437 (N_6437,N_5870,N_5510);
nand U6438 (N_6438,N_5952,N_5770);
xnor U6439 (N_6439,N_5717,N_5527);
and U6440 (N_6440,N_5699,N_5790);
nor U6441 (N_6441,N_5794,N_5742);
nand U6442 (N_6442,N_5930,N_5536);
nand U6443 (N_6443,N_5737,N_5754);
xnor U6444 (N_6444,N_5535,N_5569);
or U6445 (N_6445,N_5975,N_5956);
xor U6446 (N_6446,N_5879,N_5718);
xor U6447 (N_6447,N_5795,N_5595);
and U6448 (N_6448,N_5614,N_5731);
nand U6449 (N_6449,N_5739,N_5748);
nor U6450 (N_6450,N_5783,N_5854);
xor U6451 (N_6451,N_5701,N_5949);
xnor U6452 (N_6452,N_5940,N_5803);
xor U6453 (N_6453,N_5936,N_5948);
nor U6454 (N_6454,N_5723,N_5795);
or U6455 (N_6455,N_5640,N_5695);
or U6456 (N_6456,N_5663,N_5619);
xnor U6457 (N_6457,N_5573,N_5995);
or U6458 (N_6458,N_5578,N_5801);
xor U6459 (N_6459,N_5700,N_5777);
or U6460 (N_6460,N_5775,N_5716);
or U6461 (N_6461,N_5922,N_5609);
nor U6462 (N_6462,N_5925,N_5510);
or U6463 (N_6463,N_5902,N_5546);
or U6464 (N_6464,N_5898,N_5639);
nand U6465 (N_6465,N_5842,N_5608);
nor U6466 (N_6466,N_5866,N_5537);
nand U6467 (N_6467,N_5913,N_5810);
nor U6468 (N_6468,N_5526,N_5840);
nor U6469 (N_6469,N_5983,N_5761);
nor U6470 (N_6470,N_5852,N_5957);
nor U6471 (N_6471,N_5626,N_5646);
xnor U6472 (N_6472,N_5555,N_5996);
and U6473 (N_6473,N_5728,N_5765);
nor U6474 (N_6474,N_5874,N_5521);
and U6475 (N_6475,N_5852,N_5916);
nand U6476 (N_6476,N_5744,N_5609);
xnor U6477 (N_6477,N_5743,N_5778);
nor U6478 (N_6478,N_5782,N_5948);
xor U6479 (N_6479,N_5759,N_5829);
nor U6480 (N_6480,N_5518,N_5859);
or U6481 (N_6481,N_5704,N_5697);
or U6482 (N_6482,N_5505,N_5970);
xor U6483 (N_6483,N_5606,N_5634);
nor U6484 (N_6484,N_5605,N_5725);
or U6485 (N_6485,N_5762,N_5853);
or U6486 (N_6486,N_5518,N_5909);
nand U6487 (N_6487,N_5846,N_5717);
xnor U6488 (N_6488,N_5571,N_5921);
xor U6489 (N_6489,N_5702,N_5519);
nor U6490 (N_6490,N_5867,N_5910);
nor U6491 (N_6491,N_5860,N_5633);
xor U6492 (N_6492,N_5784,N_5968);
nor U6493 (N_6493,N_5561,N_5662);
nor U6494 (N_6494,N_5775,N_5987);
or U6495 (N_6495,N_5913,N_5783);
xnor U6496 (N_6496,N_5910,N_5943);
and U6497 (N_6497,N_5894,N_5725);
nor U6498 (N_6498,N_5749,N_5552);
or U6499 (N_6499,N_5528,N_5818);
and U6500 (N_6500,N_6111,N_6411);
nor U6501 (N_6501,N_6349,N_6163);
nand U6502 (N_6502,N_6288,N_6068);
and U6503 (N_6503,N_6298,N_6206);
and U6504 (N_6504,N_6457,N_6150);
xnor U6505 (N_6505,N_6124,N_6302);
nor U6506 (N_6506,N_6126,N_6159);
nor U6507 (N_6507,N_6433,N_6460);
nand U6508 (N_6508,N_6165,N_6406);
nand U6509 (N_6509,N_6202,N_6403);
xor U6510 (N_6510,N_6205,N_6450);
nor U6511 (N_6511,N_6451,N_6107);
nand U6512 (N_6512,N_6401,N_6213);
and U6513 (N_6513,N_6410,N_6414);
or U6514 (N_6514,N_6434,N_6086);
nand U6515 (N_6515,N_6359,N_6498);
or U6516 (N_6516,N_6475,N_6032);
nand U6517 (N_6517,N_6262,N_6191);
or U6518 (N_6518,N_6372,N_6322);
or U6519 (N_6519,N_6420,N_6218);
or U6520 (N_6520,N_6249,N_6245);
or U6521 (N_6521,N_6468,N_6492);
or U6522 (N_6522,N_6296,N_6315);
xnor U6523 (N_6523,N_6198,N_6109);
nor U6524 (N_6524,N_6131,N_6229);
or U6525 (N_6525,N_6125,N_6145);
nor U6526 (N_6526,N_6120,N_6228);
xnor U6527 (N_6527,N_6258,N_6123);
nor U6528 (N_6528,N_6478,N_6044);
or U6529 (N_6529,N_6356,N_6074);
xor U6530 (N_6530,N_6170,N_6175);
or U6531 (N_6531,N_6182,N_6419);
and U6532 (N_6532,N_6423,N_6161);
and U6533 (N_6533,N_6375,N_6248);
xnor U6534 (N_6534,N_6477,N_6392);
or U6535 (N_6535,N_6254,N_6137);
and U6536 (N_6536,N_6227,N_6330);
nand U6537 (N_6537,N_6076,N_6408);
and U6538 (N_6538,N_6116,N_6179);
or U6539 (N_6539,N_6253,N_6415);
xor U6540 (N_6540,N_6438,N_6432);
nand U6541 (N_6541,N_6130,N_6234);
nor U6542 (N_6542,N_6442,N_6223);
or U6543 (N_6543,N_6336,N_6201);
nor U6544 (N_6544,N_6448,N_6365);
nor U6545 (N_6545,N_6271,N_6097);
or U6546 (N_6546,N_6447,N_6304);
nor U6547 (N_6547,N_6291,N_6225);
or U6548 (N_6548,N_6242,N_6101);
or U6549 (N_6549,N_6113,N_6220);
nor U6550 (N_6550,N_6416,N_6270);
and U6551 (N_6551,N_6247,N_6491);
nor U6552 (N_6552,N_6476,N_6473);
or U6553 (N_6553,N_6269,N_6141);
xor U6554 (N_6554,N_6022,N_6233);
or U6555 (N_6555,N_6215,N_6338);
xor U6556 (N_6556,N_6071,N_6367);
or U6557 (N_6557,N_6065,N_6169);
and U6558 (N_6558,N_6239,N_6311);
nand U6559 (N_6559,N_6441,N_6284);
nor U6560 (N_6560,N_6287,N_6292);
or U6561 (N_6561,N_6219,N_6461);
or U6562 (N_6562,N_6045,N_6050);
and U6563 (N_6563,N_6340,N_6436);
xnor U6564 (N_6564,N_6405,N_6320);
xor U6565 (N_6565,N_6464,N_6112);
nor U6566 (N_6566,N_6014,N_6329);
nand U6567 (N_6567,N_6314,N_6023);
nand U6568 (N_6568,N_6456,N_6197);
or U6569 (N_6569,N_6466,N_6010);
and U6570 (N_6570,N_6246,N_6484);
nor U6571 (N_6571,N_6252,N_6306);
xor U6572 (N_6572,N_6199,N_6216);
xor U6573 (N_6573,N_6230,N_6232);
xor U6574 (N_6574,N_6479,N_6166);
xnor U6575 (N_6575,N_6078,N_6395);
nor U6576 (N_6576,N_6485,N_6425);
nand U6577 (N_6577,N_6042,N_6259);
and U6578 (N_6578,N_6181,N_6381);
nor U6579 (N_6579,N_6463,N_6480);
and U6580 (N_6580,N_6143,N_6482);
nand U6581 (N_6581,N_6398,N_6079);
or U6582 (N_6582,N_6424,N_6147);
nand U6583 (N_6583,N_6310,N_6110);
or U6584 (N_6584,N_6462,N_6431);
or U6585 (N_6585,N_6091,N_6487);
and U6586 (N_6586,N_6121,N_6339);
nand U6587 (N_6587,N_6290,N_6458);
or U6588 (N_6588,N_6361,N_6499);
xor U6589 (N_6589,N_6200,N_6030);
and U6590 (N_6590,N_6038,N_6203);
or U6591 (N_6591,N_6020,N_6133);
nor U6592 (N_6592,N_6303,N_6155);
nor U6593 (N_6593,N_6486,N_6388);
nand U6594 (N_6594,N_6426,N_6031);
or U6595 (N_6595,N_6049,N_6353);
nand U6596 (N_6596,N_6093,N_6374);
or U6597 (N_6597,N_6013,N_6069);
nor U6598 (N_6598,N_6039,N_6404);
xnor U6599 (N_6599,N_6019,N_6370);
nor U6600 (N_6600,N_6297,N_6236);
and U6601 (N_6601,N_6047,N_6293);
xor U6602 (N_6602,N_6312,N_6240);
xor U6603 (N_6603,N_6129,N_6055);
nor U6604 (N_6604,N_6207,N_6007);
nand U6605 (N_6605,N_6208,N_6427);
xnor U6606 (N_6606,N_6168,N_6282);
nand U6607 (N_6607,N_6469,N_6280);
and U6608 (N_6608,N_6040,N_6281);
and U6609 (N_6609,N_6052,N_6127);
nor U6610 (N_6610,N_6173,N_6265);
nand U6611 (N_6611,N_6094,N_6278);
nor U6612 (N_6612,N_6108,N_6085);
nand U6613 (N_6613,N_6313,N_6021);
nand U6614 (N_6614,N_6307,N_6128);
and U6615 (N_6615,N_6148,N_6103);
and U6616 (N_6616,N_6059,N_6394);
xnor U6617 (N_6617,N_6015,N_6017);
or U6618 (N_6618,N_6051,N_6440);
or U6619 (N_6619,N_6309,N_6053);
nand U6620 (N_6620,N_6192,N_6209);
and U6621 (N_6621,N_6080,N_6114);
or U6622 (N_6622,N_6366,N_6263);
or U6623 (N_6623,N_6204,N_6183);
nand U6624 (N_6624,N_6092,N_6088);
or U6625 (N_6625,N_6000,N_6060);
or U6626 (N_6626,N_6140,N_6283);
nand U6627 (N_6627,N_6334,N_6026);
xnor U6628 (N_6628,N_6257,N_6363);
or U6629 (N_6629,N_6289,N_6318);
or U6630 (N_6630,N_6001,N_6489);
or U6631 (N_6631,N_6177,N_6305);
xnor U6632 (N_6632,N_6099,N_6352);
nand U6633 (N_6633,N_6279,N_6494);
or U6634 (N_6634,N_6029,N_6035);
or U6635 (N_6635,N_6064,N_6308);
xnor U6636 (N_6636,N_6364,N_6324);
and U6637 (N_6637,N_6294,N_6383);
and U6638 (N_6638,N_6224,N_6326);
nor U6639 (N_6639,N_6470,N_6235);
nand U6640 (N_6640,N_6054,N_6027);
or U6641 (N_6641,N_6067,N_6034);
and U6642 (N_6642,N_6379,N_6376);
or U6643 (N_6643,N_6222,N_6012);
or U6644 (N_6644,N_6267,N_6194);
and U6645 (N_6645,N_6285,N_6057);
or U6646 (N_6646,N_6028,N_6373);
or U6647 (N_6647,N_6273,N_6316);
or U6648 (N_6648,N_6244,N_6327);
nor U6649 (N_6649,N_6146,N_6443);
xor U6650 (N_6650,N_6171,N_6009);
nand U6651 (N_6651,N_6445,N_6256);
or U6652 (N_6652,N_6011,N_6378);
xor U6653 (N_6653,N_6481,N_6272);
nor U6654 (N_6654,N_6350,N_6384);
xnor U6655 (N_6655,N_6355,N_6430);
xor U6656 (N_6656,N_6452,N_6418);
and U6657 (N_6657,N_6138,N_6328);
and U6658 (N_6658,N_6260,N_6136);
and U6659 (N_6659,N_6295,N_6139);
nand U6660 (N_6660,N_6186,N_6348);
and U6661 (N_6661,N_6048,N_6357);
xor U6662 (N_6662,N_6396,N_6033);
and U6663 (N_6663,N_6342,N_6002);
nand U6664 (N_6664,N_6286,N_6185);
and U6665 (N_6665,N_6151,N_6277);
or U6666 (N_6666,N_6167,N_6041);
nor U6667 (N_6667,N_6004,N_6439);
nand U6668 (N_6668,N_6250,N_6299);
nand U6669 (N_6669,N_6465,N_6066);
xnor U6670 (N_6670,N_6152,N_6180);
nor U6671 (N_6671,N_6488,N_6300);
nand U6672 (N_6672,N_6371,N_6453);
or U6673 (N_6673,N_6184,N_6098);
nand U6674 (N_6674,N_6474,N_6087);
xnor U6675 (N_6675,N_6188,N_6226);
and U6676 (N_6676,N_6264,N_6210);
or U6677 (N_6677,N_6082,N_6331);
nor U6678 (N_6678,N_6333,N_6358);
or U6679 (N_6679,N_6446,N_6362);
or U6680 (N_6680,N_6073,N_6455);
nor U6681 (N_6681,N_6435,N_6325);
nand U6682 (N_6682,N_6368,N_6400);
nand U6683 (N_6683,N_6268,N_6118);
or U6684 (N_6684,N_6360,N_6117);
or U6685 (N_6685,N_6119,N_6238);
or U6686 (N_6686,N_6421,N_6106);
or U6687 (N_6687,N_6422,N_6058);
nor U6688 (N_6688,N_6495,N_6266);
nand U6689 (N_6689,N_6385,N_6483);
and U6690 (N_6690,N_6190,N_6391);
and U6691 (N_6691,N_6341,N_6193);
nand U6692 (N_6692,N_6301,N_6459);
or U6693 (N_6693,N_6231,N_6090);
nor U6694 (N_6694,N_6196,N_6115);
nor U6695 (N_6695,N_6428,N_6255);
and U6696 (N_6696,N_6241,N_6351);
nand U6697 (N_6697,N_6237,N_6162);
or U6698 (N_6698,N_6397,N_6081);
xor U6699 (N_6699,N_6008,N_6454);
and U6700 (N_6700,N_6195,N_6402);
xor U6701 (N_6701,N_6345,N_6343);
nor U6702 (N_6702,N_6444,N_6062);
nand U6703 (N_6703,N_6153,N_6321);
or U6704 (N_6704,N_6134,N_6157);
or U6705 (N_6705,N_6025,N_6100);
xnor U6706 (N_6706,N_6437,N_6075);
or U6707 (N_6707,N_6046,N_6024);
nor U6708 (N_6708,N_6417,N_6149);
and U6709 (N_6709,N_6084,N_6344);
and U6710 (N_6710,N_6072,N_6122);
and U6711 (N_6711,N_6037,N_6174);
xor U6712 (N_6712,N_6036,N_6346);
and U6713 (N_6713,N_6164,N_6382);
nor U6714 (N_6714,N_6154,N_6471);
and U6715 (N_6715,N_6160,N_6056);
nand U6716 (N_6716,N_6319,N_6335);
nor U6717 (N_6717,N_6490,N_6409);
or U6718 (N_6718,N_6275,N_6429);
nand U6719 (N_6719,N_6413,N_6187);
or U6720 (N_6720,N_6472,N_6212);
and U6721 (N_6721,N_6323,N_6070);
nand U6722 (N_6722,N_6214,N_6018);
and U6723 (N_6723,N_6096,N_6083);
nor U6724 (N_6724,N_6211,N_6105);
or U6725 (N_6725,N_6005,N_6387);
nand U6726 (N_6726,N_6332,N_6135);
xnor U6727 (N_6727,N_6393,N_6189);
nor U6728 (N_6728,N_6354,N_6016);
or U6729 (N_6729,N_6156,N_6132);
and U6730 (N_6730,N_6178,N_6317);
nor U6731 (N_6731,N_6243,N_6144);
and U6732 (N_6732,N_6412,N_6497);
or U6733 (N_6733,N_6221,N_6172);
xnor U6734 (N_6734,N_6102,N_6377);
xnor U6735 (N_6735,N_6043,N_6369);
xor U6736 (N_6736,N_6077,N_6386);
or U6737 (N_6737,N_6061,N_6217);
or U6738 (N_6738,N_6493,N_6276);
nand U6739 (N_6739,N_6390,N_6089);
or U6740 (N_6740,N_6158,N_6251);
nand U6741 (N_6741,N_6407,N_6006);
nor U6742 (N_6742,N_6063,N_6449);
nor U6743 (N_6743,N_6274,N_6347);
and U6744 (N_6744,N_6380,N_6003);
or U6745 (N_6745,N_6389,N_6261);
nand U6746 (N_6746,N_6104,N_6496);
and U6747 (N_6747,N_6142,N_6399);
nor U6748 (N_6748,N_6176,N_6467);
xor U6749 (N_6749,N_6337,N_6095);
and U6750 (N_6750,N_6160,N_6023);
or U6751 (N_6751,N_6276,N_6274);
nor U6752 (N_6752,N_6325,N_6262);
and U6753 (N_6753,N_6036,N_6347);
and U6754 (N_6754,N_6199,N_6361);
or U6755 (N_6755,N_6452,N_6014);
nand U6756 (N_6756,N_6203,N_6027);
and U6757 (N_6757,N_6109,N_6418);
and U6758 (N_6758,N_6330,N_6113);
xnor U6759 (N_6759,N_6389,N_6412);
nor U6760 (N_6760,N_6386,N_6202);
xor U6761 (N_6761,N_6212,N_6434);
xor U6762 (N_6762,N_6482,N_6087);
and U6763 (N_6763,N_6155,N_6498);
nand U6764 (N_6764,N_6189,N_6039);
nand U6765 (N_6765,N_6003,N_6118);
nand U6766 (N_6766,N_6366,N_6131);
and U6767 (N_6767,N_6075,N_6324);
and U6768 (N_6768,N_6104,N_6388);
nor U6769 (N_6769,N_6192,N_6361);
nor U6770 (N_6770,N_6063,N_6019);
or U6771 (N_6771,N_6122,N_6272);
or U6772 (N_6772,N_6439,N_6360);
nor U6773 (N_6773,N_6472,N_6281);
xnor U6774 (N_6774,N_6076,N_6053);
xor U6775 (N_6775,N_6199,N_6140);
and U6776 (N_6776,N_6045,N_6135);
xnor U6777 (N_6777,N_6210,N_6475);
nand U6778 (N_6778,N_6184,N_6131);
or U6779 (N_6779,N_6222,N_6022);
nand U6780 (N_6780,N_6171,N_6189);
xor U6781 (N_6781,N_6493,N_6475);
and U6782 (N_6782,N_6018,N_6380);
nand U6783 (N_6783,N_6268,N_6144);
or U6784 (N_6784,N_6208,N_6224);
xnor U6785 (N_6785,N_6194,N_6160);
nand U6786 (N_6786,N_6107,N_6461);
nor U6787 (N_6787,N_6268,N_6079);
nor U6788 (N_6788,N_6478,N_6098);
xor U6789 (N_6789,N_6275,N_6079);
or U6790 (N_6790,N_6095,N_6443);
nand U6791 (N_6791,N_6113,N_6123);
nor U6792 (N_6792,N_6262,N_6205);
xnor U6793 (N_6793,N_6363,N_6351);
nand U6794 (N_6794,N_6449,N_6339);
xnor U6795 (N_6795,N_6151,N_6390);
or U6796 (N_6796,N_6086,N_6229);
or U6797 (N_6797,N_6070,N_6218);
xor U6798 (N_6798,N_6091,N_6330);
xnor U6799 (N_6799,N_6324,N_6306);
nand U6800 (N_6800,N_6174,N_6339);
nand U6801 (N_6801,N_6362,N_6186);
or U6802 (N_6802,N_6238,N_6191);
xnor U6803 (N_6803,N_6105,N_6018);
or U6804 (N_6804,N_6166,N_6287);
xnor U6805 (N_6805,N_6031,N_6386);
nor U6806 (N_6806,N_6097,N_6456);
and U6807 (N_6807,N_6173,N_6233);
nor U6808 (N_6808,N_6324,N_6422);
and U6809 (N_6809,N_6355,N_6499);
nand U6810 (N_6810,N_6397,N_6312);
and U6811 (N_6811,N_6232,N_6459);
nand U6812 (N_6812,N_6254,N_6499);
nand U6813 (N_6813,N_6361,N_6446);
or U6814 (N_6814,N_6325,N_6294);
xnor U6815 (N_6815,N_6423,N_6036);
xnor U6816 (N_6816,N_6397,N_6430);
xnor U6817 (N_6817,N_6417,N_6057);
xnor U6818 (N_6818,N_6375,N_6018);
xnor U6819 (N_6819,N_6155,N_6399);
and U6820 (N_6820,N_6025,N_6436);
and U6821 (N_6821,N_6154,N_6067);
and U6822 (N_6822,N_6428,N_6085);
nor U6823 (N_6823,N_6125,N_6277);
xnor U6824 (N_6824,N_6065,N_6057);
and U6825 (N_6825,N_6023,N_6045);
xnor U6826 (N_6826,N_6338,N_6397);
xnor U6827 (N_6827,N_6303,N_6232);
xor U6828 (N_6828,N_6380,N_6136);
xor U6829 (N_6829,N_6075,N_6287);
nor U6830 (N_6830,N_6371,N_6185);
nor U6831 (N_6831,N_6059,N_6323);
nand U6832 (N_6832,N_6027,N_6418);
nor U6833 (N_6833,N_6282,N_6002);
xnor U6834 (N_6834,N_6362,N_6382);
and U6835 (N_6835,N_6188,N_6008);
nand U6836 (N_6836,N_6068,N_6062);
or U6837 (N_6837,N_6431,N_6430);
nand U6838 (N_6838,N_6471,N_6008);
nor U6839 (N_6839,N_6394,N_6223);
nor U6840 (N_6840,N_6403,N_6351);
xnor U6841 (N_6841,N_6389,N_6073);
and U6842 (N_6842,N_6168,N_6001);
xor U6843 (N_6843,N_6204,N_6161);
nand U6844 (N_6844,N_6327,N_6104);
or U6845 (N_6845,N_6403,N_6360);
nand U6846 (N_6846,N_6195,N_6166);
nor U6847 (N_6847,N_6444,N_6306);
or U6848 (N_6848,N_6058,N_6114);
nand U6849 (N_6849,N_6201,N_6451);
or U6850 (N_6850,N_6494,N_6453);
xnor U6851 (N_6851,N_6174,N_6412);
xnor U6852 (N_6852,N_6016,N_6477);
xor U6853 (N_6853,N_6323,N_6098);
and U6854 (N_6854,N_6000,N_6173);
nand U6855 (N_6855,N_6314,N_6105);
or U6856 (N_6856,N_6237,N_6286);
nor U6857 (N_6857,N_6133,N_6275);
or U6858 (N_6858,N_6333,N_6215);
xnor U6859 (N_6859,N_6291,N_6472);
and U6860 (N_6860,N_6347,N_6435);
or U6861 (N_6861,N_6453,N_6471);
nand U6862 (N_6862,N_6331,N_6236);
and U6863 (N_6863,N_6026,N_6299);
or U6864 (N_6864,N_6113,N_6073);
xnor U6865 (N_6865,N_6179,N_6498);
or U6866 (N_6866,N_6327,N_6289);
and U6867 (N_6867,N_6447,N_6055);
xor U6868 (N_6868,N_6183,N_6353);
and U6869 (N_6869,N_6430,N_6051);
xor U6870 (N_6870,N_6290,N_6132);
or U6871 (N_6871,N_6082,N_6170);
xnor U6872 (N_6872,N_6261,N_6290);
nor U6873 (N_6873,N_6326,N_6465);
or U6874 (N_6874,N_6076,N_6049);
nand U6875 (N_6875,N_6229,N_6247);
and U6876 (N_6876,N_6496,N_6417);
nand U6877 (N_6877,N_6414,N_6105);
nor U6878 (N_6878,N_6136,N_6261);
or U6879 (N_6879,N_6376,N_6177);
nor U6880 (N_6880,N_6431,N_6124);
and U6881 (N_6881,N_6360,N_6050);
and U6882 (N_6882,N_6109,N_6308);
or U6883 (N_6883,N_6196,N_6298);
and U6884 (N_6884,N_6267,N_6026);
xnor U6885 (N_6885,N_6185,N_6492);
nor U6886 (N_6886,N_6160,N_6053);
nand U6887 (N_6887,N_6059,N_6251);
and U6888 (N_6888,N_6357,N_6312);
xnor U6889 (N_6889,N_6278,N_6034);
xnor U6890 (N_6890,N_6414,N_6088);
xnor U6891 (N_6891,N_6151,N_6110);
nor U6892 (N_6892,N_6087,N_6133);
nand U6893 (N_6893,N_6330,N_6274);
xor U6894 (N_6894,N_6405,N_6400);
nor U6895 (N_6895,N_6043,N_6295);
and U6896 (N_6896,N_6430,N_6470);
xor U6897 (N_6897,N_6101,N_6453);
xor U6898 (N_6898,N_6364,N_6158);
nor U6899 (N_6899,N_6322,N_6191);
nand U6900 (N_6900,N_6054,N_6035);
nor U6901 (N_6901,N_6239,N_6185);
nand U6902 (N_6902,N_6184,N_6414);
xnor U6903 (N_6903,N_6344,N_6470);
and U6904 (N_6904,N_6003,N_6134);
or U6905 (N_6905,N_6418,N_6441);
nor U6906 (N_6906,N_6165,N_6415);
nor U6907 (N_6907,N_6202,N_6076);
or U6908 (N_6908,N_6080,N_6361);
xnor U6909 (N_6909,N_6322,N_6211);
or U6910 (N_6910,N_6286,N_6373);
and U6911 (N_6911,N_6293,N_6401);
and U6912 (N_6912,N_6181,N_6150);
nand U6913 (N_6913,N_6011,N_6039);
or U6914 (N_6914,N_6314,N_6116);
or U6915 (N_6915,N_6348,N_6046);
or U6916 (N_6916,N_6307,N_6113);
xnor U6917 (N_6917,N_6339,N_6133);
nor U6918 (N_6918,N_6153,N_6309);
nand U6919 (N_6919,N_6444,N_6128);
or U6920 (N_6920,N_6496,N_6163);
or U6921 (N_6921,N_6048,N_6058);
nand U6922 (N_6922,N_6313,N_6116);
xnor U6923 (N_6923,N_6459,N_6478);
xor U6924 (N_6924,N_6438,N_6494);
nor U6925 (N_6925,N_6484,N_6198);
nand U6926 (N_6926,N_6392,N_6494);
and U6927 (N_6927,N_6049,N_6278);
xor U6928 (N_6928,N_6189,N_6255);
xnor U6929 (N_6929,N_6225,N_6256);
or U6930 (N_6930,N_6391,N_6477);
or U6931 (N_6931,N_6015,N_6250);
nor U6932 (N_6932,N_6391,N_6396);
nand U6933 (N_6933,N_6467,N_6215);
nor U6934 (N_6934,N_6472,N_6443);
nor U6935 (N_6935,N_6485,N_6402);
or U6936 (N_6936,N_6010,N_6092);
and U6937 (N_6937,N_6427,N_6364);
nor U6938 (N_6938,N_6138,N_6131);
xnor U6939 (N_6939,N_6341,N_6121);
nand U6940 (N_6940,N_6106,N_6197);
and U6941 (N_6941,N_6157,N_6340);
xor U6942 (N_6942,N_6134,N_6427);
or U6943 (N_6943,N_6285,N_6091);
xor U6944 (N_6944,N_6123,N_6313);
nor U6945 (N_6945,N_6282,N_6411);
xor U6946 (N_6946,N_6317,N_6017);
nand U6947 (N_6947,N_6406,N_6220);
nand U6948 (N_6948,N_6272,N_6409);
or U6949 (N_6949,N_6414,N_6249);
nor U6950 (N_6950,N_6487,N_6168);
nand U6951 (N_6951,N_6174,N_6125);
xnor U6952 (N_6952,N_6015,N_6170);
xnor U6953 (N_6953,N_6450,N_6014);
nor U6954 (N_6954,N_6146,N_6087);
and U6955 (N_6955,N_6034,N_6487);
nor U6956 (N_6956,N_6499,N_6197);
or U6957 (N_6957,N_6450,N_6454);
nor U6958 (N_6958,N_6140,N_6097);
nand U6959 (N_6959,N_6242,N_6270);
and U6960 (N_6960,N_6228,N_6491);
nand U6961 (N_6961,N_6194,N_6462);
nor U6962 (N_6962,N_6427,N_6337);
or U6963 (N_6963,N_6377,N_6407);
and U6964 (N_6964,N_6054,N_6469);
nor U6965 (N_6965,N_6479,N_6158);
xnor U6966 (N_6966,N_6291,N_6487);
and U6967 (N_6967,N_6178,N_6314);
and U6968 (N_6968,N_6491,N_6238);
nor U6969 (N_6969,N_6114,N_6199);
and U6970 (N_6970,N_6023,N_6335);
or U6971 (N_6971,N_6397,N_6254);
nand U6972 (N_6972,N_6048,N_6474);
or U6973 (N_6973,N_6225,N_6448);
xor U6974 (N_6974,N_6254,N_6493);
and U6975 (N_6975,N_6101,N_6223);
nand U6976 (N_6976,N_6334,N_6114);
and U6977 (N_6977,N_6409,N_6027);
nand U6978 (N_6978,N_6068,N_6152);
nor U6979 (N_6979,N_6221,N_6087);
or U6980 (N_6980,N_6325,N_6338);
and U6981 (N_6981,N_6062,N_6204);
xnor U6982 (N_6982,N_6278,N_6197);
xor U6983 (N_6983,N_6390,N_6349);
xnor U6984 (N_6984,N_6152,N_6386);
or U6985 (N_6985,N_6239,N_6271);
nand U6986 (N_6986,N_6030,N_6486);
nand U6987 (N_6987,N_6310,N_6211);
nor U6988 (N_6988,N_6275,N_6236);
nor U6989 (N_6989,N_6406,N_6035);
nor U6990 (N_6990,N_6471,N_6226);
nor U6991 (N_6991,N_6358,N_6322);
or U6992 (N_6992,N_6187,N_6242);
or U6993 (N_6993,N_6055,N_6398);
xnor U6994 (N_6994,N_6339,N_6329);
nor U6995 (N_6995,N_6481,N_6416);
or U6996 (N_6996,N_6429,N_6034);
and U6997 (N_6997,N_6043,N_6438);
or U6998 (N_6998,N_6470,N_6320);
and U6999 (N_6999,N_6250,N_6233);
or U7000 (N_7000,N_6703,N_6636);
xnor U7001 (N_7001,N_6578,N_6801);
nor U7002 (N_7002,N_6978,N_6585);
and U7003 (N_7003,N_6524,N_6822);
nand U7004 (N_7004,N_6715,N_6544);
or U7005 (N_7005,N_6571,N_6840);
or U7006 (N_7006,N_6883,N_6714);
xor U7007 (N_7007,N_6958,N_6873);
nor U7008 (N_7008,N_6891,N_6887);
nor U7009 (N_7009,N_6751,N_6541);
or U7010 (N_7010,N_6909,N_6825);
xnor U7011 (N_7011,N_6760,N_6640);
or U7012 (N_7012,N_6834,N_6947);
or U7013 (N_7013,N_6599,N_6737);
nand U7014 (N_7014,N_6881,N_6786);
nand U7015 (N_7015,N_6955,N_6692);
and U7016 (N_7016,N_6964,N_6895);
or U7017 (N_7017,N_6682,N_6773);
nor U7018 (N_7018,N_6613,N_6654);
or U7019 (N_7019,N_6962,N_6506);
xnor U7020 (N_7020,N_6618,N_6897);
or U7021 (N_7021,N_6904,N_6648);
nor U7022 (N_7022,N_6960,N_6752);
nor U7023 (N_7023,N_6782,N_6531);
xor U7024 (N_7024,N_6713,N_6527);
xor U7025 (N_7025,N_6522,N_6543);
and U7026 (N_7026,N_6770,N_6756);
xor U7027 (N_7027,N_6923,N_6879);
nand U7028 (N_7028,N_6707,N_6681);
xor U7029 (N_7029,N_6719,N_6623);
nand U7030 (N_7030,N_6657,N_6573);
or U7031 (N_7031,N_6753,N_6979);
or U7032 (N_7032,N_6841,N_6547);
or U7033 (N_7033,N_6984,N_6675);
nor U7034 (N_7034,N_6507,N_6846);
nor U7035 (N_7035,N_6723,N_6575);
or U7036 (N_7036,N_6804,N_6565);
xor U7037 (N_7037,N_6669,N_6679);
nand U7038 (N_7038,N_6534,N_6742);
and U7039 (N_7039,N_6503,N_6918);
xnor U7040 (N_7040,N_6561,N_6929);
and U7041 (N_7041,N_6901,N_6845);
nor U7042 (N_7042,N_6582,N_6676);
xor U7043 (N_7043,N_6866,N_6624);
and U7044 (N_7044,N_6698,N_6589);
or U7045 (N_7045,N_6560,N_6766);
nand U7046 (N_7046,N_6593,N_6763);
nand U7047 (N_7047,N_6793,N_6646);
or U7048 (N_7048,N_6596,N_6982);
nand U7049 (N_7049,N_6789,N_6937);
nand U7050 (N_7050,N_6933,N_6849);
or U7051 (N_7051,N_6584,N_6944);
nand U7052 (N_7052,N_6548,N_6678);
nand U7053 (N_7053,N_6890,N_6819);
nor U7054 (N_7054,N_6919,N_6581);
and U7055 (N_7055,N_6748,N_6806);
and U7056 (N_7056,N_6725,N_6871);
nand U7057 (N_7057,N_6671,N_6739);
and U7058 (N_7058,N_6785,N_6829);
or U7059 (N_7059,N_6975,N_6647);
xor U7060 (N_7060,N_6729,N_6610);
nor U7061 (N_7061,N_6824,N_6608);
nand U7062 (N_7062,N_6781,N_6970);
xnor U7063 (N_7063,N_6969,N_6697);
nand U7064 (N_7064,N_6882,N_6519);
xor U7065 (N_7065,N_6855,N_6712);
nand U7066 (N_7066,N_6907,N_6949);
and U7067 (N_7067,N_6888,N_6562);
xnor U7068 (N_7068,N_6985,N_6911);
nand U7069 (N_7069,N_6780,N_6996);
xor U7070 (N_7070,N_6659,N_6701);
xnor U7071 (N_7071,N_6778,N_6501);
or U7072 (N_7072,N_6717,N_6761);
xnor U7073 (N_7073,N_6835,N_6792);
and U7074 (N_7074,N_6848,N_6622);
nand U7075 (N_7075,N_6833,N_6767);
or U7076 (N_7076,N_6759,N_6579);
and U7077 (N_7077,N_6971,N_6851);
nor U7078 (N_7078,N_6880,N_6699);
and U7079 (N_7079,N_6619,N_6774);
nand U7080 (N_7080,N_6798,N_6525);
or U7081 (N_7081,N_6661,N_6950);
or U7082 (N_7082,N_6569,N_6885);
or U7083 (N_7083,N_6511,N_6722);
xnor U7084 (N_7084,N_6651,N_6931);
or U7085 (N_7085,N_6914,N_6601);
and U7086 (N_7086,N_6521,N_6667);
nand U7087 (N_7087,N_6546,N_6728);
or U7088 (N_7088,N_6831,N_6586);
and U7089 (N_7089,N_6554,N_6516);
or U7090 (N_7090,N_6857,N_6607);
nor U7091 (N_7091,N_6966,N_6754);
xnor U7092 (N_7092,N_6852,N_6746);
nor U7093 (N_7093,N_6967,N_6614);
nand U7094 (N_7094,N_6594,N_6952);
xor U7095 (N_7095,N_6989,N_6685);
nand U7096 (N_7096,N_6652,N_6802);
xnor U7097 (N_7097,N_6734,N_6745);
and U7098 (N_7098,N_6595,N_6823);
xor U7099 (N_7099,N_6764,N_6942);
and U7100 (N_7100,N_6509,N_6830);
and U7101 (N_7101,N_6686,N_6807);
nor U7102 (N_7102,N_6539,N_6794);
nand U7103 (N_7103,N_6542,N_6872);
xnor U7104 (N_7104,N_6644,N_6862);
nand U7105 (N_7105,N_6791,N_6821);
nand U7106 (N_7106,N_6615,N_6653);
nand U7107 (N_7107,N_6627,N_6532);
nor U7108 (N_7108,N_6567,N_6708);
or U7109 (N_7109,N_6917,N_6924);
xnor U7110 (N_7110,N_6617,N_6634);
nor U7111 (N_7111,N_6765,N_6788);
nand U7112 (N_7112,N_6564,N_6721);
and U7113 (N_7113,N_6726,N_6787);
xor U7114 (N_7114,N_6743,N_6656);
nor U7115 (N_7115,N_6811,N_6994);
and U7116 (N_7116,N_6662,N_6514);
and U7117 (N_7117,N_6987,N_6592);
and U7118 (N_7118,N_6616,N_6858);
nand U7119 (N_7119,N_6702,N_6693);
or U7120 (N_7120,N_6810,N_6817);
and U7121 (N_7121,N_6528,N_6903);
and U7122 (N_7122,N_6563,N_6672);
xnor U7123 (N_7123,N_6998,N_6876);
and U7124 (N_7124,N_6854,N_6983);
nand U7125 (N_7125,N_6570,N_6991);
or U7126 (N_7126,N_6776,N_6869);
and U7127 (N_7127,N_6666,N_6861);
xnor U7128 (N_7128,N_6733,N_6535);
xor U7129 (N_7129,N_6513,N_6859);
and U7130 (N_7130,N_6816,N_6583);
nand U7131 (N_7131,N_6938,N_6864);
nor U7132 (N_7132,N_6590,N_6916);
nor U7133 (N_7133,N_6545,N_6769);
or U7134 (N_7134,N_6797,N_6800);
nand U7135 (N_7135,N_6660,N_6956);
or U7136 (N_7136,N_6957,N_6850);
and U7137 (N_7137,N_6951,N_6557);
nor U7138 (N_7138,N_6899,N_6517);
or U7139 (N_7139,N_6603,N_6953);
nor U7140 (N_7140,N_6795,N_6526);
nor U7141 (N_7141,N_6588,N_6505);
or U7142 (N_7142,N_6665,N_6902);
nand U7143 (N_7143,N_6691,N_6632);
or U7144 (N_7144,N_6894,N_6577);
or U7145 (N_7145,N_6755,N_6921);
nand U7146 (N_7146,N_6626,N_6920);
and U7147 (N_7147,N_6633,N_6696);
xor U7148 (N_7148,N_6735,N_6597);
nor U7149 (N_7149,N_6889,N_6520);
and U7150 (N_7150,N_6912,N_6689);
xnor U7151 (N_7151,N_6551,N_6510);
xnor U7152 (N_7152,N_6684,N_6604);
or U7153 (N_7153,N_6620,N_6680);
nor U7154 (N_7154,N_6915,N_6943);
or U7155 (N_7155,N_6762,N_6538);
xnor U7156 (N_7156,N_6731,N_6704);
nand U7157 (N_7157,N_6867,N_6783);
nor U7158 (N_7158,N_6736,N_6948);
or U7159 (N_7159,N_6856,N_6874);
or U7160 (N_7160,N_6980,N_6658);
nand U7161 (N_7161,N_6504,N_6572);
nand U7162 (N_7162,N_6677,N_6965);
nor U7163 (N_7163,N_6939,N_6927);
nand U7164 (N_7164,N_6803,N_6740);
nor U7165 (N_7165,N_6536,N_6598);
nor U7166 (N_7166,N_6668,N_6805);
or U7167 (N_7167,N_6629,N_6673);
nor U7168 (N_7168,N_6941,N_6533);
nand U7169 (N_7169,N_6818,N_6730);
or U7170 (N_7170,N_6606,N_6772);
nand U7171 (N_7171,N_6625,N_6995);
nor U7172 (N_7172,N_6683,N_6757);
xor U7173 (N_7173,N_6968,N_6580);
xnor U7174 (N_7174,N_6976,N_6959);
or U7175 (N_7175,N_6926,N_6946);
and U7176 (N_7176,N_6518,N_6973);
or U7177 (N_7177,N_6552,N_6630);
and U7178 (N_7178,N_6591,N_6609);
and U7179 (N_7179,N_6724,N_6986);
nor U7180 (N_7180,N_6934,N_6650);
nand U7181 (N_7181,N_6537,N_6643);
nor U7182 (N_7182,N_6670,N_6963);
and U7183 (N_7183,N_6977,N_6711);
nand U7184 (N_7184,N_6945,N_6928);
nor U7185 (N_7185,N_6777,N_6710);
nor U7186 (N_7186,N_6906,N_6508);
or U7187 (N_7187,N_6555,N_6940);
or U7188 (N_7188,N_6700,N_6576);
and U7189 (N_7189,N_6796,N_6512);
nand U7190 (N_7190,N_6893,N_6898);
or U7191 (N_7191,N_6771,N_6992);
xor U7192 (N_7192,N_6635,N_6529);
xor U7193 (N_7193,N_6974,N_6843);
nor U7194 (N_7194,N_6611,N_6875);
xor U7195 (N_7195,N_6566,N_6990);
nor U7196 (N_7196,N_6837,N_6706);
nand U7197 (N_7197,N_6972,N_6663);
xnor U7198 (N_7198,N_6500,N_6925);
nand U7199 (N_7199,N_6910,N_6844);
nand U7200 (N_7200,N_6808,N_6727);
nor U7201 (N_7201,N_6768,N_6997);
nor U7202 (N_7202,N_6558,N_6688);
or U7203 (N_7203,N_6775,N_6639);
nand U7204 (N_7204,N_6877,N_6905);
nor U7205 (N_7205,N_6574,N_6605);
nand U7206 (N_7206,N_6587,N_6799);
or U7207 (N_7207,N_6813,N_6687);
xor U7208 (N_7208,N_6655,N_6961);
xor U7209 (N_7209,N_6884,N_6935);
or U7210 (N_7210,N_6865,N_6988);
nand U7211 (N_7211,N_6559,N_6838);
and U7212 (N_7212,N_6863,N_6853);
or U7213 (N_7213,N_6540,N_6870);
nand U7214 (N_7214,N_6621,N_6999);
or U7215 (N_7215,N_6720,N_6842);
and U7216 (N_7216,N_6832,N_6674);
nor U7217 (N_7217,N_6826,N_6758);
and U7218 (N_7218,N_6913,N_6641);
and U7219 (N_7219,N_6809,N_6820);
xnor U7220 (N_7220,N_6502,N_6900);
nor U7221 (N_7221,N_6645,N_6836);
nand U7222 (N_7222,N_6738,N_6550);
nand U7223 (N_7223,N_6690,N_6549);
xor U7224 (N_7224,N_6922,N_6628);
nand U7225 (N_7225,N_6839,N_6930);
nand U7226 (N_7226,N_6908,N_6530);
and U7227 (N_7227,N_6612,N_6936);
nor U7228 (N_7228,N_6790,N_6718);
xnor U7229 (N_7229,N_6812,N_6815);
nor U7230 (N_7230,N_6732,N_6827);
nor U7231 (N_7231,N_6892,N_6705);
or U7232 (N_7232,N_6932,N_6878);
nor U7233 (N_7233,N_6602,N_6814);
or U7234 (N_7234,N_6828,N_6868);
nor U7235 (N_7235,N_6784,N_6695);
or U7236 (N_7236,N_6631,N_6860);
nor U7237 (N_7237,N_6709,N_6600);
or U7238 (N_7238,N_6664,N_6749);
nand U7239 (N_7239,N_6954,N_6847);
nor U7240 (N_7240,N_6981,N_6694);
and U7241 (N_7241,N_6716,N_6741);
and U7242 (N_7242,N_6779,N_6637);
xnor U7243 (N_7243,N_6886,N_6556);
nor U7244 (N_7244,N_6642,N_6993);
xnor U7245 (N_7245,N_6750,N_6638);
or U7246 (N_7246,N_6896,N_6553);
nand U7247 (N_7247,N_6744,N_6515);
and U7248 (N_7248,N_6568,N_6649);
nand U7249 (N_7249,N_6523,N_6747);
nand U7250 (N_7250,N_6702,N_6503);
xor U7251 (N_7251,N_6581,N_6589);
or U7252 (N_7252,N_6858,N_6961);
nand U7253 (N_7253,N_6582,N_6760);
nor U7254 (N_7254,N_6747,N_6783);
nand U7255 (N_7255,N_6837,N_6937);
nand U7256 (N_7256,N_6538,N_6955);
and U7257 (N_7257,N_6868,N_6759);
and U7258 (N_7258,N_6686,N_6961);
nand U7259 (N_7259,N_6937,N_6773);
nand U7260 (N_7260,N_6744,N_6653);
xnor U7261 (N_7261,N_6573,N_6991);
and U7262 (N_7262,N_6960,N_6808);
nand U7263 (N_7263,N_6798,N_6814);
and U7264 (N_7264,N_6569,N_6719);
nor U7265 (N_7265,N_6879,N_6880);
and U7266 (N_7266,N_6558,N_6581);
xnor U7267 (N_7267,N_6505,N_6826);
xnor U7268 (N_7268,N_6505,N_6926);
xnor U7269 (N_7269,N_6529,N_6956);
or U7270 (N_7270,N_6698,N_6815);
nand U7271 (N_7271,N_6918,N_6959);
nor U7272 (N_7272,N_6720,N_6965);
xor U7273 (N_7273,N_6977,N_6982);
and U7274 (N_7274,N_6787,N_6503);
xnor U7275 (N_7275,N_6545,N_6549);
nand U7276 (N_7276,N_6553,N_6950);
or U7277 (N_7277,N_6690,N_6539);
and U7278 (N_7278,N_6946,N_6762);
nor U7279 (N_7279,N_6796,N_6990);
or U7280 (N_7280,N_6702,N_6711);
nor U7281 (N_7281,N_6743,N_6842);
xor U7282 (N_7282,N_6567,N_6879);
or U7283 (N_7283,N_6605,N_6791);
or U7284 (N_7284,N_6666,N_6615);
and U7285 (N_7285,N_6753,N_6823);
nand U7286 (N_7286,N_6577,N_6647);
nor U7287 (N_7287,N_6611,N_6647);
and U7288 (N_7288,N_6616,N_6940);
or U7289 (N_7289,N_6626,N_6586);
xnor U7290 (N_7290,N_6652,N_6670);
xnor U7291 (N_7291,N_6720,N_6794);
nand U7292 (N_7292,N_6647,N_6850);
nor U7293 (N_7293,N_6688,N_6925);
nand U7294 (N_7294,N_6916,N_6554);
nand U7295 (N_7295,N_6722,N_6914);
and U7296 (N_7296,N_6515,N_6774);
or U7297 (N_7297,N_6970,N_6617);
or U7298 (N_7298,N_6514,N_6671);
or U7299 (N_7299,N_6792,N_6913);
nand U7300 (N_7300,N_6810,N_6580);
nand U7301 (N_7301,N_6534,N_6815);
or U7302 (N_7302,N_6693,N_6914);
nand U7303 (N_7303,N_6993,N_6802);
or U7304 (N_7304,N_6773,N_6994);
nand U7305 (N_7305,N_6726,N_6651);
xnor U7306 (N_7306,N_6869,N_6805);
nand U7307 (N_7307,N_6940,N_6759);
and U7308 (N_7308,N_6512,N_6572);
nand U7309 (N_7309,N_6790,N_6944);
or U7310 (N_7310,N_6935,N_6655);
or U7311 (N_7311,N_6684,N_6808);
xor U7312 (N_7312,N_6724,N_6723);
xor U7313 (N_7313,N_6857,N_6822);
nor U7314 (N_7314,N_6568,N_6583);
and U7315 (N_7315,N_6888,N_6589);
nand U7316 (N_7316,N_6692,N_6972);
and U7317 (N_7317,N_6888,N_6834);
or U7318 (N_7318,N_6613,N_6739);
and U7319 (N_7319,N_6845,N_6847);
nand U7320 (N_7320,N_6867,N_6820);
nor U7321 (N_7321,N_6855,N_6555);
nor U7322 (N_7322,N_6537,N_6869);
nor U7323 (N_7323,N_6827,N_6557);
nor U7324 (N_7324,N_6911,N_6710);
or U7325 (N_7325,N_6868,N_6591);
or U7326 (N_7326,N_6717,N_6578);
and U7327 (N_7327,N_6725,N_6836);
nand U7328 (N_7328,N_6507,N_6634);
xor U7329 (N_7329,N_6576,N_6880);
nor U7330 (N_7330,N_6965,N_6502);
xnor U7331 (N_7331,N_6863,N_6619);
nor U7332 (N_7332,N_6782,N_6680);
xnor U7333 (N_7333,N_6721,N_6863);
xor U7334 (N_7334,N_6587,N_6597);
xor U7335 (N_7335,N_6508,N_6541);
nor U7336 (N_7336,N_6755,N_6694);
nor U7337 (N_7337,N_6759,N_6979);
nand U7338 (N_7338,N_6751,N_6765);
nand U7339 (N_7339,N_6748,N_6975);
nor U7340 (N_7340,N_6543,N_6546);
nand U7341 (N_7341,N_6979,N_6714);
or U7342 (N_7342,N_6689,N_6878);
and U7343 (N_7343,N_6603,N_6976);
nor U7344 (N_7344,N_6873,N_6600);
or U7345 (N_7345,N_6604,N_6519);
nand U7346 (N_7346,N_6957,N_6750);
xnor U7347 (N_7347,N_6853,N_6588);
or U7348 (N_7348,N_6918,N_6755);
nor U7349 (N_7349,N_6755,N_6648);
nor U7350 (N_7350,N_6868,N_6531);
nor U7351 (N_7351,N_6950,N_6610);
nor U7352 (N_7352,N_6655,N_6673);
xnor U7353 (N_7353,N_6969,N_6993);
and U7354 (N_7354,N_6853,N_6856);
and U7355 (N_7355,N_6768,N_6507);
xnor U7356 (N_7356,N_6736,N_6917);
nand U7357 (N_7357,N_6554,N_6642);
or U7358 (N_7358,N_6764,N_6509);
nor U7359 (N_7359,N_6798,N_6559);
or U7360 (N_7360,N_6514,N_6713);
nand U7361 (N_7361,N_6929,N_6739);
nor U7362 (N_7362,N_6865,N_6515);
xor U7363 (N_7363,N_6766,N_6509);
or U7364 (N_7364,N_6640,N_6988);
nand U7365 (N_7365,N_6759,N_6982);
or U7366 (N_7366,N_6508,N_6847);
and U7367 (N_7367,N_6778,N_6653);
nand U7368 (N_7368,N_6575,N_6738);
nor U7369 (N_7369,N_6734,N_6835);
and U7370 (N_7370,N_6678,N_6823);
xnor U7371 (N_7371,N_6953,N_6672);
xnor U7372 (N_7372,N_6729,N_6879);
nor U7373 (N_7373,N_6688,N_6505);
nor U7374 (N_7374,N_6554,N_6830);
or U7375 (N_7375,N_6526,N_6567);
xor U7376 (N_7376,N_6982,N_6720);
or U7377 (N_7377,N_6859,N_6686);
and U7378 (N_7378,N_6682,N_6956);
nand U7379 (N_7379,N_6725,N_6581);
or U7380 (N_7380,N_6586,N_6862);
or U7381 (N_7381,N_6925,N_6706);
nand U7382 (N_7382,N_6761,N_6773);
xnor U7383 (N_7383,N_6509,N_6575);
and U7384 (N_7384,N_6950,N_6990);
and U7385 (N_7385,N_6637,N_6880);
nor U7386 (N_7386,N_6686,N_6760);
nand U7387 (N_7387,N_6878,N_6595);
and U7388 (N_7388,N_6981,N_6696);
nor U7389 (N_7389,N_6721,N_6967);
or U7390 (N_7390,N_6648,N_6683);
and U7391 (N_7391,N_6915,N_6668);
nor U7392 (N_7392,N_6592,N_6985);
nor U7393 (N_7393,N_6891,N_6781);
nand U7394 (N_7394,N_6955,N_6699);
nor U7395 (N_7395,N_6564,N_6971);
nand U7396 (N_7396,N_6777,N_6671);
xnor U7397 (N_7397,N_6630,N_6612);
and U7398 (N_7398,N_6895,N_6632);
and U7399 (N_7399,N_6537,N_6903);
nor U7400 (N_7400,N_6591,N_6521);
nand U7401 (N_7401,N_6859,N_6922);
nand U7402 (N_7402,N_6690,N_6510);
nor U7403 (N_7403,N_6543,N_6922);
nor U7404 (N_7404,N_6766,N_6749);
xnor U7405 (N_7405,N_6552,N_6540);
nor U7406 (N_7406,N_6627,N_6731);
xnor U7407 (N_7407,N_6624,N_6527);
nand U7408 (N_7408,N_6927,N_6922);
or U7409 (N_7409,N_6637,N_6660);
xnor U7410 (N_7410,N_6890,N_6896);
and U7411 (N_7411,N_6943,N_6715);
xnor U7412 (N_7412,N_6877,N_6840);
nor U7413 (N_7413,N_6965,N_6928);
nand U7414 (N_7414,N_6903,N_6578);
and U7415 (N_7415,N_6957,N_6926);
xnor U7416 (N_7416,N_6552,N_6585);
nand U7417 (N_7417,N_6820,N_6614);
nor U7418 (N_7418,N_6530,N_6577);
and U7419 (N_7419,N_6764,N_6880);
nor U7420 (N_7420,N_6861,N_6637);
nand U7421 (N_7421,N_6752,N_6531);
and U7422 (N_7422,N_6790,N_6744);
or U7423 (N_7423,N_6689,N_6762);
xor U7424 (N_7424,N_6579,N_6875);
or U7425 (N_7425,N_6625,N_6905);
or U7426 (N_7426,N_6501,N_6503);
nor U7427 (N_7427,N_6962,N_6726);
or U7428 (N_7428,N_6853,N_6692);
xor U7429 (N_7429,N_6699,N_6975);
or U7430 (N_7430,N_6733,N_6879);
or U7431 (N_7431,N_6613,N_6818);
nand U7432 (N_7432,N_6691,N_6951);
xor U7433 (N_7433,N_6591,N_6757);
nor U7434 (N_7434,N_6612,N_6512);
nor U7435 (N_7435,N_6656,N_6751);
xor U7436 (N_7436,N_6636,N_6940);
xor U7437 (N_7437,N_6746,N_6931);
xnor U7438 (N_7438,N_6923,N_6565);
xnor U7439 (N_7439,N_6870,N_6839);
nor U7440 (N_7440,N_6692,N_6788);
or U7441 (N_7441,N_6519,N_6769);
or U7442 (N_7442,N_6847,N_6916);
xnor U7443 (N_7443,N_6766,N_6691);
and U7444 (N_7444,N_6977,N_6852);
and U7445 (N_7445,N_6821,N_6903);
nor U7446 (N_7446,N_6535,N_6978);
or U7447 (N_7447,N_6672,N_6833);
nor U7448 (N_7448,N_6796,N_6877);
nor U7449 (N_7449,N_6855,N_6558);
and U7450 (N_7450,N_6926,N_6885);
and U7451 (N_7451,N_6816,N_6929);
nor U7452 (N_7452,N_6961,N_6658);
nor U7453 (N_7453,N_6801,N_6674);
and U7454 (N_7454,N_6877,N_6908);
and U7455 (N_7455,N_6560,N_6746);
nand U7456 (N_7456,N_6921,N_6991);
and U7457 (N_7457,N_6634,N_6889);
nand U7458 (N_7458,N_6923,N_6556);
nor U7459 (N_7459,N_6986,N_6693);
or U7460 (N_7460,N_6659,N_6832);
and U7461 (N_7461,N_6857,N_6703);
and U7462 (N_7462,N_6796,N_6554);
xnor U7463 (N_7463,N_6638,N_6963);
or U7464 (N_7464,N_6705,N_6787);
nor U7465 (N_7465,N_6685,N_6556);
xnor U7466 (N_7466,N_6580,N_6901);
and U7467 (N_7467,N_6724,N_6775);
and U7468 (N_7468,N_6604,N_6771);
nor U7469 (N_7469,N_6509,N_6929);
and U7470 (N_7470,N_6664,N_6504);
nand U7471 (N_7471,N_6890,N_6815);
xor U7472 (N_7472,N_6722,N_6539);
nand U7473 (N_7473,N_6708,N_6912);
or U7474 (N_7474,N_6951,N_6911);
nand U7475 (N_7475,N_6614,N_6980);
or U7476 (N_7476,N_6854,N_6773);
or U7477 (N_7477,N_6794,N_6650);
nand U7478 (N_7478,N_6771,N_6709);
or U7479 (N_7479,N_6705,N_6877);
and U7480 (N_7480,N_6943,N_6755);
nor U7481 (N_7481,N_6682,N_6830);
xnor U7482 (N_7482,N_6692,N_6806);
or U7483 (N_7483,N_6812,N_6617);
and U7484 (N_7484,N_6606,N_6656);
xnor U7485 (N_7485,N_6642,N_6572);
xnor U7486 (N_7486,N_6849,N_6600);
or U7487 (N_7487,N_6650,N_6928);
nand U7488 (N_7488,N_6650,N_6867);
or U7489 (N_7489,N_6964,N_6891);
xor U7490 (N_7490,N_6561,N_6791);
nor U7491 (N_7491,N_6945,N_6522);
nand U7492 (N_7492,N_6719,N_6680);
nand U7493 (N_7493,N_6971,N_6738);
or U7494 (N_7494,N_6930,N_6561);
and U7495 (N_7495,N_6706,N_6690);
or U7496 (N_7496,N_6741,N_6985);
or U7497 (N_7497,N_6750,N_6995);
xnor U7498 (N_7498,N_6802,N_6576);
xor U7499 (N_7499,N_6611,N_6986);
or U7500 (N_7500,N_7109,N_7224);
or U7501 (N_7501,N_7152,N_7280);
and U7502 (N_7502,N_7164,N_7311);
nor U7503 (N_7503,N_7053,N_7184);
nor U7504 (N_7504,N_7299,N_7436);
xnor U7505 (N_7505,N_7340,N_7290);
and U7506 (N_7506,N_7371,N_7424);
nor U7507 (N_7507,N_7167,N_7227);
and U7508 (N_7508,N_7319,N_7172);
xnor U7509 (N_7509,N_7165,N_7293);
or U7510 (N_7510,N_7007,N_7218);
nor U7511 (N_7511,N_7325,N_7206);
nor U7512 (N_7512,N_7332,N_7470);
or U7513 (N_7513,N_7248,N_7033);
and U7514 (N_7514,N_7396,N_7479);
nand U7515 (N_7515,N_7375,N_7179);
nor U7516 (N_7516,N_7004,N_7327);
xnor U7517 (N_7517,N_7405,N_7328);
nand U7518 (N_7518,N_7409,N_7461);
or U7519 (N_7519,N_7222,N_7052);
or U7520 (N_7520,N_7485,N_7258);
nand U7521 (N_7521,N_7365,N_7130);
or U7522 (N_7522,N_7215,N_7458);
nor U7523 (N_7523,N_7068,N_7383);
and U7524 (N_7524,N_7486,N_7360);
nor U7525 (N_7525,N_7459,N_7239);
and U7526 (N_7526,N_7358,N_7372);
and U7527 (N_7527,N_7317,N_7141);
and U7528 (N_7528,N_7276,N_7469);
nor U7529 (N_7529,N_7401,N_7347);
nand U7530 (N_7530,N_7275,N_7463);
xor U7531 (N_7531,N_7450,N_7399);
nor U7532 (N_7532,N_7223,N_7140);
xor U7533 (N_7533,N_7240,N_7483);
xor U7534 (N_7534,N_7392,N_7391);
xor U7535 (N_7535,N_7185,N_7414);
and U7536 (N_7536,N_7377,N_7288);
or U7537 (N_7537,N_7342,N_7149);
or U7538 (N_7538,N_7413,N_7351);
xnor U7539 (N_7539,N_7048,N_7002);
or U7540 (N_7540,N_7335,N_7115);
nor U7541 (N_7541,N_7397,N_7416);
or U7542 (N_7542,N_7225,N_7495);
xor U7543 (N_7543,N_7482,N_7205);
and U7544 (N_7544,N_7431,N_7009);
nand U7545 (N_7545,N_7208,N_7444);
or U7546 (N_7546,N_7429,N_7013);
xnor U7547 (N_7547,N_7457,N_7281);
xnor U7548 (N_7548,N_7387,N_7354);
and U7549 (N_7549,N_7022,N_7020);
nor U7550 (N_7550,N_7092,N_7320);
nand U7551 (N_7551,N_7304,N_7237);
xor U7552 (N_7552,N_7128,N_7489);
and U7553 (N_7553,N_7419,N_7000);
or U7554 (N_7554,N_7091,N_7492);
nor U7555 (N_7555,N_7027,N_7061);
xnor U7556 (N_7556,N_7462,N_7255);
and U7557 (N_7557,N_7272,N_7267);
xnor U7558 (N_7558,N_7302,N_7361);
nand U7559 (N_7559,N_7232,N_7251);
nand U7560 (N_7560,N_7256,N_7086);
or U7561 (N_7561,N_7065,N_7193);
xor U7562 (N_7562,N_7465,N_7306);
nand U7563 (N_7563,N_7014,N_7220);
or U7564 (N_7564,N_7282,N_7199);
or U7565 (N_7565,N_7295,N_7284);
nor U7566 (N_7566,N_7338,N_7047);
nand U7567 (N_7567,N_7261,N_7379);
and U7568 (N_7568,N_7074,N_7334);
xor U7569 (N_7569,N_7161,N_7246);
and U7570 (N_7570,N_7082,N_7245);
or U7571 (N_7571,N_7169,N_7145);
or U7572 (N_7572,N_7408,N_7376);
and U7573 (N_7573,N_7430,N_7189);
nand U7574 (N_7574,N_7252,N_7034);
nor U7575 (N_7575,N_7270,N_7196);
and U7576 (N_7576,N_7229,N_7136);
nand U7577 (N_7577,N_7417,N_7072);
and U7578 (N_7578,N_7466,N_7021);
and U7579 (N_7579,N_7100,N_7129);
xnor U7580 (N_7580,N_7477,N_7207);
nor U7581 (N_7581,N_7201,N_7291);
nand U7582 (N_7582,N_7488,N_7194);
nand U7583 (N_7583,N_7312,N_7449);
nor U7584 (N_7584,N_7352,N_7031);
nand U7585 (N_7585,N_7157,N_7203);
and U7586 (N_7586,N_7118,N_7209);
xnor U7587 (N_7587,N_7353,N_7268);
nand U7588 (N_7588,N_7150,N_7238);
xnor U7589 (N_7589,N_7370,N_7442);
and U7590 (N_7590,N_7178,N_7384);
or U7591 (N_7591,N_7348,N_7487);
and U7592 (N_7592,N_7303,N_7231);
nand U7593 (N_7593,N_7181,N_7309);
and U7594 (N_7594,N_7367,N_7154);
or U7595 (N_7595,N_7337,N_7120);
nor U7596 (N_7596,N_7088,N_7471);
or U7597 (N_7597,N_7412,N_7116);
nor U7598 (N_7598,N_7012,N_7339);
nand U7599 (N_7599,N_7090,N_7380);
or U7600 (N_7600,N_7305,N_7102);
or U7601 (N_7601,N_7024,N_7108);
and U7602 (N_7602,N_7038,N_7433);
and U7603 (N_7603,N_7025,N_7478);
or U7604 (N_7604,N_7138,N_7023);
or U7605 (N_7605,N_7452,N_7067);
nor U7606 (N_7606,N_7394,N_7233);
nor U7607 (N_7607,N_7307,N_7018);
and U7608 (N_7608,N_7078,N_7467);
xnor U7609 (N_7609,N_7346,N_7273);
nor U7610 (N_7610,N_7427,N_7481);
and U7611 (N_7611,N_7491,N_7044);
nor U7612 (N_7612,N_7114,N_7146);
xnor U7613 (N_7613,N_7244,N_7214);
xor U7614 (N_7614,N_7395,N_7263);
and U7615 (N_7615,N_7075,N_7437);
or U7616 (N_7616,N_7243,N_7324);
xor U7617 (N_7617,N_7415,N_7374);
xor U7618 (N_7618,N_7366,N_7066);
xnor U7619 (N_7619,N_7310,N_7105);
nand U7620 (N_7620,N_7156,N_7418);
and U7621 (N_7621,N_7274,N_7247);
nor U7622 (N_7622,N_7122,N_7028);
nor U7623 (N_7623,N_7236,N_7070);
nor U7624 (N_7624,N_7135,N_7402);
nand U7625 (N_7625,N_7133,N_7112);
nand U7626 (N_7626,N_7095,N_7011);
or U7627 (N_7627,N_7333,N_7058);
nand U7628 (N_7628,N_7250,N_7323);
nor U7629 (N_7629,N_7390,N_7137);
nor U7630 (N_7630,N_7316,N_7084);
xnor U7631 (N_7631,N_7113,N_7125);
nor U7632 (N_7632,N_7197,N_7336);
or U7633 (N_7633,N_7453,N_7422);
and U7634 (N_7634,N_7056,N_7386);
nor U7635 (N_7635,N_7212,N_7119);
xor U7636 (N_7636,N_7005,N_7216);
nand U7637 (N_7637,N_7446,N_7057);
nor U7638 (N_7638,N_7097,N_7171);
nor U7639 (N_7639,N_7062,N_7355);
nor U7640 (N_7640,N_7104,N_7144);
nor U7641 (N_7641,N_7180,N_7287);
nand U7642 (N_7642,N_7123,N_7314);
nor U7643 (N_7643,N_7087,N_7016);
nand U7644 (N_7644,N_7080,N_7176);
xnor U7645 (N_7645,N_7030,N_7110);
nand U7646 (N_7646,N_7472,N_7445);
and U7647 (N_7647,N_7443,N_7098);
nand U7648 (N_7648,N_7493,N_7079);
nand U7649 (N_7649,N_7373,N_7271);
and U7650 (N_7650,N_7032,N_7254);
xnor U7651 (N_7651,N_7037,N_7159);
and U7652 (N_7652,N_7432,N_7195);
or U7653 (N_7653,N_7266,N_7343);
or U7654 (N_7654,N_7476,N_7464);
nor U7655 (N_7655,N_7042,N_7063);
xnor U7656 (N_7656,N_7103,N_7480);
and U7657 (N_7657,N_7198,N_7089);
and U7658 (N_7658,N_7404,N_7294);
and U7659 (N_7659,N_7242,N_7318);
nand U7660 (N_7660,N_7127,N_7139);
nor U7661 (N_7661,N_7234,N_7035);
nor U7662 (N_7662,N_7474,N_7151);
xnor U7663 (N_7663,N_7441,N_7313);
xnor U7664 (N_7664,N_7393,N_7049);
nand U7665 (N_7665,N_7315,N_7279);
xor U7666 (N_7666,N_7300,N_7183);
xor U7667 (N_7667,N_7426,N_7029);
nor U7668 (N_7668,N_7060,N_7099);
nand U7669 (N_7669,N_7260,N_7188);
nand U7670 (N_7670,N_7073,N_7043);
nand U7671 (N_7671,N_7059,N_7297);
nor U7672 (N_7672,N_7096,N_7400);
or U7673 (N_7673,N_7439,N_7296);
and U7674 (N_7674,N_7363,N_7447);
nand U7675 (N_7675,N_7359,N_7093);
nor U7676 (N_7676,N_7301,N_7289);
xor U7677 (N_7677,N_7264,N_7175);
and U7678 (N_7678,N_7036,N_7153);
xor U7679 (N_7679,N_7111,N_7055);
nand U7680 (N_7680,N_7191,N_7162);
xor U7681 (N_7681,N_7388,N_7454);
and U7682 (N_7682,N_7158,N_7221);
and U7683 (N_7683,N_7045,N_7496);
nand U7684 (N_7684,N_7076,N_7019);
and U7685 (N_7685,N_7085,N_7168);
or U7686 (N_7686,N_7143,N_7345);
nor U7687 (N_7687,N_7142,N_7262);
nand U7688 (N_7688,N_7200,N_7051);
and U7689 (N_7689,N_7407,N_7278);
nor U7690 (N_7690,N_7226,N_7434);
nand U7691 (N_7691,N_7132,N_7241);
and U7692 (N_7692,N_7131,N_7054);
nor U7693 (N_7693,N_7253,N_7040);
xnor U7694 (N_7694,N_7050,N_7475);
nand U7695 (N_7695,N_7259,N_7451);
nand U7696 (N_7696,N_7428,N_7438);
and U7697 (N_7697,N_7330,N_7326);
nand U7698 (N_7698,N_7106,N_7101);
xnor U7699 (N_7699,N_7389,N_7217);
xor U7700 (N_7700,N_7468,N_7499);
nor U7701 (N_7701,N_7331,N_7349);
xnor U7702 (N_7702,N_7230,N_7174);
or U7703 (N_7703,N_7003,N_7435);
xnor U7704 (N_7704,N_7046,N_7277);
nand U7705 (N_7705,N_7292,N_7213);
nor U7706 (N_7706,N_7155,N_7160);
nor U7707 (N_7707,N_7192,N_7117);
xnor U7708 (N_7708,N_7006,N_7440);
xor U7709 (N_7709,N_7382,N_7490);
and U7710 (N_7710,N_7202,N_7460);
xnor U7711 (N_7711,N_7473,N_7147);
xnor U7712 (N_7712,N_7420,N_7381);
nor U7713 (N_7713,N_7494,N_7170);
xnor U7714 (N_7714,N_7177,N_7017);
nand U7715 (N_7715,N_7456,N_7071);
or U7716 (N_7716,N_7321,N_7134);
nor U7717 (N_7717,N_7001,N_7219);
nand U7718 (N_7718,N_7356,N_7187);
nor U7719 (N_7719,N_7008,N_7368);
nand U7720 (N_7720,N_7322,N_7362);
nor U7721 (N_7721,N_7484,N_7448);
or U7722 (N_7722,N_7406,N_7369);
or U7723 (N_7723,N_7269,N_7357);
xor U7724 (N_7724,N_7211,N_7283);
xnor U7725 (N_7725,N_7015,N_7204);
xnor U7726 (N_7726,N_7286,N_7378);
xor U7727 (N_7727,N_7124,N_7235);
nor U7728 (N_7728,N_7411,N_7210);
nand U7729 (N_7729,N_7364,N_7069);
nand U7730 (N_7730,N_7398,N_7308);
xor U7731 (N_7731,N_7298,N_7249);
nor U7732 (N_7732,N_7039,N_7421);
nor U7733 (N_7733,N_7341,N_7257);
nor U7734 (N_7734,N_7182,N_7107);
nand U7735 (N_7735,N_7228,N_7344);
nor U7736 (N_7736,N_7163,N_7498);
nand U7737 (N_7737,N_7077,N_7121);
or U7738 (N_7738,N_7148,N_7026);
and U7739 (N_7739,N_7126,N_7186);
nand U7740 (N_7740,N_7455,N_7329);
or U7741 (N_7741,N_7173,N_7385);
nor U7742 (N_7742,N_7041,N_7285);
nor U7743 (N_7743,N_7350,N_7064);
or U7744 (N_7744,N_7423,N_7094);
xnor U7745 (N_7745,N_7081,N_7190);
xor U7746 (N_7746,N_7403,N_7083);
and U7747 (N_7747,N_7265,N_7166);
and U7748 (N_7748,N_7497,N_7410);
xor U7749 (N_7749,N_7425,N_7010);
and U7750 (N_7750,N_7285,N_7004);
nand U7751 (N_7751,N_7475,N_7160);
xnor U7752 (N_7752,N_7329,N_7418);
or U7753 (N_7753,N_7492,N_7093);
or U7754 (N_7754,N_7425,N_7100);
nor U7755 (N_7755,N_7387,N_7408);
and U7756 (N_7756,N_7278,N_7223);
and U7757 (N_7757,N_7173,N_7462);
nand U7758 (N_7758,N_7152,N_7195);
xor U7759 (N_7759,N_7297,N_7283);
and U7760 (N_7760,N_7323,N_7288);
xor U7761 (N_7761,N_7462,N_7165);
nor U7762 (N_7762,N_7206,N_7000);
and U7763 (N_7763,N_7248,N_7393);
or U7764 (N_7764,N_7325,N_7000);
xor U7765 (N_7765,N_7428,N_7343);
nand U7766 (N_7766,N_7429,N_7153);
nand U7767 (N_7767,N_7052,N_7089);
or U7768 (N_7768,N_7294,N_7008);
xnor U7769 (N_7769,N_7352,N_7062);
nor U7770 (N_7770,N_7413,N_7024);
or U7771 (N_7771,N_7356,N_7391);
xnor U7772 (N_7772,N_7221,N_7131);
or U7773 (N_7773,N_7456,N_7370);
xnor U7774 (N_7774,N_7220,N_7368);
or U7775 (N_7775,N_7187,N_7034);
xor U7776 (N_7776,N_7094,N_7350);
or U7777 (N_7777,N_7155,N_7285);
nand U7778 (N_7778,N_7470,N_7299);
or U7779 (N_7779,N_7123,N_7365);
or U7780 (N_7780,N_7228,N_7060);
nand U7781 (N_7781,N_7030,N_7166);
nor U7782 (N_7782,N_7405,N_7261);
or U7783 (N_7783,N_7355,N_7332);
or U7784 (N_7784,N_7320,N_7479);
and U7785 (N_7785,N_7085,N_7227);
or U7786 (N_7786,N_7398,N_7245);
xor U7787 (N_7787,N_7066,N_7154);
and U7788 (N_7788,N_7043,N_7141);
nand U7789 (N_7789,N_7390,N_7485);
nor U7790 (N_7790,N_7259,N_7458);
nor U7791 (N_7791,N_7105,N_7152);
and U7792 (N_7792,N_7058,N_7246);
nor U7793 (N_7793,N_7015,N_7016);
or U7794 (N_7794,N_7431,N_7301);
and U7795 (N_7795,N_7160,N_7252);
and U7796 (N_7796,N_7442,N_7423);
or U7797 (N_7797,N_7173,N_7426);
nand U7798 (N_7798,N_7001,N_7280);
nand U7799 (N_7799,N_7398,N_7481);
nand U7800 (N_7800,N_7395,N_7205);
or U7801 (N_7801,N_7081,N_7139);
nor U7802 (N_7802,N_7015,N_7238);
or U7803 (N_7803,N_7012,N_7179);
nor U7804 (N_7804,N_7278,N_7383);
nor U7805 (N_7805,N_7293,N_7290);
nor U7806 (N_7806,N_7366,N_7471);
and U7807 (N_7807,N_7340,N_7284);
or U7808 (N_7808,N_7106,N_7470);
xor U7809 (N_7809,N_7342,N_7469);
and U7810 (N_7810,N_7386,N_7026);
and U7811 (N_7811,N_7389,N_7231);
nand U7812 (N_7812,N_7145,N_7062);
nor U7813 (N_7813,N_7327,N_7336);
and U7814 (N_7814,N_7460,N_7074);
nor U7815 (N_7815,N_7082,N_7253);
and U7816 (N_7816,N_7284,N_7281);
xor U7817 (N_7817,N_7024,N_7406);
nor U7818 (N_7818,N_7047,N_7301);
xor U7819 (N_7819,N_7359,N_7237);
nor U7820 (N_7820,N_7285,N_7157);
nor U7821 (N_7821,N_7330,N_7230);
nor U7822 (N_7822,N_7317,N_7468);
and U7823 (N_7823,N_7455,N_7324);
or U7824 (N_7824,N_7021,N_7314);
xnor U7825 (N_7825,N_7436,N_7111);
xnor U7826 (N_7826,N_7204,N_7045);
nor U7827 (N_7827,N_7190,N_7386);
nand U7828 (N_7828,N_7222,N_7377);
nor U7829 (N_7829,N_7486,N_7309);
or U7830 (N_7830,N_7270,N_7469);
or U7831 (N_7831,N_7194,N_7049);
nor U7832 (N_7832,N_7008,N_7091);
nor U7833 (N_7833,N_7212,N_7470);
nor U7834 (N_7834,N_7418,N_7043);
xor U7835 (N_7835,N_7318,N_7255);
nand U7836 (N_7836,N_7492,N_7409);
and U7837 (N_7837,N_7424,N_7154);
and U7838 (N_7838,N_7071,N_7032);
and U7839 (N_7839,N_7334,N_7126);
nand U7840 (N_7840,N_7259,N_7408);
and U7841 (N_7841,N_7108,N_7151);
nor U7842 (N_7842,N_7331,N_7032);
and U7843 (N_7843,N_7401,N_7295);
and U7844 (N_7844,N_7281,N_7383);
or U7845 (N_7845,N_7441,N_7112);
nand U7846 (N_7846,N_7055,N_7091);
and U7847 (N_7847,N_7277,N_7488);
or U7848 (N_7848,N_7125,N_7242);
nor U7849 (N_7849,N_7229,N_7279);
xnor U7850 (N_7850,N_7343,N_7005);
and U7851 (N_7851,N_7022,N_7424);
or U7852 (N_7852,N_7140,N_7233);
or U7853 (N_7853,N_7149,N_7239);
nand U7854 (N_7854,N_7136,N_7205);
nand U7855 (N_7855,N_7129,N_7196);
nand U7856 (N_7856,N_7205,N_7469);
nor U7857 (N_7857,N_7309,N_7132);
or U7858 (N_7858,N_7320,N_7432);
nor U7859 (N_7859,N_7394,N_7443);
and U7860 (N_7860,N_7127,N_7243);
xnor U7861 (N_7861,N_7323,N_7442);
xor U7862 (N_7862,N_7087,N_7154);
or U7863 (N_7863,N_7181,N_7048);
and U7864 (N_7864,N_7247,N_7130);
nand U7865 (N_7865,N_7037,N_7076);
nor U7866 (N_7866,N_7121,N_7415);
or U7867 (N_7867,N_7007,N_7170);
xor U7868 (N_7868,N_7115,N_7272);
nand U7869 (N_7869,N_7238,N_7290);
or U7870 (N_7870,N_7238,N_7151);
nor U7871 (N_7871,N_7024,N_7411);
nand U7872 (N_7872,N_7140,N_7246);
nor U7873 (N_7873,N_7407,N_7057);
or U7874 (N_7874,N_7035,N_7268);
nor U7875 (N_7875,N_7375,N_7048);
nor U7876 (N_7876,N_7494,N_7254);
nand U7877 (N_7877,N_7384,N_7313);
xor U7878 (N_7878,N_7439,N_7092);
and U7879 (N_7879,N_7338,N_7034);
nor U7880 (N_7880,N_7309,N_7270);
and U7881 (N_7881,N_7416,N_7112);
xor U7882 (N_7882,N_7198,N_7497);
nor U7883 (N_7883,N_7306,N_7056);
or U7884 (N_7884,N_7223,N_7322);
and U7885 (N_7885,N_7422,N_7066);
and U7886 (N_7886,N_7270,N_7429);
or U7887 (N_7887,N_7150,N_7213);
xor U7888 (N_7888,N_7006,N_7127);
xor U7889 (N_7889,N_7195,N_7453);
xor U7890 (N_7890,N_7476,N_7451);
nand U7891 (N_7891,N_7482,N_7367);
nor U7892 (N_7892,N_7228,N_7048);
and U7893 (N_7893,N_7278,N_7476);
and U7894 (N_7894,N_7048,N_7235);
nand U7895 (N_7895,N_7096,N_7258);
nand U7896 (N_7896,N_7463,N_7431);
nand U7897 (N_7897,N_7029,N_7005);
xor U7898 (N_7898,N_7351,N_7099);
nor U7899 (N_7899,N_7361,N_7326);
or U7900 (N_7900,N_7161,N_7478);
nand U7901 (N_7901,N_7111,N_7282);
nand U7902 (N_7902,N_7139,N_7483);
or U7903 (N_7903,N_7042,N_7289);
or U7904 (N_7904,N_7406,N_7416);
nand U7905 (N_7905,N_7065,N_7132);
or U7906 (N_7906,N_7380,N_7282);
nor U7907 (N_7907,N_7070,N_7199);
and U7908 (N_7908,N_7391,N_7299);
and U7909 (N_7909,N_7132,N_7485);
nand U7910 (N_7910,N_7126,N_7318);
or U7911 (N_7911,N_7001,N_7399);
nor U7912 (N_7912,N_7014,N_7358);
or U7913 (N_7913,N_7175,N_7008);
nor U7914 (N_7914,N_7232,N_7298);
or U7915 (N_7915,N_7354,N_7498);
xnor U7916 (N_7916,N_7189,N_7389);
nand U7917 (N_7917,N_7410,N_7043);
nand U7918 (N_7918,N_7316,N_7044);
xor U7919 (N_7919,N_7065,N_7304);
nor U7920 (N_7920,N_7239,N_7371);
nor U7921 (N_7921,N_7046,N_7365);
xor U7922 (N_7922,N_7338,N_7156);
xor U7923 (N_7923,N_7295,N_7269);
or U7924 (N_7924,N_7397,N_7251);
or U7925 (N_7925,N_7356,N_7139);
and U7926 (N_7926,N_7057,N_7182);
nor U7927 (N_7927,N_7441,N_7065);
and U7928 (N_7928,N_7275,N_7056);
or U7929 (N_7929,N_7279,N_7211);
xor U7930 (N_7930,N_7459,N_7293);
xor U7931 (N_7931,N_7018,N_7036);
nor U7932 (N_7932,N_7335,N_7476);
nand U7933 (N_7933,N_7055,N_7325);
and U7934 (N_7934,N_7150,N_7358);
or U7935 (N_7935,N_7230,N_7352);
nor U7936 (N_7936,N_7231,N_7336);
xor U7937 (N_7937,N_7003,N_7223);
and U7938 (N_7938,N_7181,N_7191);
nor U7939 (N_7939,N_7173,N_7380);
nor U7940 (N_7940,N_7365,N_7341);
and U7941 (N_7941,N_7360,N_7419);
nand U7942 (N_7942,N_7105,N_7488);
xor U7943 (N_7943,N_7319,N_7351);
xnor U7944 (N_7944,N_7057,N_7017);
nand U7945 (N_7945,N_7325,N_7263);
and U7946 (N_7946,N_7300,N_7406);
and U7947 (N_7947,N_7400,N_7185);
or U7948 (N_7948,N_7486,N_7473);
nand U7949 (N_7949,N_7133,N_7093);
nor U7950 (N_7950,N_7408,N_7070);
or U7951 (N_7951,N_7085,N_7011);
or U7952 (N_7952,N_7366,N_7082);
xor U7953 (N_7953,N_7261,N_7094);
and U7954 (N_7954,N_7100,N_7043);
and U7955 (N_7955,N_7098,N_7408);
nand U7956 (N_7956,N_7267,N_7198);
nand U7957 (N_7957,N_7293,N_7174);
xor U7958 (N_7958,N_7201,N_7313);
and U7959 (N_7959,N_7352,N_7362);
and U7960 (N_7960,N_7070,N_7393);
nor U7961 (N_7961,N_7204,N_7489);
and U7962 (N_7962,N_7382,N_7055);
nand U7963 (N_7963,N_7450,N_7295);
xor U7964 (N_7964,N_7388,N_7018);
nand U7965 (N_7965,N_7414,N_7239);
and U7966 (N_7966,N_7481,N_7353);
or U7967 (N_7967,N_7486,N_7380);
xor U7968 (N_7968,N_7206,N_7150);
or U7969 (N_7969,N_7136,N_7347);
nor U7970 (N_7970,N_7423,N_7384);
and U7971 (N_7971,N_7216,N_7464);
nand U7972 (N_7972,N_7476,N_7229);
or U7973 (N_7973,N_7210,N_7233);
and U7974 (N_7974,N_7331,N_7362);
nor U7975 (N_7975,N_7213,N_7060);
xnor U7976 (N_7976,N_7084,N_7486);
nand U7977 (N_7977,N_7116,N_7211);
xnor U7978 (N_7978,N_7480,N_7157);
nand U7979 (N_7979,N_7174,N_7309);
xor U7980 (N_7980,N_7363,N_7116);
nand U7981 (N_7981,N_7326,N_7258);
xnor U7982 (N_7982,N_7183,N_7441);
and U7983 (N_7983,N_7087,N_7161);
nand U7984 (N_7984,N_7191,N_7143);
nor U7985 (N_7985,N_7101,N_7085);
xor U7986 (N_7986,N_7029,N_7054);
nor U7987 (N_7987,N_7246,N_7325);
nand U7988 (N_7988,N_7219,N_7269);
and U7989 (N_7989,N_7116,N_7436);
xnor U7990 (N_7990,N_7011,N_7301);
nand U7991 (N_7991,N_7003,N_7440);
or U7992 (N_7992,N_7308,N_7192);
and U7993 (N_7993,N_7405,N_7191);
nand U7994 (N_7994,N_7449,N_7325);
nand U7995 (N_7995,N_7133,N_7377);
xor U7996 (N_7996,N_7413,N_7089);
nand U7997 (N_7997,N_7060,N_7258);
or U7998 (N_7998,N_7365,N_7445);
nor U7999 (N_7999,N_7333,N_7422);
or U8000 (N_8000,N_7786,N_7572);
or U8001 (N_8001,N_7884,N_7540);
and U8002 (N_8002,N_7985,N_7817);
or U8003 (N_8003,N_7861,N_7908);
nand U8004 (N_8004,N_7671,N_7663);
or U8005 (N_8005,N_7839,N_7791);
or U8006 (N_8006,N_7926,N_7684);
xor U8007 (N_8007,N_7525,N_7758);
xor U8008 (N_8008,N_7611,N_7629);
xor U8009 (N_8009,N_7954,N_7746);
and U8010 (N_8010,N_7559,N_7959);
xnor U8011 (N_8011,N_7705,N_7974);
or U8012 (N_8012,N_7837,N_7711);
or U8013 (N_8013,N_7858,N_7813);
or U8014 (N_8014,N_7585,N_7823);
and U8015 (N_8015,N_7722,N_7683);
and U8016 (N_8016,N_7595,N_7770);
xnor U8017 (N_8017,N_7635,N_7565);
nor U8018 (N_8018,N_7987,N_7831);
and U8019 (N_8019,N_7665,N_7804);
nand U8020 (N_8020,N_7556,N_7912);
nand U8021 (N_8021,N_7668,N_7507);
and U8022 (N_8022,N_7606,N_7570);
xor U8023 (N_8023,N_7951,N_7883);
nand U8024 (N_8024,N_7851,N_7661);
nand U8025 (N_8025,N_7560,N_7502);
nand U8026 (N_8026,N_7516,N_7631);
nand U8027 (N_8027,N_7679,N_7744);
xor U8028 (N_8028,N_7872,N_7821);
and U8029 (N_8029,N_7520,N_7816);
nor U8030 (N_8030,N_7793,N_7524);
and U8031 (N_8031,N_7539,N_7917);
or U8032 (N_8032,N_7736,N_7913);
nor U8033 (N_8033,N_7914,N_7757);
nand U8034 (N_8034,N_7965,N_7939);
nor U8035 (N_8035,N_7810,N_7607);
nand U8036 (N_8036,N_7782,N_7933);
and U8037 (N_8037,N_7971,N_7656);
xor U8038 (N_8038,N_7522,N_7742);
and U8039 (N_8039,N_7827,N_7873);
xnor U8040 (N_8040,N_7836,N_7899);
or U8041 (N_8041,N_7709,N_7894);
xor U8042 (N_8042,N_7593,N_7584);
nor U8043 (N_8043,N_7530,N_7728);
xor U8044 (N_8044,N_7689,N_7515);
or U8045 (N_8045,N_7692,N_7698);
and U8046 (N_8046,N_7915,N_7561);
xor U8047 (N_8047,N_7680,N_7503);
and U8048 (N_8048,N_7976,N_7551);
or U8049 (N_8049,N_7845,N_7569);
nor U8050 (N_8050,N_7775,N_7592);
or U8051 (N_8051,N_7521,N_7970);
xor U8052 (N_8052,N_7903,N_7865);
xor U8053 (N_8053,N_7527,N_7989);
or U8054 (N_8054,N_7760,N_7616);
and U8055 (N_8055,N_7552,N_7844);
nor U8056 (N_8056,N_7734,N_7920);
nand U8057 (N_8057,N_7573,N_7938);
nor U8058 (N_8058,N_7774,N_7532);
and U8059 (N_8059,N_7519,N_7510);
xnor U8060 (N_8060,N_7598,N_7928);
nor U8061 (N_8061,N_7640,N_7935);
or U8062 (N_8062,N_7764,N_7518);
and U8063 (N_8063,N_7719,N_7644);
or U8064 (N_8064,N_7687,N_7988);
or U8065 (N_8065,N_7898,N_7832);
and U8066 (N_8066,N_7646,N_7927);
or U8067 (N_8067,N_7769,N_7923);
nor U8068 (N_8068,N_7922,N_7643);
and U8069 (N_8069,N_7534,N_7651);
and U8070 (N_8070,N_7547,N_7567);
xor U8071 (N_8071,N_7703,N_7797);
nor U8072 (N_8072,N_7800,N_7768);
and U8073 (N_8073,N_7608,N_7937);
nor U8074 (N_8074,N_7685,N_7716);
or U8075 (N_8075,N_7733,N_7767);
and U8076 (N_8076,N_7612,N_7802);
and U8077 (N_8077,N_7513,N_7747);
or U8078 (N_8078,N_7819,N_7980);
xnor U8079 (N_8079,N_7655,N_7968);
or U8080 (N_8080,N_7755,N_7712);
or U8081 (N_8081,N_7801,N_7619);
and U8082 (N_8082,N_7740,N_7849);
nand U8083 (N_8083,N_7864,N_7597);
or U8084 (N_8084,N_7627,N_7977);
xor U8085 (N_8085,N_7526,N_7895);
or U8086 (N_8086,N_7662,N_7785);
or U8087 (N_8087,N_7888,N_7523);
and U8088 (N_8088,N_7720,N_7967);
nor U8089 (N_8089,N_7596,N_7602);
or U8090 (N_8090,N_7856,N_7780);
and U8091 (N_8091,N_7590,N_7583);
xor U8092 (N_8092,N_7803,N_7549);
xor U8093 (N_8093,N_7706,N_7932);
and U8094 (N_8094,N_7792,N_7695);
nor U8095 (N_8095,N_7718,N_7529);
and U8096 (N_8096,N_7779,N_7838);
and U8097 (N_8097,N_7702,N_7991);
nor U8098 (N_8098,N_7541,N_7852);
xor U8099 (N_8099,N_7741,N_7835);
and U8100 (N_8100,N_7924,N_7633);
xnor U8101 (N_8101,N_7778,N_7958);
nand U8102 (N_8102,N_7807,N_7843);
and U8103 (N_8103,N_7670,N_7860);
xnor U8104 (N_8104,N_7833,N_7512);
nor U8105 (N_8105,N_7509,N_7617);
and U8106 (N_8106,N_7604,N_7754);
or U8107 (N_8107,N_7880,N_7535);
and U8108 (N_8108,N_7790,N_7881);
and U8109 (N_8109,N_7647,N_7870);
xnor U8110 (N_8110,N_7669,N_7739);
xor U8111 (N_8111,N_7961,N_7943);
and U8112 (N_8112,N_7936,N_7586);
and U8113 (N_8113,N_7842,N_7996);
nand U8114 (N_8114,N_7956,N_7505);
xnor U8115 (N_8115,N_7511,N_7855);
xor U8116 (N_8116,N_7528,N_7942);
and U8117 (N_8117,N_7994,N_7641);
xor U8118 (N_8118,N_7981,N_7879);
or U8119 (N_8119,N_7504,N_7745);
nand U8120 (N_8120,N_7723,N_7724);
nand U8121 (N_8121,N_7808,N_7568);
nor U8122 (N_8122,N_7892,N_7548);
nor U8123 (N_8123,N_7546,N_7834);
and U8124 (N_8124,N_7978,N_7626);
nor U8125 (N_8125,N_7624,N_7566);
nand U8126 (N_8126,N_7649,N_7576);
or U8127 (N_8127,N_7998,N_7866);
nor U8128 (N_8128,N_7918,N_7642);
and U8129 (N_8129,N_7882,N_7654);
xnor U8130 (N_8130,N_7621,N_7587);
xnor U8131 (N_8131,N_7652,N_7964);
and U8132 (N_8132,N_7953,N_7678);
xor U8133 (N_8133,N_7645,N_7979);
or U8134 (N_8134,N_7850,N_7876);
and U8135 (N_8135,N_7811,N_7916);
xor U8136 (N_8136,N_7787,N_7847);
xor U8137 (N_8137,N_7658,N_7925);
nand U8138 (N_8138,N_7634,N_7773);
or U8139 (N_8139,N_7885,N_7601);
and U8140 (N_8140,N_7829,N_7944);
and U8141 (N_8141,N_7828,N_7575);
xnor U8142 (N_8142,N_7948,N_7848);
and U8143 (N_8143,N_7579,N_7660);
or U8144 (N_8144,N_7657,N_7743);
xnor U8145 (N_8145,N_7675,N_7999);
nand U8146 (N_8146,N_7605,N_7506);
nor U8147 (N_8147,N_7867,N_7713);
xnor U8148 (N_8148,N_7542,N_7581);
or U8149 (N_8149,N_7940,N_7558);
and U8150 (N_8150,N_7783,N_7729);
or U8151 (N_8151,N_7906,N_7690);
and U8152 (N_8152,N_7955,N_7699);
nor U8153 (N_8153,N_7982,N_7929);
or U8154 (N_8154,N_7557,N_7615);
xor U8155 (N_8155,N_7667,N_7517);
or U8156 (N_8156,N_7550,N_7500);
xnor U8157 (N_8157,N_7806,N_7952);
nand U8158 (N_8158,N_7632,N_7708);
nor U8159 (N_8159,N_7578,N_7777);
nor U8160 (N_8160,N_7907,N_7763);
nand U8161 (N_8161,N_7911,N_7761);
or U8162 (N_8162,N_7600,N_7571);
nor U8163 (N_8163,N_7962,N_7853);
nand U8164 (N_8164,N_7580,N_7622);
and U8165 (N_8165,N_7805,N_7648);
nor U8166 (N_8166,N_7941,N_7676);
nor U8167 (N_8167,N_7891,N_7696);
or U8168 (N_8168,N_7704,N_7756);
nand U8169 (N_8169,N_7886,N_7666);
and U8170 (N_8170,N_7950,N_7609);
or U8171 (N_8171,N_7751,N_7825);
xnor U8172 (N_8172,N_7610,N_7591);
nand U8173 (N_8173,N_7904,N_7674);
xor U8174 (N_8174,N_7715,N_7931);
or U8175 (N_8175,N_7795,N_7840);
nand U8176 (N_8176,N_7772,N_7614);
nor U8177 (N_8177,N_7963,N_7983);
xor U8178 (N_8178,N_7677,N_7691);
and U8179 (N_8179,N_7620,N_7784);
nor U8180 (N_8180,N_7599,N_7721);
or U8181 (N_8181,N_7564,N_7887);
and U8182 (N_8182,N_7628,N_7582);
nand U8183 (N_8183,N_7700,N_7545);
nand U8184 (N_8184,N_7625,N_7863);
xor U8185 (N_8185,N_7543,N_7949);
and U8186 (N_8186,N_7533,N_7636);
xnor U8187 (N_8187,N_7794,N_7749);
nor U8188 (N_8188,N_7637,N_7613);
and U8189 (N_8189,N_7818,N_7969);
nand U8190 (N_8190,N_7889,N_7707);
xor U8191 (N_8191,N_7781,N_7947);
or U8192 (N_8192,N_7562,N_7650);
and U8193 (N_8193,N_7826,N_7897);
or U8194 (N_8194,N_7553,N_7623);
xnor U8195 (N_8195,N_7946,N_7859);
or U8196 (N_8196,N_7577,N_7701);
or U8197 (N_8197,N_7555,N_7789);
nor U8198 (N_8198,N_7750,N_7997);
and U8199 (N_8199,N_7846,N_7588);
and U8200 (N_8200,N_7673,N_7603);
xor U8201 (N_8201,N_7759,N_7735);
nand U8202 (N_8202,N_7544,N_7841);
nor U8203 (N_8203,N_7890,N_7896);
or U8204 (N_8204,N_7830,N_7815);
xor U8205 (N_8205,N_7871,N_7905);
nor U8206 (N_8206,N_7960,N_7752);
nand U8207 (N_8207,N_7869,N_7714);
and U8208 (N_8208,N_7984,N_7538);
xor U8209 (N_8209,N_7737,N_7659);
and U8210 (N_8210,N_7877,N_7738);
and U8211 (N_8211,N_7554,N_7874);
xnor U8212 (N_8212,N_7814,N_7725);
or U8213 (N_8213,N_7682,N_7717);
or U8214 (N_8214,N_7776,N_7796);
xor U8215 (N_8215,N_7730,N_7630);
or U8216 (N_8216,N_7653,N_7930);
or U8217 (N_8217,N_7875,N_7893);
or U8218 (N_8218,N_7710,N_7798);
or U8219 (N_8219,N_7788,N_7594);
nor U8220 (N_8220,N_7681,N_7639);
or U8221 (N_8221,N_7686,N_7694);
or U8222 (N_8222,N_7992,N_7731);
and U8223 (N_8223,N_7986,N_7868);
nand U8224 (N_8224,N_7766,N_7514);
nand U8225 (N_8225,N_7688,N_7857);
or U8226 (N_8226,N_7574,N_7824);
or U8227 (N_8227,N_7672,N_7799);
nor U8228 (N_8228,N_7854,N_7902);
nand U8229 (N_8229,N_7921,N_7771);
or U8230 (N_8230,N_7966,N_7753);
and U8231 (N_8231,N_7563,N_7638);
nand U8232 (N_8232,N_7910,N_7993);
nor U8233 (N_8233,N_7762,N_7972);
nand U8234 (N_8234,N_7531,N_7862);
nor U8235 (N_8235,N_7748,N_7901);
nor U8236 (N_8236,N_7693,N_7919);
nand U8237 (N_8237,N_7501,N_7934);
nor U8238 (N_8238,N_7726,N_7973);
and U8239 (N_8239,N_7975,N_7508);
and U8240 (N_8240,N_7909,N_7664);
nor U8241 (N_8241,N_7727,N_7812);
xor U8242 (N_8242,N_7900,N_7809);
xnor U8243 (N_8243,N_7822,N_7618);
and U8244 (N_8244,N_7537,N_7878);
and U8245 (N_8245,N_7945,N_7990);
xnor U8246 (N_8246,N_7536,N_7697);
nand U8247 (N_8247,N_7995,N_7732);
and U8248 (N_8248,N_7957,N_7589);
or U8249 (N_8249,N_7820,N_7765);
nand U8250 (N_8250,N_7773,N_7727);
or U8251 (N_8251,N_7943,N_7518);
xnor U8252 (N_8252,N_7783,N_7666);
and U8253 (N_8253,N_7738,N_7855);
and U8254 (N_8254,N_7637,N_7630);
and U8255 (N_8255,N_7799,N_7564);
xnor U8256 (N_8256,N_7772,N_7895);
nor U8257 (N_8257,N_7674,N_7777);
nand U8258 (N_8258,N_7631,N_7802);
xnor U8259 (N_8259,N_7954,N_7676);
xnor U8260 (N_8260,N_7962,N_7738);
nand U8261 (N_8261,N_7615,N_7703);
nand U8262 (N_8262,N_7723,N_7965);
or U8263 (N_8263,N_7869,N_7893);
nand U8264 (N_8264,N_7583,N_7753);
nor U8265 (N_8265,N_7738,N_7646);
xor U8266 (N_8266,N_7522,N_7787);
nand U8267 (N_8267,N_7526,N_7620);
or U8268 (N_8268,N_7728,N_7992);
and U8269 (N_8269,N_7862,N_7532);
nand U8270 (N_8270,N_7613,N_7720);
nor U8271 (N_8271,N_7864,N_7784);
or U8272 (N_8272,N_7549,N_7914);
nor U8273 (N_8273,N_7918,N_7872);
and U8274 (N_8274,N_7676,N_7584);
or U8275 (N_8275,N_7871,N_7765);
and U8276 (N_8276,N_7705,N_7956);
nand U8277 (N_8277,N_7656,N_7529);
or U8278 (N_8278,N_7633,N_7974);
nand U8279 (N_8279,N_7748,N_7977);
and U8280 (N_8280,N_7759,N_7700);
nand U8281 (N_8281,N_7683,N_7791);
or U8282 (N_8282,N_7929,N_7955);
nand U8283 (N_8283,N_7966,N_7731);
or U8284 (N_8284,N_7508,N_7911);
xnor U8285 (N_8285,N_7702,N_7577);
xnor U8286 (N_8286,N_7689,N_7953);
nor U8287 (N_8287,N_7847,N_7718);
or U8288 (N_8288,N_7822,N_7770);
xnor U8289 (N_8289,N_7840,N_7876);
and U8290 (N_8290,N_7994,N_7942);
and U8291 (N_8291,N_7979,N_7989);
xor U8292 (N_8292,N_7959,N_7968);
nor U8293 (N_8293,N_7878,N_7791);
xnor U8294 (N_8294,N_7778,N_7717);
or U8295 (N_8295,N_7987,N_7924);
or U8296 (N_8296,N_7717,N_7996);
nor U8297 (N_8297,N_7876,N_7685);
nor U8298 (N_8298,N_7899,N_7680);
xnor U8299 (N_8299,N_7881,N_7998);
xor U8300 (N_8300,N_7525,N_7713);
nand U8301 (N_8301,N_7866,N_7649);
xnor U8302 (N_8302,N_7750,N_7720);
or U8303 (N_8303,N_7586,N_7608);
and U8304 (N_8304,N_7781,N_7710);
and U8305 (N_8305,N_7847,N_7618);
xor U8306 (N_8306,N_7709,N_7531);
xnor U8307 (N_8307,N_7511,N_7929);
or U8308 (N_8308,N_7880,N_7707);
nand U8309 (N_8309,N_7551,N_7910);
xor U8310 (N_8310,N_7869,N_7544);
and U8311 (N_8311,N_7807,N_7932);
and U8312 (N_8312,N_7540,N_7969);
and U8313 (N_8313,N_7612,N_7559);
nor U8314 (N_8314,N_7832,N_7995);
nand U8315 (N_8315,N_7604,N_7636);
or U8316 (N_8316,N_7699,N_7570);
nand U8317 (N_8317,N_7915,N_7593);
and U8318 (N_8318,N_7714,N_7936);
nor U8319 (N_8319,N_7775,N_7937);
and U8320 (N_8320,N_7553,N_7693);
or U8321 (N_8321,N_7770,N_7549);
and U8322 (N_8322,N_7912,N_7536);
nor U8323 (N_8323,N_7539,N_7876);
nand U8324 (N_8324,N_7917,N_7838);
nor U8325 (N_8325,N_7706,N_7948);
xor U8326 (N_8326,N_7996,N_7570);
or U8327 (N_8327,N_7898,N_7839);
or U8328 (N_8328,N_7685,N_7833);
nand U8329 (N_8329,N_7624,N_7651);
or U8330 (N_8330,N_7960,N_7729);
nor U8331 (N_8331,N_7537,N_7656);
or U8332 (N_8332,N_7962,N_7610);
or U8333 (N_8333,N_7754,N_7536);
xor U8334 (N_8334,N_7697,N_7901);
or U8335 (N_8335,N_7668,N_7919);
nor U8336 (N_8336,N_7751,N_7938);
xnor U8337 (N_8337,N_7775,N_7890);
nand U8338 (N_8338,N_7904,N_7653);
nor U8339 (N_8339,N_7752,N_7817);
nor U8340 (N_8340,N_7897,N_7557);
xnor U8341 (N_8341,N_7938,N_7758);
nand U8342 (N_8342,N_7848,N_7554);
nor U8343 (N_8343,N_7511,N_7816);
nand U8344 (N_8344,N_7734,N_7963);
and U8345 (N_8345,N_7511,N_7641);
nor U8346 (N_8346,N_7737,N_7878);
or U8347 (N_8347,N_7608,N_7896);
xor U8348 (N_8348,N_7546,N_7758);
nand U8349 (N_8349,N_7787,N_7634);
nand U8350 (N_8350,N_7705,N_7606);
xor U8351 (N_8351,N_7941,N_7622);
and U8352 (N_8352,N_7727,N_7921);
nor U8353 (N_8353,N_7869,N_7958);
and U8354 (N_8354,N_7646,N_7907);
xor U8355 (N_8355,N_7839,N_7658);
nor U8356 (N_8356,N_7688,N_7579);
xor U8357 (N_8357,N_7732,N_7681);
nor U8358 (N_8358,N_7727,N_7591);
or U8359 (N_8359,N_7775,N_7851);
or U8360 (N_8360,N_7829,N_7638);
nand U8361 (N_8361,N_7700,N_7690);
nor U8362 (N_8362,N_7606,N_7557);
nand U8363 (N_8363,N_7973,N_7756);
xnor U8364 (N_8364,N_7756,N_7749);
xnor U8365 (N_8365,N_7966,N_7696);
nand U8366 (N_8366,N_7908,N_7511);
nand U8367 (N_8367,N_7780,N_7732);
or U8368 (N_8368,N_7812,N_7956);
and U8369 (N_8369,N_7646,N_7786);
nand U8370 (N_8370,N_7734,N_7961);
or U8371 (N_8371,N_7729,N_7962);
and U8372 (N_8372,N_7633,N_7854);
nand U8373 (N_8373,N_7936,N_7654);
or U8374 (N_8374,N_7751,N_7927);
or U8375 (N_8375,N_7876,N_7797);
or U8376 (N_8376,N_7743,N_7709);
nor U8377 (N_8377,N_7981,N_7656);
nor U8378 (N_8378,N_7816,N_7674);
and U8379 (N_8379,N_7574,N_7817);
or U8380 (N_8380,N_7827,N_7745);
nand U8381 (N_8381,N_7773,N_7980);
xor U8382 (N_8382,N_7768,N_7631);
and U8383 (N_8383,N_7666,N_7764);
and U8384 (N_8384,N_7630,N_7869);
and U8385 (N_8385,N_7675,N_7855);
and U8386 (N_8386,N_7825,N_7511);
nand U8387 (N_8387,N_7712,N_7620);
or U8388 (N_8388,N_7876,N_7503);
nand U8389 (N_8389,N_7774,N_7668);
nor U8390 (N_8390,N_7863,N_7563);
or U8391 (N_8391,N_7776,N_7722);
or U8392 (N_8392,N_7587,N_7669);
or U8393 (N_8393,N_7767,N_7709);
nand U8394 (N_8394,N_7565,N_7849);
and U8395 (N_8395,N_7765,N_7725);
and U8396 (N_8396,N_7988,N_7963);
or U8397 (N_8397,N_7527,N_7593);
nand U8398 (N_8398,N_7725,N_7975);
or U8399 (N_8399,N_7919,N_7524);
nor U8400 (N_8400,N_7846,N_7844);
and U8401 (N_8401,N_7927,N_7814);
and U8402 (N_8402,N_7991,N_7712);
and U8403 (N_8403,N_7728,N_7670);
nor U8404 (N_8404,N_7798,N_7728);
xnor U8405 (N_8405,N_7968,N_7517);
or U8406 (N_8406,N_7978,N_7803);
nand U8407 (N_8407,N_7795,N_7584);
and U8408 (N_8408,N_7870,N_7554);
and U8409 (N_8409,N_7933,N_7636);
nand U8410 (N_8410,N_7675,N_7548);
nor U8411 (N_8411,N_7753,N_7817);
xnor U8412 (N_8412,N_7961,N_7864);
or U8413 (N_8413,N_7936,N_7881);
xnor U8414 (N_8414,N_7633,N_7862);
nor U8415 (N_8415,N_7764,N_7865);
nor U8416 (N_8416,N_7977,N_7919);
nor U8417 (N_8417,N_7851,N_7681);
nand U8418 (N_8418,N_7885,N_7515);
or U8419 (N_8419,N_7824,N_7747);
xnor U8420 (N_8420,N_7601,N_7703);
nor U8421 (N_8421,N_7660,N_7628);
nor U8422 (N_8422,N_7987,N_7969);
xnor U8423 (N_8423,N_7880,N_7897);
or U8424 (N_8424,N_7874,N_7767);
or U8425 (N_8425,N_7530,N_7570);
and U8426 (N_8426,N_7683,N_7821);
xor U8427 (N_8427,N_7752,N_7593);
xor U8428 (N_8428,N_7833,N_7502);
nand U8429 (N_8429,N_7749,N_7732);
and U8430 (N_8430,N_7654,N_7713);
xor U8431 (N_8431,N_7552,N_7734);
nand U8432 (N_8432,N_7732,N_7736);
or U8433 (N_8433,N_7594,N_7509);
nand U8434 (N_8434,N_7691,N_7569);
nor U8435 (N_8435,N_7684,N_7894);
and U8436 (N_8436,N_7644,N_7706);
and U8437 (N_8437,N_7871,N_7554);
or U8438 (N_8438,N_7815,N_7604);
nand U8439 (N_8439,N_7753,N_7826);
or U8440 (N_8440,N_7659,N_7870);
nor U8441 (N_8441,N_7703,N_7552);
xor U8442 (N_8442,N_7706,N_7802);
and U8443 (N_8443,N_7557,N_7640);
or U8444 (N_8444,N_7753,N_7774);
and U8445 (N_8445,N_7898,N_7674);
xnor U8446 (N_8446,N_7803,N_7698);
or U8447 (N_8447,N_7830,N_7805);
xnor U8448 (N_8448,N_7886,N_7754);
or U8449 (N_8449,N_7879,N_7749);
xnor U8450 (N_8450,N_7798,N_7618);
or U8451 (N_8451,N_7838,N_7766);
and U8452 (N_8452,N_7564,N_7861);
and U8453 (N_8453,N_7506,N_7874);
nand U8454 (N_8454,N_7816,N_7647);
or U8455 (N_8455,N_7633,N_7629);
or U8456 (N_8456,N_7964,N_7537);
and U8457 (N_8457,N_7652,N_7949);
nor U8458 (N_8458,N_7819,N_7924);
or U8459 (N_8459,N_7833,N_7861);
nor U8460 (N_8460,N_7708,N_7860);
or U8461 (N_8461,N_7915,N_7966);
and U8462 (N_8462,N_7677,N_7823);
or U8463 (N_8463,N_7949,N_7691);
nor U8464 (N_8464,N_7750,N_7879);
and U8465 (N_8465,N_7721,N_7646);
nand U8466 (N_8466,N_7780,N_7887);
nor U8467 (N_8467,N_7508,N_7745);
nor U8468 (N_8468,N_7796,N_7984);
or U8469 (N_8469,N_7831,N_7751);
nand U8470 (N_8470,N_7935,N_7966);
nor U8471 (N_8471,N_7620,N_7951);
nand U8472 (N_8472,N_7846,N_7641);
nand U8473 (N_8473,N_7630,N_7559);
and U8474 (N_8474,N_7592,N_7983);
nor U8475 (N_8475,N_7788,N_7770);
nand U8476 (N_8476,N_7503,N_7746);
nor U8477 (N_8477,N_7971,N_7673);
or U8478 (N_8478,N_7796,N_7734);
xnor U8479 (N_8479,N_7955,N_7794);
or U8480 (N_8480,N_7591,N_7975);
or U8481 (N_8481,N_7623,N_7962);
xnor U8482 (N_8482,N_7717,N_7969);
or U8483 (N_8483,N_7770,N_7954);
xor U8484 (N_8484,N_7571,N_7722);
nor U8485 (N_8485,N_7920,N_7724);
and U8486 (N_8486,N_7759,N_7719);
nand U8487 (N_8487,N_7880,N_7753);
xnor U8488 (N_8488,N_7765,N_7707);
xor U8489 (N_8489,N_7622,N_7819);
and U8490 (N_8490,N_7822,N_7800);
xnor U8491 (N_8491,N_7744,N_7933);
nor U8492 (N_8492,N_7959,N_7847);
nand U8493 (N_8493,N_7604,N_7764);
and U8494 (N_8494,N_7943,N_7718);
and U8495 (N_8495,N_7905,N_7679);
xor U8496 (N_8496,N_7645,N_7997);
nand U8497 (N_8497,N_7561,N_7504);
and U8498 (N_8498,N_7855,N_7956);
or U8499 (N_8499,N_7820,N_7595);
or U8500 (N_8500,N_8237,N_8415);
and U8501 (N_8501,N_8168,N_8108);
or U8502 (N_8502,N_8428,N_8445);
or U8503 (N_8503,N_8223,N_8332);
nor U8504 (N_8504,N_8242,N_8377);
nand U8505 (N_8505,N_8158,N_8388);
nand U8506 (N_8506,N_8055,N_8310);
xor U8507 (N_8507,N_8100,N_8249);
nor U8508 (N_8508,N_8451,N_8162);
or U8509 (N_8509,N_8203,N_8058);
and U8510 (N_8510,N_8008,N_8328);
nand U8511 (N_8511,N_8190,N_8319);
nand U8512 (N_8512,N_8116,N_8066);
nand U8513 (N_8513,N_8414,N_8441);
or U8514 (N_8514,N_8124,N_8085);
or U8515 (N_8515,N_8060,N_8012);
nand U8516 (N_8516,N_8307,N_8404);
xor U8517 (N_8517,N_8245,N_8474);
or U8518 (N_8518,N_8061,N_8457);
or U8519 (N_8519,N_8102,N_8042);
nand U8520 (N_8520,N_8296,N_8326);
or U8521 (N_8521,N_8356,N_8001);
nand U8522 (N_8522,N_8215,N_8490);
and U8523 (N_8523,N_8460,N_8040);
or U8524 (N_8524,N_8391,N_8226);
nor U8525 (N_8525,N_8435,N_8436);
nand U8526 (N_8526,N_8094,N_8260);
nand U8527 (N_8527,N_8238,N_8021);
nor U8528 (N_8528,N_8165,N_8313);
nor U8529 (N_8529,N_8454,N_8253);
nor U8530 (N_8530,N_8230,N_8396);
or U8531 (N_8531,N_8473,N_8375);
or U8532 (N_8532,N_8355,N_8430);
nand U8533 (N_8533,N_8202,N_8269);
and U8534 (N_8534,N_8321,N_8188);
nor U8535 (N_8535,N_8185,N_8106);
nand U8536 (N_8536,N_8438,N_8411);
and U8537 (N_8537,N_8329,N_8099);
or U8538 (N_8538,N_8285,N_8265);
xor U8539 (N_8539,N_8292,N_8330);
nor U8540 (N_8540,N_8154,N_8323);
and U8541 (N_8541,N_8484,N_8127);
or U8542 (N_8542,N_8264,N_8191);
xnor U8543 (N_8543,N_8224,N_8125);
xnor U8544 (N_8544,N_8469,N_8337);
nor U8545 (N_8545,N_8029,N_8229);
nor U8546 (N_8546,N_8358,N_8405);
nand U8547 (N_8547,N_8302,N_8131);
and U8548 (N_8548,N_8416,N_8347);
and U8549 (N_8549,N_8344,N_8462);
nor U8550 (N_8550,N_8135,N_8240);
or U8551 (N_8551,N_8065,N_8104);
and U8552 (N_8552,N_8498,N_8286);
or U8553 (N_8553,N_8172,N_8367);
nand U8554 (N_8554,N_8376,N_8175);
or U8555 (N_8555,N_8161,N_8197);
or U8556 (N_8556,N_8251,N_8281);
and U8557 (N_8557,N_8045,N_8049);
or U8558 (N_8558,N_8083,N_8256);
or U8559 (N_8559,N_8290,N_8088);
xor U8560 (N_8560,N_8424,N_8426);
xnor U8561 (N_8561,N_8018,N_8220);
nor U8562 (N_8562,N_8013,N_8015);
xor U8563 (N_8563,N_8231,N_8455);
nand U8564 (N_8564,N_8280,N_8246);
nor U8565 (N_8565,N_8317,N_8263);
and U8566 (N_8566,N_8216,N_8222);
and U8567 (N_8567,N_8077,N_8174);
or U8568 (N_8568,N_8079,N_8316);
nand U8569 (N_8569,N_8402,N_8442);
or U8570 (N_8570,N_8343,N_8335);
nand U8571 (N_8571,N_8312,N_8348);
nor U8572 (N_8572,N_8373,N_8069);
and U8573 (N_8573,N_8132,N_8417);
nand U8574 (N_8574,N_8288,N_8480);
and U8575 (N_8575,N_8467,N_8090);
and U8576 (N_8576,N_8299,N_8204);
nor U8577 (N_8577,N_8005,N_8393);
or U8578 (N_8578,N_8047,N_8142);
and U8579 (N_8579,N_8051,N_8297);
xor U8580 (N_8580,N_8212,N_8091);
nand U8581 (N_8581,N_8019,N_8437);
xnor U8582 (N_8582,N_8499,N_8050);
and U8583 (N_8583,N_8118,N_8087);
or U8584 (N_8584,N_8293,N_8398);
or U8585 (N_8585,N_8192,N_8144);
nand U8586 (N_8586,N_8233,N_8456);
and U8587 (N_8587,N_8159,N_8370);
and U8588 (N_8588,N_8177,N_8225);
nand U8589 (N_8589,N_8123,N_8443);
xor U8590 (N_8590,N_8447,N_8383);
and U8591 (N_8591,N_8073,N_8007);
and U8592 (N_8592,N_8227,N_8180);
and U8593 (N_8593,N_8327,N_8493);
nor U8594 (N_8594,N_8481,N_8147);
xor U8595 (N_8595,N_8272,N_8163);
and U8596 (N_8596,N_8401,N_8022);
or U8597 (N_8597,N_8208,N_8394);
nor U8598 (N_8598,N_8410,N_8362);
nand U8599 (N_8599,N_8440,N_8365);
or U8600 (N_8600,N_8390,N_8363);
nor U8601 (N_8601,N_8076,N_8193);
xor U8602 (N_8602,N_8194,N_8145);
nor U8603 (N_8603,N_8221,N_8063);
xor U8604 (N_8604,N_8494,N_8214);
nand U8605 (N_8605,N_8030,N_8234);
xnor U8606 (N_8606,N_8271,N_8488);
nor U8607 (N_8607,N_8448,N_8181);
xnor U8608 (N_8608,N_8252,N_8418);
nand U8609 (N_8609,N_8122,N_8120);
and U8610 (N_8610,N_8157,N_8075);
and U8611 (N_8611,N_8399,N_8305);
xor U8612 (N_8612,N_8346,N_8107);
xnor U8613 (N_8613,N_8384,N_8115);
and U8614 (N_8614,N_8352,N_8217);
nor U8615 (N_8615,N_8336,N_8136);
xor U8616 (N_8616,N_8150,N_8366);
xnor U8617 (N_8617,N_8339,N_8156);
nand U8618 (N_8618,N_8259,N_8155);
nor U8619 (N_8619,N_8121,N_8138);
nand U8620 (N_8620,N_8206,N_8450);
and U8621 (N_8621,N_8446,N_8274);
or U8622 (N_8622,N_8479,N_8146);
and U8623 (N_8623,N_8432,N_8403);
nand U8624 (N_8624,N_8002,N_8137);
or U8625 (N_8625,N_8357,N_8017);
or U8626 (N_8626,N_8248,N_8482);
xnor U8627 (N_8627,N_8475,N_8064);
nand U8628 (N_8628,N_8109,N_8128);
and U8629 (N_8629,N_8184,N_8354);
nor U8630 (N_8630,N_8320,N_8491);
nor U8631 (N_8631,N_8232,N_8444);
and U8632 (N_8632,N_8054,N_8112);
or U8633 (N_8633,N_8291,N_8173);
xor U8634 (N_8634,N_8067,N_8186);
nand U8635 (N_8635,N_8408,N_8371);
and U8636 (N_8636,N_8287,N_8074);
or U8637 (N_8637,N_8089,N_8010);
nand U8638 (N_8638,N_8304,N_8166);
nor U8639 (N_8639,N_8470,N_8353);
and U8640 (N_8640,N_8477,N_8038);
xnor U8641 (N_8641,N_8036,N_8023);
or U8642 (N_8642,N_8277,N_8458);
and U8643 (N_8643,N_8325,N_8046);
nand U8644 (N_8644,N_8476,N_8345);
nor U8645 (N_8645,N_8306,N_8322);
xnor U8646 (N_8646,N_8176,N_8431);
or U8647 (N_8647,N_8011,N_8400);
nor U8648 (N_8648,N_8141,N_8392);
nor U8649 (N_8649,N_8301,N_8200);
nor U8650 (N_8650,N_8409,N_8461);
or U8651 (N_8651,N_8084,N_8338);
or U8652 (N_8652,N_8318,N_8062);
nand U8653 (N_8653,N_8465,N_8149);
nor U8654 (N_8654,N_8183,N_8093);
xor U8655 (N_8655,N_8459,N_8201);
nand U8656 (N_8656,N_8098,N_8374);
or U8657 (N_8657,N_8129,N_8284);
nor U8658 (N_8658,N_8210,N_8169);
nor U8659 (N_8659,N_8195,N_8235);
and U8660 (N_8660,N_8283,N_8315);
and U8661 (N_8661,N_8198,N_8261);
xnor U8662 (N_8662,N_8092,N_8031);
or U8663 (N_8663,N_8368,N_8387);
or U8664 (N_8664,N_8364,N_8407);
xor U8665 (N_8665,N_8349,N_8495);
nor U8666 (N_8666,N_8097,N_8333);
or U8667 (N_8667,N_8103,N_8453);
or U8668 (N_8668,N_8427,N_8369);
nand U8669 (N_8669,N_8267,N_8420);
xnor U8670 (N_8670,N_8026,N_8170);
nand U8671 (N_8671,N_8119,N_8489);
nor U8672 (N_8672,N_8207,N_8496);
nand U8673 (N_8673,N_8072,N_8360);
nand U8674 (N_8674,N_8134,N_8258);
nor U8675 (N_8675,N_8359,N_8492);
or U8676 (N_8676,N_8101,N_8449);
nor U8677 (N_8677,N_8487,N_8276);
nand U8678 (N_8678,N_8209,N_8110);
and U8679 (N_8679,N_8171,N_8334);
nor U8680 (N_8680,N_8041,N_8068);
and U8681 (N_8681,N_8389,N_8372);
xor U8682 (N_8682,N_8160,N_8429);
or U8683 (N_8683,N_8351,N_8000);
nor U8684 (N_8684,N_8035,N_8052);
and U8685 (N_8685,N_8303,N_8199);
nor U8686 (N_8686,N_8213,N_8324);
xnor U8687 (N_8687,N_8032,N_8178);
xor U8688 (N_8688,N_8406,N_8308);
nor U8689 (N_8689,N_8081,N_8148);
and U8690 (N_8690,N_8275,N_8314);
nand U8691 (N_8691,N_8250,N_8086);
xor U8692 (N_8692,N_8027,N_8028);
or U8693 (N_8693,N_8059,N_8434);
nand U8694 (N_8694,N_8361,N_8255);
nor U8695 (N_8695,N_8257,N_8298);
nor U8696 (N_8696,N_8382,N_8105);
nand U8697 (N_8697,N_8179,N_8006);
nand U8698 (N_8698,N_8020,N_8114);
xnor U8699 (N_8699,N_8289,N_8080);
nand U8700 (N_8700,N_8056,N_8472);
xor U8701 (N_8701,N_8048,N_8262);
and U8702 (N_8702,N_8196,N_8497);
xnor U8703 (N_8703,N_8009,N_8113);
nor U8704 (N_8704,N_8486,N_8471);
or U8705 (N_8705,N_8053,N_8243);
or U8706 (N_8706,N_8439,N_8140);
and U8707 (N_8707,N_8096,N_8167);
and U8708 (N_8708,N_8385,N_8311);
nand U8709 (N_8709,N_8139,N_8033);
nand U8710 (N_8710,N_8219,N_8413);
or U8711 (N_8711,N_8037,N_8247);
nand U8712 (N_8712,N_8025,N_8143);
xor U8713 (N_8713,N_8340,N_8386);
and U8714 (N_8714,N_8421,N_8350);
and U8715 (N_8715,N_8228,N_8419);
nor U8716 (N_8716,N_8133,N_8078);
nor U8717 (N_8717,N_8187,N_8433);
xor U8718 (N_8718,N_8082,N_8423);
nor U8719 (N_8719,N_8239,N_8266);
xor U8720 (N_8720,N_8483,N_8024);
nor U8721 (N_8721,N_8381,N_8071);
nor U8722 (N_8722,N_8095,N_8270);
or U8723 (N_8723,N_8044,N_8273);
nand U8724 (N_8724,N_8016,N_8463);
xnor U8725 (N_8725,N_8014,N_8282);
xor U8726 (N_8726,N_8378,N_8464);
nor U8727 (N_8727,N_8468,N_8452);
or U8728 (N_8728,N_8153,N_8254);
or U8729 (N_8729,N_8004,N_8039);
xnor U8730 (N_8730,N_8342,N_8279);
nand U8731 (N_8731,N_8003,N_8164);
and U8732 (N_8732,N_8211,N_8412);
nor U8733 (N_8733,N_8034,N_8111);
and U8734 (N_8734,N_8395,N_8236);
and U8735 (N_8735,N_8478,N_8152);
xor U8736 (N_8736,N_8397,N_8309);
nor U8737 (N_8737,N_8043,N_8205);
nor U8738 (N_8738,N_8241,N_8070);
and U8739 (N_8739,N_8331,N_8295);
nor U8740 (N_8740,N_8422,N_8057);
nand U8741 (N_8741,N_8341,N_8379);
and U8742 (N_8742,N_8485,N_8126);
or U8743 (N_8743,N_8151,N_8466);
nand U8744 (N_8744,N_8182,N_8130);
and U8745 (N_8745,N_8425,N_8117);
nor U8746 (N_8746,N_8244,N_8268);
and U8747 (N_8747,N_8189,N_8278);
and U8748 (N_8748,N_8380,N_8300);
or U8749 (N_8749,N_8294,N_8218);
and U8750 (N_8750,N_8269,N_8251);
nand U8751 (N_8751,N_8422,N_8356);
or U8752 (N_8752,N_8045,N_8318);
nor U8753 (N_8753,N_8357,N_8302);
or U8754 (N_8754,N_8187,N_8275);
xnor U8755 (N_8755,N_8231,N_8059);
xnor U8756 (N_8756,N_8179,N_8380);
xnor U8757 (N_8757,N_8322,N_8139);
xor U8758 (N_8758,N_8326,N_8245);
nand U8759 (N_8759,N_8116,N_8426);
or U8760 (N_8760,N_8418,N_8309);
and U8761 (N_8761,N_8424,N_8483);
xnor U8762 (N_8762,N_8454,N_8313);
xor U8763 (N_8763,N_8415,N_8333);
nor U8764 (N_8764,N_8479,N_8062);
nand U8765 (N_8765,N_8420,N_8184);
and U8766 (N_8766,N_8456,N_8081);
and U8767 (N_8767,N_8303,N_8305);
and U8768 (N_8768,N_8104,N_8010);
nand U8769 (N_8769,N_8469,N_8031);
or U8770 (N_8770,N_8261,N_8383);
or U8771 (N_8771,N_8281,N_8324);
or U8772 (N_8772,N_8120,N_8058);
xnor U8773 (N_8773,N_8259,N_8006);
nand U8774 (N_8774,N_8306,N_8115);
nand U8775 (N_8775,N_8276,N_8359);
nand U8776 (N_8776,N_8070,N_8395);
or U8777 (N_8777,N_8421,N_8218);
nor U8778 (N_8778,N_8402,N_8152);
nor U8779 (N_8779,N_8488,N_8254);
nor U8780 (N_8780,N_8328,N_8325);
nand U8781 (N_8781,N_8475,N_8072);
or U8782 (N_8782,N_8473,N_8340);
nand U8783 (N_8783,N_8376,N_8046);
or U8784 (N_8784,N_8236,N_8167);
xnor U8785 (N_8785,N_8373,N_8079);
nor U8786 (N_8786,N_8266,N_8111);
or U8787 (N_8787,N_8154,N_8490);
and U8788 (N_8788,N_8082,N_8402);
xor U8789 (N_8789,N_8246,N_8413);
and U8790 (N_8790,N_8209,N_8178);
or U8791 (N_8791,N_8099,N_8245);
and U8792 (N_8792,N_8131,N_8079);
nor U8793 (N_8793,N_8424,N_8175);
and U8794 (N_8794,N_8137,N_8070);
and U8795 (N_8795,N_8012,N_8319);
xor U8796 (N_8796,N_8001,N_8430);
and U8797 (N_8797,N_8168,N_8369);
nor U8798 (N_8798,N_8325,N_8279);
nand U8799 (N_8799,N_8034,N_8333);
or U8800 (N_8800,N_8361,N_8222);
xor U8801 (N_8801,N_8246,N_8448);
and U8802 (N_8802,N_8238,N_8257);
or U8803 (N_8803,N_8086,N_8062);
or U8804 (N_8804,N_8258,N_8137);
and U8805 (N_8805,N_8210,N_8306);
nor U8806 (N_8806,N_8289,N_8439);
and U8807 (N_8807,N_8379,N_8055);
and U8808 (N_8808,N_8182,N_8453);
nor U8809 (N_8809,N_8017,N_8362);
nor U8810 (N_8810,N_8064,N_8044);
and U8811 (N_8811,N_8119,N_8067);
nand U8812 (N_8812,N_8131,N_8452);
xnor U8813 (N_8813,N_8248,N_8461);
xor U8814 (N_8814,N_8429,N_8401);
nor U8815 (N_8815,N_8227,N_8184);
and U8816 (N_8816,N_8347,N_8056);
and U8817 (N_8817,N_8119,N_8463);
nand U8818 (N_8818,N_8008,N_8308);
nor U8819 (N_8819,N_8364,N_8325);
or U8820 (N_8820,N_8070,N_8200);
nand U8821 (N_8821,N_8146,N_8281);
or U8822 (N_8822,N_8051,N_8056);
or U8823 (N_8823,N_8028,N_8279);
nor U8824 (N_8824,N_8411,N_8217);
nand U8825 (N_8825,N_8085,N_8305);
and U8826 (N_8826,N_8128,N_8234);
and U8827 (N_8827,N_8214,N_8022);
nor U8828 (N_8828,N_8498,N_8224);
nand U8829 (N_8829,N_8143,N_8197);
or U8830 (N_8830,N_8370,N_8222);
and U8831 (N_8831,N_8167,N_8117);
nor U8832 (N_8832,N_8437,N_8057);
nor U8833 (N_8833,N_8032,N_8177);
or U8834 (N_8834,N_8499,N_8232);
xnor U8835 (N_8835,N_8089,N_8301);
and U8836 (N_8836,N_8275,N_8492);
nor U8837 (N_8837,N_8385,N_8161);
and U8838 (N_8838,N_8428,N_8194);
nand U8839 (N_8839,N_8051,N_8423);
and U8840 (N_8840,N_8033,N_8467);
and U8841 (N_8841,N_8096,N_8175);
nand U8842 (N_8842,N_8282,N_8126);
xor U8843 (N_8843,N_8334,N_8446);
or U8844 (N_8844,N_8319,N_8296);
nor U8845 (N_8845,N_8275,N_8306);
nand U8846 (N_8846,N_8126,N_8433);
nand U8847 (N_8847,N_8388,N_8363);
or U8848 (N_8848,N_8307,N_8224);
nand U8849 (N_8849,N_8397,N_8225);
xnor U8850 (N_8850,N_8034,N_8072);
nor U8851 (N_8851,N_8413,N_8442);
xor U8852 (N_8852,N_8296,N_8293);
or U8853 (N_8853,N_8204,N_8138);
nand U8854 (N_8854,N_8112,N_8456);
xnor U8855 (N_8855,N_8151,N_8337);
nor U8856 (N_8856,N_8204,N_8234);
nor U8857 (N_8857,N_8390,N_8236);
xor U8858 (N_8858,N_8040,N_8061);
and U8859 (N_8859,N_8474,N_8099);
nand U8860 (N_8860,N_8251,N_8274);
and U8861 (N_8861,N_8208,N_8036);
or U8862 (N_8862,N_8162,N_8035);
and U8863 (N_8863,N_8187,N_8212);
or U8864 (N_8864,N_8320,N_8180);
or U8865 (N_8865,N_8462,N_8076);
and U8866 (N_8866,N_8042,N_8489);
nand U8867 (N_8867,N_8218,N_8390);
xnor U8868 (N_8868,N_8264,N_8355);
and U8869 (N_8869,N_8211,N_8039);
and U8870 (N_8870,N_8102,N_8277);
or U8871 (N_8871,N_8276,N_8178);
or U8872 (N_8872,N_8356,N_8474);
or U8873 (N_8873,N_8458,N_8227);
or U8874 (N_8874,N_8034,N_8247);
nand U8875 (N_8875,N_8396,N_8062);
nor U8876 (N_8876,N_8347,N_8476);
nand U8877 (N_8877,N_8381,N_8124);
nand U8878 (N_8878,N_8498,N_8075);
and U8879 (N_8879,N_8401,N_8076);
nand U8880 (N_8880,N_8009,N_8489);
or U8881 (N_8881,N_8045,N_8355);
and U8882 (N_8882,N_8342,N_8375);
nand U8883 (N_8883,N_8069,N_8021);
nand U8884 (N_8884,N_8366,N_8011);
and U8885 (N_8885,N_8211,N_8329);
nand U8886 (N_8886,N_8489,N_8071);
nor U8887 (N_8887,N_8471,N_8265);
xnor U8888 (N_8888,N_8392,N_8109);
nor U8889 (N_8889,N_8162,N_8308);
nand U8890 (N_8890,N_8373,N_8432);
nand U8891 (N_8891,N_8388,N_8258);
nand U8892 (N_8892,N_8160,N_8047);
or U8893 (N_8893,N_8103,N_8387);
and U8894 (N_8894,N_8186,N_8057);
nor U8895 (N_8895,N_8394,N_8335);
nand U8896 (N_8896,N_8440,N_8279);
nor U8897 (N_8897,N_8026,N_8131);
and U8898 (N_8898,N_8496,N_8166);
or U8899 (N_8899,N_8085,N_8120);
or U8900 (N_8900,N_8049,N_8295);
xnor U8901 (N_8901,N_8349,N_8337);
and U8902 (N_8902,N_8113,N_8233);
or U8903 (N_8903,N_8393,N_8434);
or U8904 (N_8904,N_8162,N_8345);
and U8905 (N_8905,N_8275,N_8323);
nor U8906 (N_8906,N_8408,N_8281);
nand U8907 (N_8907,N_8036,N_8152);
xor U8908 (N_8908,N_8004,N_8403);
nand U8909 (N_8909,N_8409,N_8171);
or U8910 (N_8910,N_8228,N_8283);
xnor U8911 (N_8911,N_8371,N_8347);
nor U8912 (N_8912,N_8226,N_8249);
xor U8913 (N_8913,N_8307,N_8021);
nor U8914 (N_8914,N_8131,N_8195);
xnor U8915 (N_8915,N_8366,N_8179);
xor U8916 (N_8916,N_8380,N_8216);
or U8917 (N_8917,N_8481,N_8290);
nand U8918 (N_8918,N_8334,N_8161);
nor U8919 (N_8919,N_8167,N_8422);
nor U8920 (N_8920,N_8260,N_8076);
or U8921 (N_8921,N_8044,N_8087);
and U8922 (N_8922,N_8489,N_8257);
or U8923 (N_8923,N_8388,N_8425);
nand U8924 (N_8924,N_8056,N_8329);
xor U8925 (N_8925,N_8225,N_8398);
xnor U8926 (N_8926,N_8136,N_8252);
nor U8927 (N_8927,N_8239,N_8310);
nor U8928 (N_8928,N_8364,N_8028);
nand U8929 (N_8929,N_8024,N_8049);
or U8930 (N_8930,N_8390,N_8240);
xor U8931 (N_8931,N_8043,N_8388);
and U8932 (N_8932,N_8253,N_8408);
and U8933 (N_8933,N_8149,N_8474);
xor U8934 (N_8934,N_8222,N_8138);
nor U8935 (N_8935,N_8429,N_8289);
xnor U8936 (N_8936,N_8408,N_8470);
xor U8937 (N_8937,N_8048,N_8016);
or U8938 (N_8938,N_8453,N_8279);
nand U8939 (N_8939,N_8144,N_8357);
nand U8940 (N_8940,N_8458,N_8091);
nor U8941 (N_8941,N_8146,N_8191);
or U8942 (N_8942,N_8342,N_8237);
or U8943 (N_8943,N_8141,N_8145);
and U8944 (N_8944,N_8035,N_8346);
or U8945 (N_8945,N_8155,N_8230);
xnor U8946 (N_8946,N_8443,N_8228);
xnor U8947 (N_8947,N_8284,N_8454);
or U8948 (N_8948,N_8297,N_8017);
or U8949 (N_8949,N_8406,N_8141);
nand U8950 (N_8950,N_8119,N_8370);
xor U8951 (N_8951,N_8358,N_8167);
or U8952 (N_8952,N_8000,N_8029);
nor U8953 (N_8953,N_8488,N_8265);
or U8954 (N_8954,N_8032,N_8357);
xor U8955 (N_8955,N_8144,N_8222);
nor U8956 (N_8956,N_8340,N_8141);
nand U8957 (N_8957,N_8368,N_8291);
or U8958 (N_8958,N_8268,N_8119);
and U8959 (N_8959,N_8411,N_8289);
or U8960 (N_8960,N_8404,N_8113);
and U8961 (N_8961,N_8325,N_8403);
nand U8962 (N_8962,N_8130,N_8454);
nand U8963 (N_8963,N_8378,N_8208);
xor U8964 (N_8964,N_8012,N_8267);
nor U8965 (N_8965,N_8004,N_8485);
or U8966 (N_8966,N_8079,N_8223);
xor U8967 (N_8967,N_8412,N_8037);
nand U8968 (N_8968,N_8428,N_8330);
nor U8969 (N_8969,N_8469,N_8116);
or U8970 (N_8970,N_8035,N_8307);
xnor U8971 (N_8971,N_8435,N_8401);
and U8972 (N_8972,N_8485,N_8254);
nor U8973 (N_8973,N_8163,N_8085);
or U8974 (N_8974,N_8207,N_8053);
and U8975 (N_8975,N_8008,N_8379);
or U8976 (N_8976,N_8361,N_8358);
or U8977 (N_8977,N_8061,N_8316);
nand U8978 (N_8978,N_8425,N_8021);
and U8979 (N_8979,N_8373,N_8225);
or U8980 (N_8980,N_8309,N_8381);
nand U8981 (N_8981,N_8435,N_8039);
nand U8982 (N_8982,N_8007,N_8132);
nor U8983 (N_8983,N_8440,N_8367);
nor U8984 (N_8984,N_8033,N_8205);
xnor U8985 (N_8985,N_8297,N_8391);
and U8986 (N_8986,N_8446,N_8460);
nor U8987 (N_8987,N_8146,N_8062);
nor U8988 (N_8988,N_8296,N_8226);
or U8989 (N_8989,N_8041,N_8128);
nor U8990 (N_8990,N_8122,N_8481);
xnor U8991 (N_8991,N_8232,N_8106);
nor U8992 (N_8992,N_8003,N_8422);
nor U8993 (N_8993,N_8209,N_8106);
xor U8994 (N_8994,N_8462,N_8082);
and U8995 (N_8995,N_8022,N_8305);
xnor U8996 (N_8996,N_8109,N_8001);
and U8997 (N_8997,N_8104,N_8387);
xnor U8998 (N_8998,N_8376,N_8087);
or U8999 (N_8999,N_8027,N_8295);
and U9000 (N_9000,N_8882,N_8838);
and U9001 (N_9001,N_8949,N_8896);
nor U9002 (N_9002,N_8737,N_8871);
xor U9003 (N_9003,N_8521,N_8576);
and U9004 (N_9004,N_8705,N_8651);
or U9005 (N_9005,N_8557,N_8850);
nand U9006 (N_9006,N_8534,N_8506);
and U9007 (N_9007,N_8726,N_8797);
nor U9008 (N_9008,N_8591,N_8806);
xnor U9009 (N_9009,N_8599,N_8607);
and U9010 (N_9010,N_8768,N_8745);
or U9011 (N_9011,N_8809,N_8958);
xnor U9012 (N_9012,N_8878,N_8728);
nor U9013 (N_9013,N_8953,N_8652);
or U9014 (N_9014,N_8743,N_8614);
nor U9015 (N_9015,N_8761,N_8841);
and U9016 (N_9016,N_8788,N_8787);
and U9017 (N_9017,N_8957,N_8682);
or U9018 (N_9018,N_8702,N_8596);
xnor U9019 (N_9019,N_8538,N_8644);
and U9020 (N_9020,N_8764,N_8843);
nand U9021 (N_9021,N_8823,N_8588);
nor U9022 (N_9022,N_8869,N_8713);
xnor U9023 (N_9023,N_8872,N_8844);
xnor U9024 (N_9024,N_8803,N_8573);
or U9025 (N_9025,N_8912,N_8877);
or U9026 (N_9026,N_8560,N_8537);
nand U9027 (N_9027,N_8839,N_8733);
xor U9028 (N_9028,N_8974,N_8720);
nor U9029 (N_9029,N_8827,N_8902);
or U9030 (N_9030,N_8561,N_8815);
nand U9031 (N_9031,N_8566,N_8837);
xor U9032 (N_9032,N_8884,N_8829);
and U9033 (N_9033,N_8893,N_8834);
and U9034 (N_9034,N_8621,N_8615);
nand U9035 (N_9035,N_8629,N_8890);
and U9036 (N_9036,N_8666,N_8980);
and U9037 (N_9037,N_8865,N_8796);
or U9038 (N_9038,N_8710,N_8555);
or U9039 (N_9039,N_8821,N_8805);
or U9040 (N_9040,N_8680,N_8904);
or U9041 (N_9041,N_8687,N_8747);
nand U9042 (N_9042,N_8985,N_8715);
xnor U9043 (N_9043,N_8751,N_8598);
and U9044 (N_9044,N_8739,N_8723);
and U9045 (N_9045,N_8766,N_8583);
xor U9046 (N_9046,N_8888,N_8785);
nand U9047 (N_9047,N_8669,N_8595);
or U9048 (N_9048,N_8870,N_8661);
and U9049 (N_9049,N_8756,N_8918);
nand U9050 (N_9050,N_8721,N_8714);
or U9051 (N_9051,N_8757,N_8531);
xnor U9052 (N_9052,N_8848,N_8759);
nand U9053 (N_9053,N_8584,N_8618);
nor U9054 (N_9054,N_8678,N_8916);
or U9055 (N_9055,N_8986,N_8933);
and U9056 (N_9056,N_8536,N_8836);
nand U9057 (N_9057,N_8518,N_8697);
nor U9058 (N_9058,N_8601,N_8558);
xnor U9059 (N_9059,N_8993,N_8820);
or U9060 (N_9060,N_8660,N_8541);
nor U9061 (N_9061,N_8992,N_8662);
xnor U9062 (N_9062,N_8817,N_8683);
and U9063 (N_9063,N_8990,N_8559);
and U9064 (N_9064,N_8753,N_8690);
and U9065 (N_9065,N_8971,N_8794);
or U9066 (N_9066,N_8771,N_8590);
or U9067 (N_9067,N_8845,N_8866);
xnor U9068 (N_9068,N_8623,N_8847);
or U9069 (N_9069,N_8988,N_8909);
nand U9070 (N_9070,N_8706,N_8592);
xnor U9071 (N_9071,N_8998,N_8552);
nand U9072 (N_9072,N_8926,N_8956);
and U9073 (N_9073,N_8649,N_8906);
xnor U9074 (N_9074,N_8528,N_8892);
or U9075 (N_9075,N_8711,N_8999);
xnor U9076 (N_9076,N_8655,N_8594);
and U9077 (N_9077,N_8658,N_8966);
and U9078 (N_9078,N_8790,N_8860);
nand U9079 (N_9079,N_8968,N_8638);
xnor U9080 (N_9080,N_8522,N_8754);
and U9081 (N_9081,N_8931,N_8670);
and U9082 (N_9082,N_8626,N_8873);
or U9083 (N_9083,N_8502,N_8619);
nand U9084 (N_9084,N_8948,N_8840);
nand U9085 (N_9085,N_8556,N_8671);
or U9086 (N_9086,N_8608,N_8944);
and U9087 (N_9087,N_8709,N_8819);
nand U9088 (N_9088,N_8852,N_8548);
nor U9089 (N_9089,N_8940,N_8786);
and U9090 (N_9090,N_8507,N_8693);
xor U9091 (N_9091,N_8574,N_8734);
and U9092 (N_9092,N_8738,N_8854);
or U9093 (N_9093,N_8910,N_8879);
and U9094 (N_9094,N_8579,N_8960);
xor U9095 (N_9095,N_8544,N_8587);
and U9096 (N_9096,N_8859,N_8874);
xnor U9097 (N_9097,N_8970,N_8719);
xor U9098 (N_9098,N_8630,N_8965);
nand U9099 (N_9099,N_8939,N_8774);
xor U9100 (N_9100,N_8832,N_8791);
xnor U9101 (N_9101,N_8984,N_8928);
and U9102 (N_9102,N_8616,N_8523);
or U9103 (N_9103,N_8744,N_8602);
nor U9104 (N_9104,N_8569,N_8604);
and U9105 (N_9105,N_8934,N_8914);
xnor U9106 (N_9106,N_8593,N_8898);
xor U9107 (N_9107,N_8762,N_8831);
xnor U9108 (N_9108,N_8810,N_8643);
nor U9109 (N_9109,N_8826,N_8677);
nand U9110 (N_9110,N_8636,N_8514);
xnor U9111 (N_9111,N_8818,N_8936);
nor U9112 (N_9112,N_8853,N_8704);
xnor U9113 (N_9113,N_8802,N_8695);
or U9114 (N_9114,N_8937,N_8770);
nor U9115 (N_9115,N_8779,N_8943);
xnor U9116 (N_9116,N_8858,N_8568);
xnor U9117 (N_9117,N_8967,N_8765);
nor U9118 (N_9118,N_8927,N_8606);
or U9119 (N_9119,N_8816,N_8505);
or U9120 (N_9120,N_8625,N_8775);
xor U9121 (N_9121,N_8907,N_8567);
and U9122 (N_9122,N_8730,N_8500);
nand U9123 (N_9123,N_8688,N_8897);
nand U9124 (N_9124,N_8922,N_8947);
and U9125 (N_9125,N_8707,N_8863);
xnor U9126 (N_9126,N_8696,N_8613);
nor U9127 (N_9127,N_8763,N_8700);
xnor U9128 (N_9128,N_8830,N_8855);
and U9129 (N_9129,N_8641,N_8981);
nor U9130 (N_9130,N_8777,N_8868);
or U9131 (N_9131,N_8609,N_8814);
nand U9132 (N_9132,N_8575,N_8982);
or U9133 (N_9133,N_8973,N_8637);
nand U9134 (N_9134,N_8674,N_8824);
nand U9135 (N_9135,N_8708,N_8659);
xnor U9136 (N_9136,N_8955,N_8813);
nand U9137 (N_9137,N_8656,N_8749);
or U9138 (N_9138,N_8856,N_8640);
nor U9139 (N_9139,N_8952,N_8520);
nor U9140 (N_9140,N_8510,N_8935);
and U9141 (N_9141,N_8822,N_8772);
and U9142 (N_9142,N_8800,N_8736);
xor U9143 (N_9143,N_8976,N_8735);
or U9144 (N_9144,N_8894,N_8972);
nor U9145 (N_9145,N_8833,N_8954);
xor U9146 (N_9146,N_8672,N_8673);
xnor U9147 (N_9147,N_8792,N_8938);
and U9148 (N_9148,N_8929,N_8741);
or U9149 (N_9149,N_8582,N_8610);
or U9150 (N_9150,N_8701,N_8513);
or U9151 (N_9151,N_8950,N_8646);
xor U9152 (N_9152,N_8798,N_8703);
nand U9153 (N_9153,N_8554,N_8901);
or U9154 (N_9154,N_8501,N_8789);
xor U9155 (N_9155,N_8645,N_8729);
or U9156 (N_9156,N_8540,N_8812);
nor U9157 (N_9157,N_8851,N_8577);
nor U9158 (N_9158,N_8570,N_8908);
xor U9159 (N_9159,N_8517,N_8628);
or U9160 (N_9160,N_8564,N_8899);
or U9161 (N_9161,N_8755,N_8919);
xor U9162 (N_9162,N_8781,N_8750);
xnor U9163 (N_9163,N_8597,N_8905);
or U9164 (N_9164,N_8565,N_8808);
nor U9165 (N_9165,N_8586,N_8539);
nand U9166 (N_9166,N_8684,N_8795);
nand U9167 (N_9167,N_8699,N_8722);
xor U9168 (N_9168,N_8642,N_8535);
nor U9169 (N_9169,N_8600,N_8553);
nor U9170 (N_9170,N_8532,N_8545);
nand U9171 (N_9171,N_8605,N_8758);
nand U9172 (N_9172,N_8867,N_8585);
xnor U9173 (N_9173,N_8941,N_8718);
or U9174 (N_9174,N_8634,N_8917);
nand U9175 (N_9175,N_8508,N_8793);
xor U9176 (N_9176,N_8691,N_8686);
nand U9177 (N_9177,N_8681,N_8978);
and U9178 (N_9178,N_8524,N_8846);
nor U9179 (N_9179,N_8503,N_8530);
nand U9180 (N_9180,N_8664,N_8886);
or U9181 (N_9181,N_8861,N_8546);
or U9182 (N_9182,N_8946,N_8782);
xnor U9183 (N_9183,N_8675,N_8977);
or U9184 (N_9184,N_8667,N_8983);
xnor U9185 (N_9185,N_8987,N_8945);
nand U9186 (N_9186,N_8525,N_8516);
xnor U9187 (N_9187,N_8911,N_8969);
or U9188 (N_9188,N_8889,N_8549);
xnor U9189 (N_9189,N_8580,N_8875);
and U9190 (N_9190,N_8835,N_8880);
or U9191 (N_9191,N_8589,N_8891);
and U9192 (N_9192,N_8930,N_8663);
xor U9193 (N_9193,N_8581,N_8519);
nand U9194 (N_9194,N_8620,N_8769);
and U9195 (N_9195,N_8746,N_8921);
or U9196 (N_9196,N_8533,N_8685);
nor U9197 (N_9197,N_8679,N_8612);
and U9198 (N_9198,N_8784,N_8924);
or U9199 (N_9199,N_8676,N_8961);
and U9200 (N_9200,N_8920,N_8780);
or U9201 (N_9201,N_8694,N_8962);
or U9202 (N_9202,N_8883,N_8627);
and U9203 (N_9203,N_8740,N_8509);
or U9204 (N_9204,N_8542,N_8975);
xor U9205 (N_9205,N_8724,N_8932);
nor U9206 (N_9206,N_8716,N_8842);
nor U9207 (N_9207,N_8731,N_8783);
or U9208 (N_9208,N_8571,N_8997);
nor U9209 (N_9209,N_8773,N_8903);
and U9210 (N_9210,N_8752,N_8633);
nand U9211 (N_9211,N_8923,N_8825);
nor U9212 (N_9212,N_8611,N_8578);
xnor U9213 (N_9213,N_8653,N_8547);
xor U9214 (N_9214,N_8742,N_8900);
nor U9215 (N_9215,N_8635,N_8563);
or U9216 (N_9216,N_8632,N_8959);
nor U9217 (N_9217,N_8515,N_8915);
xor U9218 (N_9218,N_8748,N_8648);
or U9219 (N_9219,N_8727,N_8807);
and U9220 (N_9220,N_8964,N_8698);
and U9221 (N_9221,N_8725,N_8994);
nand U9222 (N_9222,N_8996,N_8864);
xnor U9223 (N_9223,N_8951,N_8654);
and U9224 (N_9224,N_8527,N_8828);
xor U9225 (N_9225,N_8562,N_8804);
and U9226 (N_9226,N_8551,N_8778);
nor U9227 (N_9227,N_8767,N_8991);
nor U9228 (N_9228,N_8512,N_8572);
nand U9229 (N_9229,N_8760,N_8995);
or U9230 (N_9230,N_8862,N_8963);
or U9231 (N_9231,N_8799,N_8887);
nor U9232 (N_9232,N_8529,N_8624);
nand U9233 (N_9233,N_8603,N_8504);
and U9234 (N_9234,N_8732,N_8543);
and U9235 (N_9235,N_8650,N_8617);
and U9236 (N_9236,N_8913,N_8692);
or U9237 (N_9237,N_8876,N_8885);
nand U9238 (N_9238,N_8622,N_8857);
nor U9239 (N_9239,N_8647,N_8639);
nor U9240 (N_9240,N_8665,N_8550);
nor U9241 (N_9241,N_8895,N_8511);
or U9242 (N_9242,N_8689,N_8631);
and U9243 (N_9243,N_8989,N_8979);
nand U9244 (N_9244,N_8668,N_8776);
nor U9245 (N_9245,N_8811,N_8801);
and U9246 (N_9246,N_8717,N_8925);
or U9247 (N_9247,N_8657,N_8526);
nor U9248 (N_9248,N_8712,N_8881);
and U9249 (N_9249,N_8942,N_8849);
nor U9250 (N_9250,N_8997,N_8998);
nand U9251 (N_9251,N_8919,N_8931);
nand U9252 (N_9252,N_8604,N_8808);
and U9253 (N_9253,N_8573,N_8969);
nor U9254 (N_9254,N_8570,N_8910);
nand U9255 (N_9255,N_8690,N_8682);
xnor U9256 (N_9256,N_8531,N_8994);
nand U9257 (N_9257,N_8875,N_8802);
and U9258 (N_9258,N_8595,N_8770);
nand U9259 (N_9259,N_8698,N_8903);
nand U9260 (N_9260,N_8897,N_8800);
and U9261 (N_9261,N_8830,N_8803);
or U9262 (N_9262,N_8715,N_8638);
nand U9263 (N_9263,N_8679,N_8658);
and U9264 (N_9264,N_8882,N_8844);
and U9265 (N_9265,N_8688,N_8964);
nor U9266 (N_9266,N_8905,N_8935);
xor U9267 (N_9267,N_8723,N_8531);
nand U9268 (N_9268,N_8570,N_8895);
or U9269 (N_9269,N_8538,N_8638);
xor U9270 (N_9270,N_8969,N_8619);
nand U9271 (N_9271,N_8978,N_8713);
nand U9272 (N_9272,N_8630,N_8738);
nor U9273 (N_9273,N_8866,N_8970);
xnor U9274 (N_9274,N_8822,N_8880);
or U9275 (N_9275,N_8713,N_8706);
nor U9276 (N_9276,N_8980,N_8582);
nand U9277 (N_9277,N_8611,N_8530);
nor U9278 (N_9278,N_8892,N_8793);
nand U9279 (N_9279,N_8527,N_8552);
nor U9280 (N_9280,N_8660,N_8641);
or U9281 (N_9281,N_8563,N_8933);
or U9282 (N_9282,N_8579,N_8953);
xor U9283 (N_9283,N_8880,N_8827);
xor U9284 (N_9284,N_8930,N_8864);
nor U9285 (N_9285,N_8877,N_8575);
xor U9286 (N_9286,N_8519,N_8640);
and U9287 (N_9287,N_8841,N_8771);
nor U9288 (N_9288,N_8570,N_8905);
nand U9289 (N_9289,N_8710,N_8790);
and U9290 (N_9290,N_8971,N_8846);
nor U9291 (N_9291,N_8781,N_8985);
and U9292 (N_9292,N_8683,N_8580);
xor U9293 (N_9293,N_8636,N_8836);
nor U9294 (N_9294,N_8628,N_8851);
nand U9295 (N_9295,N_8721,N_8650);
xor U9296 (N_9296,N_8516,N_8669);
and U9297 (N_9297,N_8854,N_8507);
or U9298 (N_9298,N_8627,N_8523);
and U9299 (N_9299,N_8838,N_8815);
or U9300 (N_9300,N_8913,N_8897);
nand U9301 (N_9301,N_8882,N_8754);
nor U9302 (N_9302,N_8555,N_8759);
or U9303 (N_9303,N_8956,N_8775);
nor U9304 (N_9304,N_8988,N_8822);
nand U9305 (N_9305,N_8654,N_8784);
or U9306 (N_9306,N_8986,N_8851);
nand U9307 (N_9307,N_8673,N_8995);
nor U9308 (N_9308,N_8817,N_8754);
xor U9309 (N_9309,N_8553,N_8709);
and U9310 (N_9310,N_8664,N_8514);
nor U9311 (N_9311,N_8517,N_8721);
and U9312 (N_9312,N_8924,N_8596);
and U9313 (N_9313,N_8961,N_8716);
nand U9314 (N_9314,N_8712,N_8709);
and U9315 (N_9315,N_8931,N_8912);
nor U9316 (N_9316,N_8936,N_8945);
xnor U9317 (N_9317,N_8816,N_8536);
nand U9318 (N_9318,N_8523,N_8858);
nor U9319 (N_9319,N_8511,N_8942);
xnor U9320 (N_9320,N_8956,N_8852);
xor U9321 (N_9321,N_8599,N_8680);
nand U9322 (N_9322,N_8724,N_8756);
nand U9323 (N_9323,N_8509,N_8575);
nor U9324 (N_9324,N_8570,N_8806);
nor U9325 (N_9325,N_8805,N_8642);
and U9326 (N_9326,N_8534,N_8784);
or U9327 (N_9327,N_8512,N_8755);
nor U9328 (N_9328,N_8909,N_8507);
nor U9329 (N_9329,N_8838,N_8813);
or U9330 (N_9330,N_8684,N_8660);
and U9331 (N_9331,N_8844,N_8757);
and U9332 (N_9332,N_8956,N_8999);
and U9333 (N_9333,N_8918,N_8729);
nand U9334 (N_9334,N_8968,N_8659);
nor U9335 (N_9335,N_8947,N_8928);
nor U9336 (N_9336,N_8925,N_8978);
and U9337 (N_9337,N_8968,N_8953);
or U9338 (N_9338,N_8884,N_8873);
or U9339 (N_9339,N_8604,N_8595);
and U9340 (N_9340,N_8638,N_8919);
nand U9341 (N_9341,N_8989,N_8866);
xor U9342 (N_9342,N_8627,N_8997);
nand U9343 (N_9343,N_8980,N_8694);
nand U9344 (N_9344,N_8515,N_8599);
xnor U9345 (N_9345,N_8705,N_8810);
or U9346 (N_9346,N_8809,N_8530);
and U9347 (N_9347,N_8855,N_8588);
xor U9348 (N_9348,N_8884,N_8624);
nand U9349 (N_9349,N_8855,N_8825);
and U9350 (N_9350,N_8753,N_8956);
xor U9351 (N_9351,N_8838,N_8730);
xnor U9352 (N_9352,N_8633,N_8786);
xor U9353 (N_9353,N_8521,N_8946);
nor U9354 (N_9354,N_8634,N_8691);
nor U9355 (N_9355,N_8837,N_8985);
nand U9356 (N_9356,N_8909,N_8745);
xnor U9357 (N_9357,N_8699,N_8587);
and U9358 (N_9358,N_8740,N_8545);
nand U9359 (N_9359,N_8524,N_8695);
or U9360 (N_9360,N_8653,N_8790);
xnor U9361 (N_9361,N_8782,N_8896);
nand U9362 (N_9362,N_8599,N_8954);
or U9363 (N_9363,N_8511,N_8906);
or U9364 (N_9364,N_8695,N_8717);
nand U9365 (N_9365,N_8539,N_8971);
or U9366 (N_9366,N_8511,N_8717);
and U9367 (N_9367,N_8593,N_8990);
xnor U9368 (N_9368,N_8695,N_8729);
xor U9369 (N_9369,N_8936,N_8686);
nand U9370 (N_9370,N_8775,N_8535);
nor U9371 (N_9371,N_8550,N_8718);
or U9372 (N_9372,N_8789,N_8850);
nor U9373 (N_9373,N_8995,N_8581);
and U9374 (N_9374,N_8513,N_8883);
nor U9375 (N_9375,N_8786,N_8971);
or U9376 (N_9376,N_8634,N_8794);
nand U9377 (N_9377,N_8637,N_8988);
or U9378 (N_9378,N_8977,N_8841);
nor U9379 (N_9379,N_8667,N_8656);
nand U9380 (N_9380,N_8945,N_8720);
and U9381 (N_9381,N_8922,N_8711);
xnor U9382 (N_9382,N_8591,N_8644);
and U9383 (N_9383,N_8788,N_8705);
or U9384 (N_9384,N_8573,N_8527);
xnor U9385 (N_9385,N_8503,N_8934);
nor U9386 (N_9386,N_8552,N_8578);
xor U9387 (N_9387,N_8626,N_8652);
xor U9388 (N_9388,N_8691,N_8900);
and U9389 (N_9389,N_8806,N_8600);
xor U9390 (N_9390,N_8545,N_8554);
nand U9391 (N_9391,N_8980,N_8885);
nand U9392 (N_9392,N_8695,N_8881);
and U9393 (N_9393,N_8834,N_8517);
xor U9394 (N_9394,N_8596,N_8532);
xor U9395 (N_9395,N_8698,N_8921);
and U9396 (N_9396,N_8931,N_8589);
xnor U9397 (N_9397,N_8699,N_8819);
nand U9398 (N_9398,N_8983,N_8505);
or U9399 (N_9399,N_8736,N_8529);
nor U9400 (N_9400,N_8946,N_8952);
xnor U9401 (N_9401,N_8711,N_8956);
and U9402 (N_9402,N_8668,N_8563);
or U9403 (N_9403,N_8793,N_8585);
nor U9404 (N_9404,N_8613,N_8824);
and U9405 (N_9405,N_8556,N_8854);
nand U9406 (N_9406,N_8820,N_8774);
nor U9407 (N_9407,N_8816,N_8838);
xnor U9408 (N_9408,N_8575,N_8562);
nor U9409 (N_9409,N_8626,N_8784);
nor U9410 (N_9410,N_8772,N_8926);
or U9411 (N_9411,N_8882,N_8898);
and U9412 (N_9412,N_8578,N_8998);
nand U9413 (N_9413,N_8931,N_8539);
and U9414 (N_9414,N_8874,N_8688);
or U9415 (N_9415,N_8889,N_8537);
or U9416 (N_9416,N_8612,N_8834);
nand U9417 (N_9417,N_8937,N_8515);
nand U9418 (N_9418,N_8657,N_8867);
nor U9419 (N_9419,N_8716,N_8715);
or U9420 (N_9420,N_8758,N_8850);
xor U9421 (N_9421,N_8665,N_8613);
or U9422 (N_9422,N_8911,N_8663);
nand U9423 (N_9423,N_8572,N_8601);
nor U9424 (N_9424,N_8915,N_8774);
or U9425 (N_9425,N_8587,N_8516);
nand U9426 (N_9426,N_8664,N_8605);
or U9427 (N_9427,N_8953,N_8689);
nand U9428 (N_9428,N_8699,N_8744);
nor U9429 (N_9429,N_8974,N_8906);
or U9430 (N_9430,N_8730,N_8717);
and U9431 (N_9431,N_8562,N_8604);
nor U9432 (N_9432,N_8816,N_8902);
and U9433 (N_9433,N_8838,N_8581);
nand U9434 (N_9434,N_8612,N_8688);
or U9435 (N_9435,N_8966,N_8544);
nand U9436 (N_9436,N_8949,N_8655);
and U9437 (N_9437,N_8792,N_8543);
and U9438 (N_9438,N_8753,N_8712);
nand U9439 (N_9439,N_8928,N_8638);
nor U9440 (N_9440,N_8604,N_8516);
or U9441 (N_9441,N_8694,N_8898);
nor U9442 (N_9442,N_8878,N_8779);
nand U9443 (N_9443,N_8895,N_8539);
and U9444 (N_9444,N_8878,N_8783);
or U9445 (N_9445,N_8606,N_8997);
nand U9446 (N_9446,N_8770,N_8846);
nand U9447 (N_9447,N_8864,N_8721);
xnor U9448 (N_9448,N_8970,N_8924);
nand U9449 (N_9449,N_8605,N_8678);
nor U9450 (N_9450,N_8754,N_8607);
nand U9451 (N_9451,N_8574,N_8746);
nor U9452 (N_9452,N_8558,N_8664);
nor U9453 (N_9453,N_8708,N_8517);
nor U9454 (N_9454,N_8848,N_8597);
nand U9455 (N_9455,N_8771,N_8744);
and U9456 (N_9456,N_8892,N_8702);
nor U9457 (N_9457,N_8527,N_8629);
and U9458 (N_9458,N_8936,N_8735);
or U9459 (N_9459,N_8672,N_8733);
and U9460 (N_9460,N_8847,N_8975);
and U9461 (N_9461,N_8760,N_8780);
or U9462 (N_9462,N_8745,N_8625);
nand U9463 (N_9463,N_8674,N_8929);
or U9464 (N_9464,N_8673,N_8539);
or U9465 (N_9465,N_8586,N_8732);
nand U9466 (N_9466,N_8919,N_8640);
nor U9467 (N_9467,N_8814,N_8522);
nand U9468 (N_9468,N_8757,N_8625);
xor U9469 (N_9469,N_8581,N_8969);
xnor U9470 (N_9470,N_8744,N_8925);
nor U9471 (N_9471,N_8622,N_8763);
nor U9472 (N_9472,N_8783,N_8838);
nand U9473 (N_9473,N_8673,N_8892);
nor U9474 (N_9474,N_8742,N_8684);
xor U9475 (N_9475,N_8565,N_8693);
nor U9476 (N_9476,N_8801,N_8814);
xnor U9477 (N_9477,N_8978,N_8795);
nor U9478 (N_9478,N_8703,N_8637);
nor U9479 (N_9479,N_8736,N_8717);
or U9480 (N_9480,N_8717,N_8817);
nand U9481 (N_9481,N_8640,N_8888);
nand U9482 (N_9482,N_8979,N_8777);
nor U9483 (N_9483,N_8948,N_8535);
and U9484 (N_9484,N_8757,N_8832);
or U9485 (N_9485,N_8836,N_8720);
nor U9486 (N_9486,N_8567,N_8911);
nand U9487 (N_9487,N_8988,N_8504);
xor U9488 (N_9488,N_8793,N_8648);
nand U9489 (N_9489,N_8581,N_8545);
nor U9490 (N_9490,N_8753,N_8656);
and U9491 (N_9491,N_8717,N_8845);
nand U9492 (N_9492,N_8846,N_8783);
nand U9493 (N_9493,N_8699,N_8663);
and U9494 (N_9494,N_8620,N_8913);
and U9495 (N_9495,N_8669,N_8580);
nand U9496 (N_9496,N_8748,N_8900);
nor U9497 (N_9497,N_8987,N_8767);
and U9498 (N_9498,N_8726,N_8507);
nor U9499 (N_9499,N_8862,N_8907);
nor U9500 (N_9500,N_9328,N_9336);
nand U9501 (N_9501,N_9280,N_9379);
and U9502 (N_9502,N_9143,N_9162);
nand U9503 (N_9503,N_9092,N_9137);
xnor U9504 (N_9504,N_9145,N_9176);
nand U9505 (N_9505,N_9397,N_9108);
nand U9506 (N_9506,N_9148,N_9307);
nand U9507 (N_9507,N_9495,N_9332);
and U9508 (N_9508,N_9300,N_9412);
or U9509 (N_9509,N_9022,N_9353);
xor U9510 (N_9510,N_9260,N_9270);
xnor U9511 (N_9511,N_9301,N_9457);
and U9512 (N_9512,N_9334,N_9481);
and U9513 (N_9513,N_9019,N_9103);
or U9514 (N_9514,N_9093,N_9211);
xor U9515 (N_9515,N_9393,N_9361);
xor U9516 (N_9516,N_9290,N_9335);
nor U9517 (N_9517,N_9321,N_9253);
xor U9518 (N_9518,N_9070,N_9207);
or U9519 (N_9519,N_9248,N_9487);
and U9520 (N_9520,N_9465,N_9198);
or U9521 (N_9521,N_9292,N_9446);
nand U9522 (N_9522,N_9122,N_9175);
or U9523 (N_9523,N_9043,N_9042);
nor U9524 (N_9524,N_9343,N_9217);
xnor U9525 (N_9525,N_9499,N_9383);
xor U9526 (N_9526,N_9144,N_9247);
or U9527 (N_9527,N_9045,N_9249);
nor U9528 (N_9528,N_9064,N_9405);
nor U9529 (N_9529,N_9391,N_9479);
nand U9530 (N_9530,N_9406,N_9413);
nor U9531 (N_9531,N_9432,N_9411);
or U9532 (N_9532,N_9297,N_9053);
and U9533 (N_9533,N_9483,N_9130);
or U9534 (N_9534,N_9165,N_9371);
and U9535 (N_9535,N_9470,N_9235);
and U9536 (N_9536,N_9017,N_9200);
or U9537 (N_9537,N_9267,N_9416);
and U9538 (N_9538,N_9478,N_9206);
and U9539 (N_9539,N_9132,N_9273);
or U9540 (N_9540,N_9239,N_9427);
nand U9541 (N_9541,N_9255,N_9288);
nor U9542 (N_9542,N_9490,N_9046);
and U9543 (N_9543,N_9475,N_9011);
nand U9544 (N_9544,N_9072,N_9403);
nand U9545 (N_9545,N_9073,N_9319);
xnor U9546 (N_9546,N_9453,N_9456);
nor U9547 (N_9547,N_9348,N_9068);
nor U9548 (N_9548,N_9090,N_9396);
nor U9549 (N_9549,N_9149,N_9473);
or U9550 (N_9550,N_9182,N_9197);
nor U9551 (N_9551,N_9357,N_9250);
xnor U9552 (N_9552,N_9298,N_9408);
nand U9553 (N_9553,N_9430,N_9060);
nand U9554 (N_9554,N_9223,N_9291);
or U9555 (N_9555,N_9238,N_9049);
nand U9556 (N_9556,N_9443,N_9189);
or U9557 (N_9557,N_9299,N_9016);
and U9558 (N_9558,N_9415,N_9477);
or U9559 (N_9559,N_9180,N_9256);
nor U9560 (N_9560,N_9054,N_9215);
nand U9561 (N_9561,N_9059,N_9057);
nand U9562 (N_9562,N_9114,N_9433);
xor U9563 (N_9563,N_9376,N_9174);
and U9564 (N_9564,N_9034,N_9095);
nand U9565 (N_9565,N_9214,N_9099);
xnor U9566 (N_9566,N_9218,N_9106);
nor U9567 (N_9567,N_9467,N_9442);
or U9568 (N_9568,N_9313,N_9401);
and U9569 (N_9569,N_9326,N_9121);
nand U9570 (N_9570,N_9362,N_9126);
and U9571 (N_9571,N_9240,N_9025);
or U9572 (N_9572,N_9212,N_9370);
nor U9573 (N_9573,N_9316,N_9233);
xnor U9574 (N_9574,N_9493,N_9167);
and U9575 (N_9575,N_9242,N_9344);
or U9576 (N_9576,N_9436,N_9489);
nor U9577 (N_9577,N_9262,N_9040);
nand U9578 (N_9578,N_9410,N_9252);
nand U9579 (N_9579,N_9423,N_9384);
or U9580 (N_9580,N_9354,N_9352);
nand U9581 (N_9581,N_9277,N_9205);
nand U9582 (N_9582,N_9373,N_9210);
nand U9583 (N_9583,N_9086,N_9098);
and U9584 (N_9584,N_9220,N_9044);
and U9585 (N_9585,N_9461,N_9380);
nand U9586 (N_9586,N_9107,N_9105);
xnor U9587 (N_9587,N_9278,N_9439);
and U9588 (N_9588,N_9026,N_9183);
or U9589 (N_9589,N_9450,N_9331);
or U9590 (N_9590,N_9261,N_9437);
and U9591 (N_9591,N_9279,N_9209);
nor U9592 (N_9592,N_9010,N_9399);
or U9593 (N_9593,N_9431,N_9056);
nor U9594 (N_9594,N_9081,N_9458);
nor U9595 (N_9595,N_9468,N_9360);
or U9596 (N_9596,N_9318,N_9116);
and U9597 (N_9597,N_9322,N_9346);
or U9598 (N_9598,N_9077,N_9033);
nand U9599 (N_9599,N_9089,N_9041);
xor U9600 (N_9600,N_9364,N_9094);
xnor U9601 (N_9601,N_9150,N_9381);
nor U9602 (N_9602,N_9039,N_9320);
xor U9603 (N_9603,N_9296,N_9258);
and U9604 (N_9604,N_9002,N_9448);
and U9605 (N_9605,N_9003,N_9190);
nand U9606 (N_9606,N_9271,N_9225);
nor U9607 (N_9607,N_9498,N_9356);
or U9608 (N_9608,N_9492,N_9272);
nor U9609 (N_9609,N_9484,N_9440);
nand U9610 (N_9610,N_9324,N_9111);
or U9611 (N_9611,N_9164,N_9204);
xor U9612 (N_9612,N_9485,N_9452);
nand U9613 (N_9613,N_9222,N_9259);
and U9614 (N_9614,N_9203,N_9055);
or U9615 (N_9615,N_9141,N_9323);
or U9616 (N_9616,N_9173,N_9066);
nor U9617 (N_9617,N_9177,N_9192);
or U9618 (N_9618,N_9385,N_9382);
nor U9619 (N_9619,N_9251,N_9163);
nand U9620 (N_9620,N_9065,N_9418);
nand U9621 (N_9621,N_9110,N_9422);
or U9622 (N_9622,N_9109,N_9372);
and U9623 (N_9623,N_9306,N_9063);
xor U9624 (N_9624,N_9369,N_9265);
or U9625 (N_9625,N_9359,N_9085);
nor U9626 (N_9626,N_9023,N_9184);
and U9627 (N_9627,N_9230,N_9229);
or U9628 (N_9628,N_9488,N_9133);
or U9629 (N_9629,N_9069,N_9181);
and U9630 (N_9630,N_9154,N_9394);
nand U9631 (N_9631,N_9274,N_9425);
and U9632 (N_9632,N_9367,N_9084);
xnor U9633 (N_9633,N_9135,N_9191);
xnor U9634 (N_9634,N_9139,N_9464);
xor U9635 (N_9635,N_9158,N_9285);
or U9636 (N_9636,N_9339,N_9409);
and U9637 (N_9637,N_9426,N_9294);
nand U9638 (N_9638,N_9263,N_9000);
xor U9639 (N_9639,N_9459,N_9429);
nand U9640 (N_9640,N_9358,N_9172);
and U9641 (N_9641,N_9028,N_9146);
and U9642 (N_9642,N_9337,N_9314);
xor U9643 (N_9643,N_9208,N_9414);
and U9644 (N_9644,N_9398,N_9170);
and U9645 (N_9645,N_9350,N_9035);
nor U9646 (N_9646,N_9067,N_9071);
and U9647 (N_9647,N_9341,N_9213);
nor U9648 (N_9648,N_9236,N_9195);
and U9649 (N_9649,N_9275,N_9009);
nor U9650 (N_9650,N_9377,N_9389);
xor U9651 (N_9651,N_9365,N_9245);
nor U9652 (N_9652,N_9325,N_9131);
nor U9653 (N_9653,N_9268,N_9005);
nand U9654 (N_9654,N_9123,N_9395);
or U9655 (N_9655,N_9438,N_9082);
and U9656 (N_9656,N_9368,N_9168);
or U9657 (N_9657,N_9315,N_9283);
xnor U9658 (N_9658,N_9312,N_9058);
nand U9659 (N_9659,N_9140,N_9047);
and U9660 (N_9660,N_9386,N_9241);
xnor U9661 (N_9661,N_9232,N_9125);
nor U9662 (N_9662,N_9329,N_9061);
nand U9663 (N_9663,N_9342,N_9088);
nor U9664 (N_9664,N_9243,N_9454);
and U9665 (N_9665,N_9157,N_9118);
or U9666 (N_9666,N_9194,N_9091);
xor U9667 (N_9667,N_9472,N_9015);
xnor U9668 (N_9668,N_9345,N_9100);
nand U9669 (N_9669,N_9226,N_9295);
nor U9670 (N_9670,N_9078,N_9387);
nor U9671 (N_9671,N_9102,N_9449);
or U9672 (N_9672,N_9032,N_9392);
nor U9673 (N_9673,N_9480,N_9330);
xor U9674 (N_9674,N_9124,N_9417);
and U9675 (N_9675,N_9117,N_9079);
nor U9676 (N_9676,N_9421,N_9020);
nand U9677 (N_9677,N_9228,N_9347);
nor U9678 (N_9678,N_9282,N_9496);
or U9679 (N_9679,N_9134,N_9246);
nand U9680 (N_9680,N_9445,N_9289);
nor U9681 (N_9681,N_9327,N_9281);
nor U9682 (N_9682,N_9466,N_9287);
nand U9683 (N_9683,N_9224,N_9469);
nand U9684 (N_9684,N_9029,N_9169);
and U9685 (N_9685,N_9013,N_9463);
and U9686 (N_9686,N_9428,N_9424);
or U9687 (N_9687,N_9187,N_9216);
xnor U9688 (N_9688,N_9338,N_9115);
nand U9689 (N_9689,N_9447,N_9462);
or U9690 (N_9690,N_9083,N_9199);
or U9691 (N_9691,N_9001,N_9151);
xnor U9692 (N_9692,N_9024,N_9062);
and U9693 (N_9693,N_9113,N_9101);
and U9694 (N_9694,N_9471,N_9284);
xnor U9695 (N_9695,N_9491,N_9264);
nor U9696 (N_9696,N_9349,N_9455);
xor U9697 (N_9697,N_9419,N_9402);
nor U9698 (N_9698,N_9155,N_9257);
or U9699 (N_9699,N_9112,N_9374);
nor U9700 (N_9700,N_9075,N_9136);
nor U9701 (N_9701,N_9014,N_9006);
nand U9702 (N_9702,N_9244,N_9388);
nand U9703 (N_9703,N_9156,N_9482);
xnor U9704 (N_9704,N_9050,N_9021);
nor U9705 (N_9705,N_9497,N_9012);
and U9706 (N_9706,N_9269,N_9311);
nor U9707 (N_9707,N_9004,N_9036);
nand U9708 (N_9708,N_9201,N_9404);
or U9709 (N_9709,N_9400,N_9052);
xor U9710 (N_9710,N_9178,N_9008);
or U9711 (N_9711,N_9193,N_9051);
or U9712 (N_9712,N_9147,N_9460);
and U9713 (N_9713,N_9444,N_9310);
or U9714 (N_9714,N_9420,N_9351);
xor U9715 (N_9715,N_9254,N_9286);
and U9716 (N_9716,N_9185,N_9080);
and U9717 (N_9717,N_9031,N_9152);
nor U9718 (N_9718,N_9104,N_9097);
or U9719 (N_9719,N_9119,N_9048);
nand U9720 (N_9720,N_9142,N_9378);
xor U9721 (N_9721,N_9434,N_9304);
and U9722 (N_9722,N_9293,N_9037);
nor U9723 (N_9723,N_9366,N_9390);
nor U9724 (N_9724,N_9486,N_9179);
and U9725 (N_9725,N_9196,N_9227);
nand U9726 (N_9726,N_9234,N_9221);
and U9727 (N_9727,N_9087,N_9407);
nor U9728 (N_9728,N_9166,N_9333);
xnor U9729 (N_9729,N_9018,N_9340);
nand U9730 (N_9730,N_9303,N_9266);
nand U9731 (N_9731,N_9138,N_9309);
or U9732 (N_9732,N_9074,N_9441);
nand U9733 (N_9733,N_9128,N_9474);
nand U9734 (N_9734,N_9308,N_9129);
xor U9735 (N_9735,N_9435,N_9096);
nand U9736 (N_9736,N_9038,N_9120);
or U9737 (N_9737,N_9494,N_9153);
or U9738 (N_9738,N_9027,N_9363);
nand U9739 (N_9739,N_9030,N_9127);
or U9740 (N_9740,N_9302,N_9076);
or U9741 (N_9741,N_9317,N_9171);
nand U9742 (N_9742,N_9159,N_9160);
and U9743 (N_9743,N_9375,N_9476);
and U9744 (N_9744,N_9202,N_9451);
or U9745 (N_9745,N_9007,N_9355);
xor U9746 (N_9746,N_9305,N_9186);
nand U9747 (N_9747,N_9237,N_9231);
xnor U9748 (N_9748,N_9219,N_9276);
or U9749 (N_9749,N_9161,N_9188);
nand U9750 (N_9750,N_9171,N_9335);
nor U9751 (N_9751,N_9038,N_9162);
nor U9752 (N_9752,N_9115,N_9074);
or U9753 (N_9753,N_9342,N_9035);
nor U9754 (N_9754,N_9298,N_9110);
nor U9755 (N_9755,N_9044,N_9007);
nand U9756 (N_9756,N_9277,N_9204);
nor U9757 (N_9757,N_9326,N_9018);
nand U9758 (N_9758,N_9229,N_9064);
xor U9759 (N_9759,N_9072,N_9032);
or U9760 (N_9760,N_9129,N_9164);
xnor U9761 (N_9761,N_9175,N_9199);
and U9762 (N_9762,N_9475,N_9487);
xor U9763 (N_9763,N_9128,N_9201);
nor U9764 (N_9764,N_9202,N_9160);
or U9765 (N_9765,N_9148,N_9138);
xor U9766 (N_9766,N_9327,N_9050);
nand U9767 (N_9767,N_9039,N_9458);
nand U9768 (N_9768,N_9284,N_9480);
nor U9769 (N_9769,N_9400,N_9331);
xor U9770 (N_9770,N_9102,N_9012);
nor U9771 (N_9771,N_9346,N_9106);
xnor U9772 (N_9772,N_9162,N_9196);
nor U9773 (N_9773,N_9027,N_9441);
or U9774 (N_9774,N_9462,N_9326);
xnor U9775 (N_9775,N_9362,N_9363);
and U9776 (N_9776,N_9145,N_9042);
or U9777 (N_9777,N_9449,N_9148);
xor U9778 (N_9778,N_9024,N_9232);
xor U9779 (N_9779,N_9218,N_9086);
xor U9780 (N_9780,N_9406,N_9147);
nand U9781 (N_9781,N_9385,N_9020);
nor U9782 (N_9782,N_9299,N_9239);
nand U9783 (N_9783,N_9067,N_9288);
nor U9784 (N_9784,N_9282,N_9056);
nor U9785 (N_9785,N_9371,N_9242);
xnor U9786 (N_9786,N_9234,N_9231);
nor U9787 (N_9787,N_9219,N_9095);
nand U9788 (N_9788,N_9150,N_9411);
or U9789 (N_9789,N_9372,N_9257);
xor U9790 (N_9790,N_9430,N_9119);
nand U9791 (N_9791,N_9208,N_9345);
xor U9792 (N_9792,N_9246,N_9175);
or U9793 (N_9793,N_9458,N_9010);
or U9794 (N_9794,N_9356,N_9190);
xnor U9795 (N_9795,N_9237,N_9378);
xor U9796 (N_9796,N_9282,N_9101);
and U9797 (N_9797,N_9136,N_9308);
nor U9798 (N_9798,N_9203,N_9498);
xnor U9799 (N_9799,N_9215,N_9387);
xnor U9800 (N_9800,N_9319,N_9402);
and U9801 (N_9801,N_9305,N_9406);
and U9802 (N_9802,N_9346,N_9031);
nand U9803 (N_9803,N_9326,N_9339);
and U9804 (N_9804,N_9300,N_9380);
nor U9805 (N_9805,N_9431,N_9191);
and U9806 (N_9806,N_9084,N_9246);
nor U9807 (N_9807,N_9337,N_9090);
and U9808 (N_9808,N_9017,N_9336);
nor U9809 (N_9809,N_9217,N_9335);
nand U9810 (N_9810,N_9027,N_9224);
xnor U9811 (N_9811,N_9224,N_9396);
and U9812 (N_9812,N_9000,N_9328);
nor U9813 (N_9813,N_9341,N_9496);
nor U9814 (N_9814,N_9331,N_9144);
nand U9815 (N_9815,N_9441,N_9377);
or U9816 (N_9816,N_9382,N_9169);
nor U9817 (N_9817,N_9461,N_9165);
nand U9818 (N_9818,N_9216,N_9337);
and U9819 (N_9819,N_9028,N_9054);
nand U9820 (N_9820,N_9180,N_9063);
nand U9821 (N_9821,N_9019,N_9013);
nand U9822 (N_9822,N_9435,N_9355);
and U9823 (N_9823,N_9196,N_9028);
nand U9824 (N_9824,N_9475,N_9397);
xor U9825 (N_9825,N_9270,N_9282);
nor U9826 (N_9826,N_9419,N_9285);
or U9827 (N_9827,N_9395,N_9057);
or U9828 (N_9828,N_9171,N_9447);
xor U9829 (N_9829,N_9173,N_9351);
xnor U9830 (N_9830,N_9178,N_9260);
nor U9831 (N_9831,N_9111,N_9318);
xor U9832 (N_9832,N_9303,N_9325);
and U9833 (N_9833,N_9485,N_9386);
nand U9834 (N_9834,N_9478,N_9285);
and U9835 (N_9835,N_9196,N_9354);
and U9836 (N_9836,N_9494,N_9365);
nor U9837 (N_9837,N_9414,N_9174);
or U9838 (N_9838,N_9365,N_9166);
or U9839 (N_9839,N_9215,N_9398);
nand U9840 (N_9840,N_9459,N_9013);
or U9841 (N_9841,N_9474,N_9472);
xnor U9842 (N_9842,N_9120,N_9148);
nand U9843 (N_9843,N_9245,N_9434);
nor U9844 (N_9844,N_9142,N_9120);
nor U9845 (N_9845,N_9105,N_9261);
and U9846 (N_9846,N_9444,N_9405);
and U9847 (N_9847,N_9487,N_9082);
nor U9848 (N_9848,N_9416,N_9075);
or U9849 (N_9849,N_9361,N_9424);
nand U9850 (N_9850,N_9393,N_9380);
and U9851 (N_9851,N_9040,N_9344);
nand U9852 (N_9852,N_9041,N_9326);
or U9853 (N_9853,N_9208,N_9419);
xor U9854 (N_9854,N_9013,N_9187);
or U9855 (N_9855,N_9438,N_9222);
nand U9856 (N_9856,N_9481,N_9420);
nor U9857 (N_9857,N_9046,N_9103);
or U9858 (N_9858,N_9487,N_9443);
xnor U9859 (N_9859,N_9285,N_9160);
nand U9860 (N_9860,N_9433,N_9406);
or U9861 (N_9861,N_9459,N_9079);
and U9862 (N_9862,N_9224,N_9449);
nor U9863 (N_9863,N_9492,N_9279);
xor U9864 (N_9864,N_9203,N_9033);
nor U9865 (N_9865,N_9042,N_9343);
nand U9866 (N_9866,N_9458,N_9001);
and U9867 (N_9867,N_9121,N_9321);
xor U9868 (N_9868,N_9005,N_9261);
xnor U9869 (N_9869,N_9148,N_9102);
xnor U9870 (N_9870,N_9200,N_9321);
or U9871 (N_9871,N_9032,N_9281);
and U9872 (N_9872,N_9209,N_9200);
xnor U9873 (N_9873,N_9195,N_9225);
nor U9874 (N_9874,N_9307,N_9291);
xnor U9875 (N_9875,N_9129,N_9416);
or U9876 (N_9876,N_9263,N_9302);
nor U9877 (N_9877,N_9112,N_9337);
or U9878 (N_9878,N_9311,N_9232);
xnor U9879 (N_9879,N_9268,N_9214);
and U9880 (N_9880,N_9161,N_9192);
nor U9881 (N_9881,N_9251,N_9041);
and U9882 (N_9882,N_9023,N_9093);
and U9883 (N_9883,N_9048,N_9111);
and U9884 (N_9884,N_9032,N_9444);
nand U9885 (N_9885,N_9230,N_9221);
or U9886 (N_9886,N_9100,N_9333);
or U9887 (N_9887,N_9364,N_9372);
nor U9888 (N_9888,N_9352,N_9016);
or U9889 (N_9889,N_9359,N_9356);
xnor U9890 (N_9890,N_9187,N_9346);
or U9891 (N_9891,N_9495,N_9073);
nor U9892 (N_9892,N_9067,N_9489);
and U9893 (N_9893,N_9092,N_9029);
xor U9894 (N_9894,N_9343,N_9028);
and U9895 (N_9895,N_9239,N_9159);
or U9896 (N_9896,N_9315,N_9162);
xor U9897 (N_9897,N_9434,N_9378);
xor U9898 (N_9898,N_9499,N_9393);
and U9899 (N_9899,N_9100,N_9316);
nor U9900 (N_9900,N_9183,N_9010);
and U9901 (N_9901,N_9196,N_9261);
nor U9902 (N_9902,N_9227,N_9370);
nand U9903 (N_9903,N_9006,N_9209);
nor U9904 (N_9904,N_9022,N_9476);
nand U9905 (N_9905,N_9058,N_9242);
nor U9906 (N_9906,N_9273,N_9068);
nor U9907 (N_9907,N_9250,N_9428);
or U9908 (N_9908,N_9281,N_9191);
or U9909 (N_9909,N_9391,N_9001);
xor U9910 (N_9910,N_9074,N_9435);
and U9911 (N_9911,N_9421,N_9473);
nor U9912 (N_9912,N_9121,N_9098);
nand U9913 (N_9913,N_9323,N_9181);
nor U9914 (N_9914,N_9049,N_9365);
and U9915 (N_9915,N_9131,N_9420);
or U9916 (N_9916,N_9080,N_9358);
xor U9917 (N_9917,N_9252,N_9103);
and U9918 (N_9918,N_9427,N_9218);
nand U9919 (N_9919,N_9464,N_9044);
nor U9920 (N_9920,N_9008,N_9495);
or U9921 (N_9921,N_9253,N_9219);
xor U9922 (N_9922,N_9304,N_9126);
or U9923 (N_9923,N_9232,N_9398);
and U9924 (N_9924,N_9242,N_9173);
nor U9925 (N_9925,N_9153,N_9224);
xnor U9926 (N_9926,N_9454,N_9409);
and U9927 (N_9927,N_9032,N_9001);
and U9928 (N_9928,N_9481,N_9020);
xnor U9929 (N_9929,N_9095,N_9210);
xnor U9930 (N_9930,N_9159,N_9299);
or U9931 (N_9931,N_9157,N_9115);
xor U9932 (N_9932,N_9347,N_9422);
nand U9933 (N_9933,N_9193,N_9415);
and U9934 (N_9934,N_9380,N_9460);
and U9935 (N_9935,N_9380,N_9478);
nand U9936 (N_9936,N_9202,N_9016);
xor U9937 (N_9937,N_9442,N_9487);
or U9938 (N_9938,N_9301,N_9200);
xor U9939 (N_9939,N_9162,N_9337);
and U9940 (N_9940,N_9138,N_9104);
nor U9941 (N_9941,N_9232,N_9340);
xnor U9942 (N_9942,N_9088,N_9294);
and U9943 (N_9943,N_9477,N_9205);
nor U9944 (N_9944,N_9348,N_9361);
or U9945 (N_9945,N_9463,N_9215);
or U9946 (N_9946,N_9036,N_9427);
or U9947 (N_9947,N_9125,N_9395);
nand U9948 (N_9948,N_9263,N_9444);
and U9949 (N_9949,N_9226,N_9012);
xor U9950 (N_9950,N_9088,N_9276);
or U9951 (N_9951,N_9306,N_9344);
nor U9952 (N_9952,N_9120,N_9029);
nor U9953 (N_9953,N_9147,N_9127);
and U9954 (N_9954,N_9113,N_9490);
and U9955 (N_9955,N_9149,N_9087);
and U9956 (N_9956,N_9012,N_9480);
or U9957 (N_9957,N_9022,N_9432);
xnor U9958 (N_9958,N_9336,N_9498);
or U9959 (N_9959,N_9034,N_9067);
nand U9960 (N_9960,N_9489,N_9449);
xnor U9961 (N_9961,N_9294,N_9429);
nand U9962 (N_9962,N_9104,N_9388);
and U9963 (N_9963,N_9139,N_9146);
nand U9964 (N_9964,N_9129,N_9065);
and U9965 (N_9965,N_9195,N_9241);
nand U9966 (N_9966,N_9147,N_9308);
and U9967 (N_9967,N_9182,N_9360);
nor U9968 (N_9968,N_9158,N_9464);
or U9969 (N_9969,N_9490,N_9084);
or U9970 (N_9970,N_9112,N_9409);
nand U9971 (N_9971,N_9158,N_9127);
or U9972 (N_9972,N_9112,N_9147);
and U9973 (N_9973,N_9390,N_9016);
or U9974 (N_9974,N_9314,N_9164);
nor U9975 (N_9975,N_9044,N_9497);
xnor U9976 (N_9976,N_9320,N_9073);
nand U9977 (N_9977,N_9018,N_9369);
and U9978 (N_9978,N_9427,N_9103);
or U9979 (N_9979,N_9333,N_9158);
xnor U9980 (N_9980,N_9243,N_9141);
and U9981 (N_9981,N_9252,N_9232);
xor U9982 (N_9982,N_9293,N_9123);
nor U9983 (N_9983,N_9017,N_9240);
nor U9984 (N_9984,N_9147,N_9369);
xnor U9985 (N_9985,N_9319,N_9347);
nor U9986 (N_9986,N_9477,N_9281);
xor U9987 (N_9987,N_9377,N_9250);
nand U9988 (N_9988,N_9145,N_9038);
and U9989 (N_9989,N_9228,N_9036);
nand U9990 (N_9990,N_9196,N_9268);
nand U9991 (N_9991,N_9452,N_9292);
nand U9992 (N_9992,N_9069,N_9317);
nand U9993 (N_9993,N_9413,N_9376);
xor U9994 (N_9994,N_9425,N_9216);
nand U9995 (N_9995,N_9222,N_9140);
or U9996 (N_9996,N_9115,N_9006);
xnor U9997 (N_9997,N_9351,N_9090);
xor U9998 (N_9998,N_9300,N_9075);
nor U9999 (N_9999,N_9460,N_9309);
or U10000 (N_10000,N_9508,N_9979);
nor U10001 (N_10001,N_9983,N_9779);
nand U10002 (N_10002,N_9907,N_9861);
or U10003 (N_10003,N_9692,N_9858);
xnor U10004 (N_10004,N_9984,N_9518);
xor U10005 (N_10005,N_9723,N_9596);
or U10006 (N_10006,N_9856,N_9994);
nand U10007 (N_10007,N_9580,N_9737);
xnor U10008 (N_10008,N_9604,N_9756);
and U10009 (N_10009,N_9838,N_9965);
nor U10010 (N_10010,N_9662,N_9993);
or U10011 (N_10011,N_9587,N_9699);
nand U10012 (N_10012,N_9786,N_9813);
xnor U10013 (N_10013,N_9908,N_9682);
or U10014 (N_10014,N_9768,N_9828);
or U10015 (N_10015,N_9539,N_9797);
nor U10016 (N_10016,N_9741,N_9793);
nor U10017 (N_10017,N_9796,N_9778);
nor U10018 (N_10018,N_9640,N_9873);
nor U10019 (N_10019,N_9666,N_9591);
xor U10020 (N_10020,N_9749,N_9782);
nand U10021 (N_10021,N_9601,N_9523);
nand U10022 (N_10022,N_9857,N_9981);
and U10023 (N_10023,N_9693,N_9829);
or U10024 (N_10024,N_9930,N_9760);
or U10025 (N_10025,N_9509,N_9597);
xnor U10026 (N_10026,N_9775,N_9663);
nand U10027 (N_10027,N_9744,N_9568);
nor U10028 (N_10028,N_9678,N_9985);
nor U10029 (N_10029,N_9649,N_9854);
or U10030 (N_10030,N_9578,N_9641);
or U10031 (N_10031,N_9689,N_9690);
and U10032 (N_10032,N_9761,N_9524);
xnor U10033 (N_10033,N_9812,N_9927);
nor U10034 (N_10034,N_9842,N_9619);
and U10035 (N_10035,N_9996,N_9574);
nor U10036 (N_10036,N_9819,N_9680);
nand U10037 (N_10037,N_9999,N_9872);
nand U10038 (N_10038,N_9507,N_9977);
and U10039 (N_10039,N_9562,N_9814);
and U10040 (N_10040,N_9738,N_9705);
and U10041 (N_10041,N_9918,N_9841);
xnor U10042 (N_10042,N_9948,N_9939);
or U10043 (N_10043,N_9957,N_9708);
nor U10044 (N_10044,N_9929,N_9638);
or U10045 (N_10045,N_9909,N_9825);
or U10046 (N_10046,N_9516,N_9694);
xnor U10047 (N_10047,N_9946,N_9544);
or U10048 (N_10048,N_9571,N_9794);
nand U10049 (N_10049,N_9631,N_9664);
and U10050 (N_10050,N_9774,N_9679);
nand U10051 (N_10051,N_9661,N_9792);
nand U10052 (N_10052,N_9754,N_9955);
or U10053 (N_10053,N_9890,N_9790);
or U10054 (N_10054,N_9731,N_9942);
xnor U10055 (N_10055,N_9881,N_9968);
xor U10056 (N_10056,N_9743,N_9709);
nor U10057 (N_10057,N_9729,N_9555);
or U10058 (N_10058,N_9520,N_9755);
xor U10059 (N_10059,N_9765,N_9733);
xnor U10060 (N_10060,N_9644,N_9506);
nand U10061 (N_10061,N_9855,N_9657);
and U10062 (N_10062,N_9916,N_9952);
nand U10063 (N_10063,N_9982,N_9620);
nor U10064 (N_10064,N_9746,N_9800);
nand U10065 (N_10065,N_9944,N_9906);
nand U10066 (N_10066,N_9951,N_9630);
nor U10067 (N_10067,N_9770,N_9845);
or U10068 (N_10068,N_9933,N_9889);
nor U10069 (N_10069,N_9833,N_9914);
xor U10070 (N_10070,N_9608,N_9745);
nand U10071 (N_10071,N_9931,N_9712);
or U10072 (N_10072,N_9700,N_9886);
nor U10073 (N_10073,N_9972,N_9964);
and U10074 (N_10074,N_9599,N_9923);
nand U10075 (N_10075,N_9553,N_9725);
nand U10076 (N_10076,N_9541,N_9691);
or U10077 (N_10077,N_9766,N_9896);
nor U10078 (N_10078,N_9522,N_9538);
nor U10079 (N_10079,N_9818,N_9799);
xnor U10080 (N_10080,N_9897,N_9710);
or U10081 (N_10081,N_9980,N_9988);
nand U10082 (N_10082,N_9787,N_9877);
xor U10083 (N_10083,N_9767,N_9559);
nand U10084 (N_10084,N_9961,N_9667);
nand U10085 (N_10085,N_9827,N_9598);
and U10086 (N_10086,N_9875,N_9997);
or U10087 (N_10087,N_9688,N_9515);
xor U10088 (N_10088,N_9922,N_9893);
nor U10089 (N_10089,N_9910,N_9502);
xnor U10090 (N_10090,N_9764,N_9973);
xnor U10091 (N_10091,N_9891,N_9917);
xor U10092 (N_10092,N_9780,N_9565);
nand U10093 (N_10093,N_9773,N_9570);
nand U10094 (N_10094,N_9535,N_9521);
nand U10095 (N_10095,N_9730,N_9592);
and U10096 (N_10096,N_9703,N_9920);
and U10097 (N_10097,N_9593,N_9724);
nand U10098 (N_10098,N_9898,N_9995);
nand U10099 (N_10099,N_9880,N_9668);
and U10100 (N_10100,N_9545,N_9576);
xor U10101 (N_10101,N_9614,N_9823);
and U10102 (N_10102,N_9788,N_9647);
or U10103 (N_10103,N_9938,N_9659);
or U10104 (N_10104,N_9622,N_9525);
and U10105 (N_10105,N_9573,N_9528);
nand U10106 (N_10106,N_9653,N_9763);
xnor U10107 (N_10107,N_9721,N_9899);
xor U10108 (N_10108,N_9505,N_9816);
nor U10109 (N_10109,N_9696,N_9554);
nand U10110 (N_10110,N_9637,N_9950);
nor U10111 (N_10111,N_9656,N_9707);
nor U10112 (N_10112,N_9966,N_9847);
or U10113 (N_10113,N_9783,N_9830);
or U10114 (N_10114,N_9815,N_9956);
xor U10115 (N_10115,N_9990,N_9808);
and U10116 (N_10116,N_9824,N_9903);
and U10117 (N_10117,N_9963,N_9804);
or U10118 (N_10118,N_9697,N_9879);
xnor U10119 (N_10119,N_9626,N_9716);
xor U10120 (N_10120,N_9671,N_9998);
or U10121 (N_10121,N_9711,N_9684);
xnor U10122 (N_10122,N_9600,N_9660);
xnor U10123 (N_10123,N_9549,N_9581);
nand U10124 (N_10124,N_9953,N_9967);
and U10125 (N_10125,N_9962,N_9567);
and U10126 (N_10126,N_9915,N_9747);
nor U10127 (N_10127,N_9894,N_9859);
xnor U10128 (N_10128,N_9695,N_9655);
and U10129 (N_10129,N_9844,N_9865);
and U10130 (N_10130,N_9577,N_9586);
nor U10131 (N_10131,N_9551,N_9607);
or U10132 (N_10132,N_9878,N_9902);
nand U10133 (N_10133,N_9612,N_9905);
xnor U10134 (N_10134,N_9613,N_9552);
or U10135 (N_10135,N_9719,N_9795);
nand U10136 (N_10136,N_9532,N_9750);
nand U10137 (N_10137,N_9851,N_9685);
or U10138 (N_10138,N_9687,N_9978);
nor U10139 (N_10139,N_9513,N_9821);
and U10140 (N_10140,N_9740,N_9869);
nor U10141 (N_10141,N_9739,N_9771);
and U10142 (N_10142,N_9543,N_9540);
xnor U10143 (N_10143,N_9868,N_9807);
nor U10144 (N_10144,N_9588,N_9843);
or U10145 (N_10145,N_9860,N_9569);
and U10146 (N_10146,N_9585,N_9547);
xor U10147 (N_10147,N_9548,N_9820);
xnor U10148 (N_10148,N_9706,N_9654);
xnor U10149 (N_10149,N_9672,N_9883);
nand U10150 (N_10150,N_9840,N_9866);
or U10151 (N_10151,N_9803,N_9987);
xor U10152 (N_10152,N_9633,N_9558);
xor U10153 (N_10153,N_9960,N_9514);
or U10154 (N_10154,N_9769,N_9701);
or U10155 (N_10155,N_9669,N_9752);
xnor U10156 (N_10156,N_9628,N_9992);
xor U10157 (N_10157,N_9512,N_9947);
or U10158 (N_10158,N_9674,N_9564);
xor U10159 (N_10159,N_9623,N_9718);
or U10160 (N_10160,N_9913,N_9853);
or U10161 (N_10161,N_9615,N_9537);
or U10162 (N_10162,N_9959,N_9584);
and U10163 (N_10163,N_9651,N_9810);
and U10164 (N_10164,N_9885,N_9791);
or U10165 (N_10165,N_9609,N_9734);
nand U10166 (N_10166,N_9645,N_9610);
or U10167 (N_10167,N_9757,N_9759);
xnor U10168 (N_10168,N_9686,N_9876);
or U10169 (N_10169,N_9676,N_9949);
nor U10170 (N_10170,N_9556,N_9811);
nand U10171 (N_10171,N_9579,N_9753);
and U10172 (N_10172,N_9937,N_9683);
and U10173 (N_10173,N_9904,N_9673);
xor U10174 (N_10174,N_9932,N_9594);
xnor U10175 (N_10175,N_9720,N_9958);
nor U10176 (N_10176,N_9789,N_9943);
nor U10177 (N_10177,N_9945,N_9919);
and U10178 (N_10178,N_9636,N_9777);
nand U10179 (N_10179,N_9561,N_9560);
nand U10180 (N_10180,N_9715,N_9975);
and U10181 (N_10181,N_9895,N_9971);
xor U10182 (N_10182,N_9642,N_9940);
nand U10183 (N_10183,N_9806,N_9846);
nand U10184 (N_10184,N_9563,N_9530);
xor U10185 (N_10185,N_9801,N_9665);
and U10186 (N_10186,N_9590,N_9546);
nor U10187 (N_10187,N_9617,N_9802);
nand U10188 (N_10188,N_9582,N_9575);
xnor U10189 (N_10189,N_9618,N_9698);
xnor U10190 (N_10190,N_9536,N_9643);
and U10191 (N_10191,N_9650,N_9784);
xor U10192 (N_10192,N_9924,N_9837);
nand U10193 (N_10193,N_9510,N_9928);
nor U10194 (N_10194,N_9798,N_9911);
nor U10195 (N_10195,N_9751,N_9542);
or U10196 (N_10196,N_9602,N_9566);
nand U10197 (N_10197,N_9834,N_9503);
nor U10198 (N_10198,N_9635,N_9864);
xor U10199 (N_10199,N_9557,N_9519);
nand U10200 (N_10200,N_9921,N_9627);
xnor U10201 (N_10201,N_9974,N_9785);
nor U10202 (N_10202,N_9531,N_9595);
and U10203 (N_10203,N_9926,N_9836);
nand U10204 (N_10204,N_9639,N_9986);
or U10205 (N_10205,N_9871,N_9634);
or U10206 (N_10206,N_9742,N_9714);
and U10207 (N_10207,N_9629,N_9605);
xor U10208 (N_10208,N_9572,N_9772);
nand U10209 (N_10209,N_9735,N_9658);
or U10210 (N_10210,N_9504,N_9762);
and U10211 (N_10211,N_9511,N_9648);
nand U10212 (N_10212,N_9781,N_9934);
nor U10213 (N_10213,N_9884,N_9526);
nor U10214 (N_10214,N_9809,N_9500);
and U10215 (N_10215,N_9728,N_9862);
nor U10216 (N_10216,N_9534,N_9870);
nor U10217 (N_10217,N_9941,N_9533);
nor U10218 (N_10218,N_9727,N_9702);
xnor U10219 (N_10219,N_9874,N_9849);
nor U10220 (N_10220,N_9970,N_9646);
nand U10221 (N_10221,N_9529,N_9887);
or U10222 (N_10222,N_9776,N_9826);
nor U10223 (N_10223,N_9863,N_9748);
nand U10224 (N_10224,N_9758,N_9722);
nor U10225 (N_10225,N_9589,N_9717);
nand U10226 (N_10226,N_9912,N_9832);
and U10227 (N_10227,N_9583,N_9527);
or U10228 (N_10228,N_9704,N_9892);
nand U10229 (N_10229,N_9611,N_9850);
xor U10230 (N_10230,N_9675,N_9839);
nand U10231 (N_10231,N_9726,N_9848);
xor U10232 (N_10232,N_9991,N_9831);
nand U10233 (N_10233,N_9736,N_9817);
nor U10234 (N_10234,N_9805,N_9901);
nor U10235 (N_10235,N_9517,N_9835);
nand U10236 (N_10236,N_9550,N_9616);
and U10237 (N_10237,N_9925,N_9732);
or U10238 (N_10238,N_9677,N_9900);
xor U10239 (N_10239,N_9935,N_9822);
xnor U10240 (N_10240,N_9976,N_9713);
and U10241 (N_10241,N_9625,N_9621);
and U10242 (N_10242,N_9969,N_9670);
and U10243 (N_10243,N_9624,N_9867);
nand U10244 (N_10244,N_9888,N_9501);
or U10245 (N_10245,N_9606,N_9954);
nand U10246 (N_10246,N_9989,N_9681);
or U10247 (N_10247,N_9936,N_9882);
or U10248 (N_10248,N_9852,N_9603);
and U10249 (N_10249,N_9632,N_9652);
or U10250 (N_10250,N_9780,N_9625);
or U10251 (N_10251,N_9756,N_9534);
or U10252 (N_10252,N_9884,N_9506);
nor U10253 (N_10253,N_9757,N_9755);
xor U10254 (N_10254,N_9642,N_9973);
xnor U10255 (N_10255,N_9874,N_9721);
nor U10256 (N_10256,N_9995,N_9996);
nor U10257 (N_10257,N_9765,N_9609);
xnor U10258 (N_10258,N_9751,N_9975);
nand U10259 (N_10259,N_9554,N_9505);
or U10260 (N_10260,N_9691,N_9854);
or U10261 (N_10261,N_9867,N_9884);
and U10262 (N_10262,N_9587,N_9950);
and U10263 (N_10263,N_9647,N_9925);
and U10264 (N_10264,N_9693,N_9676);
or U10265 (N_10265,N_9591,N_9765);
nor U10266 (N_10266,N_9900,N_9505);
xor U10267 (N_10267,N_9809,N_9768);
and U10268 (N_10268,N_9602,N_9648);
and U10269 (N_10269,N_9984,N_9719);
nand U10270 (N_10270,N_9996,N_9910);
xnor U10271 (N_10271,N_9530,N_9965);
and U10272 (N_10272,N_9657,N_9928);
xnor U10273 (N_10273,N_9637,N_9985);
or U10274 (N_10274,N_9645,N_9891);
and U10275 (N_10275,N_9506,N_9648);
nor U10276 (N_10276,N_9839,N_9832);
xnor U10277 (N_10277,N_9732,N_9991);
and U10278 (N_10278,N_9583,N_9743);
nand U10279 (N_10279,N_9546,N_9691);
or U10280 (N_10280,N_9556,N_9673);
nor U10281 (N_10281,N_9983,N_9584);
or U10282 (N_10282,N_9816,N_9869);
or U10283 (N_10283,N_9781,N_9850);
nand U10284 (N_10284,N_9508,N_9929);
nand U10285 (N_10285,N_9977,N_9645);
nor U10286 (N_10286,N_9698,N_9846);
nand U10287 (N_10287,N_9925,N_9566);
xor U10288 (N_10288,N_9795,N_9811);
xnor U10289 (N_10289,N_9607,N_9585);
and U10290 (N_10290,N_9900,N_9873);
nand U10291 (N_10291,N_9869,N_9936);
and U10292 (N_10292,N_9670,N_9728);
xor U10293 (N_10293,N_9801,N_9659);
nor U10294 (N_10294,N_9795,N_9618);
nand U10295 (N_10295,N_9679,N_9507);
and U10296 (N_10296,N_9554,N_9851);
nand U10297 (N_10297,N_9856,N_9761);
nand U10298 (N_10298,N_9598,N_9968);
nand U10299 (N_10299,N_9965,N_9920);
xnor U10300 (N_10300,N_9518,N_9557);
nand U10301 (N_10301,N_9622,N_9978);
xor U10302 (N_10302,N_9837,N_9912);
nand U10303 (N_10303,N_9869,N_9917);
or U10304 (N_10304,N_9879,N_9514);
nor U10305 (N_10305,N_9895,N_9966);
or U10306 (N_10306,N_9570,N_9590);
nor U10307 (N_10307,N_9794,N_9757);
or U10308 (N_10308,N_9999,N_9861);
nand U10309 (N_10309,N_9612,N_9832);
and U10310 (N_10310,N_9803,N_9820);
or U10311 (N_10311,N_9835,N_9647);
xnor U10312 (N_10312,N_9917,N_9728);
nand U10313 (N_10313,N_9875,N_9859);
or U10314 (N_10314,N_9671,N_9667);
nand U10315 (N_10315,N_9591,N_9584);
or U10316 (N_10316,N_9610,N_9990);
or U10317 (N_10317,N_9597,N_9810);
or U10318 (N_10318,N_9809,N_9886);
nand U10319 (N_10319,N_9868,N_9942);
nor U10320 (N_10320,N_9533,N_9539);
nand U10321 (N_10321,N_9983,N_9822);
and U10322 (N_10322,N_9534,N_9862);
or U10323 (N_10323,N_9972,N_9676);
or U10324 (N_10324,N_9689,N_9826);
or U10325 (N_10325,N_9676,N_9833);
nor U10326 (N_10326,N_9617,N_9845);
and U10327 (N_10327,N_9531,N_9750);
nand U10328 (N_10328,N_9535,N_9675);
and U10329 (N_10329,N_9608,N_9964);
and U10330 (N_10330,N_9802,N_9583);
or U10331 (N_10331,N_9613,N_9621);
and U10332 (N_10332,N_9678,N_9785);
xnor U10333 (N_10333,N_9674,N_9802);
or U10334 (N_10334,N_9718,N_9770);
nand U10335 (N_10335,N_9961,N_9639);
and U10336 (N_10336,N_9739,N_9939);
xnor U10337 (N_10337,N_9601,N_9737);
xnor U10338 (N_10338,N_9961,N_9590);
and U10339 (N_10339,N_9559,N_9877);
and U10340 (N_10340,N_9878,N_9818);
xor U10341 (N_10341,N_9801,N_9903);
nand U10342 (N_10342,N_9713,N_9685);
or U10343 (N_10343,N_9891,N_9949);
nor U10344 (N_10344,N_9880,N_9778);
xor U10345 (N_10345,N_9552,N_9566);
or U10346 (N_10346,N_9588,N_9555);
or U10347 (N_10347,N_9566,N_9949);
and U10348 (N_10348,N_9621,N_9880);
xnor U10349 (N_10349,N_9877,N_9746);
xnor U10350 (N_10350,N_9647,N_9779);
and U10351 (N_10351,N_9557,N_9610);
nand U10352 (N_10352,N_9888,N_9570);
nand U10353 (N_10353,N_9934,N_9942);
nand U10354 (N_10354,N_9871,N_9509);
or U10355 (N_10355,N_9595,N_9680);
or U10356 (N_10356,N_9913,N_9575);
or U10357 (N_10357,N_9751,N_9533);
and U10358 (N_10358,N_9610,N_9981);
xnor U10359 (N_10359,N_9604,N_9905);
nor U10360 (N_10360,N_9884,N_9960);
nor U10361 (N_10361,N_9643,N_9770);
nor U10362 (N_10362,N_9594,N_9651);
nand U10363 (N_10363,N_9506,N_9921);
nor U10364 (N_10364,N_9559,N_9830);
and U10365 (N_10365,N_9626,N_9581);
and U10366 (N_10366,N_9977,N_9777);
or U10367 (N_10367,N_9514,N_9905);
nor U10368 (N_10368,N_9638,N_9697);
xor U10369 (N_10369,N_9773,N_9896);
or U10370 (N_10370,N_9596,N_9985);
or U10371 (N_10371,N_9878,N_9791);
xnor U10372 (N_10372,N_9972,N_9815);
or U10373 (N_10373,N_9614,N_9943);
nand U10374 (N_10374,N_9898,N_9996);
and U10375 (N_10375,N_9613,N_9834);
or U10376 (N_10376,N_9830,N_9881);
nor U10377 (N_10377,N_9945,N_9785);
and U10378 (N_10378,N_9741,N_9715);
or U10379 (N_10379,N_9727,N_9716);
nand U10380 (N_10380,N_9740,N_9894);
xor U10381 (N_10381,N_9873,N_9542);
and U10382 (N_10382,N_9947,N_9905);
nand U10383 (N_10383,N_9906,N_9782);
xor U10384 (N_10384,N_9756,N_9645);
or U10385 (N_10385,N_9647,N_9923);
and U10386 (N_10386,N_9848,N_9967);
or U10387 (N_10387,N_9611,N_9830);
and U10388 (N_10388,N_9814,N_9632);
xor U10389 (N_10389,N_9846,N_9624);
and U10390 (N_10390,N_9737,N_9597);
nor U10391 (N_10391,N_9599,N_9730);
xor U10392 (N_10392,N_9803,N_9611);
nand U10393 (N_10393,N_9715,N_9982);
and U10394 (N_10394,N_9557,N_9536);
and U10395 (N_10395,N_9529,N_9705);
or U10396 (N_10396,N_9729,N_9917);
nand U10397 (N_10397,N_9799,N_9777);
and U10398 (N_10398,N_9520,N_9869);
or U10399 (N_10399,N_9932,N_9939);
or U10400 (N_10400,N_9704,N_9732);
and U10401 (N_10401,N_9959,N_9756);
nor U10402 (N_10402,N_9927,N_9961);
nand U10403 (N_10403,N_9571,N_9721);
xor U10404 (N_10404,N_9500,N_9934);
and U10405 (N_10405,N_9953,N_9545);
xnor U10406 (N_10406,N_9942,N_9902);
nand U10407 (N_10407,N_9792,N_9659);
xnor U10408 (N_10408,N_9605,N_9792);
xnor U10409 (N_10409,N_9694,N_9596);
nand U10410 (N_10410,N_9509,N_9816);
nor U10411 (N_10411,N_9870,N_9837);
xnor U10412 (N_10412,N_9848,N_9604);
nor U10413 (N_10413,N_9891,N_9757);
nor U10414 (N_10414,N_9966,N_9528);
or U10415 (N_10415,N_9811,N_9608);
nand U10416 (N_10416,N_9656,N_9658);
nor U10417 (N_10417,N_9504,N_9734);
or U10418 (N_10418,N_9745,N_9740);
xnor U10419 (N_10419,N_9872,N_9541);
xnor U10420 (N_10420,N_9932,N_9683);
and U10421 (N_10421,N_9548,N_9813);
nand U10422 (N_10422,N_9659,N_9929);
or U10423 (N_10423,N_9759,N_9585);
nand U10424 (N_10424,N_9502,N_9505);
nand U10425 (N_10425,N_9646,N_9980);
and U10426 (N_10426,N_9674,N_9687);
nand U10427 (N_10427,N_9674,N_9636);
nor U10428 (N_10428,N_9999,N_9728);
nor U10429 (N_10429,N_9870,N_9617);
nand U10430 (N_10430,N_9644,N_9714);
or U10431 (N_10431,N_9595,N_9808);
or U10432 (N_10432,N_9865,N_9775);
or U10433 (N_10433,N_9543,N_9913);
or U10434 (N_10434,N_9649,N_9650);
xnor U10435 (N_10435,N_9577,N_9506);
xnor U10436 (N_10436,N_9576,N_9652);
nor U10437 (N_10437,N_9718,N_9889);
nor U10438 (N_10438,N_9910,N_9703);
xor U10439 (N_10439,N_9538,N_9637);
nand U10440 (N_10440,N_9794,N_9864);
or U10441 (N_10441,N_9618,N_9803);
nand U10442 (N_10442,N_9973,N_9550);
xor U10443 (N_10443,N_9511,N_9748);
xnor U10444 (N_10444,N_9582,N_9508);
and U10445 (N_10445,N_9958,N_9896);
nand U10446 (N_10446,N_9684,N_9759);
xor U10447 (N_10447,N_9986,N_9876);
or U10448 (N_10448,N_9607,N_9625);
xor U10449 (N_10449,N_9725,N_9703);
or U10450 (N_10450,N_9971,N_9511);
nor U10451 (N_10451,N_9979,N_9677);
xnor U10452 (N_10452,N_9771,N_9992);
or U10453 (N_10453,N_9924,N_9869);
nand U10454 (N_10454,N_9991,N_9759);
nor U10455 (N_10455,N_9675,N_9506);
or U10456 (N_10456,N_9770,N_9938);
nor U10457 (N_10457,N_9567,N_9615);
or U10458 (N_10458,N_9973,N_9575);
nand U10459 (N_10459,N_9861,N_9791);
or U10460 (N_10460,N_9504,N_9519);
xnor U10461 (N_10461,N_9761,N_9719);
xor U10462 (N_10462,N_9705,N_9761);
or U10463 (N_10463,N_9975,N_9942);
nand U10464 (N_10464,N_9981,N_9930);
or U10465 (N_10465,N_9532,N_9802);
xnor U10466 (N_10466,N_9822,N_9806);
and U10467 (N_10467,N_9678,N_9868);
nor U10468 (N_10468,N_9829,N_9609);
and U10469 (N_10469,N_9667,N_9793);
nand U10470 (N_10470,N_9655,N_9901);
xor U10471 (N_10471,N_9529,N_9716);
nor U10472 (N_10472,N_9851,N_9803);
nand U10473 (N_10473,N_9900,N_9952);
or U10474 (N_10474,N_9668,N_9508);
and U10475 (N_10475,N_9742,N_9933);
nor U10476 (N_10476,N_9667,N_9620);
nand U10477 (N_10477,N_9986,N_9660);
nor U10478 (N_10478,N_9583,N_9922);
xor U10479 (N_10479,N_9940,N_9732);
and U10480 (N_10480,N_9958,N_9838);
nor U10481 (N_10481,N_9929,N_9627);
or U10482 (N_10482,N_9750,N_9636);
nand U10483 (N_10483,N_9566,N_9998);
xor U10484 (N_10484,N_9619,N_9761);
nand U10485 (N_10485,N_9697,N_9636);
or U10486 (N_10486,N_9658,N_9964);
or U10487 (N_10487,N_9621,N_9572);
nor U10488 (N_10488,N_9852,N_9502);
and U10489 (N_10489,N_9584,N_9996);
xor U10490 (N_10490,N_9573,N_9713);
xor U10491 (N_10491,N_9822,N_9650);
or U10492 (N_10492,N_9796,N_9758);
nor U10493 (N_10493,N_9833,N_9685);
xnor U10494 (N_10494,N_9773,N_9724);
nor U10495 (N_10495,N_9614,N_9519);
or U10496 (N_10496,N_9565,N_9813);
or U10497 (N_10497,N_9894,N_9806);
nand U10498 (N_10498,N_9892,N_9718);
xnor U10499 (N_10499,N_9603,N_9845);
xnor U10500 (N_10500,N_10226,N_10231);
nor U10501 (N_10501,N_10160,N_10434);
xor U10502 (N_10502,N_10118,N_10284);
xnor U10503 (N_10503,N_10474,N_10204);
nor U10504 (N_10504,N_10283,N_10042);
nor U10505 (N_10505,N_10223,N_10206);
or U10506 (N_10506,N_10190,N_10041);
nand U10507 (N_10507,N_10117,N_10458);
nand U10508 (N_10508,N_10378,N_10103);
or U10509 (N_10509,N_10060,N_10000);
xnor U10510 (N_10510,N_10498,N_10374);
or U10511 (N_10511,N_10282,N_10407);
and U10512 (N_10512,N_10119,N_10074);
nand U10513 (N_10513,N_10279,N_10011);
nor U10514 (N_10514,N_10270,N_10006);
nor U10515 (N_10515,N_10201,N_10216);
nand U10516 (N_10516,N_10063,N_10161);
nor U10517 (N_10517,N_10124,N_10017);
xor U10518 (N_10518,N_10172,N_10392);
and U10519 (N_10519,N_10315,N_10435);
nor U10520 (N_10520,N_10157,N_10427);
nor U10521 (N_10521,N_10256,N_10246);
nand U10522 (N_10522,N_10235,N_10421);
nand U10523 (N_10523,N_10010,N_10258);
xor U10524 (N_10524,N_10189,N_10410);
or U10525 (N_10525,N_10304,N_10228);
nor U10526 (N_10526,N_10243,N_10209);
nor U10527 (N_10527,N_10364,N_10014);
nand U10528 (N_10528,N_10207,N_10142);
and U10529 (N_10529,N_10497,N_10092);
and U10530 (N_10530,N_10131,N_10170);
nand U10531 (N_10531,N_10477,N_10121);
and U10532 (N_10532,N_10397,N_10449);
or U10533 (N_10533,N_10199,N_10369);
and U10534 (N_10534,N_10286,N_10416);
or U10535 (N_10535,N_10049,N_10450);
or U10536 (N_10536,N_10318,N_10081);
xor U10537 (N_10537,N_10330,N_10229);
nand U10538 (N_10538,N_10217,N_10418);
nand U10539 (N_10539,N_10431,N_10068);
nand U10540 (N_10540,N_10316,N_10347);
and U10541 (N_10541,N_10461,N_10048);
nor U10542 (N_10542,N_10070,N_10383);
or U10543 (N_10543,N_10134,N_10287);
and U10544 (N_10544,N_10038,N_10150);
nor U10545 (N_10545,N_10173,N_10003);
nand U10546 (N_10546,N_10472,N_10454);
nand U10547 (N_10547,N_10423,N_10093);
xor U10548 (N_10548,N_10085,N_10455);
or U10549 (N_10549,N_10395,N_10137);
or U10550 (N_10550,N_10184,N_10263);
xor U10551 (N_10551,N_10175,N_10156);
nor U10552 (N_10552,N_10188,N_10419);
nand U10553 (N_10553,N_10381,N_10260);
nand U10554 (N_10554,N_10032,N_10391);
nor U10555 (N_10555,N_10023,N_10112);
or U10556 (N_10556,N_10313,N_10333);
nand U10557 (N_10557,N_10297,N_10192);
and U10558 (N_10558,N_10194,N_10130);
xor U10559 (N_10559,N_10125,N_10197);
xnor U10560 (N_10560,N_10295,N_10225);
and U10561 (N_10561,N_10336,N_10035);
and U10562 (N_10562,N_10087,N_10205);
and U10563 (N_10563,N_10016,N_10101);
nand U10564 (N_10564,N_10185,N_10453);
nor U10565 (N_10565,N_10230,N_10490);
xor U10566 (N_10566,N_10499,N_10005);
nand U10567 (N_10567,N_10020,N_10098);
and U10568 (N_10568,N_10417,N_10191);
and U10569 (N_10569,N_10106,N_10187);
or U10570 (N_10570,N_10213,N_10211);
nor U10571 (N_10571,N_10236,N_10430);
nor U10572 (N_10572,N_10466,N_10470);
nor U10573 (N_10573,N_10399,N_10266);
xor U10574 (N_10574,N_10310,N_10342);
nand U10575 (N_10575,N_10232,N_10350);
xnor U10576 (N_10576,N_10344,N_10055);
xor U10577 (N_10577,N_10238,N_10349);
nor U10578 (N_10578,N_10467,N_10019);
nand U10579 (N_10579,N_10234,N_10433);
xor U10580 (N_10580,N_10355,N_10451);
or U10581 (N_10581,N_10319,N_10129);
or U10582 (N_10582,N_10276,N_10412);
and U10583 (N_10583,N_10366,N_10045);
nand U10584 (N_10584,N_10460,N_10224);
xor U10585 (N_10585,N_10377,N_10024);
nor U10586 (N_10586,N_10296,N_10114);
or U10587 (N_10587,N_10116,N_10271);
nor U10588 (N_10588,N_10328,N_10312);
xnor U10589 (N_10589,N_10179,N_10051);
and U10590 (N_10590,N_10273,N_10075);
nor U10591 (N_10591,N_10385,N_10208);
nand U10592 (N_10592,N_10127,N_10200);
or U10593 (N_10593,N_10182,N_10360);
xnor U10594 (N_10594,N_10067,N_10110);
nor U10595 (N_10595,N_10348,N_10241);
nand U10596 (N_10596,N_10008,N_10305);
xnor U10597 (N_10597,N_10135,N_10329);
nor U10598 (N_10598,N_10442,N_10196);
xor U10599 (N_10599,N_10317,N_10043);
nand U10600 (N_10600,N_10496,N_10428);
nor U10601 (N_10601,N_10069,N_10332);
nor U10602 (N_10602,N_10322,N_10462);
or U10603 (N_10603,N_10298,N_10036);
xnor U10604 (N_10604,N_10480,N_10218);
nor U10605 (N_10605,N_10289,N_10169);
xor U10606 (N_10606,N_10227,N_10440);
nand U10607 (N_10607,N_10126,N_10058);
xnor U10608 (N_10608,N_10375,N_10326);
and U10609 (N_10609,N_10459,N_10484);
and U10610 (N_10610,N_10468,N_10202);
and U10611 (N_10611,N_10148,N_10111);
and U10612 (N_10612,N_10141,N_10278);
nand U10613 (N_10613,N_10033,N_10327);
and U10614 (N_10614,N_10183,N_10285);
xnor U10615 (N_10615,N_10052,N_10341);
xnor U10616 (N_10616,N_10086,N_10088);
and U10617 (N_10617,N_10351,N_10039);
nor U10618 (N_10618,N_10394,N_10210);
and U10619 (N_10619,N_10425,N_10193);
nand U10620 (N_10620,N_10186,N_10162);
or U10621 (N_10621,N_10483,N_10149);
nor U10622 (N_10622,N_10143,N_10083);
nand U10623 (N_10623,N_10138,N_10082);
nand U10624 (N_10624,N_10105,N_10398);
and U10625 (N_10625,N_10439,N_10424);
xor U10626 (N_10626,N_10252,N_10294);
xnor U10627 (N_10627,N_10307,N_10053);
and U10628 (N_10628,N_10233,N_10221);
and U10629 (N_10629,N_10097,N_10331);
or U10630 (N_10630,N_10065,N_10379);
nor U10631 (N_10631,N_10174,N_10007);
nor U10632 (N_10632,N_10390,N_10476);
nor U10633 (N_10633,N_10489,N_10494);
nor U10634 (N_10634,N_10465,N_10047);
xnor U10635 (N_10635,N_10203,N_10456);
xnor U10636 (N_10636,N_10422,N_10415);
nor U10637 (N_10637,N_10096,N_10432);
xor U10638 (N_10638,N_10314,N_10357);
nor U10639 (N_10639,N_10146,N_10090);
xnor U10640 (N_10640,N_10109,N_10255);
nand U10641 (N_10641,N_10178,N_10250);
nand U10642 (N_10642,N_10359,N_10158);
nand U10643 (N_10643,N_10361,N_10122);
nor U10644 (N_10644,N_10436,N_10219);
or U10645 (N_10645,N_10066,N_10240);
nor U10646 (N_10646,N_10429,N_10237);
and U10647 (N_10647,N_10413,N_10277);
xor U10648 (N_10648,N_10247,N_10139);
or U10649 (N_10649,N_10242,N_10245);
nand U10650 (N_10650,N_10414,N_10325);
and U10651 (N_10651,N_10300,N_10491);
xnor U10652 (N_10652,N_10473,N_10059);
and U10653 (N_10653,N_10064,N_10057);
xor U10654 (N_10654,N_10373,N_10457);
and U10655 (N_10655,N_10072,N_10015);
nor U10656 (N_10656,N_10324,N_10486);
or U10657 (N_10657,N_10303,N_10257);
or U10658 (N_10658,N_10107,N_10387);
xor U10659 (N_10659,N_10406,N_10249);
or U10660 (N_10660,N_10198,N_10363);
and U10661 (N_10661,N_10140,N_10168);
or U10662 (N_10662,N_10040,N_10031);
and U10663 (N_10663,N_10444,N_10401);
nand U10664 (N_10664,N_10448,N_10446);
and U10665 (N_10665,N_10478,N_10251);
or U10666 (N_10666,N_10411,N_10254);
and U10667 (N_10667,N_10370,N_10469);
or U10668 (N_10668,N_10013,N_10420);
or U10669 (N_10669,N_10408,N_10153);
and U10670 (N_10670,N_10180,N_10291);
xnor U10671 (N_10671,N_10272,N_10362);
and U10672 (N_10672,N_10471,N_10274);
xnor U10673 (N_10673,N_10308,N_10147);
or U10674 (N_10674,N_10267,N_10405);
xnor U10675 (N_10675,N_10292,N_10028);
and U10676 (N_10676,N_10076,N_10367);
or U10677 (N_10677,N_10441,N_10113);
xnor U10678 (N_10678,N_10046,N_10262);
or U10679 (N_10679,N_10004,N_10365);
and U10680 (N_10680,N_10386,N_10080);
and U10681 (N_10681,N_10248,N_10022);
nor U10682 (N_10682,N_10393,N_10154);
nor U10683 (N_10683,N_10094,N_10152);
nor U10684 (N_10684,N_10050,N_10288);
or U10685 (N_10685,N_10320,N_10062);
nand U10686 (N_10686,N_10214,N_10293);
or U10687 (N_10687,N_10337,N_10089);
nor U10688 (N_10688,N_10071,N_10136);
nor U10689 (N_10689,N_10115,N_10027);
or U10690 (N_10690,N_10264,N_10222);
or U10691 (N_10691,N_10488,N_10438);
nor U10692 (N_10692,N_10120,N_10353);
or U10693 (N_10693,N_10380,N_10371);
nor U10694 (N_10694,N_10025,N_10078);
nand U10695 (N_10695,N_10382,N_10463);
xnor U10696 (N_10696,N_10492,N_10340);
nand U10697 (N_10697,N_10012,N_10321);
nor U10698 (N_10698,N_10487,N_10475);
or U10699 (N_10699,N_10177,N_10220);
nand U10700 (N_10700,N_10334,N_10306);
nand U10701 (N_10701,N_10482,N_10054);
xnor U10702 (N_10702,N_10163,N_10485);
and U10703 (N_10703,N_10268,N_10084);
or U10704 (N_10704,N_10244,N_10166);
nor U10705 (N_10705,N_10352,N_10396);
xor U10706 (N_10706,N_10159,N_10100);
and U10707 (N_10707,N_10037,N_10493);
xor U10708 (N_10708,N_10171,N_10167);
nor U10709 (N_10709,N_10384,N_10128);
nand U10710 (N_10710,N_10029,N_10343);
nand U10711 (N_10711,N_10102,N_10132);
or U10712 (N_10712,N_10079,N_10002);
nor U10713 (N_10713,N_10338,N_10151);
xnor U10714 (N_10714,N_10402,N_10261);
nor U10715 (N_10715,N_10345,N_10108);
nor U10716 (N_10716,N_10452,N_10215);
and U10717 (N_10717,N_10346,N_10144);
and U10718 (N_10718,N_10044,N_10239);
xnor U10719 (N_10719,N_10356,N_10133);
xnor U10720 (N_10720,N_10404,N_10056);
and U10721 (N_10721,N_10309,N_10176);
xnor U10722 (N_10722,N_10445,N_10253);
xnor U10723 (N_10723,N_10265,N_10358);
and U10724 (N_10724,N_10409,N_10376);
or U10725 (N_10725,N_10368,N_10481);
nand U10726 (N_10726,N_10335,N_10073);
and U10727 (N_10727,N_10299,N_10212);
or U10728 (N_10728,N_10155,N_10034);
nor U10729 (N_10729,N_10030,N_10290);
xor U10730 (N_10730,N_10389,N_10026);
nor U10731 (N_10731,N_10061,N_10447);
nand U10732 (N_10732,N_10301,N_10323);
and U10733 (N_10733,N_10354,N_10021);
xor U10734 (N_10734,N_10280,N_10339);
nor U10735 (N_10735,N_10311,N_10372);
nand U10736 (N_10736,N_10269,N_10165);
or U10737 (N_10737,N_10495,N_10009);
or U10738 (N_10738,N_10195,N_10388);
xor U10739 (N_10739,N_10181,N_10281);
and U10740 (N_10740,N_10091,N_10302);
and U10741 (N_10741,N_10123,N_10275);
nand U10742 (N_10742,N_10095,N_10464);
nor U10743 (N_10743,N_10018,N_10164);
or U10744 (N_10744,N_10001,N_10104);
nor U10745 (N_10745,N_10099,N_10259);
nand U10746 (N_10746,N_10403,N_10437);
xor U10747 (N_10747,N_10479,N_10145);
nand U10748 (N_10748,N_10443,N_10426);
and U10749 (N_10749,N_10077,N_10400);
and U10750 (N_10750,N_10229,N_10195);
nand U10751 (N_10751,N_10086,N_10160);
nor U10752 (N_10752,N_10140,N_10172);
nand U10753 (N_10753,N_10080,N_10417);
xor U10754 (N_10754,N_10031,N_10033);
xnor U10755 (N_10755,N_10307,N_10227);
and U10756 (N_10756,N_10319,N_10451);
and U10757 (N_10757,N_10488,N_10094);
or U10758 (N_10758,N_10258,N_10061);
xor U10759 (N_10759,N_10192,N_10091);
nand U10760 (N_10760,N_10093,N_10043);
xor U10761 (N_10761,N_10286,N_10374);
xor U10762 (N_10762,N_10147,N_10121);
nor U10763 (N_10763,N_10087,N_10237);
or U10764 (N_10764,N_10438,N_10426);
nand U10765 (N_10765,N_10205,N_10171);
and U10766 (N_10766,N_10406,N_10382);
nor U10767 (N_10767,N_10411,N_10443);
and U10768 (N_10768,N_10121,N_10462);
or U10769 (N_10769,N_10155,N_10249);
and U10770 (N_10770,N_10141,N_10232);
or U10771 (N_10771,N_10090,N_10082);
nor U10772 (N_10772,N_10083,N_10313);
xor U10773 (N_10773,N_10349,N_10067);
nand U10774 (N_10774,N_10341,N_10070);
nand U10775 (N_10775,N_10279,N_10446);
nor U10776 (N_10776,N_10377,N_10007);
or U10777 (N_10777,N_10466,N_10407);
and U10778 (N_10778,N_10243,N_10189);
and U10779 (N_10779,N_10483,N_10287);
and U10780 (N_10780,N_10199,N_10097);
xnor U10781 (N_10781,N_10392,N_10468);
or U10782 (N_10782,N_10382,N_10384);
and U10783 (N_10783,N_10254,N_10155);
or U10784 (N_10784,N_10276,N_10485);
xor U10785 (N_10785,N_10182,N_10039);
and U10786 (N_10786,N_10207,N_10032);
nor U10787 (N_10787,N_10338,N_10110);
xnor U10788 (N_10788,N_10200,N_10233);
and U10789 (N_10789,N_10070,N_10406);
nand U10790 (N_10790,N_10254,N_10307);
nand U10791 (N_10791,N_10480,N_10133);
and U10792 (N_10792,N_10246,N_10226);
and U10793 (N_10793,N_10123,N_10142);
nand U10794 (N_10794,N_10460,N_10425);
xnor U10795 (N_10795,N_10179,N_10386);
and U10796 (N_10796,N_10195,N_10126);
nand U10797 (N_10797,N_10270,N_10186);
nand U10798 (N_10798,N_10392,N_10445);
nor U10799 (N_10799,N_10407,N_10365);
nand U10800 (N_10800,N_10209,N_10348);
nand U10801 (N_10801,N_10276,N_10333);
xor U10802 (N_10802,N_10374,N_10394);
nor U10803 (N_10803,N_10390,N_10197);
nor U10804 (N_10804,N_10435,N_10388);
or U10805 (N_10805,N_10120,N_10063);
and U10806 (N_10806,N_10297,N_10106);
and U10807 (N_10807,N_10030,N_10226);
and U10808 (N_10808,N_10416,N_10008);
nor U10809 (N_10809,N_10247,N_10499);
nor U10810 (N_10810,N_10338,N_10345);
nand U10811 (N_10811,N_10116,N_10351);
and U10812 (N_10812,N_10350,N_10020);
nor U10813 (N_10813,N_10338,N_10108);
xor U10814 (N_10814,N_10217,N_10054);
or U10815 (N_10815,N_10247,N_10133);
xor U10816 (N_10816,N_10360,N_10320);
nand U10817 (N_10817,N_10043,N_10028);
and U10818 (N_10818,N_10086,N_10282);
nand U10819 (N_10819,N_10303,N_10205);
or U10820 (N_10820,N_10242,N_10044);
nor U10821 (N_10821,N_10311,N_10174);
nor U10822 (N_10822,N_10447,N_10335);
nor U10823 (N_10823,N_10080,N_10482);
nor U10824 (N_10824,N_10394,N_10142);
xnor U10825 (N_10825,N_10243,N_10363);
nand U10826 (N_10826,N_10333,N_10202);
and U10827 (N_10827,N_10457,N_10153);
nor U10828 (N_10828,N_10078,N_10035);
nor U10829 (N_10829,N_10401,N_10331);
and U10830 (N_10830,N_10219,N_10176);
nand U10831 (N_10831,N_10047,N_10199);
nor U10832 (N_10832,N_10363,N_10492);
or U10833 (N_10833,N_10025,N_10214);
nor U10834 (N_10834,N_10347,N_10007);
or U10835 (N_10835,N_10436,N_10421);
nand U10836 (N_10836,N_10339,N_10342);
xor U10837 (N_10837,N_10227,N_10044);
or U10838 (N_10838,N_10162,N_10461);
or U10839 (N_10839,N_10219,N_10059);
xnor U10840 (N_10840,N_10052,N_10171);
nand U10841 (N_10841,N_10284,N_10337);
and U10842 (N_10842,N_10313,N_10135);
nor U10843 (N_10843,N_10162,N_10160);
and U10844 (N_10844,N_10348,N_10184);
nand U10845 (N_10845,N_10495,N_10240);
xor U10846 (N_10846,N_10206,N_10449);
nor U10847 (N_10847,N_10493,N_10364);
nor U10848 (N_10848,N_10096,N_10000);
and U10849 (N_10849,N_10151,N_10378);
xnor U10850 (N_10850,N_10461,N_10428);
and U10851 (N_10851,N_10464,N_10418);
and U10852 (N_10852,N_10003,N_10396);
xnor U10853 (N_10853,N_10080,N_10075);
xnor U10854 (N_10854,N_10017,N_10320);
xnor U10855 (N_10855,N_10000,N_10304);
and U10856 (N_10856,N_10015,N_10430);
nor U10857 (N_10857,N_10027,N_10119);
and U10858 (N_10858,N_10338,N_10336);
nor U10859 (N_10859,N_10201,N_10285);
and U10860 (N_10860,N_10430,N_10341);
nor U10861 (N_10861,N_10279,N_10100);
xnor U10862 (N_10862,N_10474,N_10254);
or U10863 (N_10863,N_10280,N_10220);
nand U10864 (N_10864,N_10173,N_10185);
and U10865 (N_10865,N_10452,N_10356);
nand U10866 (N_10866,N_10412,N_10117);
xnor U10867 (N_10867,N_10047,N_10207);
or U10868 (N_10868,N_10464,N_10462);
nand U10869 (N_10869,N_10327,N_10151);
xnor U10870 (N_10870,N_10339,N_10086);
nand U10871 (N_10871,N_10110,N_10126);
nor U10872 (N_10872,N_10147,N_10410);
xnor U10873 (N_10873,N_10337,N_10241);
or U10874 (N_10874,N_10466,N_10070);
xor U10875 (N_10875,N_10095,N_10169);
and U10876 (N_10876,N_10332,N_10110);
and U10877 (N_10877,N_10364,N_10210);
nor U10878 (N_10878,N_10124,N_10392);
nand U10879 (N_10879,N_10411,N_10096);
and U10880 (N_10880,N_10451,N_10426);
and U10881 (N_10881,N_10186,N_10055);
nand U10882 (N_10882,N_10425,N_10445);
or U10883 (N_10883,N_10208,N_10350);
or U10884 (N_10884,N_10013,N_10150);
nor U10885 (N_10885,N_10223,N_10317);
and U10886 (N_10886,N_10449,N_10134);
or U10887 (N_10887,N_10062,N_10453);
xor U10888 (N_10888,N_10064,N_10216);
and U10889 (N_10889,N_10419,N_10024);
nor U10890 (N_10890,N_10434,N_10276);
nand U10891 (N_10891,N_10323,N_10413);
or U10892 (N_10892,N_10432,N_10021);
and U10893 (N_10893,N_10345,N_10371);
nor U10894 (N_10894,N_10488,N_10329);
or U10895 (N_10895,N_10135,N_10252);
or U10896 (N_10896,N_10163,N_10155);
and U10897 (N_10897,N_10245,N_10362);
nor U10898 (N_10898,N_10364,N_10430);
and U10899 (N_10899,N_10333,N_10134);
xor U10900 (N_10900,N_10428,N_10213);
xor U10901 (N_10901,N_10157,N_10159);
nand U10902 (N_10902,N_10207,N_10384);
and U10903 (N_10903,N_10454,N_10221);
nor U10904 (N_10904,N_10288,N_10230);
and U10905 (N_10905,N_10485,N_10062);
or U10906 (N_10906,N_10265,N_10108);
nor U10907 (N_10907,N_10063,N_10146);
and U10908 (N_10908,N_10487,N_10119);
nand U10909 (N_10909,N_10349,N_10057);
nor U10910 (N_10910,N_10282,N_10335);
and U10911 (N_10911,N_10074,N_10103);
nand U10912 (N_10912,N_10399,N_10314);
nor U10913 (N_10913,N_10440,N_10222);
or U10914 (N_10914,N_10035,N_10143);
nor U10915 (N_10915,N_10153,N_10171);
and U10916 (N_10916,N_10054,N_10112);
nand U10917 (N_10917,N_10168,N_10400);
nand U10918 (N_10918,N_10366,N_10115);
xor U10919 (N_10919,N_10090,N_10167);
nand U10920 (N_10920,N_10451,N_10125);
xor U10921 (N_10921,N_10196,N_10003);
nor U10922 (N_10922,N_10288,N_10418);
and U10923 (N_10923,N_10258,N_10064);
or U10924 (N_10924,N_10327,N_10138);
nor U10925 (N_10925,N_10422,N_10284);
xor U10926 (N_10926,N_10073,N_10499);
and U10927 (N_10927,N_10002,N_10110);
and U10928 (N_10928,N_10453,N_10260);
and U10929 (N_10929,N_10335,N_10349);
and U10930 (N_10930,N_10242,N_10404);
nor U10931 (N_10931,N_10147,N_10267);
or U10932 (N_10932,N_10322,N_10235);
or U10933 (N_10933,N_10165,N_10255);
and U10934 (N_10934,N_10162,N_10310);
xor U10935 (N_10935,N_10214,N_10154);
and U10936 (N_10936,N_10328,N_10251);
and U10937 (N_10937,N_10385,N_10447);
or U10938 (N_10938,N_10493,N_10028);
nor U10939 (N_10939,N_10093,N_10329);
xor U10940 (N_10940,N_10383,N_10276);
xnor U10941 (N_10941,N_10099,N_10085);
xnor U10942 (N_10942,N_10464,N_10230);
xor U10943 (N_10943,N_10017,N_10401);
xnor U10944 (N_10944,N_10163,N_10136);
xnor U10945 (N_10945,N_10498,N_10160);
and U10946 (N_10946,N_10062,N_10249);
and U10947 (N_10947,N_10302,N_10146);
xor U10948 (N_10948,N_10248,N_10039);
and U10949 (N_10949,N_10455,N_10295);
or U10950 (N_10950,N_10390,N_10469);
or U10951 (N_10951,N_10089,N_10245);
and U10952 (N_10952,N_10273,N_10306);
or U10953 (N_10953,N_10356,N_10488);
nor U10954 (N_10954,N_10131,N_10406);
nand U10955 (N_10955,N_10459,N_10192);
or U10956 (N_10956,N_10441,N_10487);
xnor U10957 (N_10957,N_10454,N_10203);
or U10958 (N_10958,N_10301,N_10103);
and U10959 (N_10959,N_10462,N_10022);
nand U10960 (N_10960,N_10275,N_10460);
nand U10961 (N_10961,N_10432,N_10044);
nand U10962 (N_10962,N_10076,N_10025);
and U10963 (N_10963,N_10271,N_10227);
nor U10964 (N_10964,N_10099,N_10187);
or U10965 (N_10965,N_10134,N_10451);
xor U10966 (N_10966,N_10230,N_10404);
nand U10967 (N_10967,N_10388,N_10053);
nor U10968 (N_10968,N_10192,N_10209);
or U10969 (N_10969,N_10451,N_10496);
and U10970 (N_10970,N_10084,N_10413);
nand U10971 (N_10971,N_10003,N_10387);
nand U10972 (N_10972,N_10179,N_10431);
and U10973 (N_10973,N_10132,N_10166);
and U10974 (N_10974,N_10232,N_10464);
nand U10975 (N_10975,N_10237,N_10297);
and U10976 (N_10976,N_10222,N_10414);
nand U10977 (N_10977,N_10368,N_10076);
or U10978 (N_10978,N_10226,N_10045);
xor U10979 (N_10979,N_10420,N_10186);
xor U10980 (N_10980,N_10231,N_10237);
and U10981 (N_10981,N_10448,N_10132);
xnor U10982 (N_10982,N_10485,N_10493);
xor U10983 (N_10983,N_10151,N_10010);
nor U10984 (N_10984,N_10173,N_10243);
or U10985 (N_10985,N_10488,N_10033);
and U10986 (N_10986,N_10213,N_10201);
xor U10987 (N_10987,N_10166,N_10426);
and U10988 (N_10988,N_10464,N_10455);
and U10989 (N_10989,N_10308,N_10099);
xnor U10990 (N_10990,N_10079,N_10462);
or U10991 (N_10991,N_10449,N_10116);
and U10992 (N_10992,N_10035,N_10113);
nor U10993 (N_10993,N_10394,N_10344);
nor U10994 (N_10994,N_10045,N_10203);
and U10995 (N_10995,N_10391,N_10341);
xor U10996 (N_10996,N_10350,N_10334);
nor U10997 (N_10997,N_10313,N_10365);
nor U10998 (N_10998,N_10352,N_10299);
or U10999 (N_10999,N_10198,N_10183);
and U11000 (N_11000,N_10550,N_10865);
nand U11001 (N_11001,N_10624,N_10759);
and U11002 (N_11002,N_10555,N_10900);
nor U11003 (N_11003,N_10753,N_10642);
xnor U11004 (N_11004,N_10841,N_10594);
nor U11005 (N_11005,N_10811,N_10991);
and U11006 (N_11006,N_10846,N_10765);
and U11007 (N_11007,N_10596,N_10576);
xor U11008 (N_11008,N_10844,N_10728);
nor U11009 (N_11009,N_10791,N_10534);
nand U11010 (N_11010,N_10872,N_10561);
xor U11011 (N_11011,N_10814,N_10907);
nand U11012 (N_11012,N_10780,N_10587);
xor U11013 (N_11013,N_10834,N_10639);
xnor U11014 (N_11014,N_10793,N_10700);
xor U11015 (N_11015,N_10833,N_10884);
nand U11016 (N_11016,N_10953,N_10645);
nor U11017 (N_11017,N_10828,N_10852);
xor U11018 (N_11018,N_10946,N_10966);
nand U11019 (N_11019,N_10813,N_10644);
or U11020 (N_11020,N_10942,N_10837);
nor U11021 (N_11021,N_10971,N_10520);
nand U11022 (N_11022,N_10689,N_10960);
or U11023 (N_11023,N_10980,N_10735);
xor U11024 (N_11024,N_10731,N_10674);
nor U11025 (N_11025,N_10881,N_10693);
nor U11026 (N_11026,N_10636,N_10663);
nand U11027 (N_11027,N_10789,N_10940);
xor U11028 (N_11028,N_10653,N_10826);
nand U11029 (N_11029,N_10818,N_10547);
or U11030 (N_11030,N_10709,N_10599);
and U11031 (N_11031,N_10912,N_10694);
xor U11032 (N_11032,N_10832,N_10947);
or U11033 (N_11033,N_10609,N_10713);
nor U11034 (N_11034,N_10562,N_10514);
or U11035 (N_11035,N_10879,N_10752);
xor U11036 (N_11036,N_10761,N_10661);
nor U11037 (N_11037,N_10896,N_10679);
nand U11038 (N_11038,N_10558,N_10979);
xor U11039 (N_11039,N_10816,N_10533);
nand U11040 (N_11040,N_10899,N_10598);
nand U11041 (N_11041,N_10937,N_10540);
and U11042 (N_11042,N_10666,N_10740);
or U11043 (N_11043,N_10554,N_10741);
nand U11044 (N_11044,N_10917,N_10866);
nor U11045 (N_11045,N_10830,N_10508);
and U11046 (N_11046,N_10821,N_10795);
xor U11047 (N_11047,N_10678,N_10578);
or U11048 (N_11048,N_10726,N_10994);
or U11049 (N_11049,N_10707,N_10608);
nand U11050 (N_11050,N_10929,N_10559);
xnor U11051 (N_11051,N_10870,N_10840);
nand U11052 (N_11052,N_10506,N_10503);
xor U11053 (N_11053,N_10756,N_10986);
xor U11054 (N_11054,N_10683,N_10716);
nand U11055 (N_11055,N_10792,N_10972);
nand U11056 (N_11056,N_10908,N_10664);
and U11057 (N_11057,N_10968,N_10887);
nor U11058 (N_11058,N_10623,N_10571);
nor U11059 (N_11059,N_10861,N_10688);
nand U11060 (N_11060,N_10770,N_10543);
xor U11061 (N_11061,N_10626,N_10775);
xor U11062 (N_11062,N_10781,N_10746);
and U11063 (N_11063,N_10779,N_10806);
and U11064 (N_11064,N_10748,N_10737);
xor U11065 (N_11065,N_10502,N_10631);
and U11066 (N_11066,N_10904,N_10668);
nand U11067 (N_11067,N_10563,N_10815);
nor U11068 (N_11068,N_10725,N_10703);
or U11069 (N_11069,N_10911,N_10685);
nand U11070 (N_11070,N_10662,N_10938);
nor U11071 (N_11071,N_10771,N_10876);
nor U11072 (N_11072,N_10714,N_10595);
and U11073 (N_11073,N_10982,N_10794);
or U11074 (N_11074,N_10922,N_10560);
or U11075 (N_11075,N_10999,N_10641);
xor U11076 (N_11076,N_10500,N_10601);
nand U11077 (N_11077,N_10807,N_10751);
and U11078 (N_11078,N_10646,N_10656);
or U11079 (N_11079,N_10600,N_10909);
nor U11080 (N_11080,N_10548,N_10566);
xor U11081 (N_11081,N_10916,N_10574);
or U11082 (N_11082,N_10621,N_10579);
and U11083 (N_11083,N_10724,N_10627);
or U11084 (N_11084,N_10886,N_10750);
or U11085 (N_11085,N_10858,N_10640);
nand U11086 (N_11086,N_10605,N_10787);
nor U11087 (N_11087,N_10827,N_10706);
or U11088 (N_11088,N_10754,N_10874);
xnor U11089 (N_11089,N_10913,N_10965);
nand U11090 (N_11090,N_10531,N_10897);
nor U11091 (N_11091,N_10584,N_10905);
xor U11092 (N_11092,N_10831,N_10878);
nand U11093 (N_11093,N_10854,N_10802);
nor U11094 (N_11094,N_10755,N_10658);
or U11095 (N_11095,N_10810,N_10931);
or U11096 (N_11096,N_10962,N_10682);
nor U11097 (N_11097,N_10629,N_10949);
xor U11098 (N_11098,N_10718,N_10567);
nand U11099 (N_11099,N_10860,N_10801);
or U11100 (N_11100,N_10970,N_10546);
xnor U11101 (N_11101,N_10528,N_10501);
nor U11102 (N_11102,N_10914,N_10710);
xor U11103 (N_11103,N_10720,N_10610);
or U11104 (N_11104,N_10691,N_10655);
or U11105 (N_11105,N_10936,N_10894);
nor U11106 (N_11106,N_10635,N_10538);
nor U11107 (N_11107,N_10512,N_10575);
nor U11108 (N_11108,N_10989,N_10696);
nand U11109 (N_11109,N_10783,N_10612);
nor U11110 (N_11110,N_10869,N_10733);
nor U11111 (N_11111,N_10786,N_10808);
nand U11112 (N_11112,N_10829,N_10880);
or U11113 (N_11113,N_10680,N_10855);
or U11114 (N_11114,N_10988,N_10935);
xor U11115 (N_11115,N_10769,N_10684);
and U11116 (N_11116,N_10542,N_10715);
xnor U11117 (N_11117,N_10941,N_10618);
or U11118 (N_11118,N_10997,N_10875);
xnor U11119 (N_11119,N_10788,N_10637);
and U11120 (N_11120,N_10730,N_10934);
nand U11121 (N_11121,N_10647,N_10863);
or U11122 (N_11122,N_10614,N_10686);
nand U11123 (N_11123,N_10836,N_10958);
nand U11124 (N_11124,N_10975,N_10711);
nand U11125 (N_11125,N_10532,N_10749);
and U11126 (N_11126,N_10513,N_10985);
or U11127 (N_11127,N_10853,N_10944);
nor U11128 (N_11128,N_10604,N_10620);
xor U11129 (N_11129,N_10704,N_10950);
nand U11130 (N_11130,N_10504,N_10606);
nor U11131 (N_11131,N_10822,N_10505);
nand U11132 (N_11132,N_10910,N_10964);
nor U11133 (N_11133,N_10898,N_10745);
nor U11134 (N_11134,N_10993,N_10580);
xnor U11135 (N_11135,N_10742,N_10734);
and U11136 (N_11136,N_10565,N_10615);
nand U11137 (N_11137,N_10712,N_10592);
and U11138 (N_11138,N_10885,N_10665);
nor U11139 (N_11139,N_10611,N_10516);
nand U11140 (N_11140,N_10676,N_10868);
nand U11141 (N_11141,N_10586,N_10613);
nor U11142 (N_11142,N_10569,N_10643);
nand U11143 (N_11143,N_10996,N_10521);
nor U11144 (N_11144,N_10955,N_10864);
and U11145 (N_11145,N_10622,N_10892);
nand U11146 (N_11146,N_10654,N_10539);
nand U11147 (N_11147,N_10638,N_10895);
and U11148 (N_11148,N_10681,N_10697);
or U11149 (N_11149,N_10952,N_10782);
and U11150 (N_11150,N_10757,N_10933);
nor U11151 (N_11151,N_10768,N_10590);
and U11152 (N_11152,N_10695,N_10617);
xor U11153 (N_11153,N_10535,N_10650);
or U11154 (N_11154,N_10702,N_10803);
and U11155 (N_11155,N_10785,N_10859);
or U11156 (N_11156,N_10509,N_10925);
nor U11157 (N_11157,N_10848,N_10893);
xor U11158 (N_11158,N_10570,N_10772);
xnor U11159 (N_11159,N_10763,N_10552);
nor U11160 (N_11160,N_10657,N_10890);
and U11161 (N_11161,N_10519,N_10823);
nand U11162 (N_11162,N_10847,N_10800);
and U11163 (N_11163,N_10951,N_10632);
or U11164 (N_11164,N_10867,N_10923);
xnor U11165 (N_11165,N_10723,N_10536);
xnor U11166 (N_11166,N_10969,N_10767);
nor U11167 (N_11167,N_10797,N_10777);
nand U11168 (N_11168,N_10582,N_10729);
xnor U11169 (N_11169,N_10577,N_10820);
and U11170 (N_11170,N_10591,N_10778);
or U11171 (N_11171,N_10659,N_10523);
nor U11172 (N_11172,N_10776,N_10545);
or U11173 (N_11173,N_10717,N_10926);
or U11174 (N_11174,N_10557,N_10541);
nor U11175 (N_11175,N_10549,N_10669);
xor U11176 (N_11176,N_10526,N_10974);
xor U11177 (N_11177,N_10903,N_10995);
nand U11178 (N_11178,N_10630,N_10888);
xnor U11179 (N_11179,N_10524,N_10551);
nand U11180 (N_11180,N_10698,N_10882);
nor U11181 (N_11181,N_10625,N_10928);
nor U11182 (N_11182,N_10992,N_10809);
xnor U11183 (N_11183,N_10959,N_10784);
and U11184 (N_11184,N_10977,N_10510);
nor U11185 (N_11185,N_10798,N_10648);
nor U11186 (N_11186,N_10774,N_10819);
nor U11187 (N_11187,N_10652,N_10984);
nor U11188 (N_11188,N_10553,N_10845);
nand U11189 (N_11189,N_10877,N_10825);
nor U11190 (N_11190,N_10515,N_10727);
nand U11191 (N_11191,N_10633,N_10883);
or U11192 (N_11192,N_10998,N_10517);
and U11193 (N_11193,N_10593,N_10919);
or U11194 (N_11194,N_10701,N_10619);
and U11195 (N_11195,N_10961,N_10842);
nor U11196 (N_11196,N_10747,N_10871);
and U11197 (N_11197,N_10773,N_10744);
nor U11198 (N_11198,N_10760,N_10585);
or U11199 (N_11199,N_10839,N_10602);
nand U11200 (N_11200,N_10804,N_10901);
nand U11201 (N_11201,N_10849,N_10738);
nor U11202 (N_11202,N_10889,N_10963);
or U11203 (N_11203,N_10568,N_10556);
or U11204 (N_11204,N_10722,N_10527);
and U11205 (N_11205,N_10564,N_10954);
xor U11206 (N_11206,N_10597,N_10672);
and U11207 (N_11207,N_10607,N_10537);
nand U11208 (N_11208,N_10719,N_10812);
xor U11209 (N_11209,N_10511,N_10824);
or U11210 (N_11210,N_10507,N_10956);
nand U11211 (N_11211,N_10943,N_10939);
nand U11212 (N_11212,N_10589,N_10790);
xnor U11213 (N_11213,N_10634,N_10687);
and U11214 (N_11214,N_10976,N_10670);
xor U11215 (N_11215,N_10692,N_10529);
nor U11216 (N_11216,N_10805,N_10649);
or U11217 (N_11217,N_10736,N_10708);
nand U11218 (N_11218,N_10851,N_10973);
or U11219 (N_11219,N_10573,N_10583);
nand U11220 (N_11220,N_10906,N_10660);
and U11221 (N_11221,N_10799,N_10675);
xnor U11222 (N_11222,N_10699,N_10677);
xor U11223 (N_11223,N_10856,N_10987);
nand U11224 (N_11224,N_10930,N_10690);
nor U11225 (N_11225,N_10628,N_10732);
nor U11226 (N_11226,N_10902,N_10518);
or U11227 (N_11227,N_10603,N_10957);
or U11228 (N_11228,N_10983,N_10673);
nor U11229 (N_11229,N_10764,N_10932);
nand U11230 (N_11230,N_10530,N_10857);
nand U11231 (N_11231,N_10838,N_10981);
nand U11232 (N_11232,N_10945,N_10921);
xnor U11233 (N_11233,N_10616,N_10525);
xor U11234 (N_11234,N_10651,N_10924);
nor U11235 (N_11235,N_10967,N_10850);
xor U11236 (N_11236,N_10705,N_10835);
nor U11237 (N_11237,N_10873,N_10758);
nand U11238 (N_11238,N_10948,N_10843);
or U11239 (N_11239,N_10739,N_10743);
and U11240 (N_11240,N_10920,N_10766);
nor U11241 (N_11241,N_10762,N_10544);
nor U11242 (N_11242,N_10918,N_10817);
nand U11243 (N_11243,N_10588,N_10978);
xnor U11244 (N_11244,N_10927,N_10522);
nor U11245 (N_11245,N_10667,N_10796);
nand U11246 (N_11246,N_10721,N_10915);
nand U11247 (N_11247,N_10891,N_10671);
nor U11248 (N_11248,N_10572,N_10990);
nand U11249 (N_11249,N_10862,N_10581);
or U11250 (N_11250,N_10675,N_10828);
xor U11251 (N_11251,N_10859,N_10645);
or U11252 (N_11252,N_10732,N_10829);
or U11253 (N_11253,N_10703,N_10802);
nand U11254 (N_11254,N_10740,N_10762);
nand U11255 (N_11255,N_10753,N_10879);
or U11256 (N_11256,N_10813,N_10663);
and U11257 (N_11257,N_10705,N_10771);
or U11258 (N_11258,N_10657,N_10686);
and U11259 (N_11259,N_10504,N_10684);
nand U11260 (N_11260,N_10721,N_10922);
or U11261 (N_11261,N_10707,N_10635);
xnor U11262 (N_11262,N_10561,N_10878);
nand U11263 (N_11263,N_10637,N_10882);
nor U11264 (N_11264,N_10792,N_10854);
nor U11265 (N_11265,N_10521,N_10509);
nand U11266 (N_11266,N_10709,N_10552);
nand U11267 (N_11267,N_10623,N_10500);
xnor U11268 (N_11268,N_10689,N_10664);
nand U11269 (N_11269,N_10674,N_10728);
nand U11270 (N_11270,N_10655,N_10806);
nand U11271 (N_11271,N_10546,N_10820);
or U11272 (N_11272,N_10543,N_10571);
nor U11273 (N_11273,N_10820,N_10579);
and U11274 (N_11274,N_10643,N_10988);
or U11275 (N_11275,N_10777,N_10505);
or U11276 (N_11276,N_10514,N_10753);
xor U11277 (N_11277,N_10839,N_10899);
and U11278 (N_11278,N_10961,N_10743);
xor U11279 (N_11279,N_10815,N_10584);
nand U11280 (N_11280,N_10548,N_10923);
or U11281 (N_11281,N_10988,N_10978);
or U11282 (N_11282,N_10915,N_10876);
xnor U11283 (N_11283,N_10635,N_10927);
and U11284 (N_11284,N_10588,N_10645);
and U11285 (N_11285,N_10964,N_10933);
nand U11286 (N_11286,N_10540,N_10845);
or U11287 (N_11287,N_10755,N_10889);
nand U11288 (N_11288,N_10734,N_10645);
or U11289 (N_11289,N_10515,N_10644);
nand U11290 (N_11290,N_10690,N_10676);
or U11291 (N_11291,N_10908,N_10965);
and U11292 (N_11292,N_10503,N_10608);
nand U11293 (N_11293,N_10863,N_10979);
xnor U11294 (N_11294,N_10962,N_10885);
or U11295 (N_11295,N_10500,N_10824);
nand U11296 (N_11296,N_10910,N_10545);
and U11297 (N_11297,N_10915,N_10894);
nor U11298 (N_11298,N_10575,N_10664);
nor U11299 (N_11299,N_10846,N_10568);
xnor U11300 (N_11300,N_10562,N_10830);
and U11301 (N_11301,N_10593,N_10957);
nand U11302 (N_11302,N_10589,N_10617);
nor U11303 (N_11303,N_10782,N_10675);
nand U11304 (N_11304,N_10876,N_10530);
nor U11305 (N_11305,N_10635,N_10598);
nor U11306 (N_11306,N_10682,N_10708);
nor U11307 (N_11307,N_10884,N_10613);
or U11308 (N_11308,N_10877,N_10880);
nor U11309 (N_11309,N_10794,N_10771);
nor U11310 (N_11310,N_10909,N_10739);
nor U11311 (N_11311,N_10519,N_10708);
and U11312 (N_11312,N_10673,N_10749);
nor U11313 (N_11313,N_10798,N_10765);
nor U11314 (N_11314,N_10812,N_10656);
and U11315 (N_11315,N_10958,N_10639);
nor U11316 (N_11316,N_10606,N_10736);
or U11317 (N_11317,N_10582,N_10930);
xnor U11318 (N_11318,N_10886,N_10877);
and U11319 (N_11319,N_10605,N_10528);
or U11320 (N_11320,N_10635,N_10671);
nor U11321 (N_11321,N_10712,N_10882);
nand U11322 (N_11322,N_10779,N_10535);
nor U11323 (N_11323,N_10648,N_10950);
or U11324 (N_11324,N_10631,N_10962);
xor U11325 (N_11325,N_10733,N_10522);
or U11326 (N_11326,N_10801,N_10624);
nor U11327 (N_11327,N_10961,N_10716);
nor U11328 (N_11328,N_10709,N_10572);
nor U11329 (N_11329,N_10880,N_10870);
and U11330 (N_11330,N_10867,N_10697);
or U11331 (N_11331,N_10534,N_10514);
xnor U11332 (N_11332,N_10942,N_10672);
xor U11333 (N_11333,N_10776,N_10675);
or U11334 (N_11334,N_10641,N_10802);
nor U11335 (N_11335,N_10703,N_10931);
nand U11336 (N_11336,N_10592,N_10519);
nand U11337 (N_11337,N_10719,N_10800);
xnor U11338 (N_11338,N_10985,N_10781);
nand U11339 (N_11339,N_10926,N_10653);
nand U11340 (N_11340,N_10759,N_10920);
or U11341 (N_11341,N_10808,N_10906);
nand U11342 (N_11342,N_10924,N_10817);
nand U11343 (N_11343,N_10891,N_10720);
nor U11344 (N_11344,N_10657,N_10976);
xnor U11345 (N_11345,N_10820,N_10781);
nor U11346 (N_11346,N_10717,N_10640);
xor U11347 (N_11347,N_10605,N_10877);
nand U11348 (N_11348,N_10840,N_10661);
xor U11349 (N_11349,N_10508,N_10915);
xnor U11350 (N_11350,N_10901,N_10701);
xor U11351 (N_11351,N_10989,N_10631);
nor U11352 (N_11352,N_10576,N_10959);
and U11353 (N_11353,N_10708,N_10689);
nand U11354 (N_11354,N_10611,N_10884);
or U11355 (N_11355,N_10525,N_10878);
nor U11356 (N_11356,N_10792,N_10924);
or U11357 (N_11357,N_10800,N_10977);
and U11358 (N_11358,N_10502,N_10795);
nor U11359 (N_11359,N_10847,N_10816);
and U11360 (N_11360,N_10830,N_10788);
nand U11361 (N_11361,N_10629,N_10970);
xor U11362 (N_11362,N_10599,N_10908);
xnor U11363 (N_11363,N_10892,N_10704);
nand U11364 (N_11364,N_10708,N_10889);
or U11365 (N_11365,N_10640,N_10513);
and U11366 (N_11366,N_10531,N_10902);
or U11367 (N_11367,N_10738,N_10748);
or U11368 (N_11368,N_10695,N_10715);
nor U11369 (N_11369,N_10680,N_10633);
xor U11370 (N_11370,N_10926,N_10639);
or U11371 (N_11371,N_10803,N_10648);
nand U11372 (N_11372,N_10934,N_10985);
nand U11373 (N_11373,N_10682,N_10891);
or U11374 (N_11374,N_10590,N_10739);
nor U11375 (N_11375,N_10788,N_10588);
and U11376 (N_11376,N_10560,N_10524);
xnor U11377 (N_11377,N_10511,N_10509);
and U11378 (N_11378,N_10972,N_10537);
xor U11379 (N_11379,N_10989,N_10521);
xnor U11380 (N_11380,N_10821,N_10995);
and U11381 (N_11381,N_10509,N_10858);
xor U11382 (N_11382,N_10746,N_10972);
and U11383 (N_11383,N_10570,N_10982);
nand U11384 (N_11384,N_10831,N_10655);
and U11385 (N_11385,N_10639,N_10917);
nor U11386 (N_11386,N_10791,N_10995);
xnor U11387 (N_11387,N_10592,N_10747);
and U11388 (N_11388,N_10518,N_10771);
xor U11389 (N_11389,N_10640,N_10952);
nand U11390 (N_11390,N_10852,N_10532);
xor U11391 (N_11391,N_10782,N_10687);
nand U11392 (N_11392,N_10508,N_10693);
nor U11393 (N_11393,N_10702,N_10529);
nand U11394 (N_11394,N_10960,N_10687);
nand U11395 (N_11395,N_10670,N_10679);
xnor U11396 (N_11396,N_10816,N_10780);
nor U11397 (N_11397,N_10798,N_10839);
nor U11398 (N_11398,N_10945,N_10898);
or U11399 (N_11399,N_10505,N_10863);
or U11400 (N_11400,N_10940,N_10888);
xnor U11401 (N_11401,N_10605,N_10738);
and U11402 (N_11402,N_10976,N_10787);
xor U11403 (N_11403,N_10517,N_10940);
and U11404 (N_11404,N_10922,N_10943);
and U11405 (N_11405,N_10502,N_10731);
nand U11406 (N_11406,N_10509,N_10751);
and U11407 (N_11407,N_10613,N_10602);
nand U11408 (N_11408,N_10554,N_10539);
and U11409 (N_11409,N_10592,N_10967);
nor U11410 (N_11410,N_10576,N_10624);
nor U11411 (N_11411,N_10583,N_10927);
xnor U11412 (N_11412,N_10755,N_10890);
nor U11413 (N_11413,N_10818,N_10879);
nand U11414 (N_11414,N_10745,N_10822);
xnor U11415 (N_11415,N_10528,N_10798);
and U11416 (N_11416,N_10918,N_10859);
and U11417 (N_11417,N_10712,N_10650);
or U11418 (N_11418,N_10903,N_10600);
nand U11419 (N_11419,N_10505,N_10957);
xor U11420 (N_11420,N_10806,N_10840);
or U11421 (N_11421,N_10509,N_10594);
and U11422 (N_11422,N_10628,N_10564);
xor U11423 (N_11423,N_10532,N_10970);
and U11424 (N_11424,N_10805,N_10591);
xor U11425 (N_11425,N_10810,N_10797);
nor U11426 (N_11426,N_10552,N_10982);
or U11427 (N_11427,N_10784,N_10702);
nor U11428 (N_11428,N_10518,N_10661);
and U11429 (N_11429,N_10991,N_10964);
xnor U11430 (N_11430,N_10847,N_10762);
nand U11431 (N_11431,N_10500,N_10613);
nor U11432 (N_11432,N_10780,N_10591);
xor U11433 (N_11433,N_10601,N_10623);
nand U11434 (N_11434,N_10907,N_10767);
xor U11435 (N_11435,N_10574,N_10955);
nand U11436 (N_11436,N_10726,N_10907);
nor U11437 (N_11437,N_10531,N_10967);
nor U11438 (N_11438,N_10735,N_10550);
nand U11439 (N_11439,N_10726,N_10649);
nor U11440 (N_11440,N_10777,N_10761);
and U11441 (N_11441,N_10774,N_10931);
nor U11442 (N_11442,N_10504,N_10797);
nor U11443 (N_11443,N_10977,N_10686);
or U11444 (N_11444,N_10832,N_10877);
xnor U11445 (N_11445,N_10602,N_10768);
nand U11446 (N_11446,N_10916,N_10544);
and U11447 (N_11447,N_10578,N_10697);
and U11448 (N_11448,N_10536,N_10591);
nor U11449 (N_11449,N_10636,N_10932);
nor U11450 (N_11450,N_10501,N_10742);
nand U11451 (N_11451,N_10873,N_10701);
or U11452 (N_11452,N_10910,N_10604);
xor U11453 (N_11453,N_10773,N_10887);
nor U11454 (N_11454,N_10586,N_10553);
nand U11455 (N_11455,N_10728,N_10630);
and U11456 (N_11456,N_10628,N_10744);
xnor U11457 (N_11457,N_10917,N_10684);
nor U11458 (N_11458,N_10773,N_10700);
and U11459 (N_11459,N_10756,N_10524);
nor U11460 (N_11460,N_10513,N_10768);
and U11461 (N_11461,N_10893,N_10763);
nor U11462 (N_11462,N_10831,N_10844);
and U11463 (N_11463,N_10706,N_10586);
xnor U11464 (N_11464,N_10725,N_10914);
nand U11465 (N_11465,N_10776,N_10595);
xnor U11466 (N_11466,N_10623,N_10581);
and U11467 (N_11467,N_10546,N_10826);
or U11468 (N_11468,N_10824,N_10751);
xnor U11469 (N_11469,N_10881,N_10922);
xor U11470 (N_11470,N_10696,N_10855);
xnor U11471 (N_11471,N_10510,N_10824);
and U11472 (N_11472,N_10556,N_10833);
xor U11473 (N_11473,N_10853,N_10622);
and U11474 (N_11474,N_10718,N_10912);
xnor U11475 (N_11475,N_10748,N_10909);
nand U11476 (N_11476,N_10940,N_10956);
and U11477 (N_11477,N_10675,N_10808);
and U11478 (N_11478,N_10543,N_10581);
or U11479 (N_11479,N_10905,N_10571);
nor U11480 (N_11480,N_10644,N_10801);
xnor U11481 (N_11481,N_10692,N_10625);
or U11482 (N_11482,N_10989,N_10667);
nand U11483 (N_11483,N_10796,N_10616);
and U11484 (N_11484,N_10790,N_10535);
nand U11485 (N_11485,N_10882,N_10501);
and U11486 (N_11486,N_10557,N_10579);
and U11487 (N_11487,N_10637,N_10706);
or U11488 (N_11488,N_10987,N_10500);
nand U11489 (N_11489,N_10962,N_10774);
or U11490 (N_11490,N_10703,N_10825);
or U11491 (N_11491,N_10520,N_10543);
nor U11492 (N_11492,N_10852,N_10554);
xor U11493 (N_11493,N_10866,N_10635);
nor U11494 (N_11494,N_10571,N_10738);
and U11495 (N_11495,N_10647,N_10539);
and U11496 (N_11496,N_10803,N_10649);
or U11497 (N_11497,N_10955,N_10850);
nor U11498 (N_11498,N_10794,N_10983);
nor U11499 (N_11499,N_10820,N_10720);
xnor U11500 (N_11500,N_11332,N_11484);
nand U11501 (N_11501,N_11005,N_11325);
nor U11502 (N_11502,N_11369,N_11212);
nor U11503 (N_11503,N_11255,N_11219);
nor U11504 (N_11504,N_11376,N_11179);
xor U11505 (N_11505,N_11455,N_11430);
or U11506 (N_11506,N_11440,N_11390);
or U11507 (N_11507,N_11481,N_11000);
nor U11508 (N_11508,N_11446,N_11347);
or U11509 (N_11509,N_11428,N_11343);
xnor U11510 (N_11510,N_11175,N_11061);
nand U11511 (N_11511,N_11068,N_11327);
or U11512 (N_11512,N_11195,N_11261);
or U11513 (N_11513,N_11322,N_11177);
xor U11514 (N_11514,N_11112,N_11458);
nor U11515 (N_11515,N_11391,N_11135);
xnor U11516 (N_11516,N_11030,N_11095);
nor U11517 (N_11517,N_11365,N_11114);
nand U11518 (N_11518,N_11364,N_11190);
xnor U11519 (N_11519,N_11259,N_11292);
nor U11520 (N_11520,N_11013,N_11144);
xor U11521 (N_11521,N_11379,N_11444);
or U11522 (N_11522,N_11375,N_11449);
nor U11523 (N_11523,N_11054,N_11227);
nand U11524 (N_11524,N_11386,N_11394);
and U11525 (N_11525,N_11451,N_11252);
nor U11526 (N_11526,N_11492,N_11439);
xnor U11527 (N_11527,N_11027,N_11208);
and U11528 (N_11528,N_11249,N_11371);
xnor U11529 (N_11529,N_11334,N_11064);
xnor U11530 (N_11530,N_11395,N_11337);
nor U11531 (N_11531,N_11370,N_11240);
xor U11532 (N_11532,N_11459,N_11271);
and U11533 (N_11533,N_11268,N_11281);
nand U11534 (N_11534,N_11265,N_11433);
nor U11535 (N_11535,N_11010,N_11091);
xnor U11536 (N_11536,N_11045,N_11183);
nand U11537 (N_11537,N_11423,N_11304);
nand U11538 (N_11538,N_11210,N_11125);
xnor U11539 (N_11539,N_11388,N_11174);
xor U11540 (N_11540,N_11431,N_11075);
or U11541 (N_11541,N_11079,N_11130);
nand U11542 (N_11542,N_11434,N_11059);
nor U11543 (N_11543,N_11341,N_11497);
and U11544 (N_11544,N_11124,N_11493);
nand U11545 (N_11545,N_11129,N_11184);
xor U11546 (N_11546,N_11299,N_11397);
or U11547 (N_11547,N_11254,N_11169);
xnor U11548 (N_11548,N_11466,N_11310);
xor U11549 (N_11549,N_11321,N_11160);
nor U11550 (N_11550,N_11146,N_11137);
and U11551 (N_11551,N_11153,N_11499);
nor U11552 (N_11552,N_11140,N_11479);
or U11553 (N_11553,N_11089,N_11467);
and U11554 (N_11554,N_11462,N_11486);
and U11555 (N_11555,N_11171,N_11076);
and U11556 (N_11556,N_11131,N_11009);
nor U11557 (N_11557,N_11495,N_11498);
and U11558 (N_11558,N_11173,N_11478);
or U11559 (N_11559,N_11052,N_11436);
or U11560 (N_11560,N_11057,N_11096);
nand U11561 (N_11561,N_11127,N_11288);
nand U11562 (N_11562,N_11239,N_11488);
xnor U11563 (N_11563,N_11474,N_11480);
nor U11564 (N_11564,N_11026,N_11279);
or U11565 (N_11565,N_11245,N_11251);
nand U11566 (N_11566,N_11333,N_11264);
and U11567 (N_11567,N_11329,N_11411);
xnor U11568 (N_11568,N_11046,N_11258);
nand U11569 (N_11569,N_11232,N_11063);
and U11570 (N_11570,N_11263,N_11378);
xor U11571 (N_11571,N_11012,N_11283);
or U11572 (N_11572,N_11018,N_11412);
or U11573 (N_11573,N_11448,N_11351);
or U11574 (N_11574,N_11469,N_11342);
nand U11575 (N_11575,N_11143,N_11401);
nor U11576 (N_11576,N_11218,N_11485);
xor U11577 (N_11577,N_11354,N_11119);
nor U11578 (N_11578,N_11093,N_11402);
nor U11579 (N_11579,N_11470,N_11189);
xnor U11580 (N_11580,N_11036,N_11083);
or U11581 (N_11581,N_11250,N_11122);
nand U11582 (N_11582,N_11217,N_11424);
and U11583 (N_11583,N_11330,N_11353);
nand U11584 (N_11584,N_11286,N_11396);
nor U11585 (N_11585,N_11235,N_11496);
or U11586 (N_11586,N_11032,N_11269);
xor U11587 (N_11587,N_11198,N_11348);
and U11588 (N_11588,N_11142,N_11350);
or U11589 (N_11589,N_11319,N_11120);
nand U11590 (N_11590,N_11367,N_11253);
nand U11591 (N_11591,N_11199,N_11085);
nand U11592 (N_11592,N_11324,N_11138);
and U11593 (N_11593,N_11180,N_11416);
nand U11594 (N_11594,N_11105,N_11004);
or U11595 (N_11595,N_11489,N_11023);
nand U11596 (N_11596,N_11355,N_11475);
xor U11597 (N_11597,N_11233,N_11311);
nor U11598 (N_11598,N_11461,N_11368);
and U11599 (N_11599,N_11077,N_11037);
or U11600 (N_11600,N_11298,N_11117);
xnor U11601 (N_11601,N_11302,N_11092);
xor U11602 (N_11602,N_11072,N_11331);
nor U11603 (N_11603,N_11038,N_11274);
nor U11604 (N_11604,N_11405,N_11228);
or U11605 (N_11605,N_11049,N_11362);
or U11606 (N_11606,N_11011,N_11154);
nor U11607 (N_11607,N_11164,N_11290);
xor U11608 (N_11608,N_11115,N_11192);
or U11609 (N_11609,N_11284,N_11050);
xor U11610 (N_11610,N_11377,N_11187);
or U11611 (N_11611,N_11088,N_11081);
nor U11612 (N_11612,N_11483,N_11150);
or U11613 (N_11613,N_11460,N_11197);
nor U11614 (N_11614,N_11016,N_11415);
nand U11615 (N_11615,N_11024,N_11222);
nor U11616 (N_11616,N_11074,N_11028);
nor U11617 (N_11617,N_11019,N_11248);
and U11618 (N_11618,N_11069,N_11214);
or U11619 (N_11619,N_11270,N_11136);
xor U11620 (N_11620,N_11312,N_11313);
xor U11621 (N_11621,N_11361,N_11307);
or U11622 (N_11622,N_11422,N_11099);
or U11623 (N_11623,N_11058,N_11380);
or U11624 (N_11624,N_11225,N_11297);
or U11625 (N_11625,N_11001,N_11078);
xnor U11626 (N_11626,N_11166,N_11477);
nand U11627 (N_11627,N_11106,N_11360);
and U11628 (N_11628,N_11409,N_11213);
nor U11629 (N_11629,N_11326,N_11314);
or U11630 (N_11630,N_11285,N_11170);
or U11631 (N_11631,N_11418,N_11246);
nor U11632 (N_11632,N_11055,N_11158);
nand U11633 (N_11633,N_11111,N_11168);
nand U11634 (N_11634,N_11244,N_11102);
nand U11635 (N_11635,N_11103,N_11303);
xnor U11636 (N_11636,N_11182,N_11065);
nand U11637 (N_11637,N_11456,N_11029);
or U11638 (N_11638,N_11257,N_11188);
and U11639 (N_11639,N_11108,N_11389);
or U11640 (N_11640,N_11305,N_11100);
xor U11641 (N_11641,N_11134,N_11204);
nor U11642 (N_11642,N_11098,N_11482);
nor U11643 (N_11643,N_11003,N_11031);
nor U11644 (N_11644,N_11382,N_11410);
and U11645 (N_11645,N_11186,N_11359);
and U11646 (N_11646,N_11487,N_11398);
and U11647 (N_11647,N_11300,N_11464);
or U11648 (N_11648,N_11205,N_11420);
and U11649 (N_11649,N_11087,N_11155);
or U11650 (N_11650,N_11006,N_11080);
nor U11651 (N_11651,N_11033,N_11231);
or U11652 (N_11652,N_11280,N_11128);
or U11653 (N_11653,N_11211,N_11071);
xnor U11654 (N_11654,N_11275,N_11308);
nor U11655 (N_11655,N_11453,N_11392);
or U11656 (N_11656,N_11357,N_11471);
and U11657 (N_11657,N_11193,N_11441);
or U11658 (N_11658,N_11419,N_11181);
and U11659 (N_11659,N_11294,N_11387);
or U11660 (N_11660,N_11295,N_11406);
xor U11661 (N_11661,N_11309,N_11172);
nand U11662 (N_11662,N_11425,N_11349);
nor U11663 (N_11663,N_11040,N_11047);
nand U11664 (N_11664,N_11306,N_11034);
xnor U11665 (N_11665,N_11393,N_11163);
and U11666 (N_11666,N_11162,N_11476);
nor U11667 (N_11667,N_11452,N_11443);
or U11668 (N_11668,N_11256,N_11336);
nand U11669 (N_11669,N_11021,N_11346);
nor U11670 (N_11670,N_11133,N_11316);
nor U11671 (N_11671,N_11008,N_11039);
or U11672 (N_11672,N_11490,N_11109);
nand U11673 (N_11673,N_11421,N_11427);
or U11674 (N_11674,N_11082,N_11017);
xor U11675 (N_11675,N_11317,N_11159);
nor U11676 (N_11676,N_11273,N_11472);
nor U11677 (N_11677,N_11053,N_11201);
nor U11678 (N_11678,N_11110,N_11293);
nand U11679 (N_11679,N_11296,N_11118);
xor U11680 (N_11680,N_11442,N_11301);
nor U11681 (N_11681,N_11149,N_11178);
nand U11682 (N_11682,N_11236,N_11056);
and U11683 (N_11683,N_11363,N_11438);
or U11684 (N_11684,N_11282,N_11242);
xnor U11685 (N_11685,N_11215,N_11203);
nor U11686 (N_11686,N_11450,N_11260);
nor U11687 (N_11687,N_11426,N_11191);
nand U11688 (N_11688,N_11126,N_11206);
or U11689 (N_11689,N_11044,N_11196);
or U11690 (N_11690,N_11167,N_11086);
nor U11691 (N_11691,N_11042,N_11408);
or U11692 (N_11692,N_11400,N_11151);
and U11693 (N_11693,N_11247,N_11414);
xnor U11694 (N_11694,N_11352,N_11457);
and U11695 (N_11695,N_11277,N_11226);
and U11696 (N_11696,N_11404,N_11454);
and U11697 (N_11697,N_11339,N_11060);
and U11698 (N_11698,N_11356,N_11022);
xnor U11699 (N_11699,N_11373,N_11289);
and U11700 (N_11700,N_11385,N_11156);
nand U11701 (N_11701,N_11015,N_11344);
and U11702 (N_11702,N_11437,N_11291);
nand U11703 (N_11703,N_11051,N_11220);
nand U11704 (N_11704,N_11468,N_11267);
and U11705 (N_11705,N_11335,N_11116);
and U11706 (N_11706,N_11328,N_11463);
or U11707 (N_11707,N_11223,N_11073);
nand U11708 (N_11708,N_11340,N_11157);
nor U11709 (N_11709,N_11374,N_11224);
or U11710 (N_11710,N_11465,N_11216);
nor U11711 (N_11711,N_11221,N_11320);
nor U11712 (N_11712,N_11200,N_11473);
nor U11713 (N_11713,N_11007,N_11121);
nor U11714 (N_11714,N_11209,N_11381);
nor U11715 (N_11715,N_11366,N_11104);
nand U11716 (N_11716,N_11161,N_11084);
nand U11717 (N_11717,N_11237,N_11262);
nor U11718 (N_11718,N_11383,N_11272);
and U11719 (N_11719,N_11407,N_11432);
xnor U11720 (N_11720,N_11278,N_11241);
and U11721 (N_11721,N_11276,N_11429);
nand U11722 (N_11722,N_11043,N_11358);
or U11723 (N_11723,N_11345,N_11107);
and U11724 (N_11724,N_11147,N_11323);
xor U11725 (N_11725,N_11141,N_11384);
nand U11726 (N_11726,N_11152,N_11041);
nor U11727 (N_11727,N_11266,N_11101);
nand U11728 (N_11728,N_11194,N_11148);
or U11729 (N_11729,N_11176,N_11048);
and U11730 (N_11730,N_11067,N_11287);
or U11731 (N_11731,N_11230,N_11066);
or U11732 (N_11732,N_11185,N_11229);
and U11733 (N_11733,N_11315,N_11002);
and U11734 (N_11734,N_11445,N_11123);
nor U11735 (N_11735,N_11318,N_11234);
xor U11736 (N_11736,N_11145,N_11399);
xor U11737 (N_11737,N_11090,N_11097);
nand U11738 (N_11738,N_11035,N_11447);
and U11739 (N_11739,N_11025,N_11139);
xnor U11740 (N_11740,N_11062,N_11338);
xor U11741 (N_11741,N_11070,N_11491);
nand U11742 (N_11742,N_11417,N_11243);
xnor U11743 (N_11743,N_11165,N_11020);
or U11744 (N_11744,N_11094,N_11132);
nor U11745 (N_11745,N_11207,N_11413);
xor U11746 (N_11746,N_11435,N_11113);
xor U11747 (N_11747,N_11238,N_11202);
nand U11748 (N_11748,N_11494,N_11372);
and U11749 (N_11749,N_11403,N_11014);
nor U11750 (N_11750,N_11111,N_11292);
or U11751 (N_11751,N_11268,N_11038);
or U11752 (N_11752,N_11165,N_11157);
xor U11753 (N_11753,N_11391,N_11409);
and U11754 (N_11754,N_11079,N_11399);
nor U11755 (N_11755,N_11268,N_11048);
nand U11756 (N_11756,N_11465,N_11474);
xnor U11757 (N_11757,N_11116,N_11422);
nor U11758 (N_11758,N_11172,N_11435);
nor U11759 (N_11759,N_11342,N_11014);
xnor U11760 (N_11760,N_11289,N_11460);
and U11761 (N_11761,N_11064,N_11292);
and U11762 (N_11762,N_11478,N_11428);
xnor U11763 (N_11763,N_11105,N_11252);
or U11764 (N_11764,N_11146,N_11002);
and U11765 (N_11765,N_11312,N_11403);
xnor U11766 (N_11766,N_11116,N_11282);
or U11767 (N_11767,N_11196,N_11444);
nand U11768 (N_11768,N_11268,N_11156);
nand U11769 (N_11769,N_11479,N_11093);
nor U11770 (N_11770,N_11422,N_11252);
or U11771 (N_11771,N_11324,N_11392);
xnor U11772 (N_11772,N_11138,N_11191);
nor U11773 (N_11773,N_11112,N_11218);
and U11774 (N_11774,N_11338,N_11378);
and U11775 (N_11775,N_11342,N_11184);
and U11776 (N_11776,N_11088,N_11435);
nand U11777 (N_11777,N_11403,N_11414);
nor U11778 (N_11778,N_11232,N_11102);
and U11779 (N_11779,N_11274,N_11262);
xor U11780 (N_11780,N_11430,N_11458);
nand U11781 (N_11781,N_11499,N_11182);
nor U11782 (N_11782,N_11382,N_11436);
xor U11783 (N_11783,N_11417,N_11098);
nand U11784 (N_11784,N_11124,N_11427);
xnor U11785 (N_11785,N_11088,N_11462);
xor U11786 (N_11786,N_11438,N_11445);
xor U11787 (N_11787,N_11038,N_11292);
nand U11788 (N_11788,N_11285,N_11374);
xnor U11789 (N_11789,N_11483,N_11012);
xnor U11790 (N_11790,N_11011,N_11318);
xnor U11791 (N_11791,N_11049,N_11374);
xor U11792 (N_11792,N_11433,N_11309);
and U11793 (N_11793,N_11363,N_11226);
and U11794 (N_11794,N_11248,N_11392);
xnor U11795 (N_11795,N_11222,N_11231);
nand U11796 (N_11796,N_11414,N_11183);
or U11797 (N_11797,N_11300,N_11433);
or U11798 (N_11798,N_11307,N_11137);
or U11799 (N_11799,N_11095,N_11187);
nor U11800 (N_11800,N_11351,N_11395);
or U11801 (N_11801,N_11361,N_11143);
and U11802 (N_11802,N_11479,N_11429);
nor U11803 (N_11803,N_11459,N_11286);
nand U11804 (N_11804,N_11425,N_11158);
nor U11805 (N_11805,N_11268,N_11206);
nor U11806 (N_11806,N_11279,N_11277);
or U11807 (N_11807,N_11244,N_11466);
nand U11808 (N_11808,N_11017,N_11215);
nand U11809 (N_11809,N_11367,N_11187);
nor U11810 (N_11810,N_11046,N_11455);
nor U11811 (N_11811,N_11382,N_11105);
and U11812 (N_11812,N_11282,N_11347);
xnor U11813 (N_11813,N_11103,N_11176);
nand U11814 (N_11814,N_11414,N_11268);
nor U11815 (N_11815,N_11279,N_11388);
nor U11816 (N_11816,N_11467,N_11412);
nor U11817 (N_11817,N_11099,N_11146);
and U11818 (N_11818,N_11165,N_11391);
and U11819 (N_11819,N_11227,N_11250);
or U11820 (N_11820,N_11280,N_11204);
and U11821 (N_11821,N_11426,N_11258);
and U11822 (N_11822,N_11144,N_11002);
nor U11823 (N_11823,N_11355,N_11399);
xnor U11824 (N_11824,N_11373,N_11384);
nand U11825 (N_11825,N_11433,N_11278);
and U11826 (N_11826,N_11002,N_11317);
and U11827 (N_11827,N_11398,N_11168);
and U11828 (N_11828,N_11243,N_11290);
and U11829 (N_11829,N_11312,N_11212);
or U11830 (N_11830,N_11241,N_11001);
nor U11831 (N_11831,N_11481,N_11351);
nand U11832 (N_11832,N_11241,N_11491);
nand U11833 (N_11833,N_11197,N_11171);
nand U11834 (N_11834,N_11065,N_11334);
and U11835 (N_11835,N_11430,N_11095);
and U11836 (N_11836,N_11373,N_11102);
xor U11837 (N_11837,N_11057,N_11350);
nor U11838 (N_11838,N_11217,N_11292);
xor U11839 (N_11839,N_11417,N_11163);
nor U11840 (N_11840,N_11183,N_11186);
xor U11841 (N_11841,N_11449,N_11377);
and U11842 (N_11842,N_11409,N_11038);
nand U11843 (N_11843,N_11060,N_11075);
nand U11844 (N_11844,N_11359,N_11378);
and U11845 (N_11845,N_11025,N_11090);
xor U11846 (N_11846,N_11305,N_11112);
nand U11847 (N_11847,N_11366,N_11276);
and U11848 (N_11848,N_11313,N_11378);
and U11849 (N_11849,N_11114,N_11425);
xnor U11850 (N_11850,N_11055,N_11415);
nand U11851 (N_11851,N_11374,N_11128);
or U11852 (N_11852,N_11473,N_11489);
or U11853 (N_11853,N_11232,N_11182);
nand U11854 (N_11854,N_11343,N_11141);
or U11855 (N_11855,N_11259,N_11216);
nand U11856 (N_11856,N_11369,N_11246);
nand U11857 (N_11857,N_11246,N_11126);
nor U11858 (N_11858,N_11484,N_11109);
or U11859 (N_11859,N_11318,N_11488);
or U11860 (N_11860,N_11348,N_11420);
or U11861 (N_11861,N_11143,N_11465);
or U11862 (N_11862,N_11250,N_11080);
or U11863 (N_11863,N_11073,N_11379);
nor U11864 (N_11864,N_11158,N_11296);
or U11865 (N_11865,N_11058,N_11231);
and U11866 (N_11866,N_11047,N_11126);
xor U11867 (N_11867,N_11091,N_11435);
nand U11868 (N_11868,N_11250,N_11254);
and U11869 (N_11869,N_11139,N_11053);
and U11870 (N_11870,N_11491,N_11051);
or U11871 (N_11871,N_11305,N_11176);
nand U11872 (N_11872,N_11041,N_11115);
and U11873 (N_11873,N_11395,N_11010);
and U11874 (N_11874,N_11241,N_11444);
nor U11875 (N_11875,N_11131,N_11241);
or U11876 (N_11876,N_11255,N_11234);
nand U11877 (N_11877,N_11408,N_11430);
or U11878 (N_11878,N_11147,N_11453);
and U11879 (N_11879,N_11064,N_11134);
nand U11880 (N_11880,N_11306,N_11185);
and U11881 (N_11881,N_11149,N_11169);
nor U11882 (N_11882,N_11218,N_11037);
and U11883 (N_11883,N_11116,N_11330);
nand U11884 (N_11884,N_11210,N_11306);
nor U11885 (N_11885,N_11366,N_11199);
and U11886 (N_11886,N_11084,N_11460);
nor U11887 (N_11887,N_11219,N_11211);
and U11888 (N_11888,N_11318,N_11224);
xor U11889 (N_11889,N_11041,N_11029);
and U11890 (N_11890,N_11361,N_11138);
nand U11891 (N_11891,N_11350,N_11303);
and U11892 (N_11892,N_11030,N_11494);
xnor U11893 (N_11893,N_11011,N_11281);
and U11894 (N_11894,N_11321,N_11330);
and U11895 (N_11895,N_11310,N_11331);
xor U11896 (N_11896,N_11067,N_11417);
and U11897 (N_11897,N_11123,N_11026);
xor U11898 (N_11898,N_11135,N_11472);
or U11899 (N_11899,N_11382,N_11193);
nor U11900 (N_11900,N_11370,N_11211);
or U11901 (N_11901,N_11384,N_11320);
and U11902 (N_11902,N_11060,N_11317);
xnor U11903 (N_11903,N_11437,N_11232);
and U11904 (N_11904,N_11383,N_11157);
xor U11905 (N_11905,N_11106,N_11221);
nor U11906 (N_11906,N_11280,N_11064);
and U11907 (N_11907,N_11221,N_11375);
nand U11908 (N_11908,N_11041,N_11190);
and U11909 (N_11909,N_11340,N_11167);
or U11910 (N_11910,N_11137,N_11216);
nor U11911 (N_11911,N_11416,N_11421);
nor U11912 (N_11912,N_11453,N_11238);
xor U11913 (N_11913,N_11159,N_11384);
or U11914 (N_11914,N_11354,N_11016);
xor U11915 (N_11915,N_11093,N_11019);
nor U11916 (N_11916,N_11306,N_11013);
nor U11917 (N_11917,N_11193,N_11199);
or U11918 (N_11918,N_11018,N_11251);
and U11919 (N_11919,N_11132,N_11355);
or U11920 (N_11920,N_11474,N_11070);
xor U11921 (N_11921,N_11109,N_11027);
xnor U11922 (N_11922,N_11216,N_11377);
nor U11923 (N_11923,N_11189,N_11097);
or U11924 (N_11924,N_11225,N_11232);
xor U11925 (N_11925,N_11322,N_11040);
and U11926 (N_11926,N_11212,N_11111);
and U11927 (N_11927,N_11153,N_11329);
nand U11928 (N_11928,N_11237,N_11200);
nor U11929 (N_11929,N_11435,N_11454);
nand U11930 (N_11930,N_11119,N_11182);
nand U11931 (N_11931,N_11409,N_11449);
and U11932 (N_11932,N_11101,N_11236);
or U11933 (N_11933,N_11294,N_11445);
nand U11934 (N_11934,N_11094,N_11170);
nor U11935 (N_11935,N_11422,N_11377);
nor U11936 (N_11936,N_11172,N_11426);
and U11937 (N_11937,N_11406,N_11369);
nor U11938 (N_11938,N_11265,N_11372);
or U11939 (N_11939,N_11384,N_11018);
xnor U11940 (N_11940,N_11300,N_11057);
and U11941 (N_11941,N_11297,N_11216);
nor U11942 (N_11942,N_11221,N_11147);
nor U11943 (N_11943,N_11448,N_11469);
nand U11944 (N_11944,N_11182,N_11349);
and U11945 (N_11945,N_11202,N_11059);
or U11946 (N_11946,N_11135,N_11294);
xnor U11947 (N_11947,N_11326,N_11381);
or U11948 (N_11948,N_11179,N_11363);
or U11949 (N_11949,N_11472,N_11163);
xnor U11950 (N_11950,N_11118,N_11364);
or U11951 (N_11951,N_11176,N_11245);
or U11952 (N_11952,N_11467,N_11250);
nor U11953 (N_11953,N_11072,N_11198);
nor U11954 (N_11954,N_11406,N_11012);
and U11955 (N_11955,N_11460,N_11338);
xor U11956 (N_11956,N_11427,N_11407);
or U11957 (N_11957,N_11416,N_11060);
and U11958 (N_11958,N_11279,N_11400);
nand U11959 (N_11959,N_11212,N_11249);
xnor U11960 (N_11960,N_11194,N_11142);
nor U11961 (N_11961,N_11308,N_11204);
nand U11962 (N_11962,N_11371,N_11226);
nand U11963 (N_11963,N_11077,N_11007);
or U11964 (N_11964,N_11204,N_11270);
or U11965 (N_11965,N_11038,N_11304);
nor U11966 (N_11966,N_11386,N_11485);
xnor U11967 (N_11967,N_11330,N_11429);
and U11968 (N_11968,N_11420,N_11158);
nand U11969 (N_11969,N_11278,N_11185);
or U11970 (N_11970,N_11492,N_11407);
or U11971 (N_11971,N_11384,N_11238);
and U11972 (N_11972,N_11353,N_11032);
xnor U11973 (N_11973,N_11190,N_11315);
nor U11974 (N_11974,N_11458,N_11052);
or U11975 (N_11975,N_11004,N_11122);
nor U11976 (N_11976,N_11189,N_11263);
and U11977 (N_11977,N_11421,N_11384);
nor U11978 (N_11978,N_11338,N_11352);
nor U11979 (N_11979,N_11467,N_11238);
nor U11980 (N_11980,N_11362,N_11002);
and U11981 (N_11981,N_11249,N_11071);
xnor U11982 (N_11982,N_11385,N_11180);
nor U11983 (N_11983,N_11075,N_11017);
and U11984 (N_11984,N_11107,N_11401);
or U11985 (N_11985,N_11377,N_11072);
xnor U11986 (N_11986,N_11288,N_11241);
nor U11987 (N_11987,N_11479,N_11179);
and U11988 (N_11988,N_11076,N_11262);
and U11989 (N_11989,N_11412,N_11167);
or U11990 (N_11990,N_11442,N_11289);
nand U11991 (N_11991,N_11241,N_11005);
nor U11992 (N_11992,N_11459,N_11268);
and U11993 (N_11993,N_11001,N_11134);
nand U11994 (N_11994,N_11251,N_11086);
nor U11995 (N_11995,N_11362,N_11178);
nand U11996 (N_11996,N_11417,N_11109);
nor U11997 (N_11997,N_11485,N_11031);
nand U11998 (N_11998,N_11186,N_11033);
nor U11999 (N_11999,N_11082,N_11345);
nand U12000 (N_12000,N_11678,N_11598);
or U12001 (N_12001,N_11961,N_11763);
or U12002 (N_12002,N_11797,N_11707);
nor U12003 (N_12003,N_11889,N_11700);
or U12004 (N_12004,N_11987,N_11990);
xnor U12005 (N_12005,N_11999,N_11551);
and U12006 (N_12006,N_11932,N_11603);
and U12007 (N_12007,N_11582,N_11680);
or U12008 (N_12008,N_11936,N_11625);
and U12009 (N_12009,N_11703,N_11920);
nand U12010 (N_12010,N_11535,N_11697);
or U12011 (N_12011,N_11996,N_11600);
or U12012 (N_12012,N_11871,N_11578);
xnor U12013 (N_12013,N_11839,N_11562);
and U12014 (N_12014,N_11682,N_11812);
or U12015 (N_12015,N_11943,N_11514);
or U12016 (N_12016,N_11685,N_11615);
nor U12017 (N_12017,N_11732,N_11907);
nor U12018 (N_12018,N_11923,N_11553);
xnor U12019 (N_12019,N_11838,N_11569);
and U12020 (N_12020,N_11610,N_11765);
nand U12021 (N_12021,N_11588,N_11762);
nand U12022 (N_12022,N_11970,N_11733);
nand U12023 (N_12023,N_11856,N_11575);
and U12024 (N_12024,N_11712,N_11816);
and U12025 (N_12025,N_11721,N_11817);
nor U12026 (N_12026,N_11946,N_11580);
nor U12027 (N_12027,N_11719,N_11767);
nor U12028 (N_12028,N_11888,N_11847);
xor U12029 (N_12029,N_11823,N_11964);
or U12030 (N_12030,N_11628,N_11583);
and U12031 (N_12031,N_11858,N_11820);
and U12032 (N_12032,N_11892,N_11750);
nor U12033 (N_12033,N_11941,N_11660);
and U12034 (N_12034,N_11821,N_11806);
nand U12035 (N_12035,N_11908,N_11554);
or U12036 (N_12036,N_11813,N_11541);
and U12037 (N_12037,N_11503,N_11691);
and U12038 (N_12038,N_11877,N_11559);
nand U12039 (N_12039,N_11737,N_11925);
or U12040 (N_12040,N_11619,N_11741);
or U12041 (N_12041,N_11656,N_11959);
xor U12042 (N_12042,N_11924,N_11798);
nor U12043 (N_12043,N_11713,N_11543);
and U12044 (N_12044,N_11523,N_11525);
and U12045 (N_12045,N_11881,N_11804);
nor U12046 (N_12046,N_11853,N_11507);
nand U12047 (N_12047,N_11770,N_11533);
nand U12048 (N_12048,N_11571,N_11743);
xor U12049 (N_12049,N_11612,N_11702);
and U12050 (N_12050,N_11926,N_11893);
or U12051 (N_12051,N_11601,N_11793);
and U12052 (N_12052,N_11659,N_11865);
nand U12053 (N_12053,N_11945,N_11686);
nor U12054 (N_12054,N_11909,N_11758);
nand U12055 (N_12055,N_11662,N_11940);
and U12056 (N_12056,N_11657,N_11969);
nand U12057 (N_12057,N_11784,N_11792);
xor U12058 (N_12058,N_11992,N_11833);
xor U12059 (N_12059,N_11783,N_11772);
nand U12060 (N_12060,N_11555,N_11540);
and U12061 (N_12061,N_11661,N_11529);
nand U12062 (N_12062,N_11720,N_11501);
or U12063 (N_12063,N_11903,N_11854);
and U12064 (N_12064,N_11708,N_11550);
and U12065 (N_12065,N_11519,N_11761);
nand U12066 (N_12066,N_11753,N_11664);
and U12067 (N_12067,N_11887,N_11728);
nor U12068 (N_12068,N_11778,N_11746);
and U12069 (N_12069,N_11984,N_11912);
xnor U12070 (N_12070,N_11641,N_11734);
nor U12071 (N_12071,N_11542,N_11973);
or U12072 (N_12072,N_11972,N_11749);
nand U12073 (N_12073,N_11826,N_11511);
or U12074 (N_12074,N_11631,N_11790);
nor U12075 (N_12075,N_11819,N_11614);
or U12076 (N_12076,N_11704,N_11827);
or U12077 (N_12077,N_11736,N_11671);
nor U12078 (N_12078,N_11568,N_11979);
or U12079 (N_12079,N_11930,N_11563);
xnor U12080 (N_12080,N_11739,N_11836);
or U12081 (N_12081,N_11683,N_11870);
and U12082 (N_12082,N_11735,N_11620);
or U12083 (N_12083,N_11531,N_11611);
xnor U12084 (N_12084,N_11729,N_11693);
or U12085 (N_12085,N_11950,N_11808);
nand U12086 (N_12086,N_11803,N_11844);
nand U12087 (N_12087,N_11645,N_11592);
xnor U12088 (N_12088,N_11991,N_11876);
xnor U12089 (N_12089,N_11998,N_11597);
nor U12090 (N_12090,N_11957,N_11521);
nand U12091 (N_12091,N_11584,N_11599);
xor U12092 (N_12092,N_11769,N_11850);
nor U12093 (N_12093,N_11560,N_11883);
or U12094 (N_12094,N_11518,N_11755);
nor U12095 (N_12095,N_11648,N_11787);
xnor U12096 (N_12096,N_11670,N_11629);
and U12097 (N_12097,N_11723,N_11647);
nor U12098 (N_12098,N_11633,N_11825);
or U12099 (N_12099,N_11891,N_11919);
and U12100 (N_12100,N_11849,N_11727);
and U12101 (N_12101,N_11801,N_11902);
nor U12102 (N_12102,N_11897,N_11944);
nor U12103 (N_12103,N_11677,N_11570);
or U12104 (N_12104,N_11818,N_11658);
or U12105 (N_12105,N_11933,N_11526);
and U12106 (N_12106,N_11985,N_11567);
nand U12107 (N_12107,N_11795,N_11617);
xnor U12108 (N_12108,N_11829,N_11627);
or U12109 (N_12109,N_11634,N_11502);
xnor U12110 (N_12110,N_11982,N_11807);
or U12111 (N_12111,N_11914,N_11799);
nand U12112 (N_12112,N_11766,N_11794);
or U12113 (N_12113,N_11744,N_11717);
nand U12114 (N_12114,N_11952,N_11968);
and U12115 (N_12115,N_11824,N_11832);
and U12116 (N_12116,N_11642,N_11556);
xnor U12117 (N_12117,N_11949,N_11710);
nand U12118 (N_12118,N_11725,N_11637);
nand U12119 (N_12119,N_11815,N_11626);
nor U12120 (N_12120,N_11840,N_11831);
xnor U12121 (N_12121,N_11586,N_11978);
and U12122 (N_12122,N_11921,N_11724);
xnor U12123 (N_12123,N_11546,N_11545);
and U12124 (N_12124,N_11557,N_11951);
nor U12125 (N_12125,N_11915,N_11731);
xor U12126 (N_12126,N_11880,N_11948);
and U12127 (N_12127,N_11768,N_11929);
and U12128 (N_12128,N_11864,N_11975);
and U12129 (N_12129,N_11796,N_11852);
nand U12130 (N_12130,N_11669,N_11809);
or U12131 (N_12131,N_11916,N_11938);
nand U12132 (N_12132,N_11869,N_11564);
nand U12133 (N_12133,N_11937,N_11576);
nor U12134 (N_12134,N_11995,N_11913);
or U12135 (N_12135,N_11747,N_11667);
nor U12136 (N_12136,N_11591,N_11956);
or U12137 (N_12137,N_11742,N_11547);
or U12138 (N_12138,N_11757,N_11623);
and U12139 (N_12139,N_11609,N_11911);
or U12140 (N_12140,N_11654,N_11530);
nor U12141 (N_12141,N_11810,N_11834);
nand U12142 (N_12142,N_11608,N_11607);
or U12143 (N_12143,N_11885,N_11756);
or U12144 (N_12144,N_11500,N_11851);
nor U12145 (N_12145,N_11989,N_11552);
and U12146 (N_12146,N_11986,N_11775);
xor U12147 (N_12147,N_11878,N_11706);
nand U12148 (N_12148,N_11745,N_11934);
and U12149 (N_12149,N_11699,N_11997);
and U12150 (N_12150,N_11845,N_11760);
xnor U12151 (N_12151,N_11726,N_11635);
nand U12152 (N_12152,N_11701,N_11574);
and U12153 (N_12153,N_11896,N_11522);
nand U12154 (N_12154,N_11917,N_11638);
or U12155 (N_12155,N_11947,N_11566);
nor U12156 (N_12156,N_11565,N_11788);
or U12157 (N_12157,N_11898,N_11528);
nand U12158 (N_12158,N_11587,N_11841);
and U12159 (N_12159,N_11505,N_11630);
and U12160 (N_12160,N_11536,N_11874);
xor U12161 (N_12161,N_11651,N_11695);
xnor U12162 (N_12162,N_11718,N_11860);
xnor U12163 (N_12163,N_11558,N_11595);
xor U12164 (N_12164,N_11855,N_11859);
and U12165 (N_12165,N_11520,N_11513);
nand U12166 (N_12166,N_11901,N_11527);
nand U12167 (N_12167,N_11974,N_11585);
and U12168 (N_12168,N_11976,N_11684);
and U12169 (N_12169,N_11894,N_11716);
xor U12170 (N_12170,N_11646,N_11605);
nor U12171 (N_12171,N_11879,N_11900);
or U12172 (N_12172,N_11666,N_11581);
or U12173 (N_12173,N_11590,N_11643);
or U12174 (N_12174,N_11604,N_11754);
nor U12175 (N_12175,N_11875,N_11649);
nand U12176 (N_12176,N_11621,N_11977);
or U12177 (N_12177,N_11675,N_11785);
nand U12178 (N_12178,N_11539,N_11506);
nor U12179 (N_12179,N_11764,N_11953);
and U12180 (N_12180,N_11679,N_11942);
nor U12181 (N_12181,N_11512,N_11906);
nand U12182 (N_12182,N_11805,N_11689);
nand U12183 (N_12183,N_11709,N_11759);
nor U12184 (N_12184,N_11960,N_11594);
xnor U12185 (N_12185,N_11613,N_11668);
nand U12186 (N_12186,N_11927,N_11866);
or U12187 (N_12187,N_11549,N_11516);
nor U12188 (N_12188,N_11655,N_11508);
or U12189 (N_12189,N_11884,N_11782);
and U12190 (N_12190,N_11673,N_11781);
and U12191 (N_12191,N_11882,N_11993);
or U12192 (N_12192,N_11994,N_11835);
nand U12193 (N_12193,N_11577,N_11644);
and U12194 (N_12194,N_11857,N_11789);
nor U12195 (N_12195,N_11905,N_11517);
and U12196 (N_12196,N_11939,N_11748);
nor U12197 (N_12197,N_11837,N_11663);
nand U12198 (N_12198,N_11814,N_11624);
xnor U12199 (N_12199,N_11504,N_11830);
and U12200 (N_12200,N_11509,N_11722);
or U12201 (N_12201,N_11714,N_11983);
nand U12202 (N_12202,N_11593,N_11665);
nand U12203 (N_12203,N_11606,N_11848);
nor U12204 (N_12204,N_11918,N_11861);
and U12205 (N_12205,N_11981,N_11715);
nand U12206 (N_12206,N_11910,N_11672);
or U12207 (N_12207,N_11618,N_11524);
nand U12208 (N_12208,N_11776,N_11653);
or U12209 (N_12209,N_11800,N_11904);
and U12210 (N_12210,N_11751,N_11544);
nand U12211 (N_12211,N_11573,N_11740);
or U12212 (N_12212,N_11738,N_11867);
nor U12213 (N_12213,N_11873,N_11676);
or U12214 (N_12214,N_11863,N_11534);
xor U12215 (N_12215,N_11935,N_11872);
or U12216 (N_12216,N_11842,N_11538);
nor U12217 (N_12217,N_11966,N_11636);
and U12218 (N_12218,N_11802,N_11640);
nand U12219 (N_12219,N_11688,N_11537);
nor U12220 (N_12220,N_11773,N_11868);
xnor U12221 (N_12221,N_11922,N_11828);
nor U12222 (N_12222,N_11862,N_11639);
and U12223 (N_12223,N_11572,N_11931);
nor U12224 (N_12224,N_11811,N_11650);
nor U12225 (N_12225,N_11955,N_11692);
nand U12226 (N_12226,N_11786,N_11777);
nand U12227 (N_12227,N_11954,N_11886);
or U12228 (N_12228,N_11843,N_11698);
and U12229 (N_12229,N_11771,N_11971);
and U12230 (N_12230,N_11962,N_11967);
nor U12231 (N_12231,N_11652,N_11681);
nand U12232 (N_12232,N_11616,N_11705);
xnor U12233 (N_12233,N_11690,N_11510);
xnor U12234 (N_12234,N_11890,N_11752);
and U12235 (N_12235,N_11965,N_11711);
xor U12236 (N_12236,N_11589,N_11730);
and U12237 (N_12237,N_11928,N_11687);
or U12238 (N_12238,N_11532,N_11846);
or U12239 (N_12239,N_11515,N_11988);
xnor U12240 (N_12240,N_11779,N_11899);
and U12241 (N_12241,N_11622,N_11780);
and U12242 (N_12242,N_11791,N_11963);
xor U12243 (N_12243,N_11548,N_11774);
and U12244 (N_12244,N_11579,N_11822);
or U12245 (N_12245,N_11602,N_11696);
nor U12246 (N_12246,N_11895,N_11632);
and U12247 (N_12247,N_11958,N_11561);
nand U12248 (N_12248,N_11674,N_11980);
xnor U12249 (N_12249,N_11694,N_11596);
xnor U12250 (N_12250,N_11963,N_11995);
and U12251 (N_12251,N_11924,N_11827);
or U12252 (N_12252,N_11747,N_11964);
or U12253 (N_12253,N_11701,N_11677);
and U12254 (N_12254,N_11819,N_11838);
and U12255 (N_12255,N_11717,N_11814);
nand U12256 (N_12256,N_11508,N_11554);
and U12257 (N_12257,N_11967,N_11711);
nand U12258 (N_12258,N_11803,N_11945);
or U12259 (N_12259,N_11974,N_11877);
nand U12260 (N_12260,N_11567,N_11805);
or U12261 (N_12261,N_11806,N_11538);
nor U12262 (N_12262,N_11843,N_11816);
nor U12263 (N_12263,N_11713,N_11964);
nor U12264 (N_12264,N_11557,N_11614);
nor U12265 (N_12265,N_11818,N_11616);
nor U12266 (N_12266,N_11915,N_11590);
and U12267 (N_12267,N_11709,N_11775);
and U12268 (N_12268,N_11649,N_11908);
xor U12269 (N_12269,N_11760,N_11518);
nand U12270 (N_12270,N_11733,N_11866);
and U12271 (N_12271,N_11643,N_11731);
and U12272 (N_12272,N_11705,N_11946);
nand U12273 (N_12273,N_11507,N_11720);
or U12274 (N_12274,N_11640,N_11636);
xnor U12275 (N_12275,N_11854,N_11945);
or U12276 (N_12276,N_11612,N_11792);
or U12277 (N_12277,N_11582,N_11690);
or U12278 (N_12278,N_11976,N_11549);
or U12279 (N_12279,N_11610,N_11969);
xor U12280 (N_12280,N_11666,N_11909);
or U12281 (N_12281,N_11802,N_11619);
and U12282 (N_12282,N_11522,N_11523);
and U12283 (N_12283,N_11961,N_11879);
nand U12284 (N_12284,N_11824,N_11674);
or U12285 (N_12285,N_11515,N_11953);
nand U12286 (N_12286,N_11550,N_11874);
nand U12287 (N_12287,N_11720,N_11787);
xor U12288 (N_12288,N_11821,N_11959);
nand U12289 (N_12289,N_11681,N_11792);
xnor U12290 (N_12290,N_11535,N_11828);
or U12291 (N_12291,N_11640,N_11511);
and U12292 (N_12292,N_11839,N_11805);
nor U12293 (N_12293,N_11974,N_11825);
nor U12294 (N_12294,N_11734,N_11652);
nand U12295 (N_12295,N_11557,N_11935);
nor U12296 (N_12296,N_11518,N_11594);
nor U12297 (N_12297,N_11989,N_11888);
nand U12298 (N_12298,N_11939,N_11775);
nor U12299 (N_12299,N_11866,N_11643);
or U12300 (N_12300,N_11982,N_11745);
or U12301 (N_12301,N_11806,N_11950);
nand U12302 (N_12302,N_11693,N_11736);
or U12303 (N_12303,N_11835,N_11761);
and U12304 (N_12304,N_11993,N_11573);
nand U12305 (N_12305,N_11801,N_11508);
xor U12306 (N_12306,N_11688,N_11968);
or U12307 (N_12307,N_11629,N_11686);
nor U12308 (N_12308,N_11864,N_11820);
nand U12309 (N_12309,N_11866,N_11783);
and U12310 (N_12310,N_11808,N_11578);
and U12311 (N_12311,N_11729,N_11758);
xnor U12312 (N_12312,N_11766,N_11629);
xor U12313 (N_12313,N_11697,N_11523);
nand U12314 (N_12314,N_11641,N_11504);
nand U12315 (N_12315,N_11846,N_11504);
xnor U12316 (N_12316,N_11797,N_11638);
xor U12317 (N_12317,N_11936,N_11594);
or U12318 (N_12318,N_11558,N_11537);
and U12319 (N_12319,N_11998,N_11866);
xnor U12320 (N_12320,N_11952,N_11766);
or U12321 (N_12321,N_11630,N_11749);
or U12322 (N_12322,N_11514,N_11508);
or U12323 (N_12323,N_11853,N_11855);
nor U12324 (N_12324,N_11635,N_11641);
xor U12325 (N_12325,N_11821,N_11706);
xnor U12326 (N_12326,N_11894,N_11896);
xnor U12327 (N_12327,N_11814,N_11747);
nand U12328 (N_12328,N_11852,N_11691);
or U12329 (N_12329,N_11697,N_11633);
nand U12330 (N_12330,N_11833,N_11577);
nor U12331 (N_12331,N_11960,N_11604);
and U12332 (N_12332,N_11747,N_11857);
nand U12333 (N_12333,N_11569,N_11551);
or U12334 (N_12334,N_11504,N_11532);
nor U12335 (N_12335,N_11617,N_11605);
and U12336 (N_12336,N_11884,N_11524);
xnor U12337 (N_12337,N_11782,N_11524);
and U12338 (N_12338,N_11745,N_11563);
nor U12339 (N_12339,N_11777,N_11700);
nor U12340 (N_12340,N_11678,N_11724);
or U12341 (N_12341,N_11777,N_11837);
and U12342 (N_12342,N_11783,N_11807);
xnor U12343 (N_12343,N_11744,N_11767);
xor U12344 (N_12344,N_11839,N_11738);
nand U12345 (N_12345,N_11920,N_11803);
or U12346 (N_12346,N_11675,N_11733);
nor U12347 (N_12347,N_11856,N_11881);
and U12348 (N_12348,N_11797,N_11798);
or U12349 (N_12349,N_11542,N_11630);
and U12350 (N_12350,N_11538,N_11800);
xor U12351 (N_12351,N_11559,N_11753);
and U12352 (N_12352,N_11581,N_11866);
xor U12353 (N_12353,N_11908,N_11539);
nand U12354 (N_12354,N_11568,N_11835);
and U12355 (N_12355,N_11865,N_11682);
or U12356 (N_12356,N_11538,N_11643);
nor U12357 (N_12357,N_11951,N_11856);
xnor U12358 (N_12358,N_11956,N_11985);
and U12359 (N_12359,N_11932,N_11923);
xor U12360 (N_12360,N_11890,N_11663);
nor U12361 (N_12361,N_11504,N_11507);
xnor U12362 (N_12362,N_11965,N_11769);
nor U12363 (N_12363,N_11700,N_11918);
xor U12364 (N_12364,N_11968,N_11662);
and U12365 (N_12365,N_11784,N_11519);
or U12366 (N_12366,N_11894,N_11889);
nand U12367 (N_12367,N_11737,N_11619);
and U12368 (N_12368,N_11603,N_11966);
xnor U12369 (N_12369,N_11537,N_11595);
xnor U12370 (N_12370,N_11878,N_11863);
xnor U12371 (N_12371,N_11728,N_11798);
nand U12372 (N_12372,N_11970,N_11561);
or U12373 (N_12373,N_11507,N_11907);
xnor U12374 (N_12374,N_11567,N_11891);
nor U12375 (N_12375,N_11826,N_11859);
and U12376 (N_12376,N_11923,N_11751);
nand U12377 (N_12377,N_11705,N_11791);
nor U12378 (N_12378,N_11624,N_11881);
nand U12379 (N_12379,N_11667,N_11673);
nand U12380 (N_12380,N_11904,N_11885);
or U12381 (N_12381,N_11707,N_11853);
xor U12382 (N_12382,N_11849,N_11877);
or U12383 (N_12383,N_11906,N_11893);
and U12384 (N_12384,N_11556,N_11571);
nor U12385 (N_12385,N_11963,N_11733);
nand U12386 (N_12386,N_11666,N_11826);
and U12387 (N_12387,N_11590,N_11917);
nor U12388 (N_12388,N_11615,N_11810);
or U12389 (N_12389,N_11519,N_11999);
and U12390 (N_12390,N_11870,N_11906);
nor U12391 (N_12391,N_11886,N_11618);
nor U12392 (N_12392,N_11908,N_11641);
nor U12393 (N_12393,N_11659,N_11686);
nor U12394 (N_12394,N_11575,N_11526);
or U12395 (N_12395,N_11733,N_11973);
nor U12396 (N_12396,N_11554,N_11729);
xor U12397 (N_12397,N_11582,N_11912);
xnor U12398 (N_12398,N_11631,N_11559);
and U12399 (N_12399,N_11586,N_11832);
xnor U12400 (N_12400,N_11724,N_11792);
nor U12401 (N_12401,N_11552,N_11526);
and U12402 (N_12402,N_11602,N_11640);
or U12403 (N_12403,N_11969,N_11980);
and U12404 (N_12404,N_11638,N_11918);
or U12405 (N_12405,N_11672,N_11929);
nand U12406 (N_12406,N_11603,N_11755);
xnor U12407 (N_12407,N_11729,N_11999);
nand U12408 (N_12408,N_11892,N_11916);
and U12409 (N_12409,N_11738,N_11939);
xor U12410 (N_12410,N_11783,N_11574);
nand U12411 (N_12411,N_11736,N_11786);
or U12412 (N_12412,N_11565,N_11626);
and U12413 (N_12413,N_11728,N_11538);
nand U12414 (N_12414,N_11755,N_11746);
xor U12415 (N_12415,N_11820,N_11504);
or U12416 (N_12416,N_11648,N_11599);
and U12417 (N_12417,N_11530,N_11500);
or U12418 (N_12418,N_11509,N_11862);
xor U12419 (N_12419,N_11888,N_11788);
or U12420 (N_12420,N_11768,N_11856);
nor U12421 (N_12421,N_11636,N_11615);
nor U12422 (N_12422,N_11850,N_11976);
or U12423 (N_12423,N_11946,N_11632);
and U12424 (N_12424,N_11741,N_11767);
nor U12425 (N_12425,N_11984,N_11742);
and U12426 (N_12426,N_11569,N_11801);
nor U12427 (N_12427,N_11776,N_11504);
nor U12428 (N_12428,N_11895,N_11928);
and U12429 (N_12429,N_11940,N_11683);
xor U12430 (N_12430,N_11511,N_11949);
and U12431 (N_12431,N_11620,N_11886);
nand U12432 (N_12432,N_11969,N_11784);
or U12433 (N_12433,N_11626,N_11951);
nand U12434 (N_12434,N_11504,N_11720);
or U12435 (N_12435,N_11547,N_11953);
or U12436 (N_12436,N_11873,N_11733);
and U12437 (N_12437,N_11981,N_11717);
nand U12438 (N_12438,N_11704,N_11513);
and U12439 (N_12439,N_11774,N_11563);
nand U12440 (N_12440,N_11530,N_11971);
and U12441 (N_12441,N_11615,N_11503);
nand U12442 (N_12442,N_11746,N_11762);
nor U12443 (N_12443,N_11526,N_11535);
or U12444 (N_12444,N_11857,N_11757);
nand U12445 (N_12445,N_11609,N_11557);
and U12446 (N_12446,N_11864,N_11676);
or U12447 (N_12447,N_11695,N_11871);
and U12448 (N_12448,N_11691,N_11673);
nor U12449 (N_12449,N_11914,N_11944);
nor U12450 (N_12450,N_11821,N_11809);
nand U12451 (N_12451,N_11509,N_11743);
and U12452 (N_12452,N_11517,N_11815);
or U12453 (N_12453,N_11600,N_11673);
xor U12454 (N_12454,N_11521,N_11574);
and U12455 (N_12455,N_11689,N_11841);
nor U12456 (N_12456,N_11730,N_11727);
xor U12457 (N_12457,N_11808,N_11947);
xor U12458 (N_12458,N_11736,N_11879);
and U12459 (N_12459,N_11603,N_11847);
nand U12460 (N_12460,N_11689,N_11591);
and U12461 (N_12461,N_11731,N_11735);
nand U12462 (N_12462,N_11557,N_11836);
nand U12463 (N_12463,N_11660,N_11904);
nor U12464 (N_12464,N_11553,N_11698);
nor U12465 (N_12465,N_11971,N_11878);
nand U12466 (N_12466,N_11988,N_11922);
nand U12467 (N_12467,N_11973,N_11731);
nor U12468 (N_12468,N_11738,N_11883);
nor U12469 (N_12469,N_11973,N_11662);
xor U12470 (N_12470,N_11770,N_11619);
nand U12471 (N_12471,N_11912,N_11845);
nor U12472 (N_12472,N_11920,N_11998);
and U12473 (N_12473,N_11503,N_11767);
nand U12474 (N_12474,N_11767,N_11670);
or U12475 (N_12475,N_11994,N_11823);
or U12476 (N_12476,N_11938,N_11565);
nor U12477 (N_12477,N_11698,N_11615);
xor U12478 (N_12478,N_11777,N_11793);
or U12479 (N_12479,N_11894,N_11500);
nand U12480 (N_12480,N_11529,N_11930);
or U12481 (N_12481,N_11652,N_11711);
xnor U12482 (N_12482,N_11517,N_11866);
xor U12483 (N_12483,N_11820,N_11765);
nand U12484 (N_12484,N_11585,N_11531);
nand U12485 (N_12485,N_11961,N_11798);
nand U12486 (N_12486,N_11534,N_11541);
xnor U12487 (N_12487,N_11548,N_11780);
nor U12488 (N_12488,N_11537,N_11511);
nor U12489 (N_12489,N_11893,N_11817);
nand U12490 (N_12490,N_11980,N_11960);
nand U12491 (N_12491,N_11745,N_11987);
nor U12492 (N_12492,N_11635,N_11786);
or U12493 (N_12493,N_11778,N_11582);
or U12494 (N_12494,N_11748,N_11666);
or U12495 (N_12495,N_11872,N_11927);
and U12496 (N_12496,N_11733,N_11992);
nand U12497 (N_12497,N_11814,N_11873);
and U12498 (N_12498,N_11802,N_11523);
xnor U12499 (N_12499,N_11769,N_11573);
or U12500 (N_12500,N_12098,N_12458);
and U12501 (N_12501,N_12114,N_12288);
or U12502 (N_12502,N_12083,N_12011);
and U12503 (N_12503,N_12322,N_12303);
nand U12504 (N_12504,N_12053,N_12172);
and U12505 (N_12505,N_12398,N_12418);
nand U12506 (N_12506,N_12313,N_12162);
nand U12507 (N_12507,N_12478,N_12327);
or U12508 (N_12508,N_12422,N_12173);
and U12509 (N_12509,N_12015,N_12268);
or U12510 (N_12510,N_12022,N_12308);
nand U12511 (N_12511,N_12437,N_12430);
nor U12512 (N_12512,N_12254,N_12000);
nor U12513 (N_12513,N_12006,N_12450);
nand U12514 (N_12514,N_12289,N_12052);
or U12515 (N_12515,N_12257,N_12387);
nor U12516 (N_12516,N_12104,N_12129);
xor U12517 (N_12517,N_12379,N_12390);
nand U12518 (N_12518,N_12385,N_12323);
nor U12519 (N_12519,N_12446,N_12448);
xnor U12520 (N_12520,N_12463,N_12138);
nor U12521 (N_12521,N_12306,N_12147);
or U12522 (N_12522,N_12141,N_12126);
nand U12523 (N_12523,N_12210,N_12130);
xnor U12524 (N_12524,N_12324,N_12045);
nor U12525 (N_12525,N_12449,N_12163);
xor U12526 (N_12526,N_12346,N_12034);
and U12527 (N_12527,N_12444,N_12490);
nand U12528 (N_12528,N_12486,N_12166);
nor U12529 (N_12529,N_12188,N_12187);
xnor U12530 (N_12530,N_12435,N_12179);
and U12531 (N_12531,N_12017,N_12095);
xnor U12532 (N_12532,N_12493,N_12117);
xnor U12533 (N_12533,N_12497,N_12315);
or U12534 (N_12534,N_12499,N_12487);
and U12535 (N_12535,N_12230,N_12122);
xor U12536 (N_12536,N_12231,N_12408);
nor U12537 (N_12537,N_12321,N_12229);
nor U12538 (N_12538,N_12338,N_12194);
and U12539 (N_12539,N_12201,N_12206);
nand U12540 (N_12540,N_12027,N_12372);
nand U12541 (N_12541,N_12089,N_12073);
xor U12542 (N_12542,N_12169,N_12029);
nand U12543 (N_12543,N_12247,N_12090);
nor U12544 (N_12544,N_12363,N_12415);
xor U12545 (N_12545,N_12472,N_12165);
xor U12546 (N_12546,N_12036,N_12423);
nor U12547 (N_12547,N_12185,N_12439);
xor U12548 (N_12548,N_12263,N_12170);
or U12549 (N_12549,N_12361,N_12399);
xnor U12550 (N_12550,N_12284,N_12436);
nand U12551 (N_12551,N_12107,N_12051);
and U12552 (N_12552,N_12014,N_12309);
xnor U12553 (N_12553,N_12055,N_12181);
nor U12554 (N_12554,N_12214,N_12208);
xor U12555 (N_12555,N_12211,N_12271);
and U12556 (N_12556,N_12237,N_12146);
and U12557 (N_12557,N_12496,N_12222);
xnor U12558 (N_12558,N_12156,N_12153);
xnor U12559 (N_12559,N_12016,N_12360);
nand U12560 (N_12560,N_12047,N_12252);
and U12561 (N_12561,N_12245,N_12364);
nor U12562 (N_12562,N_12485,N_12186);
nand U12563 (N_12563,N_12110,N_12457);
xor U12564 (N_12564,N_12295,N_12150);
nand U12565 (N_12565,N_12154,N_12330);
or U12566 (N_12566,N_12427,N_12175);
and U12567 (N_12567,N_12224,N_12275);
nor U12568 (N_12568,N_12101,N_12099);
or U12569 (N_12569,N_12196,N_12420);
nand U12570 (N_12570,N_12035,N_12351);
xor U12571 (N_12571,N_12269,N_12386);
and U12572 (N_12572,N_12270,N_12197);
or U12573 (N_12573,N_12125,N_12343);
and U12574 (N_12574,N_12426,N_12023);
and U12575 (N_12575,N_12241,N_12442);
or U12576 (N_12576,N_12026,N_12007);
and U12577 (N_12577,N_12137,N_12223);
xor U12578 (N_12578,N_12039,N_12183);
or U12579 (N_12579,N_12178,N_12447);
xnor U12580 (N_12580,N_12302,N_12464);
nand U12581 (N_12581,N_12108,N_12212);
nor U12582 (N_12582,N_12168,N_12082);
or U12583 (N_12583,N_12260,N_12461);
and U12584 (N_12584,N_12093,N_12180);
nand U12585 (N_12585,N_12282,N_12074);
nand U12586 (N_12586,N_12339,N_12228);
or U12587 (N_12587,N_12374,N_12251);
nand U12588 (N_12588,N_12454,N_12318);
nor U12589 (N_12589,N_12362,N_12355);
and U12590 (N_12590,N_12042,N_12468);
and U12591 (N_12591,N_12305,N_12127);
nor U12592 (N_12592,N_12382,N_12492);
and U12593 (N_12593,N_12060,N_12072);
and U12594 (N_12594,N_12349,N_12294);
nand U12595 (N_12595,N_12280,N_12103);
xnor U12596 (N_12596,N_12193,N_12118);
xnor U12597 (N_12597,N_12249,N_12003);
xor U12598 (N_12598,N_12266,N_12480);
xnor U12599 (N_12599,N_12238,N_12044);
nand U12600 (N_12600,N_12264,N_12253);
nor U12601 (N_12601,N_12031,N_12205);
xor U12602 (N_12602,N_12411,N_12344);
and U12603 (N_12603,N_12373,N_12226);
nor U12604 (N_12604,N_12236,N_12317);
and U12605 (N_12605,N_12258,N_12190);
nor U12606 (N_12606,N_12128,N_12337);
nor U12607 (N_12607,N_12043,N_12477);
nor U12608 (N_12608,N_12100,N_12389);
nor U12609 (N_12609,N_12380,N_12164);
nand U12610 (N_12610,N_12445,N_12354);
nand U12611 (N_12611,N_12394,N_12353);
and U12612 (N_12612,N_12091,N_12397);
or U12613 (N_12613,N_12069,N_12184);
nor U12614 (N_12614,N_12123,N_12061);
nand U12615 (N_12615,N_12476,N_12299);
or U12616 (N_12616,N_12075,N_12005);
nor U12617 (N_12617,N_12151,N_12046);
or U12618 (N_12618,N_12310,N_12417);
or U12619 (N_12619,N_12056,N_12024);
nand U12620 (N_12620,N_12157,N_12097);
or U12621 (N_12621,N_12155,N_12388);
and U12622 (N_12622,N_12200,N_12105);
xor U12623 (N_12623,N_12234,N_12347);
or U12624 (N_12624,N_12037,N_12142);
or U12625 (N_12625,N_12067,N_12272);
and U12626 (N_12626,N_12081,N_12058);
nand U12627 (N_12627,N_12265,N_12498);
xor U12628 (N_12628,N_12124,N_12475);
and U12629 (N_12629,N_12048,N_12032);
xor U12630 (N_12630,N_12356,N_12277);
and U12631 (N_12631,N_12391,N_12336);
or U12632 (N_12632,N_12434,N_12012);
or U12633 (N_12633,N_12202,N_12488);
nand U12634 (N_12634,N_12064,N_12413);
nand U12635 (N_12635,N_12033,N_12287);
or U12636 (N_12636,N_12304,N_12131);
nor U12637 (N_12637,N_12297,N_12329);
xor U12638 (N_12638,N_12376,N_12063);
xnor U12639 (N_12639,N_12471,N_12451);
nand U12640 (N_12640,N_12358,N_12174);
or U12641 (N_12641,N_12334,N_12456);
and U12642 (N_12642,N_12484,N_12213);
xnor U12643 (N_12643,N_12176,N_12407);
or U12644 (N_12644,N_12301,N_12009);
nor U12645 (N_12645,N_12331,N_12352);
or U12646 (N_12646,N_12189,N_12167);
nand U12647 (N_12647,N_12158,N_12481);
nand U12648 (N_12648,N_12215,N_12144);
or U12649 (N_12649,N_12119,N_12041);
and U12650 (N_12650,N_12332,N_12218);
nor U12651 (N_12651,N_12261,N_12291);
and U12652 (N_12652,N_12460,N_12019);
nand U12653 (N_12653,N_12465,N_12049);
or U12654 (N_12654,N_12474,N_12292);
nand U12655 (N_12655,N_12143,N_12283);
nor U12656 (N_12656,N_12357,N_12160);
xor U12657 (N_12657,N_12370,N_12491);
and U12658 (N_12658,N_12298,N_12395);
nor U12659 (N_12659,N_12065,N_12133);
or U12660 (N_12660,N_12320,N_12396);
and U12661 (N_12661,N_12429,N_12112);
xnor U12662 (N_12662,N_12350,N_12025);
nand U12663 (N_12663,N_12433,N_12120);
and U12664 (N_12664,N_12239,N_12495);
and U12665 (N_12665,N_12021,N_12182);
xor U12666 (N_12666,N_12207,N_12038);
nor U12667 (N_12667,N_12384,N_12462);
nor U12668 (N_12668,N_12377,N_12115);
and U12669 (N_12669,N_12013,N_12113);
xor U12670 (N_12670,N_12405,N_12345);
nand U12671 (N_12671,N_12001,N_12087);
nor U12672 (N_12672,N_12084,N_12159);
nor U12673 (N_12673,N_12066,N_12078);
nand U12674 (N_12674,N_12220,N_12217);
or U12675 (N_12675,N_12225,N_12401);
or U12676 (N_12676,N_12102,N_12195);
or U12677 (N_12677,N_12018,N_12191);
nor U12678 (N_12678,N_12094,N_12010);
and U12679 (N_12679,N_12470,N_12262);
or U12680 (N_12680,N_12059,N_12088);
nor U12681 (N_12681,N_12077,N_12421);
or U12682 (N_12682,N_12096,N_12335);
or U12683 (N_12683,N_12371,N_12348);
nor U12684 (N_12684,N_12243,N_12242);
nor U12685 (N_12685,N_12341,N_12489);
xnor U12686 (N_12686,N_12040,N_12004);
and U12687 (N_12687,N_12080,N_12199);
nor U12688 (N_12688,N_12057,N_12145);
nand U12689 (N_12689,N_12256,N_12248);
and U12690 (N_12690,N_12425,N_12375);
or U12691 (N_12691,N_12232,N_12455);
nor U12692 (N_12692,N_12227,N_12203);
nand U12693 (N_12693,N_12216,N_12177);
nor U12694 (N_12694,N_12255,N_12367);
nand U12695 (N_12695,N_12325,N_12319);
and U12696 (N_12696,N_12432,N_12274);
or U12697 (N_12697,N_12136,N_12290);
nor U12698 (N_12698,N_12293,N_12393);
nor U12699 (N_12699,N_12092,N_12244);
and U12700 (N_12700,N_12219,N_12412);
nor U12701 (N_12701,N_12273,N_12392);
or U12702 (N_12702,N_12473,N_12281);
and U12703 (N_12703,N_12076,N_12221);
nor U12704 (N_12704,N_12483,N_12198);
nor U12705 (N_12705,N_12431,N_12479);
nor U12706 (N_12706,N_12149,N_12139);
and U12707 (N_12707,N_12482,N_12328);
or U12708 (N_12708,N_12410,N_12116);
nand U12709 (N_12709,N_12246,N_12459);
nor U12710 (N_12710,N_12312,N_12404);
nor U12711 (N_12711,N_12400,N_12326);
xnor U12712 (N_12712,N_12440,N_12453);
nand U12713 (N_12713,N_12452,N_12494);
nand U12714 (N_12714,N_12286,N_12368);
xor U12715 (N_12715,N_12240,N_12403);
and U12716 (N_12716,N_12068,N_12054);
xor U12717 (N_12717,N_12414,N_12278);
and U12718 (N_12718,N_12030,N_12209);
nor U12719 (N_12719,N_12106,N_12416);
xor U12720 (N_12720,N_12134,N_12071);
nand U12721 (N_12721,N_12028,N_12109);
or U12722 (N_12722,N_12002,N_12152);
xnor U12723 (N_12723,N_12161,N_12235);
xnor U12724 (N_12724,N_12342,N_12311);
xnor U12725 (N_12725,N_12424,N_12340);
nand U12726 (N_12726,N_12419,N_12050);
or U12727 (N_12727,N_12135,N_12469);
nand U12728 (N_12728,N_12365,N_12307);
and U12729 (N_12729,N_12020,N_12148);
nor U12730 (N_12730,N_12008,N_12279);
nor U12731 (N_12731,N_12233,N_12314);
and U12732 (N_12732,N_12111,N_12086);
nand U12733 (N_12733,N_12276,N_12369);
nand U12734 (N_12734,N_12409,N_12316);
and U12735 (N_12735,N_12259,N_12467);
or U12736 (N_12736,N_12466,N_12171);
xnor U12737 (N_12737,N_12085,N_12443);
xnor U12738 (N_12738,N_12062,N_12070);
or U12739 (N_12739,N_12132,N_12250);
and U12740 (N_12740,N_12359,N_12441);
nor U12741 (N_12741,N_12121,N_12300);
xnor U12742 (N_12742,N_12428,N_12285);
or U12743 (N_12743,N_12079,N_12378);
nand U12744 (N_12744,N_12383,N_12406);
nor U12745 (N_12745,N_12381,N_12333);
nand U12746 (N_12746,N_12402,N_12204);
and U12747 (N_12747,N_12192,N_12296);
xor U12748 (N_12748,N_12366,N_12267);
and U12749 (N_12749,N_12438,N_12140);
and U12750 (N_12750,N_12315,N_12283);
nor U12751 (N_12751,N_12128,N_12019);
or U12752 (N_12752,N_12033,N_12285);
nor U12753 (N_12753,N_12455,N_12410);
nand U12754 (N_12754,N_12219,N_12444);
or U12755 (N_12755,N_12041,N_12393);
xor U12756 (N_12756,N_12320,N_12337);
xor U12757 (N_12757,N_12158,N_12478);
or U12758 (N_12758,N_12303,N_12430);
nand U12759 (N_12759,N_12391,N_12059);
or U12760 (N_12760,N_12411,N_12040);
nor U12761 (N_12761,N_12346,N_12039);
xor U12762 (N_12762,N_12219,N_12220);
nor U12763 (N_12763,N_12265,N_12264);
and U12764 (N_12764,N_12223,N_12321);
nor U12765 (N_12765,N_12135,N_12143);
nand U12766 (N_12766,N_12256,N_12067);
xnor U12767 (N_12767,N_12262,N_12339);
nor U12768 (N_12768,N_12248,N_12323);
xnor U12769 (N_12769,N_12038,N_12492);
nand U12770 (N_12770,N_12014,N_12305);
xor U12771 (N_12771,N_12178,N_12438);
or U12772 (N_12772,N_12112,N_12493);
xnor U12773 (N_12773,N_12099,N_12356);
xnor U12774 (N_12774,N_12121,N_12487);
nor U12775 (N_12775,N_12239,N_12202);
and U12776 (N_12776,N_12108,N_12075);
nand U12777 (N_12777,N_12172,N_12089);
or U12778 (N_12778,N_12247,N_12245);
nor U12779 (N_12779,N_12185,N_12265);
nand U12780 (N_12780,N_12132,N_12097);
or U12781 (N_12781,N_12436,N_12208);
nand U12782 (N_12782,N_12441,N_12498);
and U12783 (N_12783,N_12420,N_12000);
nor U12784 (N_12784,N_12045,N_12059);
nand U12785 (N_12785,N_12122,N_12111);
and U12786 (N_12786,N_12367,N_12275);
nor U12787 (N_12787,N_12120,N_12150);
nor U12788 (N_12788,N_12031,N_12145);
nand U12789 (N_12789,N_12092,N_12213);
and U12790 (N_12790,N_12273,N_12209);
and U12791 (N_12791,N_12125,N_12438);
nor U12792 (N_12792,N_12277,N_12428);
xnor U12793 (N_12793,N_12486,N_12308);
or U12794 (N_12794,N_12489,N_12264);
nor U12795 (N_12795,N_12320,N_12118);
nand U12796 (N_12796,N_12236,N_12233);
nand U12797 (N_12797,N_12478,N_12025);
or U12798 (N_12798,N_12039,N_12208);
nor U12799 (N_12799,N_12416,N_12154);
nand U12800 (N_12800,N_12076,N_12292);
and U12801 (N_12801,N_12177,N_12296);
or U12802 (N_12802,N_12254,N_12474);
nand U12803 (N_12803,N_12250,N_12108);
and U12804 (N_12804,N_12433,N_12474);
and U12805 (N_12805,N_12248,N_12159);
nor U12806 (N_12806,N_12138,N_12369);
nand U12807 (N_12807,N_12431,N_12273);
or U12808 (N_12808,N_12428,N_12291);
xnor U12809 (N_12809,N_12112,N_12356);
nor U12810 (N_12810,N_12100,N_12367);
xor U12811 (N_12811,N_12185,N_12299);
xor U12812 (N_12812,N_12039,N_12235);
xor U12813 (N_12813,N_12122,N_12288);
xor U12814 (N_12814,N_12425,N_12073);
nand U12815 (N_12815,N_12204,N_12483);
xnor U12816 (N_12816,N_12049,N_12109);
and U12817 (N_12817,N_12247,N_12451);
and U12818 (N_12818,N_12217,N_12142);
nor U12819 (N_12819,N_12275,N_12234);
or U12820 (N_12820,N_12308,N_12312);
nor U12821 (N_12821,N_12025,N_12060);
xnor U12822 (N_12822,N_12476,N_12380);
or U12823 (N_12823,N_12200,N_12435);
nor U12824 (N_12824,N_12067,N_12455);
nor U12825 (N_12825,N_12092,N_12316);
xnor U12826 (N_12826,N_12093,N_12411);
nor U12827 (N_12827,N_12081,N_12202);
xor U12828 (N_12828,N_12164,N_12363);
or U12829 (N_12829,N_12133,N_12021);
and U12830 (N_12830,N_12260,N_12360);
or U12831 (N_12831,N_12016,N_12165);
or U12832 (N_12832,N_12030,N_12052);
nand U12833 (N_12833,N_12022,N_12252);
nand U12834 (N_12834,N_12127,N_12180);
xnor U12835 (N_12835,N_12122,N_12212);
and U12836 (N_12836,N_12488,N_12472);
nor U12837 (N_12837,N_12147,N_12143);
xor U12838 (N_12838,N_12250,N_12042);
nand U12839 (N_12839,N_12265,N_12497);
nor U12840 (N_12840,N_12177,N_12360);
nor U12841 (N_12841,N_12133,N_12398);
nand U12842 (N_12842,N_12472,N_12494);
or U12843 (N_12843,N_12188,N_12409);
or U12844 (N_12844,N_12141,N_12212);
and U12845 (N_12845,N_12467,N_12291);
or U12846 (N_12846,N_12146,N_12286);
nand U12847 (N_12847,N_12030,N_12081);
xnor U12848 (N_12848,N_12378,N_12085);
nor U12849 (N_12849,N_12379,N_12165);
nand U12850 (N_12850,N_12084,N_12167);
nor U12851 (N_12851,N_12252,N_12473);
nand U12852 (N_12852,N_12019,N_12377);
or U12853 (N_12853,N_12368,N_12166);
nor U12854 (N_12854,N_12126,N_12187);
and U12855 (N_12855,N_12338,N_12252);
and U12856 (N_12856,N_12454,N_12031);
nand U12857 (N_12857,N_12441,N_12330);
and U12858 (N_12858,N_12256,N_12167);
and U12859 (N_12859,N_12237,N_12161);
xor U12860 (N_12860,N_12264,N_12275);
xor U12861 (N_12861,N_12201,N_12354);
or U12862 (N_12862,N_12410,N_12001);
or U12863 (N_12863,N_12001,N_12407);
or U12864 (N_12864,N_12138,N_12337);
nand U12865 (N_12865,N_12136,N_12347);
or U12866 (N_12866,N_12212,N_12078);
and U12867 (N_12867,N_12452,N_12346);
nor U12868 (N_12868,N_12091,N_12177);
or U12869 (N_12869,N_12441,N_12014);
or U12870 (N_12870,N_12033,N_12434);
xnor U12871 (N_12871,N_12090,N_12089);
and U12872 (N_12872,N_12147,N_12172);
xor U12873 (N_12873,N_12470,N_12148);
and U12874 (N_12874,N_12066,N_12457);
and U12875 (N_12875,N_12195,N_12457);
xnor U12876 (N_12876,N_12078,N_12016);
and U12877 (N_12877,N_12045,N_12267);
nor U12878 (N_12878,N_12179,N_12053);
nand U12879 (N_12879,N_12233,N_12388);
nor U12880 (N_12880,N_12073,N_12276);
xor U12881 (N_12881,N_12312,N_12434);
xor U12882 (N_12882,N_12359,N_12448);
and U12883 (N_12883,N_12306,N_12218);
or U12884 (N_12884,N_12072,N_12029);
or U12885 (N_12885,N_12182,N_12020);
or U12886 (N_12886,N_12115,N_12005);
xor U12887 (N_12887,N_12198,N_12389);
nor U12888 (N_12888,N_12363,N_12441);
xnor U12889 (N_12889,N_12022,N_12314);
and U12890 (N_12890,N_12294,N_12461);
xnor U12891 (N_12891,N_12284,N_12233);
and U12892 (N_12892,N_12051,N_12234);
nor U12893 (N_12893,N_12408,N_12388);
and U12894 (N_12894,N_12103,N_12270);
xor U12895 (N_12895,N_12372,N_12397);
nor U12896 (N_12896,N_12309,N_12193);
and U12897 (N_12897,N_12170,N_12105);
and U12898 (N_12898,N_12232,N_12349);
nor U12899 (N_12899,N_12430,N_12061);
and U12900 (N_12900,N_12346,N_12487);
xnor U12901 (N_12901,N_12460,N_12401);
nand U12902 (N_12902,N_12281,N_12062);
nand U12903 (N_12903,N_12301,N_12048);
nand U12904 (N_12904,N_12154,N_12099);
or U12905 (N_12905,N_12177,N_12323);
nor U12906 (N_12906,N_12195,N_12429);
and U12907 (N_12907,N_12294,N_12219);
xor U12908 (N_12908,N_12175,N_12266);
or U12909 (N_12909,N_12459,N_12284);
and U12910 (N_12910,N_12087,N_12012);
nor U12911 (N_12911,N_12393,N_12172);
or U12912 (N_12912,N_12035,N_12196);
xnor U12913 (N_12913,N_12134,N_12206);
and U12914 (N_12914,N_12349,N_12391);
and U12915 (N_12915,N_12446,N_12135);
nor U12916 (N_12916,N_12067,N_12276);
or U12917 (N_12917,N_12435,N_12101);
and U12918 (N_12918,N_12378,N_12331);
nor U12919 (N_12919,N_12407,N_12026);
xor U12920 (N_12920,N_12243,N_12056);
and U12921 (N_12921,N_12457,N_12232);
nor U12922 (N_12922,N_12186,N_12195);
and U12923 (N_12923,N_12328,N_12203);
or U12924 (N_12924,N_12278,N_12466);
nand U12925 (N_12925,N_12484,N_12168);
nor U12926 (N_12926,N_12446,N_12264);
xor U12927 (N_12927,N_12148,N_12414);
nor U12928 (N_12928,N_12363,N_12130);
nor U12929 (N_12929,N_12037,N_12186);
or U12930 (N_12930,N_12319,N_12496);
xnor U12931 (N_12931,N_12060,N_12097);
nand U12932 (N_12932,N_12261,N_12396);
and U12933 (N_12933,N_12353,N_12079);
or U12934 (N_12934,N_12332,N_12258);
or U12935 (N_12935,N_12341,N_12183);
nor U12936 (N_12936,N_12208,N_12223);
xnor U12937 (N_12937,N_12415,N_12407);
xor U12938 (N_12938,N_12173,N_12470);
nor U12939 (N_12939,N_12022,N_12357);
and U12940 (N_12940,N_12374,N_12271);
nand U12941 (N_12941,N_12316,N_12238);
nand U12942 (N_12942,N_12002,N_12174);
and U12943 (N_12943,N_12050,N_12001);
and U12944 (N_12944,N_12082,N_12182);
nand U12945 (N_12945,N_12476,N_12472);
nand U12946 (N_12946,N_12134,N_12253);
or U12947 (N_12947,N_12492,N_12404);
xnor U12948 (N_12948,N_12017,N_12337);
or U12949 (N_12949,N_12426,N_12103);
xnor U12950 (N_12950,N_12288,N_12264);
nand U12951 (N_12951,N_12206,N_12361);
and U12952 (N_12952,N_12280,N_12221);
and U12953 (N_12953,N_12428,N_12217);
nand U12954 (N_12954,N_12077,N_12303);
and U12955 (N_12955,N_12387,N_12464);
nor U12956 (N_12956,N_12064,N_12260);
nand U12957 (N_12957,N_12271,N_12225);
or U12958 (N_12958,N_12101,N_12450);
nor U12959 (N_12959,N_12271,N_12072);
or U12960 (N_12960,N_12478,N_12107);
and U12961 (N_12961,N_12488,N_12172);
or U12962 (N_12962,N_12190,N_12298);
nor U12963 (N_12963,N_12189,N_12498);
or U12964 (N_12964,N_12284,N_12127);
or U12965 (N_12965,N_12044,N_12444);
or U12966 (N_12966,N_12402,N_12397);
nand U12967 (N_12967,N_12042,N_12274);
xnor U12968 (N_12968,N_12221,N_12464);
and U12969 (N_12969,N_12372,N_12380);
and U12970 (N_12970,N_12327,N_12390);
nor U12971 (N_12971,N_12282,N_12053);
or U12972 (N_12972,N_12093,N_12323);
nor U12973 (N_12973,N_12274,N_12183);
nand U12974 (N_12974,N_12270,N_12325);
and U12975 (N_12975,N_12108,N_12028);
nor U12976 (N_12976,N_12448,N_12198);
and U12977 (N_12977,N_12475,N_12266);
xnor U12978 (N_12978,N_12297,N_12499);
or U12979 (N_12979,N_12039,N_12468);
and U12980 (N_12980,N_12223,N_12253);
nor U12981 (N_12981,N_12204,N_12328);
xor U12982 (N_12982,N_12034,N_12079);
xnor U12983 (N_12983,N_12382,N_12145);
xnor U12984 (N_12984,N_12099,N_12129);
or U12985 (N_12985,N_12089,N_12470);
xnor U12986 (N_12986,N_12263,N_12364);
nor U12987 (N_12987,N_12253,N_12305);
nor U12988 (N_12988,N_12437,N_12191);
or U12989 (N_12989,N_12263,N_12151);
xnor U12990 (N_12990,N_12077,N_12334);
or U12991 (N_12991,N_12471,N_12342);
and U12992 (N_12992,N_12183,N_12472);
xor U12993 (N_12993,N_12001,N_12412);
nand U12994 (N_12994,N_12445,N_12411);
and U12995 (N_12995,N_12465,N_12417);
or U12996 (N_12996,N_12184,N_12365);
and U12997 (N_12997,N_12089,N_12058);
nor U12998 (N_12998,N_12336,N_12305);
or U12999 (N_12999,N_12383,N_12272);
xnor U13000 (N_13000,N_12570,N_12571);
or U13001 (N_13001,N_12553,N_12951);
nand U13002 (N_13002,N_12893,N_12639);
nor U13003 (N_13003,N_12766,N_12798);
nor U13004 (N_13004,N_12719,N_12908);
xor U13005 (N_13005,N_12802,N_12751);
xor U13006 (N_13006,N_12747,N_12632);
xor U13007 (N_13007,N_12787,N_12651);
or U13008 (N_13008,N_12997,N_12931);
xor U13009 (N_13009,N_12611,N_12677);
nor U13010 (N_13010,N_12772,N_12656);
and U13011 (N_13011,N_12644,N_12635);
nand U13012 (N_13012,N_12636,N_12525);
and U13013 (N_13013,N_12717,N_12946);
and U13014 (N_13014,N_12838,N_12898);
xnor U13015 (N_13015,N_12740,N_12590);
nor U13016 (N_13016,N_12586,N_12830);
nor U13017 (N_13017,N_12616,N_12837);
or U13018 (N_13018,N_12732,N_12736);
and U13019 (N_13019,N_12863,N_12791);
nand U13020 (N_13020,N_12615,N_12793);
nor U13021 (N_13021,N_12701,N_12536);
xor U13022 (N_13022,N_12652,N_12914);
nor U13023 (N_13023,N_12592,N_12682);
xor U13024 (N_13024,N_12731,N_12851);
nand U13025 (N_13025,N_12771,N_12547);
or U13026 (N_13026,N_12862,N_12780);
and U13027 (N_13027,N_12587,N_12937);
nand U13028 (N_13028,N_12777,N_12819);
and U13029 (N_13029,N_12742,N_12961);
and U13030 (N_13030,N_12530,N_12900);
or U13031 (N_13031,N_12988,N_12704);
and U13032 (N_13032,N_12597,N_12550);
or U13033 (N_13033,N_12510,N_12964);
xor U13034 (N_13034,N_12853,N_12580);
nand U13035 (N_13035,N_12660,N_12657);
and U13036 (N_13036,N_12994,N_12733);
or U13037 (N_13037,N_12750,N_12519);
nor U13038 (N_13038,N_12715,N_12794);
xnor U13039 (N_13039,N_12993,N_12722);
nand U13040 (N_13040,N_12546,N_12641);
and U13041 (N_13041,N_12552,N_12601);
and U13042 (N_13042,N_12516,N_12775);
xor U13043 (N_13043,N_12557,N_12690);
or U13044 (N_13044,N_12642,N_12583);
and U13045 (N_13045,N_12844,N_12696);
nand U13046 (N_13046,N_12818,N_12860);
and U13047 (N_13047,N_12948,N_12610);
and U13048 (N_13048,N_12539,N_12779);
xnor U13049 (N_13049,N_12558,N_12581);
or U13050 (N_13050,N_12943,N_12541);
nor U13051 (N_13051,N_12883,N_12889);
xor U13052 (N_13052,N_12620,N_12739);
nand U13053 (N_13053,N_12672,N_12649);
nand U13054 (N_13054,N_12782,N_12855);
xor U13055 (N_13055,N_12500,N_12512);
and U13056 (N_13056,N_12882,N_12990);
and U13057 (N_13057,N_12626,N_12591);
nand U13058 (N_13058,N_12673,N_12506);
nand U13059 (N_13059,N_12650,N_12892);
nor U13060 (N_13060,N_12671,N_12816);
xnor U13061 (N_13061,N_12926,N_12891);
xnor U13062 (N_13062,N_12599,N_12524);
and U13063 (N_13063,N_12934,N_12606);
or U13064 (N_13064,N_12746,N_12797);
xnor U13065 (N_13065,N_12795,N_12637);
or U13066 (N_13066,N_12752,N_12758);
nand U13067 (N_13067,N_12634,N_12630);
xor U13068 (N_13068,N_12562,N_12669);
nand U13069 (N_13069,N_12666,N_12605);
or U13070 (N_13070,N_12609,N_12854);
and U13071 (N_13071,N_12683,N_12728);
or U13072 (N_13072,N_12848,N_12527);
nand U13073 (N_13073,N_12560,N_12589);
nand U13074 (N_13074,N_12573,N_12809);
and U13075 (N_13075,N_12582,N_12958);
nor U13076 (N_13076,N_12959,N_12691);
or U13077 (N_13077,N_12658,N_12999);
nor U13078 (N_13078,N_12577,N_12845);
or U13079 (N_13079,N_12594,N_12832);
nor U13080 (N_13080,N_12874,N_12738);
nand U13081 (N_13081,N_12852,N_12971);
xnor U13082 (N_13082,N_12505,N_12901);
and U13083 (N_13083,N_12697,N_12761);
nand U13084 (N_13084,N_12680,N_12531);
and U13085 (N_13085,N_12684,N_12607);
nor U13086 (N_13086,N_12785,N_12859);
nand U13087 (N_13087,N_12694,N_12538);
or U13088 (N_13088,N_12842,N_12790);
nor U13089 (N_13089,N_12975,N_12815);
xor U13090 (N_13090,N_12501,N_12783);
nor U13091 (N_13091,N_12803,N_12619);
nand U13092 (N_13092,N_12973,N_12757);
xnor U13093 (N_13093,N_12665,N_12850);
or U13094 (N_13094,N_12814,N_12957);
nor U13095 (N_13095,N_12511,N_12831);
and U13096 (N_13096,N_12817,N_12950);
nand U13097 (N_13097,N_12521,N_12847);
nand U13098 (N_13098,N_12907,N_12712);
xnor U13099 (N_13099,N_12678,N_12828);
and U13100 (N_13100,N_12910,N_12861);
xor U13101 (N_13101,N_12767,N_12593);
and U13102 (N_13102,N_12754,N_12698);
nor U13103 (N_13103,N_12935,N_12781);
and U13104 (N_13104,N_12799,N_12764);
xor U13105 (N_13105,N_12743,N_12878);
nand U13106 (N_13106,N_12936,N_12915);
and U13107 (N_13107,N_12695,N_12588);
or U13108 (N_13108,N_12895,N_12595);
nor U13109 (N_13109,N_12822,N_12612);
and U13110 (N_13110,N_12839,N_12692);
and U13111 (N_13111,N_12904,N_12890);
and U13112 (N_13112,N_12744,N_12759);
nor U13113 (N_13113,N_12789,N_12718);
xor U13114 (N_13114,N_12614,N_12663);
xnor U13115 (N_13115,N_12730,N_12982);
nand U13116 (N_13116,N_12792,N_12617);
and U13117 (N_13117,N_12768,N_12956);
nand U13118 (N_13118,N_12824,N_12543);
nor U13119 (N_13119,N_12629,N_12886);
xnor U13120 (N_13120,N_12667,N_12523);
xnor U13121 (N_13121,N_12535,N_12834);
nor U13122 (N_13122,N_12945,N_12645);
and U13123 (N_13123,N_12654,N_12776);
nand U13124 (N_13124,N_12638,N_12579);
nor U13125 (N_13125,N_12709,N_12821);
and U13126 (N_13126,N_12840,N_12986);
and U13127 (N_13127,N_12627,N_12940);
or U13128 (N_13128,N_12784,N_12796);
nand U13129 (N_13129,N_12801,N_12548);
or U13130 (N_13130,N_12966,N_12917);
xnor U13131 (N_13131,N_12554,N_12544);
xnor U13132 (N_13132,N_12858,N_12676);
and U13133 (N_13133,N_12778,N_12923);
or U13134 (N_13134,N_12760,N_12773);
xor U13135 (N_13135,N_12864,N_12963);
xnor U13136 (N_13136,N_12603,N_12625);
xnor U13137 (N_13137,N_12867,N_12880);
and U13138 (N_13138,N_12515,N_12574);
or U13139 (N_13139,N_12911,N_12706);
and U13140 (N_13140,N_12741,N_12970);
nor U13141 (N_13141,N_12913,N_12974);
nand U13142 (N_13142,N_12938,N_12526);
nor U13143 (N_13143,N_12542,N_12856);
and U13144 (N_13144,N_12668,N_12930);
nor U13145 (N_13145,N_12748,N_12517);
xnor U13146 (N_13146,N_12662,N_12756);
nor U13147 (N_13147,N_12769,N_12502);
or U13148 (N_13148,N_12567,N_12735);
or U13149 (N_13149,N_12920,N_12540);
or U13150 (N_13150,N_12813,N_12976);
nand U13151 (N_13151,N_12804,N_12685);
xor U13152 (N_13152,N_12984,N_12763);
nor U13153 (N_13153,N_12969,N_12623);
nor U13154 (N_13154,N_12723,N_12563);
nor U13155 (N_13155,N_12846,N_12545);
or U13156 (N_13156,N_12962,N_12716);
xor U13157 (N_13157,N_12869,N_12879);
xor U13158 (N_13158,N_12871,N_12721);
nor U13159 (N_13159,N_12520,N_12933);
nor U13160 (N_13160,N_12823,N_12674);
xor U13161 (N_13161,N_12841,N_12836);
nor U13162 (N_13162,N_12843,N_12528);
nand U13163 (N_13163,N_12877,N_12928);
or U13164 (N_13164,N_12575,N_12737);
or U13165 (N_13165,N_12774,N_12693);
and U13166 (N_13166,N_12921,N_12724);
nand U13167 (N_13167,N_12905,N_12624);
nand U13168 (N_13168,N_12947,N_12826);
nor U13169 (N_13169,N_12870,N_12873);
nand U13170 (N_13170,N_12664,N_12829);
or U13171 (N_13171,N_12995,N_12786);
and U13172 (N_13172,N_12618,N_12670);
xor U13173 (N_13173,N_12518,N_12522);
and U13174 (N_13174,N_12944,N_12968);
nand U13175 (N_13175,N_12640,N_12655);
nand U13176 (N_13176,N_12849,N_12504);
nand U13177 (N_13177,N_12875,N_12953);
nor U13178 (N_13178,N_12903,N_12688);
and U13179 (N_13179,N_12702,N_12902);
nand U13180 (N_13180,N_12762,N_12646);
nand U13181 (N_13181,N_12725,N_12942);
xor U13182 (N_13182,N_12631,N_12749);
nor U13183 (N_13183,N_12927,N_12965);
nor U13184 (N_13184,N_12967,N_12810);
and U13185 (N_13185,N_12549,N_12578);
nor U13186 (N_13186,N_12566,N_12897);
nor U13187 (N_13187,N_12924,N_12508);
nor U13188 (N_13188,N_12894,N_12628);
nor U13189 (N_13189,N_12833,N_12699);
nand U13190 (N_13190,N_12952,N_12745);
xor U13191 (N_13191,N_12866,N_12812);
and U13192 (N_13192,N_12529,N_12687);
and U13193 (N_13193,N_12600,N_12753);
or U13194 (N_13194,N_12734,N_12765);
or U13195 (N_13195,N_12613,N_12534);
nand U13196 (N_13196,N_12977,N_12983);
nand U13197 (N_13197,N_12925,N_12564);
nand U13198 (N_13198,N_12513,N_12514);
or U13199 (N_13199,N_12568,N_12949);
xor U13200 (N_13200,N_12608,N_12980);
nand U13201 (N_13201,N_12909,N_12503);
xnor U13202 (N_13202,N_12705,N_12598);
nand U13203 (N_13203,N_12827,N_12710);
or U13204 (N_13204,N_12621,N_12711);
and U13205 (N_13205,N_12572,N_12551);
and U13206 (N_13206,N_12929,N_12806);
or U13207 (N_13207,N_12916,N_12919);
nor U13208 (N_13208,N_12960,N_12537);
and U13209 (N_13209,N_12679,N_12906);
nor U13210 (N_13210,N_12675,N_12992);
or U13211 (N_13211,N_12912,N_12708);
xor U13212 (N_13212,N_12585,N_12714);
and U13213 (N_13213,N_12569,N_12835);
nor U13214 (N_13214,N_12556,N_12533);
xnor U13215 (N_13215,N_12955,N_12918);
xor U13216 (N_13216,N_12559,N_12643);
nor U13217 (N_13217,N_12979,N_12561);
and U13218 (N_13218,N_12884,N_12987);
nand U13219 (N_13219,N_12888,N_12647);
and U13220 (N_13220,N_12507,N_12807);
nand U13221 (N_13221,N_12868,N_12703);
nor U13222 (N_13222,N_12881,N_12991);
nor U13223 (N_13223,N_12820,N_12941);
and U13224 (N_13224,N_12985,N_12576);
nor U13225 (N_13225,N_12932,N_12825);
or U13226 (N_13226,N_12726,N_12686);
or U13227 (N_13227,N_12805,N_12689);
xnor U13228 (N_13228,N_12707,N_12998);
nand U13229 (N_13229,N_12954,N_12857);
or U13230 (N_13230,N_12596,N_12532);
xor U13231 (N_13231,N_12865,N_12800);
and U13232 (N_13232,N_12727,N_12887);
nand U13233 (N_13233,N_12648,N_12978);
nor U13234 (N_13234,N_12811,N_12808);
nand U13235 (N_13235,N_12899,N_12972);
nand U13236 (N_13236,N_12713,N_12584);
xor U13237 (N_13237,N_12659,N_12622);
and U13238 (N_13238,N_12896,N_12788);
xor U13239 (N_13239,N_12565,N_12989);
xor U13240 (N_13240,N_12602,N_12604);
or U13241 (N_13241,N_12509,N_12729);
xor U13242 (N_13242,N_12661,N_12770);
xnor U13243 (N_13243,N_12922,N_12720);
nor U13244 (N_13244,N_12555,N_12872);
and U13245 (N_13245,N_12755,N_12653);
nand U13246 (N_13246,N_12876,N_12996);
or U13247 (N_13247,N_12700,N_12939);
or U13248 (N_13248,N_12885,N_12681);
or U13249 (N_13249,N_12981,N_12633);
and U13250 (N_13250,N_12690,N_12550);
nand U13251 (N_13251,N_12985,N_12683);
nand U13252 (N_13252,N_12856,N_12676);
and U13253 (N_13253,N_12776,N_12850);
and U13254 (N_13254,N_12593,N_12875);
xnor U13255 (N_13255,N_12577,N_12848);
nand U13256 (N_13256,N_12706,N_12606);
nand U13257 (N_13257,N_12618,N_12810);
nor U13258 (N_13258,N_12990,N_12783);
nand U13259 (N_13259,N_12618,N_12792);
nand U13260 (N_13260,N_12616,N_12943);
and U13261 (N_13261,N_12991,N_12835);
nor U13262 (N_13262,N_12591,N_12928);
nand U13263 (N_13263,N_12580,N_12697);
and U13264 (N_13264,N_12877,N_12687);
or U13265 (N_13265,N_12860,N_12595);
xor U13266 (N_13266,N_12748,N_12687);
xor U13267 (N_13267,N_12750,N_12927);
or U13268 (N_13268,N_12678,N_12501);
nor U13269 (N_13269,N_12671,N_12859);
nand U13270 (N_13270,N_12820,N_12701);
or U13271 (N_13271,N_12684,N_12537);
nand U13272 (N_13272,N_12804,N_12864);
nor U13273 (N_13273,N_12752,N_12892);
or U13274 (N_13274,N_12949,N_12631);
and U13275 (N_13275,N_12712,N_12764);
and U13276 (N_13276,N_12611,N_12807);
and U13277 (N_13277,N_12930,N_12792);
or U13278 (N_13278,N_12742,N_12968);
nor U13279 (N_13279,N_12948,N_12595);
nand U13280 (N_13280,N_12695,N_12820);
nand U13281 (N_13281,N_12861,N_12821);
xnor U13282 (N_13282,N_12872,N_12999);
nand U13283 (N_13283,N_12998,N_12865);
and U13284 (N_13284,N_12585,N_12771);
nor U13285 (N_13285,N_12549,N_12778);
nand U13286 (N_13286,N_12828,N_12925);
or U13287 (N_13287,N_12509,N_12866);
nor U13288 (N_13288,N_12798,N_12848);
or U13289 (N_13289,N_12781,N_12540);
xor U13290 (N_13290,N_12843,N_12826);
and U13291 (N_13291,N_12549,N_12680);
xor U13292 (N_13292,N_12924,N_12709);
nor U13293 (N_13293,N_12866,N_12612);
nor U13294 (N_13294,N_12522,N_12538);
nand U13295 (N_13295,N_12642,N_12838);
nor U13296 (N_13296,N_12579,N_12636);
nand U13297 (N_13297,N_12985,N_12848);
and U13298 (N_13298,N_12634,N_12530);
xor U13299 (N_13299,N_12810,N_12960);
or U13300 (N_13300,N_12969,N_12636);
xor U13301 (N_13301,N_12737,N_12924);
nor U13302 (N_13302,N_12988,N_12966);
or U13303 (N_13303,N_12796,N_12714);
xnor U13304 (N_13304,N_12833,N_12585);
nor U13305 (N_13305,N_12930,N_12639);
or U13306 (N_13306,N_12783,N_12734);
xor U13307 (N_13307,N_12733,N_12937);
nor U13308 (N_13308,N_12787,N_12761);
and U13309 (N_13309,N_12810,N_12805);
nor U13310 (N_13310,N_12795,N_12563);
xnor U13311 (N_13311,N_12528,N_12819);
xnor U13312 (N_13312,N_12809,N_12901);
and U13313 (N_13313,N_12694,N_12859);
nor U13314 (N_13314,N_12591,N_12815);
and U13315 (N_13315,N_12708,N_12999);
nand U13316 (N_13316,N_12535,N_12621);
or U13317 (N_13317,N_12742,N_12863);
nand U13318 (N_13318,N_12873,N_12506);
nor U13319 (N_13319,N_12696,N_12752);
nor U13320 (N_13320,N_12681,N_12992);
nand U13321 (N_13321,N_12526,N_12522);
or U13322 (N_13322,N_12557,N_12964);
nor U13323 (N_13323,N_12656,N_12742);
nor U13324 (N_13324,N_12693,N_12819);
xnor U13325 (N_13325,N_12704,N_12614);
xnor U13326 (N_13326,N_12542,N_12669);
nor U13327 (N_13327,N_12679,N_12950);
nor U13328 (N_13328,N_12803,N_12919);
nand U13329 (N_13329,N_12970,N_12532);
or U13330 (N_13330,N_12912,N_12909);
xor U13331 (N_13331,N_12903,N_12836);
and U13332 (N_13332,N_12863,N_12934);
nor U13333 (N_13333,N_12682,N_12509);
or U13334 (N_13334,N_12696,N_12746);
or U13335 (N_13335,N_12953,N_12723);
or U13336 (N_13336,N_12840,N_12851);
or U13337 (N_13337,N_12766,N_12690);
or U13338 (N_13338,N_12826,N_12592);
and U13339 (N_13339,N_12817,N_12546);
nand U13340 (N_13340,N_12756,N_12897);
xnor U13341 (N_13341,N_12732,N_12718);
xor U13342 (N_13342,N_12797,N_12807);
xnor U13343 (N_13343,N_12690,N_12714);
and U13344 (N_13344,N_12555,N_12994);
xnor U13345 (N_13345,N_12684,N_12780);
xor U13346 (N_13346,N_12918,N_12669);
nand U13347 (N_13347,N_12733,N_12621);
and U13348 (N_13348,N_12967,N_12700);
nand U13349 (N_13349,N_12596,N_12628);
nand U13350 (N_13350,N_12835,N_12578);
or U13351 (N_13351,N_12877,N_12541);
nand U13352 (N_13352,N_12758,N_12852);
and U13353 (N_13353,N_12755,N_12685);
or U13354 (N_13354,N_12966,N_12987);
or U13355 (N_13355,N_12737,N_12962);
xnor U13356 (N_13356,N_12587,N_12521);
xnor U13357 (N_13357,N_12718,N_12740);
nor U13358 (N_13358,N_12641,N_12797);
xor U13359 (N_13359,N_12573,N_12906);
nand U13360 (N_13360,N_12920,N_12786);
or U13361 (N_13361,N_12965,N_12609);
nor U13362 (N_13362,N_12654,N_12767);
or U13363 (N_13363,N_12655,N_12947);
and U13364 (N_13364,N_12679,N_12987);
xnor U13365 (N_13365,N_12739,N_12582);
and U13366 (N_13366,N_12738,N_12816);
xor U13367 (N_13367,N_12865,N_12787);
xnor U13368 (N_13368,N_12573,N_12982);
xor U13369 (N_13369,N_12509,N_12515);
or U13370 (N_13370,N_12937,N_12638);
nand U13371 (N_13371,N_12656,N_12874);
or U13372 (N_13372,N_12751,N_12761);
and U13373 (N_13373,N_12704,N_12899);
xor U13374 (N_13374,N_12913,N_12559);
nor U13375 (N_13375,N_12534,N_12895);
nor U13376 (N_13376,N_12961,N_12600);
and U13377 (N_13377,N_12813,N_12921);
nor U13378 (N_13378,N_12884,N_12551);
xor U13379 (N_13379,N_12846,N_12931);
xnor U13380 (N_13380,N_12549,N_12713);
nand U13381 (N_13381,N_12729,N_12947);
and U13382 (N_13382,N_12763,N_12956);
or U13383 (N_13383,N_12755,N_12851);
or U13384 (N_13384,N_12566,N_12673);
or U13385 (N_13385,N_12678,N_12664);
xor U13386 (N_13386,N_12660,N_12670);
nor U13387 (N_13387,N_12808,N_12636);
and U13388 (N_13388,N_12513,N_12990);
nor U13389 (N_13389,N_12660,N_12585);
xor U13390 (N_13390,N_12607,N_12985);
xor U13391 (N_13391,N_12579,N_12677);
nor U13392 (N_13392,N_12705,N_12534);
nor U13393 (N_13393,N_12875,N_12569);
nand U13394 (N_13394,N_12582,N_12715);
nor U13395 (N_13395,N_12764,N_12931);
xnor U13396 (N_13396,N_12816,N_12867);
xnor U13397 (N_13397,N_12552,N_12638);
nor U13398 (N_13398,N_12756,N_12694);
xor U13399 (N_13399,N_12647,N_12653);
nor U13400 (N_13400,N_12844,N_12726);
nand U13401 (N_13401,N_12873,N_12735);
or U13402 (N_13402,N_12764,N_12590);
and U13403 (N_13403,N_12838,N_12717);
nand U13404 (N_13404,N_12822,N_12791);
and U13405 (N_13405,N_12996,N_12636);
and U13406 (N_13406,N_12964,N_12994);
nor U13407 (N_13407,N_12655,N_12662);
nand U13408 (N_13408,N_12815,N_12796);
and U13409 (N_13409,N_12996,N_12869);
xnor U13410 (N_13410,N_12524,N_12602);
nor U13411 (N_13411,N_12696,N_12869);
xnor U13412 (N_13412,N_12814,N_12904);
xor U13413 (N_13413,N_12676,N_12719);
or U13414 (N_13414,N_12542,N_12528);
and U13415 (N_13415,N_12908,N_12724);
xor U13416 (N_13416,N_12514,N_12594);
xor U13417 (N_13417,N_12946,N_12983);
xor U13418 (N_13418,N_12645,N_12872);
and U13419 (N_13419,N_12947,N_12687);
nor U13420 (N_13420,N_12809,N_12951);
and U13421 (N_13421,N_12948,N_12688);
and U13422 (N_13422,N_12725,N_12946);
nor U13423 (N_13423,N_12800,N_12937);
nor U13424 (N_13424,N_12894,N_12643);
xor U13425 (N_13425,N_12987,N_12893);
nor U13426 (N_13426,N_12755,N_12785);
nand U13427 (N_13427,N_12934,N_12837);
nor U13428 (N_13428,N_12503,N_12522);
and U13429 (N_13429,N_12662,N_12539);
nor U13430 (N_13430,N_12601,N_12982);
xnor U13431 (N_13431,N_12933,N_12500);
nand U13432 (N_13432,N_12729,N_12658);
and U13433 (N_13433,N_12600,N_12840);
xnor U13434 (N_13434,N_12658,N_12722);
xor U13435 (N_13435,N_12762,N_12854);
xnor U13436 (N_13436,N_12688,N_12844);
nand U13437 (N_13437,N_12812,N_12834);
and U13438 (N_13438,N_12582,N_12706);
nand U13439 (N_13439,N_12999,N_12965);
xor U13440 (N_13440,N_12894,N_12925);
nor U13441 (N_13441,N_12510,N_12587);
nand U13442 (N_13442,N_12837,N_12680);
xnor U13443 (N_13443,N_12618,N_12953);
nor U13444 (N_13444,N_12951,N_12865);
nand U13445 (N_13445,N_12566,N_12761);
nor U13446 (N_13446,N_12862,N_12730);
and U13447 (N_13447,N_12860,N_12740);
nor U13448 (N_13448,N_12935,N_12853);
or U13449 (N_13449,N_12900,N_12603);
xor U13450 (N_13450,N_12560,N_12919);
nor U13451 (N_13451,N_12838,N_12556);
nand U13452 (N_13452,N_12729,N_12820);
xnor U13453 (N_13453,N_12607,N_12669);
nor U13454 (N_13454,N_12794,N_12811);
xor U13455 (N_13455,N_12670,N_12979);
or U13456 (N_13456,N_12720,N_12719);
xnor U13457 (N_13457,N_12960,N_12528);
nand U13458 (N_13458,N_12550,N_12754);
or U13459 (N_13459,N_12572,N_12926);
and U13460 (N_13460,N_12551,N_12503);
nor U13461 (N_13461,N_12516,N_12512);
and U13462 (N_13462,N_12776,N_12800);
and U13463 (N_13463,N_12912,N_12841);
nor U13464 (N_13464,N_12738,N_12916);
or U13465 (N_13465,N_12842,N_12997);
nor U13466 (N_13466,N_12517,N_12827);
or U13467 (N_13467,N_12643,N_12718);
and U13468 (N_13468,N_12525,N_12502);
nor U13469 (N_13469,N_12779,N_12915);
nand U13470 (N_13470,N_12617,N_12669);
or U13471 (N_13471,N_12552,N_12919);
xor U13472 (N_13472,N_12543,N_12908);
nor U13473 (N_13473,N_12785,N_12550);
xnor U13474 (N_13474,N_12872,N_12739);
nor U13475 (N_13475,N_12577,N_12647);
and U13476 (N_13476,N_12570,N_12554);
or U13477 (N_13477,N_12620,N_12902);
or U13478 (N_13478,N_12941,N_12611);
and U13479 (N_13479,N_12606,N_12967);
nor U13480 (N_13480,N_12746,N_12922);
nor U13481 (N_13481,N_12684,N_12804);
or U13482 (N_13482,N_12524,N_12607);
nor U13483 (N_13483,N_12515,N_12709);
nor U13484 (N_13484,N_12935,N_12970);
nand U13485 (N_13485,N_12531,N_12734);
or U13486 (N_13486,N_12793,N_12803);
and U13487 (N_13487,N_12912,N_12567);
xnor U13488 (N_13488,N_12864,N_12510);
nand U13489 (N_13489,N_12513,N_12953);
or U13490 (N_13490,N_12912,N_12636);
or U13491 (N_13491,N_12601,N_12793);
nand U13492 (N_13492,N_12549,N_12710);
nor U13493 (N_13493,N_12636,N_12855);
nor U13494 (N_13494,N_12858,N_12942);
and U13495 (N_13495,N_12907,N_12981);
or U13496 (N_13496,N_12704,N_12517);
nor U13497 (N_13497,N_12831,N_12964);
nor U13498 (N_13498,N_12648,N_12569);
nor U13499 (N_13499,N_12852,N_12627);
xor U13500 (N_13500,N_13195,N_13022);
xnor U13501 (N_13501,N_13310,N_13163);
and U13502 (N_13502,N_13235,N_13350);
and U13503 (N_13503,N_13026,N_13048);
xor U13504 (N_13504,N_13442,N_13066);
nand U13505 (N_13505,N_13327,N_13402);
nor U13506 (N_13506,N_13352,N_13485);
and U13507 (N_13507,N_13256,N_13435);
and U13508 (N_13508,N_13103,N_13076);
nor U13509 (N_13509,N_13030,N_13390);
nor U13510 (N_13510,N_13481,N_13252);
and U13511 (N_13511,N_13192,N_13112);
xor U13512 (N_13512,N_13108,N_13330);
and U13513 (N_13513,N_13216,N_13148);
xor U13514 (N_13514,N_13271,N_13362);
nor U13515 (N_13515,N_13068,N_13196);
xor U13516 (N_13516,N_13110,N_13170);
xor U13517 (N_13517,N_13198,N_13044);
or U13518 (N_13518,N_13418,N_13344);
xnor U13519 (N_13519,N_13345,N_13420);
nor U13520 (N_13520,N_13028,N_13392);
xnor U13521 (N_13521,N_13070,N_13241);
and U13522 (N_13522,N_13228,N_13100);
or U13523 (N_13523,N_13062,N_13398);
and U13524 (N_13524,N_13126,N_13449);
nor U13525 (N_13525,N_13171,N_13412);
and U13526 (N_13526,N_13224,N_13272);
and U13527 (N_13527,N_13024,N_13492);
nor U13528 (N_13528,N_13243,N_13475);
and U13529 (N_13529,N_13354,N_13431);
nand U13530 (N_13530,N_13031,N_13166);
and U13531 (N_13531,N_13490,N_13169);
or U13532 (N_13532,N_13416,N_13270);
xor U13533 (N_13533,N_13225,N_13489);
nand U13534 (N_13534,N_13377,N_13125);
xnor U13535 (N_13535,N_13358,N_13432);
or U13536 (N_13536,N_13079,N_13214);
and U13537 (N_13537,N_13251,N_13367);
nor U13538 (N_13538,N_13208,N_13237);
and U13539 (N_13539,N_13427,N_13054);
nor U13540 (N_13540,N_13080,N_13133);
and U13541 (N_13541,N_13380,N_13387);
xor U13542 (N_13542,N_13211,N_13356);
or U13543 (N_13543,N_13283,N_13290);
nor U13544 (N_13544,N_13307,N_13257);
xnor U13545 (N_13545,N_13494,N_13471);
nor U13546 (N_13546,N_13353,N_13071);
or U13547 (N_13547,N_13084,N_13274);
nor U13548 (N_13548,N_13246,N_13113);
xnor U13549 (N_13549,N_13312,N_13083);
or U13550 (N_13550,N_13158,N_13462);
or U13551 (N_13551,N_13222,N_13029);
or U13552 (N_13552,N_13458,N_13324);
or U13553 (N_13553,N_13127,N_13003);
xnor U13554 (N_13554,N_13314,N_13039);
xor U13555 (N_13555,N_13315,N_13207);
or U13556 (N_13556,N_13326,N_13154);
nor U13557 (N_13557,N_13182,N_13351);
xor U13558 (N_13558,N_13409,N_13428);
or U13559 (N_13559,N_13000,N_13088);
or U13560 (N_13560,N_13036,N_13093);
nand U13561 (N_13561,N_13499,N_13020);
or U13562 (N_13562,N_13332,N_13346);
nor U13563 (N_13563,N_13366,N_13466);
xor U13564 (N_13564,N_13253,N_13321);
nand U13565 (N_13565,N_13201,N_13065);
nor U13566 (N_13566,N_13189,N_13450);
xor U13567 (N_13567,N_13419,N_13160);
and U13568 (N_13568,N_13111,N_13331);
or U13569 (N_13569,N_13049,N_13372);
xor U13570 (N_13570,N_13035,N_13284);
nor U13571 (N_13571,N_13027,N_13212);
nor U13572 (N_13572,N_13259,N_13102);
nand U13573 (N_13573,N_13297,N_13313);
or U13574 (N_13574,N_13109,N_13338);
nor U13575 (N_13575,N_13437,N_13286);
nand U13576 (N_13576,N_13115,N_13339);
nand U13577 (N_13577,N_13004,N_13382);
nor U13578 (N_13578,N_13242,N_13269);
or U13579 (N_13579,N_13145,N_13064);
and U13580 (N_13580,N_13384,N_13091);
nor U13581 (N_13581,N_13082,N_13188);
nand U13582 (N_13582,N_13142,N_13299);
xor U13583 (N_13583,N_13470,N_13176);
and U13584 (N_13584,N_13230,N_13368);
nor U13585 (N_13585,N_13441,N_13119);
nor U13586 (N_13586,N_13168,N_13317);
or U13587 (N_13587,N_13484,N_13394);
or U13588 (N_13588,N_13060,N_13033);
nand U13589 (N_13589,N_13149,N_13130);
xnor U13590 (N_13590,N_13407,N_13135);
nor U13591 (N_13591,N_13165,N_13401);
nand U13592 (N_13592,N_13151,N_13092);
or U13593 (N_13593,N_13177,N_13159);
nor U13594 (N_13594,N_13219,N_13006);
nor U13595 (N_13595,N_13138,N_13063);
nor U13596 (N_13596,N_13194,N_13280);
nor U13597 (N_13597,N_13282,N_13478);
or U13598 (N_13598,N_13007,N_13287);
nor U13599 (N_13599,N_13175,N_13476);
nand U13600 (N_13600,N_13129,N_13231);
xor U13601 (N_13601,N_13337,N_13061);
and U13602 (N_13602,N_13204,N_13279);
nor U13603 (N_13603,N_13429,N_13482);
nand U13604 (N_13604,N_13370,N_13185);
xnor U13605 (N_13605,N_13005,N_13278);
and U13606 (N_13606,N_13468,N_13069);
and U13607 (N_13607,N_13008,N_13364);
or U13608 (N_13608,N_13172,N_13474);
nor U13609 (N_13609,N_13067,N_13463);
nor U13610 (N_13610,N_13303,N_13452);
xor U13611 (N_13611,N_13085,N_13023);
and U13612 (N_13612,N_13203,N_13221);
nand U13613 (N_13613,N_13388,N_13098);
or U13614 (N_13614,N_13335,N_13050);
xnor U13615 (N_13615,N_13086,N_13021);
xor U13616 (N_13616,N_13493,N_13001);
nor U13617 (N_13617,N_13247,N_13043);
nand U13618 (N_13618,N_13360,N_13379);
xor U13619 (N_13619,N_13376,N_13487);
nor U13620 (N_13620,N_13095,N_13164);
and U13621 (N_13621,N_13014,N_13465);
nor U13622 (N_13622,N_13396,N_13381);
nand U13623 (N_13623,N_13446,N_13473);
xnor U13624 (N_13624,N_13461,N_13025);
nor U13625 (N_13625,N_13190,N_13105);
nand U13626 (N_13626,N_13017,N_13155);
or U13627 (N_13627,N_13180,N_13289);
xor U13628 (N_13628,N_13308,N_13209);
xor U13629 (N_13629,N_13359,N_13268);
and U13630 (N_13630,N_13161,N_13288);
nor U13631 (N_13631,N_13264,N_13137);
or U13632 (N_13632,N_13117,N_13052);
nor U13633 (N_13633,N_13144,N_13174);
and U13634 (N_13634,N_13275,N_13298);
and U13635 (N_13635,N_13425,N_13496);
and U13636 (N_13636,N_13254,N_13019);
and U13637 (N_13637,N_13232,N_13213);
nor U13638 (N_13638,N_13248,N_13229);
or U13639 (N_13639,N_13267,N_13236);
xor U13640 (N_13640,N_13143,N_13118);
nand U13641 (N_13641,N_13097,N_13488);
xor U13642 (N_13642,N_13385,N_13460);
or U13643 (N_13643,N_13319,N_13122);
xor U13644 (N_13644,N_13276,N_13309);
nor U13645 (N_13645,N_13002,N_13106);
xor U13646 (N_13646,N_13051,N_13032);
nor U13647 (N_13647,N_13059,N_13277);
or U13648 (N_13648,N_13491,N_13405);
or U13649 (N_13649,N_13438,N_13316);
or U13650 (N_13650,N_13453,N_13467);
nand U13651 (N_13651,N_13087,N_13389);
nand U13652 (N_13652,N_13311,N_13245);
and U13653 (N_13653,N_13220,N_13325);
nand U13654 (N_13654,N_13090,N_13451);
or U13655 (N_13655,N_13104,N_13294);
xor U13656 (N_13656,N_13304,N_13393);
nand U13657 (N_13657,N_13016,N_13322);
nand U13658 (N_13658,N_13415,N_13058);
or U13659 (N_13659,N_13413,N_13469);
and U13660 (N_13660,N_13099,N_13479);
and U13661 (N_13661,N_13053,N_13472);
or U13662 (N_13662,N_13012,N_13357);
or U13663 (N_13663,N_13217,N_13340);
or U13664 (N_13664,N_13375,N_13408);
nor U13665 (N_13665,N_13013,N_13300);
and U13666 (N_13666,N_13434,N_13101);
nand U13667 (N_13667,N_13009,N_13261);
nor U13668 (N_13668,N_13329,N_13038);
xnor U13669 (N_13669,N_13223,N_13081);
xor U13670 (N_13670,N_13342,N_13128);
nor U13671 (N_13671,N_13162,N_13191);
nand U13672 (N_13672,N_13404,N_13439);
nand U13673 (N_13673,N_13226,N_13328);
xnor U13674 (N_13674,N_13459,N_13197);
nor U13675 (N_13675,N_13255,N_13132);
nand U13676 (N_13676,N_13395,N_13134);
nor U13677 (N_13677,N_13077,N_13089);
xor U13678 (N_13678,N_13378,N_13424);
xor U13679 (N_13679,N_13301,N_13262);
nor U13680 (N_13680,N_13187,N_13260);
xor U13681 (N_13681,N_13233,N_13045);
nand U13682 (N_13682,N_13399,N_13239);
xnor U13683 (N_13683,N_13373,N_13445);
nor U13684 (N_13684,N_13293,N_13422);
or U13685 (N_13685,N_13285,N_13140);
xnor U13686 (N_13686,N_13041,N_13363);
nor U13687 (N_13687,N_13464,N_13440);
and U13688 (N_13688,N_13250,N_13010);
nor U13689 (N_13689,N_13107,N_13075);
or U13690 (N_13690,N_13047,N_13056);
nand U13691 (N_13691,N_13347,N_13249);
nand U13692 (N_13692,N_13200,N_13057);
xnor U13693 (N_13693,N_13240,N_13486);
or U13694 (N_13694,N_13199,N_13495);
nor U13695 (N_13695,N_13034,N_13391);
nand U13696 (N_13696,N_13234,N_13258);
nor U13697 (N_13697,N_13114,N_13320);
nand U13698 (N_13698,N_13406,N_13497);
xor U13699 (N_13699,N_13266,N_13210);
or U13700 (N_13700,N_13073,N_13131);
and U13701 (N_13701,N_13433,N_13281);
nand U13702 (N_13702,N_13193,N_13349);
nor U13703 (N_13703,N_13265,N_13318);
or U13704 (N_13704,N_13116,N_13238);
xor U13705 (N_13705,N_13123,N_13343);
or U13706 (N_13706,N_13120,N_13410);
xor U13707 (N_13707,N_13386,N_13477);
or U13708 (N_13708,N_13206,N_13157);
xor U13709 (N_13709,N_13306,N_13423);
nand U13710 (N_13710,N_13295,N_13178);
nand U13711 (N_13711,N_13333,N_13417);
xor U13712 (N_13712,N_13454,N_13152);
or U13713 (N_13713,N_13096,N_13218);
nor U13714 (N_13714,N_13444,N_13397);
and U13715 (N_13715,N_13323,N_13167);
and U13716 (N_13716,N_13150,N_13121);
xnor U13717 (N_13717,N_13436,N_13400);
and U13718 (N_13718,N_13273,N_13348);
nor U13719 (N_13719,N_13336,N_13365);
xor U13720 (N_13720,N_13205,N_13074);
or U13721 (N_13721,N_13186,N_13173);
nor U13722 (N_13722,N_13046,N_13341);
nand U13723 (N_13723,N_13456,N_13072);
nor U13724 (N_13724,N_13296,N_13302);
nand U13725 (N_13725,N_13139,N_13227);
and U13726 (N_13726,N_13037,N_13153);
xor U13727 (N_13727,N_13443,N_13430);
or U13728 (N_13728,N_13078,N_13011);
xnor U13729 (N_13729,N_13136,N_13371);
xor U13730 (N_13730,N_13291,N_13403);
or U13731 (N_13731,N_13498,N_13355);
xnor U13732 (N_13732,N_13215,N_13179);
nand U13733 (N_13733,N_13369,N_13124);
nand U13734 (N_13734,N_13202,N_13414);
xor U13735 (N_13735,N_13244,N_13292);
xnor U13736 (N_13736,N_13042,N_13305);
nand U13737 (N_13737,N_13146,N_13015);
nor U13738 (N_13738,N_13181,N_13455);
and U13739 (N_13739,N_13184,N_13263);
and U13740 (N_13740,N_13040,N_13018);
xor U13741 (N_13741,N_13426,N_13334);
xor U13742 (N_13742,N_13483,N_13421);
nor U13743 (N_13743,N_13457,N_13383);
xor U13744 (N_13744,N_13447,N_13480);
xnor U13745 (N_13745,N_13156,N_13374);
nand U13746 (N_13746,N_13411,N_13055);
xor U13747 (N_13747,N_13141,N_13448);
and U13748 (N_13748,N_13183,N_13094);
nor U13749 (N_13749,N_13147,N_13361);
nor U13750 (N_13750,N_13409,N_13417);
and U13751 (N_13751,N_13309,N_13280);
nand U13752 (N_13752,N_13154,N_13433);
xor U13753 (N_13753,N_13464,N_13091);
and U13754 (N_13754,N_13231,N_13086);
nor U13755 (N_13755,N_13243,N_13372);
xor U13756 (N_13756,N_13160,N_13271);
nor U13757 (N_13757,N_13092,N_13283);
or U13758 (N_13758,N_13150,N_13073);
xnor U13759 (N_13759,N_13446,N_13090);
and U13760 (N_13760,N_13005,N_13092);
or U13761 (N_13761,N_13453,N_13137);
xnor U13762 (N_13762,N_13349,N_13152);
and U13763 (N_13763,N_13147,N_13314);
and U13764 (N_13764,N_13128,N_13477);
and U13765 (N_13765,N_13193,N_13181);
and U13766 (N_13766,N_13013,N_13080);
nand U13767 (N_13767,N_13040,N_13127);
nand U13768 (N_13768,N_13021,N_13429);
nand U13769 (N_13769,N_13453,N_13478);
nand U13770 (N_13770,N_13160,N_13262);
or U13771 (N_13771,N_13336,N_13192);
and U13772 (N_13772,N_13046,N_13249);
nand U13773 (N_13773,N_13310,N_13364);
nor U13774 (N_13774,N_13018,N_13246);
xnor U13775 (N_13775,N_13168,N_13233);
or U13776 (N_13776,N_13255,N_13016);
and U13777 (N_13777,N_13337,N_13212);
nand U13778 (N_13778,N_13022,N_13226);
or U13779 (N_13779,N_13161,N_13177);
and U13780 (N_13780,N_13133,N_13444);
nor U13781 (N_13781,N_13348,N_13013);
and U13782 (N_13782,N_13044,N_13087);
or U13783 (N_13783,N_13261,N_13118);
xor U13784 (N_13784,N_13124,N_13022);
xor U13785 (N_13785,N_13451,N_13147);
nand U13786 (N_13786,N_13404,N_13051);
nand U13787 (N_13787,N_13216,N_13199);
nand U13788 (N_13788,N_13028,N_13083);
or U13789 (N_13789,N_13145,N_13104);
or U13790 (N_13790,N_13228,N_13345);
and U13791 (N_13791,N_13430,N_13108);
and U13792 (N_13792,N_13491,N_13056);
and U13793 (N_13793,N_13307,N_13248);
and U13794 (N_13794,N_13066,N_13027);
xor U13795 (N_13795,N_13386,N_13400);
xor U13796 (N_13796,N_13488,N_13076);
nand U13797 (N_13797,N_13205,N_13365);
nand U13798 (N_13798,N_13119,N_13453);
xnor U13799 (N_13799,N_13286,N_13440);
nor U13800 (N_13800,N_13274,N_13163);
nand U13801 (N_13801,N_13465,N_13367);
or U13802 (N_13802,N_13046,N_13317);
or U13803 (N_13803,N_13459,N_13436);
xnor U13804 (N_13804,N_13144,N_13307);
or U13805 (N_13805,N_13054,N_13196);
xor U13806 (N_13806,N_13056,N_13452);
nor U13807 (N_13807,N_13165,N_13106);
xor U13808 (N_13808,N_13349,N_13442);
xnor U13809 (N_13809,N_13308,N_13051);
nor U13810 (N_13810,N_13266,N_13324);
nor U13811 (N_13811,N_13372,N_13026);
nand U13812 (N_13812,N_13144,N_13325);
and U13813 (N_13813,N_13165,N_13351);
nor U13814 (N_13814,N_13402,N_13394);
nor U13815 (N_13815,N_13033,N_13163);
nand U13816 (N_13816,N_13102,N_13493);
and U13817 (N_13817,N_13204,N_13112);
and U13818 (N_13818,N_13249,N_13214);
and U13819 (N_13819,N_13042,N_13358);
nor U13820 (N_13820,N_13087,N_13162);
and U13821 (N_13821,N_13205,N_13126);
nor U13822 (N_13822,N_13177,N_13003);
and U13823 (N_13823,N_13062,N_13238);
nor U13824 (N_13824,N_13344,N_13470);
and U13825 (N_13825,N_13258,N_13215);
nor U13826 (N_13826,N_13068,N_13487);
or U13827 (N_13827,N_13084,N_13068);
nand U13828 (N_13828,N_13148,N_13091);
nand U13829 (N_13829,N_13172,N_13487);
nor U13830 (N_13830,N_13358,N_13192);
nand U13831 (N_13831,N_13423,N_13470);
nand U13832 (N_13832,N_13184,N_13343);
or U13833 (N_13833,N_13104,N_13197);
or U13834 (N_13834,N_13281,N_13259);
and U13835 (N_13835,N_13032,N_13228);
and U13836 (N_13836,N_13376,N_13443);
and U13837 (N_13837,N_13007,N_13163);
and U13838 (N_13838,N_13135,N_13148);
or U13839 (N_13839,N_13106,N_13083);
xnor U13840 (N_13840,N_13254,N_13343);
or U13841 (N_13841,N_13039,N_13262);
nand U13842 (N_13842,N_13323,N_13059);
xor U13843 (N_13843,N_13268,N_13128);
nand U13844 (N_13844,N_13086,N_13413);
and U13845 (N_13845,N_13413,N_13329);
nand U13846 (N_13846,N_13106,N_13345);
nand U13847 (N_13847,N_13216,N_13240);
nor U13848 (N_13848,N_13237,N_13235);
xnor U13849 (N_13849,N_13122,N_13224);
nor U13850 (N_13850,N_13005,N_13373);
nand U13851 (N_13851,N_13362,N_13413);
nor U13852 (N_13852,N_13073,N_13151);
nor U13853 (N_13853,N_13245,N_13338);
or U13854 (N_13854,N_13060,N_13389);
or U13855 (N_13855,N_13371,N_13419);
xor U13856 (N_13856,N_13289,N_13275);
nand U13857 (N_13857,N_13486,N_13471);
or U13858 (N_13858,N_13400,N_13178);
xor U13859 (N_13859,N_13133,N_13482);
nor U13860 (N_13860,N_13359,N_13005);
or U13861 (N_13861,N_13288,N_13323);
nor U13862 (N_13862,N_13291,N_13136);
nor U13863 (N_13863,N_13045,N_13310);
or U13864 (N_13864,N_13473,N_13479);
and U13865 (N_13865,N_13385,N_13328);
or U13866 (N_13866,N_13252,N_13409);
nand U13867 (N_13867,N_13227,N_13338);
and U13868 (N_13868,N_13187,N_13007);
nor U13869 (N_13869,N_13299,N_13230);
nor U13870 (N_13870,N_13484,N_13458);
or U13871 (N_13871,N_13368,N_13254);
and U13872 (N_13872,N_13047,N_13232);
xor U13873 (N_13873,N_13255,N_13368);
nor U13874 (N_13874,N_13349,N_13329);
or U13875 (N_13875,N_13173,N_13475);
xor U13876 (N_13876,N_13426,N_13261);
or U13877 (N_13877,N_13102,N_13106);
xnor U13878 (N_13878,N_13034,N_13275);
or U13879 (N_13879,N_13038,N_13056);
or U13880 (N_13880,N_13139,N_13270);
nor U13881 (N_13881,N_13222,N_13172);
or U13882 (N_13882,N_13012,N_13137);
nand U13883 (N_13883,N_13317,N_13305);
nor U13884 (N_13884,N_13287,N_13116);
and U13885 (N_13885,N_13183,N_13277);
and U13886 (N_13886,N_13400,N_13285);
nor U13887 (N_13887,N_13235,N_13169);
and U13888 (N_13888,N_13460,N_13136);
xor U13889 (N_13889,N_13188,N_13291);
and U13890 (N_13890,N_13328,N_13066);
nand U13891 (N_13891,N_13279,N_13436);
xor U13892 (N_13892,N_13072,N_13302);
nor U13893 (N_13893,N_13236,N_13478);
nand U13894 (N_13894,N_13330,N_13201);
xor U13895 (N_13895,N_13446,N_13475);
xnor U13896 (N_13896,N_13390,N_13011);
or U13897 (N_13897,N_13284,N_13393);
nor U13898 (N_13898,N_13050,N_13228);
nand U13899 (N_13899,N_13224,N_13368);
and U13900 (N_13900,N_13074,N_13161);
xnor U13901 (N_13901,N_13433,N_13429);
and U13902 (N_13902,N_13014,N_13016);
nor U13903 (N_13903,N_13274,N_13168);
and U13904 (N_13904,N_13482,N_13162);
and U13905 (N_13905,N_13290,N_13103);
nor U13906 (N_13906,N_13347,N_13071);
nor U13907 (N_13907,N_13381,N_13003);
and U13908 (N_13908,N_13158,N_13197);
or U13909 (N_13909,N_13004,N_13226);
nand U13910 (N_13910,N_13145,N_13417);
nor U13911 (N_13911,N_13244,N_13297);
xnor U13912 (N_13912,N_13483,N_13248);
or U13913 (N_13913,N_13376,N_13433);
xnor U13914 (N_13914,N_13010,N_13141);
or U13915 (N_13915,N_13072,N_13373);
nand U13916 (N_13916,N_13254,N_13218);
nor U13917 (N_13917,N_13421,N_13144);
xnor U13918 (N_13918,N_13390,N_13181);
nand U13919 (N_13919,N_13382,N_13411);
and U13920 (N_13920,N_13458,N_13031);
or U13921 (N_13921,N_13143,N_13132);
and U13922 (N_13922,N_13285,N_13089);
nand U13923 (N_13923,N_13274,N_13400);
and U13924 (N_13924,N_13007,N_13073);
or U13925 (N_13925,N_13395,N_13185);
or U13926 (N_13926,N_13100,N_13282);
nand U13927 (N_13927,N_13026,N_13488);
xor U13928 (N_13928,N_13031,N_13401);
nand U13929 (N_13929,N_13355,N_13143);
xnor U13930 (N_13930,N_13267,N_13220);
xnor U13931 (N_13931,N_13226,N_13366);
nor U13932 (N_13932,N_13148,N_13289);
and U13933 (N_13933,N_13094,N_13420);
nor U13934 (N_13934,N_13021,N_13289);
nor U13935 (N_13935,N_13191,N_13106);
and U13936 (N_13936,N_13243,N_13301);
and U13937 (N_13937,N_13167,N_13493);
nor U13938 (N_13938,N_13256,N_13180);
and U13939 (N_13939,N_13024,N_13068);
or U13940 (N_13940,N_13372,N_13157);
xor U13941 (N_13941,N_13017,N_13442);
nand U13942 (N_13942,N_13350,N_13134);
xnor U13943 (N_13943,N_13124,N_13499);
or U13944 (N_13944,N_13361,N_13239);
nor U13945 (N_13945,N_13158,N_13414);
or U13946 (N_13946,N_13486,N_13390);
nand U13947 (N_13947,N_13038,N_13289);
nand U13948 (N_13948,N_13344,N_13162);
or U13949 (N_13949,N_13398,N_13471);
or U13950 (N_13950,N_13152,N_13496);
xor U13951 (N_13951,N_13245,N_13278);
and U13952 (N_13952,N_13183,N_13262);
and U13953 (N_13953,N_13089,N_13315);
or U13954 (N_13954,N_13333,N_13493);
nor U13955 (N_13955,N_13349,N_13133);
nand U13956 (N_13956,N_13011,N_13475);
and U13957 (N_13957,N_13296,N_13141);
nand U13958 (N_13958,N_13356,N_13422);
or U13959 (N_13959,N_13264,N_13489);
or U13960 (N_13960,N_13028,N_13431);
or U13961 (N_13961,N_13448,N_13244);
and U13962 (N_13962,N_13266,N_13226);
and U13963 (N_13963,N_13442,N_13141);
nor U13964 (N_13964,N_13291,N_13112);
xor U13965 (N_13965,N_13049,N_13074);
nor U13966 (N_13966,N_13206,N_13067);
and U13967 (N_13967,N_13458,N_13312);
and U13968 (N_13968,N_13265,N_13195);
nor U13969 (N_13969,N_13064,N_13189);
nor U13970 (N_13970,N_13474,N_13140);
nand U13971 (N_13971,N_13138,N_13041);
xnor U13972 (N_13972,N_13105,N_13122);
and U13973 (N_13973,N_13261,N_13226);
or U13974 (N_13974,N_13477,N_13322);
or U13975 (N_13975,N_13308,N_13278);
nand U13976 (N_13976,N_13471,N_13390);
nand U13977 (N_13977,N_13459,N_13476);
and U13978 (N_13978,N_13420,N_13090);
or U13979 (N_13979,N_13023,N_13185);
and U13980 (N_13980,N_13372,N_13368);
or U13981 (N_13981,N_13125,N_13010);
xnor U13982 (N_13982,N_13481,N_13017);
or U13983 (N_13983,N_13227,N_13133);
or U13984 (N_13984,N_13241,N_13485);
xor U13985 (N_13985,N_13176,N_13379);
nand U13986 (N_13986,N_13499,N_13245);
or U13987 (N_13987,N_13018,N_13394);
and U13988 (N_13988,N_13143,N_13282);
or U13989 (N_13989,N_13257,N_13415);
nor U13990 (N_13990,N_13278,N_13286);
and U13991 (N_13991,N_13301,N_13273);
nand U13992 (N_13992,N_13376,N_13316);
nand U13993 (N_13993,N_13305,N_13075);
or U13994 (N_13994,N_13433,N_13208);
nand U13995 (N_13995,N_13236,N_13461);
nor U13996 (N_13996,N_13074,N_13261);
nand U13997 (N_13997,N_13196,N_13310);
nor U13998 (N_13998,N_13130,N_13013);
xnor U13999 (N_13999,N_13368,N_13376);
and U14000 (N_14000,N_13534,N_13936);
nand U14001 (N_14001,N_13915,N_13700);
or U14002 (N_14002,N_13984,N_13814);
and U14003 (N_14003,N_13985,N_13543);
nand U14004 (N_14004,N_13580,N_13591);
and U14005 (N_14005,N_13917,N_13747);
nor U14006 (N_14006,N_13903,N_13940);
nand U14007 (N_14007,N_13756,N_13832);
nand U14008 (N_14008,N_13722,N_13744);
xor U14009 (N_14009,N_13567,N_13675);
nand U14010 (N_14010,N_13688,N_13759);
nand U14011 (N_14011,N_13930,N_13801);
xor U14012 (N_14012,N_13879,N_13853);
and U14013 (N_14013,N_13625,N_13515);
nand U14014 (N_14014,N_13926,N_13527);
nor U14015 (N_14015,N_13731,N_13523);
or U14016 (N_14016,N_13568,N_13566);
nand U14017 (N_14017,N_13957,N_13989);
and U14018 (N_14018,N_13648,N_13739);
nor U14019 (N_14019,N_13766,N_13774);
xnor U14020 (N_14020,N_13729,N_13737);
or U14021 (N_14021,N_13782,N_13871);
nor U14022 (N_14022,N_13861,N_13525);
nor U14023 (N_14023,N_13736,N_13696);
xnor U14024 (N_14024,N_13786,N_13891);
xor U14025 (N_14025,N_13843,N_13512);
nor U14026 (N_14026,N_13797,N_13862);
or U14027 (N_14027,N_13702,N_13829);
xnor U14028 (N_14028,N_13844,N_13845);
nand U14029 (N_14029,N_13539,N_13849);
nor U14030 (N_14030,N_13794,N_13790);
nor U14031 (N_14031,N_13995,N_13603);
nor U14032 (N_14032,N_13847,N_13518);
nand U14033 (N_14033,N_13890,N_13990);
nand U14034 (N_14034,N_13939,N_13927);
nor U14035 (N_14035,N_13994,N_13901);
and U14036 (N_14036,N_13654,N_13916);
xor U14037 (N_14037,N_13532,N_13511);
nand U14038 (N_14038,N_13595,N_13530);
xnor U14039 (N_14039,N_13502,N_13676);
or U14040 (N_14040,N_13909,N_13841);
and U14041 (N_14041,N_13979,N_13992);
xnor U14042 (N_14042,N_13577,N_13955);
or U14043 (N_14043,N_13682,N_13725);
nand U14044 (N_14044,N_13639,N_13818);
or U14045 (N_14045,N_13770,N_13937);
nand U14046 (N_14046,N_13520,N_13852);
xnor U14047 (N_14047,N_13694,N_13644);
xor U14048 (N_14048,N_13629,N_13711);
or U14049 (N_14049,N_13602,N_13635);
or U14050 (N_14050,N_13810,N_13627);
nor U14051 (N_14051,N_13870,N_13552);
xor U14052 (N_14052,N_13562,N_13953);
nand U14053 (N_14053,N_13628,N_13604);
or U14054 (N_14054,N_13811,N_13899);
or U14055 (N_14055,N_13524,N_13519);
and U14056 (N_14056,N_13689,N_13652);
nor U14057 (N_14057,N_13968,N_13948);
and U14058 (N_14058,N_13606,N_13695);
xnor U14059 (N_14059,N_13768,N_13560);
xor U14060 (N_14060,N_13618,N_13670);
nor U14061 (N_14061,N_13545,N_13834);
nand U14062 (N_14062,N_13872,N_13906);
and U14063 (N_14063,N_13723,N_13658);
nor U14064 (N_14064,N_13967,N_13503);
nor U14065 (N_14065,N_13724,N_13646);
or U14066 (N_14066,N_13703,N_13836);
nor U14067 (N_14067,N_13954,N_13765);
nand U14068 (N_14068,N_13971,N_13815);
nand U14069 (N_14069,N_13581,N_13505);
and U14070 (N_14070,N_13791,N_13544);
and U14071 (N_14071,N_13709,N_13900);
and U14072 (N_14072,N_13718,N_13687);
xor U14073 (N_14073,N_13809,N_13970);
nor U14074 (N_14074,N_13565,N_13526);
nor U14075 (N_14075,N_13943,N_13907);
nand U14076 (N_14076,N_13589,N_13986);
nor U14077 (N_14077,N_13828,N_13949);
nand U14078 (N_14078,N_13674,N_13691);
xnor U14079 (N_14079,N_13780,N_13745);
nor U14080 (N_14080,N_13800,N_13888);
xor U14081 (N_14081,N_13666,N_13905);
nor U14082 (N_14082,N_13886,N_13662);
nand U14083 (N_14083,N_13776,N_13594);
or U14084 (N_14084,N_13657,N_13787);
or U14085 (N_14085,N_13660,N_13698);
xnor U14086 (N_14086,N_13501,N_13650);
or U14087 (N_14087,N_13582,N_13740);
and U14088 (N_14088,N_13964,N_13704);
and U14089 (N_14089,N_13669,N_13798);
and U14090 (N_14090,N_13822,N_13713);
and U14091 (N_14091,N_13935,N_13751);
nor U14092 (N_14092,N_13858,N_13923);
and U14093 (N_14093,N_13997,N_13500);
and U14094 (N_14094,N_13509,N_13981);
xor U14095 (N_14095,N_13781,N_13732);
nand U14096 (N_14096,N_13912,N_13622);
and U14097 (N_14097,N_13777,N_13680);
and U14098 (N_14098,N_13920,N_13571);
or U14099 (N_14099,N_13902,N_13649);
and U14100 (N_14100,N_13656,N_13645);
nand U14101 (N_14101,N_13504,N_13588);
nand U14102 (N_14102,N_13621,N_13898);
or U14103 (N_14103,N_13869,N_13750);
xnor U14104 (N_14104,N_13510,N_13708);
nor U14105 (N_14105,N_13816,N_13758);
xor U14106 (N_14106,N_13956,N_13827);
nor U14107 (N_14107,N_13742,N_13804);
xor U14108 (N_14108,N_13941,N_13579);
nand U14109 (N_14109,N_13963,N_13638);
xor U14110 (N_14110,N_13878,N_13553);
nor U14111 (N_14111,N_13817,N_13730);
or U14112 (N_14112,N_13607,N_13641);
nor U14113 (N_14113,N_13664,N_13507);
xnor U14114 (N_14114,N_13640,N_13671);
nor U14115 (N_14115,N_13746,N_13880);
or U14116 (N_14116,N_13895,N_13554);
nand U14117 (N_14117,N_13548,N_13719);
and U14118 (N_14118,N_13881,N_13668);
nor U14119 (N_14119,N_13913,N_13788);
and U14120 (N_14120,N_13633,N_13616);
nor U14121 (N_14121,N_13529,N_13587);
or U14122 (N_14122,N_13617,N_13599);
nor U14123 (N_14123,N_13585,N_13726);
nand U14124 (N_14124,N_13556,N_13763);
nor U14125 (N_14125,N_13609,N_13772);
nand U14126 (N_14126,N_13896,N_13767);
xor U14127 (N_14127,N_13559,N_13743);
or U14128 (N_14128,N_13690,N_13842);
nand U14129 (N_14129,N_13848,N_13717);
and U14130 (N_14130,N_13821,N_13555);
nor U14131 (N_14131,N_13993,N_13813);
nor U14132 (N_14132,N_13535,N_13928);
nor U14133 (N_14133,N_13651,N_13933);
and U14134 (N_14134,N_13733,N_13569);
nor U14135 (N_14135,N_13864,N_13875);
or U14136 (N_14136,N_13793,N_13647);
nor U14137 (N_14137,N_13549,N_13681);
or U14138 (N_14138,N_13812,N_13974);
or U14139 (N_14139,N_13914,N_13803);
nor U14140 (N_14140,N_13988,N_13942);
xor U14141 (N_14141,N_13802,N_13752);
xor U14142 (N_14142,N_13659,N_13982);
nor U14143 (N_14143,N_13685,N_13672);
nor U14144 (N_14144,N_13998,N_13830);
or U14145 (N_14145,N_13973,N_13760);
nor U14146 (N_14146,N_13908,N_13710);
and U14147 (N_14147,N_13865,N_13643);
xnor U14148 (N_14148,N_13820,N_13558);
xnor U14149 (N_14149,N_13684,N_13761);
nand U14150 (N_14150,N_13897,N_13833);
nand U14151 (N_14151,N_13661,N_13508);
xor U14152 (N_14152,N_13838,N_13976);
or U14153 (N_14153,N_13944,N_13721);
xnor U14154 (N_14154,N_13596,N_13945);
and U14155 (N_14155,N_13655,N_13614);
xor U14156 (N_14156,N_13679,N_13550);
xor U14157 (N_14157,N_13826,N_13665);
nand U14158 (N_14158,N_13792,N_13572);
or U14159 (N_14159,N_13855,N_13540);
nand U14160 (N_14160,N_13699,N_13578);
nand U14161 (N_14161,N_13958,N_13769);
and U14162 (N_14162,N_13678,N_13859);
xnor U14163 (N_14163,N_13775,N_13686);
or U14164 (N_14164,N_13590,N_13860);
nor U14165 (N_14165,N_13626,N_13934);
xnor U14166 (N_14166,N_13608,N_13546);
or U14167 (N_14167,N_13796,N_13653);
or U14168 (N_14168,N_13570,N_13734);
or U14169 (N_14169,N_13831,N_13806);
or U14170 (N_14170,N_13789,N_13991);
and U14171 (N_14171,N_13877,N_13701);
xor U14172 (N_14172,N_13592,N_13846);
nor U14173 (N_14173,N_13922,N_13716);
nand U14174 (N_14174,N_13521,N_13887);
and U14175 (N_14175,N_13961,N_13637);
nand U14176 (N_14176,N_13612,N_13921);
or U14177 (N_14177,N_13754,N_13522);
nand U14178 (N_14178,N_13966,N_13683);
nor U14179 (N_14179,N_13598,N_13863);
or U14180 (N_14180,N_13919,N_13642);
or U14181 (N_14181,N_13514,N_13741);
nand U14182 (N_14182,N_13835,N_13778);
and U14183 (N_14183,N_13692,N_13996);
nand U14184 (N_14184,N_13611,N_13575);
nand U14185 (N_14185,N_13506,N_13677);
and U14186 (N_14186,N_13856,N_13975);
or U14187 (N_14187,N_13904,N_13715);
xnor U14188 (N_14188,N_13840,N_13632);
or U14189 (N_14189,N_13925,N_13946);
or U14190 (N_14190,N_13727,N_13938);
and U14191 (N_14191,N_13972,N_13805);
nor U14192 (N_14192,N_13728,N_13712);
and U14193 (N_14193,N_13753,N_13574);
xnor U14194 (N_14194,N_13932,N_13876);
xnor U14195 (N_14195,N_13673,N_13551);
xor U14196 (N_14196,N_13837,N_13962);
nor U14197 (N_14197,N_13541,N_13613);
nand U14198 (N_14198,N_13882,N_13951);
and U14199 (N_14199,N_13952,N_13885);
nand U14200 (N_14200,N_13576,N_13911);
nor U14201 (N_14201,N_13987,N_13857);
nor U14202 (N_14202,N_13630,N_13610);
nor U14203 (N_14203,N_13960,N_13850);
nor U14204 (N_14204,N_13531,N_13573);
or U14205 (N_14205,N_13563,N_13892);
nor U14206 (N_14206,N_13714,N_13980);
and U14207 (N_14207,N_13823,N_13873);
or U14208 (N_14208,N_13866,N_13623);
or U14209 (N_14209,N_13605,N_13593);
nor U14210 (N_14210,N_13738,N_13583);
nand U14211 (N_14211,N_13773,N_13516);
nand U14212 (N_14212,N_13839,N_13693);
and U14213 (N_14213,N_13884,N_13667);
xnor U14214 (N_14214,N_13918,N_13874);
or U14215 (N_14215,N_13924,N_13536);
or U14216 (N_14216,N_13983,N_13619);
nand U14217 (N_14217,N_13624,N_13779);
xor U14218 (N_14218,N_13634,N_13620);
and U14219 (N_14219,N_13969,N_13513);
or U14220 (N_14220,N_13597,N_13615);
nand U14221 (N_14221,N_13584,N_13557);
and U14222 (N_14222,N_13929,N_13947);
and U14223 (N_14223,N_13783,N_13720);
nor U14224 (N_14224,N_13528,N_13824);
and U14225 (N_14225,N_13600,N_13819);
nor U14226 (N_14226,N_13631,N_13851);
nor U14227 (N_14227,N_13663,N_13762);
xnor U14228 (N_14228,N_13950,N_13517);
nor U14229 (N_14229,N_13735,N_13799);
xnor U14230 (N_14230,N_13764,N_13749);
xor U14231 (N_14231,N_13785,N_13978);
nand U14232 (N_14232,N_13586,N_13795);
or U14233 (N_14233,N_13883,N_13867);
or U14234 (N_14234,N_13807,N_13755);
xnor U14235 (N_14235,N_13538,N_13697);
and U14236 (N_14236,N_13893,N_13910);
nor U14237 (N_14237,N_13748,N_13757);
nand U14238 (N_14238,N_13977,N_13999);
nor U14239 (N_14239,N_13808,N_13965);
nor U14240 (N_14240,N_13706,N_13601);
nand U14241 (N_14241,N_13894,N_13564);
xor U14242 (N_14242,N_13561,N_13784);
xnor U14243 (N_14243,N_13542,N_13854);
xor U14244 (N_14244,N_13825,N_13771);
and U14245 (N_14245,N_13707,N_13705);
or U14246 (N_14246,N_13547,N_13533);
and U14247 (N_14247,N_13636,N_13959);
or U14248 (N_14248,N_13889,N_13931);
nor U14249 (N_14249,N_13537,N_13868);
or U14250 (N_14250,N_13878,N_13910);
nor U14251 (N_14251,N_13968,N_13865);
nor U14252 (N_14252,N_13659,N_13782);
nand U14253 (N_14253,N_13588,N_13532);
and U14254 (N_14254,N_13663,N_13727);
and U14255 (N_14255,N_13868,N_13948);
xor U14256 (N_14256,N_13751,N_13817);
nor U14257 (N_14257,N_13767,N_13821);
or U14258 (N_14258,N_13708,N_13796);
nor U14259 (N_14259,N_13612,N_13776);
or U14260 (N_14260,N_13599,N_13984);
nor U14261 (N_14261,N_13893,N_13699);
and U14262 (N_14262,N_13524,N_13877);
nand U14263 (N_14263,N_13821,N_13786);
and U14264 (N_14264,N_13721,N_13685);
and U14265 (N_14265,N_13980,N_13838);
or U14266 (N_14266,N_13929,N_13844);
xor U14267 (N_14267,N_13659,N_13627);
xnor U14268 (N_14268,N_13686,N_13859);
nand U14269 (N_14269,N_13867,N_13527);
and U14270 (N_14270,N_13992,N_13931);
nand U14271 (N_14271,N_13547,N_13777);
or U14272 (N_14272,N_13642,N_13654);
xnor U14273 (N_14273,N_13977,N_13972);
nor U14274 (N_14274,N_13785,N_13527);
xnor U14275 (N_14275,N_13525,N_13825);
xnor U14276 (N_14276,N_13672,N_13828);
nand U14277 (N_14277,N_13969,N_13834);
nand U14278 (N_14278,N_13518,N_13567);
or U14279 (N_14279,N_13779,N_13739);
and U14280 (N_14280,N_13835,N_13543);
xnor U14281 (N_14281,N_13768,N_13570);
and U14282 (N_14282,N_13855,N_13979);
nand U14283 (N_14283,N_13983,N_13999);
nand U14284 (N_14284,N_13856,N_13530);
xor U14285 (N_14285,N_13926,N_13865);
or U14286 (N_14286,N_13768,N_13989);
or U14287 (N_14287,N_13846,N_13787);
xor U14288 (N_14288,N_13514,N_13863);
or U14289 (N_14289,N_13787,N_13638);
xnor U14290 (N_14290,N_13718,N_13701);
or U14291 (N_14291,N_13591,N_13747);
nand U14292 (N_14292,N_13906,N_13543);
nand U14293 (N_14293,N_13941,N_13513);
nor U14294 (N_14294,N_13726,N_13753);
xnor U14295 (N_14295,N_13563,N_13635);
nand U14296 (N_14296,N_13594,N_13623);
or U14297 (N_14297,N_13832,N_13931);
xnor U14298 (N_14298,N_13909,N_13616);
xnor U14299 (N_14299,N_13686,N_13547);
nand U14300 (N_14300,N_13514,N_13977);
nor U14301 (N_14301,N_13964,N_13725);
xor U14302 (N_14302,N_13952,N_13751);
and U14303 (N_14303,N_13629,N_13544);
xor U14304 (N_14304,N_13951,N_13905);
and U14305 (N_14305,N_13559,N_13545);
or U14306 (N_14306,N_13555,N_13745);
nand U14307 (N_14307,N_13559,N_13983);
or U14308 (N_14308,N_13985,N_13885);
and U14309 (N_14309,N_13636,N_13564);
nor U14310 (N_14310,N_13636,N_13722);
or U14311 (N_14311,N_13569,N_13833);
xor U14312 (N_14312,N_13992,N_13675);
xor U14313 (N_14313,N_13633,N_13525);
nor U14314 (N_14314,N_13923,N_13904);
or U14315 (N_14315,N_13653,N_13836);
xor U14316 (N_14316,N_13819,N_13583);
and U14317 (N_14317,N_13973,N_13806);
nor U14318 (N_14318,N_13860,N_13770);
xor U14319 (N_14319,N_13735,N_13844);
or U14320 (N_14320,N_13787,N_13823);
and U14321 (N_14321,N_13865,N_13704);
or U14322 (N_14322,N_13682,N_13644);
xnor U14323 (N_14323,N_13733,N_13581);
xor U14324 (N_14324,N_13864,N_13599);
xnor U14325 (N_14325,N_13578,N_13755);
or U14326 (N_14326,N_13764,N_13914);
nand U14327 (N_14327,N_13947,N_13976);
xor U14328 (N_14328,N_13987,N_13933);
and U14329 (N_14329,N_13831,N_13529);
xor U14330 (N_14330,N_13929,N_13691);
and U14331 (N_14331,N_13572,N_13763);
and U14332 (N_14332,N_13959,N_13899);
or U14333 (N_14333,N_13935,N_13923);
and U14334 (N_14334,N_13529,N_13702);
and U14335 (N_14335,N_13553,N_13707);
and U14336 (N_14336,N_13519,N_13702);
or U14337 (N_14337,N_13867,N_13891);
nor U14338 (N_14338,N_13965,N_13856);
and U14339 (N_14339,N_13544,N_13885);
nor U14340 (N_14340,N_13569,N_13868);
and U14341 (N_14341,N_13718,N_13954);
or U14342 (N_14342,N_13968,N_13989);
nor U14343 (N_14343,N_13831,N_13837);
nor U14344 (N_14344,N_13667,N_13504);
or U14345 (N_14345,N_13724,N_13714);
and U14346 (N_14346,N_13610,N_13960);
xnor U14347 (N_14347,N_13608,N_13901);
nand U14348 (N_14348,N_13528,N_13859);
nor U14349 (N_14349,N_13547,N_13975);
or U14350 (N_14350,N_13540,N_13861);
nor U14351 (N_14351,N_13514,N_13805);
or U14352 (N_14352,N_13827,N_13529);
or U14353 (N_14353,N_13532,N_13899);
nand U14354 (N_14354,N_13999,N_13771);
and U14355 (N_14355,N_13930,N_13942);
nor U14356 (N_14356,N_13767,N_13781);
xnor U14357 (N_14357,N_13519,N_13505);
nand U14358 (N_14358,N_13544,N_13525);
nand U14359 (N_14359,N_13873,N_13889);
nor U14360 (N_14360,N_13600,N_13698);
and U14361 (N_14361,N_13555,N_13879);
nand U14362 (N_14362,N_13588,N_13694);
or U14363 (N_14363,N_13581,N_13676);
nand U14364 (N_14364,N_13831,N_13593);
nand U14365 (N_14365,N_13746,N_13887);
xnor U14366 (N_14366,N_13866,N_13993);
nor U14367 (N_14367,N_13565,N_13890);
nand U14368 (N_14368,N_13685,N_13944);
and U14369 (N_14369,N_13541,N_13829);
nand U14370 (N_14370,N_13863,N_13540);
nand U14371 (N_14371,N_13956,N_13814);
nand U14372 (N_14372,N_13579,N_13852);
xor U14373 (N_14373,N_13609,N_13532);
nand U14374 (N_14374,N_13919,N_13708);
nand U14375 (N_14375,N_13520,N_13997);
nor U14376 (N_14376,N_13887,N_13714);
and U14377 (N_14377,N_13776,N_13915);
or U14378 (N_14378,N_13596,N_13892);
or U14379 (N_14379,N_13740,N_13946);
and U14380 (N_14380,N_13790,N_13779);
or U14381 (N_14381,N_13754,N_13739);
xnor U14382 (N_14382,N_13804,N_13799);
nand U14383 (N_14383,N_13869,N_13981);
nor U14384 (N_14384,N_13846,N_13721);
or U14385 (N_14385,N_13646,N_13947);
or U14386 (N_14386,N_13840,N_13828);
or U14387 (N_14387,N_13520,N_13752);
nand U14388 (N_14388,N_13502,N_13960);
xnor U14389 (N_14389,N_13892,N_13877);
and U14390 (N_14390,N_13538,N_13622);
nor U14391 (N_14391,N_13580,N_13571);
nand U14392 (N_14392,N_13783,N_13799);
or U14393 (N_14393,N_13952,N_13593);
nand U14394 (N_14394,N_13501,N_13930);
or U14395 (N_14395,N_13791,N_13520);
or U14396 (N_14396,N_13595,N_13913);
nor U14397 (N_14397,N_13711,N_13544);
nor U14398 (N_14398,N_13754,N_13747);
nand U14399 (N_14399,N_13831,N_13629);
nand U14400 (N_14400,N_13727,N_13994);
nor U14401 (N_14401,N_13649,N_13570);
nor U14402 (N_14402,N_13666,N_13654);
nand U14403 (N_14403,N_13995,N_13746);
or U14404 (N_14404,N_13667,N_13983);
nand U14405 (N_14405,N_13737,N_13629);
nor U14406 (N_14406,N_13978,N_13740);
nand U14407 (N_14407,N_13913,N_13626);
or U14408 (N_14408,N_13865,N_13579);
or U14409 (N_14409,N_13716,N_13635);
nand U14410 (N_14410,N_13542,N_13767);
or U14411 (N_14411,N_13865,N_13504);
and U14412 (N_14412,N_13770,N_13721);
nand U14413 (N_14413,N_13588,N_13601);
nand U14414 (N_14414,N_13884,N_13904);
nand U14415 (N_14415,N_13616,N_13906);
or U14416 (N_14416,N_13633,N_13961);
xnor U14417 (N_14417,N_13803,N_13610);
and U14418 (N_14418,N_13889,N_13677);
nand U14419 (N_14419,N_13700,N_13944);
xnor U14420 (N_14420,N_13985,N_13692);
nand U14421 (N_14421,N_13651,N_13895);
and U14422 (N_14422,N_13978,N_13852);
nor U14423 (N_14423,N_13744,N_13813);
and U14424 (N_14424,N_13659,N_13893);
nor U14425 (N_14425,N_13796,N_13721);
or U14426 (N_14426,N_13649,N_13808);
and U14427 (N_14427,N_13664,N_13866);
and U14428 (N_14428,N_13947,N_13737);
nor U14429 (N_14429,N_13972,N_13692);
and U14430 (N_14430,N_13959,N_13787);
and U14431 (N_14431,N_13528,N_13884);
or U14432 (N_14432,N_13548,N_13542);
nor U14433 (N_14433,N_13500,N_13519);
nand U14434 (N_14434,N_13667,N_13812);
and U14435 (N_14435,N_13741,N_13944);
xor U14436 (N_14436,N_13553,N_13770);
nand U14437 (N_14437,N_13746,N_13610);
or U14438 (N_14438,N_13725,N_13567);
or U14439 (N_14439,N_13871,N_13868);
nand U14440 (N_14440,N_13678,N_13524);
and U14441 (N_14441,N_13686,N_13872);
nand U14442 (N_14442,N_13533,N_13684);
and U14443 (N_14443,N_13755,N_13738);
nand U14444 (N_14444,N_13923,N_13831);
and U14445 (N_14445,N_13597,N_13756);
nand U14446 (N_14446,N_13808,N_13962);
nand U14447 (N_14447,N_13598,N_13802);
or U14448 (N_14448,N_13661,N_13620);
and U14449 (N_14449,N_13844,N_13988);
xnor U14450 (N_14450,N_13638,N_13864);
and U14451 (N_14451,N_13663,N_13860);
or U14452 (N_14452,N_13548,N_13645);
or U14453 (N_14453,N_13613,N_13903);
nor U14454 (N_14454,N_13550,N_13625);
nand U14455 (N_14455,N_13868,N_13623);
or U14456 (N_14456,N_13702,N_13628);
nand U14457 (N_14457,N_13736,N_13524);
and U14458 (N_14458,N_13925,N_13929);
or U14459 (N_14459,N_13948,N_13599);
xor U14460 (N_14460,N_13590,N_13538);
xor U14461 (N_14461,N_13727,N_13660);
nor U14462 (N_14462,N_13621,N_13516);
and U14463 (N_14463,N_13793,N_13932);
xor U14464 (N_14464,N_13722,N_13819);
nand U14465 (N_14465,N_13579,N_13946);
or U14466 (N_14466,N_13713,N_13792);
nand U14467 (N_14467,N_13793,N_13965);
nor U14468 (N_14468,N_13985,N_13829);
and U14469 (N_14469,N_13558,N_13994);
and U14470 (N_14470,N_13966,N_13997);
or U14471 (N_14471,N_13783,N_13530);
or U14472 (N_14472,N_13880,N_13945);
xor U14473 (N_14473,N_13980,N_13697);
nor U14474 (N_14474,N_13732,N_13710);
xor U14475 (N_14475,N_13767,N_13527);
and U14476 (N_14476,N_13849,N_13619);
xnor U14477 (N_14477,N_13712,N_13590);
and U14478 (N_14478,N_13603,N_13985);
nand U14479 (N_14479,N_13808,N_13655);
and U14480 (N_14480,N_13828,N_13816);
or U14481 (N_14481,N_13984,N_13652);
xnor U14482 (N_14482,N_13949,N_13948);
or U14483 (N_14483,N_13647,N_13645);
nand U14484 (N_14484,N_13657,N_13718);
or U14485 (N_14485,N_13754,N_13604);
xnor U14486 (N_14486,N_13809,N_13742);
xnor U14487 (N_14487,N_13793,N_13892);
xor U14488 (N_14488,N_13935,N_13679);
nand U14489 (N_14489,N_13878,N_13754);
or U14490 (N_14490,N_13620,N_13814);
xnor U14491 (N_14491,N_13959,N_13854);
or U14492 (N_14492,N_13783,N_13762);
xnor U14493 (N_14493,N_13938,N_13921);
xnor U14494 (N_14494,N_13780,N_13526);
or U14495 (N_14495,N_13810,N_13733);
and U14496 (N_14496,N_13924,N_13985);
xnor U14497 (N_14497,N_13760,N_13748);
nor U14498 (N_14498,N_13663,N_13957);
nor U14499 (N_14499,N_13859,N_13786);
nor U14500 (N_14500,N_14088,N_14321);
nand U14501 (N_14501,N_14282,N_14498);
nor U14502 (N_14502,N_14329,N_14405);
nand U14503 (N_14503,N_14146,N_14341);
nand U14504 (N_14504,N_14445,N_14204);
or U14505 (N_14505,N_14170,N_14112);
and U14506 (N_14506,N_14378,N_14233);
nor U14507 (N_14507,N_14150,N_14049);
nor U14508 (N_14508,N_14413,N_14179);
nor U14509 (N_14509,N_14120,N_14215);
nand U14510 (N_14510,N_14254,N_14468);
nor U14511 (N_14511,N_14460,N_14349);
and U14512 (N_14512,N_14289,N_14030);
nand U14513 (N_14513,N_14382,N_14486);
and U14514 (N_14514,N_14429,N_14190);
or U14515 (N_14515,N_14350,N_14453);
nor U14516 (N_14516,N_14199,N_14247);
xnor U14517 (N_14517,N_14305,N_14416);
or U14518 (N_14518,N_14175,N_14301);
xor U14519 (N_14519,N_14411,N_14041);
and U14520 (N_14520,N_14499,N_14298);
xor U14521 (N_14521,N_14184,N_14352);
nor U14522 (N_14522,N_14493,N_14180);
and U14523 (N_14523,N_14492,N_14219);
nand U14524 (N_14524,N_14217,N_14427);
or U14525 (N_14525,N_14372,N_14358);
and U14526 (N_14526,N_14220,N_14001);
nand U14527 (N_14527,N_14064,N_14391);
and U14528 (N_14528,N_14011,N_14343);
or U14529 (N_14529,N_14024,N_14087);
xnor U14530 (N_14530,N_14478,N_14265);
nand U14531 (N_14531,N_14497,N_14419);
nor U14532 (N_14532,N_14037,N_14467);
nor U14533 (N_14533,N_14465,N_14194);
xnor U14534 (N_14534,N_14353,N_14153);
nand U14535 (N_14535,N_14266,N_14365);
nand U14536 (N_14536,N_14481,N_14241);
xnor U14537 (N_14537,N_14235,N_14161);
xnor U14538 (N_14538,N_14267,N_14008);
nand U14539 (N_14539,N_14268,N_14483);
or U14540 (N_14540,N_14263,N_14007);
nand U14541 (N_14541,N_14073,N_14316);
or U14542 (N_14542,N_14090,N_14489);
nor U14543 (N_14543,N_14068,N_14178);
nand U14544 (N_14544,N_14314,N_14361);
nor U14545 (N_14545,N_14078,N_14402);
and U14546 (N_14546,N_14061,N_14388);
xor U14547 (N_14547,N_14389,N_14224);
or U14548 (N_14548,N_14027,N_14035);
xnor U14549 (N_14549,N_14136,N_14065);
xnor U14550 (N_14550,N_14397,N_14264);
and U14551 (N_14551,N_14396,N_14022);
nor U14552 (N_14552,N_14026,N_14306);
and U14553 (N_14553,N_14177,N_14356);
and U14554 (N_14554,N_14086,N_14166);
and U14555 (N_14555,N_14318,N_14395);
or U14556 (N_14556,N_14244,N_14206);
nor U14557 (N_14557,N_14439,N_14278);
nand U14558 (N_14558,N_14374,N_14295);
and U14559 (N_14559,N_14428,N_14484);
or U14560 (N_14560,N_14012,N_14139);
xnor U14561 (N_14561,N_14440,N_14345);
or U14562 (N_14562,N_14257,N_14050);
nor U14563 (N_14563,N_14021,N_14100);
or U14564 (N_14564,N_14213,N_14149);
nor U14565 (N_14565,N_14259,N_14123);
or U14566 (N_14566,N_14317,N_14095);
xor U14567 (N_14567,N_14029,N_14243);
xor U14568 (N_14568,N_14121,N_14044);
nor U14569 (N_14569,N_14183,N_14414);
nor U14570 (N_14570,N_14127,N_14294);
nor U14571 (N_14571,N_14009,N_14325);
or U14572 (N_14572,N_14162,N_14193);
nand U14573 (N_14573,N_14451,N_14403);
nand U14574 (N_14574,N_14063,N_14198);
nand U14575 (N_14575,N_14040,N_14415);
xor U14576 (N_14576,N_14205,N_14225);
and U14577 (N_14577,N_14043,N_14300);
nand U14578 (N_14578,N_14141,N_14174);
and U14579 (N_14579,N_14185,N_14071);
nand U14580 (N_14580,N_14010,N_14116);
and U14581 (N_14581,N_14494,N_14444);
and U14582 (N_14582,N_14412,N_14135);
or U14583 (N_14583,N_14222,N_14148);
xor U14584 (N_14584,N_14031,N_14046);
nand U14585 (N_14585,N_14421,N_14401);
or U14586 (N_14586,N_14272,N_14096);
or U14587 (N_14587,N_14344,N_14239);
or U14588 (N_14588,N_14383,N_14058);
or U14589 (N_14589,N_14076,N_14209);
nor U14590 (N_14590,N_14385,N_14079);
and U14591 (N_14591,N_14060,N_14370);
nand U14592 (N_14592,N_14056,N_14191);
nand U14593 (N_14593,N_14053,N_14496);
or U14594 (N_14594,N_14407,N_14384);
and U14595 (N_14595,N_14309,N_14433);
nor U14596 (N_14596,N_14052,N_14042);
nor U14597 (N_14597,N_14034,N_14140);
or U14598 (N_14598,N_14393,N_14474);
nor U14599 (N_14599,N_14200,N_14347);
xor U14600 (N_14600,N_14181,N_14229);
nand U14601 (N_14601,N_14152,N_14125);
xor U14602 (N_14602,N_14094,N_14255);
nand U14603 (N_14603,N_14400,N_14117);
or U14604 (N_14604,N_14147,N_14057);
or U14605 (N_14605,N_14367,N_14270);
nand U14606 (N_14606,N_14342,N_14381);
and U14607 (N_14607,N_14236,N_14286);
or U14608 (N_14608,N_14473,N_14275);
nor U14609 (N_14609,N_14288,N_14080);
xnor U14610 (N_14610,N_14338,N_14277);
or U14611 (N_14611,N_14323,N_14015);
nand U14612 (N_14612,N_14490,N_14249);
or U14613 (N_14613,N_14067,N_14107);
nor U14614 (N_14614,N_14482,N_14203);
xor U14615 (N_14615,N_14488,N_14406);
or U14616 (N_14616,N_14276,N_14299);
and U14617 (N_14617,N_14122,N_14134);
nand U14618 (N_14618,N_14328,N_14327);
and U14619 (N_14619,N_14274,N_14126);
nand U14620 (N_14620,N_14452,N_14032);
and U14621 (N_14621,N_14104,N_14069);
xor U14622 (N_14622,N_14210,N_14144);
and U14623 (N_14623,N_14438,N_14005);
and U14624 (N_14624,N_14446,N_14285);
xor U14625 (N_14625,N_14366,N_14099);
or U14626 (N_14626,N_14074,N_14038);
or U14627 (N_14627,N_14431,N_14477);
or U14628 (N_14628,N_14283,N_14133);
nor U14629 (N_14629,N_14485,N_14387);
nor U14630 (N_14630,N_14129,N_14377);
and U14631 (N_14631,N_14157,N_14487);
nor U14632 (N_14632,N_14240,N_14311);
xor U14633 (N_14633,N_14420,N_14196);
or U14634 (N_14634,N_14441,N_14297);
nor U14635 (N_14635,N_14113,N_14158);
nor U14636 (N_14636,N_14048,N_14333);
and U14637 (N_14637,N_14322,N_14047);
and U14638 (N_14638,N_14337,N_14077);
nand U14639 (N_14639,N_14168,N_14340);
and U14640 (N_14640,N_14223,N_14319);
nand U14641 (N_14641,N_14256,N_14472);
xor U14642 (N_14642,N_14084,N_14106);
nor U14643 (N_14643,N_14192,N_14293);
xor U14644 (N_14644,N_14025,N_14410);
nor U14645 (N_14645,N_14459,N_14287);
xor U14646 (N_14646,N_14167,N_14218);
nand U14647 (N_14647,N_14449,N_14252);
or U14648 (N_14648,N_14368,N_14138);
nor U14649 (N_14649,N_14188,N_14262);
and U14650 (N_14650,N_14348,N_14145);
nand U14651 (N_14651,N_14160,N_14399);
xor U14652 (N_14652,N_14462,N_14111);
nand U14653 (N_14653,N_14102,N_14437);
nor U14654 (N_14654,N_14118,N_14115);
xnor U14655 (N_14655,N_14376,N_14232);
xor U14656 (N_14656,N_14119,N_14004);
nor U14657 (N_14657,N_14404,N_14002);
nor U14658 (N_14658,N_14189,N_14461);
nor U14659 (N_14659,N_14163,N_14284);
xnor U14660 (N_14660,N_14207,N_14124);
nand U14661 (N_14661,N_14466,N_14142);
nand U14662 (N_14662,N_14083,N_14426);
nor U14663 (N_14663,N_14470,N_14226);
nand U14664 (N_14664,N_14435,N_14332);
xor U14665 (N_14665,N_14003,N_14258);
or U14666 (N_14666,N_14075,N_14330);
or U14667 (N_14667,N_14172,N_14154);
nor U14668 (N_14668,N_14335,N_14130);
nand U14669 (N_14669,N_14023,N_14491);
xor U14670 (N_14670,N_14458,N_14055);
nand U14671 (N_14671,N_14221,N_14230);
nor U14672 (N_14672,N_14182,N_14019);
or U14673 (N_14673,N_14132,N_14308);
and U14674 (N_14674,N_14363,N_14418);
nand U14675 (N_14675,N_14089,N_14369);
and U14676 (N_14676,N_14279,N_14237);
and U14677 (N_14677,N_14454,N_14228);
or U14678 (N_14678,N_14434,N_14197);
nand U14679 (N_14679,N_14371,N_14131);
or U14680 (N_14680,N_14390,N_14072);
and U14681 (N_14681,N_14351,N_14151);
xor U14682 (N_14682,N_14422,N_14059);
and U14683 (N_14683,N_14290,N_14245);
or U14684 (N_14684,N_14291,N_14108);
xnor U14685 (N_14685,N_14375,N_14281);
and U14686 (N_14686,N_14475,N_14098);
or U14687 (N_14687,N_14271,N_14436);
and U14688 (N_14688,N_14360,N_14036);
nor U14689 (N_14689,N_14304,N_14457);
and U14690 (N_14690,N_14326,N_14469);
or U14691 (N_14691,N_14331,N_14234);
nor U14692 (N_14692,N_14424,N_14250);
xor U14693 (N_14693,N_14364,N_14355);
xnor U14694 (N_14694,N_14109,N_14039);
or U14695 (N_14695,N_14156,N_14315);
or U14696 (N_14696,N_14303,N_14137);
and U14697 (N_14697,N_14346,N_14379);
nor U14698 (N_14698,N_14028,N_14373);
nand U14699 (N_14699,N_14091,N_14081);
or U14700 (N_14700,N_14165,N_14013);
nand U14701 (N_14701,N_14092,N_14296);
nor U14702 (N_14702,N_14164,N_14082);
nor U14703 (N_14703,N_14159,N_14105);
or U14704 (N_14704,N_14006,N_14334);
or U14705 (N_14705,N_14128,N_14017);
nand U14706 (N_14706,N_14054,N_14292);
xnor U14707 (N_14707,N_14320,N_14430);
and U14708 (N_14708,N_14432,N_14066);
nand U14709 (N_14709,N_14216,N_14463);
nand U14710 (N_14710,N_14456,N_14339);
nor U14711 (N_14711,N_14479,N_14173);
and U14712 (N_14712,N_14307,N_14425);
and U14713 (N_14713,N_14409,N_14070);
and U14714 (N_14714,N_14423,N_14171);
nand U14715 (N_14715,N_14464,N_14242);
or U14716 (N_14716,N_14260,N_14033);
nor U14717 (N_14717,N_14211,N_14357);
nor U14718 (N_14718,N_14359,N_14020);
or U14719 (N_14719,N_14261,N_14380);
xor U14720 (N_14720,N_14212,N_14093);
or U14721 (N_14721,N_14273,N_14269);
and U14722 (N_14722,N_14302,N_14186);
nor U14723 (N_14723,N_14443,N_14103);
nand U14724 (N_14724,N_14085,N_14448);
and U14725 (N_14725,N_14354,N_14114);
nor U14726 (N_14726,N_14392,N_14480);
or U14727 (N_14727,N_14238,N_14045);
and U14728 (N_14728,N_14442,N_14495);
nand U14729 (N_14729,N_14476,N_14143);
or U14730 (N_14730,N_14208,N_14417);
xnor U14731 (N_14731,N_14214,N_14408);
xor U14732 (N_14732,N_14201,N_14231);
nand U14733 (N_14733,N_14176,N_14324);
nor U14734 (N_14734,N_14101,N_14195);
nand U14735 (N_14735,N_14398,N_14280);
or U14736 (N_14736,N_14394,N_14248);
xor U14737 (N_14737,N_14227,N_14312);
or U14738 (N_14738,N_14336,N_14016);
and U14739 (N_14739,N_14097,N_14251);
xor U14740 (N_14740,N_14471,N_14062);
nor U14741 (N_14741,N_14253,N_14000);
or U14742 (N_14742,N_14386,N_14313);
xnor U14743 (N_14743,N_14455,N_14450);
nor U14744 (N_14744,N_14310,N_14051);
nor U14745 (N_14745,N_14014,N_14169);
and U14746 (N_14746,N_14246,N_14155);
or U14747 (N_14747,N_14362,N_14202);
xor U14748 (N_14748,N_14018,N_14187);
xor U14749 (N_14749,N_14447,N_14110);
xor U14750 (N_14750,N_14439,N_14012);
nand U14751 (N_14751,N_14161,N_14130);
xnor U14752 (N_14752,N_14208,N_14364);
nor U14753 (N_14753,N_14407,N_14005);
nand U14754 (N_14754,N_14259,N_14485);
or U14755 (N_14755,N_14469,N_14484);
nor U14756 (N_14756,N_14332,N_14285);
nor U14757 (N_14757,N_14328,N_14425);
or U14758 (N_14758,N_14262,N_14090);
xor U14759 (N_14759,N_14143,N_14400);
nor U14760 (N_14760,N_14216,N_14002);
or U14761 (N_14761,N_14384,N_14284);
nor U14762 (N_14762,N_14105,N_14021);
xnor U14763 (N_14763,N_14272,N_14256);
or U14764 (N_14764,N_14454,N_14032);
nor U14765 (N_14765,N_14072,N_14440);
nand U14766 (N_14766,N_14142,N_14330);
nor U14767 (N_14767,N_14268,N_14074);
nand U14768 (N_14768,N_14308,N_14476);
xor U14769 (N_14769,N_14498,N_14245);
xnor U14770 (N_14770,N_14124,N_14208);
or U14771 (N_14771,N_14404,N_14048);
and U14772 (N_14772,N_14239,N_14438);
or U14773 (N_14773,N_14448,N_14351);
nor U14774 (N_14774,N_14490,N_14271);
nor U14775 (N_14775,N_14006,N_14320);
or U14776 (N_14776,N_14437,N_14235);
nand U14777 (N_14777,N_14443,N_14417);
xnor U14778 (N_14778,N_14359,N_14299);
xnor U14779 (N_14779,N_14363,N_14010);
nor U14780 (N_14780,N_14435,N_14041);
nand U14781 (N_14781,N_14459,N_14108);
nand U14782 (N_14782,N_14130,N_14309);
and U14783 (N_14783,N_14015,N_14204);
and U14784 (N_14784,N_14039,N_14343);
nand U14785 (N_14785,N_14070,N_14300);
nand U14786 (N_14786,N_14410,N_14443);
or U14787 (N_14787,N_14368,N_14074);
nor U14788 (N_14788,N_14088,N_14478);
nand U14789 (N_14789,N_14333,N_14246);
and U14790 (N_14790,N_14166,N_14171);
nor U14791 (N_14791,N_14318,N_14058);
or U14792 (N_14792,N_14104,N_14243);
and U14793 (N_14793,N_14226,N_14183);
and U14794 (N_14794,N_14269,N_14000);
nand U14795 (N_14795,N_14120,N_14462);
xnor U14796 (N_14796,N_14424,N_14164);
and U14797 (N_14797,N_14429,N_14031);
and U14798 (N_14798,N_14458,N_14172);
nor U14799 (N_14799,N_14000,N_14474);
xor U14800 (N_14800,N_14480,N_14133);
nand U14801 (N_14801,N_14103,N_14322);
or U14802 (N_14802,N_14181,N_14016);
or U14803 (N_14803,N_14395,N_14407);
nand U14804 (N_14804,N_14021,N_14043);
nand U14805 (N_14805,N_14167,N_14031);
nor U14806 (N_14806,N_14147,N_14368);
nand U14807 (N_14807,N_14074,N_14375);
nor U14808 (N_14808,N_14171,N_14128);
and U14809 (N_14809,N_14443,N_14307);
xnor U14810 (N_14810,N_14385,N_14468);
xor U14811 (N_14811,N_14408,N_14238);
nor U14812 (N_14812,N_14029,N_14459);
or U14813 (N_14813,N_14271,N_14188);
and U14814 (N_14814,N_14185,N_14365);
and U14815 (N_14815,N_14269,N_14319);
nor U14816 (N_14816,N_14425,N_14059);
xor U14817 (N_14817,N_14204,N_14158);
nand U14818 (N_14818,N_14228,N_14241);
nand U14819 (N_14819,N_14250,N_14023);
and U14820 (N_14820,N_14489,N_14265);
and U14821 (N_14821,N_14138,N_14471);
and U14822 (N_14822,N_14360,N_14273);
or U14823 (N_14823,N_14166,N_14454);
nand U14824 (N_14824,N_14194,N_14171);
nor U14825 (N_14825,N_14153,N_14375);
or U14826 (N_14826,N_14293,N_14423);
nor U14827 (N_14827,N_14306,N_14094);
and U14828 (N_14828,N_14029,N_14298);
nand U14829 (N_14829,N_14134,N_14233);
nand U14830 (N_14830,N_14365,N_14123);
and U14831 (N_14831,N_14409,N_14300);
or U14832 (N_14832,N_14332,N_14013);
nor U14833 (N_14833,N_14093,N_14110);
nor U14834 (N_14834,N_14065,N_14098);
or U14835 (N_14835,N_14018,N_14366);
xor U14836 (N_14836,N_14475,N_14009);
and U14837 (N_14837,N_14256,N_14454);
nor U14838 (N_14838,N_14071,N_14062);
or U14839 (N_14839,N_14242,N_14466);
xor U14840 (N_14840,N_14302,N_14362);
and U14841 (N_14841,N_14479,N_14293);
and U14842 (N_14842,N_14489,N_14031);
xor U14843 (N_14843,N_14407,N_14186);
xor U14844 (N_14844,N_14160,N_14445);
and U14845 (N_14845,N_14083,N_14489);
nor U14846 (N_14846,N_14455,N_14303);
xnor U14847 (N_14847,N_14103,N_14350);
and U14848 (N_14848,N_14079,N_14103);
or U14849 (N_14849,N_14094,N_14355);
xor U14850 (N_14850,N_14234,N_14266);
or U14851 (N_14851,N_14436,N_14306);
nand U14852 (N_14852,N_14158,N_14368);
and U14853 (N_14853,N_14261,N_14449);
or U14854 (N_14854,N_14087,N_14359);
xor U14855 (N_14855,N_14171,N_14051);
or U14856 (N_14856,N_14345,N_14277);
nor U14857 (N_14857,N_14475,N_14050);
and U14858 (N_14858,N_14331,N_14263);
or U14859 (N_14859,N_14242,N_14286);
and U14860 (N_14860,N_14316,N_14177);
or U14861 (N_14861,N_14022,N_14011);
nor U14862 (N_14862,N_14223,N_14352);
or U14863 (N_14863,N_14119,N_14167);
xor U14864 (N_14864,N_14173,N_14368);
xnor U14865 (N_14865,N_14095,N_14263);
xnor U14866 (N_14866,N_14462,N_14497);
nand U14867 (N_14867,N_14061,N_14492);
or U14868 (N_14868,N_14435,N_14250);
and U14869 (N_14869,N_14051,N_14339);
nand U14870 (N_14870,N_14263,N_14434);
xor U14871 (N_14871,N_14363,N_14125);
or U14872 (N_14872,N_14012,N_14464);
and U14873 (N_14873,N_14094,N_14008);
or U14874 (N_14874,N_14460,N_14257);
xor U14875 (N_14875,N_14126,N_14259);
and U14876 (N_14876,N_14312,N_14421);
or U14877 (N_14877,N_14073,N_14221);
nand U14878 (N_14878,N_14103,N_14234);
nor U14879 (N_14879,N_14270,N_14448);
xor U14880 (N_14880,N_14217,N_14380);
nand U14881 (N_14881,N_14293,N_14486);
nor U14882 (N_14882,N_14385,N_14390);
nor U14883 (N_14883,N_14188,N_14071);
and U14884 (N_14884,N_14359,N_14470);
and U14885 (N_14885,N_14291,N_14402);
or U14886 (N_14886,N_14217,N_14178);
or U14887 (N_14887,N_14443,N_14484);
xnor U14888 (N_14888,N_14036,N_14116);
and U14889 (N_14889,N_14333,N_14458);
nand U14890 (N_14890,N_14006,N_14011);
xor U14891 (N_14891,N_14162,N_14287);
xnor U14892 (N_14892,N_14319,N_14461);
xor U14893 (N_14893,N_14105,N_14234);
xor U14894 (N_14894,N_14178,N_14225);
xnor U14895 (N_14895,N_14494,N_14326);
or U14896 (N_14896,N_14113,N_14162);
xnor U14897 (N_14897,N_14317,N_14224);
and U14898 (N_14898,N_14150,N_14189);
xnor U14899 (N_14899,N_14361,N_14227);
nand U14900 (N_14900,N_14041,N_14419);
nor U14901 (N_14901,N_14449,N_14294);
or U14902 (N_14902,N_14140,N_14308);
and U14903 (N_14903,N_14005,N_14411);
and U14904 (N_14904,N_14078,N_14061);
nor U14905 (N_14905,N_14464,N_14367);
and U14906 (N_14906,N_14440,N_14216);
xor U14907 (N_14907,N_14108,N_14225);
nor U14908 (N_14908,N_14095,N_14091);
or U14909 (N_14909,N_14368,N_14333);
nand U14910 (N_14910,N_14125,N_14266);
nand U14911 (N_14911,N_14125,N_14206);
nor U14912 (N_14912,N_14321,N_14483);
nor U14913 (N_14913,N_14383,N_14008);
and U14914 (N_14914,N_14462,N_14389);
nor U14915 (N_14915,N_14261,N_14467);
nor U14916 (N_14916,N_14266,N_14363);
nand U14917 (N_14917,N_14278,N_14311);
or U14918 (N_14918,N_14163,N_14474);
nand U14919 (N_14919,N_14295,N_14171);
and U14920 (N_14920,N_14430,N_14175);
nand U14921 (N_14921,N_14085,N_14463);
or U14922 (N_14922,N_14296,N_14320);
xnor U14923 (N_14923,N_14134,N_14361);
or U14924 (N_14924,N_14441,N_14251);
nor U14925 (N_14925,N_14295,N_14151);
nand U14926 (N_14926,N_14030,N_14042);
or U14927 (N_14927,N_14234,N_14040);
and U14928 (N_14928,N_14204,N_14364);
xnor U14929 (N_14929,N_14245,N_14177);
xnor U14930 (N_14930,N_14416,N_14194);
or U14931 (N_14931,N_14406,N_14088);
xnor U14932 (N_14932,N_14114,N_14055);
nor U14933 (N_14933,N_14383,N_14139);
and U14934 (N_14934,N_14117,N_14333);
xor U14935 (N_14935,N_14197,N_14410);
nand U14936 (N_14936,N_14015,N_14259);
or U14937 (N_14937,N_14447,N_14104);
xnor U14938 (N_14938,N_14077,N_14095);
xor U14939 (N_14939,N_14027,N_14263);
or U14940 (N_14940,N_14233,N_14037);
nand U14941 (N_14941,N_14251,N_14132);
nor U14942 (N_14942,N_14018,N_14353);
or U14943 (N_14943,N_14117,N_14216);
xnor U14944 (N_14944,N_14218,N_14377);
nand U14945 (N_14945,N_14171,N_14103);
nor U14946 (N_14946,N_14329,N_14336);
or U14947 (N_14947,N_14038,N_14205);
or U14948 (N_14948,N_14180,N_14118);
xor U14949 (N_14949,N_14439,N_14193);
and U14950 (N_14950,N_14209,N_14199);
or U14951 (N_14951,N_14044,N_14203);
nor U14952 (N_14952,N_14474,N_14300);
xor U14953 (N_14953,N_14462,N_14038);
nand U14954 (N_14954,N_14126,N_14293);
nand U14955 (N_14955,N_14251,N_14178);
or U14956 (N_14956,N_14009,N_14238);
nand U14957 (N_14957,N_14476,N_14491);
and U14958 (N_14958,N_14357,N_14100);
nand U14959 (N_14959,N_14275,N_14213);
or U14960 (N_14960,N_14478,N_14359);
or U14961 (N_14961,N_14339,N_14345);
xor U14962 (N_14962,N_14337,N_14170);
and U14963 (N_14963,N_14046,N_14072);
nor U14964 (N_14964,N_14156,N_14236);
or U14965 (N_14965,N_14192,N_14022);
nor U14966 (N_14966,N_14143,N_14022);
nand U14967 (N_14967,N_14204,N_14411);
nand U14968 (N_14968,N_14221,N_14022);
nor U14969 (N_14969,N_14291,N_14492);
xor U14970 (N_14970,N_14082,N_14156);
or U14971 (N_14971,N_14486,N_14344);
and U14972 (N_14972,N_14266,N_14212);
and U14973 (N_14973,N_14452,N_14335);
xor U14974 (N_14974,N_14200,N_14176);
or U14975 (N_14975,N_14423,N_14420);
and U14976 (N_14976,N_14009,N_14012);
nor U14977 (N_14977,N_14374,N_14379);
nor U14978 (N_14978,N_14429,N_14257);
nor U14979 (N_14979,N_14460,N_14416);
nand U14980 (N_14980,N_14076,N_14192);
nor U14981 (N_14981,N_14192,N_14051);
xor U14982 (N_14982,N_14092,N_14169);
xnor U14983 (N_14983,N_14147,N_14227);
and U14984 (N_14984,N_14470,N_14317);
nor U14985 (N_14985,N_14322,N_14312);
nor U14986 (N_14986,N_14493,N_14219);
nand U14987 (N_14987,N_14068,N_14105);
or U14988 (N_14988,N_14386,N_14052);
nand U14989 (N_14989,N_14024,N_14011);
or U14990 (N_14990,N_14236,N_14327);
and U14991 (N_14991,N_14265,N_14361);
or U14992 (N_14992,N_14292,N_14255);
xnor U14993 (N_14993,N_14485,N_14152);
nand U14994 (N_14994,N_14483,N_14008);
xor U14995 (N_14995,N_14114,N_14231);
or U14996 (N_14996,N_14495,N_14465);
or U14997 (N_14997,N_14263,N_14202);
or U14998 (N_14998,N_14376,N_14007);
nor U14999 (N_14999,N_14104,N_14247);
or U15000 (N_15000,N_14984,N_14555);
nor U15001 (N_15001,N_14685,N_14930);
and U15002 (N_15002,N_14785,N_14514);
and U15003 (N_15003,N_14762,N_14970);
nand U15004 (N_15004,N_14730,N_14746);
xor U15005 (N_15005,N_14606,N_14946);
or U15006 (N_15006,N_14764,N_14739);
xor U15007 (N_15007,N_14879,N_14923);
or U15008 (N_15008,N_14819,N_14759);
or U15009 (N_15009,N_14605,N_14773);
nand U15010 (N_15010,N_14980,N_14848);
or U15011 (N_15011,N_14578,N_14540);
or U15012 (N_15012,N_14951,N_14736);
or U15013 (N_15013,N_14586,N_14925);
xor U15014 (N_15014,N_14654,N_14875);
nand U15015 (N_15015,N_14636,N_14818);
nand U15016 (N_15016,N_14684,N_14844);
and U15017 (N_15017,N_14884,N_14895);
nor U15018 (N_15018,N_14999,N_14571);
nor U15019 (N_15019,N_14554,N_14883);
xor U15020 (N_15020,N_14594,N_14994);
nor U15021 (N_15021,N_14691,N_14872);
or U15022 (N_15022,N_14500,N_14655);
xor U15023 (N_15023,N_14678,N_14607);
or U15024 (N_15024,N_14993,N_14790);
nor U15025 (N_15025,N_14502,N_14569);
or U15026 (N_15026,N_14885,N_14972);
nor U15027 (N_15027,N_14829,N_14513);
or U15028 (N_15028,N_14836,N_14783);
nor U15029 (N_15029,N_14711,N_14572);
and U15030 (N_15030,N_14556,N_14698);
nand U15031 (N_15031,N_14763,N_14743);
or U15032 (N_15032,N_14867,N_14646);
nor U15033 (N_15033,N_14859,N_14512);
xor U15034 (N_15034,N_14667,N_14553);
nor U15035 (N_15035,N_14516,N_14754);
or U15036 (N_15036,N_14950,N_14662);
and U15037 (N_15037,N_14893,N_14505);
and U15038 (N_15038,N_14985,N_14837);
nand U15039 (N_15039,N_14589,N_14830);
or U15040 (N_15040,N_14543,N_14682);
nand U15041 (N_15041,N_14909,N_14535);
xnor U15042 (N_15042,N_14604,N_14888);
nand U15043 (N_15043,N_14728,N_14537);
xor U15044 (N_15044,N_14780,N_14528);
nor U15045 (N_15045,N_14596,N_14561);
nand U15046 (N_15046,N_14849,N_14576);
and U15047 (N_15047,N_14842,N_14778);
xor U15048 (N_15048,N_14936,N_14597);
xnor U15049 (N_15049,N_14957,N_14622);
nand U15050 (N_15050,N_14550,N_14665);
and U15051 (N_15051,N_14916,N_14575);
nand U15052 (N_15052,N_14983,N_14737);
nor U15053 (N_15053,N_14742,N_14927);
nor U15054 (N_15054,N_14799,N_14881);
nand U15055 (N_15055,N_14988,N_14966);
nand U15056 (N_15056,N_14886,N_14542);
and U15057 (N_15057,N_14788,N_14639);
xor U15058 (N_15058,N_14979,N_14977);
nand U15059 (N_15059,N_14890,N_14536);
or U15060 (N_15060,N_14962,N_14960);
nand U15061 (N_15061,N_14861,N_14526);
xnor U15062 (N_15062,N_14769,N_14629);
nand U15063 (N_15063,N_14593,N_14928);
and U15064 (N_15064,N_14887,N_14677);
nand U15065 (N_15065,N_14720,N_14624);
nand U15066 (N_15066,N_14789,N_14915);
and U15067 (N_15067,N_14847,N_14775);
nor U15068 (N_15068,N_14545,N_14738);
xnor U15069 (N_15069,N_14715,N_14855);
nand U15070 (N_15070,N_14638,N_14515);
nand U15071 (N_15071,N_14838,N_14782);
xor U15072 (N_15072,N_14753,N_14548);
and U15073 (N_15073,N_14889,N_14748);
or U15074 (N_15074,N_14843,N_14574);
xor U15075 (N_15075,N_14852,N_14897);
xor U15076 (N_15076,N_14722,N_14801);
and U15077 (N_15077,N_14958,N_14876);
and U15078 (N_15078,N_14906,N_14940);
xor U15079 (N_15079,N_14564,N_14530);
xnor U15080 (N_15080,N_14935,N_14544);
or U15081 (N_15081,N_14995,N_14756);
xor U15082 (N_15082,N_14992,N_14534);
nand U15083 (N_15083,N_14953,N_14944);
or U15084 (N_15084,N_14527,N_14573);
xor U15085 (N_15085,N_14705,N_14912);
nor U15086 (N_15086,N_14635,N_14702);
nand U15087 (N_15087,N_14614,N_14733);
and U15088 (N_15088,N_14750,N_14856);
and U15089 (N_15089,N_14541,N_14539);
and U15090 (N_15090,N_14663,N_14834);
xnor U15091 (N_15091,N_14587,N_14922);
nor U15092 (N_15092,N_14640,N_14501);
and U15093 (N_15093,N_14652,N_14968);
xor U15094 (N_15094,N_14701,N_14904);
nor U15095 (N_15095,N_14529,N_14860);
or U15096 (N_15096,N_14615,N_14522);
nand U15097 (N_15097,N_14643,N_14786);
nand U15098 (N_15098,N_14570,N_14792);
xnor U15099 (N_15099,N_14841,N_14592);
xnor U15100 (N_15100,N_14892,N_14680);
nand U15101 (N_15101,N_14933,N_14508);
nand U15102 (N_15102,N_14880,N_14582);
and U15103 (N_15103,N_14976,N_14645);
and U15104 (N_15104,N_14523,N_14600);
or U15105 (N_15105,N_14507,N_14943);
and U15106 (N_15106,N_14598,N_14560);
nand U15107 (N_15107,N_14712,N_14812);
xnor U15108 (N_15108,N_14903,N_14531);
nand U15109 (N_15109,N_14590,N_14779);
nand U15110 (N_15110,N_14719,N_14637);
nand U15111 (N_15111,N_14520,N_14760);
nand U15112 (N_15112,N_14625,N_14709);
nand U15113 (N_15113,N_14693,N_14631);
nor U15114 (N_15114,N_14891,N_14755);
nand U15115 (N_15115,N_14749,N_14716);
and U15116 (N_15116,N_14850,N_14732);
and U15117 (N_15117,N_14621,N_14731);
or U15118 (N_15118,N_14565,N_14566);
nand U15119 (N_15119,N_14696,N_14896);
nand U15120 (N_15120,N_14681,N_14595);
xor U15121 (N_15121,N_14686,N_14692);
nor U15122 (N_15122,N_14558,N_14918);
xnor U15123 (N_15123,N_14648,N_14809);
xor U15124 (N_15124,N_14617,N_14616);
or U15125 (N_15125,N_14899,N_14557);
nand U15126 (N_15126,N_14741,N_14794);
nand U15127 (N_15127,N_14661,N_14873);
xnor U15128 (N_15128,N_14945,N_14659);
or U15129 (N_15129,N_14931,N_14929);
nand U15130 (N_15130,N_14959,N_14815);
nor U15131 (N_15131,N_14688,N_14757);
nor U15132 (N_15132,N_14632,N_14577);
or U15133 (N_15133,N_14700,N_14552);
or U15134 (N_15134,N_14651,N_14768);
nor U15135 (N_15135,N_14932,N_14986);
xor U15136 (N_15136,N_14767,N_14689);
nor U15137 (N_15137,N_14690,N_14703);
xnor U15138 (N_15138,N_14774,N_14644);
and U15139 (N_15139,N_14619,N_14997);
and U15140 (N_15140,N_14710,N_14973);
and U15141 (N_15141,N_14911,N_14770);
and U15142 (N_15142,N_14825,N_14533);
xnor U15143 (N_15143,N_14559,N_14725);
xor U15144 (N_15144,N_14562,N_14865);
or U15145 (N_15145,N_14900,N_14991);
xnor U15146 (N_15146,N_14664,N_14694);
and U15147 (N_15147,N_14580,N_14695);
nand U15148 (N_15148,N_14905,N_14870);
nand U15149 (N_15149,N_14802,N_14752);
nand U15150 (N_15150,N_14798,N_14724);
or U15151 (N_15151,N_14877,N_14969);
nand U15152 (N_15152,N_14858,N_14990);
nand U15153 (N_15153,N_14714,N_14603);
nand U15154 (N_15154,N_14823,N_14669);
or U15155 (N_15155,N_14744,N_14967);
or U15156 (N_15156,N_14766,N_14998);
nor U15157 (N_15157,N_14630,N_14921);
nand U15158 (N_15158,N_14804,N_14660);
or U15159 (N_15159,N_14729,N_14914);
nand U15160 (N_15160,N_14517,N_14941);
nand U15161 (N_15161,N_14797,N_14811);
xnor U15162 (N_15162,N_14717,N_14675);
xor U15163 (N_15163,N_14683,N_14882);
nand U15164 (N_15164,N_14924,N_14816);
nand U15165 (N_15165,N_14939,N_14869);
nand U15166 (N_15166,N_14866,N_14525);
nor U15167 (N_15167,N_14504,N_14699);
or U15168 (N_15168,N_14628,N_14735);
and U15169 (N_15169,N_14734,N_14996);
xnor U15170 (N_15170,N_14707,N_14676);
or U15171 (N_15171,N_14547,N_14673);
or U15172 (N_15172,N_14697,N_14795);
or U15173 (N_15173,N_14751,N_14926);
and U15174 (N_15174,N_14781,N_14807);
or U15175 (N_15175,N_14777,N_14828);
nor U15176 (N_15176,N_14808,N_14956);
or U15177 (N_15177,N_14568,N_14810);
nand U15178 (N_15178,N_14549,N_14671);
xor U15179 (N_15179,N_14670,N_14851);
xor U15180 (N_15180,N_14839,N_14987);
or U15181 (N_15181,N_14938,N_14955);
xnor U15182 (N_15182,N_14687,N_14832);
nand U15183 (N_15183,N_14563,N_14898);
and U15184 (N_15184,N_14620,N_14947);
nand U15185 (N_15185,N_14579,N_14796);
or U15186 (N_15186,N_14524,N_14583);
xnor U15187 (N_15187,N_14917,N_14588);
and U15188 (N_15188,N_14627,N_14942);
xor U15189 (N_15189,N_14863,N_14854);
xnor U15190 (N_15190,N_14964,N_14723);
nand U15191 (N_15191,N_14610,N_14642);
nand U15192 (N_15192,N_14846,N_14989);
or U15193 (N_15193,N_14599,N_14982);
and U15194 (N_15194,N_14845,N_14878);
nor U15195 (N_15195,N_14585,N_14765);
xor U15196 (N_15196,N_14814,N_14666);
nor U15197 (N_15197,N_14817,N_14803);
nor U15198 (N_15198,N_14668,N_14726);
nor U15199 (N_15199,N_14511,N_14641);
nand U15200 (N_15200,N_14567,N_14813);
xor U15201 (N_15201,N_14907,N_14672);
nand U15202 (N_15202,N_14840,N_14704);
and U15203 (N_15203,N_14919,N_14706);
or U15204 (N_15204,N_14902,N_14833);
nand U15205 (N_15205,N_14868,N_14713);
and U15206 (N_15206,N_14509,N_14650);
or U15207 (N_15207,N_14934,N_14747);
or U15208 (N_15208,N_14937,N_14961);
or U15209 (N_15209,N_14963,N_14784);
xnor U15210 (N_15210,N_14626,N_14975);
nand U15211 (N_15211,N_14821,N_14827);
and U15212 (N_15212,N_14824,N_14835);
and U15213 (N_15213,N_14623,N_14656);
or U15214 (N_15214,N_14581,N_14974);
nand U15215 (N_15215,N_14551,N_14674);
or U15216 (N_15216,N_14612,N_14949);
and U15217 (N_15217,N_14820,N_14679);
or U15218 (N_15218,N_14634,N_14800);
or U15219 (N_15219,N_14948,N_14793);
nor U15220 (N_15220,N_14831,N_14546);
xor U15221 (N_15221,N_14965,N_14978);
nand U15222 (N_15222,N_14971,N_14761);
xnor U15223 (N_15223,N_14658,N_14727);
or U15224 (N_15224,N_14826,N_14601);
and U15225 (N_15225,N_14805,N_14822);
or U15226 (N_15226,N_14718,N_14894);
xnor U15227 (N_15227,N_14874,N_14721);
nor U15228 (N_15228,N_14871,N_14521);
xnor U15229 (N_15229,N_14864,N_14538);
xor U15230 (N_15230,N_14901,N_14758);
nand U15231 (N_15231,N_14776,N_14952);
and U15232 (N_15232,N_14613,N_14602);
nand U15233 (N_15233,N_14745,N_14772);
xnor U15234 (N_15234,N_14708,N_14857);
xor U15235 (N_15235,N_14611,N_14771);
xor U15236 (N_15236,N_14787,N_14532);
or U15237 (N_15237,N_14853,N_14647);
nand U15238 (N_15238,N_14649,N_14519);
and U15239 (N_15239,N_14633,N_14740);
nor U15240 (N_15240,N_14913,N_14908);
nand U15241 (N_15241,N_14584,N_14981);
xnor U15242 (N_15242,N_14591,N_14806);
nand U15243 (N_15243,N_14608,N_14653);
xor U15244 (N_15244,N_14510,N_14657);
nor U15245 (N_15245,N_14618,N_14862);
nor U15246 (N_15246,N_14503,N_14954);
nand U15247 (N_15247,N_14506,N_14920);
xnor U15248 (N_15248,N_14791,N_14910);
xor U15249 (N_15249,N_14518,N_14609);
nand U15250 (N_15250,N_14810,N_14749);
nand U15251 (N_15251,N_14760,N_14876);
nand U15252 (N_15252,N_14554,N_14800);
nor U15253 (N_15253,N_14712,N_14652);
and U15254 (N_15254,N_14685,N_14580);
and U15255 (N_15255,N_14920,N_14951);
nor U15256 (N_15256,N_14635,N_14831);
or U15257 (N_15257,N_14676,N_14752);
and U15258 (N_15258,N_14718,N_14994);
and U15259 (N_15259,N_14958,N_14950);
xor U15260 (N_15260,N_14521,N_14872);
and U15261 (N_15261,N_14894,N_14640);
nor U15262 (N_15262,N_14989,N_14912);
nand U15263 (N_15263,N_14942,N_14717);
or U15264 (N_15264,N_14509,N_14667);
nand U15265 (N_15265,N_14853,N_14799);
xor U15266 (N_15266,N_14848,N_14923);
or U15267 (N_15267,N_14603,N_14938);
nand U15268 (N_15268,N_14955,N_14888);
xnor U15269 (N_15269,N_14885,N_14535);
nor U15270 (N_15270,N_14779,N_14843);
xnor U15271 (N_15271,N_14554,N_14982);
nor U15272 (N_15272,N_14639,N_14871);
nand U15273 (N_15273,N_14870,N_14639);
nor U15274 (N_15274,N_14733,N_14744);
nand U15275 (N_15275,N_14734,N_14746);
nand U15276 (N_15276,N_14635,N_14753);
xor U15277 (N_15277,N_14670,N_14773);
xor U15278 (N_15278,N_14679,N_14547);
nand U15279 (N_15279,N_14541,N_14771);
nor U15280 (N_15280,N_14716,N_14906);
and U15281 (N_15281,N_14998,N_14980);
nand U15282 (N_15282,N_14551,N_14953);
xor U15283 (N_15283,N_14591,N_14848);
xnor U15284 (N_15284,N_14798,N_14556);
or U15285 (N_15285,N_14532,N_14652);
nand U15286 (N_15286,N_14546,N_14850);
or U15287 (N_15287,N_14751,N_14589);
or U15288 (N_15288,N_14996,N_14889);
nand U15289 (N_15289,N_14640,N_14910);
nand U15290 (N_15290,N_14531,N_14737);
nand U15291 (N_15291,N_14615,N_14653);
nand U15292 (N_15292,N_14780,N_14828);
nor U15293 (N_15293,N_14944,N_14661);
or U15294 (N_15294,N_14695,N_14620);
nand U15295 (N_15295,N_14649,N_14787);
or U15296 (N_15296,N_14675,N_14680);
nand U15297 (N_15297,N_14504,N_14901);
and U15298 (N_15298,N_14544,N_14511);
or U15299 (N_15299,N_14985,N_14505);
nor U15300 (N_15300,N_14524,N_14951);
or U15301 (N_15301,N_14627,N_14733);
or U15302 (N_15302,N_14840,N_14906);
and U15303 (N_15303,N_14705,N_14723);
nor U15304 (N_15304,N_14671,N_14633);
xnor U15305 (N_15305,N_14829,N_14703);
and U15306 (N_15306,N_14543,N_14629);
nand U15307 (N_15307,N_14819,N_14761);
or U15308 (N_15308,N_14542,N_14808);
or U15309 (N_15309,N_14669,N_14591);
xor U15310 (N_15310,N_14818,N_14815);
and U15311 (N_15311,N_14631,N_14605);
xnor U15312 (N_15312,N_14907,N_14842);
xor U15313 (N_15313,N_14961,N_14900);
xnor U15314 (N_15314,N_14598,N_14567);
and U15315 (N_15315,N_14726,N_14967);
nand U15316 (N_15316,N_14799,N_14506);
nor U15317 (N_15317,N_14952,N_14519);
xor U15318 (N_15318,N_14557,N_14765);
xor U15319 (N_15319,N_14750,N_14606);
and U15320 (N_15320,N_14899,N_14742);
or U15321 (N_15321,N_14902,N_14939);
and U15322 (N_15322,N_14795,N_14912);
xnor U15323 (N_15323,N_14625,N_14681);
xor U15324 (N_15324,N_14922,N_14939);
xor U15325 (N_15325,N_14653,N_14613);
nand U15326 (N_15326,N_14509,N_14741);
or U15327 (N_15327,N_14606,N_14837);
nor U15328 (N_15328,N_14693,N_14551);
or U15329 (N_15329,N_14801,N_14786);
nor U15330 (N_15330,N_14560,N_14573);
nand U15331 (N_15331,N_14701,N_14950);
xor U15332 (N_15332,N_14978,N_14794);
nor U15333 (N_15333,N_14510,N_14955);
nor U15334 (N_15334,N_14548,N_14799);
nand U15335 (N_15335,N_14515,N_14547);
nand U15336 (N_15336,N_14933,N_14877);
nand U15337 (N_15337,N_14832,N_14530);
and U15338 (N_15338,N_14511,N_14900);
xnor U15339 (N_15339,N_14767,N_14965);
and U15340 (N_15340,N_14584,N_14677);
and U15341 (N_15341,N_14752,N_14700);
nor U15342 (N_15342,N_14905,N_14831);
nor U15343 (N_15343,N_14844,N_14592);
xnor U15344 (N_15344,N_14720,N_14865);
nor U15345 (N_15345,N_14690,N_14901);
nand U15346 (N_15346,N_14572,N_14933);
xor U15347 (N_15347,N_14660,N_14927);
xnor U15348 (N_15348,N_14598,N_14890);
nor U15349 (N_15349,N_14691,N_14624);
nor U15350 (N_15350,N_14694,N_14643);
nor U15351 (N_15351,N_14857,N_14673);
or U15352 (N_15352,N_14558,N_14512);
or U15353 (N_15353,N_14531,N_14860);
nor U15354 (N_15354,N_14542,N_14853);
or U15355 (N_15355,N_14917,N_14506);
or U15356 (N_15356,N_14631,N_14772);
or U15357 (N_15357,N_14920,N_14675);
nor U15358 (N_15358,N_14591,N_14503);
nor U15359 (N_15359,N_14975,N_14776);
and U15360 (N_15360,N_14946,N_14687);
nor U15361 (N_15361,N_14753,N_14824);
or U15362 (N_15362,N_14577,N_14803);
and U15363 (N_15363,N_14598,N_14896);
nor U15364 (N_15364,N_14713,N_14956);
xnor U15365 (N_15365,N_14814,N_14535);
nor U15366 (N_15366,N_14779,N_14881);
nor U15367 (N_15367,N_14815,N_14870);
and U15368 (N_15368,N_14971,N_14810);
nand U15369 (N_15369,N_14970,N_14830);
or U15370 (N_15370,N_14734,N_14682);
and U15371 (N_15371,N_14744,N_14704);
or U15372 (N_15372,N_14812,N_14636);
nand U15373 (N_15373,N_14557,N_14686);
or U15374 (N_15374,N_14623,N_14977);
or U15375 (N_15375,N_14807,N_14677);
nand U15376 (N_15376,N_14602,N_14644);
nor U15377 (N_15377,N_14803,N_14729);
or U15378 (N_15378,N_14805,N_14712);
nor U15379 (N_15379,N_14777,N_14594);
xnor U15380 (N_15380,N_14993,N_14739);
nand U15381 (N_15381,N_14623,N_14680);
or U15382 (N_15382,N_14706,N_14579);
nand U15383 (N_15383,N_14862,N_14649);
or U15384 (N_15384,N_14540,N_14759);
nand U15385 (N_15385,N_14983,N_14930);
nand U15386 (N_15386,N_14949,N_14641);
or U15387 (N_15387,N_14800,N_14673);
nand U15388 (N_15388,N_14755,N_14886);
nand U15389 (N_15389,N_14888,N_14689);
and U15390 (N_15390,N_14799,N_14679);
nand U15391 (N_15391,N_14809,N_14766);
xnor U15392 (N_15392,N_14975,N_14791);
nor U15393 (N_15393,N_14853,N_14708);
xor U15394 (N_15394,N_14746,N_14562);
nand U15395 (N_15395,N_14759,N_14754);
nand U15396 (N_15396,N_14637,N_14703);
and U15397 (N_15397,N_14849,N_14749);
nor U15398 (N_15398,N_14659,N_14751);
or U15399 (N_15399,N_14590,N_14529);
nand U15400 (N_15400,N_14778,N_14606);
xnor U15401 (N_15401,N_14959,N_14908);
and U15402 (N_15402,N_14589,N_14692);
xor U15403 (N_15403,N_14692,N_14562);
and U15404 (N_15404,N_14528,N_14544);
or U15405 (N_15405,N_14846,N_14643);
nor U15406 (N_15406,N_14834,N_14830);
xnor U15407 (N_15407,N_14620,N_14530);
nand U15408 (N_15408,N_14922,N_14522);
nor U15409 (N_15409,N_14809,N_14570);
and U15410 (N_15410,N_14944,N_14630);
xnor U15411 (N_15411,N_14990,N_14908);
nor U15412 (N_15412,N_14777,N_14952);
nor U15413 (N_15413,N_14625,N_14946);
xor U15414 (N_15414,N_14813,N_14640);
and U15415 (N_15415,N_14603,N_14972);
and U15416 (N_15416,N_14666,N_14712);
or U15417 (N_15417,N_14764,N_14614);
and U15418 (N_15418,N_14707,N_14841);
nand U15419 (N_15419,N_14674,N_14828);
and U15420 (N_15420,N_14976,N_14992);
nand U15421 (N_15421,N_14681,N_14701);
and U15422 (N_15422,N_14733,N_14804);
and U15423 (N_15423,N_14885,N_14850);
and U15424 (N_15424,N_14735,N_14575);
nand U15425 (N_15425,N_14598,N_14738);
and U15426 (N_15426,N_14624,N_14636);
nor U15427 (N_15427,N_14964,N_14610);
nand U15428 (N_15428,N_14932,N_14741);
nand U15429 (N_15429,N_14513,N_14518);
xor U15430 (N_15430,N_14742,N_14834);
and U15431 (N_15431,N_14724,N_14999);
and U15432 (N_15432,N_14959,N_14593);
and U15433 (N_15433,N_14707,N_14577);
nand U15434 (N_15434,N_14854,N_14951);
nand U15435 (N_15435,N_14881,N_14915);
nand U15436 (N_15436,N_14997,N_14757);
nand U15437 (N_15437,N_14546,N_14507);
and U15438 (N_15438,N_14803,N_14847);
or U15439 (N_15439,N_14527,N_14663);
or U15440 (N_15440,N_14591,N_14609);
and U15441 (N_15441,N_14740,N_14657);
nand U15442 (N_15442,N_14971,N_14616);
xor U15443 (N_15443,N_14991,N_14954);
or U15444 (N_15444,N_14836,N_14699);
nand U15445 (N_15445,N_14965,N_14545);
xor U15446 (N_15446,N_14690,N_14547);
and U15447 (N_15447,N_14754,N_14544);
or U15448 (N_15448,N_14755,N_14560);
and U15449 (N_15449,N_14996,N_14719);
or U15450 (N_15450,N_14584,N_14924);
nor U15451 (N_15451,N_14622,N_14847);
or U15452 (N_15452,N_14676,N_14985);
or U15453 (N_15453,N_14769,N_14848);
nand U15454 (N_15454,N_14533,N_14665);
or U15455 (N_15455,N_14775,N_14885);
nand U15456 (N_15456,N_14621,N_14976);
xor U15457 (N_15457,N_14586,N_14679);
and U15458 (N_15458,N_14581,N_14663);
xnor U15459 (N_15459,N_14736,N_14536);
and U15460 (N_15460,N_14759,N_14756);
nand U15461 (N_15461,N_14593,N_14996);
or U15462 (N_15462,N_14922,N_14925);
nand U15463 (N_15463,N_14602,N_14897);
xnor U15464 (N_15464,N_14984,N_14720);
or U15465 (N_15465,N_14722,N_14695);
nand U15466 (N_15466,N_14671,N_14524);
xor U15467 (N_15467,N_14798,N_14895);
or U15468 (N_15468,N_14980,N_14881);
nand U15469 (N_15469,N_14588,N_14628);
or U15470 (N_15470,N_14614,N_14876);
nand U15471 (N_15471,N_14671,N_14990);
nor U15472 (N_15472,N_14585,N_14635);
nand U15473 (N_15473,N_14808,N_14718);
nand U15474 (N_15474,N_14611,N_14912);
or U15475 (N_15475,N_14658,N_14928);
or U15476 (N_15476,N_14597,N_14912);
xor U15477 (N_15477,N_14840,N_14539);
xor U15478 (N_15478,N_14940,N_14826);
nand U15479 (N_15479,N_14663,N_14761);
or U15480 (N_15480,N_14729,N_14561);
xnor U15481 (N_15481,N_14780,N_14567);
xnor U15482 (N_15482,N_14809,N_14710);
nor U15483 (N_15483,N_14693,N_14740);
xor U15484 (N_15484,N_14602,N_14798);
nor U15485 (N_15485,N_14530,N_14758);
or U15486 (N_15486,N_14685,N_14898);
nor U15487 (N_15487,N_14898,N_14734);
and U15488 (N_15488,N_14707,N_14711);
nor U15489 (N_15489,N_14523,N_14693);
and U15490 (N_15490,N_14653,N_14595);
or U15491 (N_15491,N_14631,N_14624);
xor U15492 (N_15492,N_14998,N_14947);
nor U15493 (N_15493,N_14900,N_14724);
nor U15494 (N_15494,N_14857,N_14937);
xor U15495 (N_15495,N_14981,N_14516);
xor U15496 (N_15496,N_14511,N_14525);
nor U15497 (N_15497,N_14686,N_14629);
or U15498 (N_15498,N_14634,N_14877);
nor U15499 (N_15499,N_14776,N_14524);
nor U15500 (N_15500,N_15205,N_15103);
nand U15501 (N_15501,N_15319,N_15123);
nor U15502 (N_15502,N_15067,N_15152);
nor U15503 (N_15503,N_15132,N_15447);
and U15504 (N_15504,N_15015,N_15478);
nor U15505 (N_15505,N_15204,N_15337);
xor U15506 (N_15506,N_15266,N_15270);
and U15507 (N_15507,N_15332,N_15434);
nor U15508 (N_15508,N_15182,N_15353);
and U15509 (N_15509,N_15267,N_15079);
nand U15510 (N_15510,N_15364,N_15209);
xnor U15511 (N_15511,N_15352,N_15148);
or U15512 (N_15512,N_15240,N_15495);
and U15513 (N_15513,N_15170,N_15494);
xor U15514 (N_15514,N_15375,N_15039);
xor U15515 (N_15515,N_15143,N_15177);
and U15516 (N_15516,N_15395,N_15409);
nand U15517 (N_15517,N_15211,N_15051);
or U15518 (N_15518,N_15093,N_15191);
or U15519 (N_15519,N_15194,N_15292);
xor U15520 (N_15520,N_15066,N_15073);
and U15521 (N_15521,N_15376,N_15316);
nor U15522 (N_15522,N_15385,N_15324);
nand U15523 (N_15523,N_15308,N_15336);
xor U15524 (N_15524,N_15206,N_15176);
nor U15525 (N_15525,N_15305,N_15120);
xnor U15526 (N_15526,N_15081,N_15481);
xor U15527 (N_15527,N_15440,N_15471);
nand U15528 (N_15528,N_15338,N_15371);
xnor U15529 (N_15529,N_15411,N_15210);
or U15530 (N_15530,N_15173,N_15078);
nor U15531 (N_15531,N_15278,N_15091);
or U15532 (N_15532,N_15068,N_15055);
and U15533 (N_15533,N_15180,N_15219);
and U15534 (N_15534,N_15432,N_15258);
nand U15535 (N_15535,N_15181,N_15313);
nor U15536 (N_15536,N_15282,N_15442);
xnor U15537 (N_15537,N_15358,N_15228);
nor U15538 (N_15538,N_15381,N_15394);
or U15539 (N_15539,N_15168,N_15496);
nor U15540 (N_15540,N_15160,N_15196);
or U15541 (N_15541,N_15095,N_15377);
or U15542 (N_15542,N_15435,N_15455);
and U15543 (N_15543,N_15135,N_15074);
nor U15544 (N_15544,N_15264,N_15480);
nor U15545 (N_15545,N_15118,N_15053);
xor U15546 (N_15546,N_15001,N_15243);
or U15547 (N_15547,N_15167,N_15460);
nor U15548 (N_15548,N_15233,N_15226);
xnor U15549 (N_15549,N_15075,N_15320);
and U15550 (N_15550,N_15430,N_15198);
and U15551 (N_15551,N_15046,N_15351);
or U15552 (N_15552,N_15369,N_15466);
nand U15553 (N_15553,N_15248,N_15298);
nor U15554 (N_15554,N_15080,N_15229);
nand U15555 (N_15555,N_15145,N_15252);
or U15556 (N_15556,N_15222,N_15179);
or U15557 (N_15557,N_15098,N_15087);
or U15558 (N_15558,N_15431,N_15490);
or U15559 (N_15559,N_15105,N_15307);
xnor U15560 (N_15560,N_15311,N_15407);
nand U15561 (N_15561,N_15380,N_15201);
nand U15562 (N_15562,N_15279,N_15059);
xor U15563 (N_15563,N_15329,N_15467);
or U15564 (N_15564,N_15461,N_15464);
and U15565 (N_15565,N_15356,N_15048);
xor U15566 (N_15566,N_15111,N_15345);
xor U15567 (N_15567,N_15454,N_15134);
or U15568 (N_15568,N_15357,N_15388);
or U15569 (N_15569,N_15361,N_15330);
or U15570 (N_15570,N_15058,N_15367);
xnor U15571 (N_15571,N_15484,N_15296);
and U15572 (N_15572,N_15419,N_15485);
xor U15573 (N_15573,N_15005,N_15190);
xor U15574 (N_15574,N_15004,N_15113);
nand U15575 (N_15575,N_15343,N_15139);
and U15576 (N_15576,N_15444,N_15340);
nor U15577 (N_15577,N_15418,N_15421);
nor U15578 (N_15578,N_15011,N_15295);
xor U15579 (N_15579,N_15030,N_15404);
xor U15580 (N_15580,N_15085,N_15162);
or U15581 (N_15581,N_15112,N_15406);
or U15582 (N_15582,N_15144,N_15323);
or U15583 (N_15583,N_15374,N_15116);
nor U15584 (N_15584,N_15479,N_15086);
or U15585 (N_15585,N_15246,N_15497);
or U15586 (N_15586,N_15276,N_15433);
or U15587 (N_15587,N_15036,N_15187);
nor U15588 (N_15588,N_15293,N_15257);
nand U15589 (N_15589,N_15197,N_15477);
nor U15590 (N_15590,N_15038,N_15090);
xnor U15591 (N_15591,N_15334,N_15408);
and U15592 (N_15592,N_15403,N_15449);
or U15593 (N_15593,N_15268,N_15493);
nor U15594 (N_15594,N_15498,N_15189);
or U15595 (N_15595,N_15489,N_15284);
and U15596 (N_15596,N_15227,N_15096);
and U15597 (N_15597,N_15106,N_15032);
nand U15598 (N_15598,N_15070,N_15450);
or U15599 (N_15599,N_15328,N_15089);
nand U15600 (N_15600,N_15163,N_15384);
or U15601 (N_15601,N_15169,N_15373);
nand U15602 (N_15602,N_15127,N_15410);
nor U15603 (N_15603,N_15137,N_15186);
or U15604 (N_15604,N_15231,N_15425);
nand U15605 (N_15605,N_15441,N_15468);
and U15606 (N_15606,N_15473,N_15216);
or U15607 (N_15607,N_15289,N_15025);
and U15608 (N_15608,N_15138,N_15463);
xor U15609 (N_15609,N_15234,N_15288);
or U15610 (N_15610,N_15446,N_15420);
nor U15611 (N_15611,N_15133,N_15261);
nand U15612 (N_15612,N_15443,N_15347);
xnor U15613 (N_15613,N_15149,N_15126);
nor U15614 (N_15614,N_15237,N_15462);
xor U15615 (N_15615,N_15346,N_15301);
and U15616 (N_15616,N_15062,N_15034);
and U15617 (N_15617,N_15012,N_15023);
nor U15618 (N_15618,N_15212,N_15183);
nor U15619 (N_15619,N_15256,N_15459);
xnor U15620 (N_15620,N_15304,N_15457);
nand U15621 (N_15621,N_15448,N_15014);
nand U15622 (N_15622,N_15031,N_15124);
xnor U15623 (N_15623,N_15016,N_15121);
xor U15624 (N_15624,N_15047,N_15043);
nand U15625 (N_15625,N_15286,N_15220);
nor U15626 (N_15626,N_15392,N_15018);
nand U15627 (N_15627,N_15499,N_15341);
nand U15628 (N_15628,N_15439,N_15214);
or U15629 (N_15629,N_15315,N_15389);
nor U15630 (N_15630,N_15057,N_15063);
and U15631 (N_15631,N_15002,N_15064);
nand U15632 (N_15632,N_15291,N_15365);
or U15633 (N_15633,N_15396,N_15339);
nor U15634 (N_15634,N_15265,N_15076);
nand U15635 (N_15635,N_15154,N_15151);
and U15636 (N_15636,N_15129,N_15269);
xor U15637 (N_15637,N_15049,N_15317);
nand U15638 (N_15638,N_15263,N_15245);
xnor U15639 (N_15639,N_15028,N_15037);
xnor U15640 (N_15640,N_15101,N_15108);
nor U15641 (N_15641,N_15280,N_15000);
and U15642 (N_15642,N_15155,N_15349);
and U15643 (N_15643,N_15241,N_15363);
xor U15644 (N_15644,N_15094,N_15107);
nor U15645 (N_15645,N_15122,N_15322);
nand U15646 (N_15646,N_15232,N_15429);
nor U15647 (N_15647,N_15368,N_15125);
xnor U15648 (N_15648,N_15017,N_15156);
nand U15649 (N_15649,N_15050,N_15483);
or U15650 (N_15650,N_15221,N_15208);
xnor U15651 (N_15651,N_15027,N_15109);
nand U15652 (N_15652,N_15119,N_15488);
nand U15653 (N_15653,N_15042,N_15294);
nand U15654 (N_15654,N_15486,N_15424);
nor U15655 (N_15655,N_15146,N_15150);
and U15656 (N_15656,N_15013,N_15274);
or U15657 (N_15657,N_15006,N_15475);
or U15658 (N_15658,N_15161,N_15283);
nor U15659 (N_15659,N_15297,N_15456);
or U15660 (N_15660,N_15236,N_15366);
or U15661 (N_15661,N_15142,N_15092);
nand U15662 (N_15662,N_15326,N_15044);
nand U15663 (N_15663,N_15303,N_15415);
xnor U15664 (N_15664,N_15071,N_15040);
or U15665 (N_15665,N_15230,N_15223);
nand U15666 (N_15666,N_15195,N_15215);
and U15667 (N_15667,N_15166,N_15321);
or U15668 (N_15668,N_15354,N_15250);
or U15669 (N_15669,N_15312,N_15262);
or U15670 (N_15670,N_15438,N_15359);
xor U15671 (N_15671,N_15008,N_15054);
nand U15672 (N_15672,N_15147,N_15387);
or U15673 (N_15673,N_15379,N_15188);
nand U15674 (N_15674,N_15414,N_15199);
and U15675 (N_15675,N_15383,N_15386);
and U15676 (N_15676,N_15178,N_15117);
nor U15677 (N_15677,N_15203,N_15140);
nor U15678 (N_15678,N_15281,N_15325);
and U15679 (N_15679,N_15458,N_15172);
nor U15680 (N_15680,N_15225,N_15021);
and U15681 (N_15681,N_15104,N_15165);
nand U15682 (N_15682,N_15218,N_15242);
xor U15683 (N_15683,N_15402,N_15024);
nand U15684 (N_15684,N_15290,N_15007);
xor U15685 (N_15685,N_15251,N_15088);
nand U15686 (N_15686,N_15476,N_15390);
nor U15687 (N_15687,N_15399,N_15072);
xor U15688 (N_15688,N_15253,N_15193);
and U15689 (N_15689,N_15249,N_15041);
nor U15690 (N_15690,N_15426,N_15436);
nand U15691 (N_15691,N_15158,N_15254);
or U15692 (N_15692,N_15184,N_15022);
nor U15693 (N_15693,N_15200,N_15318);
nor U15694 (N_15694,N_15427,N_15393);
xnor U15695 (N_15695,N_15026,N_15437);
or U15696 (N_15696,N_15300,N_15192);
nand U15697 (N_15697,N_15342,N_15082);
xnor U15698 (N_15698,N_15077,N_15131);
or U15699 (N_15699,N_15314,N_15451);
nor U15700 (N_15700,N_15136,N_15465);
nor U15701 (N_15701,N_15056,N_15235);
nor U15702 (N_15702,N_15083,N_15115);
nor U15703 (N_15703,N_15114,N_15202);
nor U15704 (N_15704,N_15185,N_15259);
xnor U15705 (N_15705,N_15247,N_15159);
or U15706 (N_15706,N_15272,N_15416);
xor U15707 (N_15707,N_15405,N_15310);
nand U15708 (N_15708,N_15331,N_15174);
and U15709 (N_15709,N_15275,N_15061);
nand U15710 (N_15710,N_15299,N_15487);
and U15711 (N_15711,N_15382,N_15472);
or U15712 (N_15712,N_15302,N_15401);
xor U15713 (N_15713,N_15065,N_15445);
nand U15714 (N_15714,N_15400,N_15164);
xor U15715 (N_15715,N_15355,N_15099);
xnor U15716 (N_15716,N_15128,N_15045);
or U15717 (N_15717,N_15175,N_15474);
nor U15718 (N_15718,N_15255,N_15452);
nand U15719 (N_15719,N_15372,N_15453);
nand U15720 (N_15720,N_15239,N_15130);
xnor U15721 (N_15721,N_15271,N_15060);
or U15722 (N_15722,N_15217,N_15350);
nor U15723 (N_15723,N_15360,N_15009);
xor U15724 (N_15724,N_15428,N_15141);
xor U15725 (N_15725,N_15224,N_15470);
or U15726 (N_15726,N_15370,N_15348);
and U15727 (N_15727,N_15035,N_15260);
or U15728 (N_15728,N_15412,N_15423);
or U15729 (N_15729,N_15422,N_15207);
or U15730 (N_15730,N_15153,N_15287);
nand U15731 (N_15731,N_15362,N_15306);
nand U15732 (N_15732,N_15157,N_15052);
and U15733 (N_15733,N_15344,N_15391);
xnor U15734 (N_15734,N_15097,N_15285);
nor U15735 (N_15735,N_15238,N_15110);
and U15736 (N_15736,N_15102,N_15084);
nor U15737 (N_15737,N_15020,N_15273);
xnor U15738 (N_15738,N_15019,N_15333);
and U15739 (N_15739,N_15327,N_15213);
nand U15740 (N_15740,N_15378,N_15417);
or U15741 (N_15741,N_15469,N_15335);
or U15742 (N_15742,N_15100,N_15069);
or U15743 (N_15743,N_15033,N_15398);
and U15744 (N_15744,N_15397,N_15171);
or U15745 (N_15745,N_15482,N_15244);
or U15746 (N_15746,N_15491,N_15309);
and U15747 (N_15747,N_15010,N_15003);
or U15748 (N_15748,N_15492,N_15413);
nand U15749 (N_15749,N_15277,N_15029);
or U15750 (N_15750,N_15080,N_15048);
nand U15751 (N_15751,N_15266,N_15284);
nor U15752 (N_15752,N_15350,N_15049);
xor U15753 (N_15753,N_15175,N_15263);
and U15754 (N_15754,N_15215,N_15281);
or U15755 (N_15755,N_15214,N_15490);
nand U15756 (N_15756,N_15434,N_15116);
or U15757 (N_15757,N_15072,N_15352);
and U15758 (N_15758,N_15088,N_15446);
xor U15759 (N_15759,N_15383,N_15105);
xor U15760 (N_15760,N_15187,N_15438);
nand U15761 (N_15761,N_15363,N_15387);
nor U15762 (N_15762,N_15369,N_15436);
xnor U15763 (N_15763,N_15290,N_15097);
or U15764 (N_15764,N_15448,N_15025);
and U15765 (N_15765,N_15097,N_15292);
nand U15766 (N_15766,N_15148,N_15169);
or U15767 (N_15767,N_15317,N_15246);
nor U15768 (N_15768,N_15293,N_15496);
nor U15769 (N_15769,N_15289,N_15151);
and U15770 (N_15770,N_15356,N_15256);
nor U15771 (N_15771,N_15441,N_15156);
nor U15772 (N_15772,N_15472,N_15128);
nor U15773 (N_15773,N_15010,N_15493);
or U15774 (N_15774,N_15200,N_15015);
or U15775 (N_15775,N_15193,N_15467);
nand U15776 (N_15776,N_15239,N_15164);
xor U15777 (N_15777,N_15073,N_15339);
nand U15778 (N_15778,N_15488,N_15106);
nor U15779 (N_15779,N_15239,N_15038);
and U15780 (N_15780,N_15034,N_15028);
or U15781 (N_15781,N_15383,N_15412);
xor U15782 (N_15782,N_15127,N_15191);
or U15783 (N_15783,N_15023,N_15431);
nand U15784 (N_15784,N_15499,N_15243);
xor U15785 (N_15785,N_15359,N_15101);
and U15786 (N_15786,N_15474,N_15093);
nand U15787 (N_15787,N_15248,N_15085);
nand U15788 (N_15788,N_15490,N_15015);
nand U15789 (N_15789,N_15329,N_15048);
nor U15790 (N_15790,N_15352,N_15487);
nor U15791 (N_15791,N_15252,N_15480);
nand U15792 (N_15792,N_15369,N_15309);
and U15793 (N_15793,N_15273,N_15365);
and U15794 (N_15794,N_15463,N_15161);
nand U15795 (N_15795,N_15497,N_15045);
nor U15796 (N_15796,N_15150,N_15400);
xor U15797 (N_15797,N_15401,N_15195);
or U15798 (N_15798,N_15494,N_15467);
nand U15799 (N_15799,N_15407,N_15390);
and U15800 (N_15800,N_15279,N_15142);
or U15801 (N_15801,N_15393,N_15241);
nor U15802 (N_15802,N_15146,N_15238);
xnor U15803 (N_15803,N_15084,N_15250);
nand U15804 (N_15804,N_15270,N_15025);
nand U15805 (N_15805,N_15167,N_15442);
and U15806 (N_15806,N_15245,N_15184);
or U15807 (N_15807,N_15091,N_15230);
and U15808 (N_15808,N_15365,N_15341);
and U15809 (N_15809,N_15382,N_15309);
and U15810 (N_15810,N_15495,N_15025);
xnor U15811 (N_15811,N_15189,N_15382);
xor U15812 (N_15812,N_15142,N_15428);
and U15813 (N_15813,N_15217,N_15207);
xnor U15814 (N_15814,N_15210,N_15023);
nor U15815 (N_15815,N_15282,N_15074);
nand U15816 (N_15816,N_15102,N_15435);
xnor U15817 (N_15817,N_15456,N_15347);
nand U15818 (N_15818,N_15477,N_15055);
nor U15819 (N_15819,N_15401,N_15459);
or U15820 (N_15820,N_15112,N_15037);
xnor U15821 (N_15821,N_15430,N_15491);
nor U15822 (N_15822,N_15140,N_15328);
nor U15823 (N_15823,N_15284,N_15055);
or U15824 (N_15824,N_15110,N_15268);
and U15825 (N_15825,N_15114,N_15086);
nor U15826 (N_15826,N_15109,N_15304);
and U15827 (N_15827,N_15044,N_15199);
nand U15828 (N_15828,N_15062,N_15444);
and U15829 (N_15829,N_15016,N_15238);
xor U15830 (N_15830,N_15000,N_15066);
or U15831 (N_15831,N_15109,N_15236);
xnor U15832 (N_15832,N_15156,N_15380);
nor U15833 (N_15833,N_15011,N_15366);
nor U15834 (N_15834,N_15075,N_15255);
xnor U15835 (N_15835,N_15221,N_15123);
xor U15836 (N_15836,N_15273,N_15419);
or U15837 (N_15837,N_15017,N_15402);
xor U15838 (N_15838,N_15327,N_15057);
or U15839 (N_15839,N_15449,N_15323);
and U15840 (N_15840,N_15435,N_15080);
or U15841 (N_15841,N_15262,N_15178);
or U15842 (N_15842,N_15159,N_15201);
nand U15843 (N_15843,N_15431,N_15099);
nand U15844 (N_15844,N_15033,N_15221);
or U15845 (N_15845,N_15140,N_15176);
xor U15846 (N_15846,N_15012,N_15076);
or U15847 (N_15847,N_15475,N_15154);
and U15848 (N_15848,N_15016,N_15422);
and U15849 (N_15849,N_15207,N_15197);
nand U15850 (N_15850,N_15390,N_15027);
or U15851 (N_15851,N_15380,N_15418);
nand U15852 (N_15852,N_15253,N_15338);
nand U15853 (N_15853,N_15448,N_15469);
nand U15854 (N_15854,N_15010,N_15143);
and U15855 (N_15855,N_15033,N_15027);
nor U15856 (N_15856,N_15220,N_15242);
nand U15857 (N_15857,N_15097,N_15183);
and U15858 (N_15858,N_15297,N_15202);
or U15859 (N_15859,N_15466,N_15159);
nor U15860 (N_15860,N_15017,N_15331);
xnor U15861 (N_15861,N_15482,N_15412);
nor U15862 (N_15862,N_15472,N_15108);
nand U15863 (N_15863,N_15467,N_15286);
nand U15864 (N_15864,N_15272,N_15244);
or U15865 (N_15865,N_15048,N_15166);
and U15866 (N_15866,N_15126,N_15429);
nand U15867 (N_15867,N_15228,N_15241);
nor U15868 (N_15868,N_15422,N_15008);
xnor U15869 (N_15869,N_15194,N_15479);
nor U15870 (N_15870,N_15268,N_15351);
and U15871 (N_15871,N_15337,N_15181);
nand U15872 (N_15872,N_15093,N_15455);
nand U15873 (N_15873,N_15102,N_15027);
xor U15874 (N_15874,N_15211,N_15261);
xor U15875 (N_15875,N_15156,N_15273);
and U15876 (N_15876,N_15244,N_15339);
xnor U15877 (N_15877,N_15118,N_15038);
nor U15878 (N_15878,N_15265,N_15497);
xor U15879 (N_15879,N_15485,N_15213);
or U15880 (N_15880,N_15207,N_15004);
nor U15881 (N_15881,N_15326,N_15045);
nand U15882 (N_15882,N_15398,N_15478);
xnor U15883 (N_15883,N_15085,N_15252);
nor U15884 (N_15884,N_15059,N_15271);
nor U15885 (N_15885,N_15136,N_15011);
or U15886 (N_15886,N_15305,N_15008);
and U15887 (N_15887,N_15048,N_15246);
xnor U15888 (N_15888,N_15434,N_15047);
nor U15889 (N_15889,N_15382,N_15362);
nand U15890 (N_15890,N_15468,N_15266);
nor U15891 (N_15891,N_15445,N_15253);
nand U15892 (N_15892,N_15331,N_15437);
nor U15893 (N_15893,N_15395,N_15383);
xor U15894 (N_15894,N_15298,N_15477);
and U15895 (N_15895,N_15224,N_15352);
nor U15896 (N_15896,N_15270,N_15362);
or U15897 (N_15897,N_15380,N_15473);
or U15898 (N_15898,N_15268,N_15422);
or U15899 (N_15899,N_15438,N_15097);
and U15900 (N_15900,N_15060,N_15344);
xor U15901 (N_15901,N_15198,N_15477);
nand U15902 (N_15902,N_15223,N_15431);
or U15903 (N_15903,N_15366,N_15081);
nand U15904 (N_15904,N_15367,N_15317);
nand U15905 (N_15905,N_15082,N_15322);
xor U15906 (N_15906,N_15368,N_15043);
and U15907 (N_15907,N_15203,N_15250);
or U15908 (N_15908,N_15491,N_15144);
xnor U15909 (N_15909,N_15376,N_15495);
nand U15910 (N_15910,N_15106,N_15258);
or U15911 (N_15911,N_15253,N_15482);
xnor U15912 (N_15912,N_15272,N_15287);
xor U15913 (N_15913,N_15079,N_15308);
xor U15914 (N_15914,N_15434,N_15041);
nor U15915 (N_15915,N_15221,N_15433);
nor U15916 (N_15916,N_15402,N_15137);
nand U15917 (N_15917,N_15209,N_15016);
xnor U15918 (N_15918,N_15432,N_15317);
nor U15919 (N_15919,N_15290,N_15343);
nor U15920 (N_15920,N_15378,N_15496);
or U15921 (N_15921,N_15341,N_15019);
and U15922 (N_15922,N_15191,N_15126);
nand U15923 (N_15923,N_15146,N_15048);
xnor U15924 (N_15924,N_15248,N_15225);
nand U15925 (N_15925,N_15498,N_15206);
nand U15926 (N_15926,N_15212,N_15396);
and U15927 (N_15927,N_15475,N_15179);
nor U15928 (N_15928,N_15220,N_15233);
nand U15929 (N_15929,N_15067,N_15495);
and U15930 (N_15930,N_15083,N_15367);
nor U15931 (N_15931,N_15317,N_15161);
nor U15932 (N_15932,N_15000,N_15444);
xor U15933 (N_15933,N_15247,N_15194);
and U15934 (N_15934,N_15489,N_15169);
or U15935 (N_15935,N_15293,N_15192);
xnor U15936 (N_15936,N_15486,N_15341);
nand U15937 (N_15937,N_15081,N_15095);
and U15938 (N_15938,N_15340,N_15346);
xor U15939 (N_15939,N_15387,N_15262);
and U15940 (N_15940,N_15349,N_15443);
xor U15941 (N_15941,N_15128,N_15234);
or U15942 (N_15942,N_15218,N_15159);
and U15943 (N_15943,N_15490,N_15091);
nor U15944 (N_15944,N_15058,N_15465);
xnor U15945 (N_15945,N_15358,N_15414);
nand U15946 (N_15946,N_15392,N_15330);
xor U15947 (N_15947,N_15319,N_15414);
xor U15948 (N_15948,N_15333,N_15057);
nand U15949 (N_15949,N_15379,N_15289);
nor U15950 (N_15950,N_15488,N_15310);
xor U15951 (N_15951,N_15235,N_15400);
xor U15952 (N_15952,N_15228,N_15364);
or U15953 (N_15953,N_15147,N_15199);
or U15954 (N_15954,N_15344,N_15329);
and U15955 (N_15955,N_15444,N_15497);
and U15956 (N_15956,N_15396,N_15257);
nor U15957 (N_15957,N_15347,N_15300);
or U15958 (N_15958,N_15200,N_15487);
nor U15959 (N_15959,N_15008,N_15083);
nand U15960 (N_15960,N_15073,N_15368);
xnor U15961 (N_15961,N_15213,N_15492);
or U15962 (N_15962,N_15296,N_15474);
nor U15963 (N_15963,N_15494,N_15370);
or U15964 (N_15964,N_15439,N_15012);
nor U15965 (N_15965,N_15014,N_15106);
or U15966 (N_15966,N_15457,N_15046);
or U15967 (N_15967,N_15320,N_15488);
xnor U15968 (N_15968,N_15464,N_15240);
or U15969 (N_15969,N_15275,N_15482);
and U15970 (N_15970,N_15147,N_15079);
nor U15971 (N_15971,N_15212,N_15443);
or U15972 (N_15972,N_15172,N_15493);
xnor U15973 (N_15973,N_15294,N_15084);
xor U15974 (N_15974,N_15395,N_15190);
xor U15975 (N_15975,N_15013,N_15069);
nand U15976 (N_15976,N_15084,N_15413);
nand U15977 (N_15977,N_15374,N_15212);
or U15978 (N_15978,N_15248,N_15127);
xor U15979 (N_15979,N_15020,N_15308);
or U15980 (N_15980,N_15270,N_15349);
or U15981 (N_15981,N_15067,N_15442);
xnor U15982 (N_15982,N_15467,N_15029);
xnor U15983 (N_15983,N_15383,N_15283);
and U15984 (N_15984,N_15134,N_15090);
nand U15985 (N_15985,N_15313,N_15273);
and U15986 (N_15986,N_15217,N_15000);
and U15987 (N_15987,N_15415,N_15079);
nor U15988 (N_15988,N_15220,N_15180);
nor U15989 (N_15989,N_15390,N_15418);
and U15990 (N_15990,N_15005,N_15100);
and U15991 (N_15991,N_15179,N_15077);
nand U15992 (N_15992,N_15232,N_15150);
nor U15993 (N_15993,N_15003,N_15146);
nand U15994 (N_15994,N_15087,N_15162);
or U15995 (N_15995,N_15301,N_15472);
nor U15996 (N_15996,N_15450,N_15286);
xor U15997 (N_15997,N_15105,N_15333);
and U15998 (N_15998,N_15414,N_15405);
xor U15999 (N_15999,N_15017,N_15408);
nand U16000 (N_16000,N_15703,N_15964);
nand U16001 (N_16001,N_15979,N_15831);
or U16002 (N_16002,N_15578,N_15756);
nor U16003 (N_16003,N_15673,N_15502);
nor U16004 (N_16004,N_15670,N_15882);
xor U16005 (N_16005,N_15766,N_15661);
nand U16006 (N_16006,N_15637,N_15878);
nor U16007 (N_16007,N_15729,N_15892);
or U16008 (N_16008,N_15746,N_15697);
xnor U16009 (N_16009,N_15823,N_15995);
nand U16010 (N_16010,N_15508,N_15859);
and U16011 (N_16011,N_15903,N_15998);
and U16012 (N_16012,N_15790,N_15512);
nor U16013 (N_16013,N_15632,N_15686);
xnor U16014 (N_16014,N_15540,N_15574);
or U16015 (N_16015,N_15700,N_15664);
nand U16016 (N_16016,N_15658,N_15924);
and U16017 (N_16017,N_15590,N_15691);
nand U16018 (N_16018,N_15877,N_15610);
xor U16019 (N_16019,N_15707,N_15806);
xor U16020 (N_16020,N_15532,N_15941);
or U16021 (N_16021,N_15934,N_15730);
xnor U16022 (N_16022,N_15606,N_15744);
xor U16023 (N_16023,N_15844,N_15567);
xor U16024 (N_16024,N_15556,N_15526);
xnor U16025 (N_16025,N_15883,N_15791);
nand U16026 (N_16026,N_15951,N_15890);
and U16027 (N_16027,N_15737,N_15980);
and U16028 (N_16028,N_15856,N_15946);
and U16029 (N_16029,N_15555,N_15865);
and U16030 (N_16030,N_15937,N_15705);
nand U16031 (N_16031,N_15566,N_15564);
nand U16032 (N_16032,N_15679,N_15528);
nand U16033 (N_16033,N_15699,N_15863);
or U16034 (N_16034,N_15957,N_15548);
nor U16035 (N_16035,N_15602,N_15690);
xnor U16036 (N_16036,N_15503,N_15634);
or U16037 (N_16037,N_15816,N_15544);
and U16038 (N_16038,N_15620,N_15727);
nor U16039 (N_16039,N_15684,N_15666);
nor U16040 (N_16040,N_15693,N_15748);
nand U16041 (N_16041,N_15662,N_15994);
and U16042 (N_16042,N_15983,N_15612);
nor U16043 (N_16043,N_15820,N_15988);
and U16044 (N_16044,N_15802,N_15573);
nand U16045 (N_16045,N_15622,N_15971);
and U16046 (N_16046,N_15561,N_15959);
or U16047 (N_16047,N_15552,N_15507);
or U16048 (N_16048,N_15547,N_15631);
nand U16049 (N_16049,N_15529,N_15513);
or U16050 (N_16050,N_15663,N_15641);
or U16051 (N_16051,N_15696,N_15913);
and U16052 (N_16052,N_15589,N_15930);
and U16053 (N_16053,N_15685,N_15799);
and U16054 (N_16054,N_15682,N_15991);
nand U16055 (N_16055,N_15582,N_15519);
xor U16056 (N_16056,N_15769,N_15990);
or U16057 (N_16057,N_15947,N_15809);
and U16058 (N_16058,N_15617,N_15783);
nor U16059 (N_16059,N_15857,N_15592);
and U16060 (N_16060,N_15608,N_15553);
nor U16061 (N_16061,N_15905,N_15972);
or U16062 (N_16062,N_15710,N_15862);
or U16063 (N_16063,N_15948,N_15619);
and U16064 (N_16064,N_15889,N_15698);
nor U16065 (N_16065,N_15726,N_15918);
or U16066 (N_16066,N_15888,N_15736);
nand U16067 (N_16067,N_15757,N_15753);
xor U16068 (N_16068,N_15536,N_15542);
nor U16069 (N_16069,N_15656,N_15876);
nor U16070 (N_16070,N_15935,N_15628);
and U16071 (N_16071,N_15752,N_15843);
xnor U16072 (N_16072,N_15762,N_15525);
xnor U16073 (N_16073,N_15648,N_15909);
and U16074 (N_16074,N_15623,N_15600);
nand U16075 (N_16075,N_15928,N_15813);
or U16076 (N_16076,N_15694,N_15767);
nor U16077 (N_16077,N_15801,N_15645);
nor U16078 (N_16078,N_15789,N_15825);
or U16079 (N_16079,N_15683,N_15771);
xor U16080 (N_16080,N_15676,N_15961);
xnor U16081 (N_16081,N_15765,N_15659);
nand U16082 (N_16082,N_15982,N_15958);
xnor U16083 (N_16083,N_15939,N_15893);
nor U16084 (N_16084,N_15761,N_15795);
xor U16085 (N_16085,N_15524,N_15866);
nor U16086 (N_16086,N_15598,N_15772);
xnor U16087 (N_16087,N_15973,N_15559);
nand U16088 (N_16088,N_15601,N_15675);
xor U16089 (N_16089,N_15721,N_15792);
nand U16090 (N_16090,N_15635,N_15720);
xnor U16091 (N_16091,N_15902,N_15775);
xnor U16092 (N_16092,N_15840,N_15904);
and U16093 (N_16093,N_15569,N_15841);
or U16094 (N_16094,N_15558,N_15724);
and U16095 (N_16095,N_15560,N_15885);
nor U16096 (N_16096,N_15758,N_15846);
nand U16097 (N_16097,N_15695,N_15940);
nor U16098 (N_16098,N_15581,N_15916);
nor U16099 (N_16099,N_15618,N_15974);
and U16100 (N_16100,N_15510,N_15861);
or U16101 (N_16101,N_15504,N_15740);
and U16102 (N_16102,N_15652,N_15718);
and U16103 (N_16103,N_15938,N_15630);
and U16104 (N_16104,N_15917,N_15759);
or U16105 (N_16105,N_15845,N_15835);
nor U16106 (N_16106,N_15899,N_15749);
nor U16107 (N_16107,N_15599,N_15949);
nor U16108 (N_16108,N_15956,N_15945);
nand U16109 (N_16109,N_15704,N_15596);
or U16110 (N_16110,N_15836,N_15711);
and U16111 (N_16111,N_15869,N_15605);
nor U16112 (N_16112,N_15774,N_15760);
xor U16113 (N_16113,N_15797,N_15523);
nand U16114 (N_16114,N_15912,N_15807);
nand U16115 (N_16115,N_15960,N_15687);
and U16116 (N_16116,N_15585,N_15966);
and U16117 (N_16117,N_15868,N_15577);
nand U16118 (N_16118,N_15651,N_15516);
nor U16119 (N_16119,N_15588,N_15625);
xnor U16120 (N_16120,N_15531,N_15828);
nor U16121 (N_16121,N_15776,N_15576);
nand U16122 (N_16122,N_15665,N_15535);
nand U16123 (N_16123,N_15702,N_15647);
nor U16124 (N_16124,N_15901,N_15963);
xnor U16125 (N_16125,N_15847,N_15734);
xnor U16126 (N_16126,N_15900,N_15853);
nor U16127 (N_16127,N_15922,N_15688);
xor U16128 (N_16128,N_15713,N_15541);
and U16129 (N_16129,N_15874,N_15927);
and U16130 (N_16130,N_15739,N_15773);
nor U16131 (N_16131,N_15615,N_15650);
xnor U16132 (N_16132,N_15714,N_15796);
xnor U16133 (N_16133,N_15975,N_15649);
or U16134 (N_16134,N_15879,N_15978);
xor U16135 (N_16135,N_15591,N_15537);
xor U16136 (N_16136,N_15817,N_15826);
nor U16137 (N_16137,N_15921,N_15839);
nor U16138 (N_16138,N_15954,N_15914);
nand U16139 (N_16139,N_15613,N_15616);
and U16140 (N_16140,N_15514,N_15538);
and U16141 (N_16141,N_15875,N_15603);
or U16142 (N_16142,N_15633,N_15787);
xnor U16143 (N_16143,N_15587,N_15580);
and U16144 (N_16144,N_15763,N_15747);
or U16145 (N_16145,N_15815,N_15741);
nor U16146 (N_16146,N_15655,N_15554);
and U16147 (N_16147,N_15984,N_15867);
xnor U16148 (N_16148,N_15784,N_15669);
or U16149 (N_16149,N_15583,N_15881);
xor U16150 (N_16150,N_15723,N_15910);
nor U16151 (N_16151,N_15764,N_15621);
nor U16152 (N_16152,N_15584,N_15830);
nand U16153 (N_16153,N_15768,N_15906);
xor U16154 (N_16154,N_15855,N_15575);
and U16155 (N_16155,N_15919,N_15607);
xnor U16156 (N_16156,N_15871,N_15848);
nand U16157 (N_16157,N_15911,N_15672);
nand U16158 (N_16158,N_15572,N_15586);
nor U16159 (N_16159,N_15818,N_15798);
or U16160 (N_16160,N_15886,N_15829);
xor U16161 (N_16161,N_15671,N_15657);
nand U16162 (N_16162,N_15579,N_15770);
xnor U16163 (N_16163,N_15870,N_15933);
xnor U16164 (N_16164,N_15604,N_15880);
xor U16165 (N_16165,N_15915,N_15923);
and U16166 (N_16166,N_15745,N_15932);
or U16167 (N_16167,N_15895,N_15896);
xnor U16168 (N_16168,N_15668,N_15653);
and U16169 (N_16169,N_15522,N_15595);
or U16170 (N_16170,N_15725,N_15944);
xor U16171 (N_16171,N_15642,N_15987);
nand U16172 (N_16172,N_15810,N_15568);
or U16173 (N_16173,N_15680,N_15743);
or U16174 (N_16174,N_15955,N_15950);
or U16175 (N_16175,N_15952,N_15985);
nand U16176 (N_16176,N_15709,N_15969);
xnor U16177 (N_16177,N_15533,N_15785);
xnor U16178 (N_16178,N_15565,N_15786);
nor U16179 (N_16179,N_15640,N_15943);
or U16180 (N_16180,N_15735,N_15993);
and U16181 (N_16181,N_15803,N_15908);
and U16182 (N_16182,N_15965,N_15864);
or U16183 (N_16183,N_15543,N_15717);
and U16184 (N_16184,N_15728,N_15549);
or U16185 (N_16185,N_15624,N_15678);
nand U16186 (N_16186,N_15733,N_15997);
nand U16187 (N_16187,N_15755,N_15926);
or U16188 (N_16188,N_15777,N_15808);
xor U16189 (N_16189,N_15639,N_15722);
xor U16190 (N_16190,N_15597,N_15780);
nor U16191 (N_16191,N_15804,N_15731);
nor U16192 (N_16192,N_15689,N_15894);
nand U16193 (N_16193,N_15563,N_15692);
nor U16194 (N_16194,N_15636,N_15887);
xnor U16195 (N_16195,N_15819,N_15611);
nor U16196 (N_16196,N_15837,N_15550);
nor U16197 (N_16197,N_15712,N_15858);
xor U16198 (N_16198,N_15925,N_15701);
and U16199 (N_16199,N_15626,N_15931);
or U16200 (N_16200,N_15968,N_15842);
xor U16201 (N_16201,N_15517,N_15854);
nand U16202 (N_16202,N_15667,N_15833);
and U16203 (N_16203,N_15800,N_15545);
nor U16204 (N_16204,N_15838,N_15646);
nand U16205 (N_16205,N_15570,N_15614);
nor U16206 (N_16206,N_15505,N_15849);
nor U16207 (N_16207,N_15970,N_15716);
xnor U16208 (N_16208,N_15706,N_15509);
nand U16209 (N_16209,N_15778,N_15781);
and U16210 (N_16210,N_15521,N_15812);
nor U16211 (N_16211,N_15518,N_15821);
xnor U16212 (N_16212,N_15506,N_15681);
xor U16213 (N_16213,N_15793,N_15860);
or U16214 (N_16214,N_15738,N_15751);
or U16215 (N_16215,N_15593,N_15992);
or U16216 (N_16216,N_15708,N_15782);
nand U16217 (N_16217,N_15929,N_15873);
xnor U16218 (N_16218,N_15660,N_15557);
xor U16219 (N_16219,N_15609,N_15546);
and U16220 (N_16220,N_15967,N_15977);
nand U16221 (N_16221,N_15805,N_15907);
xor U16222 (N_16222,N_15539,N_15897);
nand U16223 (N_16223,N_15884,N_15953);
nand U16224 (N_16224,N_15515,N_15527);
and U16225 (N_16225,N_15822,N_15750);
or U16226 (N_16226,N_15824,N_15898);
or U16227 (N_16227,N_15936,N_15788);
nand U16228 (N_16228,N_15501,N_15534);
and U16229 (N_16229,N_15962,N_15571);
nor U16230 (N_16230,N_15779,N_15551);
or U16231 (N_16231,N_15719,N_15996);
and U16232 (N_16232,N_15794,N_15814);
xor U16233 (N_16233,N_15732,N_15638);
or U16234 (N_16234,N_15594,N_15999);
and U16235 (N_16235,N_15827,N_15643);
nor U16236 (N_16236,N_15715,N_15986);
nand U16237 (N_16237,N_15872,N_15742);
or U16238 (N_16238,N_15850,N_15852);
or U16239 (N_16239,N_15942,N_15976);
nor U16240 (N_16240,N_15832,N_15981);
or U16241 (N_16241,N_15754,N_15500);
or U16242 (N_16242,N_15834,N_15644);
nor U16243 (N_16243,N_15851,N_15511);
nor U16244 (N_16244,N_15891,N_15520);
nand U16245 (N_16245,N_15989,N_15654);
nor U16246 (N_16246,N_15674,N_15627);
xor U16247 (N_16247,N_15530,N_15629);
nor U16248 (N_16248,N_15677,N_15811);
nor U16249 (N_16249,N_15920,N_15562);
or U16250 (N_16250,N_15814,N_15907);
nand U16251 (N_16251,N_15661,N_15518);
and U16252 (N_16252,N_15987,N_15969);
nand U16253 (N_16253,N_15984,N_15838);
nor U16254 (N_16254,N_15827,N_15662);
or U16255 (N_16255,N_15707,N_15788);
nand U16256 (N_16256,N_15811,N_15931);
xor U16257 (N_16257,N_15510,N_15964);
or U16258 (N_16258,N_15795,N_15530);
and U16259 (N_16259,N_15986,N_15500);
xnor U16260 (N_16260,N_15876,N_15753);
nand U16261 (N_16261,N_15529,N_15868);
nor U16262 (N_16262,N_15737,N_15803);
or U16263 (N_16263,N_15823,N_15774);
xor U16264 (N_16264,N_15799,N_15742);
nor U16265 (N_16265,N_15728,N_15689);
and U16266 (N_16266,N_15990,N_15938);
nor U16267 (N_16267,N_15891,N_15680);
and U16268 (N_16268,N_15595,N_15978);
nand U16269 (N_16269,N_15534,N_15503);
and U16270 (N_16270,N_15794,N_15676);
and U16271 (N_16271,N_15705,N_15667);
and U16272 (N_16272,N_15692,N_15611);
nand U16273 (N_16273,N_15571,N_15760);
xor U16274 (N_16274,N_15589,N_15654);
or U16275 (N_16275,N_15533,N_15719);
nand U16276 (N_16276,N_15643,N_15587);
nand U16277 (N_16277,N_15779,N_15909);
and U16278 (N_16278,N_15779,N_15671);
or U16279 (N_16279,N_15657,N_15938);
or U16280 (N_16280,N_15808,N_15843);
nor U16281 (N_16281,N_15664,N_15651);
xor U16282 (N_16282,N_15535,N_15959);
or U16283 (N_16283,N_15522,N_15954);
or U16284 (N_16284,N_15813,N_15799);
or U16285 (N_16285,N_15701,N_15913);
nand U16286 (N_16286,N_15561,N_15992);
xor U16287 (N_16287,N_15576,N_15910);
xor U16288 (N_16288,N_15887,N_15513);
xor U16289 (N_16289,N_15918,N_15745);
and U16290 (N_16290,N_15862,N_15681);
nor U16291 (N_16291,N_15631,N_15538);
or U16292 (N_16292,N_15734,N_15677);
nand U16293 (N_16293,N_15923,N_15832);
nand U16294 (N_16294,N_15982,N_15984);
or U16295 (N_16295,N_15726,N_15777);
or U16296 (N_16296,N_15595,N_15720);
nor U16297 (N_16297,N_15782,N_15599);
nand U16298 (N_16298,N_15788,N_15950);
and U16299 (N_16299,N_15553,N_15765);
and U16300 (N_16300,N_15752,N_15523);
or U16301 (N_16301,N_15559,N_15697);
nor U16302 (N_16302,N_15924,N_15790);
nor U16303 (N_16303,N_15823,N_15700);
or U16304 (N_16304,N_15774,N_15532);
nor U16305 (N_16305,N_15845,N_15998);
and U16306 (N_16306,N_15825,N_15964);
nand U16307 (N_16307,N_15581,N_15530);
nor U16308 (N_16308,N_15625,N_15667);
and U16309 (N_16309,N_15515,N_15671);
and U16310 (N_16310,N_15631,N_15792);
xnor U16311 (N_16311,N_15623,N_15682);
xnor U16312 (N_16312,N_15651,N_15576);
nand U16313 (N_16313,N_15999,N_15795);
nand U16314 (N_16314,N_15701,N_15611);
xnor U16315 (N_16315,N_15854,N_15972);
and U16316 (N_16316,N_15546,N_15503);
xnor U16317 (N_16317,N_15551,N_15898);
nand U16318 (N_16318,N_15785,N_15830);
xnor U16319 (N_16319,N_15643,N_15978);
and U16320 (N_16320,N_15506,N_15891);
nor U16321 (N_16321,N_15930,N_15647);
nand U16322 (N_16322,N_15509,N_15977);
nand U16323 (N_16323,N_15973,N_15659);
xor U16324 (N_16324,N_15530,N_15977);
xor U16325 (N_16325,N_15679,N_15630);
or U16326 (N_16326,N_15659,N_15997);
nand U16327 (N_16327,N_15934,N_15700);
or U16328 (N_16328,N_15745,N_15674);
and U16329 (N_16329,N_15874,N_15627);
xor U16330 (N_16330,N_15803,N_15955);
nand U16331 (N_16331,N_15585,N_15718);
nand U16332 (N_16332,N_15529,N_15824);
or U16333 (N_16333,N_15956,N_15735);
nor U16334 (N_16334,N_15747,N_15506);
nor U16335 (N_16335,N_15912,N_15756);
xnor U16336 (N_16336,N_15850,N_15994);
nand U16337 (N_16337,N_15576,N_15719);
or U16338 (N_16338,N_15684,N_15695);
and U16339 (N_16339,N_15620,N_15907);
xor U16340 (N_16340,N_15679,N_15562);
nand U16341 (N_16341,N_15958,N_15822);
nor U16342 (N_16342,N_15523,N_15899);
xor U16343 (N_16343,N_15798,N_15676);
or U16344 (N_16344,N_15804,N_15672);
nand U16345 (N_16345,N_15678,N_15882);
and U16346 (N_16346,N_15621,N_15853);
nand U16347 (N_16347,N_15678,N_15516);
nand U16348 (N_16348,N_15805,N_15564);
nand U16349 (N_16349,N_15685,N_15862);
and U16350 (N_16350,N_15850,N_15795);
nor U16351 (N_16351,N_15843,N_15688);
and U16352 (N_16352,N_15777,N_15571);
or U16353 (N_16353,N_15992,N_15662);
nand U16354 (N_16354,N_15549,N_15599);
or U16355 (N_16355,N_15560,N_15805);
or U16356 (N_16356,N_15926,N_15533);
and U16357 (N_16357,N_15507,N_15854);
nand U16358 (N_16358,N_15755,N_15573);
or U16359 (N_16359,N_15661,N_15695);
and U16360 (N_16360,N_15594,N_15567);
and U16361 (N_16361,N_15515,N_15582);
and U16362 (N_16362,N_15783,N_15520);
xnor U16363 (N_16363,N_15945,N_15530);
or U16364 (N_16364,N_15635,N_15657);
and U16365 (N_16365,N_15691,N_15986);
xor U16366 (N_16366,N_15685,N_15980);
xor U16367 (N_16367,N_15881,N_15843);
and U16368 (N_16368,N_15706,N_15525);
xor U16369 (N_16369,N_15718,N_15940);
xor U16370 (N_16370,N_15885,N_15538);
nand U16371 (N_16371,N_15514,N_15686);
nor U16372 (N_16372,N_15915,N_15611);
xnor U16373 (N_16373,N_15814,N_15660);
and U16374 (N_16374,N_15523,N_15846);
nor U16375 (N_16375,N_15503,N_15984);
or U16376 (N_16376,N_15614,N_15897);
nand U16377 (N_16377,N_15574,N_15905);
nor U16378 (N_16378,N_15998,N_15718);
xnor U16379 (N_16379,N_15984,N_15888);
or U16380 (N_16380,N_15556,N_15615);
nand U16381 (N_16381,N_15616,N_15564);
nand U16382 (N_16382,N_15810,N_15933);
and U16383 (N_16383,N_15844,N_15924);
nor U16384 (N_16384,N_15550,N_15674);
xor U16385 (N_16385,N_15568,N_15500);
and U16386 (N_16386,N_15543,N_15599);
or U16387 (N_16387,N_15636,N_15695);
nand U16388 (N_16388,N_15959,N_15807);
or U16389 (N_16389,N_15734,N_15631);
nor U16390 (N_16390,N_15862,N_15572);
nand U16391 (N_16391,N_15834,N_15596);
xor U16392 (N_16392,N_15830,N_15904);
nor U16393 (N_16393,N_15804,N_15510);
nand U16394 (N_16394,N_15670,N_15909);
nand U16395 (N_16395,N_15600,N_15624);
xor U16396 (N_16396,N_15836,N_15799);
nor U16397 (N_16397,N_15651,N_15901);
and U16398 (N_16398,N_15519,N_15710);
and U16399 (N_16399,N_15736,N_15563);
and U16400 (N_16400,N_15695,N_15909);
nand U16401 (N_16401,N_15737,N_15853);
nor U16402 (N_16402,N_15553,N_15607);
or U16403 (N_16403,N_15868,N_15517);
and U16404 (N_16404,N_15542,N_15968);
nand U16405 (N_16405,N_15614,N_15982);
and U16406 (N_16406,N_15875,N_15876);
nand U16407 (N_16407,N_15721,N_15550);
nor U16408 (N_16408,N_15641,N_15705);
and U16409 (N_16409,N_15818,N_15566);
nor U16410 (N_16410,N_15762,N_15798);
nor U16411 (N_16411,N_15532,N_15947);
nand U16412 (N_16412,N_15684,N_15926);
nand U16413 (N_16413,N_15864,N_15760);
or U16414 (N_16414,N_15798,N_15989);
nand U16415 (N_16415,N_15852,N_15778);
xnor U16416 (N_16416,N_15819,N_15547);
and U16417 (N_16417,N_15783,N_15848);
and U16418 (N_16418,N_15901,N_15840);
and U16419 (N_16419,N_15514,N_15652);
nor U16420 (N_16420,N_15643,N_15814);
xnor U16421 (N_16421,N_15909,N_15855);
or U16422 (N_16422,N_15717,N_15826);
nand U16423 (N_16423,N_15654,N_15934);
and U16424 (N_16424,N_15777,N_15504);
nand U16425 (N_16425,N_15518,N_15857);
or U16426 (N_16426,N_15906,N_15970);
nand U16427 (N_16427,N_15977,N_15741);
or U16428 (N_16428,N_15653,N_15769);
nand U16429 (N_16429,N_15706,N_15942);
and U16430 (N_16430,N_15784,N_15906);
and U16431 (N_16431,N_15756,N_15555);
nor U16432 (N_16432,N_15780,N_15526);
or U16433 (N_16433,N_15758,N_15811);
nand U16434 (N_16434,N_15722,N_15809);
nor U16435 (N_16435,N_15895,N_15615);
and U16436 (N_16436,N_15817,N_15608);
or U16437 (N_16437,N_15584,N_15653);
and U16438 (N_16438,N_15610,N_15509);
or U16439 (N_16439,N_15936,N_15776);
nor U16440 (N_16440,N_15981,N_15756);
or U16441 (N_16441,N_15591,N_15989);
nor U16442 (N_16442,N_15664,N_15744);
and U16443 (N_16443,N_15526,N_15557);
nand U16444 (N_16444,N_15718,N_15653);
nand U16445 (N_16445,N_15720,N_15514);
nand U16446 (N_16446,N_15857,N_15657);
nor U16447 (N_16447,N_15670,N_15915);
or U16448 (N_16448,N_15630,N_15684);
xor U16449 (N_16449,N_15798,N_15698);
and U16450 (N_16450,N_15791,N_15821);
xor U16451 (N_16451,N_15780,N_15625);
and U16452 (N_16452,N_15999,N_15816);
xor U16453 (N_16453,N_15529,N_15676);
nand U16454 (N_16454,N_15501,N_15874);
xor U16455 (N_16455,N_15818,N_15626);
xnor U16456 (N_16456,N_15805,N_15634);
xor U16457 (N_16457,N_15734,N_15852);
nand U16458 (N_16458,N_15690,N_15736);
nand U16459 (N_16459,N_15993,N_15830);
xnor U16460 (N_16460,N_15600,N_15986);
and U16461 (N_16461,N_15713,N_15970);
xor U16462 (N_16462,N_15524,N_15785);
nand U16463 (N_16463,N_15758,N_15747);
or U16464 (N_16464,N_15712,N_15619);
nand U16465 (N_16465,N_15529,N_15723);
nand U16466 (N_16466,N_15827,N_15712);
nand U16467 (N_16467,N_15713,N_15654);
and U16468 (N_16468,N_15901,N_15835);
nand U16469 (N_16469,N_15669,N_15563);
nand U16470 (N_16470,N_15851,N_15799);
nand U16471 (N_16471,N_15811,N_15961);
xnor U16472 (N_16472,N_15641,N_15958);
and U16473 (N_16473,N_15977,N_15736);
and U16474 (N_16474,N_15946,N_15916);
nor U16475 (N_16475,N_15917,N_15774);
xnor U16476 (N_16476,N_15796,N_15711);
or U16477 (N_16477,N_15930,N_15870);
xor U16478 (N_16478,N_15724,N_15726);
nand U16479 (N_16479,N_15680,N_15580);
nand U16480 (N_16480,N_15999,N_15938);
and U16481 (N_16481,N_15832,N_15705);
nor U16482 (N_16482,N_15619,N_15682);
or U16483 (N_16483,N_15576,N_15760);
or U16484 (N_16484,N_15973,N_15758);
or U16485 (N_16485,N_15687,N_15500);
and U16486 (N_16486,N_15875,N_15640);
and U16487 (N_16487,N_15662,N_15544);
or U16488 (N_16488,N_15644,N_15761);
nor U16489 (N_16489,N_15654,N_15825);
or U16490 (N_16490,N_15639,N_15801);
nor U16491 (N_16491,N_15923,N_15699);
xnor U16492 (N_16492,N_15622,N_15802);
nor U16493 (N_16493,N_15881,N_15556);
and U16494 (N_16494,N_15713,N_15721);
nor U16495 (N_16495,N_15648,N_15890);
xnor U16496 (N_16496,N_15520,N_15525);
xor U16497 (N_16497,N_15820,N_15754);
and U16498 (N_16498,N_15840,N_15742);
or U16499 (N_16499,N_15842,N_15901);
nor U16500 (N_16500,N_16442,N_16486);
and U16501 (N_16501,N_16487,N_16025);
and U16502 (N_16502,N_16199,N_16120);
nand U16503 (N_16503,N_16488,N_16311);
nand U16504 (N_16504,N_16047,N_16080);
nand U16505 (N_16505,N_16164,N_16127);
or U16506 (N_16506,N_16467,N_16017);
or U16507 (N_16507,N_16182,N_16014);
and U16508 (N_16508,N_16102,N_16084);
and U16509 (N_16509,N_16307,N_16011);
or U16510 (N_16510,N_16093,N_16185);
xnor U16511 (N_16511,N_16172,N_16347);
xnor U16512 (N_16512,N_16207,N_16278);
nand U16513 (N_16513,N_16065,N_16188);
xor U16514 (N_16514,N_16323,N_16392);
nand U16515 (N_16515,N_16183,N_16063);
xor U16516 (N_16516,N_16133,N_16478);
xnor U16517 (N_16517,N_16411,N_16479);
nor U16518 (N_16518,N_16282,N_16138);
nand U16519 (N_16519,N_16213,N_16494);
nand U16520 (N_16520,N_16385,N_16053);
nand U16521 (N_16521,N_16175,N_16493);
nor U16522 (N_16522,N_16381,N_16137);
nor U16523 (N_16523,N_16443,N_16201);
xnor U16524 (N_16524,N_16285,N_16452);
nand U16525 (N_16525,N_16155,N_16372);
xnor U16526 (N_16526,N_16094,N_16167);
nand U16527 (N_16527,N_16223,N_16248);
nor U16528 (N_16528,N_16271,N_16058);
xnor U16529 (N_16529,N_16472,N_16499);
or U16530 (N_16530,N_16476,N_16444);
nor U16531 (N_16531,N_16163,N_16399);
xnor U16532 (N_16532,N_16460,N_16211);
or U16533 (N_16533,N_16422,N_16284);
and U16534 (N_16534,N_16024,N_16306);
nor U16535 (N_16535,N_16325,N_16335);
and U16536 (N_16536,N_16060,N_16121);
and U16537 (N_16537,N_16348,N_16131);
nor U16538 (N_16538,N_16032,N_16286);
nor U16539 (N_16539,N_16077,N_16222);
nor U16540 (N_16540,N_16464,N_16089);
nor U16541 (N_16541,N_16255,N_16148);
or U16542 (N_16542,N_16169,N_16268);
nor U16543 (N_16543,N_16289,N_16283);
nor U16544 (N_16544,N_16226,N_16152);
xor U16545 (N_16545,N_16237,N_16219);
or U16546 (N_16546,N_16018,N_16404);
xor U16547 (N_16547,N_16429,N_16477);
or U16548 (N_16548,N_16083,N_16132);
and U16549 (N_16549,N_16441,N_16022);
nand U16550 (N_16550,N_16458,N_16012);
xor U16551 (N_16551,N_16139,N_16350);
xnor U16552 (N_16552,N_16364,N_16468);
and U16553 (N_16553,N_16107,N_16326);
nor U16554 (N_16554,N_16100,N_16232);
nand U16555 (N_16555,N_16010,N_16360);
nor U16556 (N_16556,N_16426,N_16250);
and U16557 (N_16557,N_16016,N_16115);
or U16558 (N_16558,N_16075,N_16216);
or U16559 (N_16559,N_16496,N_16340);
and U16560 (N_16560,N_16143,N_16064);
nor U16561 (N_16561,N_16156,N_16240);
xor U16562 (N_16562,N_16407,N_16085);
nor U16563 (N_16563,N_16149,N_16346);
xor U16564 (N_16564,N_16124,N_16315);
nand U16565 (N_16565,N_16398,N_16170);
or U16566 (N_16566,N_16321,N_16101);
and U16567 (N_16567,N_16105,N_16489);
nand U16568 (N_16568,N_16186,N_16375);
xnor U16569 (N_16569,N_16179,N_16337);
and U16570 (N_16570,N_16174,N_16228);
nor U16571 (N_16571,N_16113,N_16136);
or U16572 (N_16572,N_16383,N_16266);
nor U16573 (N_16573,N_16056,N_16088);
or U16574 (N_16574,N_16313,N_16144);
or U16575 (N_16575,N_16236,N_16433);
nor U16576 (N_16576,N_16261,N_16153);
xnor U16577 (N_16577,N_16263,N_16424);
nand U16578 (N_16578,N_16081,N_16070);
or U16579 (N_16579,N_16457,N_16425);
or U16580 (N_16580,N_16427,N_16395);
nand U16581 (N_16581,N_16382,N_16449);
or U16582 (N_16582,N_16001,N_16008);
nand U16583 (N_16583,N_16078,N_16417);
and U16584 (N_16584,N_16006,N_16051);
nand U16585 (N_16585,N_16270,N_16414);
xnor U16586 (N_16586,N_16308,N_16106);
and U16587 (N_16587,N_16267,N_16480);
nor U16588 (N_16588,N_16402,N_16108);
nor U16589 (N_16589,N_16055,N_16459);
nor U16590 (N_16590,N_16481,N_16358);
nand U16591 (N_16591,N_16229,N_16123);
or U16592 (N_16592,N_16281,N_16320);
and U16593 (N_16593,N_16243,N_16303);
xnor U16594 (N_16594,N_16003,N_16373);
nor U16595 (N_16595,N_16082,N_16324);
and U16596 (N_16596,N_16187,N_16171);
nor U16597 (N_16597,N_16380,N_16387);
or U16598 (N_16598,N_16474,N_16368);
or U16599 (N_16599,N_16412,N_16419);
nor U16600 (N_16600,N_16334,N_16300);
nand U16601 (N_16601,N_16146,N_16463);
and U16602 (N_16602,N_16209,N_16439);
xnor U16603 (N_16603,N_16394,N_16142);
or U16604 (N_16604,N_16351,N_16379);
or U16605 (N_16605,N_16023,N_16341);
nand U16606 (N_16606,N_16253,N_16020);
nand U16607 (N_16607,N_16453,N_16231);
nand U16608 (N_16608,N_16297,N_16438);
or U16609 (N_16609,N_16252,N_16111);
xor U16610 (N_16610,N_16262,N_16114);
xnor U16611 (N_16611,N_16273,N_16059);
nand U16612 (N_16612,N_16147,N_16076);
and U16613 (N_16613,N_16196,N_16045);
nand U16614 (N_16614,N_16165,N_16052);
xnor U16615 (N_16615,N_16403,N_16420);
nor U16616 (N_16616,N_16469,N_16048);
and U16617 (N_16617,N_16354,N_16462);
xor U16618 (N_16618,N_16482,N_16450);
xnor U16619 (N_16619,N_16161,N_16362);
and U16620 (N_16620,N_16135,N_16004);
or U16621 (N_16621,N_16026,N_16035);
or U16622 (N_16622,N_16331,N_16365);
nand U16623 (N_16623,N_16272,N_16200);
nand U16624 (N_16624,N_16039,N_16212);
or U16625 (N_16625,N_16305,N_16432);
nand U16626 (N_16626,N_16269,N_16490);
and U16627 (N_16627,N_16409,N_16239);
and U16628 (N_16628,N_16396,N_16330);
nand U16629 (N_16629,N_16180,N_16233);
and U16630 (N_16630,N_16044,N_16030);
nand U16631 (N_16631,N_16264,N_16041);
and U16632 (N_16632,N_16062,N_16309);
xor U16633 (N_16633,N_16220,N_16069);
nand U16634 (N_16634,N_16483,N_16296);
nand U16635 (N_16635,N_16343,N_16224);
nor U16636 (N_16636,N_16314,N_16145);
and U16637 (N_16637,N_16386,N_16061);
xor U16638 (N_16638,N_16336,N_16319);
or U16639 (N_16639,N_16355,N_16430);
xnor U16640 (N_16640,N_16317,N_16234);
or U16641 (N_16641,N_16225,N_16254);
or U16642 (N_16642,N_16125,N_16349);
or U16643 (N_16643,N_16461,N_16166);
nand U16644 (N_16644,N_16293,N_16290);
nor U16645 (N_16645,N_16019,N_16318);
xor U16646 (N_16646,N_16190,N_16446);
and U16647 (N_16647,N_16130,N_16276);
or U16648 (N_16648,N_16208,N_16184);
and U16649 (N_16649,N_16277,N_16217);
or U16650 (N_16650,N_16162,N_16007);
xor U16651 (N_16651,N_16241,N_16181);
and U16652 (N_16652,N_16095,N_16333);
xnor U16653 (N_16653,N_16249,N_16344);
or U16654 (N_16654,N_16497,N_16258);
or U16655 (N_16655,N_16400,N_16377);
nor U16656 (N_16656,N_16265,N_16103);
nand U16657 (N_16657,N_16129,N_16040);
xnor U16658 (N_16658,N_16043,N_16384);
nand U16659 (N_16659,N_16000,N_16256);
xor U16660 (N_16660,N_16128,N_16310);
nor U16661 (N_16661,N_16072,N_16189);
nand U16662 (N_16662,N_16485,N_16437);
xor U16663 (N_16663,N_16339,N_16410);
or U16664 (N_16664,N_16436,N_16074);
nor U16665 (N_16665,N_16416,N_16110);
nand U16666 (N_16666,N_16079,N_16206);
nor U16667 (N_16667,N_16194,N_16345);
nor U16668 (N_16668,N_16096,N_16413);
xor U16669 (N_16669,N_16491,N_16238);
and U16670 (N_16670,N_16021,N_16098);
xor U16671 (N_16671,N_16423,N_16087);
nand U16672 (N_16672,N_16245,N_16328);
and U16673 (N_16673,N_16302,N_16291);
nand U16674 (N_16674,N_16119,N_16359);
or U16675 (N_16675,N_16140,N_16118);
and U16676 (N_16676,N_16090,N_16168);
xor U16677 (N_16677,N_16192,N_16390);
nor U16678 (N_16678,N_16104,N_16214);
xor U16679 (N_16679,N_16031,N_16203);
xor U16680 (N_16680,N_16246,N_16312);
or U16681 (N_16681,N_16455,N_16492);
xnor U16682 (N_16682,N_16391,N_16134);
nand U16683 (N_16683,N_16316,N_16299);
nand U16684 (N_16684,N_16401,N_16274);
nand U16685 (N_16685,N_16193,N_16295);
nand U16686 (N_16686,N_16397,N_16434);
nand U16687 (N_16687,N_16178,N_16498);
xnor U16688 (N_16688,N_16370,N_16050);
and U16689 (N_16689,N_16369,N_16091);
nor U16690 (N_16690,N_16418,N_16221);
or U16691 (N_16691,N_16099,N_16028);
and U16692 (N_16692,N_16210,N_16456);
or U16693 (N_16693,N_16197,N_16352);
and U16694 (N_16694,N_16366,N_16202);
nor U16695 (N_16695,N_16473,N_16195);
nand U16696 (N_16696,N_16475,N_16158);
nor U16697 (N_16697,N_16247,N_16154);
nor U16698 (N_16698,N_16205,N_16288);
nor U16699 (N_16699,N_16009,N_16371);
or U16700 (N_16700,N_16126,N_16471);
or U16701 (N_16701,N_16304,N_16329);
xnor U16702 (N_16702,N_16066,N_16431);
xnor U16703 (N_16703,N_16141,N_16160);
xor U16704 (N_16704,N_16036,N_16068);
xnor U16705 (N_16705,N_16374,N_16176);
nor U16706 (N_16706,N_16235,N_16367);
xnor U16707 (N_16707,N_16054,N_16279);
nand U16708 (N_16708,N_16071,N_16097);
nor U16709 (N_16709,N_16465,N_16230);
nand U16710 (N_16710,N_16405,N_16005);
nand U16711 (N_16711,N_16260,N_16173);
or U16712 (N_16712,N_16357,N_16033);
nor U16713 (N_16713,N_16151,N_16280);
xor U16714 (N_16714,N_16435,N_16198);
or U16715 (N_16715,N_16244,N_16484);
nor U16716 (N_16716,N_16092,N_16447);
or U16717 (N_16717,N_16159,N_16242);
and U16718 (N_16718,N_16013,N_16122);
or U16719 (N_16719,N_16037,N_16389);
and U16720 (N_16720,N_16470,N_16356);
nor U16721 (N_16721,N_16204,N_16495);
nor U16722 (N_16722,N_16448,N_16451);
nand U16723 (N_16723,N_16275,N_16428);
and U16724 (N_16724,N_16057,N_16322);
and U16725 (N_16725,N_16073,N_16257);
or U16726 (N_16726,N_16342,N_16116);
and U16727 (N_16727,N_16361,N_16421);
or U16728 (N_16728,N_16086,N_16287);
and U16729 (N_16729,N_16067,N_16015);
nor U16730 (N_16730,N_16406,N_16415);
and U16731 (N_16731,N_16027,N_16338);
and U16732 (N_16732,N_16046,N_16150);
xor U16733 (N_16733,N_16466,N_16294);
nand U16734 (N_16734,N_16112,N_16251);
or U16735 (N_16735,N_16049,N_16218);
or U16736 (N_16736,N_16227,N_16408);
or U16737 (N_16737,N_16215,N_16109);
and U16738 (N_16738,N_16292,N_16440);
xor U16739 (N_16739,N_16042,N_16301);
or U16740 (N_16740,N_16388,N_16454);
xnor U16741 (N_16741,N_16363,N_16445);
xnor U16742 (N_16742,N_16191,N_16378);
or U16743 (N_16743,N_16029,N_16332);
nand U16744 (N_16744,N_16177,N_16259);
xnor U16745 (N_16745,N_16002,N_16298);
xor U16746 (N_16746,N_16353,N_16038);
and U16747 (N_16747,N_16034,N_16117);
nand U16748 (N_16748,N_16327,N_16376);
nor U16749 (N_16749,N_16157,N_16393);
and U16750 (N_16750,N_16308,N_16280);
xnor U16751 (N_16751,N_16205,N_16442);
or U16752 (N_16752,N_16459,N_16222);
and U16753 (N_16753,N_16055,N_16023);
nor U16754 (N_16754,N_16023,N_16110);
or U16755 (N_16755,N_16156,N_16089);
or U16756 (N_16756,N_16291,N_16296);
and U16757 (N_16757,N_16347,N_16042);
nor U16758 (N_16758,N_16325,N_16113);
nor U16759 (N_16759,N_16173,N_16433);
and U16760 (N_16760,N_16225,N_16439);
nor U16761 (N_16761,N_16427,N_16011);
nor U16762 (N_16762,N_16483,N_16281);
and U16763 (N_16763,N_16016,N_16490);
or U16764 (N_16764,N_16213,N_16146);
xor U16765 (N_16765,N_16208,N_16163);
nand U16766 (N_16766,N_16378,N_16145);
xor U16767 (N_16767,N_16336,N_16146);
and U16768 (N_16768,N_16016,N_16485);
xor U16769 (N_16769,N_16446,N_16143);
xnor U16770 (N_16770,N_16461,N_16239);
nand U16771 (N_16771,N_16093,N_16159);
xnor U16772 (N_16772,N_16277,N_16043);
nor U16773 (N_16773,N_16194,N_16410);
xor U16774 (N_16774,N_16230,N_16193);
nand U16775 (N_16775,N_16149,N_16104);
nand U16776 (N_16776,N_16195,N_16461);
xor U16777 (N_16777,N_16255,N_16454);
and U16778 (N_16778,N_16064,N_16059);
and U16779 (N_16779,N_16270,N_16057);
or U16780 (N_16780,N_16073,N_16211);
or U16781 (N_16781,N_16219,N_16287);
nor U16782 (N_16782,N_16125,N_16422);
and U16783 (N_16783,N_16060,N_16011);
nand U16784 (N_16784,N_16287,N_16137);
or U16785 (N_16785,N_16489,N_16118);
and U16786 (N_16786,N_16293,N_16219);
xnor U16787 (N_16787,N_16101,N_16121);
nand U16788 (N_16788,N_16288,N_16282);
nor U16789 (N_16789,N_16093,N_16336);
xor U16790 (N_16790,N_16494,N_16205);
or U16791 (N_16791,N_16062,N_16230);
xor U16792 (N_16792,N_16329,N_16308);
nand U16793 (N_16793,N_16376,N_16072);
or U16794 (N_16794,N_16289,N_16374);
nand U16795 (N_16795,N_16021,N_16311);
nand U16796 (N_16796,N_16197,N_16003);
nand U16797 (N_16797,N_16352,N_16465);
nand U16798 (N_16798,N_16485,N_16214);
or U16799 (N_16799,N_16374,N_16462);
and U16800 (N_16800,N_16346,N_16150);
xor U16801 (N_16801,N_16169,N_16112);
xnor U16802 (N_16802,N_16448,N_16099);
nor U16803 (N_16803,N_16489,N_16325);
and U16804 (N_16804,N_16110,N_16392);
nand U16805 (N_16805,N_16192,N_16222);
nor U16806 (N_16806,N_16492,N_16486);
and U16807 (N_16807,N_16312,N_16370);
xnor U16808 (N_16808,N_16305,N_16395);
and U16809 (N_16809,N_16403,N_16152);
and U16810 (N_16810,N_16149,N_16427);
xnor U16811 (N_16811,N_16084,N_16260);
xor U16812 (N_16812,N_16289,N_16366);
or U16813 (N_16813,N_16099,N_16135);
xnor U16814 (N_16814,N_16421,N_16319);
xnor U16815 (N_16815,N_16062,N_16045);
xnor U16816 (N_16816,N_16104,N_16150);
xnor U16817 (N_16817,N_16079,N_16322);
nor U16818 (N_16818,N_16467,N_16273);
nand U16819 (N_16819,N_16494,N_16087);
and U16820 (N_16820,N_16432,N_16028);
and U16821 (N_16821,N_16208,N_16444);
and U16822 (N_16822,N_16017,N_16407);
nand U16823 (N_16823,N_16471,N_16448);
xnor U16824 (N_16824,N_16106,N_16175);
nand U16825 (N_16825,N_16105,N_16212);
or U16826 (N_16826,N_16189,N_16125);
nand U16827 (N_16827,N_16340,N_16326);
or U16828 (N_16828,N_16087,N_16093);
nor U16829 (N_16829,N_16408,N_16328);
nand U16830 (N_16830,N_16346,N_16355);
xor U16831 (N_16831,N_16041,N_16488);
or U16832 (N_16832,N_16271,N_16474);
nand U16833 (N_16833,N_16293,N_16042);
and U16834 (N_16834,N_16491,N_16269);
xor U16835 (N_16835,N_16162,N_16176);
xor U16836 (N_16836,N_16116,N_16480);
nor U16837 (N_16837,N_16492,N_16208);
xnor U16838 (N_16838,N_16432,N_16473);
xor U16839 (N_16839,N_16086,N_16293);
nand U16840 (N_16840,N_16054,N_16497);
nand U16841 (N_16841,N_16428,N_16097);
xor U16842 (N_16842,N_16223,N_16310);
xor U16843 (N_16843,N_16151,N_16138);
or U16844 (N_16844,N_16156,N_16182);
and U16845 (N_16845,N_16363,N_16047);
and U16846 (N_16846,N_16263,N_16422);
nand U16847 (N_16847,N_16164,N_16029);
or U16848 (N_16848,N_16481,N_16178);
or U16849 (N_16849,N_16427,N_16226);
nand U16850 (N_16850,N_16192,N_16422);
xnor U16851 (N_16851,N_16344,N_16486);
nand U16852 (N_16852,N_16404,N_16373);
and U16853 (N_16853,N_16085,N_16470);
nand U16854 (N_16854,N_16112,N_16247);
or U16855 (N_16855,N_16028,N_16304);
or U16856 (N_16856,N_16297,N_16395);
or U16857 (N_16857,N_16473,N_16154);
nand U16858 (N_16858,N_16115,N_16251);
or U16859 (N_16859,N_16329,N_16273);
xnor U16860 (N_16860,N_16259,N_16485);
nor U16861 (N_16861,N_16215,N_16488);
and U16862 (N_16862,N_16211,N_16035);
nor U16863 (N_16863,N_16161,N_16077);
or U16864 (N_16864,N_16018,N_16294);
or U16865 (N_16865,N_16071,N_16409);
nand U16866 (N_16866,N_16022,N_16272);
and U16867 (N_16867,N_16169,N_16391);
nor U16868 (N_16868,N_16377,N_16019);
nor U16869 (N_16869,N_16383,N_16028);
xor U16870 (N_16870,N_16017,N_16491);
xnor U16871 (N_16871,N_16087,N_16490);
xnor U16872 (N_16872,N_16392,N_16211);
xnor U16873 (N_16873,N_16243,N_16370);
xor U16874 (N_16874,N_16084,N_16473);
or U16875 (N_16875,N_16403,N_16053);
and U16876 (N_16876,N_16189,N_16291);
nor U16877 (N_16877,N_16390,N_16037);
or U16878 (N_16878,N_16167,N_16156);
or U16879 (N_16879,N_16291,N_16142);
and U16880 (N_16880,N_16185,N_16023);
and U16881 (N_16881,N_16448,N_16114);
or U16882 (N_16882,N_16036,N_16273);
nor U16883 (N_16883,N_16086,N_16084);
and U16884 (N_16884,N_16239,N_16355);
and U16885 (N_16885,N_16454,N_16445);
or U16886 (N_16886,N_16253,N_16091);
xnor U16887 (N_16887,N_16250,N_16463);
or U16888 (N_16888,N_16225,N_16445);
or U16889 (N_16889,N_16166,N_16418);
and U16890 (N_16890,N_16488,N_16418);
xnor U16891 (N_16891,N_16320,N_16232);
nand U16892 (N_16892,N_16095,N_16404);
nand U16893 (N_16893,N_16295,N_16276);
nor U16894 (N_16894,N_16118,N_16405);
xnor U16895 (N_16895,N_16164,N_16316);
or U16896 (N_16896,N_16384,N_16161);
xnor U16897 (N_16897,N_16353,N_16067);
or U16898 (N_16898,N_16187,N_16483);
nor U16899 (N_16899,N_16150,N_16085);
and U16900 (N_16900,N_16443,N_16410);
and U16901 (N_16901,N_16366,N_16276);
or U16902 (N_16902,N_16027,N_16444);
or U16903 (N_16903,N_16145,N_16170);
or U16904 (N_16904,N_16033,N_16025);
xnor U16905 (N_16905,N_16175,N_16480);
and U16906 (N_16906,N_16150,N_16024);
or U16907 (N_16907,N_16126,N_16468);
and U16908 (N_16908,N_16480,N_16039);
or U16909 (N_16909,N_16406,N_16445);
or U16910 (N_16910,N_16284,N_16403);
nor U16911 (N_16911,N_16037,N_16252);
nand U16912 (N_16912,N_16138,N_16025);
xnor U16913 (N_16913,N_16011,N_16461);
and U16914 (N_16914,N_16458,N_16110);
xnor U16915 (N_16915,N_16347,N_16230);
and U16916 (N_16916,N_16276,N_16193);
nand U16917 (N_16917,N_16415,N_16007);
nand U16918 (N_16918,N_16173,N_16215);
and U16919 (N_16919,N_16125,N_16382);
and U16920 (N_16920,N_16263,N_16477);
nand U16921 (N_16921,N_16110,N_16319);
nand U16922 (N_16922,N_16027,N_16340);
xor U16923 (N_16923,N_16484,N_16263);
nor U16924 (N_16924,N_16178,N_16148);
and U16925 (N_16925,N_16486,N_16428);
nor U16926 (N_16926,N_16363,N_16349);
or U16927 (N_16927,N_16228,N_16001);
or U16928 (N_16928,N_16210,N_16319);
xor U16929 (N_16929,N_16113,N_16370);
nand U16930 (N_16930,N_16336,N_16044);
and U16931 (N_16931,N_16373,N_16120);
nand U16932 (N_16932,N_16165,N_16203);
nor U16933 (N_16933,N_16041,N_16025);
nor U16934 (N_16934,N_16247,N_16130);
nor U16935 (N_16935,N_16449,N_16478);
and U16936 (N_16936,N_16307,N_16317);
nor U16937 (N_16937,N_16467,N_16176);
nand U16938 (N_16938,N_16167,N_16375);
or U16939 (N_16939,N_16089,N_16123);
nand U16940 (N_16940,N_16035,N_16304);
or U16941 (N_16941,N_16477,N_16086);
or U16942 (N_16942,N_16031,N_16320);
nor U16943 (N_16943,N_16242,N_16186);
nand U16944 (N_16944,N_16194,N_16100);
xnor U16945 (N_16945,N_16332,N_16180);
nor U16946 (N_16946,N_16119,N_16154);
or U16947 (N_16947,N_16160,N_16318);
and U16948 (N_16948,N_16236,N_16388);
nor U16949 (N_16949,N_16290,N_16440);
and U16950 (N_16950,N_16369,N_16056);
xor U16951 (N_16951,N_16479,N_16482);
nand U16952 (N_16952,N_16135,N_16286);
nand U16953 (N_16953,N_16084,N_16241);
and U16954 (N_16954,N_16048,N_16068);
nor U16955 (N_16955,N_16287,N_16292);
nand U16956 (N_16956,N_16384,N_16284);
xnor U16957 (N_16957,N_16395,N_16462);
and U16958 (N_16958,N_16381,N_16385);
nand U16959 (N_16959,N_16359,N_16214);
xnor U16960 (N_16960,N_16371,N_16361);
xor U16961 (N_16961,N_16101,N_16009);
or U16962 (N_16962,N_16215,N_16004);
and U16963 (N_16963,N_16329,N_16376);
nor U16964 (N_16964,N_16479,N_16477);
nor U16965 (N_16965,N_16378,N_16007);
or U16966 (N_16966,N_16493,N_16191);
xnor U16967 (N_16967,N_16253,N_16015);
or U16968 (N_16968,N_16312,N_16341);
xor U16969 (N_16969,N_16072,N_16006);
or U16970 (N_16970,N_16313,N_16152);
nand U16971 (N_16971,N_16175,N_16208);
and U16972 (N_16972,N_16126,N_16403);
and U16973 (N_16973,N_16426,N_16181);
nor U16974 (N_16974,N_16086,N_16325);
or U16975 (N_16975,N_16416,N_16137);
or U16976 (N_16976,N_16282,N_16073);
and U16977 (N_16977,N_16169,N_16087);
and U16978 (N_16978,N_16153,N_16097);
xor U16979 (N_16979,N_16285,N_16255);
xor U16980 (N_16980,N_16382,N_16160);
or U16981 (N_16981,N_16176,N_16297);
nor U16982 (N_16982,N_16198,N_16387);
nor U16983 (N_16983,N_16356,N_16397);
nand U16984 (N_16984,N_16160,N_16196);
nor U16985 (N_16985,N_16078,N_16330);
xor U16986 (N_16986,N_16246,N_16089);
nand U16987 (N_16987,N_16260,N_16073);
nor U16988 (N_16988,N_16453,N_16016);
nand U16989 (N_16989,N_16312,N_16159);
nor U16990 (N_16990,N_16187,N_16271);
nor U16991 (N_16991,N_16333,N_16316);
nand U16992 (N_16992,N_16207,N_16391);
xor U16993 (N_16993,N_16196,N_16301);
and U16994 (N_16994,N_16109,N_16308);
nor U16995 (N_16995,N_16491,N_16439);
nand U16996 (N_16996,N_16292,N_16488);
and U16997 (N_16997,N_16021,N_16235);
nor U16998 (N_16998,N_16127,N_16182);
or U16999 (N_16999,N_16184,N_16439);
nand U17000 (N_17000,N_16796,N_16857);
and U17001 (N_17001,N_16696,N_16587);
and U17002 (N_17002,N_16554,N_16647);
nand U17003 (N_17003,N_16518,N_16788);
nor U17004 (N_17004,N_16506,N_16827);
nand U17005 (N_17005,N_16598,N_16714);
nand U17006 (N_17006,N_16921,N_16502);
and U17007 (N_17007,N_16627,N_16971);
nor U17008 (N_17008,N_16586,N_16637);
nand U17009 (N_17009,N_16806,N_16922);
xor U17010 (N_17010,N_16540,N_16764);
nand U17011 (N_17011,N_16625,N_16626);
or U17012 (N_17012,N_16617,N_16869);
nand U17013 (N_17013,N_16670,N_16831);
nand U17014 (N_17014,N_16526,N_16679);
nand U17015 (N_17015,N_16755,N_16507);
and U17016 (N_17016,N_16754,N_16903);
nor U17017 (N_17017,N_16577,N_16636);
nand U17018 (N_17018,N_16673,N_16988);
and U17019 (N_17019,N_16942,N_16720);
nand U17020 (N_17020,N_16646,N_16551);
nor U17021 (N_17021,N_16773,N_16835);
xnor U17022 (N_17022,N_16578,N_16564);
xor U17023 (N_17023,N_16735,N_16889);
and U17024 (N_17024,N_16633,N_16976);
and U17025 (N_17025,N_16628,N_16880);
nand U17026 (N_17026,N_16571,N_16594);
nand U17027 (N_17027,N_16907,N_16891);
or U17028 (N_17028,N_16836,N_16730);
nand U17029 (N_17029,N_16808,N_16757);
xor U17030 (N_17030,N_16860,N_16684);
nand U17031 (N_17031,N_16810,N_16814);
nor U17032 (N_17032,N_16709,N_16590);
nand U17033 (N_17033,N_16951,N_16722);
or U17034 (N_17034,N_16794,N_16665);
nand U17035 (N_17035,N_16917,N_16803);
nor U17036 (N_17036,N_16642,N_16568);
nand U17037 (N_17037,N_16800,N_16783);
and U17038 (N_17038,N_16592,N_16708);
and U17039 (N_17039,N_16556,N_16525);
xnor U17040 (N_17040,N_16731,N_16542);
nor U17041 (N_17041,N_16774,N_16639);
and U17042 (N_17042,N_16521,N_16789);
nor U17043 (N_17043,N_16572,N_16842);
or U17044 (N_17044,N_16919,N_16671);
nor U17045 (N_17045,N_16759,N_16784);
and U17046 (N_17046,N_16999,N_16772);
xor U17047 (N_17047,N_16563,N_16741);
nor U17048 (N_17048,N_16736,N_16823);
nor U17049 (N_17049,N_16828,N_16939);
or U17050 (N_17050,N_16574,N_16591);
xnor U17051 (N_17051,N_16698,N_16729);
and U17052 (N_17052,N_16538,N_16992);
nand U17053 (N_17053,N_16977,N_16983);
nand U17054 (N_17054,N_16516,N_16885);
nand U17055 (N_17055,N_16858,N_16848);
nor U17056 (N_17056,N_16900,N_16974);
or U17057 (N_17057,N_16717,N_16593);
and U17058 (N_17058,N_16995,N_16632);
nor U17059 (N_17059,N_16712,N_16896);
and U17060 (N_17060,N_16873,N_16524);
and U17061 (N_17061,N_16600,N_16535);
nand U17062 (N_17062,N_16685,N_16510);
or U17063 (N_17063,N_16547,N_16982);
nand U17064 (N_17064,N_16514,N_16719);
nand U17065 (N_17065,N_16887,N_16747);
xor U17066 (N_17066,N_16513,N_16654);
xnor U17067 (N_17067,N_16904,N_16641);
or U17068 (N_17068,N_16902,N_16840);
or U17069 (N_17069,N_16989,N_16689);
and U17070 (N_17070,N_16865,N_16669);
xor U17071 (N_17071,N_16854,N_16649);
or U17072 (N_17072,N_16519,N_16924);
or U17073 (N_17073,N_16933,N_16692);
and U17074 (N_17074,N_16541,N_16972);
nand U17075 (N_17075,N_16565,N_16753);
nor U17076 (N_17076,N_16718,N_16527);
and U17077 (N_17077,N_16737,N_16756);
and U17078 (N_17078,N_16648,N_16997);
and U17079 (N_17079,N_16686,N_16599);
nor U17080 (N_17080,N_16515,N_16804);
xor U17081 (N_17081,N_16931,N_16560);
nand U17082 (N_17082,N_16875,N_16769);
nor U17083 (N_17083,N_16603,N_16812);
or U17084 (N_17084,N_16901,N_16844);
nor U17085 (N_17085,N_16793,N_16726);
nand U17086 (N_17086,N_16613,N_16956);
nor U17087 (N_17087,N_16978,N_16659);
nor U17088 (N_17088,N_16782,N_16611);
and U17089 (N_17089,N_16703,N_16706);
xnor U17090 (N_17090,N_16604,N_16734);
nand U17091 (N_17091,N_16792,N_16853);
or U17092 (N_17092,N_16781,N_16713);
xor U17093 (N_17093,N_16601,N_16512);
nor U17094 (N_17094,N_16596,N_16877);
nand U17095 (N_17095,N_16771,N_16915);
nor U17096 (N_17096,N_16562,N_16655);
xnor U17097 (N_17097,N_16935,N_16605);
and U17098 (N_17098,N_16878,N_16528);
nor U17099 (N_17099,N_16602,N_16711);
or U17100 (N_17100,N_16850,N_16943);
or U17101 (N_17101,N_16595,N_16573);
and U17102 (N_17102,N_16728,N_16807);
or U17103 (N_17103,N_16813,N_16855);
xor U17104 (N_17104,N_16621,N_16926);
and U17105 (N_17105,N_16966,N_16797);
xnor U17106 (N_17106,N_16824,N_16895);
and U17107 (N_17107,N_16536,N_16707);
or U17108 (N_17108,N_16964,N_16624);
xnor U17109 (N_17109,N_16969,N_16583);
or U17110 (N_17110,N_16963,N_16959);
nand U17111 (N_17111,N_16911,N_16868);
and U17112 (N_17112,N_16748,N_16843);
nand U17113 (N_17113,N_16890,N_16623);
xor U17114 (N_17114,N_16745,N_16967);
or U17115 (N_17115,N_16746,N_16763);
nand U17116 (N_17116,N_16805,N_16677);
or U17117 (N_17117,N_16545,N_16606);
xor U17118 (N_17118,N_16879,N_16607);
xor U17119 (N_17119,N_16790,N_16761);
or U17120 (N_17120,N_16973,N_16894);
or U17121 (N_17121,N_16682,N_16704);
nand U17122 (N_17122,N_16996,N_16899);
xor U17123 (N_17123,N_16775,N_16839);
xnor U17124 (N_17124,N_16653,N_16630);
xnor U17125 (N_17125,N_16744,N_16916);
nand U17126 (N_17126,N_16762,N_16866);
nand U17127 (N_17127,N_16936,N_16576);
xnor U17128 (N_17128,N_16534,N_16662);
nor U17129 (N_17129,N_16929,N_16768);
and U17130 (N_17130,N_16791,N_16566);
nor U17131 (N_17131,N_16511,N_16913);
nor U17132 (N_17132,N_16851,N_16838);
or U17133 (N_17133,N_16680,N_16867);
xor U17134 (N_17134,N_16618,N_16888);
and U17135 (N_17135,N_16520,N_16581);
nor U17136 (N_17136,N_16892,N_16683);
nor U17137 (N_17137,N_16923,N_16897);
nor U17138 (N_17138,N_16691,N_16883);
nand U17139 (N_17139,N_16819,N_16862);
and U17140 (N_17140,N_16643,N_16955);
and U17141 (N_17141,N_16946,N_16693);
xnor U17142 (N_17142,N_16588,N_16553);
xor U17143 (N_17143,N_16993,N_16830);
or U17144 (N_17144,N_16767,N_16950);
or U17145 (N_17145,N_16652,N_16859);
xnor U17146 (N_17146,N_16597,N_16622);
and U17147 (N_17147,N_16635,N_16777);
xnor U17148 (N_17148,N_16700,N_16531);
nor U17149 (N_17149,N_16539,N_16998);
or U17150 (N_17150,N_16817,N_16522);
xnor U17151 (N_17151,N_16620,N_16871);
nand U17152 (N_17152,N_16905,N_16750);
nor U17153 (N_17153,N_16957,N_16953);
nor U17154 (N_17154,N_16954,N_16852);
nor U17155 (N_17155,N_16765,N_16561);
nor U17156 (N_17156,N_16987,N_16668);
or U17157 (N_17157,N_16616,N_16508);
nand U17158 (N_17158,N_16610,N_16766);
and U17159 (N_17159,N_16811,N_16650);
and U17160 (N_17160,N_16886,N_16723);
or U17161 (N_17161,N_16785,N_16544);
nand U17162 (N_17162,N_16701,N_16920);
nand U17163 (N_17163,N_16975,N_16795);
and U17164 (N_17164,N_16697,N_16930);
nand U17165 (N_17165,N_16970,N_16820);
and U17166 (N_17166,N_16874,N_16845);
xor U17167 (N_17167,N_16501,N_16629);
and U17168 (N_17168,N_16825,N_16779);
xnor U17169 (N_17169,N_16558,N_16523);
xor U17170 (N_17170,N_16833,N_16965);
and U17171 (N_17171,N_16517,N_16849);
xor U17172 (N_17172,N_16914,N_16674);
xor U17173 (N_17173,N_16826,N_16656);
or U17174 (N_17174,N_16552,N_16958);
and U17175 (N_17175,N_16509,N_16580);
or U17176 (N_17176,N_16944,N_16631);
nand U17177 (N_17177,N_16529,N_16846);
xor U17178 (N_17178,N_16898,N_16615);
nand U17179 (N_17179,N_16694,N_16612);
nor U17180 (N_17180,N_16688,N_16585);
and U17181 (N_17181,N_16818,N_16881);
nand U17182 (N_17182,N_16530,N_16861);
or U17183 (N_17183,N_16947,N_16678);
xnor U17184 (N_17184,N_16733,N_16945);
nand U17185 (N_17185,N_16882,N_16934);
or U17186 (N_17186,N_16909,N_16687);
and U17187 (N_17187,N_16780,N_16822);
xor U17188 (N_17188,N_16608,N_16940);
and U17189 (N_17189,N_16856,N_16742);
nand U17190 (N_17190,N_16990,N_16546);
xnor U17191 (N_17191,N_16979,N_16918);
and U17192 (N_17192,N_16725,N_16864);
and U17193 (N_17193,N_16834,N_16821);
xor U17194 (N_17194,N_16815,N_16681);
and U17195 (N_17195,N_16863,N_16575);
xnor U17196 (N_17196,N_16644,N_16645);
nand U17197 (N_17197,N_16938,N_16609);
or U17198 (N_17198,N_16941,N_16787);
and U17199 (N_17199,N_16666,N_16980);
or U17200 (N_17200,N_16500,N_16721);
nand U17201 (N_17201,N_16724,N_16664);
nand U17202 (N_17202,N_16567,N_16555);
and U17203 (N_17203,N_16778,N_16799);
nand U17204 (N_17204,N_16960,N_16657);
nor U17205 (N_17205,N_16695,N_16537);
or U17206 (N_17206,N_16760,N_16893);
nor U17207 (N_17207,N_16816,N_16504);
or U17208 (N_17208,N_16667,N_16925);
nand U17209 (N_17209,N_16569,N_16749);
nand U17210 (N_17210,N_16829,N_16884);
or U17211 (N_17211,N_16675,N_16710);
and U17212 (N_17212,N_16985,N_16906);
nand U17213 (N_17213,N_16699,N_16876);
and U17214 (N_17214,N_16705,N_16532);
nand U17215 (N_17215,N_16870,N_16550);
and U17216 (N_17216,N_16740,N_16751);
or U17217 (N_17217,N_16533,N_16847);
nand U17218 (N_17218,N_16994,N_16658);
or U17219 (N_17219,N_16543,N_16968);
or U17220 (N_17220,N_16548,N_16984);
xnor U17221 (N_17221,N_16752,N_16802);
nand U17222 (N_17222,N_16928,N_16770);
and U17223 (N_17223,N_16937,N_16732);
nand U17224 (N_17224,N_16676,N_16584);
and U17225 (N_17225,N_16837,N_16981);
and U17226 (N_17226,N_16738,N_16932);
and U17227 (N_17227,N_16640,N_16663);
nor U17228 (N_17228,N_16809,N_16619);
and U17229 (N_17229,N_16702,N_16961);
and U17230 (N_17230,N_16582,N_16661);
nor U17231 (N_17231,N_16986,N_16912);
or U17232 (N_17232,N_16727,N_16949);
nand U17233 (N_17233,N_16948,N_16952);
nor U17234 (N_17234,N_16801,N_16690);
nor U17235 (N_17235,N_16910,N_16786);
or U17236 (N_17236,N_16841,N_16503);
xnor U17237 (N_17237,N_16557,N_16672);
nand U17238 (N_17238,N_16651,N_16614);
xor U17239 (N_17239,N_16743,N_16660);
nor U17240 (N_17240,N_16739,N_16798);
or U17241 (N_17241,N_16570,N_16908);
xor U17242 (N_17242,N_16758,N_16716);
nand U17243 (N_17243,N_16638,N_16634);
nor U17244 (N_17244,N_16927,N_16991);
and U17245 (N_17245,N_16579,N_16589);
nor U17246 (N_17246,N_16715,N_16872);
and U17247 (N_17247,N_16962,N_16832);
nand U17248 (N_17248,N_16505,N_16776);
or U17249 (N_17249,N_16549,N_16559);
nand U17250 (N_17250,N_16838,N_16561);
or U17251 (N_17251,N_16635,N_16892);
xor U17252 (N_17252,N_16745,N_16686);
or U17253 (N_17253,N_16941,N_16522);
and U17254 (N_17254,N_16845,N_16814);
nor U17255 (N_17255,N_16595,N_16522);
and U17256 (N_17256,N_16791,N_16823);
nor U17257 (N_17257,N_16625,N_16863);
and U17258 (N_17258,N_16989,N_16771);
nand U17259 (N_17259,N_16681,N_16990);
and U17260 (N_17260,N_16870,N_16947);
or U17261 (N_17261,N_16572,N_16768);
xnor U17262 (N_17262,N_16647,N_16539);
nor U17263 (N_17263,N_16535,N_16825);
or U17264 (N_17264,N_16577,N_16579);
nand U17265 (N_17265,N_16872,N_16592);
nand U17266 (N_17266,N_16756,N_16747);
or U17267 (N_17267,N_16911,N_16935);
xnor U17268 (N_17268,N_16869,N_16840);
nand U17269 (N_17269,N_16580,N_16876);
and U17270 (N_17270,N_16857,N_16900);
nand U17271 (N_17271,N_16526,N_16674);
nor U17272 (N_17272,N_16551,N_16750);
nor U17273 (N_17273,N_16747,N_16946);
nor U17274 (N_17274,N_16513,N_16605);
or U17275 (N_17275,N_16696,N_16567);
nor U17276 (N_17276,N_16827,N_16982);
and U17277 (N_17277,N_16745,N_16579);
nor U17278 (N_17278,N_16799,N_16997);
or U17279 (N_17279,N_16971,N_16690);
and U17280 (N_17280,N_16861,N_16852);
and U17281 (N_17281,N_16512,N_16546);
or U17282 (N_17282,N_16745,N_16821);
or U17283 (N_17283,N_16624,N_16948);
xnor U17284 (N_17284,N_16663,N_16578);
or U17285 (N_17285,N_16706,N_16921);
or U17286 (N_17286,N_16914,N_16701);
or U17287 (N_17287,N_16565,N_16776);
nand U17288 (N_17288,N_16610,N_16758);
or U17289 (N_17289,N_16965,N_16968);
or U17290 (N_17290,N_16863,N_16692);
nand U17291 (N_17291,N_16816,N_16525);
xnor U17292 (N_17292,N_16881,N_16608);
nand U17293 (N_17293,N_16654,N_16508);
nand U17294 (N_17294,N_16829,N_16813);
xor U17295 (N_17295,N_16737,N_16508);
xor U17296 (N_17296,N_16563,N_16914);
or U17297 (N_17297,N_16624,N_16865);
and U17298 (N_17298,N_16818,N_16787);
nand U17299 (N_17299,N_16500,N_16608);
nand U17300 (N_17300,N_16699,N_16919);
xor U17301 (N_17301,N_16946,N_16695);
xor U17302 (N_17302,N_16546,N_16717);
and U17303 (N_17303,N_16640,N_16811);
nand U17304 (N_17304,N_16970,N_16876);
or U17305 (N_17305,N_16682,N_16589);
or U17306 (N_17306,N_16879,N_16988);
nor U17307 (N_17307,N_16776,N_16588);
nor U17308 (N_17308,N_16747,N_16581);
and U17309 (N_17309,N_16692,N_16970);
and U17310 (N_17310,N_16777,N_16651);
or U17311 (N_17311,N_16941,N_16895);
and U17312 (N_17312,N_16609,N_16895);
xnor U17313 (N_17313,N_16966,N_16831);
and U17314 (N_17314,N_16999,N_16932);
nor U17315 (N_17315,N_16944,N_16639);
nand U17316 (N_17316,N_16888,N_16560);
or U17317 (N_17317,N_16748,N_16806);
and U17318 (N_17318,N_16556,N_16835);
and U17319 (N_17319,N_16632,N_16910);
and U17320 (N_17320,N_16918,N_16982);
and U17321 (N_17321,N_16617,N_16635);
or U17322 (N_17322,N_16519,N_16781);
xnor U17323 (N_17323,N_16635,N_16518);
nand U17324 (N_17324,N_16896,N_16950);
and U17325 (N_17325,N_16810,N_16872);
nand U17326 (N_17326,N_16679,N_16549);
xnor U17327 (N_17327,N_16772,N_16835);
and U17328 (N_17328,N_16833,N_16835);
and U17329 (N_17329,N_16816,N_16712);
and U17330 (N_17330,N_16672,N_16694);
and U17331 (N_17331,N_16661,N_16620);
nand U17332 (N_17332,N_16594,N_16900);
nand U17333 (N_17333,N_16768,N_16957);
and U17334 (N_17334,N_16717,N_16832);
nand U17335 (N_17335,N_16586,N_16679);
nand U17336 (N_17336,N_16565,N_16623);
or U17337 (N_17337,N_16606,N_16768);
or U17338 (N_17338,N_16562,N_16865);
xnor U17339 (N_17339,N_16952,N_16644);
nor U17340 (N_17340,N_16640,N_16575);
nor U17341 (N_17341,N_16927,N_16683);
nand U17342 (N_17342,N_16509,N_16992);
and U17343 (N_17343,N_16934,N_16916);
nor U17344 (N_17344,N_16787,N_16964);
and U17345 (N_17345,N_16644,N_16823);
nand U17346 (N_17346,N_16981,N_16804);
and U17347 (N_17347,N_16927,N_16854);
or U17348 (N_17348,N_16501,N_16728);
nor U17349 (N_17349,N_16772,N_16716);
and U17350 (N_17350,N_16532,N_16634);
or U17351 (N_17351,N_16606,N_16553);
nand U17352 (N_17352,N_16556,N_16907);
xor U17353 (N_17353,N_16841,N_16980);
and U17354 (N_17354,N_16502,N_16939);
and U17355 (N_17355,N_16634,N_16652);
or U17356 (N_17356,N_16798,N_16758);
xnor U17357 (N_17357,N_16926,N_16934);
nand U17358 (N_17358,N_16507,N_16816);
and U17359 (N_17359,N_16841,N_16989);
xor U17360 (N_17360,N_16656,N_16552);
and U17361 (N_17361,N_16840,N_16717);
and U17362 (N_17362,N_16508,N_16797);
and U17363 (N_17363,N_16612,N_16783);
or U17364 (N_17364,N_16907,N_16708);
or U17365 (N_17365,N_16946,N_16942);
and U17366 (N_17366,N_16554,N_16626);
or U17367 (N_17367,N_16732,N_16725);
xnor U17368 (N_17368,N_16757,N_16700);
or U17369 (N_17369,N_16706,N_16683);
and U17370 (N_17370,N_16563,N_16609);
xor U17371 (N_17371,N_16887,N_16736);
or U17372 (N_17372,N_16813,N_16891);
and U17373 (N_17373,N_16522,N_16986);
nand U17374 (N_17374,N_16885,N_16804);
or U17375 (N_17375,N_16535,N_16989);
and U17376 (N_17376,N_16606,N_16914);
or U17377 (N_17377,N_16550,N_16937);
xnor U17378 (N_17378,N_16933,N_16861);
or U17379 (N_17379,N_16997,N_16870);
or U17380 (N_17380,N_16927,N_16965);
nor U17381 (N_17381,N_16801,N_16703);
nor U17382 (N_17382,N_16805,N_16848);
and U17383 (N_17383,N_16991,N_16742);
nand U17384 (N_17384,N_16558,N_16885);
and U17385 (N_17385,N_16993,N_16506);
xnor U17386 (N_17386,N_16836,N_16891);
or U17387 (N_17387,N_16721,N_16957);
or U17388 (N_17388,N_16930,N_16896);
or U17389 (N_17389,N_16966,N_16986);
and U17390 (N_17390,N_16792,N_16770);
or U17391 (N_17391,N_16801,N_16934);
xor U17392 (N_17392,N_16952,N_16735);
xor U17393 (N_17393,N_16638,N_16566);
nor U17394 (N_17394,N_16759,N_16509);
nor U17395 (N_17395,N_16801,N_16691);
nand U17396 (N_17396,N_16795,N_16911);
and U17397 (N_17397,N_16803,N_16890);
nor U17398 (N_17398,N_16773,N_16764);
and U17399 (N_17399,N_16897,N_16752);
or U17400 (N_17400,N_16648,N_16785);
xnor U17401 (N_17401,N_16789,N_16643);
nor U17402 (N_17402,N_16967,N_16916);
or U17403 (N_17403,N_16979,N_16925);
or U17404 (N_17404,N_16721,N_16731);
xor U17405 (N_17405,N_16867,N_16745);
and U17406 (N_17406,N_16917,N_16609);
or U17407 (N_17407,N_16773,N_16786);
or U17408 (N_17408,N_16868,N_16844);
nor U17409 (N_17409,N_16802,N_16933);
nand U17410 (N_17410,N_16733,N_16948);
nand U17411 (N_17411,N_16870,N_16513);
or U17412 (N_17412,N_16657,N_16786);
nor U17413 (N_17413,N_16745,N_16839);
nor U17414 (N_17414,N_16604,N_16774);
nand U17415 (N_17415,N_16549,N_16665);
xor U17416 (N_17416,N_16855,N_16839);
nor U17417 (N_17417,N_16525,N_16636);
nand U17418 (N_17418,N_16641,N_16782);
or U17419 (N_17419,N_16957,N_16997);
nand U17420 (N_17420,N_16769,N_16599);
or U17421 (N_17421,N_16546,N_16610);
and U17422 (N_17422,N_16760,N_16699);
nor U17423 (N_17423,N_16799,N_16621);
and U17424 (N_17424,N_16856,N_16586);
nor U17425 (N_17425,N_16841,N_16888);
or U17426 (N_17426,N_16783,N_16965);
xnor U17427 (N_17427,N_16833,N_16885);
nand U17428 (N_17428,N_16669,N_16764);
xnor U17429 (N_17429,N_16506,N_16677);
nand U17430 (N_17430,N_16769,N_16578);
xnor U17431 (N_17431,N_16652,N_16518);
or U17432 (N_17432,N_16577,N_16691);
and U17433 (N_17433,N_16669,N_16633);
and U17434 (N_17434,N_16674,N_16918);
nor U17435 (N_17435,N_16709,N_16773);
and U17436 (N_17436,N_16639,N_16679);
nand U17437 (N_17437,N_16596,N_16749);
xor U17438 (N_17438,N_16931,N_16508);
xnor U17439 (N_17439,N_16829,N_16857);
nor U17440 (N_17440,N_16586,N_16935);
nand U17441 (N_17441,N_16871,N_16609);
nand U17442 (N_17442,N_16542,N_16576);
or U17443 (N_17443,N_16563,N_16778);
xor U17444 (N_17444,N_16867,N_16632);
or U17445 (N_17445,N_16629,N_16798);
or U17446 (N_17446,N_16859,N_16519);
nor U17447 (N_17447,N_16601,N_16688);
or U17448 (N_17448,N_16531,N_16652);
nand U17449 (N_17449,N_16808,N_16509);
and U17450 (N_17450,N_16968,N_16746);
xnor U17451 (N_17451,N_16869,N_16873);
and U17452 (N_17452,N_16976,N_16690);
nor U17453 (N_17453,N_16976,N_16823);
or U17454 (N_17454,N_16752,N_16631);
nand U17455 (N_17455,N_16931,N_16884);
nor U17456 (N_17456,N_16910,N_16538);
or U17457 (N_17457,N_16812,N_16710);
or U17458 (N_17458,N_16714,N_16995);
nor U17459 (N_17459,N_16926,N_16683);
xnor U17460 (N_17460,N_16929,N_16507);
nor U17461 (N_17461,N_16734,N_16659);
nand U17462 (N_17462,N_16789,N_16747);
and U17463 (N_17463,N_16742,N_16854);
or U17464 (N_17464,N_16775,N_16625);
nand U17465 (N_17465,N_16579,N_16961);
and U17466 (N_17466,N_16916,N_16631);
nand U17467 (N_17467,N_16888,N_16991);
nand U17468 (N_17468,N_16834,N_16742);
or U17469 (N_17469,N_16969,N_16652);
nand U17470 (N_17470,N_16854,N_16678);
or U17471 (N_17471,N_16785,N_16894);
or U17472 (N_17472,N_16989,N_16987);
and U17473 (N_17473,N_16709,N_16558);
nor U17474 (N_17474,N_16731,N_16651);
xor U17475 (N_17475,N_16639,N_16732);
nand U17476 (N_17476,N_16916,N_16973);
xor U17477 (N_17477,N_16980,N_16546);
nand U17478 (N_17478,N_16868,N_16526);
or U17479 (N_17479,N_16605,N_16868);
xnor U17480 (N_17480,N_16810,N_16850);
nand U17481 (N_17481,N_16847,N_16620);
or U17482 (N_17482,N_16766,N_16574);
xor U17483 (N_17483,N_16810,N_16885);
and U17484 (N_17484,N_16776,N_16701);
nor U17485 (N_17485,N_16871,N_16798);
and U17486 (N_17486,N_16915,N_16804);
nand U17487 (N_17487,N_16668,N_16715);
nand U17488 (N_17488,N_16603,N_16948);
nand U17489 (N_17489,N_16665,N_16769);
xor U17490 (N_17490,N_16537,N_16550);
nand U17491 (N_17491,N_16860,N_16761);
nor U17492 (N_17492,N_16748,N_16877);
nor U17493 (N_17493,N_16588,N_16662);
or U17494 (N_17494,N_16782,N_16996);
nand U17495 (N_17495,N_16919,N_16705);
and U17496 (N_17496,N_16571,N_16893);
or U17497 (N_17497,N_16841,N_16730);
or U17498 (N_17498,N_16812,N_16790);
nand U17499 (N_17499,N_16674,N_16855);
or U17500 (N_17500,N_17274,N_17100);
or U17501 (N_17501,N_17073,N_17030);
and U17502 (N_17502,N_17383,N_17219);
xnor U17503 (N_17503,N_17349,N_17482);
xnor U17504 (N_17504,N_17236,N_17089);
and U17505 (N_17505,N_17156,N_17101);
xnor U17506 (N_17506,N_17483,N_17427);
nand U17507 (N_17507,N_17471,N_17259);
or U17508 (N_17508,N_17064,N_17114);
nor U17509 (N_17509,N_17110,N_17258);
and U17510 (N_17510,N_17282,N_17496);
and U17511 (N_17511,N_17240,N_17308);
nand U17512 (N_17512,N_17499,N_17480);
nand U17513 (N_17513,N_17466,N_17304);
xor U17514 (N_17514,N_17205,N_17302);
nand U17515 (N_17515,N_17194,N_17199);
or U17516 (N_17516,N_17084,N_17394);
and U17517 (N_17517,N_17347,N_17370);
and U17518 (N_17518,N_17005,N_17348);
xnor U17519 (N_17519,N_17458,N_17147);
nand U17520 (N_17520,N_17315,N_17485);
or U17521 (N_17521,N_17031,N_17405);
xnor U17522 (N_17522,N_17452,N_17432);
xnor U17523 (N_17523,N_17209,N_17299);
or U17524 (N_17524,N_17008,N_17185);
and U17525 (N_17525,N_17234,N_17392);
nand U17526 (N_17526,N_17036,N_17342);
and U17527 (N_17527,N_17306,N_17275);
nor U17528 (N_17528,N_17099,N_17389);
and U17529 (N_17529,N_17495,N_17492);
nand U17530 (N_17530,N_17182,N_17243);
or U17531 (N_17531,N_17415,N_17417);
or U17532 (N_17532,N_17378,N_17037);
nor U17533 (N_17533,N_17293,N_17113);
nor U17534 (N_17534,N_17312,N_17157);
nor U17535 (N_17535,N_17134,N_17352);
nor U17536 (N_17536,N_17333,N_17374);
xor U17537 (N_17537,N_17484,N_17358);
nand U17538 (N_17538,N_17404,N_17455);
and U17539 (N_17539,N_17400,N_17192);
and U17540 (N_17540,N_17323,N_17246);
xnor U17541 (N_17541,N_17053,N_17191);
xor U17542 (N_17542,N_17138,N_17310);
xor U17543 (N_17543,N_17414,N_17411);
xor U17544 (N_17544,N_17057,N_17011);
nand U17545 (N_17545,N_17367,N_17369);
nand U17546 (N_17546,N_17339,N_17060);
xnor U17547 (N_17547,N_17211,N_17033);
nor U17548 (N_17548,N_17317,N_17289);
nor U17549 (N_17549,N_17026,N_17094);
nor U17550 (N_17550,N_17437,N_17221);
xnor U17551 (N_17551,N_17150,N_17050);
and U17552 (N_17552,N_17255,N_17195);
xnor U17553 (N_17553,N_17272,N_17158);
and U17554 (N_17554,N_17001,N_17264);
nor U17555 (N_17555,N_17167,N_17168);
or U17556 (N_17556,N_17468,N_17295);
nand U17557 (N_17557,N_17314,N_17444);
nor U17558 (N_17558,N_17297,N_17334);
nor U17559 (N_17559,N_17397,N_17111);
nor U17560 (N_17560,N_17474,N_17149);
nor U17561 (N_17561,N_17395,N_17430);
xnor U17562 (N_17562,N_17388,N_17385);
and U17563 (N_17563,N_17039,N_17386);
xnor U17564 (N_17564,N_17305,N_17004);
nor U17565 (N_17565,N_17269,N_17017);
or U17566 (N_17566,N_17467,N_17301);
nor U17567 (N_17567,N_17038,N_17248);
nand U17568 (N_17568,N_17140,N_17164);
xor U17569 (N_17569,N_17375,N_17095);
or U17570 (N_17570,N_17316,N_17445);
nand U17571 (N_17571,N_17131,N_17279);
nor U17572 (N_17572,N_17242,N_17262);
nor U17573 (N_17573,N_17051,N_17252);
or U17574 (N_17574,N_17090,N_17022);
or U17575 (N_17575,N_17398,N_17442);
nor U17576 (N_17576,N_17227,N_17337);
xnor U17577 (N_17577,N_17244,N_17451);
nand U17578 (N_17578,N_17491,N_17062);
xnor U17579 (N_17579,N_17103,N_17307);
nor U17580 (N_17580,N_17351,N_17019);
nor U17581 (N_17581,N_17379,N_17124);
xor U17582 (N_17582,N_17329,N_17224);
and U17583 (N_17583,N_17215,N_17396);
nand U17584 (N_17584,N_17024,N_17043);
and U17585 (N_17585,N_17159,N_17436);
and U17586 (N_17586,N_17145,N_17146);
nand U17587 (N_17587,N_17280,N_17237);
and U17588 (N_17588,N_17254,N_17230);
xor U17589 (N_17589,N_17179,N_17406);
xor U17590 (N_17590,N_17488,N_17420);
nand U17591 (N_17591,N_17371,N_17076);
or U17592 (N_17592,N_17440,N_17122);
xnor U17593 (N_17593,N_17197,N_17129);
xnor U17594 (N_17594,N_17216,N_17335);
and U17595 (N_17595,N_17384,N_17341);
nand U17596 (N_17596,N_17006,N_17196);
nand U17597 (N_17597,N_17018,N_17402);
and U17598 (N_17598,N_17476,N_17273);
nor U17599 (N_17599,N_17020,N_17190);
xnor U17600 (N_17600,N_17261,N_17487);
or U17601 (N_17601,N_17325,N_17490);
nor U17602 (N_17602,N_17169,N_17127);
or U17603 (N_17603,N_17231,N_17340);
and U17604 (N_17604,N_17220,N_17447);
nor U17605 (N_17605,N_17413,N_17013);
xnor U17606 (N_17606,N_17377,N_17330);
xnor U17607 (N_17607,N_17429,N_17373);
or U17608 (N_17608,N_17034,N_17331);
and U17609 (N_17609,N_17067,N_17403);
nor U17610 (N_17610,N_17443,N_17338);
nand U17611 (N_17611,N_17498,N_17065);
nor U17612 (N_17612,N_17015,N_17213);
nand U17613 (N_17613,N_17345,N_17118);
nand U17614 (N_17614,N_17016,N_17357);
nor U17615 (N_17615,N_17207,N_17281);
nor U17616 (N_17616,N_17108,N_17470);
xnor U17617 (N_17617,N_17233,N_17407);
xor U17618 (N_17618,N_17446,N_17290);
xnor U17619 (N_17619,N_17346,N_17174);
or U17620 (N_17620,N_17217,N_17071);
and U17621 (N_17621,N_17418,N_17105);
nand U17622 (N_17622,N_17098,N_17046);
and U17623 (N_17623,N_17126,N_17355);
nor U17624 (N_17624,N_17165,N_17226);
xnor U17625 (N_17625,N_17133,N_17336);
nor U17626 (N_17626,N_17303,N_17266);
nand U17627 (N_17627,N_17080,N_17286);
xnor U17628 (N_17628,N_17287,N_17000);
or U17629 (N_17629,N_17296,N_17072);
and U17630 (N_17630,N_17202,N_17225);
or U17631 (N_17631,N_17184,N_17428);
and U17632 (N_17632,N_17453,N_17441);
nor U17633 (N_17633,N_17271,N_17125);
nand U17634 (N_17634,N_17069,N_17093);
nor U17635 (N_17635,N_17381,N_17390);
xor U17636 (N_17636,N_17241,N_17088);
nor U17637 (N_17637,N_17267,N_17180);
nand U17638 (N_17638,N_17327,N_17232);
or U17639 (N_17639,N_17494,N_17223);
xnor U17640 (N_17640,N_17035,N_17063);
nor U17641 (N_17641,N_17462,N_17078);
or U17642 (N_17642,N_17218,N_17040);
nor U17643 (N_17643,N_17363,N_17387);
nand U17644 (N_17644,N_17083,N_17068);
nand U17645 (N_17645,N_17059,N_17077);
or U17646 (N_17646,N_17278,N_17300);
and U17647 (N_17647,N_17200,N_17176);
and U17648 (N_17648,N_17343,N_17141);
xor U17649 (N_17649,N_17364,N_17356);
nor U17650 (N_17650,N_17438,N_17028);
nor U17651 (N_17651,N_17171,N_17204);
and U17652 (N_17652,N_17136,N_17132);
xnor U17653 (N_17653,N_17142,N_17206);
nor U17654 (N_17654,N_17092,N_17464);
xor U17655 (N_17655,N_17419,N_17066);
nand U17656 (N_17656,N_17313,N_17048);
nor U17657 (N_17657,N_17439,N_17450);
or U17658 (N_17658,N_17409,N_17479);
xor U17659 (N_17659,N_17320,N_17493);
nand U17660 (N_17660,N_17049,N_17014);
nor U17661 (N_17661,N_17044,N_17459);
nand U17662 (N_17662,N_17096,N_17189);
xor U17663 (N_17663,N_17311,N_17294);
nor U17664 (N_17664,N_17298,N_17250);
or U17665 (N_17665,N_17023,N_17270);
and U17666 (N_17666,N_17319,N_17449);
and U17667 (N_17667,N_17128,N_17010);
xor U17668 (N_17668,N_17143,N_17139);
and U17669 (N_17669,N_17042,N_17332);
and U17670 (N_17670,N_17309,N_17082);
or U17671 (N_17671,N_17257,N_17475);
or U17672 (N_17672,N_17123,N_17291);
and U17673 (N_17673,N_17201,N_17235);
or U17674 (N_17674,N_17362,N_17193);
and U17675 (N_17675,N_17009,N_17360);
nand U17676 (N_17676,N_17086,N_17324);
and U17677 (N_17677,N_17353,N_17391);
and U17678 (N_17678,N_17457,N_17328);
xnor U17679 (N_17679,N_17135,N_17172);
and U17680 (N_17680,N_17003,N_17203);
nor U17681 (N_17681,N_17107,N_17055);
nor U17682 (N_17682,N_17032,N_17175);
nor U17683 (N_17683,N_17116,N_17115);
and U17684 (N_17684,N_17228,N_17151);
xor U17685 (N_17685,N_17460,N_17277);
nor U17686 (N_17686,N_17399,N_17166);
xnor U17687 (N_17687,N_17421,N_17401);
xor U17688 (N_17688,N_17104,N_17393);
nor U17689 (N_17689,N_17412,N_17117);
xor U17690 (N_17690,N_17148,N_17170);
nand U17691 (N_17691,N_17497,N_17045);
nand U17692 (N_17692,N_17276,N_17292);
nor U17693 (N_17693,N_17408,N_17431);
xnor U17694 (N_17694,N_17247,N_17489);
nor U17695 (N_17695,N_17075,N_17473);
nor U17696 (N_17696,N_17283,N_17463);
or U17697 (N_17697,N_17119,N_17188);
or U17698 (N_17698,N_17326,N_17144);
nand U17699 (N_17699,N_17288,N_17154);
xnor U17700 (N_17700,N_17178,N_17183);
or U17701 (N_17701,N_17198,N_17249);
and U17702 (N_17702,N_17162,N_17376);
and U17703 (N_17703,N_17021,N_17187);
nor U17704 (N_17704,N_17285,N_17321);
or U17705 (N_17705,N_17054,N_17186);
and U17706 (N_17706,N_17469,N_17041);
xnor U17707 (N_17707,N_17268,N_17425);
nor U17708 (N_17708,N_17210,N_17130);
or U17709 (N_17709,N_17424,N_17365);
and U17710 (N_17710,N_17012,N_17079);
nor U17711 (N_17711,N_17465,N_17251);
xnor U17712 (N_17712,N_17007,N_17097);
nor U17713 (N_17713,N_17222,N_17354);
nand U17714 (N_17714,N_17047,N_17173);
nor U17715 (N_17715,N_17461,N_17106);
or U17716 (N_17716,N_17410,N_17229);
and U17717 (N_17717,N_17260,N_17163);
xnor U17718 (N_17718,N_17366,N_17155);
nand U17719 (N_17719,N_17161,N_17433);
nor U17720 (N_17720,N_17120,N_17208);
or U17721 (N_17721,N_17085,N_17029);
nand U17722 (N_17722,N_17284,N_17102);
nor U17723 (N_17723,N_17472,N_17074);
nand U17724 (N_17724,N_17027,N_17058);
nand U17725 (N_17725,N_17214,N_17344);
nor U17726 (N_17726,N_17212,N_17056);
nor U17727 (N_17727,N_17477,N_17121);
and U17728 (N_17728,N_17025,N_17256);
xnor U17729 (N_17729,N_17153,N_17322);
or U17730 (N_17730,N_17109,N_17160);
nand U17731 (N_17731,N_17112,N_17434);
nand U17732 (N_17732,N_17239,N_17238);
or U17733 (N_17733,N_17181,N_17423);
and U17734 (N_17734,N_17478,N_17081);
and U17735 (N_17735,N_17091,N_17361);
or U17736 (N_17736,N_17435,N_17137);
nand U17737 (N_17737,N_17061,N_17382);
or U17738 (N_17738,N_17318,N_17486);
or U17739 (N_17739,N_17245,N_17372);
and U17740 (N_17740,N_17177,N_17263);
xor U17741 (N_17741,N_17253,N_17448);
nor U17742 (N_17742,N_17052,N_17454);
nor U17743 (N_17743,N_17380,N_17368);
nand U17744 (N_17744,N_17456,N_17426);
or U17745 (N_17745,N_17002,N_17265);
and U17746 (N_17746,N_17481,N_17087);
and U17747 (N_17747,N_17359,N_17070);
and U17748 (N_17748,N_17416,N_17350);
or U17749 (N_17749,N_17152,N_17422);
and U17750 (N_17750,N_17333,N_17168);
or U17751 (N_17751,N_17426,N_17246);
or U17752 (N_17752,N_17232,N_17177);
xor U17753 (N_17753,N_17494,N_17475);
nor U17754 (N_17754,N_17301,N_17314);
and U17755 (N_17755,N_17065,N_17336);
or U17756 (N_17756,N_17185,N_17159);
nor U17757 (N_17757,N_17391,N_17040);
and U17758 (N_17758,N_17451,N_17113);
nand U17759 (N_17759,N_17013,N_17359);
or U17760 (N_17760,N_17123,N_17116);
and U17761 (N_17761,N_17225,N_17319);
and U17762 (N_17762,N_17388,N_17374);
or U17763 (N_17763,N_17180,N_17288);
nor U17764 (N_17764,N_17151,N_17395);
or U17765 (N_17765,N_17481,N_17340);
and U17766 (N_17766,N_17248,N_17275);
nor U17767 (N_17767,N_17404,N_17060);
xnor U17768 (N_17768,N_17403,N_17460);
xor U17769 (N_17769,N_17451,N_17389);
and U17770 (N_17770,N_17059,N_17016);
and U17771 (N_17771,N_17339,N_17407);
and U17772 (N_17772,N_17495,N_17242);
or U17773 (N_17773,N_17014,N_17342);
nor U17774 (N_17774,N_17334,N_17451);
nand U17775 (N_17775,N_17371,N_17259);
nand U17776 (N_17776,N_17167,N_17161);
nand U17777 (N_17777,N_17037,N_17316);
nand U17778 (N_17778,N_17399,N_17104);
or U17779 (N_17779,N_17052,N_17183);
nand U17780 (N_17780,N_17483,N_17266);
nor U17781 (N_17781,N_17082,N_17316);
nand U17782 (N_17782,N_17140,N_17206);
nor U17783 (N_17783,N_17369,N_17395);
nand U17784 (N_17784,N_17118,N_17420);
xnor U17785 (N_17785,N_17322,N_17394);
and U17786 (N_17786,N_17253,N_17405);
nand U17787 (N_17787,N_17093,N_17167);
and U17788 (N_17788,N_17497,N_17241);
nand U17789 (N_17789,N_17470,N_17415);
nand U17790 (N_17790,N_17192,N_17061);
nor U17791 (N_17791,N_17051,N_17467);
and U17792 (N_17792,N_17499,N_17016);
nor U17793 (N_17793,N_17062,N_17239);
nand U17794 (N_17794,N_17341,N_17162);
nor U17795 (N_17795,N_17208,N_17306);
and U17796 (N_17796,N_17280,N_17188);
nand U17797 (N_17797,N_17382,N_17227);
and U17798 (N_17798,N_17358,N_17209);
xnor U17799 (N_17799,N_17196,N_17154);
nand U17800 (N_17800,N_17325,N_17170);
nor U17801 (N_17801,N_17107,N_17074);
nor U17802 (N_17802,N_17367,N_17058);
and U17803 (N_17803,N_17420,N_17194);
nor U17804 (N_17804,N_17062,N_17237);
nand U17805 (N_17805,N_17397,N_17317);
nor U17806 (N_17806,N_17342,N_17331);
xor U17807 (N_17807,N_17330,N_17151);
nor U17808 (N_17808,N_17091,N_17407);
nand U17809 (N_17809,N_17079,N_17250);
xor U17810 (N_17810,N_17108,N_17076);
nand U17811 (N_17811,N_17200,N_17179);
or U17812 (N_17812,N_17199,N_17461);
and U17813 (N_17813,N_17443,N_17367);
nor U17814 (N_17814,N_17094,N_17086);
nor U17815 (N_17815,N_17297,N_17317);
and U17816 (N_17816,N_17110,N_17352);
and U17817 (N_17817,N_17414,N_17211);
and U17818 (N_17818,N_17489,N_17352);
and U17819 (N_17819,N_17015,N_17283);
and U17820 (N_17820,N_17000,N_17338);
nand U17821 (N_17821,N_17159,N_17081);
nor U17822 (N_17822,N_17042,N_17209);
and U17823 (N_17823,N_17199,N_17270);
nand U17824 (N_17824,N_17073,N_17399);
and U17825 (N_17825,N_17427,N_17322);
nand U17826 (N_17826,N_17301,N_17127);
and U17827 (N_17827,N_17103,N_17135);
nand U17828 (N_17828,N_17309,N_17172);
nor U17829 (N_17829,N_17373,N_17207);
nor U17830 (N_17830,N_17447,N_17415);
nor U17831 (N_17831,N_17367,N_17272);
and U17832 (N_17832,N_17410,N_17443);
and U17833 (N_17833,N_17213,N_17247);
or U17834 (N_17834,N_17205,N_17125);
nand U17835 (N_17835,N_17147,N_17472);
and U17836 (N_17836,N_17341,N_17440);
nor U17837 (N_17837,N_17193,N_17408);
nand U17838 (N_17838,N_17319,N_17185);
nand U17839 (N_17839,N_17084,N_17317);
nand U17840 (N_17840,N_17229,N_17227);
and U17841 (N_17841,N_17129,N_17315);
nand U17842 (N_17842,N_17190,N_17024);
nand U17843 (N_17843,N_17145,N_17454);
and U17844 (N_17844,N_17035,N_17485);
nor U17845 (N_17845,N_17350,N_17292);
or U17846 (N_17846,N_17473,N_17497);
nand U17847 (N_17847,N_17447,N_17423);
and U17848 (N_17848,N_17359,N_17043);
or U17849 (N_17849,N_17048,N_17126);
xnor U17850 (N_17850,N_17227,N_17143);
xnor U17851 (N_17851,N_17138,N_17249);
and U17852 (N_17852,N_17264,N_17357);
and U17853 (N_17853,N_17272,N_17330);
and U17854 (N_17854,N_17461,N_17163);
xor U17855 (N_17855,N_17271,N_17052);
xnor U17856 (N_17856,N_17496,N_17034);
or U17857 (N_17857,N_17361,N_17450);
and U17858 (N_17858,N_17019,N_17355);
nor U17859 (N_17859,N_17137,N_17465);
or U17860 (N_17860,N_17272,N_17104);
nand U17861 (N_17861,N_17364,N_17417);
nand U17862 (N_17862,N_17184,N_17072);
and U17863 (N_17863,N_17199,N_17471);
nor U17864 (N_17864,N_17225,N_17390);
or U17865 (N_17865,N_17156,N_17131);
xnor U17866 (N_17866,N_17115,N_17282);
and U17867 (N_17867,N_17182,N_17462);
nor U17868 (N_17868,N_17022,N_17406);
xor U17869 (N_17869,N_17336,N_17050);
xor U17870 (N_17870,N_17432,N_17226);
xnor U17871 (N_17871,N_17054,N_17319);
nand U17872 (N_17872,N_17269,N_17313);
nor U17873 (N_17873,N_17499,N_17229);
xnor U17874 (N_17874,N_17211,N_17278);
nor U17875 (N_17875,N_17024,N_17069);
nor U17876 (N_17876,N_17148,N_17449);
or U17877 (N_17877,N_17156,N_17053);
xor U17878 (N_17878,N_17041,N_17208);
nor U17879 (N_17879,N_17186,N_17166);
xnor U17880 (N_17880,N_17234,N_17412);
xor U17881 (N_17881,N_17039,N_17123);
xor U17882 (N_17882,N_17019,N_17451);
nand U17883 (N_17883,N_17202,N_17004);
or U17884 (N_17884,N_17193,N_17309);
and U17885 (N_17885,N_17077,N_17326);
or U17886 (N_17886,N_17369,N_17261);
nand U17887 (N_17887,N_17441,N_17131);
nand U17888 (N_17888,N_17190,N_17228);
xor U17889 (N_17889,N_17389,N_17453);
or U17890 (N_17890,N_17388,N_17204);
nand U17891 (N_17891,N_17125,N_17046);
or U17892 (N_17892,N_17140,N_17443);
nor U17893 (N_17893,N_17453,N_17334);
nor U17894 (N_17894,N_17164,N_17326);
or U17895 (N_17895,N_17322,N_17132);
and U17896 (N_17896,N_17193,N_17425);
nand U17897 (N_17897,N_17179,N_17237);
nor U17898 (N_17898,N_17354,N_17177);
xnor U17899 (N_17899,N_17306,N_17205);
nor U17900 (N_17900,N_17014,N_17040);
or U17901 (N_17901,N_17355,N_17002);
and U17902 (N_17902,N_17217,N_17307);
and U17903 (N_17903,N_17456,N_17195);
nand U17904 (N_17904,N_17253,N_17438);
or U17905 (N_17905,N_17375,N_17118);
nor U17906 (N_17906,N_17029,N_17394);
nor U17907 (N_17907,N_17365,N_17348);
xnor U17908 (N_17908,N_17000,N_17434);
or U17909 (N_17909,N_17206,N_17340);
nor U17910 (N_17910,N_17311,N_17247);
and U17911 (N_17911,N_17010,N_17267);
or U17912 (N_17912,N_17021,N_17074);
or U17913 (N_17913,N_17495,N_17228);
and U17914 (N_17914,N_17008,N_17472);
nand U17915 (N_17915,N_17400,N_17169);
nand U17916 (N_17916,N_17137,N_17281);
or U17917 (N_17917,N_17481,N_17473);
or U17918 (N_17918,N_17218,N_17206);
and U17919 (N_17919,N_17216,N_17376);
or U17920 (N_17920,N_17475,N_17272);
and U17921 (N_17921,N_17119,N_17163);
and U17922 (N_17922,N_17303,N_17371);
nor U17923 (N_17923,N_17421,N_17309);
xnor U17924 (N_17924,N_17142,N_17052);
xor U17925 (N_17925,N_17399,N_17007);
nand U17926 (N_17926,N_17174,N_17232);
nor U17927 (N_17927,N_17427,N_17484);
or U17928 (N_17928,N_17387,N_17371);
or U17929 (N_17929,N_17193,N_17465);
and U17930 (N_17930,N_17124,N_17170);
nor U17931 (N_17931,N_17400,N_17227);
nor U17932 (N_17932,N_17096,N_17085);
xnor U17933 (N_17933,N_17282,N_17136);
xor U17934 (N_17934,N_17308,N_17338);
nor U17935 (N_17935,N_17331,N_17114);
or U17936 (N_17936,N_17167,N_17213);
or U17937 (N_17937,N_17042,N_17254);
xnor U17938 (N_17938,N_17181,N_17482);
and U17939 (N_17939,N_17200,N_17390);
xnor U17940 (N_17940,N_17280,N_17303);
xnor U17941 (N_17941,N_17283,N_17003);
and U17942 (N_17942,N_17212,N_17174);
and U17943 (N_17943,N_17191,N_17228);
nand U17944 (N_17944,N_17483,N_17019);
or U17945 (N_17945,N_17479,N_17403);
xor U17946 (N_17946,N_17147,N_17112);
nand U17947 (N_17947,N_17317,N_17241);
or U17948 (N_17948,N_17100,N_17178);
xnor U17949 (N_17949,N_17297,N_17281);
xor U17950 (N_17950,N_17377,N_17439);
xnor U17951 (N_17951,N_17435,N_17145);
xor U17952 (N_17952,N_17016,N_17102);
and U17953 (N_17953,N_17475,N_17121);
and U17954 (N_17954,N_17101,N_17286);
nor U17955 (N_17955,N_17488,N_17214);
and U17956 (N_17956,N_17370,N_17344);
xnor U17957 (N_17957,N_17186,N_17396);
nand U17958 (N_17958,N_17347,N_17480);
nand U17959 (N_17959,N_17307,N_17080);
and U17960 (N_17960,N_17219,N_17000);
nand U17961 (N_17961,N_17088,N_17286);
xor U17962 (N_17962,N_17111,N_17494);
xor U17963 (N_17963,N_17157,N_17199);
nor U17964 (N_17964,N_17009,N_17316);
nor U17965 (N_17965,N_17437,N_17030);
or U17966 (N_17966,N_17085,N_17116);
nand U17967 (N_17967,N_17098,N_17217);
and U17968 (N_17968,N_17090,N_17357);
nand U17969 (N_17969,N_17040,N_17315);
nand U17970 (N_17970,N_17400,N_17263);
or U17971 (N_17971,N_17397,N_17282);
and U17972 (N_17972,N_17108,N_17015);
nand U17973 (N_17973,N_17304,N_17039);
nand U17974 (N_17974,N_17276,N_17193);
and U17975 (N_17975,N_17466,N_17385);
nor U17976 (N_17976,N_17450,N_17043);
nor U17977 (N_17977,N_17471,N_17131);
nor U17978 (N_17978,N_17482,N_17085);
and U17979 (N_17979,N_17124,N_17105);
and U17980 (N_17980,N_17020,N_17277);
or U17981 (N_17981,N_17429,N_17273);
nor U17982 (N_17982,N_17354,N_17303);
or U17983 (N_17983,N_17187,N_17053);
or U17984 (N_17984,N_17452,N_17381);
and U17985 (N_17985,N_17348,N_17220);
nor U17986 (N_17986,N_17076,N_17272);
or U17987 (N_17987,N_17145,N_17054);
xor U17988 (N_17988,N_17021,N_17042);
nor U17989 (N_17989,N_17147,N_17379);
xnor U17990 (N_17990,N_17364,N_17039);
nand U17991 (N_17991,N_17126,N_17293);
nand U17992 (N_17992,N_17416,N_17433);
nor U17993 (N_17993,N_17175,N_17445);
xnor U17994 (N_17994,N_17222,N_17015);
or U17995 (N_17995,N_17081,N_17379);
nand U17996 (N_17996,N_17229,N_17153);
nand U17997 (N_17997,N_17169,N_17107);
and U17998 (N_17998,N_17054,N_17291);
and U17999 (N_17999,N_17170,N_17491);
and U18000 (N_18000,N_17693,N_17540);
nor U18001 (N_18001,N_17611,N_17690);
and U18002 (N_18002,N_17989,N_17701);
xor U18003 (N_18003,N_17729,N_17551);
or U18004 (N_18004,N_17728,N_17986);
or U18005 (N_18005,N_17633,N_17565);
nor U18006 (N_18006,N_17666,N_17716);
or U18007 (N_18007,N_17832,N_17634);
and U18008 (N_18008,N_17584,N_17527);
or U18009 (N_18009,N_17742,N_17833);
nor U18010 (N_18010,N_17929,N_17831);
and U18011 (N_18011,N_17965,N_17974);
nand U18012 (N_18012,N_17844,N_17776);
nor U18013 (N_18013,N_17758,N_17569);
nor U18014 (N_18014,N_17753,N_17582);
or U18015 (N_18015,N_17624,N_17916);
or U18016 (N_18016,N_17625,N_17530);
nor U18017 (N_18017,N_17902,N_17712);
and U18018 (N_18018,N_17980,N_17620);
or U18019 (N_18019,N_17834,N_17721);
and U18020 (N_18020,N_17500,N_17797);
and U18021 (N_18021,N_17763,N_17713);
and U18022 (N_18022,N_17732,N_17523);
xnor U18023 (N_18023,N_17631,N_17670);
xnor U18024 (N_18024,N_17843,N_17847);
nor U18025 (N_18025,N_17755,N_17684);
nor U18026 (N_18026,N_17999,N_17588);
and U18027 (N_18027,N_17830,N_17969);
or U18028 (N_18028,N_17703,N_17691);
nand U18029 (N_18029,N_17917,N_17737);
or U18030 (N_18030,N_17570,N_17676);
or U18031 (N_18031,N_17510,N_17984);
nor U18032 (N_18032,N_17738,N_17803);
xnor U18033 (N_18033,N_17692,N_17892);
and U18034 (N_18034,N_17535,N_17780);
nand U18035 (N_18035,N_17702,N_17931);
nor U18036 (N_18036,N_17815,N_17910);
nand U18037 (N_18037,N_17529,N_17585);
or U18038 (N_18038,N_17784,N_17814);
or U18039 (N_18039,N_17654,N_17842);
and U18040 (N_18040,N_17578,N_17733);
nor U18041 (N_18041,N_17883,N_17592);
or U18042 (N_18042,N_17757,N_17526);
xor U18043 (N_18043,N_17946,N_17586);
and U18044 (N_18044,N_17767,N_17560);
nand U18045 (N_18045,N_17508,N_17710);
nor U18046 (N_18046,N_17860,N_17517);
or U18047 (N_18047,N_17635,N_17935);
nand U18048 (N_18048,N_17900,N_17513);
or U18049 (N_18049,N_17849,N_17550);
xor U18050 (N_18050,N_17562,N_17765);
xor U18051 (N_18051,N_17736,N_17559);
or U18052 (N_18052,N_17720,N_17689);
and U18053 (N_18053,N_17786,N_17822);
or U18054 (N_18054,N_17995,N_17563);
and U18055 (N_18055,N_17516,N_17875);
nand U18056 (N_18056,N_17514,N_17991);
nor U18057 (N_18057,N_17561,N_17846);
or U18058 (N_18058,N_17744,N_17992);
or U18059 (N_18059,N_17939,N_17660);
or U18060 (N_18060,N_17557,N_17795);
nand U18061 (N_18061,N_17821,N_17714);
and U18062 (N_18062,N_17813,N_17667);
xnor U18063 (N_18063,N_17951,N_17606);
and U18064 (N_18064,N_17545,N_17699);
and U18065 (N_18065,N_17623,N_17656);
nand U18066 (N_18066,N_17683,N_17783);
nand U18067 (N_18067,N_17638,N_17807);
nor U18068 (N_18068,N_17956,N_17657);
and U18069 (N_18069,N_17750,N_17519);
xnor U18070 (N_18070,N_17687,N_17533);
nor U18071 (N_18071,N_17663,N_17773);
nand U18072 (N_18072,N_17976,N_17590);
nor U18073 (N_18073,N_17711,N_17829);
nor U18074 (N_18074,N_17983,N_17648);
nand U18075 (N_18075,N_17981,N_17665);
and U18076 (N_18076,N_17962,N_17659);
and U18077 (N_18077,N_17552,N_17791);
and U18078 (N_18078,N_17511,N_17779);
nor U18079 (N_18079,N_17885,N_17839);
nor U18080 (N_18080,N_17521,N_17769);
nand U18081 (N_18081,N_17662,N_17927);
nor U18082 (N_18082,N_17622,N_17646);
or U18083 (N_18083,N_17998,N_17942);
and U18084 (N_18084,N_17644,N_17809);
and U18085 (N_18085,N_17777,N_17906);
xor U18086 (N_18086,N_17715,N_17694);
and U18087 (N_18087,N_17655,N_17887);
nand U18088 (N_18088,N_17610,N_17515);
xor U18089 (N_18089,N_17564,N_17587);
xor U18090 (N_18090,N_17940,N_17837);
or U18091 (N_18091,N_17966,N_17840);
xor U18092 (N_18092,N_17651,N_17913);
nor U18093 (N_18093,N_17688,N_17524);
xor U18094 (N_18094,N_17658,N_17864);
or U18095 (N_18095,N_17947,N_17909);
or U18096 (N_18096,N_17677,N_17889);
nand U18097 (N_18097,N_17575,N_17705);
nor U18098 (N_18098,N_17760,N_17801);
nor U18099 (N_18099,N_17768,N_17614);
or U18100 (N_18100,N_17583,N_17754);
nand U18101 (N_18101,N_17921,N_17505);
nor U18102 (N_18102,N_17556,N_17642);
or U18103 (N_18103,N_17954,N_17781);
nor U18104 (N_18104,N_17926,N_17855);
xnor U18105 (N_18105,N_17873,N_17903);
and U18106 (N_18106,N_17888,N_17568);
nor U18107 (N_18107,N_17507,N_17593);
or U18108 (N_18108,N_17852,N_17675);
xor U18109 (N_18109,N_17718,N_17503);
or U18110 (N_18110,N_17820,N_17808);
xnor U18111 (N_18111,N_17893,N_17608);
nor U18112 (N_18112,N_17591,N_17717);
nor U18113 (N_18113,N_17993,N_17673);
nand U18114 (N_18114,N_17785,N_17601);
and U18115 (N_18115,N_17669,N_17599);
or U18116 (N_18116,N_17548,N_17982);
xor U18117 (N_18117,N_17681,N_17697);
xnor U18118 (N_18118,N_17799,N_17597);
nor U18119 (N_18119,N_17810,N_17607);
xor U18120 (N_18120,N_17971,N_17544);
xnor U18121 (N_18121,N_17868,N_17960);
or U18122 (N_18122,N_17953,N_17603);
or U18123 (N_18123,N_17706,N_17945);
nand U18124 (N_18124,N_17571,N_17871);
nor U18125 (N_18125,N_17802,N_17707);
xnor U18126 (N_18126,N_17793,N_17774);
or U18127 (N_18127,N_17896,N_17922);
xor U18128 (N_18128,N_17741,N_17841);
and U18129 (N_18129,N_17961,N_17914);
xor U18130 (N_18130,N_17941,N_17626);
and U18131 (N_18131,N_17756,N_17685);
nand U18132 (N_18132,N_17628,N_17653);
or U18133 (N_18133,N_17640,N_17778);
xor U18134 (N_18134,N_17859,N_17719);
or U18135 (N_18135,N_17747,N_17930);
and U18136 (N_18136,N_17904,N_17845);
nor U18137 (N_18137,N_17933,N_17977);
or U18138 (N_18138,N_17661,N_17766);
or U18139 (N_18139,N_17743,N_17573);
nand U18140 (N_18140,N_17862,N_17539);
and U18141 (N_18141,N_17934,N_17950);
nand U18142 (N_18142,N_17932,N_17696);
nand U18143 (N_18143,N_17549,N_17925);
nor U18144 (N_18144,N_17708,N_17730);
or U18145 (N_18145,N_17686,N_17612);
xnor U18146 (N_18146,N_17598,N_17735);
nand U18147 (N_18147,N_17895,N_17621);
and U18148 (N_18148,N_17504,N_17874);
xor U18149 (N_18149,N_17899,N_17973);
and U18150 (N_18150,N_17948,N_17905);
nor U18151 (N_18151,N_17698,N_17937);
or U18152 (N_18152,N_17745,N_17866);
and U18153 (N_18153,N_17695,N_17835);
nor U18154 (N_18154,N_17878,N_17770);
and U18155 (N_18155,N_17538,N_17805);
or U18156 (N_18156,N_17836,N_17664);
and U18157 (N_18157,N_17627,N_17674);
xor U18158 (N_18158,N_17823,N_17725);
nor U18159 (N_18159,N_17972,N_17748);
nor U18160 (N_18160,N_17877,N_17861);
xnor U18161 (N_18161,N_17547,N_17943);
or U18162 (N_18162,N_17915,N_17630);
nand U18163 (N_18163,N_17502,N_17789);
and U18164 (N_18164,N_17531,N_17751);
and U18165 (N_18165,N_17704,N_17911);
nand U18166 (N_18166,N_17850,N_17772);
xor U18167 (N_18167,N_17749,N_17632);
nand U18168 (N_18168,N_17967,N_17869);
or U18169 (N_18169,N_17812,N_17955);
nand U18170 (N_18170,N_17594,N_17901);
and U18171 (N_18171,N_17879,N_17501);
nor U18172 (N_18172,N_17589,N_17990);
xnor U18173 (N_18173,N_17816,N_17851);
nor U18174 (N_18174,N_17650,N_17898);
and U18175 (N_18175,N_17528,N_17604);
nand U18176 (N_18176,N_17907,N_17615);
or U18177 (N_18177,N_17792,N_17639);
or U18178 (N_18178,N_17897,N_17679);
nor U18179 (N_18179,N_17553,N_17572);
and U18180 (N_18180,N_17872,N_17579);
or U18181 (N_18181,N_17790,N_17682);
nand U18182 (N_18182,N_17819,N_17825);
nand U18183 (N_18183,N_17827,N_17788);
nor U18184 (N_18184,N_17576,N_17759);
or U18185 (N_18185,N_17731,N_17857);
and U18186 (N_18186,N_17923,N_17985);
and U18187 (N_18187,N_17566,N_17641);
xor U18188 (N_18188,N_17920,N_17865);
xor U18189 (N_18189,N_17863,N_17600);
nand U18190 (N_18190,N_17652,N_17645);
xor U18191 (N_18191,N_17546,N_17944);
or U18192 (N_18192,N_17806,N_17957);
nand U18193 (N_18193,N_17978,N_17709);
nand U18194 (N_18194,N_17509,N_17858);
and U18195 (N_18195,N_17678,N_17782);
nand U18196 (N_18196,N_17811,N_17596);
xnor U18197 (N_18197,N_17963,N_17854);
xnor U18198 (N_18198,N_17853,N_17908);
or U18199 (N_18199,N_17987,N_17881);
or U18200 (N_18200,N_17647,N_17964);
xor U18201 (N_18201,N_17619,N_17882);
xnor U18202 (N_18202,N_17762,N_17752);
nor U18203 (N_18203,N_17856,N_17848);
or U18204 (N_18204,N_17817,N_17649);
nor U18205 (N_18205,N_17870,N_17880);
or U18206 (N_18206,N_17746,N_17891);
nand U18207 (N_18207,N_17636,N_17609);
nand U18208 (N_18208,N_17520,N_17672);
nor U18209 (N_18209,N_17775,N_17534);
and U18210 (N_18210,N_17643,N_17787);
and U18211 (N_18211,N_17512,N_17723);
nor U18212 (N_18212,N_17886,N_17522);
nor U18213 (N_18213,N_17884,N_17518);
or U18214 (N_18214,N_17804,N_17994);
nor U18215 (N_18215,N_17567,N_17671);
nor U18216 (N_18216,N_17525,N_17574);
xor U18217 (N_18217,N_17824,N_17958);
or U18218 (N_18218,N_17542,N_17739);
or U18219 (N_18219,N_17867,N_17970);
nor U18220 (N_18220,N_17928,N_17618);
xnor U18221 (N_18221,N_17800,N_17555);
nand U18222 (N_18222,N_17771,N_17997);
nand U18223 (N_18223,N_17924,N_17764);
nand U18224 (N_18224,N_17890,N_17554);
nand U18225 (N_18225,N_17988,N_17796);
or U18226 (N_18226,N_17629,N_17506);
or U18227 (N_18227,N_17637,N_17876);
nand U18228 (N_18228,N_17949,N_17740);
nor U18229 (N_18229,N_17726,N_17541);
xor U18230 (N_18230,N_17581,N_17617);
and U18231 (N_18231,N_17919,N_17605);
nand U18232 (N_18232,N_17537,N_17952);
and U18233 (N_18233,N_17724,N_17979);
or U18234 (N_18234,N_17798,N_17577);
nand U18235 (N_18235,N_17838,N_17727);
xor U18236 (N_18236,N_17680,N_17912);
and U18237 (N_18237,N_17938,N_17828);
or U18238 (N_18238,N_17761,N_17959);
and U18239 (N_18239,N_17616,N_17818);
and U18240 (N_18240,N_17722,N_17602);
nor U18241 (N_18241,N_17595,N_17794);
nand U18242 (N_18242,N_17613,N_17996);
nor U18243 (N_18243,N_17536,N_17543);
nand U18244 (N_18244,N_17975,N_17894);
xnor U18245 (N_18245,N_17532,N_17936);
or U18246 (N_18246,N_17734,N_17700);
or U18247 (N_18247,N_17558,N_17826);
and U18248 (N_18248,N_17668,N_17918);
nand U18249 (N_18249,N_17968,N_17580);
or U18250 (N_18250,N_17697,N_17624);
or U18251 (N_18251,N_17540,N_17952);
nor U18252 (N_18252,N_17816,N_17930);
and U18253 (N_18253,N_17556,N_17529);
nor U18254 (N_18254,N_17621,N_17584);
nor U18255 (N_18255,N_17857,N_17955);
nand U18256 (N_18256,N_17964,N_17973);
or U18257 (N_18257,N_17763,N_17865);
xor U18258 (N_18258,N_17802,N_17517);
nand U18259 (N_18259,N_17700,N_17997);
and U18260 (N_18260,N_17585,N_17505);
nand U18261 (N_18261,N_17963,N_17859);
or U18262 (N_18262,N_17682,N_17888);
xnor U18263 (N_18263,N_17580,N_17616);
xnor U18264 (N_18264,N_17918,N_17869);
nor U18265 (N_18265,N_17987,N_17506);
nand U18266 (N_18266,N_17918,N_17728);
nand U18267 (N_18267,N_17926,N_17514);
xnor U18268 (N_18268,N_17546,N_17821);
nand U18269 (N_18269,N_17974,N_17862);
and U18270 (N_18270,N_17970,N_17750);
and U18271 (N_18271,N_17648,N_17581);
xor U18272 (N_18272,N_17743,N_17817);
nor U18273 (N_18273,N_17887,N_17704);
and U18274 (N_18274,N_17960,N_17667);
or U18275 (N_18275,N_17677,N_17756);
or U18276 (N_18276,N_17651,N_17535);
xor U18277 (N_18277,N_17500,N_17811);
xor U18278 (N_18278,N_17822,N_17985);
xor U18279 (N_18279,N_17718,N_17560);
or U18280 (N_18280,N_17650,N_17617);
xnor U18281 (N_18281,N_17908,N_17529);
or U18282 (N_18282,N_17834,N_17634);
xnor U18283 (N_18283,N_17790,N_17589);
and U18284 (N_18284,N_17803,N_17877);
xnor U18285 (N_18285,N_17551,N_17502);
nor U18286 (N_18286,N_17706,N_17921);
or U18287 (N_18287,N_17648,N_17889);
xor U18288 (N_18288,N_17997,N_17546);
xor U18289 (N_18289,N_17662,N_17586);
and U18290 (N_18290,N_17691,N_17560);
and U18291 (N_18291,N_17707,N_17962);
nor U18292 (N_18292,N_17939,N_17877);
and U18293 (N_18293,N_17579,N_17993);
nor U18294 (N_18294,N_17554,N_17601);
and U18295 (N_18295,N_17617,N_17766);
nand U18296 (N_18296,N_17896,N_17921);
xor U18297 (N_18297,N_17520,N_17874);
nor U18298 (N_18298,N_17651,N_17565);
or U18299 (N_18299,N_17710,N_17735);
and U18300 (N_18300,N_17704,N_17836);
nor U18301 (N_18301,N_17981,N_17530);
nor U18302 (N_18302,N_17946,N_17717);
nand U18303 (N_18303,N_17673,N_17907);
nand U18304 (N_18304,N_17666,N_17508);
xnor U18305 (N_18305,N_17726,N_17815);
or U18306 (N_18306,N_17818,N_17508);
and U18307 (N_18307,N_17673,N_17879);
or U18308 (N_18308,N_17926,N_17691);
or U18309 (N_18309,N_17661,N_17641);
or U18310 (N_18310,N_17523,N_17860);
or U18311 (N_18311,N_17908,N_17961);
and U18312 (N_18312,N_17817,N_17691);
nor U18313 (N_18313,N_17620,N_17809);
and U18314 (N_18314,N_17548,N_17936);
nand U18315 (N_18315,N_17822,N_17970);
and U18316 (N_18316,N_17862,N_17942);
nor U18317 (N_18317,N_17771,N_17502);
and U18318 (N_18318,N_17847,N_17518);
xor U18319 (N_18319,N_17610,N_17980);
nor U18320 (N_18320,N_17572,N_17946);
xor U18321 (N_18321,N_17503,N_17952);
nand U18322 (N_18322,N_17943,N_17992);
xor U18323 (N_18323,N_17614,N_17569);
xnor U18324 (N_18324,N_17528,N_17630);
nor U18325 (N_18325,N_17534,N_17702);
and U18326 (N_18326,N_17861,N_17633);
nor U18327 (N_18327,N_17858,N_17611);
xnor U18328 (N_18328,N_17658,N_17653);
xor U18329 (N_18329,N_17851,N_17786);
nand U18330 (N_18330,N_17696,N_17533);
nand U18331 (N_18331,N_17838,N_17531);
nand U18332 (N_18332,N_17606,N_17539);
nor U18333 (N_18333,N_17528,N_17658);
or U18334 (N_18334,N_17633,N_17892);
or U18335 (N_18335,N_17619,N_17808);
or U18336 (N_18336,N_17645,N_17582);
and U18337 (N_18337,N_17803,N_17668);
nand U18338 (N_18338,N_17877,N_17967);
or U18339 (N_18339,N_17961,N_17844);
or U18340 (N_18340,N_17522,N_17550);
or U18341 (N_18341,N_17983,N_17991);
nand U18342 (N_18342,N_17555,N_17699);
nand U18343 (N_18343,N_17543,N_17545);
nand U18344 (N_18344,N_17789,N_17578);
and U18345 (N_18345,N_17506,N_17592);
nor U18346 (N_18346,N_17862,N_17976);
xor U18347 (N_18347,N_17622,N_17860);
or U18348 (N_18348,N_17861,N_17945);
nor U18349 (N_18349,N_17746,N_17934);
and U18350 (N_18350,N_17745,N_17937);
xor U18351 (N_18351,N_17970,N_17861);
and U18352 (N_18352,N_17732,N_17997);
nand U18353 (N_18353,N_17652,N_17522);
and U18354 (N_18354,N_17903,N_17828);
or U18355 (N_18355,N_17551,N_17947);
or U18356 (N_18356,N_17956,N_17968);
xnor U18357 (N_18357,N_17977,N_17982);
nor U18358 (N_18358,N_17869,N_17570);
or U18359 (N_18359,N_17670,N_17549);
nor U18360 (N_18360,N_17522,N_17626);
and U18361 (N_18361,N_17554,N_17595);
nand U18362 (N_18362,N_17675,N_17597);
or U18363 (N_18363,N_17641,N_17760);
and U18364 (N_18364,N_17700,N_17693);
nand U18365 (N_18365,N_17920,N_17972);
and U18366 (N_18366,N_17684,N_17890);
nand U18367 (N_18367,N_17906,N_17578);
and U18368 (N_18368,N_17814,N_17678);
nor U18369 (N_18369,N_17981,N_17872);
or U18370 (N_18370,N_17959,N_17738);
or U18371 (N_18371,N_17863,N_17865);
or U18372 (N_18372,N_17858,N_17532);
nor U18373 (N_18373,N_17998,N_17523);
nand U18374 (N_18374,N_17631,N_17790);
and U18375 (N_18375,N_17538,N_17722);
nand U18376 (N_18376,N_17975,N_17561);
nor U18377 (N_18377,N_17748,N_17933);
nand U18378 (N_18378,N_17803,N_17521);
and U18379 (N_18379,N_17917,N_17706);
nor U18380 (N_18380,N_17762,N_17804);
nor U18381 (N_18381,N_17985,N_17735);
xnor U18382 (N_18382,N_17530,N_17918);
nor U18383 (N_18383,N_17637,N_17524);
or U18384 (N_18384,N_17537,N_17871);
nand U18385 (N_18385,N_17607,N_17688);
or U18386 (N_18386,N_17889,N_17810);
nand U18387 (N_18387,N_17717,N_17949);
xnor U18388 (N_18388,N_17762,N_17774);
or U18389 (N_18389,N_17628,N_17754);
xnor U18390 (N_18390,N_17741,N_17828);
nor U18391 (N_18391,N_17877,N_17736);
or U18392 (N_18392,N_17526,N_17949);
xor U18393 (N_18393,N_17537,N_17710);
nand U18394 (N_18394,N_17588,N_17753);
nand U18395 (N_18395,N_17924,N_17807);
or U18396 (N_18396,N_17615,N_17941);
xnor U18397 (N_18397,N_17585,N_17714);
and U18398 (N_18398,N_17868,N_17870);
nand U18399 (N_18399,N_17938,N_17594);
nor U18400 (N_18400,N_17716,N_17636);
xnor U18401 (N_18401,N_17787,N_17987);
nand U18402 (N_18402,N_17878,N_17785);
and U18403 (N_18403,N_17529,N_17573);
and U18404 (N_18404,N_17767,N_17527);
nor U18405 (N_18405,N_17711,N_17833);
or U18406 (N_18406,N_17883,N_17790);
and U18407 (N_18407,N_17509,N_17758);
nand U18408 (N_18408,N_17658,N_17532);
nand U18409 (N_18409,N_17702,N_17583);
and U18410 (N_18410,N_17832,N_17948);
and U18411 (N_18411,N_17714,N_17733);
xor U18412 (N_18412,N_17612,N_17611);
nand U18413 (N_18413,N_17635,N_17734);
and U18414 (N_18414,N_17656,N_17690);
xnor U18415 (N_18415,N_17636,N_17748);
xnor U18416 (N_18416,N_17772,N_17942);
and U18417 (N_18417,N_17514,N_17735);
and U18418 (N_18418,N_17926,N_17591);
and U18419 (N_18419,N_17780,N_17878);
xor U18420 (N_18420,N_17576,N_17715);
nor U18421 (N_18421,N_17623,N_17929);
or U18422 (N_18422,N_17943,N_17635);
nor U18423 (N_18423,N_17731,N_17764);
xor U18424 (N_18424,N_17811,N_17581);
xor U18425 (N_18425,N_17873,N_17617);
and U18426 (N_18426,N_17802,N_17698);
and U18427 (N_18427,N_17866,N_17693);
or U18428 (N_18428,N_17992,N_17668);
and U18429 (N_18429,N_17795,N_17800);
nor U18430 (N_18430,N_17629,N_17689);
or U18431 (N_18431,N_17790,N_17608);
xor U18432 (N_18432,N_17962,N_17567);
nand U18433 (N_18433,N_17965,N_17567);
xnor U18434 (N_18434,N_17572,N_17920);
and U18435 (N_18435,N_17705,N_17775);
or U18436 (N_18436,N_17507,N_17657);
nor U18437 (N_18437,N_17847,N_17713);
nor U18438 (N_18438,N_17704,N_17658);
and U18439 (N_18439,N_17833,N_17689);
and U18440 (N_18440,N_17686,N_17556);
or U18441 (N_18441,N_17942,N_17945);
and U18442 (N_18442,N_17686,N_17801);
nand U18443 (N_18443,N_17802,N_17706);
and U18444 (N_18444,N_17699,N_17905);
xor U18445 (N_18445,N_17612,N_17928);
and U18446 (N_18446,N_17535,N_17792);
and U18447 (N_18447,N_17939,N_17973);
xor U18448 (N_18448,N_17659,N_17751);
xor U18449 (N_18449,N_17610,N_17761);
or U18450 (N_18450,N_17982,N_17541);
nand U18451 (N_18451,N_17980,N_17740);
and U18452 (N_18452,N_17761,N_17570);
nand U18453 (N_18453,N_17546,N_17903);
nand U18454 (N_18454,N_17897,N_17659);
or U18455 (N_18455,N_17889,N_17990);
and U18456 (N_18456,N_17706,N_17825);
xnor U18457 (N_18457,N_17996,N_17921);
nor U18458 (N_18458,N_17847,N_17553);
xor U18459 (N_18459,N_17961,N_17571);
or U18460 (N_18460,N_17542,N_17727);
nand U18461 (N_18461,N_17686,N_17722);
or U18462 (N_18462,N_17713,N_17993);
xnor U18463 (N_18463,N_17788,N_17588);
nor U18464 (N_18464,N_17880,N_17786);
and U18465 (N_18465,N_17890,N_17607);
or U18466 (N_18466,N_17636,N_17777);
nor U18467 (N_18467,N_17724,N_17973);
and U18468 (N_18468,N_17830,N_17781);
and U18469 (N_18469,N_17856,N_17684);
or U18470 (N_18470,N_17504,N_17557);
nor U18471 (N_18471,N_17553,N_17898);
nand U18472 (N_18472,N_17993,N_17859);
or U18473 (N_18473,N_17773,N_17575);
or U18474 (N_18474,N_17837,N_17576);
nor U18475 (N_18475,N_17788,N_17611);
xnor U18476 (N_18476,N_17651,N_17939);
xor U18477 (N_18477,N_17511,N_17566);
xor U18478 (N_18478,N_17725,N_17567);
and U18479 (N_18479,N_17735,N_17990);
xnor U18480 (N_18480,N_17829,N_17880);
or U18481 (N_18481,N_17905,N_17723);
nor U18482 (N_18482,N_17605,N_17890);
nand U18483 (N_18483,N_17886,N_17573);
xor U18484 (N_18484,N_17522,N_17685);
nand U18485 (N_18485,N_17614,N_17948);
or U18486 (N_18486,N_17968,N_17925);
xor U18487 (N_18487,N_17543,N_17637);
nand U18488 (N_18488,N_17847,N_17992);
xnor U18489 (N_18489,N_17816,N_17831);
nor U18490 (N_18490,N_17559,N_17848);
xor U18491 (N_18491,N_17578,N_17769);
nand U18492 (N_18492,N_17748,N_17894);
nor U18493 (N_18493,N_17926,N_17868);
and U18494 (N_18494,N_17749,N_17868);
and U18495 (N_18495,N_17802,N_17909);
nand U18496 (N_18496,N_17815,N_17821);
or U18497 (N_18497,N_17871,N_17937);
or U18498 (N_18498,N_17578,N_17677);
or U18499 (N_18499,N_17929,N_17822);
xnor U18500 (N_18500,N_18467,N_18276);
or U18501 (N_18501,N_18056,N_18093);
and U18502 (N_18502,N_18493,N_18309);
nor U18503 (N_18503,N_18216,N_18104);
xor U18504 (N_18504,N_18453,N_18429);
nand U18505 (N_18505,N_18384,N_18103);
nand U18506 (N_18506,N_18149,N_18495);
nor U18507 (N_18507,N_18335,N_18421);
or U18508 (N_18508,N_18154,N_18360);
nor U18509 (N_18509,N_18424,N_18148);
and U18510 (N_18510,N_18333,N_18497);
nand U18511 (N_18511,N_18087,N_18465);
and U18512 (N_18512,N_18491,N_18278);
and U18513 (N_18513,N_18219,N_18184);
xor U18514 (N_18514,N_18288,N_18274);
nor U18515 (N_18515,N_18176,N_18248);
or U18516 (N_18516,N_18237,N_18372);
nor U18517 (N_18517,N_18272,N_18256);
or U18518 (N_18518,N_18064,N_18458);
xnor U18519 (N_18519,N_18426,N_18128);
and U18520 (N_18520,N_18350,N_18286);
and U18521 (N_18521,N_18224,N_18327);
and U18522 (N_18522,N_18196,N_18273);
nor U18523 (N_18523,N_18391,N_18404);
xor U18524 (N_18524,N_18410,N_18314);
nor U18525 (N_18525,N_18057,N_18137);
nor U18526 (N_18526,N_18401,N_18341);
nand U18527 (N_18527,N_18357,N_18012);
xor U18528 (N_18528,N_18270,N_18459);
nor U18529 (N_18529,N_18441,N_18030);
or U18530 (N_18530,N_18476,N_18390);
xnor U18531 (N_18531,N_18460,N_18481);
and U18532 (N_18532,N_18373,N_18385);
nor U18533 (N_18533,N_18435,N_18340);
xnor U18534 (N_18534,N_18298,N_18092);
xnor U18535 (N_18535,N_18299,N_18455);
nor U18536 (N_18536,N_18070,N_18080);
or U18537 (N_18537,N_18222,N_18046);
or U18538 (N_18538,N_18236,N_18206);
nand U18539 (N_18539,N_18017,N_18359);
nor U18540 (N_18540,N_18485,N_18312);
and U18541 (N_18541,N_18140,N_18022);
and U18542 (N_18542,N_18258,N_18339);
or U18543 (N_18543,N_18488,N_18178);
and U18544 (N_18544,N_18162,N_18132);
nand U18545 (N_18545,N_18026,N_18136);
nor U18546 (N_18546,N_18461,N_18055);
nand U18547 (N_18547,N_18448,N_18316);
nor U18548 (N_18548,N_18221,N_18079);
nor U18549 (N_18549,N_18042,N_18432);
nor U18550 (N_18550,N_18118,N_18457);
nand U18551 (N_18551,N_18254,N_18307);
nand U18552 (N_18552,N_18388,N_18439);
nand U18553 (N_18553,N_18031,N_18315);
nand U18554 (N_18554,N_18336,N_18356);
or U18555 (N_18555,N_18306,N_18076);
nand U18556 (N_18556,N_18331,N_18018);
nor U18557 (N_18557,N_18472,N_18308);
xnor U18558 (N_18558,N_18265,N_18139);
and U18559 (N_18559,N_18089,N_18067);
and U18560 (N_18560,N_18423,N_18071);
and U18561 (N_18561,N_18209,N_18004);
nor U18562 (N_18562,N_18183,N_18301);
nor U18563 (N_18563,N_18444,N_18157);
nor U18564 (N_18564,N_18257,N_18190);
or U18565 (N_18565,N_18003,N_18198);
and U18566 (N_18566,N_18297,N_18105);
xor U18567 (N_18567,N_18060,N_18201);
and U18568 (N_18568,N_18399,N_18470);
and U18569 (N_18569,N_18191,N_18440);
xnor U18570 (N_18570,N_18353,N_18121);
or U18571 (N_18571,N_18407,N_18231);
nor U18572 (N_18572,N_18217,N_18047);
nor U18573 (N_18573,N_18477,N_18235);
or U18574 (N_18574,N_18085,N_18016);
or U18575 (N_18575,N_18371,N_18084);
xnor U18576 (N_18576,N_18326,N_18434);
nor U18577 (N_18577,N_18318,N_18466);
xnor U18578 (N_18578,N_18304,N_18129);
xnor U18579 (N_18579,N_18225,N_18040);
or U18580 (N_18580,N_18468,N_18120);
or U18581 (N_18581,N_18073,N_18048);
nand U18582 (N_18582,N_18065,N_18451);
or U18583 (N_18583,N_18271,N_18358);
xor U18584 (N_18584,N_18364,N_18063);
nand U18585 (N_18585,N_18077,N_18226);
xor U18586 (N_18586,N_18486,N_18264);
or U18587 (N_18587,N_18292,N_18269);
and U18588 (N_18588,N_18430,N_18143);
or U18589 (N_18589,N_18113,N_18352);
and U18590 (N_18590,N_18066,N_18167);
nand U18591 (N_18591,N_18034,N_18054);
xnor U18592 (N_18592,N_18091,N_18395);
or U18593 (N_18593,N_18002,N_18006);
xnor U18594 (N_18594,N_18291,N_18011);
nor U18595 (N_18595,N_18379,N_18377);
and U18596 (N_18596,N_18412,N_18348);
nor U18597 (N_18597,N_18122,N_18411);
xor U18598 (N_18598,N_18069,N_18363);
and U18599 (N_18599,N_18214,N_18347);
nor U18600 (N_18600,N_18233,N_18417);
nand U18601 (N_18601,N_18409,N_18266);
nor U18602 (N_18602,N_18365,N_18096);
and U18603 (N_18603,N_18037,N_18124);
xor U18604 (N_18604,N_18294,N_18205);
or U18605 (N_18605,N_18244,N_18422);
or U18606 (N_18606,N_18389,N_18338);
xnor U18607 (N_18607,N_18160,N_18075);
or U18608 (N_18608,N_18397,N_18494);
xor U18609 (N_18609,N_18151,N_18310);
nand U18610 (N_18610,N_18199,N_18193);
nor U18611 (N_18611,N_18378,N_18419);
and U18612 (N_18612,N_18044,N_18393);
and U18613 (N_18613,N_18131,N_18249);
xor U18614 (N_18614,N_18108,N_18456);
nor U18615 (N_18615,N_18492,N_18181);
and U18616 (N_18616,N_18164,N_18452);
nor U18617 (N_18617,N_18230,N_18380);
xnor U18618 (N_18618,N_18387,N_18175);
nor U18619 (N_18619,N_18114,N_18133);
or U18620 (N_18620,N_18433,N_18496);
nand U18621 (N_18621,N_18475,N_18015);
and U18622 (N_18622,N_18437,N_18293);
nand U18623 (N_18623,N_18289,N_18130);
xor U18624 (N_18624,N_18414,N_18268);
nand U18625 (N_18625,N_18473,N_18396);
xnor U18626 (N_18626,N_18329,N_18438);
nand U18627 (N_18627,N_18058,N_18368);
and U18628 (N_18628,N_18163,N_18119);
xor U18629 (N_18629,N_18100,N_18282);
nor U18630 (N_18630,N_18462,N_18345);
xnor U18631 (N_18631,N_18285,N_18007);
nand U18632 (N_18632,N_18402,N_18499);
nor U18633 (N_18633,N_18349,N_18498);
xor U18634 (N_18634,N_18482,N_18074);
and U18635 (N_18635,N_18319,N_18279);
and U18636 (N_18636,N_18223,N_18062);
xnor U18637 (N_18637,N_18094,N_18207);
and U18638 (N_18638,N_18386,N_18204);
and U18639 (N_18639,N_18099,N_18381);
or U18640 (N_18640,N_18185,N_18019);
xor U18641 (N_18641,N_18445,N_18173);
xor U18642 (N_18642,N_18090,N_18369);
nand U18643 (N_18643,N_18262,N_18394);
xnor U18644 (N_18644,N_18382,N_18180);
xnor U18645 (N_18645,N_18246,N_18059);
or U18646 (N_18646,N_18449,N_18035);
and U18647 (N_18647,N_18227,N_18053);
xor U18648 (N_18648,N_18420,N_18251);
nand U18649 (N_18649,N_18200,N_18234);
nor U18650 (N_18650,N_18325,N_18155);
or U18651 (N_18651,N_18375,N_18068);
nand U18652 (N_18652,N_18111,N_18024);
and U18653 (N_18653,N_18186,N_18147);
nand U18654 (N_18654,N_18117,N_18480);
or U18655 (N_18655,N_18194,N_18280);
and U18656 (N_18656,N_18355,N_18436);
or U18657 (N_18657,N_18171,N_18283);
xor U18658 (N_18658,N_18328,N_18490);
xnor U18659 (N_18659,N_18195,N_18145);
and U18660 (N_18660,N_18049,N_18484);
xnor U18661 (N_18661,N_18115,N_18169);
and U18662 (N_18662,N_18259,N_18305);
nand U18663 (N_18663,N_18220,N_18045);
nand U18664 (N_18664,N_18088,N_18474);
and U18665 (N_18665,N_18478,N_18405);
and U18666 (N_18666,N_18450,N_18261);
nand U18667 (N_18667,N_18161,N_18083);
or U18668 (N_18668,N_18343,N_18317);
or U18669 (N_18669,N_18082,N_18281);
or U18670 (N_18670,N_18052,N_18241);
nand U18671 (N_18671,N_18418,N_18005);
and U18672 (N_18672,N_18142,N_18177);
xor U18673 (N_18673,N_18008,N_18416);
xnor U18674 (N_18674,N_18141,N_18218);
xor U18675 (N_18675,N_18208,N_18020);
nor U18676 (N_18676,N_18158,N_18351);
and U18677 (N_18677,N_18428,N_18028);
nand U18678 (N_18678,N_18366,N_18123);
nor U18679 (N_18679,N_18275,N_18098);
and U18680 (N_18680,N_18027,N_18392);
or U18681 (N_18681,N_18243,N_18267);
nand U18682 (N_18682,N_18144,N_18406);
nor U18683 (N_18683,N_18156,N_18346);
or U18684 (N_18684,N_18043,N_18296);
nor U18685 (N_18685,N_18361,N_18110);
or U18686 (N_18686,N_18116,N_18010);
xnor U18687 (N_18687,N_18443,N_18166);
and U18688 (N_18688,N_18039,N_18403);
or U18689 (N_18689,N_18321,N_18295);
or U18690 (N_18690,N_18000,N_18284);
nor U18691 (N_18691,N_18442,N_18081);
and U18692 (N_18692,N_18240,N_18311);
and U18693 (N_18693,N_18202,N_18138);
xor U18694 (N_18694,N_18400,N_18078);
and U18695 (N_18695,N_18165,N_18126);
nor U18696 (N_18696,N_18408,N_18242);
or U18697 (N_18697,N_18431,N_18332);
and U18698 (N_18698,N_18250,N_18300);
nand U18699 (N_18699,N_18106,N_18187);
xnor U18700 (N_18700,N_18228,N_18050);
xor U18701 (N_18701,N_18189,N_18479);
and U18702 (N_18702,N_18179,N_18029);
nand U18703 (N_18703,N_18152,N_18383);
xnor U18704 (N_18704,N_18260,N_18483);
xnor U18705 (N_18705,N_18153,N_18239);
or U18706 (N_18706,N_18324,N_18023);
nor U18707 (N_18707,N_18446,N_18303);
nand U18708 (N_18708,N_18376,N_18112);
xor U18709 (N_18709,N_18150,N_18101);
and U18710 (N_18710,N_18398,N_18255);
nand U18711 (N_18711,N_18051,N_18213);
or U18712 (N_18712,N_18302,N_18463);
xor U18713 (N_18713,N_18102,N_18447);
or U18714 (N_18714,N_18095,N_18159);
xnor U18715 (N_18715,N_18252,N_18367);
or U18716 (N_18716,N_18127,N_18182);
and U18717 (N_18717,N_18464,N_18086);
and U18718 (N_18718,N_18013,N_18320);
xnor U18719 (N_18719,N_18146,N_18097);
xor U18720 (N_18720,N_18277,N_18009);
and U18721 (N_18721,N_18203,N_18415);
nand U18722 (N_18722,N_18021,N_18174);
and U18723 (N_18723,N_18354,N_18210);
and U18724 (N_18724,N_18107,N_18229);
xor U18725 (N_18725,N_18489,N_18425);
nor U18726 (N_18726,N_18168,N_18041);
nor U18727 (N_18727,N_18427,N_18036);
or U18728 (N_18728,N_18287,N_18334);
xor U18729 (N_18729,N_18263,N_18033);
nand U18730 (N_18730,N_18362,N_18170);
nor U18731 (N_18731,N_18025,N_18038);
and U18732 (N_18732,N_18469,N_18001);
or U18733 (N_18733,N_18313,N_18061);
nor U18734 (N_18734,N_18232,N_18109);
xnor U18735 (N_18735,N_18323,N_18188);
xor U18736 (N_18736,N_18014,N_18454);
xor U18737 (N_18737,N_18212,N_18413);
or U18738 (N_18738,N_18290,N_18192);
or U18739 (N_18739,N_18370,N_18135);
and U18740 (N_18740,N_18471,N_18072);
nand U18741 (N_18741,N_18125,N_18253);
nor U18742 (N_18742,N_18197,N_18211);
nand U18743 (N_18743,N_18245,N_18247);
or U18744 (N_18744,N_18342,N_18337);
nor U18745 (N_18745,N_18215,N_18134);
xnor U18746 (N_18746,N_18032,N_18172);
nand U18747 (N_18747,N_18322,N_18374);
nor U18748 (N_18748,N_18330,N_18344);
xor U18749 (N_18749,N_18487,N_18238);
and U18750 (N_18750,N_18100,N_18419);
xnor U18751 (N_18751,N_18244,N_18337);
nor U18752 (N_18752,N_18411,N_18258);
nand U18753 (N_18753,N_18409,N_18332);
nor U18754 (N_18754,N_18017,N_18187);
and U18755 (N_18755,N_18037,N_18234);
nand U18756 (N_18756,N_18275,N_18198);
or U18757 (N_18757,N_18326,N_18458);
xnor U18758 (N_18758,N_18041,N_18305);
nand U18759 (N_18759,N_18140,N_18101);
nor U18760 (N_18760,N_18066,N_18017);
nand U18761 (N_18761,N_18024,N_18147);
nand U18762 (N_18762,N_18277,N_18139);
xor U18763 (N_18763,N_18347,N_18140);
nand U18764 (N_18764,N_18038,N_18292);
nor U18765 (N_18765,N_18416,N_18307);
xnor U18766 (N_18766,N_18324,N_18162);
xor U18767 (N_18767,N_18023,N_18362);
and U18768 (N_18768,N_18474,N_18244);
xor U18769 (N_18769,N_18343,N_18353);
xnor U18770 (N_18770,N_18139,N_18250);
nand U18771 (N_18771,N_18131,N_18224);
nand U18772 (N_18772,N_18006,N_18227);
nor U18773 (N_18773,N_18257,N_18098);
nand U18774 (N_18774,N_18163,N_18014);
xor U18775 (N_18775,N_18481,N_18295);
or U18776 (N_18776,N_18236,N_18390);
or U18777 (N_18777,N_18111,N_18389);
nand U18778 (N_18778,N_18047,N_18282);
nor U18779 (N_18779,N_18217,N_18255);
and U18780 (N_18780,N_18343,N_18330);
nand U18781 (N_18781,N_18416,N_18344);
and U18782 (N_18782,N_18352,N_18243);
or U18783 (N_18783,N_18233,N_18147);
nor U18784 (N_18784,N_18464,N_18315);
or U18785 (N_18785,N_18219,N_18015);
nor U18786 (N_18786,N_18317,N_18016);
nor U18787 (N_18787,N_18355,N_18271);
nor U18788 (N_18788,N_18237,N_18043);
or U18789 (N_18789,N_18260,N_18474);
xnor U18790 (N_18790,N_18312,N_18345);
xnor U18791 (N_18791,N_18416,N_18420);
or U18792 (N_18792,N_18075,N_18436);
xnor U18793 (N_18793,N_18107,N_18043);
nor U18794 (N_18794,N_18152,N_18433);
nand U18795 (N_18795,N_18087,N_18479);
nand U18796 (N_18796,N_18400,N_18482);
or U18797 (N_18797,N_18401,N_18018);
nand U18798 (N_18798,N_18478,N_18372);
nand U18799 (N_18799,N_18041,N_18023);
nand U18800 (N_18800,N_18104,N_18189);
xor U18801 (N_18801,N_18327,N_18188);
or U18802 (N_18802,N_18491,N_18349);
and U18803 (N_18803,N_18074,N_18131);
xnor U18804 (N_18804,N_18499,N_18185);
nand U18805 (N_18805,N_18117,N_18224);
nand U18806 (N_18806,N_18188,N_18426);
nand U18807 (N_18807,N_18172,N_18354);
xnor U18808 (N_18808,N_18023,N_18322);
and U18809 (N_18809,N_18438,N_18284);
or U18810 (N_18810,N_18077,N_18070);
xor U18811 (N_18811,N_18192,N_18278);
xor U18812 (N_18812,N_18387,N_18345);
and U18813 (N_18813,N_18236,N_18101);
xnor U18814 (N_18814,N_18189,N_18075);
xor U18815 (N_18815,N_18411,N_18441);
nand U18816 (N_18816,N_18119,N_18223);
or U18817 (N_18817,N_18368,N_18328);
xor U18818 (N_18818,N_18214,N_18406);
and U18819 (N_18819,N_18459,N_18207);
xor U18820 (N_18820,N_18298,N_18374);
nor U18821 (N_18821,N_18234,N_18034);
and U18822 (N_18822,N_18439,N_18099);
nor U18823 (N_18823,N_18199,N_18145);
xnor U18824 (N_18824,N_18230,N_18320);
nor U18825 (N_18825,N_18491,N_18221);
or U18826 (N_18826,N_18449,N_18160);
nand U18827 (N_18827,N_18416,N_18160);
nor U18828 (N_18828,N_18341,N_18440);
and U18829 (N_18829,N_18093,N_18117);
xor U18830 (N_18830,N_18113,N_18017);
and U18831 (N_18831,N_18218,N_18177);
xor U18832 (N_18832,N_18131,N_18200);
and U18833 (N_18833,N_18075,N_18296);
nand U18834 (N_18834,N_18139,N_18462);
and U18835 (N_18835,N_18419,N_18156);
nor U18836 (N_18836,N_18412,N_18103);
or U18837 (N_18837,N_18147,N_18448);
or U18838 (N_18838,N_18338,N_18063);
xnor U18839 (N_18839,N_18106,N_18479);
or U18840 (N_18840,N_18102,N_18397);
and U18841 (N_18841,N_18088,N_18471);
and U18842 (N_18842,N_18013,N_18171);
nor U18843 (N_18843,N_18356,N_18306);
or U18844 (N_18844,N_18241,N_18471);
nand U18845 (N_18845,N_18209,N_18307);
nand U18846 (N_18846,N_18334,N_18417);
nor U18847 (N_18847,N_18099,N_18361);
nor U18848 (N_18848,N_18389,N_18128);
nor U18849 (N_18849,N_18087,N_18253);
nand U18850 (N_18850,N_18259,N_18377);
nand U18851 (N_18851,N_18154,N_18243);
nand U18852 (N_18852,N_18253,N_18232);
xor U18853 (N_18853,N_18296,N_18401);
xor U18854 (N_18854,N_18357,N_18374);
and U18855 (N_18855,N_18477,N_18223);
nor U18856 (N_18856,N_18390,N_18085);
xnor U18857 (N_18857,N_18394,N_18293);
nand U18858 (N_18858,N_18377,N_18046);
nand U18859 (N_18859,N_18130,N_18444);
nand U18860 (N_18860,N_18334,N_18286);
nand U18861 (N_18861,N_18491,N_18138);
and U18862 (N_18862,N_18483,N_18490);
nand U18863 (N_18863,N_18446,N_18127);
and U18864 (N_18864,N_18171,N_18035);
and U18865 (N_18865,N_18185,N_18080);
or U18866 (N_18866,N_18499,N_18117);
or U18867 (N_18867,N_18068,N_18126);
xor U18868 (N_18868,N_18129,N_18142);
nand U18869 (N_18869,N_18410,N_18019);
nand U18870 (N_18870,N_18026,N_18091);
nor U18871 (N_18871,N_18420,N_18426);
nand U18872 (N_18872,N_18158,N_18176);
xnor U18873 (N_18873,N_18360,N_18376);
or U18874 (N_18874,N_18335,N_18266);
or U18875 (N_18875,N_18066,N_18135);
or U18876 (N_18876,N_18304,N_18371);
and U18877 (N_18877,N_18423,N_18324);
xor U18878 (N_18878,N_18015,N_18268);
xnor U18879 (N_18879,N_18103,N_18336);
xor U18880 (N_18880,N_18442,N_18438);
and U18881 (N_18881,N_18217,N_18029);
or U18882 (N_18882,N_18206,N_18411);
nor U18883 (N_18883,N_18144,N_18086);
or U18884 (N_18884,N_18256,N_18088);
or U18885 (N_18885,N_18004,N_18476);
nand U18886 (N_18886,N_18463,N_18400);
and U18887 (N_18887,N_18195,N_18487);
and U18888 (N_18888,N_18475,N_18300);
or U18889 (N_18889,N_18208,N_18180);
and U18890 (N_18890,N_18210,N_18128);
xor U18891 (N_18891,N_18076,N_18460);
nand U18892 (N_18892,N_18471,N_18025);
nor U18893 (N_18893,N_18209,N_18428);
xor U18894 (N_18894,N_18100,N_18245);
nand U18895 (N_18895,N_18310,N_18451);
and U18896 (N_18896,N_18423,N_18381);
nor U18897 (N_18897,N_18481,N_18039);
and U18898 (N_18898,N_18425,N_18273);
nor U18899 (N_18899,N_18349,N_18258);
xor U18900 (N_18900,N_18401,N_18294);
or U18901 (N_18901,N_18096,N_18293);
and U18902 (N_18902,N_18485,N_18288);
nor U18903 (N_18903,N_18232,N_18181);
or U18904 (N_18904,N_18302,N_18282);
xor U18905 (N_18905,N_18448,N_18381);
and U18906 (N_18906,N_18270,N_18479);
or U18907 (N_18907,N_18128,N_18046);
nand U18908 (N_18908,N_18138,N_18109);
and U18909 (N_18909,N_18181,N_18476);
nor U18910 (N_18910,N_18394,N_18065);
or U18911 (N_18911,N_18030,N_18452);
or U18912 (N_18912,N_18301,N_18361);
or U18913 (N_18913,N_18161,N_18022);
and U18914 (N_18914,N_18297,N_18156);
or U18915 (N_18915,N_18237,N_18119);
nand U18916 (N_18916,N_18451,N_18279);
nor U18917 (N_18917,N_18423,N_18232);
xnor U18918 (N_18918,N_18220,N_18186);
xnor U18919 (N_18919,N_18267,N_18154);
xnor U18920 (N_18920,N_18366,N_18296);
or U18921 (N_18921,N_18037,N_18130);
xor U18922 (N_18922,N_18201,N_18406);
xor U18923 (N_18923,N_18096,N_18457);
xnor U18924 (N_18924,N_18361,N_18305);
and U18925 (N_18925,N_18268,N_18201);
or U18926 (N_18926,N_18283,N_18492);
nor U18927 (N_18927,N_18127,N_18426);
nor U18928 (N_18928,N_18482,N_18068);
nand U18929 (N_18929,N_18469,N_18036);
or U18930 (N_18930,N_18486,N_18479);
and U18931 (N_18931,N_18181,N_18347);
nand U18932 (N_18932,N_18039,N_18452);
and U18933 (N_18933,N_18015,N_18484);
or U18934 (N_18934,N_18158,N_18175);
and U18935 (N_18935,N_18124,N_18253);
and U18936 (N_18936,N_18315,N_18129);
nor U18937 (N_18937,N_18265,N_18457);
or U18938 (N_18938,N_18303,N_18267);
nor U18939 (N_18939,N_18293,N_18086);
and U18940 (N_18940,N_18402,N_18070);
and U18941 (N_18941,N_18243,N_18105);
and U18942 (N_18942,N_18230,N_18128);
nand U18943 (N_18943,N_18300,N_18198);
xnor U18944 (N_18944,N_18092,N_18282);
xnor U18945 (N_18945,N_18373,N_18037);
xor U18946 (N_18946,N_18065,N_18017);
xnor U18947 (N_18947,N_18424,N_18055);
xor U18948 (N_18948,N_18134,N_18413);
nor U18949 (N_18949,N_18362,N_18229);
nand U18950 (N_18950,N_18030,N_18302);
and U18951 (N_18951,N_18081,N_18215);
and U18952 (N_18952,N_18324,N_18067);
nand U18953 (N_18953,N_18077,N_18299);
and U18954 (N_18954,N_18104,N_18202);
nand U18955 (N_18955,N_18284,N_18331);
and U18956 (N_18956,N_18363,N_18162);
and U18957 (N_18957,N_18302,N_18056);
and U18958 (N_18958,N_18055,N_18182);
nand U18959 (N_18959,N_18488,N_18149);
and U18960 (N_18960,N_18152,N_18059);
and U18961 (N_18961,N_18367,N_18219);
and U18962 (N_18962,N_18416,N_18152);
and U18963 (N_18963,N_18288,N_18013);
xor U18964 (N_18964,N_18151,N_18365);
nor U18965 (N_18965,N_18317,N_18254);
xor U18966 (N_18966,N_18451,N_18206);
or U18967 (N_18967,N_18045,N_18029);
and U18968 (N_18968,N_18174,N_18472);
and U18969 (N_18969,N_18134,N_18199);
nand U18970 (N_18970,N_18181,N_18091);
xnor U18971 (N_18971,N_18046,N_18276);
nor U18972 (N_18972,N_18045,N_18413);
nand U18973 (N_18973,N_18171,N_18311);
xor U18974 (N_18974,N_18077,N_18092);
and U18975 (N_18975,N_18271,N_18097);
xnor U18976 (N_18976,N_18304,N_18151);
and U18977 (N_18977,N_18334,N_18101);
xor U18978 (N_18978,N_18231,N_18464);
or U18979 (N_18979,N_18100,N_18425);
nand U18980 (N_18980,N_18054,N_18420);
nand U18981 (N_18981,N_18040,N_18246);
nand U18982 (N_18982,N_18042,N_18053);
or U18983 (N_18983,N_18441,N_18176);
xnor U18984 (N_18984,N_18286,N_18156);
nand U18985 (N_18985,N_18092,N_18176);
nand U18986 (N_18986,N_18013,N_18483);
and U18987 (N_18987,N_18253,N_18485);
and U18988 (N_18988,N_18400,N_18427);
xor U18989 (N_18989,N_18461,N_18270);
xor U18990 (N_18990,N_18064,N_18281);
xor U18991 (N_18991,N_18428,N_18124);
nand U18992 (N_18992,N_18477,N_18242);
and U18993 (N_18993,N_18277,N_18306);
and U18994 (N_18994,N_18092,N_18180);
xnor U18995 (N_18995,N_18410,N_18460);
and U18996 (N_18996,N_18116,N_18411);
nand U18997 (N_18997,N_18219,N_18151);
nand U18998 (N_18998,N_18171,N_18423);
xor U18999 (N_18999,N_18375,N_18366);
nand U19000 (N_19000,N_18633,N_18693);
nor U19001 (N_19001,N_18547,N_18824);
or U19002 (N_19002,N_18710,N_18570);
nor U19003 (N_19003,N_18535,N_18696);
or U19004 (N_19004,N_18516,N_18967);
or U19005 (N_19005,N_18524,N_18609);
nand U19006 (N_19006,N_18921,N_18652);
nor U19007 (N_19007,N_18725,N_18591);
nor U19008 (N_19008,N_18879,N_18762);
and U19009 (N_19009,N_18846,N_18529);
or U19010 (N_19010,N_18691,N_18690);
nand U19011 (N_19011,N_18893,N_18855);
and U19012 (N_19012,N_18955,N_18809);
xor U19013 (N_19013,N_18636,N_18913);
or U19014 (N_19014,N_18949,N_18757);
and U19015 (N_19015,N_18758,N_18706);
nand U19016 (N_19016,N_18601,N_18595);
nor U19017 (N_19017,N_18868,N_18898);
xnor U19018 (N_19018,N_18650,N_18894);
nand U19019 (N_19019,N_18683,N_18828);
or U19020 (N_19020,N_18927,N_18718);
and U19021 (N_19021,N_18843,N_18546);
xor U19022 (N_19022,N_18839,N_18986);
and U19023 (N_19023,N_18559,N_18517);
nor U19024 (N_19024,N_18996,N_18746);
and U19025 (N_19025,N_18637,N_18551);
nand U19026 (N_19026,N_18509,N_18848);
and U19027 (N_19027,N_18782,N_18643);
nor U19028 (N_19028,N_18751,N_18705);
and U19029 (N_19029,N_18803,N_18728);
nand U19030 (N_19030,N_18859,N_18656);
and U19031 (N_19031,N_18686,N_18985);
nand U19032 (N_19032,N_18947,N_18585);
nor U19033 (N_19033,N_18964,N_18805);
and U19034 (N_19034,N_18702,N_18647);
nor U19035 (N_19035,N_18765,N_18802);
or U19036 (N_19036,N_18932,N_18604);
and U19037 (N_19037,N_18826,N_18564);
and U19038 (N_19038,N_18670,N_18543);
and U19039 (N_19039,N_18588,N_18768);
xnor U19040 (N_19040,N_18612,N_18928);
and U19041 (N_19041,N_18919,N_18534);
nor U19042 (N_19042,N_18694,N_18668);
nor U19043 (N_19043,N_18922,N_18835);
or U19044 (N_19044,N_18734,N_18958);
or U19045 (N_19045,N_18811,N_18800);
and U19046 (N_19046,N_18515,N_18842);
or U19047 (N_19047,N_18605,N_18998);
xnor U19048 (N_19048,N_18733,N_18797);
and U19049 (N_19049,N_18862,N_18939);
or U19050 (N_19050,N_18885,N_18953);
nor U19051 (N_19051,N_18644,N_18738);
nand U19052 (N_19052,N_18801,N_18732);
xnor U19053 (N_19053,N_18889,N_18781);
nor U19054 (N_19054,N_18787,N_18677);
nand U19055 (N_19055,N_18852,N_18614);
nor U19056 (N_19056,N_18915,N_18657);
and U19057 (N_19057,N_18869,N_18989);
and U19058 (N_19058,N_18910,N_18825);
nand U19059 (N_19059,N_18638,N_18717);
nor U19060 (N_19060,N_18560,N_18674);
xnor U19061 (N_19061,N_18576,N_18739);
nor U19062 (N_19062,N_18945,N_18950);
xor U19063 (N_19063,N_18990,N_18908);
or U19064 (N_19064,N_18676,N_18619);
xnor U19065 (N_19065,N_18891,N_18960);
and U19066 (N_19066,N_18713,N_18844);
nand U19067 (N_19067,N_18571,N_18701);
xnor U19068 (N_19068,N_18562,N_18502);
or U19069 (N_19069,N_18769,N_18592);
and U19070 (N_19070,N_18997,N_18611);
xor U19071 (N_19071,N_18634,N_18978);
xor U19072 (N_19072,N_18533,N_18995);
or U19073 (N_19073,N_18572,N_18851);
or U19074 (N_19074,N_18749,N_18673);
or U19075 (N_19075,N_18549,N_18767);
nand U19076 (N_19076,N_18510,N_18711);
or U19077 (N_19077,N_18687,N_18622);
and U19078 (N_19078,N_18812,N_18860);
nand U19079 (N_19079,N_18902,N_18600);
nor U19080 (N_19080,N_18672,N_18658);
nand U19081 (N_19081,N_18682,N_18833);
nand U19082 (N_19082,N_18941,N_18807);
xnor U19083 (N_19083,N_18912,N_18630);
or U19084 (N_19084,N_18736,N_18943);
nor U19085 (N_19085,N_18590,N_18808);
nor U19086 (N_19086,N_18906,N_18830);
or U19087 (N_19087,N_18665,N_18987);
or U19088 (N_19088,N_18992,N_18581);
nand U19089 (N_19089,N_18936,N_18607);
and U19090 (N_19090,N_18956,N_18821);
and U19091 (N_19091,N_18961,N_18698);
or U19092 (N_19092,N_18911,N_18598);
xor U19093 (N_19093,N_18679,N_18721);
and U19094 (N_19094,N_18766,N_18895);
or U19095 (N_19095,N_18981,N_18924);
nand U19096 (N_19096,N_18608,N_18748);
and U19097 (N_19097,N_18680,N_18966);
and U19098 (N_19098,N_18525,N_18528);
nor U19099 (N_19099,N_18671,N_18730);
or U19100 (N_19100,N_18648,N_18716);
nand U19101 (N_19101,N_18849,N_18635);
nand U19102 (N_19102,N_18726,N_18715);
nor U19103 (N_19103,N_18610,N_18526);
nor U19104 (N_19104,N_18977,N_18669);
nor U19105 (N_19105,N_18583,N_18651);
nor U19106 (N_19106,N_18940,N_18937);
nor U19107 (N_19107,N_18582,N_18580);
and U19108 (N_19108,N_18503,N_18667);
nand U19109 (N_19109,N_18594,N_18563);
nor U19110 (N_19110,N_18586,N_18646);
xnor U19111 (N_19111,N_18999,N_18793);
nand U19112 (N_19112,N_18847,N_18678);
and U19113 (N_19113,N_18917,N_18541);
nand U19114 (N_19114,N_18740,N_18872);
nor U19115 (N_19115,N_18783,N_18625);
and U19116 (N_19116,N_18934,N_18786);
xor U19117 (N_19117,N_18946,N_18557);
nand U19118 (N_19118,N_18897,N_18831);
nor U19119 (N_19119,N_18756,N_18777);
nor U19120 (N_19120,N_18900,N_18500);
nand U19121 (N_19121,N_18602,N_18804);
xor U19122 (N_19122,N_18731,N_18621);
or U19123 (N_19123,N_18864,N_18511);
nor U19124 (N_19124,N_18703,N_18775);
nor U19125 (N_19125,N_18704,N_18699);
nor U19126 (N_19126,N_18615,N_18817);
nor U19127 (N_19127,N_18556,N_18791);
and U19128 (N_19128,N_18707,N_18983);
nand U19129 (N_19129,N_18880,N_18727);
nand U19130 (N_19130,N_18626,N_18501);
nor U19131 (N_19131,N_18695,N_18554);
or U19132 (N_19132,N_18861,N_18973);
nand U19133 (N_19133,N_18522,N_18976);
xnor U19134 (N_19134,N_18681,N_18640);
nor U19135 (N_19135,N_18692,N_18655);
or U19136 (N_19136,N_18870,N_18754);
nor U19137 (N_19137,N_18774,N_18606);
nor U19138 (N_19138,N_18642,N_18770);
or U19139 (N_19139,N_18834,N_18785);
nand U19140 (N_19140,N_18887,N_18752);
nand U19141 (N_19141,N_18508,N_18965);
or U19142 (N_19142,N_18935,N_18853);
nor U19143 (N_19143,N_18532,N_18603);
xnor U19144 (N_19144,N_18700,N_18764);
xor U19145 (N_19145,N_18540,N_18735);
xor U19146 (N_19146,N_18963,N_18577);
nor U19147 (N_19147,N_18761,N_18763);
and U19148 (N_19148,N_18724,N_18929);
and U19149 (N_19149,N_18794,N_18926);
and U19150 (N_19150,N_18790,N_18829);
xnor U19151 (N_19151,N_18750,N_18743);
or U19152 (N_19152,N_18579,N_18815);
nor U19153 (N_19153,N_18558,N_18971);
or U19154 (N_19154,N_18505,N_18991);
or U19155 (N_19155,N_18578,N_18575);
xor U19156 (N_19156,N_18719,N_18982);
nor U19157 (N_19157,N_18994,N_18544);
nand U19158 (N_19158,N_18530,N_18863);
and U19159 (N_19159,N_18661,N_18507);
xnor U19160 (N_19160,N_18840,N_18875);
nand U19161 (N_19161,N_18627,N_18920);
nor U19162 (N_19162,N_18841,N_18909);
nor U19163 (N_19163,N_18653,N_18660);
or U19164 (N_19164,N_18903,N_18723);
or U19165 (N_19165,N_18827,N_18742);
or U19166 (N_19166,N_18969,N_18745);
and U19167 (N_19167,N_18744,N_18988);
or U19168 (N_19168,N_18504,N_18620);
or U19169 (N_19169,N_18975,N_18587);
or U19170 (N_19170,N_18816,N_18832);
and U19171 (N_19171,N_18773,N_18788);
nand U19172 (N_19172,N_18518,N_18527);
and U19173 (N_19173,N_18873,N_18708);
and U19174 (N_19174,N_18552,N_18789);
and U19175 (N_19175,N_18675,N_18810);
xnor U19176 (N_19176,N_18741,N_18980);
and U19177 (N_19177,N_18925,N_18957);
nor U19178 (N_19178,N_18712,N_18685);
and U19179 (N_19179,N_18747,N_18931);
nand U19180 (N_19180,N_18550,N_18771);
and U19181 (N_19181,N_18818,N_18666);
nor U19182 (N_19182,N_18951,N_18918);
nor U19183 (N_19183,N_18892,N_18858);
nand U19184 (N_19184,N_18795,N_18567);
or U19185 (N_19185,N_18886,N_18792);
and U19186 (N_19186,N_18663,N_18514);
nand U19187 (N_19187,N_18865,N_18779);
nor U19188 (N_19188,N_18537,N_18520);
or U19189 (N_19189,N_18881,N_18930);
nand U19190 (N_19190,N_18573,N_18904);
and U19191 (N_19191,N_18799,N_18884);
xnor U19192 (N_19192,N_18506,N_18645);
or U19193 (N_19193,N_18798,N_18942);
xor U19194 (N_19194,N_18596,N_18542);
and U19195 (N_19195,N_18565,N_18569);
nand U19196 (N_19196,N_18566,N_18613);
nor U19197 (N_19197,N_18538,N_18968);
and U19198 (N_19198,N_18836,N_18632);
nor U19199 (N_19199,N_18954,N_18688);
nor U19200 (N_19200,N_18866,N_18684);
xor U19201 (N_19201,N_18813,N_18776);
nand U19202 (N_19202,N_18628,N_18778);
or U19203 (N_19203,N_18639,N_18623);
nand U19204 (N_19204,N_18883,N_18584);
or U19205 (N_19205,N_18948,N_18962);
nor U19206 (N_19206,N_18944,N_18933);
nand U19207 (N_19207,N_18531,N_18689);
nor U19208 (N_19208,N_18845,N_18697);
or U19209 (N_19209,N_18709,N_18722);
nor U19210 (N_19210,N_18882,N_18974);
nand U19211 (N_19211,N_18512,N_18720);
xnor U19212 (N_19212,N_18780,N_18616);
or U19213 (N_19213,N_18993,N_18772);
nor U19214 (N_19214,N_18857,N_18714);
nor U19215 (N_19215,N_18876,N_18914);
and U19216 (N_19216,N_18901,N_18753);
and U19217 (N_19217,N_18589,N_18659);
or U19218 (N_19218,N_18784,N_18959);
or U19219 (N_19219,N_18536,N_18545);
nand U19220 (N_19220,N_18760,N_18521);
or U19221 (N_19221,N_18737,N_18905);
or U19222 (N_19222,N_18561,N_18574);
and U19223 (N_19223,N_18729,N_18850);
and U19224 (N_19224,N_18871,N_18874);
nand U19225 (N_19225,N_18970,N_18599);
nor U19226 (N_19226,N_18916,N_18814);
xor U19227 (N_19227,N_18654,N_18837);
xnor U19228 (N_19228,N_18618,N_18641);
and U19229 (N_19229,N_18907,N_18593);
xnor U19230 (N_19230,N_18823,N_18822);
and U19231 (N_19231,N_18631,N_18796);
xor U19232 (N_19232,N_18662,N_18972);
nand U19233 (N_19233,N_18899,N_18984);
nor U19234 (N_19234,N_18629,N_18759);
nand U19235 (N_19235,N_18617,N_18819);
xnor U19236 (N_19236,N_18548,N_18523);
or U19237 (N_19237,N_18664,N_18896);
or U19238 (N_19238,N_18856,N_18890);
and U19239 (N_19239,N_18854,N_18878);
nor U19240 (N_19240,N_18553,N_18923);
xor U19241 (N_19241,N_18539,N_18513);
nand U19242 (N_19242,N_18838,N_18979);
nor U19243 (N_19243,N_18555,N_18820);
nand U19244 (N_19244,N_18755,N_18624);
xnor U19245 (N_19245,N_18877,N_18568);
and U19246 (N_19246,N_18952,N_18649);
or U19247 (N_19247,N_18867,N_18519);
xor U19248 (N_19248,N_18938,N_18888);
xor U19249 (N_19249,N_18806,N_18597);
xnor U19250 (N_19250,N_18644,N_18574);
nor U19251 (N_19251,N_18645,N_18734);
nor U19252 (N_19252,N_18973,N_18844);
and U19253 (N_19253,N_18798,N_18629);
nand U19254 (N_19254,N_18815,N_18973);
and U19255 (N_19255,N_18676,N_18532);
nand U19256 (N_19256,N_18790,N_18887);
and U19257 (N_19257,N_18612,N_18699);
nor U19258 (N_19258,N_18525,N_18927);
or U19259 (N_19259,N_18532,N_18951);
xnor U19260 (N_19260,N_18701,N_18933);
or U19261 (N_19261,N_18681,N_18674);
or U19262 (N_19262,N_18543,N_18770);
or U19263 (N_19263,N_18918,N_18698);
and U19264 (N_19264,N_18785,N_18694);
nor U19265 (N_19265,N_18568,N_18793);
nor U19266 (N_19266,N_18803,N_18851);
or U19267 (N_19267,N_18833,N_18805);
nand U19268 (N_19268,N_18742,N_18533);
xor U19269 (N_19269,N_18995,N_18913);
nor U19270 (N_19270,N_18848,N_18582);
nor U19271 (N_19271,N_18677,N_18564);
nand U19272 (N_19272,N_18915,N_18551);
nand U19273 (N_19273,N_18706,N_18829);
nor U19274 (N_19274,N_18574,N_18691);
and U19275 (N_19275,N_18856,N_18756);
nor U19276 (N_19276,N_18599,N_18507);
and U19277 (N_19277,N_18582,N_18852);
nand U19278 (N_19278,N_18916,N_18525);
and U19279 (N_19279,N_18640,N_18808);
nand U19280 (N_19280,N_18553,N_18956);
or U19281 (N_19281,N_18713,N_18727);
nor U19282 (N_19282,N_18904,N_18627);
and U19283 (N_19283,N_18682,N_18553);
and U19284 (N_19284,N_18528,N_18785);
nor U19285 (N_19285,N_18552,N_18966);
or U19286 (N_19286,N_18676,N_18810);
or U19287 (N_19287,N_18676,N_18817);
xnor U19288 (N_19288,N_18560,N_18791);
and U19289 (N_19289,N_18558,N_18529);
nor U19290 (N_19290,N_18866,N_18513);
nor U19291 (N_19291,N_18712,N_18704);
and U19292 (N_19292,N_18991,N_18652);
nor U19293 (N_19293,N_18967,N_18823);
nor U19294 (N_19294,N_18553,N_18835);
xor U19295 (N_19295,N_18775,N_18785);
nor U19296 (N_19296,N_18951,N_18644);
nand U19297 (N_19297,N_18727,N_18994);
and U19298 (N_19298,N_18804,N_18543);
nor U19299 (N_19299,N_18949,N_18814);
nand U19300 (N_19300,N_18991,N_18973);
and U19301 (N_19301,N_18960,N_18689);
nand U19302 (N_19302,N_18666,N_18706);
nand U19303 (N_19303,N_18644,N_18831);
or U19304 (N_19304,N_18862,N_18715);
xnor U19305 (N_19305,N_18885,N_18843);
or U19306 (N_19306,N_18786,N_18809);
nand U19307 (N_19307,N_18950,N_18845);
and U19308 (N_19308,N_18644,N_18782);
or U19309 (N_19309,N_18689,N_18774);
nand U19310 (N_19310,N_18736,N_18659);
xnor U19311 (N_19311,N_18804,N_18590);
nor U19312 (N_19312,N_18827,N_18668);
nand U19313 (N_19313,N_18969,N_18805);
or U19314 (N_19314,N_18936,N_18698);
nand U19315 (N_19315,N_18788,N_18570);
xnor U19316 (N_19316,N_18932,N_18962);
xnor U19317 (N_19317,N_18717,N_18528);
nor U19318 (N_19318,N_18805,N_18943);
xnor U19319 (N_19319,N_18994,N_18854);
nor U19320 (N_19320,N_18514,N_18729);
xnor U19321 (N_19321,N_18742,N_18576);
xnor U19322 (N_19322,N_18537,N_18623);
nor U19323 (N_19323,N_18725,N_18829);
nand U19324 (N_19324,N_18725,N_18817);
and U19325 (N_19325,N_18951,N_18513);
xnor U19326 (N_19326,N_18697,N_18973);
nor U19327 (N_19327,N_18550,N_18596);
nor U19328 (N_19328,N_18885,N_18657);
nand U19329 (N_19329,N_18746,N_18550);
and U19330 (N_19330,N_18615,N_18585);
xnor U19331 (N_19331,N_18758,N_18555);
nand U19332 (N_19332,N_18864,N_18629);
and U19333 (N_19333,N_18776,N_18814);
or U19334 (N_19334,N_18901,N_18627);
nor U19335 (N_19335,N_18556,N_18743);
nand U19336 (N_19336,N_18613,N_18667);
or U19337 (N_19337,N_18832,N_18728);
or U19338 (N_19338,N_18585,N_18894);
or U19339 (N_19339,N_18879,N_18668);
nor U19340 (N_19340,N_18988,N_18693);
and U19341 (N_19341,N_18965,N_18572);
or U19342 (N_19342,N_18513,N_18625);
nand U19343 (N_19343,N_18926,N_18779);
xor U19344 (N_19344,N_18715,N_18522);
or U19345 (N_19345,N_18616,N_18660);
and U19346 (N_19346,N_18775,N_18608);
or U19347 (N_19347,N_18727,N_18911);
or U19348 (N_19348,N_18537,N_18582);
and U19349 (N_19349,N_18632,N_18679);
nor U19350 (N_19350,N_18952,N_18980);
nor U19351 (N_19351,N_18731,N_18523);
and U19352 (N_19352,N_18674,N_18717);
xnor U19353 (N_19353,N_18761,N_18745);
or U19354 (N_19354,N_18605,N_18844);
and U19355 (N_19355,N_18679,N_18612);
xnor U19356 (N_19356,N_18540,N_18714);
nand U19357 (N_19357,N_18720,N_18697);
or U19358 (N_19358,N_18883,N_18916);
nand U19359 (N_19359,N_18906,N_18729);
or U19360 (N_19360,N_18584,N_18632);
or U19361 (N_19361,N_18785,N_18849);
nand U19362 (N_19362,N_18564,N_18789);
or U19363 (N_19363,N_18766,N_18851);
or U19364 (N_19364,N_18786,N_18839);
nand U19365 (N_19365,N_18641,N_18958);
and U19366 (N_19366,N_18794,N_18812);
nand U19367 (N_19367,N_18615,N_18686);
nand U19368 (N_19368,N_18614,N_18501);
or U19369 (N_19369,N_18760,N_18899);
xnor U19370 (N_19370,N_18625,N_18708);
and U19371 (N_19371,N_18611,N_18814);
and U19372 (N_19372,N_18919,N_18703);
or U19373 (N_19373,N_18619,N_18554);
or U19374 (N_19374,N_18629,N_18965);
and U19375 (N_19375,N_18871,N_18907);
and U19376 (N_19376,N_18780,N_18978);
or U19377 (N_19377,N_18742,N_18873);
xnor U19378 (N_19378,N_18677,N_18826);
nand U19379 (N_19379,N_18882,N_18963);
and U19380 (N_19380,N_18686,N_18554);
nand U19381 (N_19381,N_18711,N_18927);
and U19382 (N_19382,N_18992,N_18593);
xnor U19383 (N_19383,N_18547,N_18677);
and U19384 (N_19384,N_18634,N_18783);
and U19385 (N_19385,N_18678,N_18955);
xnor U19386 (N_19386,N_18635,N_18792);
xor U19387 (N_19387,N_18906,N_18650);
nand U19388 (N_19388,N_18666,N_18994);
nor U19389 (N_19389,N_18659,N_18770);
and U19390 (N_19390,N_18891,N_18944);
nand U19391 (N_19391,N_18679,N_18855);
or U19392 (N_19392,N_18802,N_18918);
or U19393 (N_19393,N_18890,N_18996);
or U19394 (N_19394,N_18791,N_18721);
nor U19395 (N_19395,N_18736,N_18781);
nand U19396 (N_19396,N_18777,N_18812);
nand U19397 (N_19397,N_18808,N_18573);
nand U19398 (N_19398,N_18754,N_18586);
or U19399 (N_19399,N_18809,N_18642);
xor U19400 (N_19400,N_18779,N_18907);
nor U19401 (N_19401,N_18613,N_18934);
nand U19402 (N_19402,N_18930,N_18816);
nor U19403 (N_19403,N_18908,N_18567);
or U19404 (N_19404,N_18717,N_18622);
xnor U19405 (N_19405,N_18877,N_18838);
nor U19406 (N_19406,N_18877,N_18812);
nand U19407 (N_19407,N_18598,N_18865);
or U19408 (N_19408,N_18717,N_18939);
and U19409 (N_19409,N_18596,N_18574);
and U19410 (N_19410,N_18965,N_18503);
nand U19411 (N_19411,N_18954,N_18769);
or U19412 (N_19412,N_18690,N_18649);
or U19413 (N_19413,N_18952,N_18509);
xor U19414 (N_19414,N_18575,N_18652);
or U19415 (N_19415,N_18883,N_18575);
or U19416 (N_19416,N_18557,N_18551);
nand U19417 (N_19417,N_18951,N_18779);
and U19418 (N_19418,N_18604,N_18805);
nor U19419 (N_19419,N_18871,N_18792);
and U19420 (N_19420,N_18741,N_18637);
or U19421 (N_19421,N_18694,N_18932);
nand U19422 (N_19422,N_18799,N_18901);
and U19423 (N_19423,N_18790,N_18651);
nor U19424 (N_19424,N_18556,N_18795);
nand U19425 (N_19425,N_18813,N_18664);
nor U19426 (N_19426,N_18629,N_18637);
and U19427 (N_19427,N_18813,N_18669);
nor U19428 (N_19428,N_18848,N_18777);
nand U19429 (N_19429,N_18805,N_18771);
xor U19430 (N_19430,N_18691,N_18787);
nor U19431 (N_19431,N_18575,N_18604);
or U19432 (N_19432,N_18720,N_18550);
nor U19433 (N_19433,N_18797,N_18885);
nor U19434 (N_19434,N_18848,N_18755);
and U19435 (N_19435,N_18540,N_18909);
or U19436 (N_19436,N_18989,N_18548);
xor U19437 (N_19437,N_18866,N_18724);
nor U19438 (N_19438,N_18914,N_18983);
and U19439 (N_19439,N_18838,N_18876);
or U19440 (N_19440,N_18728,N_18863);
xor U19441 (N_19441,N_18787,N_18979);
nor U19442 (N_19442,N_18880,N_18562);
xnor U19443 (N_19443,N_18785,N_18893);
or U19444 (N_19444,N_18903,N_18677);
nand U19445 (N_19445,N_18898,N_18875);
and U19446 (N_19446,N_18733,N_18601);
xnor U19447 (N_19447,N_18647,N_18639);
xor U19448 (N_19448,N_18771,N_18764);
nand U19449 (N_19449,N_18681,N_18882);
nor U19450 (N_19450,N_18509,N_18610);
or U19451 (N_19451,N_18755,N_18611);
or U19452 (N_19452,N_18698,N_18864);
xor U19453 (N_19453,N_18570,N_18737);
xnor U19454 (N_19454,N_18881,N_18740);
and U19455 (N_19455,N_18682,N_18837);
or U19456 (N_19456,N_18519,N_18684);
nor U19457 (N_19457,N_18963,N_18653);
or U19458 (N_19458,N_18543,N_18869);
nand U19459 (N_19459,N_18958,N_18805);
or U19460 (N_19460,N_18867,N_18979);
nand U19461 (N_19461,N_18637,N_18503);
xor U19462 (N_19462,N_18752,N_18960);
and U19463 (N_19463,N_18640,N_18688);
xor U19464 (N_19464,N_18972,N_18823);
or U19465 (N_19465,N_18696,N_18979);
xnor U19466 (N_19466,N_18997,N_18625);
nand U19467 (N_19467,N_18993,N_18748);
nor U19468 (N_19468,N_18952,N_18982);
and U19469 (N_19469,N_18956,N_18603);
or U19470 (N_19470,N_18869,N_18830);
and U19471 (N_19471,N_18772,N_18617);
or U19472 (N_19472,N_18568,N_18834);
nand U19473 (N_19473,N_18830,N_18981);
xnor U19474 (N_19474,N_18831,N_18787);
nand U19475 (N_19475,N_18692,N_18674);
xnor U19476 (N_19476,N_18687,N_18581);
nand U19477 (N_19477,N_18678,N_18529);
xor U19478 (N_19478,N_18978,N_18884);
nand U19479 (N_19479,N_18602,N_18736);
and U19480 (N_19480,N_18714,N_18818);
or U19481 (N_19481,N_18666,N_18529);
nand U19482 (N_19482,N_18875,N_18848);
or U19483 (N_19483,N_18787,N_18551);
nand U19484 (N_19484,N_18556,N_18957);
nor U19485 (N_19485,N_18764,N_18761);
nand U19486 (N_19486,N_18568,N_18598);
and U19487 (N_19487,N_18520,N_18710);
or U19488 (N_19488,N_18864,N_18937);
or U19489 (N_19489,N_18832,N_18747);
nor U19490 (N_19490,N_18794,N_18517);
and U19491 (N_19491,N_18608,N_18983);
nor U19492 (N_19492,N_18886,N_18965);
xnor U19493 (N_19493,N_18648,N_18793);
nor U19494 (N_19494,N_18685,N_18813);
nor U19495 (N_19495,N_18528,N_18851);
nor U19496 (N_19496,N_18820,N_18852);
xor U19497 (N_19497,N_18995,N_18896);
nand U19498 (N_19498,N_18775,N_18732);
nor U19499 (N_19499,N_18601,N_18655);
xor U19500 (N_19500,N_19333,N_19209);
or U19501 (N_19501,N_19498,N_19088);
or U19502 (N_19502,N_19008,N_19486);
nand U19503 (N_19503,N_19060,N_19378);
nand U19504 (N_19504,N_19258,N_19163);
or U19505 (N_19505,N_19104,N_19215);
and U19506 (N_19506,N_19266,N_19192);
xor U19507 (N_19507,N_19354,N_19186);
and U19508 (N_19508,N_19023,N_19082);
and U19509 (N_19509,N_19181,N_19496);
nor U19510 (N_19510,N_19445,N_19160);
or U19511 (N_19511,N_19447,N_19220);
nor U19512 (N_19512,N_19027,N_19430);
and U19513 (N_19513,N_19014,N_19078);
and U19514 (N_19514,N_19387,N_19157);
and U19515 (N_19515,N_19020,N_19340);
xnor U19516 (N_19516,N_19379,N_19061);
xor U19517 (N_19517,N_19065,N_19077);
nor U19518 (N_19518,N_19296,N_19221);
nor U19519 (N_19519,N_19318,N_19012);
nor U19520 (N_19520,N_19267,N_19190);
nand U19521 (N_19521,N_19396,N_19469);
nand U19522 (N_19522,N_19346,N_19177);
or U19523 (N_19523,N_19161,N_19327);
nand U19524 (N_19524,N_19265,N_19080);
and U19525 (N_19525,N_19293,N_19237);
nor U19526 (N_19526,N_19013,N_19238);
nand U19527 (N_19527,N_19417,N_19090);
xnor U19528 (N_19528,N_19336,N_19471);
nor U19529 (N_19529,N_19299,N_19337);
and U19530 (N_19530,N_19154,N_19274);
xnor U19531 (N_19531,N_19459,N_19328);
xnor U19532 (N_19532,N_19240,N_19303);
nor U19533 (N_19533,N_19149,N_19245);
and U19534 (N_19534,N_19047,N_19059);
or U19535 (N_19535,N_19432,N_19347);
and U19536 (N_19536,N_19076,N_19380);
and U19537 (N_19537,N_19195,N_19307);
and U19538 (N_19538,N_19207,N_19416);
nand U19539 (N_19539,N_19367,N_19120);
nor U19540 (N_19540,N_19365,N_19407);
xnor U19541 (N_19541,N_19398,N_19449);
nand U19542 (N_19542,N_19206,N_19199);
xor U19543 (N_19543,N_19180,N_19094);
nand U19544 (N_19544,N_19446,N_19388);
xor U19545 (N_19545,N_19089,N_19188);
or U19546 (N_19546,N_19465,N_19130);
or U19547 (N_19547,N_19382,N_19294);
nand U19548 (N_19548,N_19194,N_19034);
or U19549 (N_19549,N_19114,N_19464);
nor U19550 (N_19550,N_19042,N_19224);
nand U19551 (N_19551,N_19035,N_19068);
xor U19552 (N_19552,N_19440,N_19304);
xor U19553 (N_19553,N_19196,N_19275);
nor U19554 (N_19554,N_19234,N_19454);
nor U19555 (N_19555,N_19050,N_19159);
nor U19556 (N_19556,N_19331,N_19348);
nand U19557 (N_19557,N_19429,N_19492);
or U19558 (N_19558,N_19426,N_19376);
or U19559 (N_19559,N_19393,N_19273);
and U19560 (N_19560,N_19253,N_19063);
nor U19561 (N_19561,N_19046,N_19208);
nand U19562 (N_19562,N_19146,N_19119);
xnor U19563 (N_19563,N_19110,N_19145);
and U19564 (N_19564,N_19099,N_19103);
xnor U19565 (N_19565,N_19261,N_19249);
nand U19566 (N_19566,N_19451,N_19428);
nand U19567 (N_19567,N_19055,N_19461);
nand U19568 (N_19568,N_19412,N_19022);
nor U19569 (N_19569,N_19468,N_19197);
nand U19570 (N_19570,N_19127,N_19329);
and U19571 (N_19571,N_19437,N_19423);
nand U19572 (N_19572,N_19200,N_19455);
or U19573 (N_19573,N_19349,N_19287);
nand U19574 (N_19574,N_19394,N_19083);
xnor U19575 (N_19575,N_19124,N_19072);
xor U19576 (N_19576,N_19288,N_19374);
and U19577 (N_19577,N_19306,N_19000);
nor U19578 (N_19578,N_19286,N_19015);
or U19579 (N_19579,N_19064,N_19213);
or U19580 (N_19580,N_19176,N_19030);
nand U19581 (N_19581,N_19335,N_19268);
nor U19582 (N_19582,N_19118,N_19113);
and U19583 (N_19583,N_19325,N_19021);
or U19584 (N_19584,N_19017,N_19371);
or U19585 (N_19585,N_19372,N_19343);
and U19586 (N_19586,N_19143,N_19151);
and U19587 (N_19587,N_19310,N_19235);
xnor U19588 (N_19588,N_19230,N_19279);
xor U19589 (N_19589,N_19409,N_19352);
and U19590 (N_19590,N_19092,N_19025);
xor U19591 (N_19591,N_19375,N_19315);
or U19592 (N_19592,N_19173,N_19191);
nor U19593 (N_19593,N_19096,N_19436);
or U19594 (N_19594,N_19489,N_19026);
xnor U19595 (N_19595,N_19053,N_19048);
nand U19596 (N_19596,N_19260,N_19049);
nor U19597 (N_19597,N_19202,N_19134);
or U19598 (N_19598,N_19121,N_19247);
nand U19599 (N_19599,N_19164,N_19073);
nand U19600 (N_19600,N_19062,N_19472);
xor U19601 (N_19601,N_19165,N_19262);
and U19602 (N_19602,N_19324,N_19079);
nor U19603 (N_19603,N_19341,N_19448);
xor U19604 (N_19604,N_19236,N_19241);
nand U19605 (N_19605,N_19136,N_19497);
or U19606 (N_19606,N_19174,N_19462);
nor U19607 (N_19607,N_19431,N_19263);
or U19608 (N_19608,N_19384,N_19410);
or U19609 (N_19609,N_19087,N_19457);
and U19610 (N_19610,N_19313,N_19330);
xor U19611 (N_19611,N_19272,N_19389);
and U19612 (N_19612,N_19147,N_19250);
or U19613 (N_19613,N_19433,N_19137);
and U19614 (N_19614,N_19338,N_19128);
and U19615 (N_19615,N_19478,N_19251);
xnor U19616 (N_19616,N_19019,N_19093);
nor U19617 (N_19617,N_19298,N_19029);
or U19618 (N_19618,N_19277,N_19054);
or U19619 (N_19619,N_19182,N_19317);
xor U19620 (N_19620,N_19483,N_19123);
or U19621 (N_19621,N_19070,N_19474);
and U19622 (N_19622,N_19487,N_19381);
xnor U19623 (N_19623,N_19179,N_19283);
nand U19624 (N_19624,N_19232,N_19404);
nor U19625 (N_19625,N_19043,N_19485);
or U19626 (N_19626,N_19006,N_19133);
and U19627 (N_19627,N_19290,N_19399);
or U19628 (N_19628,N_19285,N_19052);
nor U19629 (N_19629,N_19219,N_19175);
nand U19630 (N_19630,N_19252,N_19243);
and U19631 (N_19631,N_19488,N_19040);
nand U19632 (N_19632,N_19439,N_19125);
and U19633 (N_19633,N_19218,N_19074);
and U19634 (N_19634,N_19189,N_19300);
nor U19635 (N_19635,N_19057,N_19084);
nand U19636 (N_19636,N_19494,N_19032);
nand U19637 (N_19637,N_19158,N_19463);
nor U19638 (N_19638,N_19010,N_19453);
nor U19639 (N_19639,N_19408,N_19400);
xor U19640 (N_19640,N_19355,N_19131);
nand U19641 (N_19641,N_19187,N_19255);
or U19642 (N_19642,N_19444,N_19039);
and U19643 (N_19643,N_19142,N_19001);
xor U19644 (N_19644,N_19126,N_19106);
xnor U19645 (N_19645,N_19311,N_19377);
nor U19646 (N_19646,N_19456,N_19309);
nand U19647 (N_19647,N_19415,N_19321);
nand U19648 (N_19648,N_19442,N_19112);
xnor U19649 (N_19649,N_19332,N_19427);
or U19650 (N_19650,N_19495,N_19071);
xor U19651 (N_19651,N_19210,N_19369);
and U19652 (N_19652,N_19357,N_19350);
and U19653 (N_19653,N_19401,N_19291);
xnor U19654 (N_19654,N_19222,N_19041);
and U19655 (N_19655,N_19490,N_19229);
nor U19656 (N_19656,N_19326,N_19153);
xor U19657 (N_19657,N_19166,N_19259);
xor U19658 (N_19658,N_19458,N_19156);
nand U19659 (N_19659,N_19140,N_19256);
xnor U19660 (N_19660,N_19476,N_19359);
nor U19661 (N_19661,N_19203,N_19270);
and U19662 (N_19662,N_19295,N_19011);
xnor U19663 (N_19663,N_19138,N_19257);
nor U19664 (N_19664,N_19075,N_19004);
and U19665 (N_19665,N_19002,N_19248);
xor U19666 (N_19666,N_19345,N_19193);
xor U19667 (N_19667,N_19183,N_19363);
xnor U19668 (N_19668,N_19271,N_19339);
or U19669 (N_19669,N_19480,N_19228);
nand U19670 (N_19670,N_19144,N_19434);
and U19671 (N_19671,N_19225,N_19217);
and U19672 (N_19672,N_19239,N_19028);
and U19673 (N_19673,N_19091,N_19314);
nand U19674 (N_19674,N_19212,N_19135);
xnor U19675 (N_19675,N_19491,N_19344);
or U19676 (N_19676,N_19122,N_19185);
nor U19677 (N_19677,N_19031,N_19223);
or U19678 (N_19678,N_19098,N_19081);
and U19679 (N_19679,N_19422,N_19282);
xor U19680 (N_19680,N_19264,N_19403);
nand U19681 (N_19681,N_19116,N_19095);
nand U19682 (N_19682,N_19292,N_19280);
or U19683 (N_19683,N_19305,N_19373);
or U19684 (N_19684,N_19425,N_19184);
and U19685 (N_19685,N_19391,N_19172);
or U19686 (N_19686,N_19467,N_19097);
nor U19687 (N_19687,N_19342,N_19045);
and U19688 (N_19688,N_19466,N_19281);
nand U19689 (N_19689,N_19141,N_19085);
nor U19690 (N_19690,N_19016,N_19242);
or U19691 (N_19691,N_19414,N_19470);
and U19692 (N_19692,N_19132,N_19364);
nor U19693 (N_19693,N_19056,N_19148);
nor U19694 (N_19694,N_19460,N_19441);
nand U19695 (N_19695,N_19413,N_19405);
and U19696 (N_19696,N_19007,N_19201);
nand U19697 (N_19697,N_19319,N_19421);
or U19698 (N_19698,N_19233,N_19171);
nand U19699 (N_19699,N_19051,N_19406);
nand U19700 (N_19700,N_19366,N_19108);
nand U19701 (N_19701,N_19320,N_19111);
xnor U19702 (N_19702,N_19360,N_19452);
nand U19703 (N_19703,N_19150,N_19227);
or U19704 (N_19704,N_19420,N_19368);
or U19705 (N_19705,N_19284,N_19302);
xnor U19706 (N_19706,N_19493,N_19443);
nor U19707 (N_19707,N_19038,N_19226);
and U19708 (N_19708,N_19139,N_19475);
xnor U19709 (N_19709,N_19205,N_19353);
xor U19710 (N_19710,N_19067,N_19435);
and U19711 (N_19711,N_19395,N_19036);
or U19712 (N_19712,N_19005,N_19392);
xnor U19713 (N_19713,N_19323,N_19385);
nor U19714 (N_19714,N_19482,N_19450);
and U19715 (N_19715,N_19278,N_19411);
nor U19716 (N_19716,N_19297,N_19162);
xnor U19717 (N_19717,N_19102,N_19086);
nor U19718 (N_19718,N_19316,N_19037);
and U19719 (N_19719,N_19152,N_19301);
nor U19720 (N_19720,N_19058,N_19244);
nand U19721 (N_19721,N_19419,N_19009);
nor U19722 (N_19722,N_19024,N_19362);
or U19723 (N_19723,N_19169,N_19479);
and U19724 (N_19724,N_19214,N_19390);
xor U19725 (N_19725,N_19308,N_19477);
and U19726 (N_19726,N_19198,N_19105);
xnor U19727 (N_19727,N_19178,N_19216);
xor U19728 (N_19728,N_19361,N_19115);
or U19729 (N_19729,N_19100,N_19356);
nor U19730 (N_19730,N_19117,N_19204);
xnor U19731 (N_19731,N_19018,N_19438);
nand U19732 (N_19732,N_19499,N_19170);
nand U19733 (N_19733,N_19269,N_19383);
nor U19734 (N_19734,N_19167,N_19322);
xnor U19735 (N_19735,N_19129,N_19370);
xor U19736 (N_19736,N_19334,N_19155);
and U19737 (N_19737,N_19033,N_19484);
xor U19738 (N_19738,N_19386,N_19003);
nor U19739 (N_19739,N_19418,N_19402);
nand U19740 (N_19740,N_19107,N_19397);
or U19741 (N_19741,N_19351,N_19109);
xor U19742 (N_19742,N_19231,N_19473);
or U19743 (N_19743,N_19289,N_19424);
nor U19744 (N_19744,N_19168,N_19211);
xnor U19745 (N_19745,N_19246,N_19358);
nor U19746 (N_19746,N_19481,N_19069);
or U19747 (N_19747,N_19312,N_19254);
xnor U19748 (N_19748,N_19101,N_19276);
or U19749 (N_19749,N_19066,N_19044);
nand U19750 (N_19750,N_19084,N_19174);
nor U19751 (N_19751,N_19182,N_19263);
and U19752 (N_19752,N_19354,N_19131);
xnor U19753 (N_19753,N_19136,N_19150);
xnor U19754 (N_19754,N_19452,N_19244);
nand U19755 (N_19755,N_19125,N_19003);
nor U19756 (N_19756,N_19370,N_19417);
xor U19757 (N_19757,N_19256,N_19288);
nor U19758 (N_19758,N_19407,N_19003);
nor U19759 (N_19759,N_19083,N_19472);
nand U19760 (N_19760,N_19360,N_19042);
or U19761 (N_19761,N_19356,N_19279);
nand U19762 (N_19762,N_19083,N_19246);
nand U19763 (N_19763,N_19163,N_19445);
nor U19764 (N_19764,N_19211,N_19434);
nand U19765 (N_19765,N_19306,N_19310);
and U19766 (N_19766,N_19485,N_19106);
and U19767 (N_19767,N_19115,N_19113);
nand U19768 (N_19768,N_19135,N_19238);
or U19769 (N_19769,N_19394,N_19392);
xnor U19770 (N_19770,N_19026,N_19386);
nand U19771 (N_19771,N_19364,N_19301);
nor U19772 (N_19772,N_19410,N_19474);
xnor U19773 (N_19773,N_19420,N_19424);
nor U19774 (N_19774,N_19498,N_19415);
and U19775 (N_19775,N_19395,N_19063);
xnor U19776 (N_19776,N_19115,N_19491);
xnor U19777 (N_19777,N_19034,N_19146);
and U19778 (N_19778,N_19233,N_19313);
or U19779 (N_19779,N_19079,N_19451);
nand U19780 (N_19780,N_19121,N_19125);
and U19781 (N_19781,N_19111,N_19023);
xor U19782 (N_19782,N_19073,N_19309);
xor U19783 (N_19783,N_19276,N_19024);
nor U19784 (N_19784,N_19247,N_19101);
and U19785 (N_19785,N_19271,N_19264);
or U19786 (N_19786,N_19187,N_19490);
nor U19787 (N_19787,N_19475,N_19083);
and U19788 (N_19788,N_19062,N_19112);
nand U19789 (N_19789,N_19305,N_19104);
nor U19790 (N_19790,N_19145,N_19463);
nor U19791 (N_19791,N_19374,N_19464);
and U19792 (N_19792,N_19375,N_19215);
or U19793 (N_19793,N_19419,N_19323);
nand U19794 (N_19794,N_19227,N_19239);
or U19795 (N_19795,N_19214,N_19059);
nand U19796 (N_19796,N_19277,N_19478);
nor U19797 (N_19797,N_19134,N_19311);
nand U19798 (N_19798,N_19111,N_19083);
xor U19799 (N_19799,N_19192,N_19228);
nor U19800 (N_19800,N_19387,N_19064);
nor U19801 (N_19801,N_19433,N_19045);
nand U19802 (N_19802,N_19466,N_19369);
and U19803 (N_19803,N_19316,N_19464);
and U19804 (N_19804,N_19052,N_19398);
and U19805 (N_19805,N_19499,N_19192);
and U19806 (N_19806,N_19236,N_19113);
nor U19807 (N_19807,N_19490,N_19008);
and U19808 (N_19808,N_19489,N_19041);
nor U19809 (N_19809,N_19293,N_19316);
nand U19810 (N_19810,N_19424,N_19416);
xor U19811 (N_19811,N_19340,N_19426);
or U19812 (N_19812,N_19042,N_19268);
and U19813 (N_19813,N_19424,N_19298);
or U19814 (N_19814,N_19015,N_19079);
nor U19815 (N_19815,N_19047,N_19378);
xnor U19816 (N_19816,N_19155,N_19049);
nand U19817 (N_19817,N_19153,N_19470);
nand U19818 (N_19818,N_19009,N_19003);
or U19819 (N_19819,N_19132,N_19328);
or U19820 (N_19820,N_19177,N_19383);
xnor U19821 (N_19821,N_19300,N_19261);
nand U19822 (N_19822,N_19029,N_19070);
nand U19823 (N_19823,N_19389,N_19231);
nor U19824 (N_19824,N_19476,N_19124);
and U19825 (N_19825,N_19162,N_19135);
nand U19826 (N_19826,N_19205,N_19037);
xor U19827 (N_19827,N_19069,N_19431);
nand U19828 (N_19828,N_19468,N_19320);
or U19829 (N_19829,N_19307,N_19406);
xor U19830 (N_19830,N_19450,N_19006);
and U19831 (N_19831,N_19272,N_19306);
nand U19832 (N_19832,N_19178,N_19041);
nand U19833 (N_19833,N_19400,N_19219);
nor U19834 (N_19834,N_19313,N_19002);
nor U19835 (N_19835,N_19458,N_19297);
xor U19836 (N_19836,N_19344,N_19343);
xnor U19837 (N_19837,N_19424,N_19136);
xnor U19838 (N_19838,N_19119,N_19300);
xnor U19839 (N_19839,N_19192,N_19429);
nand U19840 (N_19840,N_19195,N_19130);
xnor U19841 (N_19841,N_19279,N_19171);
nor U19842 (N_19842,N_19253,N_19076);
nand U19843 (N_19843,N_19152,N_19172);
or U19844 (N_19844,N_19164,N_19226);
and U19845 (N_19845,N_19443,N_19241);
nor U19846 (N_19846,N_19485,N_19392);
or U19847 (N_19847,N_19310,N_19082);
and U19848 (N_19848,N_19202,N_19061);
xor U19849 (N_19849,N_19170,N_19059);
xnor U19850 (N_19850,N_19068,N_19371);
nand U19851 (N_19851,N_19245,N_19338);
and U19852 (N_19852,N_19016,N_19039);
xnor U19853 (N_19853,N_19362,N_19231);
xnor U19854 (N_19854,N_19049,N_19111);
nor U19855 (N_19855,N_19005,N_19124);
and U19856 (N_19856,N_19479,N_19174);
nand U19857 (N_19857,N_19016,N_19175);
and U19858 (N_19858,N_19492,N_19037);
xnor U19859 (N_19859,N_19267,N_19098);
nand U19860 (N_19860,N_19238,N_19316);
nand U19861 (N_19861,N_19410,N_19476);
xnor U19862 (N_19862,N_19097,N_19385);
xor U19863 (N_19863,N_19347,N_19232);
nor U19864 (N_19864,N_19097,N_19417);
or U19865 (N_19865,N_19033,N_19436);
nand U19866 (N_19866,N_19102,N_19224);
and U19867 (N_19867,N_19015,N_19441);
and U19868 (N_19868,N_19295,N_19177);
xnor U19869 (N_19869,N_19402,N_19305);
nor U19870 (N_19870,N_19416,N_19323);
xnor U19871 (N_19871,N_19207,N_19459);
xnor U19872 (N_19872,N_19130,N_19000);
and U19873 (N_19873,N_19142,N_19014);
xor U19874 (N_19874,N_19042,N_19291);
and U19875 (N_19875,N_19192,N_19405);
nor U19876 (N_19876,N_19005,N_19349);
and U19877 (N_19877,N_19371,N_19406);
xnor U19878 (N_19878,N_19444,N_19053);
nand U19879 (N_19879,N_19442,N_19399);
xor U19880 (N_19880,N_19357,N_19168);
xnor U19881 (N_19881,N_19082,N_19039);
nor U19882 (N_19882,N_19446,N_19470);
nand U19883 (N_19883,N_19067,N_19413);
nor U19884 (N_19884,N_19499,N_19096);
xnor U19885 (N_19885,N_19466,N_19338);
nor U19886 (N_19886,N_19319,N_19378);
and U19887 (N_19887,N_19063,N_19025);
nor U19888 (N_19888,N_19012,N_19309);
nor U19889 (N_19889,N_19336,N_19145);
xor U19890 (N_19890,N_19394,N_19345);
nand U19891 (N_19891,N_19359,N_19005);
or U19892 (N_19892,N_19477,N_19094);
nand U19893 (N_19893,N_19318,N_19107);
xor U19894 (N_19894,N_19268,N_19208);
nand U19895 (N_19895,N_19234,N_19271);
xnor U19896 (N_19896,N_19491,N_19464);
nand U19897 (N_19897,N_19320,N_19497);
nor U19898 (N_19898,N_19472,N_19151);
and U19899 (N_19899,N_19460,N_19365);
and U19900 (N_19900,N_19286,N_19247);
nor U19901 (N_19901,N_19261,N_19272);
and U19902 (N_19902,N_19290,N_19064);
or U19903 (N_19903,N_19199,N_19040);
and U19904 (N_19904,N_19136,N_19300);
nor U19905 (N_19905,N_19226,N_19003);
and U19906 (N_19906,N_19177,N_19380);
nor U19907 (N_19907,N_19022,N_19195);
or U19908 (N_19908,N_19006,N_19073);
and U19909 (N_19909,N_19142,N_19199);
nor U19910 (N_19910,N_19018,N_19403);
nor U19911 (N_19911,N_19335,N_19049);
xor U19912 (N_19912,N_19363,N_19469);
and U19913 (N_19913,N_19135,N_19256);
nand U19914 (N_19914,N_19433,N_19110);
nand U19915 (N_19915,N_19187,N_19228);
or U19916 (N_19916,N_19104,N_19138);
nor U19917 (N_19917,N_19252,N_19420);
nand U19918 (N_19918,N_19477,N_19363);
xnor U19919 (N_19919,N_19312,N_19233);
xnor U19920 (N_19920,N_19386,N_19301);
xnor U19921 (N_19921,N_19214,N_19407);
nor U19922 (N_19922,N_19014,N_19053);
and U19923 (N_19923,N_19141,N_19252);
nand U19924 (N_19924,N_19050,N_19029);
nor U19925 (N_19925,N_19050,N_19222);
or U19926 (N_19926,N_19250,N_19308);
nor U19927 (N_19927,N_19037,N_19498);
xnor U19928 (N_19928,N_19057,N_19331);
nand U19929 (N_19929,N_19240,N_19076);
and U19930 (N_19930,N_19250,N_19048);
or U19931 (N_19931,N_19268,N_19061);
nand U19932 (N_19932,N_19359,N_19096);
or U19933 (N_19933,N_19422,N_19121);
and U19934 (N_19934,N_19314,N_19398);
and U19935 (N_19935,N_19331,N_19039);
nor U19936 (N_19936,N_19078,N_19148);
or U19937 (N_19937,N_19068,N_19145);
nand U19938 (N_19938,N_19302,N_19384);
and U19939 (N_19939,N_19169,N_19476);
nor U19940 (N_19940,N_19398,N_19390);
and U19941 (N_19941,N_19488,N_19135);
or U19942 (N_19942,N_19070,N_19166);
xnor U19943 (N_19943,N_19402,N_19194);
nor U19944 (N_19944,N_19287,N_19483);
and U19945 (N_19945,N_19074,N_19389);
nand U19946 (N_19946,N_19255,N_19082);
nor U19947 (N_19947,N_19384,N_19091);
nor U19948 (N_19948,N_19494,N_19218);
nand U19949 (N_19949,N_19201,N_19091);
nor U19950 (N_19950,N_19011,N_19374);
nor U19951 (N_19951,N_19048,N_19113);
nor U19952 (N_19952,N_19085,N_19186);
nor U19953 (N_19953,N_19223,N_19002);
nor U19954 (N_19954,N_19324,N_19007);
nand U19955 (N_19955,N_19198,N_19274);
xnor U19956 (N_19956,N_19022,N_19494);
xor U19957 (N_19957,N_19353,N_19153);
and U19958 (N_19958,N_19128,N_19004);
xor U19959 (N_19959,N_19243,N_19318);
nor U19960 (N_19960,N_19451,N_19016);
nand U19961 (N_19961,N_19322,N_19145);
nand U19962 (N_19962,N_19106,N_19281);
or U19963 (N_19963,N_19429,N_19040);
or U19964 (N_19964,N_19378,N_19430);
xnor U19965 (N_19965,N_19496,N_19086);
or U19966 (N_19966,N_19034,N_19033);
or U19967 (N_19967,N_19292,N_19258);
nor U19968 (N_19968,N_19218,N_19425);
xnor U19969 (N_19969,N_19257,N_19411);
nor U19970 (N_19970,N_19117,N_19148);
nand U19971 (N_19971,N_19213,N_19257);
or U19972 (N_19972,N_19134,N_19257);
nand U19973 (N_19973,N_19232,N_19045);
or U19974 (N_19974,N_19298,N_19456);
xor U19975 (N_19975,N_19422,N_19423);
or U19976 (N_19976,N_19271,N_19411);
nand U19977 (N_19977,N_19420,N_19498);
xor U19978 (N_19978,N_19247,N_19229);
xor U19979 (N_19979,N_19067,N_19359);
nand U19980 (N_19980,N_19322,N_19243);
nor U19981 (N_19981,N_19452,N_19293);
or U19982 (N_19982,N_19488,N_19409);
nand U19983 (N_19983,N_19270,N_19365);
and U19984 (N_19984,N_19244,N_19060);
or U19985 (N_19985,N_19420,N_19455);
nand U19986 (N_19986,N_19027,N_19169);
xnor U19987 (N_19987,N_19128,N_19035);
or U19988 (N_19988,N_19230,N_19044);
nand U19989 (N_19989,N_19358,N_19182);
nand U19990 (N_19990,N_19326,N_19278);
xnor U19991 (N_19991,N_19336,N_19436);
nor U19992 (N_19992,N_19382,N_19192);
xor U19993 (N_19993,N_19385,N_19246);
xor U19994 (N_19994,N_19306,N_19104);
nor U19995 (N_19995,N_19160,N_19405);
or U19996 (N_19996,N_19388,N_19387);
nor U19997 (N_19997,N_19249,N_19398);
and U19998 (N_19998,N_19120,N_19203);
and U19999 (N_19999,N_19308,N_19025);
xor U20000 (N_20000,N_19887,N_19603);
xor U20001 (N_20001,N_19827,N_19631);
xor U20002 (N_20002,N_19725,N_19539);
nor U20003 (N_20003,N_19519,N_19745);
xnor U20004 (N_20004,N_19811,N_19583);
nor U20005 (N_20005,N_19623,N_19975);
and U20006 (N_20006,N_19876,N_19521);
or U20007 (N_20007,N_19948,N_19943);
xor U20008 (N_20008,N_19585,N_19847);
and U20009 (N_20009,N_19930,N_19592);
nand U20010 (N_20010,N_19688,N_19541);
and U20011 (N_20011,N_19982,N_19710);
nand U20012 (N_20012,N_19879,N_19545);
or U20013 (N_20013,N_19909,N_19963);
xnor U20014 (N_20014,N_19905,N_19547);
and U20015 (N_20015,N_19752,N_19504);
or U20016 (N_20016,N_19892,N_19594);
nor U20017 (N_20017,N_19627,N_19872);
nor U20018 (N_20018,N_19924,N_19645);
or U20019 (N_20019,N_19788,N_19579);
or U20020 (N_20020,N_19736,N_19797);
nand U20021 (N_20021,N_19615,N_19964);
xnor U20022 (N_20022,N_19792,N_19514);
nor U20023 (N_20023,N_19553,N_19984);
xor U20024 (N_20024,N_19812,N_19618);
and U20025 (N_20025,N_19686,N_19965);
nor U20026 (N_20026,N_19888,N_19643);
nand U20027 (N_20027,N_19636,N_19757);
nand U20028 (N_20028,N_19974,N_19990);
and U20029 (N_20029,N_19536,N_19823);
or U20030 (N_20030,N_19906,N_19815);
nand U20031 (N_20031,N_19668,N_19743);
nand U20032 (N_20032,N_19840,N_19591);
nand U20033 (N_20033,N_19799,N_19561);
and U20034 (N_20034,N_19972,N_19667);
nor U20035 (N_20035,N_19529,N_19739);
or U20036 (N_20036,N_19582,N_19813);
or U20037 (N_20037,N_19853,N_19507);
xnor U20038 (N_20038,N_19637,N_19836);
and U20039 (N_20039,N_19932,N_19715);
xnor U20040 (N_20040,N_19896,N_19576);
nand U20041 (N_20041,N_19748,N_19895);
and U20042 (N_20042,N_19890,N_19998);
nor U20043 (N_20043,N_19968,N_19966);
xor U20044 (N_20044,N_19961,N_19852);
xor U20045 (N_20045,N_19737,N_19703);
nand U20046 (N_20046,N_19949,N_19992);
nand U20047 (N_20047,N_19729,N_19758);
nor U20048 (N_20048,N_19774,N_19789);
nor U20049 (N_20049,N_19918,N_19780);
and U20050 (N_20050,N_19628,N_19701);
nor U20051 (N_20051,N_19810,N_19566);
nor U20052 (N_20052,N_19653,N_19669);
nand U20053 (N_20053,N_19733,N_19947);
nor U20054 (N_20054,N_19958,N_19720);
and U20055 (N_20055,N_19925,N_19606);
and U20056 (N_20056,N_19995,N_19919);
nand U20057 (N_20057,N_19598,N_19915);
and U20058 (N_20058,N_19746,N_19633);
nor U20059 (N_20059,N_19663,N_19716);
or U20060 (N_20060,N_19898,N_19573);
and U20061 (N_20061,N_19534,N_19656);
nor U20062 (N_20062,N_19986,N_19540);
and U20063 (N_20063,N_19860,N_19983);
or U20064 (N_20064,N_19829,N_19988);
xor U20065 (N_20065,N_19787,N_19530);
nand U20066 (N_20066,N_19557,N_19554);
nand U20067 (N_20067,N_19546,N_19525);
nand U20068 (N_20068,N_19882,N_19850);
xnor U20069 (N_20069,N_19999,N_19770);
xor U20070 (N_20070,N_19693,N_19856);
nand U20071 (N_20071,N_19593,N_19723);
xnor U20072 (N_20072,N_19754,N_19558);
or U20073 (N_20073,N_19572,N_19819);
xnor U20074 (N_20074,N_19828,N_19768);
or U20075 (N_20075,N_19907,N_19946);
nor U20076 (N_20076,N_19611,N_19587);
or U20077 (N_20077,N_19773,N_19795);
xnor U20078 (N_20078,N_19864,N_19533);
xnor U20079 (N_20079,N_19936,N_19962);
and U20080 (N_20080,N_19769,N_19652);
nor U20081 (N_20081,N_19690,N_19979);
xnor U20082 (N_20082,N_19727,N_19845);
nand U20083 (N_20083,N_19762,N_19707);
and U20084 (N_20084,N_19711,N_19556);
and U20085 (N_20085,N_19666,N_19632);
and U20086 (N_20086,N_19674,N_19567);
xnor U20087 (N_20087,N_19781,N_19560);
xor U20088 (N_20088,N_19967,N_19692);
or U20089 (N_20089,N_19804,N_19953);
and U20090 (N_20090,N_19658,N_19698);
nand U20091 (N_20091,N_19764,N_19782);
and U20092 (N_20092,N_19894,N_19859);
and U20093 (N_20093,N_19806,N_19709);
nor U20094 (N_20094,N_19670,N_19543);
nor U20095 (N_20095,N_19803,N_19630);
xnor U20096 (N_20096,N_19518,N_19760);
nor U20097 (N_20097,N_19763,N_19708);
and U20098 (N_20098,N_19629,N_19809);
or U20099 (N_20099,N_19609,N_19904);
nor U20100 (N_20100,N_19874,N_19771);
and U20101 (N_20101,N_19677,N_19844);
or U20102 (N_20102,N_19862,N_19939);
nand U20103 (N_20103,N_19779,N_19549);
and U20104 (N_20104,N_19526,N_19916);
xnor U20105 (N_20105,N_19923,N_19646);
nand U20106 (N_20106,N_19577,N_19851);
nand U20107 (N_20107,N_19580,N_19959);
xor U20108 (N_20108,N_19713,N_19993);
and U20109 (N_20109,N_19978,N_19893);
nor U20110 (N_20110,N_19678,N_19537);
nand U20111 (N_20111,N_19857,N_19937);
xor U20112 (N_20112,N_19741,N_19548);
and U20113 (N_20113,N_19952,N_19971);
nor U20114 (N_20114,N_19734,N_19830);
nand U20115 (N_20115,N_19570,N_19866);
nor U20116 (N_20116,N_19920,N_19605);
or U20117 (N_20117,N_19502,N_19753);
and U20118 (N_20118,N_19613,N_19661);
nand U20119 (N_20119,N_19921,N_19889);
and U20120 (N_20120,N_19568,N_19601);
nor U20121 (N_20121,N_19801,N_19883);
nor U20122 (N_20122,N_19908,N_19622);
nor U20123 (N_20123,N_19755,N_19976);
or U20124 (N_20124,N_19735,N_19987);
or U20125 (N_20125,N_19927,N_19619);
and U20126 (N_20126,N_19843,N_19625);
nor U20127 (N_20127,N_19517,N_19912);
nand U20128 (N_20128,N_19522,N_19784);
nor U20129 (N_20129,N_19612,N_19863);
nand U20130 (N_20130,N_19825,N_19679);
nor U20131 (N_20131,N_19796,N_19704);
nor U20132 (N_20132,N_19858,N_19728);
nand U20133 (N_20133,N_19854,N_19726);
nand U20134 (N_20134,N_19868,N_19506);
and U20135 (N_20135,N_19621,N_19785);
or U20136 (N_20136,N_19794,N_19684);
nand U20137 (N_20137,N_19798,N_19662);
or U20138 (N_20138,N_19751,N_19740);
nor U20139 (N_20139,N_19849,N_19719);
xor U20140 (N_20140,N_19512,N_19772);
xor U20141 (N_20141,N_19875,N_19960);
nand U20142 (N_20142,N_19738,N_19586);
nand U20143 (N_20143,N_19861,N_19747);
nor U20144 (N_20144,N_19581,N_19886);
xnor U20145 (N_20145,N_19955,N_19702);
xor U20146 (N_20146,N_19913,N_19802);
nand U20147 (N_20147,N_19681,N_19538);
nor U20148 (N_20148,N_19865,N_19640);
xnor U20149 (N_20149,N_19841,N_19699);
nand U20150 (N_20150,N_19559,N_19516);
xnor U20151 (N_20151,N_19790,N_19996);
xor U20152 (N_20152,N_19911,N_19877);
or U20153 (N_20153,N_19867,N_19511);
nor U20154 (N_20154,N_19957,N_19721);
xor U20155 (N_20155,N_19808,N_19954);
nand U20156 (N_20156,N_19589,N_19838);
nor U20157 (N_20157,N_19687,N_19821);
or U20158 (N_20158,N_19878,N_19793);
and U20159 (N_20159,N_19917,N_19505);
nand U20160 (N_20160,N_19833,N_19956);
nand U20161 (N_20161,N_19578,N_19922);
and U20162 (N_20162,N_19989,N_19644);
or U20163 (N_20163,N_19528,N_19634);
and U20164 (N_20164,N_19544,N_19885);
xnor U20165 (N_20165,N_19846,N_19718);
nor U20166 (N_20166,N_19831,N_19834);
and U20167 (N_20167,N_19855,N_19820);
xnor U20168 (N_20168,N_19914,N_19783);
or U20169 (N_20169,N_19565,N_19926);
xor U20170 (N_20170,N_19664,N_19642);
or U20171 (N_20171,N_19655,N_19832);
nor U20172 (N_20172,N_19680,N_19897);
nand U20173 (N_20173,N_19510,N_19641);
nand U20174 (N_20174,N_19607,N_19750);
or U20175 (N_20175,N_19951,N_19575);
and U20176 (N_20176,N_19822,N_19997);
nand U20177 (N_20177,N_19508,N_19899);
and U20178 (N_20178,N_19839,N_19563);
xnor U20179 (N_20179,N_19730,N_19931);
xor U20180 (N_20180,N_19665,N_19654);
nand U20181 (N_20181,N_19776,N_19724);
nor U20182 (N_20182,N_19604,N_19614);
nor U20183 (N_20183,N_19891,N_19817);
nor U20184 (N_20184,N_19884,N_19527);
nor U20185 (N_20185,N_19991,N_19712);
xnor U20186 (N_20186,N_19824,N_19969);
nor U20187 (N_20187,N_19818,N_19842);
and U20188 (N_20188,N_19520,N_19938);
and U20189 (N_20189,N_19950,N_19685);
xor U20190 (N_20190,N_19610,N_19599);
nor U20191 (N_20191,N_19749,N_19695);
and U20192 (N_20192,N_19871,N_19706);
nor U20193 (N_20193,N_19555,N_19742);
nor U20194 (N_20194,N_19552,N_19985);
xor U20195 (N_20195,N_19523,N_19501);
or U20196 (N_20196,N_19659,N_19994);
nand U20197 (N_20197,N_19515,N_19869);
nor U20198 (N_20198,N_19673,N_19617);
nand U20199 (N_20199,N_19910,N_19676);
nand U20200 (N_20200,N_19531,N_19928);
and U20201 (N_20201,N_19691,N_19940);
or U20202 (N_20202,N_19602,N_19766);
nand U20203 (N_20203,N_19900,N_19778);
and U20204 (N_20204,N_19596,N_19945);
xor U20205 (N_20205,N_19714,N_19624);
nand U20206 (N_20206,N_19660,N_19597);
and U20207 (N_20207,N_19765,N_19675);
or U20208 (N_20208,N_19626,N_19584);
nand U20209 (N_20209,N_19934,N_19761);
and U20210 (N_20210,N_19616,N_19759);
xnor U20211 (N_20211,N_19980,N_19672);
or U20212 (N_20212,N_19647,N_19903);
nand U20213 (N_20213,N_19551,N_19837);
nor U20214 (N_20214,N_19542,N_19700);
nand U20215 (N_20215,N_19717,N_19807);
and U20216 (N_20216,N_19569,N_19638);
or U20217 (N_20217,N_19935,N_19564);
nor U20218 (N_20218,N_19977,N_19814);
and U20219 (N_20219,N_19513,N_19826);
nand U20220 (N_20220,N_19649,N_19791);
nor U20221 (N_20221,N_19775,N_19933);
or U20222 (N_20222,N_19744,N_19881);
or U20223 (N_20223,N_19696,N_19705);
nor U20224 (N_20224,N_19503,N_19944);
nor U20225 (N_20225,N_19595,N_19942);
or U20226 (N_20226,N_19620,N_19600);
nand U20227 (N_20227,N_19786,N_19722);
xnor U20228 (N_20228,N_19648,N_19650);
and U20229 (N_20229,N_19571,N_19509);
or U20230 (N_20230,N_19639,N_19635);
nand U20231 (N_20231,N_19732,N_19941);
and U20232 (N_20232,N_19671,N_19756);
xnor U20233 (N_20233,N_19848,N_19588);
nor U20234 (N_20234,N_19608,N_19535);
xnor U20235 (N_20235,N_19805,N_19880);
nor U20236 (N_20236,N_19777,N_19689);
nor U20237 (N_20237,N_19532,N_19901);
nor U20238 (N_20238,N_19800,N_19562);
or U20239 (N_20239,N_19590,N_19873);
nand U20240 (N_20240,N_19524,N_19970);
nor U20241 (N_20241,N_19870,N_19902);
nand U20242 (N_20242,N_19816,N_19835);
and U20243 (N_20243,N_19929,N_19657);
nand U20244 (N_20244,N_19574,N_19683);
or U20245 (N_20245,N_19550,N_19697);
or U20246 (N_20246,N_19651,N_19682);
or U20247 (N_20247,N_19500,N_19694);
xnor U20248 (N_20248,N_19767,N_19973);
or U20249 (N_20249,N_19731,N_19981);
or U20250 (N_20250,N_19880,N_19564);
nor U20251 (N_20251,N_19630,N_19987);
or U20252 (N_20252,N_19582,N_19764);
xnor U20253 (N_20253,N_19671,N_19708);
nor U20254 (N_20254,N_19832,N_19736);
xor U20255 (N_20255,N_19653,N_19784);
and U20256 (N_20256,N_19626,N_19517);
or U20257 (N_20257,N_19601,N_19821);
xnor U20258 (N_20258,N_19520,N_19535);
nand U20259 (N_20259,N_19981,N_19597);
or U20260 (N_20260,N_19711,N_19758);
or U20261 (N_20261,N_19978,N_19560);
nor U20262 (N_20262,N_19836,N_19871);
xor U20263 (N_20263,N_19838,N_19582);
or U20264 (N_20264,N_19711,N_19610);
xor U20265 (N_20265,N_19654,N_19875);
and U20266 (N_20266,N_19955,N_19744);
xnor U20267 (N_20267,N_19656,N_19626);
or U20268 (N_20268,N_19752,N_19963);
and U20269 (N_20269,N_19732,N_19813);
and U20270 (N_20270,N_19882,N_19703);
or U20271 (N_20271,N_19551,N_19515);
xor U20272 (N_20272,N_19856,N_19655);
xnor U20273 (N_20273,N_19586,N_19979);
xnor U20274 (N_20274,N_19786,N_19934);
or U20275 (N_20275,N_19731,N_19672);
nand U20276 (N_20276,N_19788,N_19624);
nor U20277 (N_20277,N_19876,N_19778);
nor U20278 (N_20278,N_19937,N_19659);
and U20279 (N_20279,N_19587,N_19800);
or U20280 (N_20280,N_19613,N_19625);
and U20281 (N_20281,N_19719,N_19507);
nor U20282 (N_20282,N_19812,N_19643);
and U20283 (N_20283,N_19599,N_19909);
and U20284 (N_20284,N_19630,N_19838);
xnor U20285 (N_20285,N_19905,N_19579);
or U20286 (N_20286,N_19874,N_19920);
or U20287 (N_20287,N_19541,N_19736);
nor U20288 (N_20288,N_19780,N_19910);
nor U20289 (N_20289,N_19989,N_19995);
nor U20290 (N_20290,N_19940,N_19563);
nor U20291 (N_20291,N_19802,N_19548);
nor U20292 (N_20292,N_19695,N_19882);
nor U20293 (N_20293,N_19607,N_19689);
xor U20294 (N_20294,N_19855,N_19726);
and U20295 (N_20295,N_19956,N_19918);
nand U20296 (N_20296,N_19983,N_19734);
nor U20297 (N_20297,N_19642,N_19849);
xor U20298 (N_20298,N_19825,N_19612);
nand U20299 (N_20299,N_19567,N_19576);
and U20300 (N_20300,N_19837,N_19623);
xor U20301 (N_20301,N_19813,N_19992);
or U20302 (N_20302,N_19701,N_19787);
nor U20303 (N_20303,N_19740,N_19536);
xnor U20304 (N_20304,N_19501,N_19668);
or U20305 (N_20305,N_19983,N_19541);
or U20306 (N_20306,N_19566,N_19957);
and U20307 (N_20307,N_19618,N_19729);
xor U20308 (N_20308,N_19687,N_19532);
xor U20309 (N_20309,N_19897,N_19777);
xor U20310 (N_20310,N_19585,N_19882);
and U20311 (N_20311,N_19533,N_19963);
and U20312 (N_20312,N_19894,N_19847);
and U20313 (N_20313,N_19510,N_19826);
nand U20314 (N_20314,N_19509,N_19782);
or U20315 (N_20315,N_19732,N_19979);
and U20316 (N_20316,N_19922,N_19668);
nor U20317 (N_20317,N_19922,N_19887);
and U20318 (N_20318,N_19596,N_19970);
or U20319 (N_20319,N_19532,N_19702);
and U20320 (N_20320,N_19819,N_19657);
and U20321 (N_20321,N_19671,N_19847);
nor U20322 (N_20322,N_19787,N_19981);
or U20323 (N_20323,N_19801,N_19627);
nor U20324 (N_20324,N_19564,N_19594);
nand U20325 (N_20325,N_19782,N_19579);
nand U20326 (N_20326,N_19973,N_19679);
and U20327 (N_20327,N_19782,N_19797);
nor U20328 (N_20328,N_19656,N_19639);
and U20329 (N_20329,N_19663,N_19938);
and U20330 (N_20330,N_19911,N_19850);
or U20331 (N_20331,N_19538,N_19778);
nor U20332 (N_20332,N_19506,N_19997);
nor U20333 (N_20333,N_19977,N_19861);
xnor U20334 (N_20334,N_19567,N_19597);
nor U20335 (N_20335,N_19763,N_19745);
xor U20336 (N_20336,N_19994,N_19786);
xnor U20337 (N_20337,N_19660,N_19756);
nor U20338 (N_20338,N_19869,N_19540);
xnor U20339 (N_20339,N_19603,N_19876);
xnor U20340 (N_20340,N_19775,N_19655);
and U20341 (N_20341,N_19970,N_19729);
and U20342 (N_20342,N_19907,N_19880);
nor U20343 (N_20343,N_19738,N_19508);
or U20344 (N_20344,N_19740,N_19693);
xor U20345 (N_20345,N_19814,N_19595);
and U20346 (N_20346,N_19914,N_19504);
xnor U20347 (N_20347,N_19578,N_19833);
or U20348 (N_20348,N_19637,N_19524);
and U20349 (N_20349,N_19991,N_19777);
and U20350 (N_20350,N_19886,N_19685);
or U20351 (N_20351,N_19769,N_19634);
xnor U20352 (N_20352,N_19501,N_19899);
or U20353 (N_20353,N_19739,N_19625);
and U20354 (N_20354,N_19671,N_19946);
xnor U20355 (N_20355,N_19872,N_19605);
xnor U20356 (N_20356,N_19654,N_19558);
xor U20357 (N_20357,N_19933,N_19733);
and U20358 (N_20358,N_19614,N_19858);
or U20359 (N_20359,N_19925,N_19614);
xnor U20360 (N_20360,N_19971,N_19522);
nor U20361 (N_20361,N_19716,N_19902);
nand U20362 (N_20362,N_19955,N_19501);
and U20363 (N_20363,N_19519,N_19780);
or U20364 (N_20364,N_19718,N_19769);
and U20365 (N_20365,N_19733,N_19786);
nor U20366 (N_20366,N_19649,N_19813);
xnor U20367 (N_20367,N_19917,N_19594);
nand U20368 (N_20368,N_19729,N_19791);
and U20369 (N_20369,N_19865,N_19953);
or U20370 (N_20370,N_19971,N_19511);
xor U20371 (N_20371,N_19812,N_19686);
or U20372 (N_20372,N_19534,N_19681);
xnor U20373 (N_20373,N_19903,N_19849);
nand U20374 (N_20374,N_19953,N_19583);
nor U20375 (N_20375,N_19789,N_19956);
nor U20376 (N_20376,N_19558,N_19537);
or U20377 (N_20377,N_19948,N_19767);
nand U20378 (N_20378,N_19616,N_19822);
nor U20379 (N_20379,N_19737,N_19671);
nor U20380 (N_20380,N_19545,N_19871);
xnor U20381 (N_20381,N_19716,N_19778);
and U20382 (N_20382,N_19783,N_19593);
xnor U20383 (N_20383,N_19967,N_19612);
nor U20384 (N_20384,N_19691,N_19728);
xnor U20385 (N_20385,N_19946,N_19605);
or U20386 (N_20386,N_19516,N_19954);
and U20387 (N_20387,N_19743,N_19918);
xor U20388 (N_20388,N_19704,N_19838);
nor U20389 (N_20389,N_19988,N_19886);
xnor U20390 (N_20390,N_19595,N_19517);
xor U20391 (N_20391,N_19568,N_19661);
nor U20392 (N_20392,N_19671,N_19571);
nor U20393 (N_20393,N_19941,N_19933);
and U20394 (N_20394,N_19590,N_19644);
nor U20395 (N_20395,N_19860,N_19639);
nand U20396 (N_20396,N_19562,N_19676);
or U20397 (N_20397,N_19903,N_19928);
xor U20398 (N_20398,N_19921,N_19871);
and U20399 (N_20399,N_19706,N_19882);
or U20400 (N_20400,N_19763,N_19721);
nand U20401 (N_20401,N_19691,N_19702);
and U20402 (N_20402,N_19899,N_19703);
nor U20403 (N_20403,N_19623,N_19538);
and U20404 (N_20404,N_19658,N_19768);
xnor U20405 (N_20405,N_19869,N_19702);
and U20406 (N_20406,N_19552,N_19995);
and U20407 (N_20407,N_19974,N_19629);
or U20408 (N_20408,N_19787,N_19690);
nand U20409 (N_20409,N_19906,N_19943);
nor U20410 (N_20410,N_19745,N_19525);
nor U20411 (N_20411,N_19913,N_19501);
nand U20412 (N_20412,N_19569,N_19549);
and U20413 (N_20413,N_19860,N_19978);
xor U20414 (N_20414,N_19876,N_19948);
and U20415 (N_20415,N_19706,N_19724);
nor U20416 (N_20416,N_19633,N_19950);
nor U20417 (N_20417,N_19954,N_19992);
nand U20418 (N_20418,N_19904,N_19559);
nand U20419 (N_20419,N_19615,N_19745);
or U20420 (N_20420,N_19927,N_19943);
and U20421 (N_20421,N_19801,N_19593);
xor U20422 (N_20422,N_19966,N_19690);
xor U20423 (N_20423,N_19947,N_19674);
nor U20424 (N_20424,N_19655,N_19850);
nor U20425 (N_20425,N_19901,N_19568);
nand U20426 (N_20426,N_19633,N_19936);
or U20427 (N_20427,N_19885,N_19549);
xor U20428 (N_20428,N_19733,N_19648);
and U20429 (N_20429,N_19736,N_19590);
or U20430 (N_20430,N_19581,N_19719);
nand U20431 (N_20431,N_19554,N_19804);
nor U20432 (N_20432,N_19839,N_19735);
or U20433 (N_20433,N_19759,N_19702);
nor U20434 (N_20434,N_19614,N_19511);
xor U20435 (N_20435,N_19800,N_19886);
nand U20436 (N_20436,N_19999,N_19979);
and U20437 (N_20437,N_19816,N_19694);
and U20438 (N_20438,N_19629,N_19702);
nor U20439 (N_20439,N_19787,N_19851);
and U20440 (N_20440,N_19946,N_19746);
and U20441 (N_20441,N_19917,N_19949);
nor U20442 (N_20442,N_19916,N_19913);
nand U20443 (N_20443,N_19966,N_19671);
or U20444 (N_20444,N_19866,N_19672);
xnor U20445 (N_20445,N_19576,N_19823);
nand U20446 (N_20446,N_19713,N_19542);
or U20447 (N_20447,N_19628,N_19934);
nand U20448 (N_20448,N_19752,N_19867);
nor U20449 (N_20449,N_19636,N_19669);
and U20450 (N_20450,N_19888,N_19684);
nor U20451 (N_20451,N_19719,N_19770);
nor U20452 (N_20452,N_19667,N_19643);
nand U20453 (N_20453,N_19685,N_19962);
or U20454 (N_20454,N_19692,N_19804);
nor U20455 (N_20455,N_19753,N_19905);
nand U20456 (N_20456,N_19793,N_19684);
and U20457 (N_20457,N_19578,N_19795);
nor U20458 (N_20458,N_19820,N_19763);
nand U20459 (N_20459,N_19594,N_19505);
or U20460 (N_20460,N_19760,N_19699);
xor U20461 (N_20461,N_19730,N_19585);
or U20462 (N_20462,N_19690,N_19534);
nand U20463 (N_20463,N_19557,N_19646);
nor U20464 (N_20464,N_19809,N_19899);
xor U20465 (N_20465,N_19561,N_19667);
or U20466 (N_20466,N_19541,N_19791);
or U20467 (N_20467,N_19825,N_19870);
and U20468 (N_20468,N_19512,N_19520);
or U20469 (N_20469,N_19759,N_19690);
or U20470 (N_20470,N_19601,N_19746);
xnor U20471 (N_20471,N_19508,N_19630);
xnor U20472 (N_20472,N_19743,N_19619);
xnor U20473 (N_20473,N_19626,N_19988);
or U20474 (N_20474,N_19612,N_19875);
or U20475 (N_20475,N_19611,N_19703);
nor U20476 (N_20476,N_19817,N_19580);
nand U20477 (N_20477,N_19872,N_19844);
xnor U20478 (N_20478,N_19583,N_19796);
and U20479 (N_20479,N_19932,N_19870);
and U20480 (N_20480,N_19824,N_19870);
xnor U20481 (N_20481,N_19641,N_19765);
xor U20482 (N_20482,N_19639,N_19894);
nand U20483 (N_20483,N_19727,N_19829);
or U20484 (N_20484,N_19766,N_19895);
nand U20485 (N_20485,N_19988,N_19765);
nor U20486 (N_20486,N_19701,N_19502);
or U20487 (N_20487,N_19870,N_19688);
nand U20488 (N_20488,N_19646,N_19958);
nand U20489 (N_20489,N_19677,N_19518);
nand U20490 (N_20490,N_19778,N_19806);
or U20491 (N_20491,N_19882,N_19522);
or U20492 (N_20492,N_19756,N_19787);
or U20493 (N_20493,N_19680,N_19788);
and U20494 (N_20494,N_19947,N_19665);
or U20495 (N_20495,N_19825,N_19919);
and U20496 (N_20496,N_19828,N_19899);
and U20497 (N_20497,N_19546,N_19531);
or U20498 (N_20498,N_19738,N_19534);
or U20499 (N_20499,N_19918,N_19975);
xor U20500 (N_20500,N_20167,N_20472);
nand U20501 (N_20501,N_20322,N_20391);
nand U20502 (N_20502,N_20325,N_20246);
or U20503 (N_20503,N_20331,N_20349);
nor U20504 (N_20504,N_20357,N_20196);
and U20505 (N_20505,N_20477,N_20224);
nor U20506 (N_20506,N_20358,N_20242);
nor U20507 (N_20507,N_20455,N_20418);
or U20508 (N_20508,N_20155,N_20465);
nand U20509 (N_20509,N_20421,N_20125);
nand U20510 (N_20510,N_20142,N_20473);
or U20511 (N_20511,N_20141,N_20347);
xor U20512 (N_20512,N_20380,N_20255);
xnor U20513 (N_20513,N_20081,N_20440);
and U20514 (N_20514,N_20361,N_20412);
nand U20515 (N_20515,N_20417,N_20199);
nand U20516 (N_20516,N_20450,N_20286);
or U20517 (N_20517,N_20041,N_20495);
and U20518 (N_20518,N_20116,N_20466);
nor U20519 (N_20519,N_20163,N_20177);
or U20520 (N_20520,N_20042,N_20399);
and U20521 (N_20521,N_20341,N_20036);
or U20522 (N_20522,N_20106,N_20335);
nand U20523 (N_20523,N_20102,N_20314);
or U20524 (N_20524,N_20205,N_20496);
or U20525 (N_20525,N_20033,N_20485);
and U20526 (N_20526,N_20103,N_20316);
nand U20527 (N_20527,N_20165,N_20187);
and U20528 (N_20528,N_20014,N_20434);
xor U20529 (N_20529,N_20161,N_20158);
nand U20530 (N_20530,N_20185,N_20258);
and U20531 (N_20531,N_20241,N_20173);
nor U20532 (N_20532,N_20071,N_20388);
nand U20533 (N_20533,N_20237,N_20323);
nor U20534 (N_20534,N_20490,N_20139);
and U20535 (N_20535,N_20453,N_20119);
xor U20536 (N_20536,N_20275,N_20423);
and U20537 (N_20537,N_20297,N_20160);
or U20538 (N_20538,N_20216,N_20193);
nand U20539 (N_20539,N_20111,N_20247);
and U20540 (N_20540,N_20148,N_20183);
and U20541 (N_20541,N_20032,N_20270);
xor U20542 (N_20542,N_20223,N_20303);
nor U20543 (N_20543,N_20488,N_20156);
nand U20544 (N_20544,N_20351,N_20336);
and U20545 (N_20545,N_20018,N_20365);
and U20546 (N_20546,N_20245,N_20019);
nand U20547 (N_20547,N_20024,N_20031);
nor U20548 (N_20548,N_20110,N_20203);
xor U20549 (N_20549,N_20372,N_20145);
or U20550 (N_20550,N_20382,N_20432);
nor U20551 (N_20551,N_20376,N_20213);
nor U20552 (N_20552,N_20211,N_20188);
xor U20553 (N_20553,N_20381,N_20257);
nand U20554 (N_20554,N_20301,N_20135);
xor U20555 (N_20555,N_20068,N_20210);
xnor U20556 (N_20556,N_20154,N_20166);
xor U20557 (N_20557,N_20047,N_20462);
or U20558 (N_20558,N_20209,N_20426);
nor U20559 (N_20559,N_20217,N_20368);
nand U20560 (N_20560,N_20099,N_20389);
or U20561 (N_20561,N_20186,N_20386);
and U20562 (N_20562,N_20494,N_20120);
xor U20563 (N_20563,N_20363,N_20044);
nand U20564 (N_20564,N_20435,N_20429);
nand U20565 (N_20565,N_20333,N_20304);
xor U20566 (N_20566,N_20202,N_20171);
nor U20567 (N_20567,N_20190,N_20457);
nand U20568 (N_20568,N_20401,N_20330);
xor U20569 (N_20569,N_20063,N_20064);
nand U20570 (N_20570,N_20084,N_20022);
nor U20571 (N_20571,N_20220,N_20164);
nand U20572 (N_20572,N_20482,N_20229);
nor U20573 (N_20573,N_20130,N_20150);
nand U20574 (N_20574,N_20373,N_20390);
and U20575 (N_20575,N_20274,N_20134);
nor U20576 (N_20576,N_20454,N_20006);
nand U20577 (N_20577,N_20384,N_20447);
nor U20578 (N_20578,N_20197,N_20452);
and U20579 (N_20579,N_20436,N_20350);
or U20580 (N_20580,N_20470,N_20419);
and U20581 (N_20581,N_20074,N_20248);
xnor U20582 (N_20582,N_20260,N_20083);
nor U20583 (N_20583,N_20309,N_20413);
and U20584 (N_20584,N_20035,N_20009);
nor U20585 (N_20585,N_20121,N_20317);
nor U20586 (N_20586,N_20463,N_20329);
nand U20587 (N_20587,N_20152,N_20222);
nand U20588 (N_20588,N_20289,N_20291);
nand U20589 (N_20589,N_20311,N_20468);
nand U20590 (N_20590,N_20027,N_20321);
nor U20591 (N_20591,N_20003,N_20402);
xor U20592 (N_20592,N_20214,N_20400);
nor U20593 (N_20593,N_20179,N_20225);
nor U20594 (N_20594,N_20305,N_20089);
and U20595 (N_20595,N_20433,N_20114);
nand U20596 (N_20596,N_20236,N_20232);
nor U20597 (N_20597,N_20374,N_20355);
xnor U20598 (N_20598,N_20095,N_20132);
and U20599 (N_20599,N_20420,N_20484);
nand U20600 (N_20600,N_20332,N_20175);
nand U20601 (N_20601,N_20097,N_20021);
and U20602 (N_20602,N_20065,N_20427);
nor U20603 (N_20603,N_20445,N_20342);
or U20604 (N_20604,N_20046,N_20327);
xnor U20605 (N_20605,N_20377,N_20218);
nor U20606 (N_20606,N_20406,N_20493);
or U20607 (N_20607,N_20446,N_20263);
and U20608 (N_20608,N_20127,N_20370);
xnor U20609 (N_20609,N_20375,N_20282);
xnor U20610 (N_20610,N_20069,N_20138);
or U20611 (N_20611,N_20499,N_20343);
nand U20612 (N_20612,N_20151,N_20198);
nor U20613 (N_20613,N_20292,N_20425);
nor U20614 (N_20614,N_20147,N_20481);
nor U20615 (N_20615,N_20475,N_20393);
nor U20616 (N_20616,N_20459,N_20379);
xnor U20617 (N_20617,N_20053,N_20040);
xnor U20618 (N_20618,N_20281,N_20029);
xnor U20619 (N_20619,N_20208,N_20367);
nand U20620 (N_20620,N_20408,N_20424);
or U20621 (N_20621,N_20228,N_20299);
or U20622 (N_20622,N_20461,N_20176);
nand U20623 (N_20623,N_20000,N_20077);
and U20624 (N_20624,N_20411,N_20431);
or U20625 (N_20625,N_20238,N_20123);
and U20626 (N_20626,N_20107,N_20091);
nand U20627 (N_20627,N_20430,N_20181);
and U20628 (N_20628,N_20078,N_20268);
xnor U20629 (N_20629,N_20359,N_20285);
nor U20630 (N_20630,N_20369,N_20170);
xnor U20631 (N_20631,N_20215,N_20479);
xnor U20632 (N_20632,N_20094,N_20293);
or U20633 (N_20633,N_20169,N_20178);
nor U20634 (N_20634,N_20030,N_20067);
and U20635 (N_20635,N_20449,N_20128);
nand U20636 (N_20636,N_20338,N_20366);
and U20637 (N_20637,N_20409,N_20007);
nor U20638 (N_20638,N_20101,N_20079);
and U20639 (N_20639,N_20448,N_20066);
or U20640 (N_20640,N_20256,N_20456);
and U20641 (N_20641,N_20356,N_20439);
nor U20642 (N_20642,N_20073,N_20273);
xor U20643 (N_20643,N_20278,N_20318);
nor U20644 (N_20644,N_20100,N_20109);
nand U20645 (N_20645,N_20276,N_20200);
or U20646 (N_20646,N_20059,N_20428);
xnor U20647 (N_20647,N_20157,N_20090);
and U20648 (N_20648,N_20354,N_20284);
nand U20649 (N_20649,N_20226,N_20131);
nand U20650 (N_20650,N_20034,N_20467);
or U20651 (N_20651,N_20234,N_20207);
or U20652 (N_20652,N_20249,N_20231);
nand U20653 (N_20653,N_20195,N_20028);
or U20654 (N_20654,N_20011,N_20016);
or U20655 (N_20655,N_20180,N_20124);
nand U20656 (N_20656,N_20113,N_20144);
nand U20657 (N_20657,N_20298,N_20204);
xnor U20658 (N_20658,N_20253,N_20339);
xnor U20659 (N_20659,N_20219,N_20153);
nand U20660 (N_20660,N_20271,N_20162);
nor U20661 (N_20661,N_20259,N_20061);
nand U20662 (N_20662,N_20397,N_20057);
or U20663 (N_20663,N_20392,N_20415);
or U20664 (N_20664,N_20239,N_20288);
nand U20665 (N_20665,N_20398,N_20407);
nor U20666 (N_20666,N_20015,N_20070);
and U20667 (N_20667,N_20050,N_20266);
or U20668 (N_20668,N_20302,N_20492);
and U20669 (N_20669,N_20476,N_20174);
nor U20670 (N_20670,N_20243,N_20300);
nand U20671 (N_20671,N_20117,N_20072);
xnor U20672 (N_20672,N_20280,N_20086);
xnor U20673 (N_20673,N_20104,N_20483);
or U20674 (N_20674,N_20037,N_20254);
xor U20675 (N_20675,N_20192,N_20096);
xor U20676 (N_20676,N_20159,N_20060);
nor U20677 (N_20677,N_20489,N_20277);
nand U20678 (N_20678,N_20039,N_20262);
nand U20679 (N_20679,N_20324,N_20189);
or U20680 (N_20680,N_20486,N_20251);
and U20681 (N_20681,N_20098,N_20056);
or U20682 (N_20682,N_20010,N_20058);
nand U20683 (N_20683,N_20227,N_20002);
xnor U20684 (N_20684,N_20026,N_20443);
xor U20685 (N_20685,N_20092,N_20126);
or U20686 (N_20686,N_20252,N_20264);
or U20687 (N_20687,N_20182,N_20149);
and U20688 (N_20688,N_20235,N_20352);
xor U20689 (N_20689,N_20410,N_20451);
nand U20690 (N_20690,N_20001,N_20055);
or U20691 (N_20691,N_20115,N_20387);
or U20692 (N_20692,N_20085,N_20320);
xor U20693 (N_20693,N_20308,N_20049);
and U20694 (N_20694,N_20296,N_20458);
and U20695 (N_20695,N_20396,N_20307);
or U20696 (N_20696,N_20005,N_20201);
and U20697 (N_20697,N_20414,N_20172);
and U20698 (N_20698,N_20017,N_20025);
and U20699 (N_20699,N_20334,N_20012);
or U20700 (N_20700,N_20080,N_20404);
xnor U20701 (N_20701,N_20441,N_20353);
xnor U20702 (N_20702,N_20474,N_20062);
nor U20703 (N_20703,N_20054,N_20498);
nor U20704 (N_20704,N_20184,N_20087);
or U20705 (N_20705,N_20075,N_20469);
nor U20706 (N_20706,N_20020,N_20140);
xnor U20707 (N_20707,N_20230,N_20405);
and U20708 (N_20708,N_20345,N_20313);
or U20709 (N_20709,N_20023,N_20269);
xnor U20710 (N_20710,N_20221,N_20112);
and U20711 (N_20711,N_20279,N_20118);
xnor U20712 (N_20712,N_20371,N_20051);
or U20713 (N_20713,N_20038,N_20326);
or U20714 (N_20714,N_20487,N_20444);
nor U20715 (N_20715,N_20129,N_20437);
and U20716 (N_20716,N_20261,N_20394);
nand U20717 (N_20717,N_20360,N_20383);
nor U20718 (N_20718,N_20122,N_20310);
nor U20719 (N_20719,N_20328,N_20480);
xnor U20720 (N_20720,N_20319,N_20287);
nor U20721 (N_20721,N_20076,N_20043);
xor U20722 (N_20722,N_20045,N_20306);
and U20723 (N_20723,N_20233,N_20416);
or U20724 (N_20724,N_20348,N_20133);
nand U20725 (N_20725,N_20422,N_20088);
or U20726 (N_20726,N_20471,N_20272);
or U20727 (N_20727,N_20194,N_20143);
xor U20728 (N_20728,N_20438,N_20008);
nand U20729 (N_20729,N_20395,N_20244);
nand U20730 (N_20730,N_20052,N_20497);
nor U20731 (N_20731,N_20478,N_20344);
and U20732 (N_20732,N_20267,N_20191);
nand U20733 (N_20733,N_20385,N_20337);
xnor U20734 (N_20734,N_20340,N_20048);
nor U20735 (N_20735,N_20082,N_20442);
nand U20736 (N_20736,N_20093,N_20346);
nand U20737 (N_20737,N_20362,N_20013);
and U20738 (N_20738,N_20378,N_20295);
xnor U20739 (N_20739,N_20364,N_20105);
or U20740 (N_20740,N_20206,N_20108);
nor U20741 (N_20741,N_20250,N_20137);
nand U20742 (N_20742,N_20315,N_20491);
nor U20743 (N_20743,N_20136,N_20240);
nand U20744 (N_20744,N_20460,N_20004);
and U20745 (N_20745,N_20265,N_20168);
nand U20746 (N_20746,N_20403,N_20294);
or U20747 (N_20747,N_20212,N_20146);
or U20748 (N_20748,N_20283,N_20290);
or U20749 (N_20749,N_20464,N_20312);
xnor U20750 (N_20750,N_20323,N_20204);
xor U20751 (N_20751,N_20435,N_20446);
xor U20752 (N_20752,N_20236,N_20380);
or U20753 (N_20753,N_20042,N_20334);
xor U20754 (N_20754,N_20154,N_20139);
and U20755 (N_20755,N_20084,N_20066);
or U20756 (N_20756,N_20155,N_20463);
nor U20757 (N_20757,N_20379,N_20195);
nand U20758 (N_20758,N_20419,N_20043);
nand U20759 (N_20759,N_20299,N_20473);
xor U20760 (N_20760,N_20239,N_20383);
or U20761 (N_20761,N_20498,N_20355);
and U20762 (N_20762,N_20309,N_20417);
xor U20763 (N_20763,N_20063,N_20495);
and U20764 (N_20764,N_20194,N_20302);
and U20765 (N_20765,N_20041,N_20224);
nor U20766 (N_20766,N_20481,N_20390);
nand U20767 (N_20767,N_20245,N_20116);
nor U20768 (N_20768,N_20389,N_20368);
nor U20769 (N_20769,N_20465,N_20098);
or U20770 (N_20770,N_20073,N_20095);
nor U20771 (N_20771,N_20177,N_20313);
or U20772 (N_20772,N_20173,N_20355);
and U20773 (N_20773,N_20089,N_20485);
xnor U20774 (N_20774,N_20337,N_20395);
xor U20775 (N_20775,N_20062,N_20063);
xor U20776 (N_20776,N_20181,N_20016);
nor U20777 (N_20777,N_20191,N_20366);
and U20778 (N_20778,N_20307,N_20197);
nor U20779 (N_20779,N_20341,N_20309);
xor U20780 (N_20780,N_20392,N_20282);
and U20781 (N_20781,N_20103,N_20327);
xnor U20782 (N_20782,N_20070,N_20289);
xor U20783 (N_20783,N_20499,N_20161);
nand U20784 (N_20784,N_20490,N_20298);
xor U20785 (N_20785,N_20436,N_20142);
and U20786 (N_20786,N_20448,N_20404);
or U20787 (N_20787,N_20423,N_20441);
nor U20788 (N_20788,N_20178,N_20266);
or U20789 (N_20789,N_20378,N_20248);
or U20790 (N_20790,N_20187,N_20421);
nor U20791 (N_20791,N_20454,N_20109);
nand U20792 (N_20792,N_20484,N_20204);
nor U20793 (N_20793,N_20331,N_20133);
or U20794 (N_20794,N_20166,N_20260);
nor U20795 (N_20795,N_20300,N_20327);
nor U20796 (N_20796,N_20089,N_20328);
xor U20797 (N_20797,N_20380,N_20102);
xor U20798 (N_20798,N_20358,N_20093);
nand U20799 (N_20799,N_20329,N_20452);
and U20800 (N_20800,N_20006,N_20189);
xnor U20801 (N_20801,N_20271,N_20275);
or U20802 (N_20802,N_20435,N_20091);
nand U20803 (N_20803,N_20071,N_20286);
and U20804 (N_20804,N_20431,N_20083);
and U20805 (N_20805,N_20103,N_20129);
xor U20806 (N_20806,N_20455,N_20460);
xnor U20807 (N_20807,N_20208,N_20406);
nor U20808 (N_20808,N_20463,N_20325);
and U20809 (N_20809,N_20264,N_20262);
nand U20810 (N_20810,N_20019,N_20443);
nand U20811 (N_20811,N_20286,N_20474);
nand U20812 (N_20812,N_20089,N_20422);
and U20813 (N_20813,N_20103,N_20367);
nand U20814 (N_20814,N_20188,N_20335);
nor U20815 (N_20815,N_20175,N_20226);
nand U20816 (N_20816,N_20306,N_20202);
nand U20817 (N_20817,N_20006,N_20310);
and U20818 (N_20818,N_20163,N_20214);
nor U20819 (N_20819,N_20299,N_20071);
xnor U20820 (N_20820,N_20155,N_20024);
and U20821 (N_20821,N_20461,N_20259);
nand U20822 (N_20822,N_20191,N_20450);
nand U20823 (N_20823,N_20077,N_20176);
xor U20824 (N_20824,N_20087,N_20141);
nor U20825 (N_20825,N_20051,N_20090);
nand U20826 (N_20826,N_20198,N_20142);
and U20827 (N_20827,N_20237,N_20332);
nor U20828 (N_20828,N_20383,N_20334);
or U20829 (N_20829,N_20147,N_20278);
xnor U20830 (N_20830,N_20407,N_20215);
or U20831 (N_20831,N_20156,N_20171);
nand U20832 (N_20832,N_20014,N_20101);
and U20833 (N_20833,N_20226,N_20220);
and U20834 (N_20834,N_20410,N_20204);
nor U20835 (N_20835,N_20046,N_20470);
and U20836 (N_20836,N_20232,N_20125);
and U20837 (N_20837,N_20389,N_20194);
and U20838 (N_20838,N_20245,N_20322);
and U20839 (N_20839,N_20484,N_20446);
or U20840 (N_20840,N_20020,N_20356);
xor U20841 (N_20841,N_20265,N_20455);
xor U20842 (N_20842,N_20443,N_20148);
nor U20843 (N_20843,N_20034,N_20290);
nor U20844 (N_20844,N_20410,N_20392);
xnor U20845 (N_20845,N_20283,N_20354);
and U20846 (N_20846,N_20070,N_20101);
nor U20847 (N_20847,N_20243,N_20066);
nor U20848 (N_20848,N_20390,N_20237);
nand U20849 (N_20849,N_20193,N_20321);
xnor U20850 (N_20850,N_20156,N_20260);
and U20851 (N_20851,N_20150,N_20387);
and U20852 (N_20852,N_20177,N_20144);
nand U20853 (N_20853,N_20286,N_20480);
xnor U20854 (N_20854,N_20250,N_20254);
or U20855 (N_20855,N_20491,N_20090);
nor U20856 (N_20856,N_20455,N_20087);
nor U20857 (N_20857,N_20456,N_20447);
and U20858 (N_20858,N_20482,N_20166);
xnor U20859 (N_20859,N_20284,N_20273);
nor U20860 (N_20860,N_20440,N_20067);
xor U20861 (N_20861,N_20301,N_20006);
and U20862 (N_20862,N_20428,N_20165);
and U20863 (N_20863,N_20480,N_20196);
and U20864 (N_20864,N_20103,N_20434);
nor U20865 (N_20865,N_20391,N_20151);
nor U20866 (N_20866,N_20292,N_20131);
nor U20867 (N_20867,N_20199,N_20385);
and U20868 (N_20868,N_20484,N_20180);
or U20869 (N_20869,N_20046,N_20349);
or U20870 (N_20870,N_20381,N_20261);
and U20871 (N_20871,N_20040,N_20311);
or U20872 (N_20872,N_20162,N_20469);
and U20873 (N_20873,N_20347,N_20000);
and U20874 (N_20874,N_20060,N_20065);
and U20875 (N_20875,N_20467,N_20405);
nor U20876 (N_20876,N_20283,N_20069);
nand U20877 (N_20877,N_20186,N_20214);
and U20878 (N_20878,N_20382,N_20336);
and U20879 (N_20879,N_20432,N_20470);
xor U20880 (N_20880,N_20051,N_20388);
and U20881 (N_20881,N_20131,N_20366);
nand U20882 (N_20882,N_20296,N_20234);
nand U20883 (N_20883,N_20293,N_20169);
xnor U20884 (N_20884,N_20373,N_20081);
nor U20885 (N_20885,N_20033,N_20124);
nor U20886 (N_20886,N_20404,N_20341);
nand U20887 (N_20887,N_20194,N_20321);
nor U20888 (N_20888,N_20190,N_20179);
or U20889 (N_20889,N_20348,N_20409);
and U20890 (N_20890,N_20080,N_20324);
xor U20891 (N_20891,N_20048,N_20381);
nor U20892 (N_20892,N_20450,N_20478);
or U20893 (N_20893,N_20232,N_20188);
and U20894 (N_20894,N_20151,N_20146);
nand U20895 (N_20895,N_20277,N_20476);
or U20896 (N_20896,N_20028,N_20323);
or U20897 (N_20897,N_20063,N_20467);
nor U20898 (N_20898,N_20473,N_20017);
nor U20899 (N_20899,N_20291,N_20321);
xnor U20900 (N_20900,N_20040,N_20498);
or U20901 (N_20901,N_20468,N_20404);
and U20902 (N_20902,N_20236,N_20132);
nor U20903 (N_20903,N_20133,N_20393);
nor U20904 (N_20904,N_20334,N_20198);
and U20905 (N_20905,N_20467,N_20340);
and U20906 (N_20906,N_20474,N_20480);
nor U20907 (N_20907,N_20388,N_20457);
nor U20908 (N_20908,N_20098,N_20438);
nand U20909 (N_20909,N_20438,N_20404);
or U20910 (N_20910,N_20440,N_20080);
xnor U20911 (N_20911,N_20471,N_20068);
and U20912 (N_20912,N_20494,N_20382);
xor U20913 (N_20913,N_20113,N_20019);
and U20914 (N_20914,N_20449,N_20291);
nand U20915 (N_20915,N_20268,N_20305);
nor U20916 (N_20916,N_20170,N_20396);
or U20917 (N_20917,N_20472,N_20234);
xor U20918 (N_20918,N_20451,N_20408);
or U20919 (N_20919,N_20323,N_20109);
or U20920 (N_20920,N_20313,N_20025);
nand U20921 (N_20921,N_20471,N_20134);
xnor U20922 (N_20922,N_20301,N_20473);
nand U20923 (N_20923,N_20285,N_20369);
xor U20924 (N_20924,N_20314,N_20244);
xnor U20925 (N_20925,N_20300,N_20480);
nor U20926 (N_20926,N_20147,N_20261);
and U20927 (N_20927,N_20074,N_20448);
or U20928 (N_20928,N_20450,N_20217);
or U20929 (N_20929,N_20022,N_20482);
xnor U20930 (N_20930,N_20476,N_20047);
nor U20931 (N_20931,N_20046,N_20405);
and U20932 (N_20932,N_20322,N_20494);
or U20933 (N_20933,N_20133,N_20111);
xnor U20934 (N_20934,N_20061,N_20237);
nor U20935 (N_20935,N_20350,N_20221);
xnor U20936 (N_20936,N_20194,N_20131);
nor U20937 (N_20937,N_20257,N_20279);
and U20938 (N_20938,N_20197,N_20375);
or U20939 (N_20939,N_20397,N_20022);
xor U20940 (N_20940,N_20014,N_20058);
and U20941 (N_20941,N_20067,N_20307);
and U20942 (N_20942,N_20453,N_20066);
or U20943 (N_20943,N_20141,N_20260);
or U20944 (N_20944,N_20443,N_20164);
and U20945 (N_20945,N_20092,N_20406);
nor U20946 (N_20946,N_20499,N_20409);
nor U20947 (N_20947,N_20170,N_20168);
xor U20948 (N_20948,N_20458,N_20242);
nand U20949 (N_20949,N_20342,N_20290);
or U20950 (N_20950,N_20454,N_20020);
nand U20951 (N_20951,N_20494,N_20499);
nand U20952 (N_20952,N_20256,N_20117);
nor U20953 (N_20953,N_20068,N_20103);
nor U20954 (N_20954,N_20213,N_20191);
nor U20955 (N_20955,N_20027,N_20042);
nand U20956 (N_20956,N_20471,N_20433);
and U20957 (N_20957,N_20283,N_20182);
xor U20958 (N_20958,N_20008,N_20219);
and U20959 (N_20959,N_20292,N_20448);
and U20960 (N_20960,N_20105,N_20201);
nand U20961 (N_20961,N_20223,N_20087);
and U20962 (N_20962,N_20282,N_20007);
xor U20963 (N_20963,N_20210,N_20251);
xnor U20964 (N_20964,N_20457,N_20427);
or U20965 (N_20965,N_20138,N_20008);
or U20966 (N_20966,N_20165,N_20167);
or U20967 (N_20967,N_20341,N_20221);
and U20968 (N_20968,N_20390,N_20158);
nand U20969 (N_20969,N_20010,N_20019);
nand U20970 (N_20970,N_20216,N_20011);
or U20971 (N_20971,N_20276,N_20003);
nor U20972 (N_20972,N_20462,N_20105);
nor U20973 (N_20973,N_20149,N_20469);
nand U20974 (N_20974,N_20337,N_20463);
or U20975 (N_20975,N_20402,N_20053);
nor U20976 (N_20976,N_20369,N_20112);
nor U20977 (N_20977,N_20171,N_20094);
and U20978 (N_20978,N_20261,N_20445);
nor U20979 (N_20979,N_20416,N_20180);
xnor U20980 (N_20980,N_20261,N_20181);
nor U20981 (N_20981,N_20246,N_20193);
or U20982 (N_20982,N_20237,N_20447);
or U20983 (N_20983,N_20331,N_20355);
or U20984 (N_20984,N_20344,N_20458);
nor U20985 (N_20985,N_20262,N_20428);
or U20986 (N_20986,N_20327,N_20264);
nor U20987 (N_20987,N_20029,N_20168);
nand U20988 (N_20988,N_20434,N_20347);
xor U20989 (N_20989,N_20034,N_20138);
xnor U20990 (N_20990,N_20189,N_20348);
xor U20991 (N_20991,N_20357,N_20150);
or U20992 (N_20992,N_20293,N_20101);
xnor U20993 (N_20993,N_20030,N_20040);
nor U20994 (N_20994,N_20010,N_20320);
xor U20995 (N_20995,N_20146,N_20465);
xor U20996 (N_20996,N_20178,N_20050);
nand U20997 (N_20997,N_20050,N_20194);
and U20998 (N_20998,N_20270,N_20240);
xor U20999 (N_20999,N_20116,N_20460);
xor U21000 (N_21000,N_20649,N_20647);
and U21001 (N_21001,N_20776,N_20597);
and U21002 (N_21002,N_20861,N_20876);
or U21003 (N_21003,N_20911,N_20917);
nand U21004 (N_21004,N_20753,N_20782);
xor U21005 (N_21005,N_20948,N_20606);
and U21006 (N_21006,N_20534,N_20660);
or U21007 (N_21007,N_20940,N_20848);
nand U21008 (N_21008,N_20902,N_20538);
and U21009 (N_21009,N_20786,N_20612);
nor U21010 (N_21010,N_20598,N_20920);
and U21011 (N_21011,N_20734,N_20966);
xor U21012 (N_21012,N_20559,N_20556);
and U21013 (N_21013,N_20619,N_20724);
and U21014 (N_21014,N_20973,N_20695);
xor U21015 (N_21015,N_20696,N_20582);
nand U21016 (N_21016,N_20555,N_20510);
nand U21017 (N_21017,N_20889,N_20603);
xnor U21018 (N_21018,N_20714,N_20543);
nor U21019 (N_21019,N_20587,N_20870);
xor U21020 (N_21020,N_20632,N_20502);
and U21021 (N_21021,N_20746,N_20872);
xor U21022 (N_21022,N_20518,N_20838);
nor U21023 (N_21023,N_20798,N_20620);
and U21024 (N_21024,N_20873,N_20816);
nor U21025 (N_21025,N_20721,N_20979);
nor U21026 (N_21026,N_20818,N_20697);
nand U21027 (N_21027,N_20933,N_20540);
nor U21028 (N_21028,N_20541,N_20953);
nor U21029 (N_21029,N_20659,N_20551);
nor U21030 (N_21030,N_20955,N_20690);
nand U21031 (N_21031,N_20744,N_20626);
or U21032 (N_21032,N_20529,N_20576);
nand U21033 (N_21033,N_20941,N_20677);
or U21034 (N_21034,N_20804,N_20894);
or U21035 (N_21035,N_20702,N_20657);
nor U21036 (N_21036,N_20977,N_20829);
nor U21037 (N_21037,N_20888,N_20665);
xor U21038 (N_21038,N_20871,N_20674);
or U21039 (N_21039,N_20661,N_20858);
nor U21040 (N_21040,N_20703,N_20519);
and U21041 (N_21041,N_20739,N_20561);
xor U21042 (N_21042,N_20994,N_20939);
xor U21043 (N_21043,N_20570,N_20947);
and U21044 (N_21044,N_20886,N_20935);
xnor U21045 (N_21045,N_20651,N_20578);
nand U21046 (N_21046,N_20532,N_20865);
nor U21047 (N_21047,N_20853,N_20964);
or U21048 (N_21048,N_20710,N_20918);
xor U21049 (N_21049,N_20595,N_20965);
xnor U21050 (N_21050,N_20704,N_20784);
or U21051 (N_21051,N_20500,N_20740);
or U21052 (N_21052,N_20914,N_20951);
nand U21053 (N_21053,N_20605,N_20859);
or U21054 (N_21054,N_20968,N_20508);
and U21055 (N_21055,N_20618,N_20879);
or U21056 (N_21056,N_20924,N_20905);
or U21057 (N_21057,N_20742,N_20516);
and U21058 (N_21058,N_20699,N_20539);
xnor U21059 (N_21059,N_20824,N_20509);
or U21060 (N_21060,N_20880,N_20883);
xor U21061 (N_21061,N_20971,N_20766);
nor U21062 (N_21062,N_20878,N_20503);
nand U21063 (N_21063,N_20814,N_20779);
or U21064 (N_21064,N_20681,N_20615);
nor U21065 (N_21065,N_20600,N_20755);
or U21066 (N_21066,N_20778,N_20921);
and U21067 (N_21067,N_20912,N_20738);
and U21068 (N_21068,N_20713,N_20528);
nand U21069 (N_21069,N_20590,N_20812);
nor U21070 (N_21070,N_20856,N_20756);
nor U21071 (N_21071,N_20643,N_20726);
nor U21072 (N_21072,N_20875,N_20944);
or U21073 (N_21073,N_20571,N_20849);
or U21074 (N_21074,N_20727,N_20560);
xor U21075 (N_21075,N_20926,N_20622);
nand U21076 (N_21076,N_20857,N_20707);
nand U21077 (N_21077,N_20970,N_20638);
xnor U21078 (N_21078,N_20767,N_20639);
nor U21079 (N_21079,N_20854,N_20799);
and U21080 (N_21080,N_20623,N_20942);
xnor U21081 (N_21081,N_20607,N_20828);
xor U21082 (N_21082,N_20811,N_20758);
xor U21083 (N_21083,N_20667,N_20736);
and U21084 (N_21084,N_20837,N_20513);
and U21085 (N_21085,N_20937,N_20771);
and U21086 (N_21086,N_20810,N_20783);
or U21087 (N_21087,N_20613,N_20760);
and U21088 (N_21088,N_20629,N_20662);
xnor U21089 (N_21089,N_20693,N_20995);
nor U21090 (N_21090,N_20827,N_20705);
or U21091 (N_21091,N_20986,N_20594);
xnor U21092 (N_21092,N_20850,N_20645);
or U21093 (N_21093,N_20761,N_20884);
and U21094 (N_21094,N_20604,N_20835);
nand U21095 (N_21095,N_20652,N_20521);
and U21096 (N_21096,N_20563,N_20715);
nand U21097 (N_21097,N_20580,N_20922);
nand U21098 (N_21098,N_20737,N_20535);
and U21099 (N_21099,N_20773,N_20903);
nand U21100 (N_21100,N_20795,N_20890);
nand U21101 (N_21101,N_20545,N_20842);
and U21102 (N_21102,N_20874,N_20774);
xor U21103 (N_21103,N_20867,N_20641);
nand U21104 (N_21104,N_20515,N_20822);
and U21105 (N_21105,N_20984,N_20862);
and U21106 (N_21106,N_20747,N_20931);
or U21107 (N_21107,N_20985,N_20684);
and U21108 (N_21108,N_20733,N_20785);
xnor U21109 (N_21109,N_20700,N_20927);
nor U21110 (N_21110,N_20946,N_20550);
nand U21111 (N_21111,N_20630,N_20511);
nand U21112 (N_21112,N_20514,N_20899);
xor U21113 (N_21113,N_20801,N_20718);
or U21114 (N_21114,N_20866,N_20698);
nand U21115 (N_21115,N_20544,N_20646);
xnor U21116 (N_21116,N_20794,N_20972);
xnor U21117 (N_21117,N_20754,N_20764);
or U21118 (N_21118,N_20789,N_20864);
or U21119 (N_21119,N_20572,N_20678);
and U21120 (N_21120,N_20893,N_20765);
nor U21121 (N_21121,N_20993,N_20844);
nor U21122 (N_21122,N_20950,N_20635);
and U21123 (N_21123,N_20839,N_20887);
nand U21124 (N_21124,N_20900,N_20983);
nand U21125 (N_21125,N_20685,N_20720);
xor U21126 (N_21126,N_20963,N_20763);
xor U21127 (N_21127,N_20666,N_20732);
nor U21128 (N_21128,N_20553,N_20974);
nor U21129 (N_21129,N_20599,N_20930);
nand U21130 (N_21130,N_20904,N_20611);
and U21131 (N_21131,N_20915,N_20554);
and U21132 (N_21132,N_20683,N_20520);
or U21133 (N_21133,N_20689,N_20506);
xnor U21134 (N_21134,N_20992,N_20601);
and U21135 (N_21135,N_20504,N_20589);
and U21136 (N_21136,N_20815,N_20910);
nor U21137 (N_21137,N_20680,N_20712);
xnor U21138 (N_21138,N_20562,N_20769);
nor U21139 (N_21139,N_20708,N_20833);
and U21140 (N_21140,N_20547,N_20564);
nand U21141 (N_21141,N_20748,N_20602);
nor U21142 (N_21142,N_20843,N_20577);
nor U21143 (N_21143,N_20803,N_20716);
xor U21144 (N_21144,N_20846,N_20749);
xor U21145 (N_21145,N_20975,N_20750);
xor U21146 (N_21146,N_20852,N_20725);
or U21147 (N_21147,N_20958,N_20791);
nand U21148 (N_21148,N_20847,N_20610);
nor U21149 (N_21149,N_20998,N_20806);
xnor U21150 (N_21150,N_20505,N_20717);
nor U21151 (N_21151,N_20722,N_20855);
nor U21152 (N_21152,N_20655,N_20731);
nand U21153 (N_21153,N_20989,N_20932);
and U21154 (N_21154,N_20885,N_20960);
nand U21155 (N_21155,N_20640,N_20530);
nand U21156 (N_21156,N_20945,N_20686);
nor U21157 (N_21157,N_20637,N_20907);
nand U21158 (N_21158,N_20593,N_20687);
xor U21159 (N_21159,N_20807,N_20790);
or U21160 (N_21160,N_20752,N_20787);
and U21161 (N_21161,N_20959,N_20581);
or U21162 (N_21162,N_20501,N_20648);
or U21163 (N_21163,N_20913,N_20719);
or U21164 (N_21164,N_20772,N_20802);
xnor U21165 (N_21165,N_20709,N_20568);
nand U21166 (N_21166,N_20831,N_20906);
and U21167 (N_21167,N_20898,N_20929);
xor U21168 (N_21168,N_20664,N_20527);
nor U21169 (N_21169,N_20569,N_20813);
nand U21170 (N_21170,N_20616,N_20588);
nor U21171 (N_21171,N_20533,N_20654);
xnor U21172 (N_21172,N_20546,N_20891);
nor U21173 (N_21173,N_20793,N_20536);
nand U21174 (N_21174,N_20729,N_20976);
or U21175 (N_21175,N_20625,N_20908);
and U21176 (N_21176,N_20676,N_20762);
or U21177 (N_21177,N_20585,N_20644);
nor U21178 (N_21178,N_20574,N_20507);
nor U21179 (N_21179,N_20658,N_20617);
nor U21180 (N_21180,N_20668,N_20670);
and U21181 (N_21181,N_20817,N_20841);
nor U21182 (N_21182,N_20781,N_20728);
nand U21183 (N_21183,N_20981,N_20621);
or U21184 (N_21184,N_20745,N_20987);
or U21185 (N_21185,N_20567,N_20624);
nand U21186 (N_21186,N_20759,N_20836);
or U21187 (N_21187,N_20851,N_20934);
nand U21188 (N_21188,N_20909,N_20628);
nor U21189 (N_21189,N_20775,N_20549);
nor U21190 (N_21190,N_20805,N_20751);
nand U21191 (N_21191,N_20996,N_20991);
or U21192 (N_21192,N_20840,N_20916);
nor U21193 (N_21193,N_20592,N_20691);
nor U21194 (N_21194,N_20777,N_20512);
and U21195 (N_21195,N_20672,N_20895);
nand U21196 (N_21196,N_20999,N_20634);
xnor U21197 (N_21197,N_20869,N_20980);
or U21198 (N_21198,N_20881,N_20819);
nand U21199 (N_21199,N_20573,N_20650);
xor U21200 (N_21200,N_20943,N_20642);
nor U21201 (N_21201,N_20990,N_20627);
and U21202 (N_21202,N_20961,N_20523);
xor U21203 (N_21203,N_20706,N_20919);
nor U21204 (N_21204,N_20524,N_20792);
and U21205 (N_21205,N_20692,N_20925);
nor U21206 (N_21206,N_20743,N_20809);
and U21207 (N_21207,N_20825,N_20531);
or U21208 (N_21208,N_20830,N_20552);
nand U21209 (N_21209,N_20936,N_20928);
nand U21210 (N_21210,N_20591,N_20688);
nor U21211 (N_21211,N_20673,N_20768);
and U21212 (N_21212,N_20845,N_20735);
nand U21213 (N_21213,N_20636,N_20957);
nand U21214 (N_21214,N_20633,N_20631);
nor U21215 (N_21215,N_20823,N_20796);
xnor U21216 (N_21216,N_20954,N_20537);
nor U21217 (N_21217,N_20757,N_20701);
and U21218 (N_21218,N_20797,N_20663);
xor U21219 (N_21219,N_20897,N_20679);
and U21220 (N_21220,N_20901,N_20860);
and U21221 (N_21221,N_20741,N_20614);
or U21222 (N_21222,N_20671,N_20653);
and U21223 (N_21223,N_20584,N_20923);
or U21224 (N_21224,N_20834,N_20949);
xnor U21225 (N_21225,N_20575,N_20788);
nand U21226 (N_21226,N_20882,N_20583);
xnor U21227 (N_21227,N_20956,N_20517);
xor U21228 (N_21228,N_20969,N_20682);
or U21229 (N_21229,N_20565,N_20694);
nand U21230 (N_21230,N_20770,N_20967);
nor U21231 (N_21231,N_20608,N_20808);
xor U21232 (N_21232,N_20982,N_20609);
xor U21233 (N_21233,N_20656,N_20821);
or U21234 (N_21234,N_20596,N_20542);
and U21235 (N_21235,N_20730,N_20892);
nor U21236 (N_21236,N_20820,N_20525);
xnor U21237 (N_21237,N_20579,N_20558);
nor U21238 (N_21238,N_20826,N_20832);
xnor U21239 (N_21239,N_20723,N_20877);
or U21240 (N_21240,N_20938,N_20675);
or U21241 (N_21241,N_20800,N_20952);
xnor U21242 (N_21242,N_20868,N_20548);
and U21243 (N_21243,N_20669,N_20526);
xor U21244 (N_21244,N_20896,N_20522);
or U21245 (N_21245,N_20978,N_20566);
nand U21246 (N_21246,N_20863,N_20557);
or U21247 (N_21247,N_20711,N_20988);
or U21248 (N_21248,N_20962,N_20586);
or U21249 (N_21249,N_20997,N_20780);
and U21250 (N_21250,N_20872,N_20793);
or U21251 (N_21251,N_20749,N_20625);
or U21252 (N_21252,N_20881,N_20713);
xor U21253 (N_21253,N_20618,N_20991);
and U21254 (N_21254,N_20965,N_20686);
nor U21255 (N_21255,N_20834,N_20642);
nand U21256 (N_21256,N_20571,N_20623);
xnor U21257 (N_21257,N_20913,N_20711);
xor U21258 (N_21258,N_20664,N_20758);
or U21259 (N_21259,N_20603,N_20564);
xnor U21260 (N_21260,N_20786,N_20788);
xor U21261 (N_21261,N_20612,N_20927);
and U21262 (N_21262,N_20926,N_20991);
xor U21263 (N_21263,N_20898,N_20502);
and U21264 (N_21264,N_20589,N_20834);
xor U21265 (N_21265,N_20777,N_20624);
nor U21266 (N_21266,N_20608,N_20888);
xor U21267 (N_21267,N_20890,N_20859);
and U21268 (N_21268,N_20916,N_20809);
xnor U21269 (N_21269,N_20763,N_20674);
nand U21270 (N_21270,N_20575,N_20526);
nand U21271 (N_21271,N_20925,N_20523);
nand U21272 (N_21272,N_20965,N_20946);
nand U21273 (N_21273,N_20857,N_20547);
nand U21274 (N_21274,N_20783,N_20925);
or U21275 (N_21275,N_20995,N_20762);
xor U21276 (N_21276,N_20521,N_20560);
nand U21277 (N_21277,N_20760,N_20783);
xnor U21278 (N_21278,N_20883,N_20554);
xor U21279 (N_21279,N_20536,N_20626);
nor U21280 (N_21280,N_20651,N_20998);
nand U21281 (N_21281,N_20501,N_20663);
nor U21282 (N_21282,N_20807,N_20582);
nor U21283 (N_21283,N_20854,N_20935);
nand U21284 (N_21284,N_20525,N_20962);
nand U21285 (N_21285,N_20669,N_20891);
nand U21286 (N_21286,N_20591,N_20515);
nand U21287 (N_21287,N_20988,N_20984);
or U21288 (N_21288,N_20807,N_20673);
or U21289 (N_21289,N_20938,N_20808);
xnor U21290 (N_21290,N_20780,N_20661);
nand U21291 (N_21291,N_20565,N_20880);
or U21292 (N_21292,N_20668,N_20525);
and U21293 (N_21293,N_20813,N_20723);
or U21294 (N_21294,N_20717,N_20610);
and U21295 (N_21295,N_20706,N_20694);
and U21296 (N_21296,N_20736,N_20823);
and U21297 (N_21297,N_20942,N_20721);
or U21298 (N_21298,N_20602,N_20607);
xor U21299 (N_21299,N_20931,N_20903);
nor U21300 (N_21300,N_20922,N_20603);
or U21301 (N_21301,N_20537,N_20603);
xor U21302 (N_21302,N_20542,N_20687);
or U21303 (N_21303,N_20669,N_20780);
nand U21304 (N_21304,N_20721,N_20972);
and U21305 (N_21305,N_20920,N_20565);
nor U21306 (N_21306,N_20894,N_20788);
nor U21307 (N_21307,N_20636,N_20585);
nand U21308 (N_21308,N_20861,N_20595);
xnor U21309 (N_21309,N_20521,N_20881);
or U21310 (N_21310,N_20662,N_20616);
or U21311 (N_21311,N_20999,N_20995);
nand U21312 (N_21312,N_20886,N_20748);
and U21313 (N_21313,N_20584,N_20929);
nor U21314 (N_21314,N_20960,N_20768);
nor U21315 (N_21315,N_20673,N_20850);
nand U21316 (N_21316,N_20815,N_20801);
xnor U21317 (N_21317,N_20594,N_20529);
or U21318 (N_21318,N_20539,N_20618);
or U21319 (N_21319,N_20940,N_20877);
nand U21320 (N_21320,N_20965,N_20885);
and U21321 (N_21321,N_20763,N_20917);
nor U21322 (N_21322,N_20555,N_20715);
nor U21323 (N_21323,N_20724,N_20855);
nor U21324 (N_21324,N_20629,N_20927);
or U21325 (N_21325,N_20657,N_20939);
and U21326 (N_21326,N_20582,N_20945);
or U21327 (N_21327,N_20683,N_20907);
xor U21328 (N_21328,N_20835,N_20983);
xnor U21329 (N_21329,N_20840,N_20838);
nand U21330 (N_21330,N_20879,N_20645);
nand U21331 (N_21331,N_20507,N_20669);
nor U21332 (N_21332,N_20747,N_20652);
xor U21333 (N_21333,N_20951,N_20805);
and U21334 (N_21334,N_20903,N_20916);
nand U21335 (N_21335,N_20868,N_20826);
xnor U21336 (N_21336,N_20905,N_20729);
nor U21337 (N_21337,N_20930,N_20581);
and U21338 (N_21338,N_20697,N_20601);
and U21339 (N_21339,N_20580,N_20965);
or U21340 (N_21340,N_20812,N_20611);
or U21341 (N_21341,N_20564,N_20500);
xor U21342 (N_21342,N_20905,N_20746);
or U21343 (N_21343,N_20700,N_20780);
xnor U21344 (N_21344,N_20762,N_20594);
and U21345 (N_21345,N_20573,N_20847);
nand U21346 (N_21346,N_20687,N_20686);
and U21347 (N_21347,N_20677,N_20649);
nor U21348 (N_21348,N_20694,N_20707);
and U21349 (N_21349,N_20830,N_20705);
xor U21350 (N_21350,N_20827,N_20548);
or U21351 (N_21351,N_20907,N_20730);
nand U21352 (N_21352,N_20861,N_20761);
or U21353 (N_21353,N_20841,N_20568);
and U21354 (N_21354,N_20796,N_20859);
or U21355 (N_21355,N_20888,N_20529);
and U21356 (N_21356,N_20627,N_20747);
or U21357 (N_21357,N_20864,N_20709);
or U21358 (N_21358,N_20644,N_20691);
xnor U21359 (N_21359,N_20681,N_20660);
nand U21360 (N_21360,N_20886,N_20781);
nor U21361 (N_21361,N_20703,N_20831);
or U21362 (N_21362,N_20684,N_20744);
and U21363 (N_21363,N_20700,N_20827);
xnor U21364 (N_21364,N_20696,N_20528);
and U21365 (N_21365,N_20533,N_20803);
nor U21366 (N_21366,N_20706,N_20723);
or U21367 (N_21367,N_20514,N_20932);
xnor U21368 (N_21368,N_20587,N_20998);
or U21369 (N_21369,N_20847,N_20930);
nand U21370 (N_21370,N_20752,N_20563);
or U21371 (N_21371,N_20782,N_20666);
nand U21372 (N_21372,N_20605,N_20981);
nor U21373 (N_21373,N_20911,N_20912);
nor U21374 (N_21374,N_20895,N_20693);
nand U21375 (N_21375,N_20718,N_20737);
nand U21376 (N_21376,N_20719,N_20995);
and U21377 (N_21377,N_20902,N_20978);
nor U21378 (N_21378,N_20654,N_20981);
nand U21379 (N_21379,N_20964,N_20771);
nor U21380 (N_21380,N_20896,N_20894);
nor U21381 (N_21381,N_20613,N_20852);
nand U21382 (N_21382,N_20626,N_20740);
nand U21383 (N_21383,N_20982,N_20561);
xor U21384 (N_21384,N_20597,N_20563);
and U21385 (N_21385,N_20933,N_20737);
nor U21386 (N_21386,N_20786,N_20883);
and U21387 (N_21387,N_20819,N_20958);
and U21388 (N_21388,N_20513,N_20609);
nand U21389 (N_21389,N_20571,N_20712);
xor U21390 (N_21390,N_20922,N_20517);
or U21391 (N_21391,N_20584,N_20808);
nor U21392 (N_21392,N_20638,N_20959);
xnor U21393 (N_21393,N_20894,N_20929);
and U21394 (N_21394,N_20714,N_20939);
and U21395 (N_21395,N_20518,N_20796);
and U21396 (N_21396,N_20571,N_20661);
nor U21397 (N_21397,N_20890,N_20964);
or U21398 (N_21398,N_20696,N_20703);
nor U21399 (N_21399,N_20804,N_20924);
or U21400 (N_21400,N_20988,N_20873);
nand U21401 (N_21401,N_20955,N_20987);
nor U21402 (N_21402,N_20972,N_20812);
and U21403 (N_21403,N_20957,N_20558);
xnor U21404 (N_21404,N_20862,N_20575);
nand U21405 (N_21405,N_20675,N_20763);
nand U21406 (N_21406,N_20946,N_20632);
and U21407 (N_21407,N_20581,N_20928);
xnor U21408 (N_21408,N_20633,N_20508);
nand U21409 (N_21409,N_20867,N_20794);
and U21410 (N_21410,N_20521,N_20868);
nand U21411 (N_21411,N_20747,N_20796);
nor U21412 (N_21412,N_20707,N_20941);
xnor U21413 (N_21413,N_20606,N_20588);
nand U21414 (N_21414,N_20696,N_20504);
xnor U21415 (N_21415,N_20521,N_20824);
nor U21416 (N_21416,N_20567,N_20643);
or U21417 (N_21417,N_20741,N_20580);
nand U21418 (N_21418,N_20713,N_20921);
nor U21419 (N_21419,N_20617,N_20900);
nand U21420 (N_21420,N_20787,N_20655);
and U21421 (N_21421,N_20992,N_20757);
xor U21422 (N_21422,N_20820,N_20843);
and U21423 (N_21423,N_20691,N_20805);
and U21424 (N_21424,N_20883,N_20753);
nor U21425 (N_21425,N_20773,N_20579);
nor U21426 (N_21426,N_20533,N_20766);
xor U21427 (N_21427,N_20619,N_20624);
xor U21428 (N_21428,N_20726,N_20571);
xor U21429 (N_21429,N_20763,N_20881);
nand U21430 (N_21430,N_20722,N_20847);
xnor U21431 (N_21431,N_20886,N_20594);
xor U21432 (N_21432,N_20664,N_20572);
xnor U21433 (N_21433,N_20759,N_20597);
xnor U21434 (N_21434,N_20866,N_20930);
nor U21435 (N_21435,N_20519,N_20972);
and U21436 (N_21436,N_20684,N_20537);
nand U21437 (N_21437,N_20517,N_20838);
or U21438 (N_21438,N_20862,N_20517);
and U21439 (N_21439,N_20544,N_20691);
and U21440 (N_21440,N_20504,N_20962);
nand U21441 (N_21441,N_20818,N_20764);
or U21442 (N_21442,N_20749,N_20693);
nor U21443 (N_21443,N_20861,N_20510);
and U21444 (N_21444,N_20677,N_20961);
nand U21445 (N_21445,N_20594,N_20591);
or U21446 (N_21446,N_20836,N_20937);
nand U21447 (N_21447,N_20848,N_20852);
xor U21448 (N_21448,N_20980,N_20688);
or U21449 (N_21449,N_20557,N_20906);
nand U21450 (N_21450,N_20868,N_20707);
nand U21451 (N_21451,N_20937,N_20899);
xnor U21452 (N_21452,N_20599,N_20947);
and U21453 (N_21453,N_20587,N_20669);
or U21454 (N_21454,N_20522,N_20777);
and U21455 (N_21455,N_20800,N_20508);
xnor U21456 (N_21456,N_20683,N_20549);
and U21457 (N_21457,N_20769,N_20582);
xor U21458 (N_21458,N_20604,N_20645);
nand U21459 (N_21459,N_20972,N_20952);
or U21460 (N_21460,N_20984,N_20829);
nand U21461 (N_21461,N_20986,N_20675);
xnor U21462 (N_21462,N_20697,N_20578);
nor U21463 (N_21463,N_20643,N_20547);
nor U21464 (N_21464,N_20638,N_20589);
nor U21465 (N_21465,N_20587,N_20560);
xor U21466 (N_21466,N_20930,N_20535);
xor U21467 (N_21467,N_20699,N_20781);
and U21468 (N_21468,N_20848,N_20571);
nor U21469 (N_21469,N_20698,N_20623);
and U21470 (N_21470,N_20582,N_20753);
nor U21471 (N_21471,N_20605,N_20621);
or U21472 (N_21472,N_20769,N_20888);
nand U21473 (N_21473,N_20777,N_20941);
or U21474 (N_21474,N_20809,N_20535);
nand U21475 (N_21475,N_20944,N_20767);
xor U21476 (N_21476,N_20583,N_20756);
nand U21477 (N_21477,N_20674,N_20583);
and U21478 (N_21478,N_20606,N_20918);
or U21479 (N_21479,N_20881,N_20983);
and U21480 (N_21480,N_20534,N_20579);
xnor U21481 (N_21481,N_20574,N_20793);
and U21482 (N_21482,N_20593,N_20536);
and U21483 (N_21483,N_20602,N_20571);
or U21484 (N_21484,N_20804,N_20806);
or U21485 (N_21485,N_20682,N_20535);
and U21486 (N_21486,N_20844,N_20642);
nand U21487 (N_21487,N_20628,N_20860);
nand U21488 (N_21488,N_20784,N_20988);
xnor U21489 (N_21489,N_20582,N_20642);
or U21490 (N_21490,N_20957,N_20502);
xor U21491 (N_21491,N_20985,N_20900);
or U21492 (N_21492,N_20642,N_20551);
or U21493 (N_21493,N_20865,N_20941);
xnor U21494 (N_21494,N_20959,N_20656);
and U21495 (N_21495,N_20958,N_20752);
nor U21496 (N_21496,N_20643,N_20757);
nand U21497 (N_21497,N_20931,N_20842);
and U21498 (N_21498,N_20707,N_20880);
or U21499 (N_21499,N_20996,N_20699);
xnor U21500 (N_21500,N_21087,N_21228);
nor U21501 (N_21501,N_21218,N_21090);
and U21502 (N_21502,N_21384,N_21476);
or U21503 (N_21503,N_21357,N_21440);
nand U21504 (N_21504,N_21400,N_21449);
and U21505 (N_21505,N_21026,N_21462);
or U21506 (N_21506,N_21349,N_21095);
nand U21507 (N_21507,N_21263,N_21229);
and U21508 (N_21508,N_21219,N_21362);
xor U21509 (N_21509,N_21408,N_21043);
xnor U21510 (N_21510,N_21497,N_21107);
nand U21511 (N_21511,N_21050,N_21429);
nor U21512 (N_21512,N_21425,N_21489);
and U21513 (N_21513,N_21366,N_21215);
or U21514 (N_21514,N_21057,N_21483);
xnor U21515 (N_21515,N_21315,N_21147);
and U21516 (N_21516,N_21352,N_21003);
xor U21517 (N_21517,N_21138,N_21376);
xnor U21518 (N_21518,N_21443,N_21073);
or U21519 (N_21519,N_21344,N_21072);
and U21520 (N_21520,N_21283,N_21000);
nand U21521 (N_21521,N_21133,N_21042);
nand U21522 (N_21522,N_21052,N_21044);
nor U21523 (N_21523,N_21447,N_21064);
and U21524 (N_21524,N_21242,N_21161);
or U21525 (N_21525,N_21297,N_21125);
nor U21526 (N_21526,N_21124,N_21296);
xnor U21527 (N_21527,N_21165,N_21067);
or U21528 (N_21528,N_21266,N_21036);
and U21529 (N_21529,N_21441,N_21198);
nand U21530 (N_21530,N_21424,N_21367);
and U21531 (N_21531,N_21231,N_21108);
nor U21532 (N_21532,N_21016,N_21484);
and U21533 (N_21533,N_21056,N_21136);
nand U21534 (N_21534,N_21088,N_21110);
nor U21535 (N_21535,N_21433,N_21285);
nand U21536 (N_21536,N_21460,N_21204);
nand U21537 (N_21537,N_21414,N_21022);
and U21538 (N_21538,N_21018,N_21160);
and U21539 (N_21539,N_21201,N_21478);
nor U21540 (N_21540,N_21093,N_21412);
nor U21541 (N_21541,N_21039,N_21370);
nor U21542 (N_21542,N_21146,N_21318);
xor U21543 (N_21543,N_21232,N_21361);
nand U21544 (N_21544,N_21438,N_21461);
or U21545 (N_21545,N_21375,N_21338);
and U21546 (N_21546,N_21121,N_21272);
nor U21547 (N_21547,N_21490,N_21031);
nand U21548 (N_21548,N_21084,N_21287);
or U21549 (N_21549,N_21221,N_21105);
and U21550 (N_21550,N_21294,N_21311);
or U21551 (N_21551,N_21451,N_21021);
xnor U21552 (N_21552,N_21098,N_21058);
or U21553 (N_21553,N_21137,N_21175);
nor U21554 (N_21554,N_21339,N_21158);
xor U21555 (N_21555,N_21379,N_21152);
or U21556 (N_21556,N_21112,N_21012);
xnor U21557 (N_21557,N_21120,N_21419);
nor U21558 (N_21558,N_21055,N_21340);
and U21559 (N_21559,N_21010,N_21322);
xor U21560 (N_21560,N_21282,N_21330);
or U21561 (N_21561,N_21019,N_21261);
and U21562 (N_21562,N_21227,N_21329);
nor U21563 (N_21563,N_21270,N_21247);
nand U21564 (N_21564,N_21312,N_21119);
xor U21565 (N_21565,N_21278,N_21196);
and U21566 (N_21566,N_21411,N_21343);
and U21567 (N_21567,N_21303,N_21331);
xnor U21568 (N_21568,N_21364,N_21033);
nand U21569 (N_21569,N_21396,N_21268);
or U21570 (N_21570,N_21001,N_21496);
nor U21571 (N_21571,N_21170,N_21390);
nand U21572 (N_21572,N_21235,N_21172);
and U21573 (N_21573,N_21060,N_21404);
xor U21574 (N_21574,N_21391,N_21399);
nor U21575 (N_21575,N_21274,N_21470);
nand U21576 (N_21576,N_21032,N_21437);
xnor U21577 (N_21577,N_21216,N_21454);
xnor U21578 (N_21578,N_21260,N_21254);
nand U21579 (N_21579,N_21080,N_21007);
nor U21580 (N_21580,N_21143,N_21486);
or U21581 (N_21581,N_21167,N_21387);
or U21582 (N_21582,N_21117,N_21104);
xor U21583 (N_21583,N_21086,N_21082);
nor U21584 (N_21584,N_21037,N_21038);
xor U21585 (N_21585,N_21488,N_21306);
or U21586 (N_21586,N_21498,N_21479);
xor U21587 (N_21587,N_21323,N_21499);
nand U21588 (N_21588,N_21079,N_21209);
nor U21589 (N_21589,N_21354,N_21074);
xnor U21590 (N_21590,N_21450,N_21275);
xnor U21591 (N_21591,N_21405,N_21421);
nand U21592 (N_21592,N_21439,N_21071);
nand U21593 (N_21593,N_21288,N_21290);
and U21594 (N_21594,N_21430,N_21264);
nand U21595 (N_21595,N_21053,N_21197);
xor U21596 (N_21596,N_21465,N_21402);
nor U21597 (N_21597,N_21314,N_21081);
nor U21598 (N_21598,N_21116,N_21214);
or U21599 (N_21599,N_21241,N_21193);
nor U21600 (N_21600,N_21213,N_21051);
nor U21601 (N_21601,N_21345,N_21406);
nand U21602 (N_21602,N_21027,N_21365);
nor U21603 (N_21603,N_21395,N_21111);
xnor U21604 (N_21604,N_21328,N_21253);
nand U21605 (N_21605,N_21385,N_21207);
nand U21606 (N_21606,N_21481,N_21122);
nand U21607 (N_21607,N_21463,N_21244);
and U21608 (N_21608,N_21100,N_21099);
nand U21609 (N_21609,N_21407,N_21166);
nand U21610 (N_21610,N_21374,N_21468);
nand U21611 (N_21611,N_21130,N_21359);
nand U21612 (N_21612,N_21135,N_21334);
nor U21613 (N_21613,N_21327,N_21205);
xnor U21614 (N_21614,N_21149,N_21348);
nand U21615 (N_21615,N_21163,N_21380);
xor U21616 (N_21616,N_21350,N_21113);
nand U21617 (N_21617,N_21427,N_21459);
and U21618 (N_21618,N_21011,N_21300);
nand U21619 (N_21619,N_21310,N_21179);
and U21620 (N_21620,N_21432,N_21302);
xnor U21621 (N_21621,N_21077,N_21417);
and U21622 (N_21622,N_21154,N_21356);
nand U21623 (N_21623,N_21203,N_21118);
xor U21624 (N_21624,N_21233,N_21292);
or U21625 (N_21625,N_21258,N_21250);
nor U21626 (N_21626,N_21492,N_21169);
nor U21627 (N_21627,N_21014,N_21182);
nor U21628 (N_21628,N_21145,N_21256);
and U21629 (N_21629,N_21369,N_21015);
xnor U21630 (N_21630,N_21393,N_21249);
nor U21631 (N_21631,N_21164,N_21075);
and U21632 (N_21632,N_21128,N_21455);
nand U21633 (N_21633,N_21185,N_21083);
xor U21634 (N_21634,N_21139,N_21148);
or U21635 (N_21635,N_21293,N_21126);
and U21636 (N_21636,N_21286,N_21453);
or U21637 (N_21637,N_21337,N_21076);
or U21638 (N_21638,N_21245,N_21190);
or U21639 (N_21639,N_21177,N_21341);
nand U21640 (N_21640,N_21251,N_21467);
or U21641 (N_21641,N_21317,N_21386);
and U21642 (N_21642,N_21176,N_21401);
and U21643 (N_21643,N_21109,N_21360);
and U21644 (N_21644,N_21381,N_21267);
nand U21645 (N_21645,N_21096,N_21153);
nor U21646 (N_21646,N_21280,N_21325);
or U21647 (N_21647,N_21040,N_21308);
nor U21648 (N_21648,N_21195,N_21223);
xnor U21649 (N_21649,N_21189,N_21141);
or U21650 (N_21650,N_21269,N_21444);
nor U21651 (N_21651,N_21240,N_21392);
and U21652 (N_21652,N_21123,N_21442);
and U21653 (N_21653,N_21236,N_21114);
nor U21654 (N_21654,N_21183,N_21262);
nor U21655 (N_21655,N_21048,N_21304);
and U21656 (N_21656,N_21485,N_21150);
and U21657 (N_21657,N_21333,N_21224);
nand U21658 (N_21658,N_21212,N_21452);
xnor U21659 (N_21659,N_21023,N_21324);
xor U21660 (N_21660,N_21326,N_21184);
nor U21661 (N_21661,N_21248,N_21456);
nand U21662 (N_21662,N_21134,N_21094);
xnor U21663 (N_21663,N_21276,N_21029);
nand U21664 (N_21664,N_21307,N_21188);
nor U21665 (N_21665,N_21085,N_21234);
nor U21666 (N_21666,N_21243,N_21445);
nor U21667 (N_21667,N_21277,N_21477);
xor U21668 (N_21668,N_21140,N_21045);
or U21669 (N_21669,N_21132,N_21473);
and U21670 (N_21670,N_21281,N_21469);
or U21671 (N_21671,N_21291,N_21259);
nand U21672 (N_21672,N_21373,N_21217);
xnor U21673 (N_21673,N_21426,N_21383);
and U21674 (N_21674,N_21159,N_21103);
or U21675 (N_21675,N_21363,N_21091);
xor U21676 (N_21676,N_21413,N_21482);
nand U21677 (N_21677,N_21377,N_21202);
or U21678 (N_21678,N_21418,N_21013);
nor U21679 (N_21679,N_21035,N_21252);
nor U21680 (N_21680,N_21480,N_21131);
and U21681 (N_21681,N_21005,N_21355);
xnor U21682 (N_21682,N_21063,N_21220);
nor U21683 (N_21683,N_21089,N_21435);
or U21684 (N_21684,N_21065,N_21279);
nand U21685 (N_21685,N_21208,N_21475);
or U21686 (N_21686,N_21006,N_21127);
or U21687 (N_21687,N_21487,N_21046);
xor U21688 (N_21688,N_21106,N_21457);
nor U21689 (N_21689,N_21246,N_21171);
or U21690 (N_21690,N_21494,N_21129);
nor U21691 (N_21691,N_21298,N_21347);
xor U21692 (N_21692,N_21472,N_21305);
or U21693 (N_21693,N_21034,N_21358);
and U21694 (N_21694,N_21410,N_21180);
and U21695 (N_21695,N_21313,N_21320);
nand U21696 (N_21696,N_21336,N_21230);
nand U21697 (N_21697,N_21194,N_21211);
and U21698 (N_21698,N_21493,N_21028);
nand U21699 (N_21699,N_21192,N_21257);
nand U21700 (N_21700,N_21353,N_21009);
nand U21701 (N_21701,N_21295,N_21319);
or U21702 (N_21702,N_21423,N_21436);
xor U21703 (N_21703,N_21059,N_21225);
or U21704 (N_21704,N_21054,N_21416);
and U21705 (N_21705,N_21210,N_21066);
xor U21706 (N_21706,N_21174,N_21335);
or U21707 (N_21707,N_21226,N_21237);
nand U21708 (N_21708,N_21162,N_21273);
or U21709 (N_21709,N_21102,N_21142);
or U21710 (N_21710,N_21378,N_21020);
nand U21711 (N_21711,N_21068,N_21398);
nand U21712 (N_21712,N_21346,N_21316);
xnor U21713 (N_21713,N_21388,N_21284);
and U21714 (N_21714,N_21025,N_21342);
nor U21715 (N_21715,N_21368,N_21178);
xnor U21716 (N_21716,N_21200,N_21092);
nand U21717 (N_21717,N_21403,N_21474);
or U21718 (N_21718,N_21041,N_21069);
nand U21719 (N_21719,N_21062,N_21255);
and U21720 (N_21720,N_21206,N_21309);
xor U21721 (N_21721,N_21332,N_21002);
or U21722 (N_21722,N_21097,N_21471);
nand U21723 (N_21723,N_21351,N_21199);
or U21724 (N_21724,N_21061,N_21415);
or U21725 (N_21725,N_21030,N_21156);
and U21726 (N_21726,N_21144,N_21428);
xor U21727 (N_21727,N_21017,N_21466);
or U21728 (N_21728,N_21409,N_21289);
nor U21729 (N_21729,N_21301,N_21397);
or U21730 (N_21730,N_21420,N_21491);
nand U21731 (N_21731,N_21495,N_21181);
or U21732 (N_21732,N_21299,N_21394);
nor U21733 (N_21733,N_21191,N_21448);
xnor U21734 (N_21734,N_21431,N_21238);
xnor U21735 (N_21735,N_21168,N_21371);
xnor U21736 (N_21736,N_21446,N_21047);
nand U21737 (N_21737,N_21422,N_21372);
or U21738 (N_21738,N_21186,N_21239);
and U21739 (N_21739,N_21271,N_21173);
xnor U21740 (N_21740,N_21004,N_21382);
xor U21741 (N_21741,N_21049,N_21265);
nor U21742 (N_21742,N_21115,N_21321);
xor U21743 (N_21743,N_21464,N_21458);
and U21744 (N_21744,N_21024,N_21151);
and U21745 (N_21745,N_21101,N_21389);
xor U21746 (N_21746,N_21434,N_21157);
xnor U21747 (N_21747,N_21222,N_21070);
nand U21748 (N_21748,N_21187,N_21008);
nor U21749 (N_21749,N_21155,N_21078);
or U21750 (N_21750,N_21139,N_21363);
or U21751 (N_21751,N_21125,N_21128);
or U21752 (N_21752,N_21131,N_21317);
or U21753 (N_21753,N_21451,N_21004);
or U21754 (N_21754,N_21135,N_21450);
or U21755 (N_21755,N_21205,N_21041);
and U21756 (N_21756,N_21489,N_21276);
nor U21757 (N_21757,N_21413,N_21103);
xnor U21758 (N_21758,N_21328,N_21121);
xor U21759 (N_21759,N_21019,N_21122);
xor U21760 (N_21760,N_21372,N_21218);
and U21761 (N_21761,N_21151,N_21075);
xnor U21762 (N_21762,N_21334,N_21327);
and U21763 (N_21763,N_21324,N_21092);
xnor U21764 (N_21764,N_21493,N_21333);
nor U21765 (N_21765,N_21336,N_21489);
nor U21766 (N_21766,N_21350,N_21294);
nor U21767 (N_21767,N_21093,N_21176);
nand U21768 (N_21768,N_21198,N_21289);
or U21769 (N_21769,N_21407,N_21014);
and U21770 (N_21770,N_21031,N_21332);
and U21771 (N_21771,N_21014,N_21024);
xor U21772 (N_21772,N_21430,N_21285);
nand U21773 (N_21773,N_21438,N_21479);
nand U21774 (N_21774,N_21117,N_21100);
nor U21775 (N_21775,N_21169,N_21079);
nor U21776 (N_21776,N_21426,N_21121);
nand U21777 (N_21777,N_21143,N_21234);
or U21778 (N_21778,N_21390,N_21067);
xnor U21779 (N_21779,N_21161,N_21128);
nand U21780 (N_21780,N_21042,N_21003);
nor U21781 (N_21781,N_21431,N_21206);
or U21782 (N_21782,N_21073,N_21294);
and U21783 (N_21783,N_21376,N_21482);
or U21784 (N_21784,N_21376,N_21092);
xnor U21785 (N_21785,N_21120,N_21203);
or U21786 (N_21786,N_21233,N_21311);
nand U21787 (N_21787,N_21404,N_21039);
or U21788 (N_21788,N_21456,N_21271);
xnor U21789 (N_21789,N_21381,N_21216);
nand U21790 (N_21790,N_21229,N_21251);
nor U21791 (N_21791,N_21132,N_21462);
nor U21792 (N_21792,N_21313,N_21204);
nor U21793 (N_21793,N_21219,N_21483);
or U21794 (N_21794,N_21438,N_21227);
xnor U21795 (N_21795,N_21272,N_21387);
or U21796 (N_21796,N_21339,N_21122);
nor U21797 (N_21797,N_21244,N_21493);
nand U21798 (N_21798,N_21071,N_21219);
or U21799 (N_21799,N_21320,N_21054);
or U21800 (N_21800,N_21282,N_21312);
nor U21801 (N_21801,N_21384,N_21075);
xor U21802 (N_21802,N_21193,N_21082);
nor U21803 (N_21803,N_21037,N_21125);
or U21804 (N_21804,N_21474,N_21460);
and U21805 (N_21805,N_21394,N_21111);
nand U21806 (N_21806,N_21327,N_21223);
and U21807 (N_21807,N_21088,N_21213);
nand U21808 (N_21808,N_21142,N_21337);
xnor U21809 (N_21809,N_21366,N_21182);
nor U21810 (N_21810,N_21010,N_21472);
xnor U21811 (N_21811,N_21237,N_21197);
or U21812 (N_21812,N_21070,N_21035);
nand U21813 (N_21813,N_21156,N_21049);
xnor U21814 (N_21814,N_21257,N_21390);
xor U21815 (N_21815,N_21193,N_21303);
xnor U21816 (N_21816,N_21393,N_21244);
nor U21817 (N_21817,N_21398,N_21102);
or U21818 (N_21818,N_21316,N_21180);
xnor U21819 (N_21819,N_21105,N_21230);
or U21820 (N_21820,N_21089,N_21415);
and U21821 (N_21821,N_21369,N_21014);
or U21822 (N_21822,N_21400,N_21259);
and U21823 (N_21823,N_21458,N_21103);
nand U21824 (N_21824,N_21064,N_21284);
nand U21825 (N_21825,N_21196,N_21185);
or U21826 (N_21826,N_21421,N_21049);
and U21827 (N_21827,N_21315,N_21350);
xnor U21828 (N_21828,N_21054,N_21150);
nand U21829 (N_21829,N_21344,N_21491);
and U21830 (N_21830,N_21066,N_21136);
nor U21831 (N_21831,N_21258,N_21367);
nor U21832 (N_21832,N_21088,N_21124);
and U21833 (N_21833,N_21432,N_21044);
and U21834 (N_21834,N_21121,N_21179);
nand U21835 (N_21835,N_21052,N_21447);
and U21836 (N_21836,N_21450,N_21423);
and U21837 (N_21837,N_21413,N_21208);
and U21838 (N_21838,N_21217,N_21380);
xor U21839 (N_21839,N_21130,N_21302);
nor U21840 (N_21840,N_21171,N_21286);
nand U21841 (N_21841,N_21148,N_21357);
nand U21842 (N_21842,N_21026,N_21195);
xnor U21843 (N_21843,N_21483,N_21264);
or U21844 (N_21844,N_21229,N_21484);
nand U21845 (N_21845,N_21323,N_21344);
xor U21846 (N_21846,N_21415,N_21023);
xnor U21847 (N_21847,N_21252,N_21327);
xor U21848 (N_21848,N_21393,N_21299);
nand U21849 (N_21849,N_21364,N_21213);
or U21850 (N_21850,N_21159,N_21326);
and U21851 (N_21851,N_21257,N_21140);
nor U21852 (N_21852,N_21437,N_21061);
nor U21853 (N_21853,N_21263,N_21338);
and U21854 (N_21854,N_21161,N_21102);
and U21855 (N_21855,N_21289,N_21406);
nor U21856 (N_21856,N_21324,N_21174);
or U21857 (N_21857,N_21350,N_21384);
xnor U21858 (N_21858,N_21342,N_21366);
nor U21859 (N_21859,N_21470,N_21479);
xor U21860 (N_21860,N_21214,N_21404);
and U21861 (N_21861,N_21323,N_21484);
and U21862 (N_21862,N_21114,N_21486);
nand U21863 (N_21863,N_21184,N_21104);
nand U21864 (N_21864,N_21343,N_21224);
or U21865 (N_21865,N_21254,N_21212);
nand U21866 (N_21866,N_21334,N_21223);
and U21867 (N_21867,N_21286,N_21351);
or U21868 (N_21868,N_21039,N_21411);
nand U21869 (N_21869,N_21152,N_21250);
or U21870 (N_21870,N_21016,N_21128);
xnor U21871 (N_21871,N_21169,N_21474);
nand U21872 (N_21872,N_21136,N_21058);
or U21873 (N_21873,N_21145,N_21370);
nor U21874 (N_21874,N_21110,N_21151);
nand U21875 (N_21875,N_21139,N_21486);
nor U21876 (N_21876,N_21129,N_21421);
nand U21877 (N_21877,N_21394,N_21090);
nor U21878 (N_21878,N_21422,N_21183);
or U21879 (N_21879,N_21042,N_21271);
nor U21880 (N_21880,N_21235,N_21490);
nand U21881 (N_21881,N_21057,N_21241);
or U21882 (N_21882,N_21318,N_21480);
nand U21883 (N_21883,N_21103,N_21203);
nand U21884 (N_21884,N_21365,N_21406);
and U21885 (N_21885,N_21429,N_21480);
nand U21886 (N_21886,N_21483,N_21428);
xor U21887 (N_21887,N_21431,N_21004);
nor U21888 (N_21888,N_21342,N_21009);
nand U21889 (N_21889,N_21294,N_21012);
xnor U21890 (N_21890,N_21213,N_21139);
nor U21891 (N_21891,N_21485,N_21413);
xor U21892 (N_21892,N_21297,N_21105);
and U21893 (N_21893,N_21140,N_21406);
nand U21894 (N_21894,N_21114,N_21142);
or U21895 (N_21895,N_21381,N_21432);
nor U21896 (N_21896,N_21341,N_21195);
or U21897 (N_21897,N_21267,N_21163);
nor U21898 (N_21898,N_21212,N_21195);
and U21899 (N_21899,N_21107,N_21391);
or U21900 (N_21900,N_21015,N_21141);
nor U21901 (N_21901,N_21388,N_21196);
nand U21902 (N_21902,N_21188,N_21375);
and U21903 (N_21903,N_21451,N_21329);
or U21904 (N_21904,N_21489,N_21403);
xor U21905 (N_21905,N_21006,N_21377);
nor U21906 (N_21906,N_21401,N_21080);
nand U21907 (N_21907,N_21234,N_21463);
and U21908 (N_21908,N_21071,N_21133);
and U21909 (N_21909,N_21410,N_21021);
and U21910 (N_21910,N_21423,N_21269);
or U21911 (N_21911,N_21348,N_21258);
nand U21912 (N_21912,N_21300,N_21319);
and U21913 (N_21913,N_21409,N_21333);
and U21914 (N_21914,N_21118,N_21342);
nor U21915 (N_21915,N_21458,N_21235);
nand U21916 (N_21916,N_21431,N_21260);
nand U21917 (N_21917,N_21193,N_21345);
nor U21918 (N_21918,N_21181,N_21384);
nand U21919 (N_21919,N_21405,N_21456);
nand U21920 (N_21920,N_21249,N_21113);
and U21921 (N_21921,N_21144,N_21181);
or U21922 (N_21922,N_21219,N_21446);
and U21923 (N_21923,N_21143,N_21375);
and U21924 (N_21924,N_21271,N_21081);
xor U21925 (N_21925,N_21003,N_21054);
nand U21926 (N_21926,N_21433,N_21477);
xnor U21927 (N_21927,N_21119,N_21397);
nand U21928 (N_21928,N_21171,N_21024);
nor U21929 (N_21929,N_21152,N_21137);
nand U21930 (N_21930,N_21143,N_21247);
or U21931 (N_21931,N_21280,N_21336);
nor U21932 (N_21932,N_21025,N_21461);
or U21933 (N_21933,N_21389,N_21050);
or U21934 (N_21934,N_21177,N_21438);
and U21935 (N_21935,N_21210,N_21056);
nand U21936 (N_21936,N_21077,N_21263);
nand U21937 (N_21937,N_21447,N_21100);
xnor U21938 (N_21938,N_21244,N_21169);
nor U21939 (N_21939,N_21343,N_21414);
nor U21940 (N_21940,N_21456,N_21356);
nand U21941 (N_21941,N_21285,N_21349);
nand U21942 (N_21942,N_21216,N_21011);
and U21943 (N_21943,N_21120,N_21187);
nand U21944 (N_21944,N_21095,N_21044);
xnor U21945 (N_21945,N_21485,N_21244);
or U21946 (N_21946,N_21289,N_21251);
nand U21947 (N_21947,N_21140,N_21272);
xor U21948 (N_21948,N_21255,N_21490);
xnor U21949 (N_21949,N_21116,N_21114);
nand U21950 (N_21950,N_21409,N_21031);
or U21951 (N_21951,N_21440,N_21231);
and U21952 (N_21952,N_21204,N_21091);
and U21953 (N_21953,N_21159,N_21325);
and U21954 (N_21954,N_21279,N_21244);
and U21955 (N_21955,N_21169,N_21252);
xnor U21956 (N_21956,N_21357,N_21317);
or U21957 (N_21957,N_21399,N_21322);
and U21958 (N_21958,N_21177,N_21012);
nor U21959 (N_21959,N_21194,N_21331);
xor U21960 (N_21960,N_21133,N_21097);
and U21961 (N_21961,N_21421,N_21391);
xor U21962 (N_21962,N_21002,N_21232);
or U21963 (N_21963,N_21384,N_21171);
nand U21964 (N_21964,N_21309,N_21438);
nor U21965 (N_21965,N_21032,N_21008);
nor U21966 (N_21966,N_21083,N_21244);
nor U21967 (N_21967,N_21011,N_21040);
nor U21968 (N_21968,N_21415,N_21476);
xnor U21969 (N_21969,N_21282,N_21431);
nor U21970 (N_21970,N_21088,N_21467);
xnor U21971 (N_21971,N_21211,N_21048);
or U21972 (N_21972,N_21123,N_21493);
and U21973 (N_21973,N_21423,N_21299);
and U21974 (N_21974,N_21177,N_21419);
xor U21975 (N_21975,N_21003,N_21315);
nand U21976 (N_21976,N_21267,N_21259);
or U21977 (N_21977,N_21190,N_21400);
and U21978 (N_21978,N_21377,N_21442);
nor U21979 (N_21979,N_21193,N_21289);
or U21980 (N_21980,N_21417,N_21069);
or U21981 (N_21981,N_21338,N_21285);
xor U21982 (N_21982,N_21075,N_21207);
nor U21983 (N_21983,N_21384,N_21051);
nand U21984 (N_21984,N_21201,N_21156);
or U21985 (N_21985,N_21155,N_21339);
or U21986 (N_21986,N_21025,N_21239);
xor U21987 (N_21987,N_21343,N_21335);
and U21988 (N_21988,N_21410,N_21071);
nor U21989 (N_21989,N_21481,N_21060);
nor U21990 (N_21990,N_21004,N_21391);
nor U21991 (N_21991,N_21254,N_21269);
and U21992 (N_21992,N_21221,N_21082);
and U21993 (N_21993,N_21302,N_21028);
and U21994 (N_21994,N_21212,N_21166);
nor U21995 (N_21995,N_21186,N_21197);
and U21996 (N_21996,N_21371,N_21209);
nand U21997 (N_21997,N_21100,N_21445);
nor U21998 (N_21998,N_21076,N_21297);
nand U21999 (N_21999,N_21493,N_21171);
and U22000 (N_22000,N_21746,N_21502);
or U22001 (N_22001,N_21928,N_21964);
nand U22002 (N_22002,N_21798,N_21622);
and U22003 (N_22003,N_21674,N_21958);
xnor U22004 (N_22004,N_21676,N_21870);
or U22005 (N_22005,N_21763,N_21857);
and U22006 (N_22006,N_21514,N_21846);
nor U22007 (N_22007,N_21861,N_21702);
and U22008 (N_22008,N_21799,N_21523);
nor U22009 (N_22009,N_21758,N_21717);
nor U22010 (N_22010,N_21696,N_21524);
nor U22011 (N_22011,N_21729,N_21781);
xnor U22012 (N_22012,N_21567,N_21780);
xnor U22013 (N_22013,N_21990,N_21645);
nand U22014 (N_22014,N_21697,N_21710);
nor U22015 (N_22015,N_21641,N_21991);
nor U22016 (N_22016,N_21621,N_21659);
and U22017 (N_22017,N_21751,N_21685);
and U22018 (N_22018,N_21898,N_21508);
or U22019 (N_22019,N_21627,N_21752);
nand U22020 (N_22020,N_21842,N_21765);
nor U22021 (N_22021,N_21698,N_21694);
or U22022 (N_22022,N_21713,N_21716);
and U22023 (N_22023,N_21580,N_21885);
nand U22024 (N_22024,N_21550,N_21691);
and U22025 (N_22025,N_21663,N_21814);
xor U22026 (N_22026,N_21932,N_21981);
nand U22027 (N_22027,N_21712,N_21644);
and U22028 (N_22028,N_21678,N_21849);
and U22029 (N_22029,N_21908,N_21989);
nor U22030 (N_22030,N_21528,N_21606);
nor U22031 (N_22031,N_21625,N_21777);
and U22032 (N_22032,N_21724,N_21655);
nand U22033 (N_22033,N_21934,N_21553);
and U22034 (N_22034,N_21791,N_21882);
xor U22035 (N_22035,N_21992,N_21608);
or U22036 (N_22036,N_21918,N_21692);
nand U22037 (N_22037,N_21688,N_21996);
nand U22038 (N_22038,N_21834,N_21795);
or U22039 (N_22039,N_21852,N_21985);
nand U22040 (N_22040,N_21792,N_21684);
nand U22041 (N_22041,N_21582,N_21821);
or U22042 (N_22042,N_21966,N_21660);
nor U22043 (N_22043,N_21703,N_21771);
nand U22044 (N_22044,N_21636,N_21920);
nor U22045 (N_22045,N_21755,N_21612);
nand U22046 (N_22046,N_21673,N_21778);
or U22047 (N_22047,N_21839,N_21914);
and U22048 (N_22048,N_21727,N_21672);
and U22049 (N_22049,N_21749,N_21573);
and U22050 (N_22050,N_21590,N_21761);
and U22051 (N_22051,N_21578,N_21706);
nand U22052 (N_22052,N_21650,N_21723);
nand U22053 (N_22053,N_21939,N_21665);
nand U22054 (N_22054,N_21824,N_21734);
nor U22055 (N_22055,N_21569,N_21828);
and U22056 (N_22056,N_21649,N_21767);
and U22057 (N_22057,N_21974,N_21630);
xor U22058 (N_22058,N_21776,N_21922);
nand U22059 (N_22059,N_21651,N_21880);
xnor U22060 (N_22060,N_21804,N_21620);
and U22061 (N_22061,N_21744,N_21613);
and U22062 (N_22062,N_21875,N_21653);
and U22063 (N_22063,N_21754,N_21813);
xor U22064 (N_22064,N_21959,N_21552);
nor U22065 (N_22065,N_21982,N_21980);
xor U22066 (N_22066,N_21519,N_21619);
nand U22067 (N_22067,N_21969,N_21575);
nand U22068 (N_22068,N_21938,N_21884);
xnor U22069 (N_22069,N_21994,N_21512);
or U22070 (N_22070,N_21815,N_21930);
nor U22071 (N_22071,N_21633,N_21785);
nor U22072 (N_22072,N_21701,N_21949);
nor U22073 (N_22073,N_21889,N_21711);
xnor U22074 (N_22074,N_21978,N_21988);
nand U22075 (N_22075,N_21681,N_21592);
nor U22076 (N_22076,N_21647,N_21566);
or U22077 (N_22077,N_21855,N_21823);
nand U22078 (N_22078,N_21586,N_21869);
nand U22079 (N_22079,N_21635,N_21944);
xor U22080 (N_22080,N_21877,N_21585);
and U22081 (N_22081,N_21549,N_21841);
and U22082 (N_22082,N_21913,N_21768);
or U22083 (N_22083,N_21505,N_21570);
xor U22084 (N_22084,N_21682,N_21967);
nand U22085 (N_22085,N_21563,N_21530);
or U22086 (N_22086,N_21733,N_21952);
xor U22087 (N_22087,N_21597,N_21794);
nor U22088 (N_22088,N_21551,N_21888);
xor U22089 (N_22089,N_21976,N_21533);
nor U22090 (N_22090,N_21793,N_21788);
xnor U22091 (N_22091,N_21854,N_21762);
or U22092 (N_22092,N_21851,N_21873);
nand U22093 (N_22093,N_21916,N_21624);
nor U22094 (N_22094,N_21693,N_21862);
nand U22095 (N_22095,N_21741,N_21829);
or U22096 (N_22096,N_21859,N_21933);
nand U22097 (N_22097,N_21720,N_21843);
or U22098 (N_22098,N_21591,N_21626);
xor U22099 (N_22099,N_21666,N_21790);
nand U22100 (N_22100,N_21912,N_21543);
nor U22101 (N_22101,N_21574,N_21929);
nand U22102 (N_22102,N_21902,N_21558);
or U22103 (N_22103,N_21517,N_21511);
or U22104 (N_22104,N_21965,N_21628);
nor U22105 (N_22105,N_21953,N_21601);
nor U22106 (N_22106,N_21501,N_21850);
and U22107 (N_22107,N_21972,N_21556);
nand U22108 (N_22108,N_21547,N_21775);
nand U22109 (N_22109,N_21560,N_21836);
and U22110 (N_22110,N_21631,N_21686);
and U22111 (N_22111,N_21867,N_21577);
xnor U22112 (N_22112,N_21652,N_21707);
and U22113 (N_22113,N_21808,N_21899);
and U22114 (N_22114,N_21516,N_21950);
nand U22115 (N_22115,N_21531,N_21943);
nand U22116 (N_22116,N_21689,N_21872);
and U22117 (N_22117,N_21871,N_21941);
xnor U22118 (N_22118,N_21787,N_21894);
or U22119 (N_22119,N_21675,N_21936);
or U22120 (N_22120,N_21866,N_21891);
or U22121 (N_22121,N_21818,N_21605);
and U22122 (N_22122,N_21838,N_21856);
nand U22123 (N_22123,N_21725,N_21748);
nor U22124 (N_22124,N_21984,N_21742);
or U22125 (N_22125,N_21957,N_21800);
and U22126 (N_22126,N_21561,N_21640);
xor U22127 (N_22127,N_21811,N_21786);
and U22128 (N_22128,N_21886,N_21895);
xor U22129 (N_22129,N_21537,N_21588);
nand U22130 (N_22130,N_21709,N_21714);
or U22131 (N_22131,N_21639,N_21518);
nand U22132 (N_22132,N_21542,N_21618);
or U22133 (N_22133,N_21648,N_21764);
and U22134 (N_22134,N_21983,N_21789);
nand U22135 (N_22135,N_21946,N_21515);
or U22136 (N_22136,N_21721,N_21921);
xnor U22137 (N_22137,N_21743,N_21832);
nand U22138 (N_22138,N_21739,N_21555);
nand U22139 (N_22139,N_21773,N_21679);
and U22140 (N_22140,N_21510,N_21812);
nand U22141 (N_22141,N_21544,N_21840);
and U22142 (N_22142,N_21683,N_21993);
nand U22143 (N_22143,N_21504,N_21760);
and U22144 (N_22144,N_21509,N_21632);
nor U22145 (N_22145,N_21925,N_21909);
nand U22146 (N_22146,N_21522,N_21817);
and U22147 (N_22147,N_21945,N_21826);
and U22148 (N_22148,N_21587,N_21593);
nand U22149 (N_22149,N_21779,N_21680);
nand U22150 (N_22150,N_21833,N_21545);
or U22151 (N_22151,N_21548,N_21796);
nor U22152 (N_22152,N_21919,N_21557);
or U22153 (N_22153,N_21878,N_21726);
nor U22154 (N_22154,N_21998,N_21503);
nor U22155 (N_22155,N_21968,N_21669);
and U22156 (N_22156,N_21735,N_21784);
xor U22157 (N_22157,N_21890,N_21745);
xnor U22158 (N_22158,N_21667,N_21687);
and U22159 (N_22159,N_21718,N_21816);
or U22160 (N_22160,N_21584,N_21797);
nand U22161 (N_22161,N_21610,N_21893);
nor U22162 (N_22162,N_21576,N_21532);
and U22163 (N_22163,N_21661,N_21642);
or U22164 (N_22164,N_21907,N_21614);
or U22165 (N_22165,N_21973,N_21772);
xor U22166 (N_22166,N_21623,N_21847);
nand U22167 (N_22167,N_21602,N_21535);
or U22168 (N_22168,N_21940,N_21534);
xor U22169 (N_22169,N_21705,N_21617);
nor U22170 (N_22170,N_21951,N_21599);
and U22171 (N_22171,N_21579,N_21960);
xnor U22172 (N_22172,N_21848,N_21737);
nand U22173 (N_22173,N_21831,N_21708);
xor U22174 (N_22174,N_21507,N_21924);
and U22175 (N_22175,N_21759,N_21520);
nand U22176 (N_22176,N_21783,N_21970);
nor U22177 (N_22177,N_21658,N_21900);
and U22178 (N_22178,N_21637,N_21883);
nand U22179 (N_22179,N_21529,N_21695);
nor U22180 (N_22180,N_21947,N_21802);
and U22181 (N_22181,N_21954,N_21564);
or U22182 (N_22182,N_21897,N_21906);
nor U22183 (N_22183,N_21677,N_21730);
nor U22184 (N_22184,N_21923,N_21948);
nor U22185 (N_22185,N_21756,N_21657);
or U22186 (N_22186,N_21589,N_21803);
nor U22187 (N_22187,N_21971,N_21917);
or U22188 (N_22188,N_21559,N_21513);
xnor U22189 (N_22189,N_21634,N_21654);
and U22190 (N_22190,N_21845,N_21874);
xor U22191 (N_22191,N_21963,N_21562);
nor U22192 (N_22192,N_21604,N_21603);
or U22193 (N_22193,N_21753,N_21671);
or U22194 (N_22194,N_21595,N_21827);
nand U22195 (N_22195,N_21807,N_21736);
or U22196 (N_22196,N_21668,N_21820);
or U22197 (N_22197,N_21805,N_21926);
nor U22198 (N_22198,N_21643,N_21616);
and U22199 (N_22199,N_21525,N_21664);
or U22200 (N_22200,N_21722,N_21809);
xor U22201 (N_22201,N_21546,N_21782);
or U22202 (N_22202,N_21868,N_21961);
or U22203 (N_22203,N_21937,N_21757);
nand U22204 (N_22204,N_21905,N_21719);
nor U22205 (N_22205,N_21987,N_21629);
nand U22206 (N_22206,N_21837,N_21738);
or U22207 (N_22207,N_21853,N_21704);
or U22208 (N_22208,N_21690,N_21931);
and U22209 (N_22209,N_21646,N_21822);
and U22210 (N_22210,N_21806,N_21801);
or U22211 (N_22211,N_21670,N_21825);
and U22212 (N_22212,N_21747,N_21609);
nand U22213 (N_22213,N_21858,N_21863);
and U22214 (N_22214,N_21770,N_21568);
nor U22215 (N_22215,N_21892,N_21810);
xor U22216 (N_22216,N_21500,N_21999);
nor U22217 (N_22217,N_21699,N_21526);
or U22218 (N_22218,N_21541,N_21750);
nand U22219 (N_22219,N_21506,N_21975);
or U22220 (N_22220,N_21977,N_21540);
xor U22221 (N_22221,N_21731,N_21881);
nor U22222 (N_22222,N_21835,N_21728);
nand U22223 (N_22223,N_21903,N_21819);
or U22224 (N_22224,N_21527,N_21774);
nand U22225 (N_22225,N_21769,N_21955);
and U22226 (N_22226,N_21732,N_21662);
nor U22227 (N_22227,N_21956,N_21554);
and U22228 (N_22228,N_21700,N_21844);
and U22229 (N_22229,N_21521,N_21638);
and U22230 (N_22230,N_21995,N_21865);
nand U22231 (N_22231,N_21997,N_21910);
nor U22232 (N_22232,N_21876,N_21860);
xor U22233 (N_22233,N_21927,N_21896);
and U22234 (N_22234,N_21571,N_21830);
and U22235 (N_22235,N_21539,N_21536);
nand U22236 (N_22236,N_21901,N_21887);
and U22237 (N_22237,N_21942,N_21565);
nor U22238 (N_22238,N_21600,N_21766);
nand U22239 (N_22239,N_21864,N_21607);
nor U22240 (N_22240,N_21715,N_21935);
nand U22241 (N_22241,N_21611,N_21656);
nor U22242 (N_22242,N_21598,N_21879);
nor U22243 (N_22243,N_21572,N_21594);
xor U22244 (N_22244,N_21979,N_21986);
nor U22245 (N_22245,N_21904,N_21615);
nor U22246 (N_22246,N_21911,N_21581);
nand U22247 (N_22247,N_21538,N_21583);
and U22248 (N_22248,N_21740,N_21962);
xnor U22249 (N_22249,N_21596,N_21915);
xnor U22250 (N_22250,N_21900,N_21772);
nor U22251 (N_22251,N_21990,N_21501);
nand U22252 (N_22252,N_21666,N_21861);
nand U22253 (N_22253,N_21722,N_21572);
or U22254 (N_22254,N_21596,N_21697);
nor U22255 (N_22255,N_21959,N_21862);
and U22256 (N_22256,N_21777,N_21727);
or U22257 (N_22257,N_21701,N_21502);
xor U22258 (N_22258,N_21995,N_21600);
and U22259 (N_22259,N_21695,N_21843);
or U22260 (N_22260,N_21596,N_21785);
nor U22261 (N_22261,N_21623,N_21678);
nor U22262 (N_22262,N_21562,N_21980);
xnor U22263 (N_22263,N_21743,N_21580);
xnor U22264 (N_22264,N_21832,N_21694);
nand U22265 (N_22265,N_21740,N_21950);
xor U22266 (N_22266,N_21809,N_21529);
and U22267 (N_22267,N_21771,N_21664);
and U22268 (N_22268,N_21606,N_21508);
xnor U22269 (N_22269,N_21781,N_21957);
or U22270 (N_22270,N_21994,N_21669);
or U22271 (N_22271,N_21938,N_21994);
nand U22272 (N_22272,N_21596,N_21549);
or U22273 (N_22273,N_21592,N_21910);
xor U22274 (N_22274,N_21746,N_21566);
nor U22275 (N_22275,N_21604,N_21722);
nand U22276 (N_22276,N_21864,N_21525);
or U22277 (N_22277,N_21771,N_21776);
and U22278 (N_22278,N_21749,N_21789);
xnor U22279 (N_22279,N_21996,N_21965);
or U22280 (N_22280,N_21738,N_21799);
or U22281 (N_22281,N_21791,N_21900);
xnor U22282 (N_22282,N_21809,N_21862);
and U22283 (N_22283,N_21587,N_21762);
xnor U22284 (N_22284,N_21697,N_21849);
nor U22285 (N_22285,N_21809,N_21587);
xnor U22286 (N_22286,N_21591,N_21643);
xor U22287 (N_22287,N_21528,N_21909);
and U22288 (N_22288,N_21953,N_21991);
xor U22289 (N_22289,N_21527,N_21804);
nand U22290 (N_22290,N_21906,N_21511);
or U22291 (N_22291,N_21966,N_21946);
or U22292 (N_22292,N_21915,N_21995);
and U22293 (N_22293,N_21675,N_21615);
nand U22294 (N_22294,N_21970,N_21733);
xnor U22295 (N_22295,N_21595,N_21907);
nor U22296 (N_22296,N_21603,N_21905);
and U22297 (N_22297,N_21560,N_21984);
nand U22298 (N_22298,N_21622,N_21942);
or U22299 (N_22299,N_21556,N_21682);
xor U22300 (N_22300,N_21737,N_21853);
or U22301 (N_22301,N_21875,N_21635);
nand U22302 (N_22302,N_21738,N_21770);
xor U22303 (N_22303,N_21872,N_21576);
xor U22304 (N_22304,N_21635,N_21725);
nor U22305 (N_22305,N_21733,N_21772);
nand U22306 (N_22306,N_21797,N_21616);
nand U22307 (N_22307,N_21538,N_21778);
or U22308 (N_22308,N_21694,N_21557);
xnor U22309 (N_22309,N_21582,N_21716);
nor U22310 (N_22310,N_21761,N_21583);
nand U22311 (N_22311,N_21809,N_21921);
and U22312 (N_22312,N_21940,N_21690);
xor U22313 (N_22313,N_21663,N_21662);
xor U22314 (N_22314,N_21717,N_21781);
nor U22315 (N_22315,N_21771,N_21874);
nand U22316 (N_22316,N_21997,N_21913);
nor U22317 (N_22317,N_21864,N_21683);
nand U22318 (N_22318,N_21809,N_21922);
and U22319 (N_22319,N_21655,N_21670);
nor U22320 (N_22320,N_21710,N_21612);
nand U22321 (N_22321,N_21838,N_21882);
nand U22322 (N_22322,N_21504,N_21633);
or U22323 (N_22323,N_21576,N_21611);
and U22324 (N_22324,N_21987,N_21628);
and U22325 (N_22325,N_21573,N_21994);
xor U22326 (N_22326,N_21837,N_21515);
nor U22327 (N_22327,N_21637,N_21818);
nand U22328 (N_22328,N_21947,N_21512);
nor U22329 (N_22329,N_21932,N_21744);
xor U22330 (N_22330,N_21989,N_21775);
xnor U22331 (N_22331,N_21883,N_21780);
or U22332 (N_22332,N_21949,N_21971);
and U22333 (N_22333,N_21744,N_21631);
or U22334 (N_22334,N_21754,N_21938);
nor U22335 (N_22335,N_21728,N_21647);
nand U22336 (N_22336,N_21680,N_21606);
nor U22337 (N_22337,N_21828,N_21509);
and U22338 (N_22338,N_21715,N_21870);
xor U22339 (N_22339,N_21801,N_21993);
or U22340 (N_22340,N_21673,N_21764);
nor U22341 (N_22341,N_21941,N_21734);
and U22342 (N_22342,N_21577,N_21789);
and U22343 (N_22343,N_21594,N_21727);
nor U22344 (N_22344,N_21825,N_21861);
nand U22345 (N_22345,N_21771,N_21561);
nand U22346 (N_22346,N_21590,N_21911);
nand U22347 (N_22347,N_21828,N_21834);
nand U22348 (N_22348,N_21982,N_21819);
xor U22349 (N_22349,N_21887,N_21872);
xnor U22350 (N_22350,N_21781,N_21502);
or U22351 (N_22351,N_21942,N_21761);
nor U22352 (N_22352,N_21594,N_21781);
and U22353 (N_22353,N_21789,N_21656);
nor U22354 (N_22354,N_21615,N_21843);
xnor U22355 (N_22355,N_21894,N_21667);
nor U22356 (N_22356,N_21823,N_21593);
and U22357 (N_22357,N_21563,N_21606);
nor U22358 (N_22358,N_21965,N_21615);
xnor U22359 (N_22359,N_21874,N_21615);
nand U22360 (N_22360,N_21771,N_21980);
or U22361 (N_22361,N_21635,N_21865);
or U22362 (N_22362,N_21929,N_21844);
nand U22363 (N_22363,N_21763,N_21546);
and U22364 (N_22364,N_21823,N_21696);
or U22365 (N_22365,N_21571,N_21697);
xor U22366 (N_22366,N_21758,N_21751);
xor U22367 (N_22367,N_21841,N_21769);
and U22368 (N_22368,N_21734,N_21582);
and U22369 (N_22369,N_21511,N_21730);
nand U22370 (N_22370,N_21666,N_21896);
and U22371 (N_22371,N_21980,N_21834);
xnor U22372 (N_22372,N_21838,N_21635);
xor U22373 (N_22373,N_21877,N_21933);
or U22374 (N_22374,N_21966,N_21836);
and U22375 (N_22375,N_21946,N_21587);
or U22376 (N_22376,N_21927,N_21593);
xnor U22377 (N_22377,N_21695,N_21591);
nand U22378 (N_22378,N_21591,N_21909);
and U22379 (N_22379,N_21778,N_21891);
or U22380 (N_22380,N_21797,N_21827);
or U22381 (N_22381,N_21751,N_21777);
nand U22382 (N_22382,N_21711,N_21639);
xor U22383 (N_22383,N_21616,N_21612);
xnor U22384 (N_22384,N_21937,N_21710);
or U22385 (N_22385,N_21606,N_21604);
nor U22386 (N_22386,N_21668,N_21718);
nor U22387 (N_22387,N_21545,N_21839);
nor U22388 (N_22388,N_21598,N_21792);
nand U22389 (N_22389,N_21857,N_21824);
and U22390 (N_22390,N_21793,N_21946);
nor U22391 (N_22391,N_21782,N_21935);
nor U22392 (N_22392,N_21776,N_21526);
or U22393 (N_22393,N_21837,N_21545);
nand U22394 (N_22394,N_21871,N_21608);
nand U22395 (N_22395,N_21830,N_21584);
nand U22396 (N_22396,N_21656,N_21555);
nand U22397 (N_22397,N_21712,N_21734);
or U22398 (N_22398,N_21530,N_21919);
or U22399 (N_22399,N_21696,N_21520);
or U22400 (N_22400,N_21749,N_21714);
nand U22401 (N_22401,N_21883,N_21723);
nand U22402 (N_22402,N_21997,N_21675);
nor U22403 (N_22403,N_21697,N_21907);
nand U22404 (N_22404,N_21656,N_21670);
xor U22405 (N_22405,N_21574,N_21738);
nand U22406 (N_22406,N_21829,N_21858);
or U22407 (N_22407,N_21873,N_21634);
xor U22408 (N_22408,N_21763,N_21785);
xnor U22409 (N_22409,N_21601,N_21724);
and U22410 (N_22410,N_21676,N_21846);
nor U22411 (N_22411,N_21615,N_21731);
nand U22412 (N_22412,N_21722,N_21856);
or U22413 (N_22413,N_21550,N_21749);
and U22414 (N_22414,N_21585,N_21947);
and U22415 (N_22415,N_21865,N_21910);
nor U22416 (N_22416,N_21889,N_21669);
xnor U22417 (N_22417,N_21676,N_21656);
nand U22418 (N_22418,N_21855,N_21554);
xnor U22419 (N_22419,N_21657,N_21603);
and U22420 (N_22420,N_21819,N_21734);
and U22421 (N_22421,N_21770,N_21614);
xor U22422 (N_22422,N_21659,N_21827);
or U22423 (N_22423,N_21895,N_21965);
and U22424 (N_22424,N_21865,N_21534);
or U22425 (N_22425,N_21737,N_21716);
and U22426 (N_22426,N_21890,N_21818);
nand U22427 (N_22427,N_21723,N_21552);
and U22428 (N_22428,N_21697,N_21846);
xor U22429 (N_22429,N_21933,N_21817);
xor U22430 (N_22430,N_21707,N_21578);
and U22431 (N_22431,N_21959,N_21991);
and U22432 (N_22432,N_21700,N_21552);
nand U22433 (N_22433,N_21993,N_21655);
or U22434 (N_22434,N_21558,N_21591);
or U22435 (N_22435,N_21924,N_21995);
nand U22436 (N_22436,N_21685,N_21509);
or U22437 (N_22437,N_21975,N_21888);
nand U22438 (N_22438,N_21853,N_21940);
xnor U22439 (N_22439,N_21738,N_21591);
or U22440 (N_22440,N_21966,N_21532);
or U22441 (N_22441,N_21812,N_21674);
nand U22442 (N_22442,N_21814,N_21778);
nor U22443 (N_22443,N_21933,N_21636);
and U22444 (N_22444,N_21888,N_21877);
xnor U22445 (N_22445,N_21699,N_21908);
nand U22446 (N_22446,N_21758,N_21523);
nor U22447 (N_22447,N_21792,N_21765);
or U22448 (N_22448,N_21610,N_21665);
xor U22449 (N_22449,N_21865,N_21943);
xor U22450 (N_22450,N_21800,N_21714);
nor U22451 (N_22451,N_21924,N_21984);
and U22452 (N_22452,N_21741,N_21567);
xor U22453 (N_22453,N_21972,N_21670);
xnor U22454 (N_22454,N_21996,N_21841);
nor U22455 (N_22455,N_21713,N_21796);
nand U22456 (N_22456,N_21515,N_21957);
and U22457 (N_22457,N_21815,N_21558);
and U22458 (N_22458,N_21693,N_21788);
and U22459 (N_22459,N_21753,N_21663);
xor U22460 (N_22460,N_21762,N_21781);
xnor U22461 (N_22461,N_21646,N_21814);
and U22462 (N_22462,N_21829,N_21544);
xor U22463 (N_22463,N_21972,N_21898);
nand U22464 (N_22464,N_21831,N_21635);
and U22465 (N_22465,N_21512,N_21951);
nand U22466 (N_22466,N_21798,N_21718);
and U22467 (N_22467,N_21713,N_21544);
nand U22468 (N_22468,N_21757,N_21640);
nand U22469 (N_22469,N_21615,N_21637);
nor U22470 (N_22470,N_21953,N_21961);
nor U22471 (N_22471,N_21650,N_21947);
xnor U22472 (N_22472,N_21732,N_21809);
nand U22473 (N_22473,N_21726,N_21939);
nor U22474 (N_22474,N_21898,N_21703);
xnor U22475 (N_22475,N_21791,N_21737);
nor U22476 (N_22476,N_21727,N_21900);
nand U22477 (N_22477,N_21848,N_21562);
nand U22478 (N_22478,N_21647,N_21617);
nor U22479 (N_22479,N_21567,N_21893);
or U22480 (N_22480,N_21816,N_21685);
nor U22481 (N_22481,N_21997,N_21669);
nor U22482 (N_22482,N_21749,N_21870);
nand U22483 (N_22483,N_21595,N_21788);
xnor U22484 (N_22484,N_21860,N_21541);
or U22485 (N_22485,N_21907,N_21977);
or U22486 (N_22486,N_21782,N_21518);
and U22487 (N_22487,N_21548,N_21794);
xor U22488 (N_22488,N_21561,N_21927);
and U22489 (N_22489,N_21665,N_21528);
or U22490 (N_22490,N_21995,N_21900);
and U22491 (N_22491,N_21562,N_21703);
nand U22492 (N_22492,N_21505,N_21843);
nor U22493 (N_22493,N_21888,N_21846);
nand U22494 (N_22494,N_21752,N_21658);
and U22495 (N_22495,N_21894,N_21741);
and U22496 (N_22496,N_21754,N_21942);
nor U22497 (N_22497,N_21685,N_21720);
nand U22498 (N_22498,N_21580,N_21659);
and U22499 (N_22499,N_21771,N_21997);
or U22500 (N_22500,N_22411,N_22474);
xnor U22501 (N_22501,N_22337,N_22428);
and U22502 (N_22502,N_22087,N_22181);
nor U22503 (N_22503,N_22231,N_22040);
xnor U22504 (N_22504,N_22435,N_22028);
and U22505 (N_22505,N_22234,N_22020);
nand U22506 (N_22506,N_22425,N_22339);
and U22507 (N_22507,N_22328,N_22356);
xnor U22508 (N_22508,N_22168,N_22045);
xnor U22509 (N_22509,N_22111,N_22324);
or U22510 (N_22510,N_22270,N_22475);
or U22511 (N_22511,N_22352,N_22497);
nor U22512 (N_22512,N_22414,N_22316);
nand U22513 (N_22513,N_22333,N_22321);
nor U22514 (N_22514,N_22467,N_22229);
xnor U22515 (N_22515,N_22479,N_22335);
nor U22516 (N_22516,N_22043,N_22495);
or U22517 (N_22517,N_22017,N_22301);
nor U22518 (N_22518,N_22484,N_22275);
nand U22519 (N_22519,N_22126,N_22355);
xnor U22520 (N_22520,N_22399,N_22451);
nor U22521 (N_22521,N_22359,N_22167);
or U22522 (N_22522,N_22032,N_22282);
or U22523 (N_22523,N_22315,N_22420);
nand U22524 (N_22524,N_22009,N_22292);
nor U22525 (N_22525,N_22320,N_22144);
nor U22526 (N_22526,N_22225,N_22308);
nand U22527 (N_22527,N_22271,N_22464);
nor U22528 (N_22528,N_22015,N_22445);
xnor U22529 (N_22529,N_22192,N_22488);
nor U22530 (N_22530,N_22120,N_22281);
nor U22531 (N_22531,N_22448,N_22358);
xnor U22532 (N_22532,N_22453,N_22329);
or U22533 (N_22533,N_22047,N_22347);
nor U22534 (N_22534,N_22389,N_22150);
nor U22535 (N_22535,N_22171,N_22143);
or U22536 (N_22536,N_22041,N_22422);
xor U22537 (N_22537,N_22002,N_22424);
and U22538 (N_22538,N_22209,N_22175);
nor U22539 (N_22539,N_22026,N_22418);
and U22540 (N_22540,N_22349,N_22460);
nor U22541 (N_22541,N_22251,N_22478);
xor U22542 (N_22542,N_22482,N_22331);
and U22543 (N_22543,N_22130,N_22343);
nand U22544 (N_22544,N_22223,N_22303);
and U22545 (N_22545,N_22403,N_22327);
or U22546 (N_22546,N_22212,N_22391);
nand U22547 (N_22547,N_22454,N_22146);
and U22548 (N_22548,N_22012,N_22363);
xnor U22549 (N_22549,N_22057,N_22361);
xnor U22550 (N_22550,N_22390,N_22011);
and U22551 (N_22551,N_22449,N_22492);
nor U22552 (N_22552,N_22293,N_22081);
or U22553 (N_22553,N_22246,N_22362);
nor U22554 (N_22554,N_22401,N_22082);
nand U22555 (N_22555,N_22240,N_22063);
nor U22556 (N_22556,N_22191,N_22396);
nor U22557 (N_22557,N_22180,N_22466);
nor U22558 (N_22558,N_22089,N_22360);
xnor U22559 (N_22559,N_22415,N_22122);
or U22560 (N_22560,N_22379,N_22119);
or U22561 (N_22561,N_22094,N_22165);
nor U22562 (N_22562,N_22006,N_22018);
nand U22563 (N_22563,N_22257,N_22097);
and U22564 (N_22564,N_22138,N_22469);
or U22565 (N_22565,N_22214,N_22436);
xnor U22566 (N_22566,N_22128,N_22357);
and U22567 (N_22567,N_22157,N_22463);
xnor U22568 (N_22568,N_22050,N_22008);
nand U22569 (N_22569,N_22326,N_22364);
nor U22570 (N_22570,N_22306,N_22105);
nand U22571 (N_22571,N_22004,N_22486);
nor U22572 (N_22572,N_22092,N_22052);
nor U22573 (N_22573,N_22049,N_22059);
nor U22574 (N_22574,N_22423,N_22172);
nor U22575 (N_22575,N_22406,N_22383);
nor U22576 (N_22576,N_22369,N_22295);
nor U22577 (N_22577,N_22099,N_22187);
nand U22578 (N_22578,N_22046,N_22048);
or U22579 (N_22579,N_22056,N_22498);
xor U22580 (N_22580,N_22493,N_22345);
nor U22581 (N_22581,N_22176,N_22330);
or U22582 (N_22582,N_22022,N_22410);
nor U22583 (N_22583,N_22136,N_22237);
or U22584 (N_22584,N_22499,N_22407);
and U22585 (N_22585,N_22074,N_22262);
xnor U22586 (N_22586,N_22434,N_22038);
nor U22587 (N_22587,N_22444,N_22433);
nor U22588 (N_22588,N_22351,N_22430);
and U22589 (N_22589,N_22164,N_22374);
nor U22590 (N_22590,N_22426,N_22005);
nand U22591 (N_22591,N_22141,N_22083);
nand U22592 (N_22592,N_22199,N_22416);
xor U22593 (N_22593,N_22166,N_22114);
or U22594 (N_22594,N_22053,N_22322);
or U22595 (N_22595,N_22121,N_22071);
and U22596 (N_22596,N_22243,N_22162);
xor U22597 (N_22597,N_22023,N_22098);
or U22598 (N_22598,N_22113,N_22373);
and U22599 (N_22599,N_22211,N_22051);
xor U22600 (N_22600,N_22093,N_22442);
nand U22601 (N_22601,N_22332,N_22135);
nand U22602 (N_22602,N_22102,N_22394);
nand U22603 (N_22603,N_22129,N_22446);
and U22604 (N_22604,N_22288,N_22266);
nor U22605 (N_22605,N_22481,N_22242);
nor U22606 (N_22606,N_22179,N_22276);
nor U22607 (N_22607,N_22380,N_22202);
and U22608 (N_22608,N_22473,N_22208);
and U22609 (N_22609,N_22066,N_22142);
nor U22610 (N_22610,N_22069,N_22215);
nor U22611 (N_22611,N_22145,N_22241);
nand U22612 (N_22612,N_22205,N_22387);
nor U22613 (N_22613,N_22117,N_22341);
nand U22614 (N_22614,N_22404,N_22402);
nand U22615 (N_22615,N_22457,N_22080);
or U22616 (N_22616,N_22297,N_22178);
or U22617 (N_22617,N_22118,N_22021);
nor U22618 (N_22618,N_22163,N_22299);
or U22619 (N_22619,N_22067,N_22054);
nor U22620 (N_22620,N_22148,N_22042);
nor U22621 (N_22621,N_22252,N_22304);
nor U22622 (N_22622,N_22203,N_22147);
or U22623 (N_22623,N_22123,N_22384);
nor U22624 (N_22624,N_22044,N_22480);
xnor U22625 (N_22625,N_22452,N_22441);
nand U22626 (N_22626,N_22393,N_22070);
and U22627 (N_22627,N_22370,N_22278);
xor U22628 (N_22628,N_22438,N_22078);
or U22629 (N_22629,N_22133,N_22095);
and U22630 (N_22630,N_22344,N_22253);
nand U22631 (N_22631,N_22279,N_22206);
nand U22632 (N_22632,N_22381,N_22264);
or U22633 (N_22633,N_22076,N_22334);
and U22634 (N_22634,N_22000,N_22222);
nor U22635 (N_22635,N_22079,N_22174);
and U22636 (N_22636,N_22200,N_22367);
or U22637 (N_22637,N_22375,N_22149);
and U22638 (N_22638,N_22058,N_22437);
or U22639 (N_22639,N_22116,N_22159);
nand U22640 (N_22640,N_22072,N_22219);
nand U22641 (N_22641,N_22489,N_22151);
nor U22642 (N_22642,N_22035,N_22198);
nor U22643 (N_22643,N_22096,N_22496);
nor U22644 (N_22644,N_22397,N_22236);
and U22645 (N_22645,N_22350,N_22227);
nand U22646 (N_22646,N_22186,N_22377);
nand U22647 (N_22647,N_22405,N_22110);
and U22648 (N_22648,N_22030,N_22112);
or U22649 (N_22649,N_22273,N_22465);
and U22650 (N_22650,N_22291,N_22213);
xor U22651 (N_22651,N_22106,N_22115);
nand U22652 (N_22652,N_22090,N_22353);
nor U22653 (N_22653,N_22016,N_22470);
or U22654 (N_22654,N_22491,N_22232);
xnor U22655 (N_22655,N_22024,N_22472);
nor U22656 (N_22656,N_22274,N_22310);
and U22657 (N_22657,N_22314,N_22001);
xnor U22658 (N_22658,N_22184,N_22443);
or U22659 (N_22659,N_22263,N_22247);
xnor U22660 (N_22660,N_22075,N_22085);
xor U22661 (N_22661,N_22400,N_22318);
or U22662 (N_22662,N_22368,N_22101);
xor U22663 (N_22663,N_22061,N_22140);
xor U22664 (N_22664,N_22007,N_22086);
xor U22665 (N_22665,N_22169,N_22037);
or U22666 (N_22666,N_22289,N_22156);
or U22667 (N_22667,N_22250,N_22027);
nor U22668 (N_22668,N_22336,N_22342);
or U22669 (N_22669,N_22338,N_22307);
nor U22670 (N_22670,N_22055,N_22183);
and U22671 (N_22671,N_22439,N_22131);
xor U22672 (N_22672,N_22248,N_22019);
nor U22673 (N_22673,N_22154,N_22152);
and U22674 (N_22674,N_22272,N_22296);
xor U22675 (N_22675,N_22195,N_22160);
or U22676 (N_22676,N_22077,N_22267);
xnor U22677 (N_22677,N_22408,N_22366);
nor U22678 (N_22678,N_22494,N_22233);
or U22679 (N_22679,N_22432,N_22003);
nand U22680 (N_22680,N_22062,N_22483);
or U22681 (N_22681,N_22204,N_22034);
xor U22682 (N_22682,N_22125,N_22309);
nand U22683 (N_22683,N_22170,N_22376);
nand U22684 (N_22684,N_22325,N_22268);
and U22685 (N_22685,N_22039,N_22447);
and U22686 (N_22686,N_22285,N_22217);
nand U22687 (N_22687,N_22259,N_22280);
and U22688 (N_22688,N_22025,N_22385);
nor U22689 (N_22689,N_22462,N_22287);
nor U22690 (N_22690,N_22300,N_22340);
and U22691 (N_22691,N_22261,N_22249);
nor U22692 (N_22692,N_22319,N_22188);
nand U22693 (N_22693,N_22283,N_22254);
and U22694 (N_22694,N_22398,N_22104);
or U22695 (N_22695,N_22036,N_22108);
or U22696 (N_22696,N_22239,N_22010);
and U22697 (N_22697,N_22155,N_22124);
and U22698 (N_22698,N_22238,N_22064);
nand U22699 (N_22699,N_22305,N_22429);
or U22700 (N_22700,N_22365,N_22256);
xnor U22701 (N_22701,N_22277,N_22456);
nor U22702 (N_22702,N_22269,N_22218);
and U22703 (N_22703,N_22193,N_22068);
and U22704 (N_22704,N_22235,N_22371);
nor U22705 (N_22705,N_22088,N_22458);
nor U22706 (N_22706,N_22348,N_22298);
nand U22707 (N_22707,N_22487,N_22476);
and U22708 (N_22708,N_22100,N_22490);
or U22709 (N_22709,N_22107,N_22103);
and U22710 (N_22710,N_22226,N_22177);
and U22711 (N_22711,N_22346,N_22033);
xor U22712 (N_22712,N_22013,N_22284);
nor U22713 (N_22713,N_22323,N_22221);
and U22714 (N_22714,N_22421,N_22290);
nand U22715 (N_22715,N_22139,N_22201);
xnor U22716 (N_22716,N_22312,N_22477);
or U22717 (N_22717,N_22065,N_22459);
xnor U22718 (N_22718,N_22431,N_22386);
nor U22719 (N_22719,N_22173,N_22210);
xor U22720 (N_22720,N_22395,N_22014);
nand U22721 (N_22721,N_22230,N_22427);
and U22722 (N_22722,N_22161,N_22412);
nor U22723 (N_22723,N_22153,N_22185);
nand U22724 (N_22724,N_22216,N_22378);
xnor U22725 (N_22725,N_22392,N_22029);
xnor U22726 (N_22726,N_22196,N_22286);
nand U22727 (N_22727,N_22244,N_22468);
xor U22728 (N_22728,N_22084,N_22265);
nand U22729 (N_22729,N_22417,N_22194);
xnor U22730 (N_22730,N_22419,N_22060);
or U22731 (N_22731,N_22471,N_22440);
or U22732 (N_22732,N_22197,N_22461);
and U22733 (N_22733,N_22311,N_22182);
or U22734 (N_22734,N_22317,N_22302);
xor U22735 (N_22735,N_22091,N_22245);
or U22736 (N_22736,N_22413,N_22255);
or U22737 (N_22737,N_22258,N_22354);
or U22738 (N_22738,N_22485,N_22409);
or U22739 (N_22739,N_22388,N_22132);
xor U22740 (N_22740,N_22372,N_22455);
nor U22741 (N_22741,N_22189,N_22313);
nor U22742 (N_22742,N_22224,N_22220);
xor U22743 (N_22743,N_22134,N_22127);
xor U22744 (N_22744,N_22158,N_22031);
and U22745 (N_22745,N_22228,N_22207);
nor U22746 (N_22746,N_22137,N_22382);
nor U22747 (N_22747,N_22260,N_22109);
and U22748 (N_22748,N_22294,N_22073);
or U22749 (N_22749,N_22190,N_22450);
and U22750 (N_22750,N_22348,N_22274);
and U22751 (N_22751,N_22181,N_22340);
nor U22752 (N_22752,N_22417,N_22424);
nand U22753 (N_22753,N_22098,N_22430);
nor U22754 (N_22754,N_22439,N_22327);
nand U22755 (N_22755,N_22291,N_22060);
or U22756 (N_22756,N_22200,N_22142);
nand U22757 (N_22757,N_22381,N_22241);
xnor U22758 (N_22758,N_22076,N_22385);
nand U22759 (N_22759,N_22389,N_22264);
or U22760 (N_22760,N_22171,N_22126);
nor U22761 (N_22761,N_22035,N_22169);
or U22762 (N_22762,N_22044,N_22237);
xnor U22763 (N_22763,N_22003,N_22228);
xnor U22764 (N_22764,N_22433,N_22398);
or U22765 (N_22765,N_22067,N_22349);
and U22766 (N_22766,N_22320,N_22175);
xor U22767 (N_22767,N_22127,N_22291);
xor U22768 (N_22768,N_22068,N_22301);
xor U22769 (N_22769,N_22279,N_22230);
nor U22770 (N_22770,N_22061,N_22097);
nor U22771 (N_22771,N_22287,N_22209);
nor U22772 (N_22772,N_22372,N_22365);
and U22773 (N_22773,N_22024,N_22276);
nand U22774 (N_22774,N_22123,N_22024);
xnor U22775 (N_22775,N_22359,N_22316);
nor U22776 (N_22776,N_22452,N_22258);
and U22777 (N_22777,N_22369,N_22055);
nand U22778 (N_22778,N_22432,N_22076);
or U22779 (N_22779,N_22206,N_22156);
xnor U22780 (N_22780,N_22135,N_22496);
nand U22781 (N_22781,N_22194,N_22242);
xor U22782 (N_22782,N_22302,N_22036);
nand U22783 (N_22783,N_22140,N_22190);
nor U22784 (N_22784,N_22156,N_22371);
nand U22785 (N_22785,N_22415,N_22375);
and U22786 (N_22786,N_22205,N_22046);
and U22787 (N_22787,N_22229,N_22094);
nor U22788 (N_22788,N_22103,N_22454);
nor U22789 (N_22789,N_22475,N_22044);
or U22790 (N_22790,N_22017,N_22205);
nand U22791 (N_22791,N_22314,N_22147);
xor U22792 (N_22792,N_22316,N_22477);
xor U22793 (N_22793,N_22366,N_22193);
or U22794 (N_22794,N_22490,N_22073);
xnor U22795 (N_22795,N_22471,N_22114);
xor U22796 (N_22796,N_22130,N_22011);
or U22797 (N_22797,N_22138,N_22460);
nor U22798 (N_22798,N_22356,N_22234);
nor U22799 (N_22799,N_22277,N_22268);
nand U22800 (N_22800,N_22320,N_22447);
and U22801 (N_22801,N_22063,N_22395);
nor U22802 (N_22802,N_22391,N_22489);
xor U22803 (N_22803,N_22372,N_22461);
nand U22804 (N_22804,N_22111,N_22342);
or U22805 (N_22805,N_22281,N_22475);
xor U22806 (N_22806,N_22488,N_22402);
and U22807 (N_22807,N_22468,N_22156);
or U22808 (N_22808,N_22156,N_22062);
xor U22809 (N_22809,N_22215,N_22402);
or U22810 (N_22810,N_22049,N_22433);
nor U22811 (N_22811,N_22470,N_22121);
or U22812 (N_22812,N_22190,N_22191);
or U22813 (N_22813,N_22012,N_22199);
and U22814 (N_22814,N_22365,N_22427);
and U22815 (N_22815,N_22232,N_22151);
and U22816 (N_22816,N_22489,N_22185);
nand U22817 (N_22817,N_22114,N_22081);
and U22818 (N_22818,N_22314,N_22326);
and U22819 (N_22819,N_22378,N_22082);
nor U22820 (N_22820,N_22384,N_22197);
or U22821 (N_22821,N_22236,N_22405);
nor U22822 (N_22822,N_22395,N_22083);
xnor U22823 (N_22823,N_22034,N_22320);
nand U22824 (N_22824,N_22180,N_22240);
or U22825 (N_22825,N_22404,N_22370);
or U22826 (N_22826,N_22175,N_22084);
nor U22827 (N_22827,N_22321,N_22136);
nand U22828 (N_22828,N_22136,N_22171);
nor U22829 (N_22829,N_22296,N_22181);
nand U22830 (N_22830,N_22097,N_22423);
xnor U22831 (N_22831,N_22323,N_22137);
and U22832 (N_22832,N_22170,N_22065);
or U22833 (N_22833,N_22268,N_22353);
and U22834 (N_22834,N_22324,N_22337);
nand U22835 (N_22835,N_22081,N_22046);
nand U22836 (N_22836,N_22300,N_22073);
xor U22837 (N_22837,N_22343,N_22229);
xor U22838 (N_22838,N_22470,N_22246);
or U22839 (N_22839,N_22055,N_22445);
nand U22840 (N_22840,N_22305,N_22434);
xnor U22841 (N_22841,N_22170,N_22438);
nand U22842 (N_22842,N_22122,N_22053);
xor U22843 (N_22843,N_22392,N_22475);
nand U22844 (N_22844,N_22274,N_22152);
and U22845 (N_22845,N_22261,N_22499);
or U22846 (N_22846,N_22040,N_22235);
and U22847 (N_22847,N_22182,N_22332);
nand U22848 (N_22848,N_22436,N_22119);
and U22849 (N_22849,N_22031,N_22100);
or U22850 (N_22850,N_22461,N_22070);
nand U22851 (N_22851,N_22338,N_22248);
nand U22852 (N_22852,N_22476,N_22478);
xnor U22853 (N_22853,N_22333,N_22247);
and U22854 (N_22854,N_22495,N_22286);
or U22855 (N_22855,N_22075,N_22359);
xnor U22856 (N_22856,N_22428,N_22078);
or U22857 (N_22857,N_22187,N_22373);
nor U22858 (N_22858,N_22179,N_22378);
xnor U22859 (N_22859,N_22101,N_22402);
or U22860 (N_22860,N_22345,N_22020);
or U22861 (N_22861,N_22083,N_22058);
nor U22862 (N_22862,N_22399,N_22393);
nor U22863 (N_22863,N_22370,N_22319);
xor U22864 (N_22864,N_22405,N_22123);
xnor U22865 (N_22865,N_22265,N_22108);
nor U22866 (N_22866,N_22349,N_22384);
xnor U22867 (N_22867,N_22320,N_22424);
and U22868 (N_22868,N_22140,N_22413);
nand U22869 (N_22869,N_22115,N_22183);
or U22870 (N_22870,N_22148,N_22473);
nand U22871 (N_22871,N_22336,N_22322);
nor U22872 (N_22872,N_22102,N_22135);
xor U22873 (N_22873,N_22081,N_22232);
nor U22874 (N_22874,N_22044,N_22029);
xnor U22875 (N_22875,N_22356,N_22165);
xnor U22876 (N_22876,N_22115,N_22464);
nand U22877 (N_22877,N_22159,N_22373);
nor U22878 (N_22878,N_22337,N_22325);
and U22879 (N_22879,N_22092,N_22412);
xor U22880 (N_22880,N_22340,N_22151);
nand U22881 (N_22881,N_22416,N_22387);
and U22882 (N_22882,N_22110,N_22440);
or U22883 (N_22883,N_22183,N_22305);
nand U22884 (N_22884,N_22405,N_22381);
and U22885 (N_22885,N_22191,N_22017);
or U22886 (N_22886,N_22058,N_22319);
xor U22887 (N_22887,N_22441,N_22338);
or U22888 (N_22888,N_22077,N_22446);
nor U22889 (N_22889,N_22186,N_22376);
xnor U22890 (N_22890,N_22050,N_22213);
and U22891 (N_22891,N_22237,N_22117);
and U22892 (N_22892,N_22435,N_22380);
nand U22893 (N_22893,N_22152,N_22391);
and U22894 (N_22894,N_22300,N_22145);
or U22895 (N_22895,N_22046,N_22294);
xor U22896 (N_22896,N_22470,N_22430);
and U22897 (N_22897,N_22233,N_22462);
nor U22898 (N_22898,N_22133,N_22344);
nor U22899 (N_22899,N_22090,N_22451);
nand U22900 (N_22900,N_22084,N_22017);
xor U22901 (N_22901,N_22367,N_22346);
or U22902 (N_22902,N_22297,N_22137);
and U22903 (N_22903,N_22044,N_22469);
nor U22904 (N_22904,N_22174,N_22186);
or U22905 (N_22905,N_22203,N_22291);
xnor U22906 (N_22906,N_22490,N_22422);
or U22907 (N_22907,N_22221,N_22448);
or U22908 (N_22908,N_22375,N_22234);
and U22909 (N_22909,N_22035,N_22155);
or U22910 (N_22910,N_22408,N_22057);
or U22911 (N_22911,N_22088,N_22382);
xor U22912 (N_22912,N_22046,N_22304);
xor U22913 (N_22913,N_22453,N_22228);
and U22914 (N_22914,N_22054,N_22031);
nor U22915 (N_22915,N_22065,N_22253);
or U22916 (N_22916,N_22444,N_22313);
or U22917 (N_22917,N_22220,N_22454);
and U22918 (N_22918,N_22016,N_22300);
nand U22919 (N_22919,N_22350,N_22283);
or U22920 (N_22920,N_22164,N_22308);
or U22921 (N_22921,N_22450,N_22055);
and U22922 (N_22922,N_22171,N_22167);
and U22923 (N_22923,N_22395,N_22293);
xor U22924 (N_22924,N_22276,N_22270);
nor U22925 (N_22925,N_22315,N_22341);
nor U22926 (N_22926,N_22438,N_22008);
and U22927 (N_22927,N_22480,N_22122);
xnor U22928 (N_22928,N_22279,N_22281);
nand U22929 (N_22929,N_22211,N_22084);
nand U22930 (N_22930,N_22156,N_22405);
and U22931 (N_22931,N_22013,N_22396);
xnor U22932 (N_22932,N_22464,N_22368);
nor U22933 (N_22933,N_22382,N_22139);
xor U22934 (N_22934,N_22054,N_22244);
and U22935 (N_22935,N_22463,N_22256);
xor U22936 (N_22936,N_22382,N_22006);
nor U22937 (N_22937,N_22295,N_22185);
or U22938 (N_22938,N_22381,N_22131);
and U22939 (N_22939,N_22427,N_22048);
xor U22940 (N_22940,N_22253,N_22322);
xnor U22941 (N_22941,N_22214,N_22493);
and U22942 (N_22942,N_22130,N_22031);
xor U22943 (N_22943,N_22157,N_22032);
nor U22944 (N_22944,N_22407,N_22477);
xnor U22945 (N_22945,N_22271,N_22036);
xor U22946 (N_22946,N_22350,N_22183);
or U22947 (N_22947,N_22015,N_22297);
nand U22948 (N_22948,N_22155,N_22021);
nand U22949 (N_22949,N_22051,N_22015);
xnor U22950 (N_22950,N_22241,N_22390);
and U22951 (N_22951,N_22299,N_22222);
nand U22952 (N_22952,N_22418,N_22324);
xor U22953 (N_22953,N_22443,N_22058);
nand U22954 (N_22954,N_22380,N_22308);
nor U22955 (N_22955,N_22278,N_22254);
or U22956 (N_22956,N_22001,N_22213);
or U22957 (N_22957,N_22032,N_22347);
or U22958 (N_22958,N_22101,N_22184);
and U22959 (N_22959,N_22190,N_22436);
or U22960 (N_22960,N_22368,N_22426);
nand U22961 (N_22961,N_22349,N_22097);
xnor U22962 (N_22962,N_22368,N_22261);
nor U22963 (N_22963,N_22189,N_22167);
nor U22964 (N_22964,N_22432,N_22162);
nand U22965 (N_22965,N_22137,N_22443);
and U22966 (N_22966,N_22346,N_22152);
and U22967 (N_22967,N_22263,N_22357);
nor U22968 (N_22968,N_22307,N_22457);
nor U22969 (N_22969,N_22466,N_22173);
nor U22970 (N_22970,N_22094,N_22402);
nor U22971 (N_22971,N_22386,N_22024);
nand U22972 (N_22972,N_22249,N_22089);
and U22973 (N_22973,N_22129,N_22153);
xnor U22974 (N_22974,N_22224,N_22168);
nand U22975 (N_22975,N_22147,N_22122);
nand U22976 (N_22976,N_22015,N_22196);
xnor U22977 (N_22977,N_22260,N_22073);
xor U22978 (N_22978,N_22429,N_22302);
nor U22979 (N_22979,N_22029,N_22322);
nor U22980 (N_22980,N_22036,N_22466);
xnor U22981 (N_22981,N_22301,N_22306);
nor U22982 (N_22982,N_22291,N_22087);
nor U22983 (N_22983,N_22482,N_22188);
xnor U22984 (N_22984,N_22162,N_22345);
nor U22985 (N_22985,N_22066,N_22289);
xnor U22986 (N_22986,N_22230,N_22070);
nand U22987 (N_22987,N_22452,N_22159);
nand U22988 (N_22988,N_22308,N_22498);
nor U22989 (N_22989,N_22195,N_22369);
and U22990 (N_22990,N_22116,N_22080);
or U22991 (N_22991,N_22147,N_22188);
and U22992 (N_22992,N_22077,N_22202);
nor U22993 (N_22993,N_22301,N_22333);
nand U22994 (N_22994,N_22312,N_22373);
nand U22995 (N_22995,N_22465,N_22198);
and U22996 (N_22996,N_22243,N_22351);
nor U22997 (N_22997,N_22378,N_22115);
nand U22998 (N_22998,N_22180,N_22001);
or U22999 (N_22999,N_22433,N_22285);
and U23000 (N_23000,N_22981,N_22855);
and U23001 (N_23001,N_22669,N_22723);
nand U23002 (N_23002,N_22829,N_22963);
xnor U23003 (N_23003,N_22954,N_22635);
xnor U23004 (N_23004,N_22557,N_22757);
nand U23005 (N_23005,N_22961,N_22902);
or U23006 (N_23006,N_22565,N_22741);
and U23007 (N_23007,N_22819,N_22670);
nor U23008 (N_23008,N_22554,N_22850);
nor U23009 (N_23009,N_22684,N_22648);
and U23010 (N_23010,N_22754,N_22881);
nor U23011 (N_23011,N_22841,N_22664);
and U23012 (N_23012,N_22667,N_22620);
nor U23013 (N_23013,N_22939,N_22671);
and U23014 (N_23014,N_22947,N_22592);
nor U23015 (N_23015,N_22583,N_22748);
nand U23016 (N_23016,N_22692,N_22873);
nand U23017 (N_23017,N_22584,N_22807);
nor U23018 (N_23018,N_22722,N_22562);
and U23019 (N_23019,N_22724,N_22989);
xor U23020 (N_23020,N_22573,N_22643);
or U23021 (N_23021,N_22708,N_22677);
nor U23022 (N_23022,N_22623,N_22535);
nand U23023 (N_23023,N_22742,N_22517);
or U23024 (N_23024,N_22884,N_22816);
and U23025 (N_23025,N_22637,N_22531);
nor U23026 (N_23026,N_22998,N_22822);
nor U23027 (N_23027,N_22821,N_22857);
xor U23028 (N_23028,N_22879,N_22705);
or U23029 (N_23029,N_22529,N_22906);
nor U23030 (N_23030,N_22527,N_22701);
nand U23031 (N_23031,N_22752,N_22540);
or U23032 (N_23032,N_22749,N_22525);
and U23033 (N_23033,N_22979,N_22951);
xor U23034 (N_23034,N_22642,N_22733);
nor U23035 (N_23035,N_22628,N_22851);
or U23036 (N_23036,N_22513,N_22767);
nor U23037 (N_23037,N_22911,N_22546);
nor U23038 (N_23038,N_22520,N_22831);
and U23039 (N_23039,N_22710,N_22920);
or U23040 (N_23040,N_22703,N_22820);
nor U23041 (N_23041,N_22709,N_22652);
nor U23042 (N_23042,N_22927,N_22561);
and U23043 (N_23043,N_22836,N_22697);
or U23044 (N_23044,N_22766,N_22897);
nor U23045 (N_23045,N_22958,N_22594);
and U23046 (N_23046,N_22859,N_22765);
nand U23047 (N_23047,N_22899,N_22640);
nand U23048 (N_23048,N_22999,N_22952);
or U23049 (N_23049,N_22833,N_22704);
and U23050 (N_23050,N_22559,N_22673);
nand U23051 (N_23051,N_22725,N_22691);
and U23052 (N_23052,N_22633,N_22696);
or U23053 (N_23053,N_22843,N_22794);
xnor U23054 (N_23054,N_22802,N_22895);
nand U23055 (N_23055,N_22904,N_22746);
xnor U23056 (N_23056,N_22738,N_22894);
nor U23057 (N_23057,N_22657,N_22682);
nor U23058 (N_23058,N_22966,N_22950);
xnor U23059 (N_23059,N_22854,N_22801);
nor U23060 (N_23060,N_22615,N_22686);
nor U23061 (N_23061,N_22534,N_22867);
and U23062 (N_23062,N_22891,N_22949);
nand U23063 (N_23063,N_22676,N_22711);
nor U23064 (N_23064,N_22769,N_22695);
nor U23065 (N_23065,N_22607,N_22515);
or U23066 (N_23066,N_22755,N_22905);
xor U23067 (N_23067,N_22878,N_22988);
xor U23068 (N_23068,N_22683,N_22768);
and U23069 (N_23069,N_22666,N_22982);
or U23070 (N_23070,N_22996,N_22596);
and U23071 (N_23071,N_22539,N_22645);
nand U23072 (N_23072,N_22886,N_22872);
xnor U23073 (N_23073,N_22582,N_22609);
xnor U23074 (N_23074,N_22991,N_22564);
nand U23075 (N_23075,N_22617,N_22745);
nand U23076 (N_23076,N_22660,N_22903);
nor U23077 (N_23077,N_22842,N_22522);
or U23078 (N_23078,N_22800,N_22786);
nor U23079 (N_23079,N_22882,N_22856);
or U23080 (N_23080,N_22980,N_22861);
nor U23081 (N_23081,N_22658,N_22622);
nand U23082 (N_23082,N_22681,N_22654);
nand U23083 (N_23083,N_22913,N_22824);
or U23084 (N_23084,N_22880,N_22675);
and U23085 (N_23085,N_22608,N_22524);
nand U23086 (N_23086,N_22544,N_22885);
and U23087 (N_23087,N_22629,N_22672);
xnor U23088 (N_23088,N_22805,N_22751);
and U23089 (N_23089,N_22631,N_22835);
or U23090 (N_23090,N_22776,N_22919);
or U23091 (N_23091,N_22815,N_22661);
xor U23092 (N_23092,N_22953,N_22781);
nor U23093 (N_23093,N_22555,N_22814);
nor U23094 (N_23094,N_22638,N_22809);
and U23095 (N_23095,N_22803,N_22685);
or U23096 (N_23096,N_22591,N_22799);
and U23097 (N_23097,N_22750,N_22798);
nor U23098 (N_23098,N_22504,N_22931);
or U23099 (N_23099,N_22945,N_22616);
nor U23100 (N_23100,N_22598,N_22626);
nor U23101 (N_23101,N_22533,N_22992);
xnor U23102 (N_23102,N_22610,N_22795);
xnor U23103 (N_23103,N_22714,N_22727);
xor U23104 (N_23104,N_22864,N_22699);
and U23105 (N_23105,N_22811,N_22706);
or U23106 (N_23106,N_22972,N_22852);
xor U23107 (N_23107,N_22935,N_22656);
or U23108 (N_23108,N_22712,N_22888);
nand U23109 (N_23109,N_22926,N_22687);
nor U23110 (N_23110,N_22537,N_22790);
or U23111 (N_23111,N_22505,N_22521);
or U23112 (N_23112,N_22550,N_22896);
xnor U23113 (N_23113,N_22764,N_22924);
nor U23114 (N_23114,N_22621,N_22548);
and U23115 (N_23115,N_22647,N_22853);
xnor U23116 (N_23116,N_22509,N_22698);
xnor U23117 (N_23117,N_22516,N_22977);
or U23118 (N_23118,N_22823,N_22870);
or U23119 (N_23119,N_22759,N_22624);
and U23120 (N_23120,N_22736,N_22549);
nor U23121 (N_23121,N_22933,N_22665);
nor U23122 (N_23122,N_22523,N_22506);
or U23123 (N_23123,N_22744,N_22789);
and U23124 (N_23124,N_22575,N_22965);
and U23125 (N_23125,N_22921,N_22530);
and U23126 (N_23126,N_22985,N_22619);
xor U23127 (N_23127,N_22604,N_22946);
and U23128 (N_23128,N_22663,N_22838);
nor U23129 (N_23129,N_22840,N_22653);
xnor U23130 (N_23130,N_22874,N_22804);
or U23131 (N_23131,N_22783,N_22987);
nor U23132 (N_23132,N_22556,N_22693);
or U23133 (N_23133,N_22956,N_22860);
nor U23134 (N_23134,N_22625,N_22892);
or U23135 (N_23135,N_22595,N_22875);
nand U23136 (N_23136,N_22771,N_22578);
nand U23137 (N_23137,N_22553,N_22649);
nor U23138 (N_23138,N_22883,N_22552);
and U23139 (N_23139,N_22818,N_22732);
and U23140 (N_23140,N_22922,N_22545);
xor U23141 (N_23141,N_22974,N_22646);
nor U23142 (N_23142,N_22774,N_22679);
and U23143 (N_23143,N_22651,N_22779);
or U23144 (N_23144,N_22976,N_22576);
and U23145 (N_23145,N_22957,N_22585);
nor U23146 (N_23146,N_22700,N_22993);
xor U23147 (N_23147,N_22541,N_22969);
xnor U23148 (N_23148,N_22678,N_22973);
nand U23149 (N_23149,N_22930,N_22934);
nand U23150 (N_23150,N_22632,N_22887);
nor U23151 (N_23151,N_22532,N_22612);
and U23152 (N_23152,N_22659,N_22674);
nor U23153 (N_23153,N_22758,N_22680);
xor U23154 (N_23154,N_22918,N_22928);
xor U23155 (N_23155,N_22605,N_22740);
or U23156 (N_23156,N_22502,N_22940);
nor U23157 (N_23157,N_22917,N_22611);
or U23158 (N_23158,N_22941,N_22915);
or U23159 (N_23159,N_22890,N_22731);
and U23160 (N_23160,N_22760,N_22912);
nor U23161 (N_23161,N_22586,N_22830);
nor U23162 (N_23162,N_22826,N_22580);
nand U23163 (N_23163,N_22787,N_22606);
nor U23164 (N_23164,N_22871,N_22542);
xor U23165 (N_23165,N_22501,N_22813);
and U23166 (N_23166,N_22869,N_22782);
nor U23167 (N_23167,N_22603,N_22942);
nand U23168 (N_23168,N_22845,N_22694);
nand U23169 (N_23169,N_22964,N_22551);
nand U23170 (N_23170,N_22614,N_22572);
or U23171 (N_23171,N_22716,N_22908);
xor U23172 (N_23172,N_22717,N_22762);
xor U23173 (N_23173,N_22512,N_22500);
or U23174 (N_23174,N_22863,N_22778);
nand U23175 (N_23175,N_22916,N_22932);
and U23176 (N_23176,N_22719,N_22994);
nand U23177 (N_23177,N_22948,N_22901);
or U23178 (N_23178,N_22862,N_22876);
or U23179 (N_23179,N_22655,N_22644);
and U23180 (N_23180,N_22567,N_22574);
nor U23181 (N_23181,N_22579,N_22599);
xnor U23182 (N_23182,N_22866,N_22514);
xor U23183 (N_23183,N_22547,N_22909);
xnor U23184 (N_23184,N_22846,N_22936);
or U23185 (N_23185,N_22662,N_22689);
nand U23186 (N_23186,N_22560,N_22832);
xor U23187 (N_23187,N_22770,N_22914);
nand U23188 (N_23188,N_22898,N_22721);
nand U23189 (N_23189,N_22639,N_22600);
nor U23190 (N_23190,N_22508,N_22877);
nor U23191 (N_23191,N_22588,N_22923);
or U23192 (N_23192,N_22938,N_22713);
nand U23193 (N_23193,N_22827,N_22907);
and U23194 (N_23194,N_22737,N_22518);
and U23195 (N_23195,N_22808,N_22970);
xnor U23196 (N_23196,N_22739,N_22849);
xor U23197 (N_23197,N_22590,N_22817);
nor U23198 (N_23198,N_22943,N_22785);
nor U23199 (N_23199,N_22761,N_22568);
nand U23200 (N_23200,N_22865,N_22889);
and U23201 (N_23201,N_22601,N_22571);
or U23202 (N_23202,N_22702,N_22834);
and U23203 (N_23203,N_22806,N_22995);
nor U23204 (N_23204,N_22791,N_22847);
nand U23205 (N_23205,N_22636,N_22780);
nand U23206 (N_23206,N_22775,N_22944);
xnor U23207 (N_23207,N_22900,N_22597);
nor U23208 (N_23208,N_22975,N_22983);
and U23209 (N_23209,N_22510,N_22997);
nor U23210 (N_23210,N_22577,N_22718);
or U23211 (N_23211,N_22747,N_22569);
or U23212 (N_23212,N_22593,N_22587);
xor U23213 (N_23213,N_22627,N_22828);
and U23214 (N_23214,N_22613,N_22729);
nand U23215 (N_23215,N_22602,N_22986);
or U23216 (N_23216,N_22868,N_22893);
or U23217 (N_23217,N_22967,N_22570);
nor U23218 (N_23218,N_22796,N_22536);
xor U23219 (N_23219,N_22734,N_22797);
nor U23220 (N_23220,N_22962,N_22715);
xor U23221 (N_23221,N_22960,N_22990);
nor U23222 (N_23222,N_22507,N_22688);
xnor U23223 (N_23223,N_22641,N_22858);
nor U23224 (N_23224,N_22792,N_22763);
and U23225 (N_23225,N_22837,N_22735);
or U23226 (N_23226,N_22788,N_22753);
nor U23227 (N_23227,N_22558,N_22793);
nand U23228 (N_23228,N_22971,N_22925);
nand U23229 (N_23229,N_22563,N_22720);
xor U23230 (N_23230,N_22511,N_22929);
xor U23231 (N_23231,N_22618,N_22726);
xor U23232 (N_23232,N_22528,N_22756);
nor U23233 (N_23233,N_22959,N_22503);
nor U23234 (N_23234,N_22784,N_22812);
and U23235 (N_23235,N_22634,N_22650);
nand U23236 (N_23236,N_22844,N_22690);
and U23237 (N_23237,N_22538,N_22728);
nor U23238 (N_23238,N_22839,N_22707);
nor U23239 (N_23239,N_22743,N_22589);
xnor U23240 (N_23240,N_22968,N_22978);
and U23241 (N_23241,N_22955,N_22777);
nand U23242 (N_23242,N_22519,N_22937);
xor U23243 (N_23243,N_22910,N_22668);
xor U23244 (N_23244,N_22526,N_22630);
or U23245 (N_23245,N_22810,N_22566);
xor U23246 (N_23246,N_22543,N_22730);
xor U23247 (N_23247,N_22984,N_22848);
and U23248 (N_23248,N_22773,N_22825);
xnor U23249 (N_23249,N_22772,N_22581);
nor U23250 (N_23250,N_22870,N_22664);
nand U23251 (N_23251,N_22860,N_22782);
xor U23252 (N_23252,N_22721,N_22790);
and U23253 (N_23253,N_22517,N_22751);
and U23254 (N_23254,N_22706,N_22748);
nor U23255 (N_23255,N_22777,N_22551);
nor U23256 (N_23256,N_22538,N_22610);
or U23257 (N_23257,N_22629,N_22992);
or U23258 (N_23258,N_22869,N_22969);
or U23259 (N_23259,N_22533,N_22902);
xnor U23260 (N_23260,N_22634,N_22864);
nor U23261 (N_23261,N_22665,N_22607);
and U23262 (N_23262,N_22932,N_22534);
or U23263 (N_23263,N_22601,N_22827);
nand U23264 (N_23264,N_22530,N_22953);
nand U23265 (N_23265,N_22517,N_22825);
nor U23266 (N_23266,N_22738,N_22727);
and U23267 (N_23267,N_22582,N_22905);
xor U23268 (N_23268,N_22627,N_22994);
or U23269 (N_23269,N_22852,N_22562);
or U23270 (N_23270,N_22994,N_22903);
nor U23271 (N_23271,N_22910,N_22581);
xor U23272 (N_23272,N_22786,N_22939);
nor U23273 (N_23273,N_22554,N_22896);
xnor U23274 (N_23274,N_22597,N_22982);
and U23275 (N_23275,N_22607,N_22706);
xor U23276 (N_23276,N_22550,N_22782);
xnor U23277 (N_23277,N_22847,N_22757);
nor U23278 (N_23278,N_22919,N_22559);
nor U23279 (N_23279,N_22816,N_22851);
or U23280 (N_23280,N_22887,N_22704);
nor U23281 (N_23281,N_22875,N_22715);
xnor U23282 (N_23282,N_22608,N_22583);
and U23283 (N_23283,N_22843,N_22531);
nor U23284 (N_23284,N_22554,N_22603);
nor U23285 (N_23285,N_22580,N_22965);
or U23286 (N_23286,N_22754,N_22736);
nor U23287 (N_23287,N_22967,N_22695);
nand U23288 (N_23288,N_22985,N_22668);
xnor U23289 (N_23289,N_22581,N_22734);
xnor U23290 (N_23290,N_22893,N_22858);
or U23291 (N_23291,N_22977,N_22996);
and U23292 (N_23292,N_22916,N_22701);
xor U23293 (N_23293,N_22628,N_22574);
nor U23294 (N_23294,N_22988,N_22941);
or U23295 (N_23295,N_22589,N_22981);
or U23296 (N_23296,N_22917,N_22720);
or U23297 (N_23297,N_22574,N_22661);
xor U23298 (N_23298,N_22746,N_22533);
nand U23299 (N_23299,N_22725,N_22899);
and U23300 (N_23300,N_22695,N_22990);
xnor U23301 (N_23301,N_22763,N_22817);
and U23302 (N_23302,N_22697,N_22745);
or U23303 (N_23303,N_22582,N_22830);
or U23304 (N_23304,N_22608,N_22622);
or U23305 (N_23305,N_22753,N_22726);
and U23306 (N_23306,N_22856,N_22567);
nor U23307 (N_23307,N_22732,N_22587);
nor U23308 (N_23308,N_22887,N_22615);
or U23309 (N_23309,N_22894,N_22509);
nor U23310 (N_23310,N_22661,N_22854);
xnor U23311 (N_23311,N_22856,N_22614);
xor U23312 (N_23312,N_22925,N_22539);
and U23313 (N_23313,N_22666,N_22898);
or U23314 (N_23314,N_22783,N_22668);
nand U23315 (N_23315,N_22564,N_22776);
nor U23316 (N_23316,N_22969,N_22993);
xnor U23317 (N_23317,N_22919,N_22520);
xor U23318 (N_23318,N_22774,N_22719);
and U23319 (N_23319,N_22956,N_22869);
nand U23320 (N_23320,N_22741,N_22626);
xnor U23321 (N_23321,N_22551,N_22967);
nor U23322 (N_23322,N_22920,N_22629);
and U23323 (N_23323,N_22825,N_22768);
nand U23324 (N_23324,N_22691,N_22687);
and U23325 (N_23325,N_22894,N_22821);
or U23326 (N_23326,N_22910,N_22796);
nand U23327 (N_23327,N_22866,N_22529);
and U23328 (N_23328,N_22597,N_22899);
nand U23329 (N_23329,N_22738,N_22715);
or U23330 (N_23330,N_22995,N_22602);
xor U23331 (N_23331,N_22842,N_22943);
nand U23332 (N_23332,N_22982,N_22862);
xor U23333 (N_23333,N_22765,N_22632);
nand U23334 (N_23334,N_22753,N_22759);
or U23335 (N_23335,N_22721,N_22863);
or U23336 (N_23336,N_22612,N_22784);
nand U23337 (N_23337,N_22761,N_22866);
and U23338 (N_23338,N_22714,N_22970);
or U23339 (N_23339,N_22874,N_22556);
xnor U23340 (N_23340,N_22891,N_22776);
xor U23341 (N_23341,N_22844,N_22899);
nand U23342 (N_23342,N_22615,N_22940);
and U23343 (N_23343,N_22712,N_22894);
nor U23344 (N_23344,N_22796,N_22906);
and U23345 (N_23345,N_22653,N_22786);
and U23346 (N_23346,N_22684,N_22996);
or U23347 (N_23347,N_22968,N_22522);
nand U23348 (N_23348,N_22617,N_22558);
nor U23349 (N_23349,N_22669,N_22738);
nand U23350 (N_23350,N_22781,N_22866);
and U23351 (N_23351,N_22929,N_22723);
nand U23352 (N_23352,N_22513,N_22764);
or U23353 (N_23353,N_22623,N_22788);
nor U23354 (N_23354,N_22865,N_22517);
nand U23355 (N_23355,N_22829,N_22803);
nor U23356 (N_23356,N_22809,N_22997);
or U23357 (N_23357,N_22584,N_22778);
nand U23358 (N_23358,N_22597,N_22845);
nor U23359 (N_23359,N_22967,N_22613);
nor U23360 (N_23360,N_22925,N_22749);
and U23361 (N_23361,N_22609,N_22563);
and U23362 (N_23362,N_22866,N_22856);
or U23363 (N_23363,N_22981,N_22678);
xnor U23364 (N_23364,N_22621,N_22501);
nor U23365 (N_23365,N_22799,N_22686);
or U23366 (N_23366,N_22557,N_22751);
nor U23367 (N_23367,N_22615,N_22595);
nor U23368 (N_23368,N_22976,N_22543);
nor U23369 (N_23369,N_22916,N_22986);
or U23370 (N_23370,N_22659,N_22731);
nor U23371 (N_23371,N_22659,N_22539);
and U23372 (N_23372,N_22575,N_22947);
and U23373 (N_23373,N_22531,N_22579);
nand U23374 (N_23374,N_22889,N_22746);
or U23375 (N_23375,N_22660,N_22965);
xnor U23376 (N_23376,N_22672,N_22873);
nand U23377 (N_23377,N_22994,N_22825);
nand U23378 (N_23378,N_22894,N_22936);
nand U23379 (N_23379,N_22566,N_22814);
nand U23380 (N_23380,N_22832,N_22984);
nand U23381 (N_23381,N_22609,N_22683);
or U23382 (N_23382,N_22608,N_22949);
and U23383 (N_23383,N_22863,N_22569);
and U23384 (N_23384,N_22869,N_22676);
and U23385 (N_23385,N_22977,N_22753);
or U23386 (N_23386,N_22706,N_22737);
and U23387 (N_23387,N_22662,N_22956);
nand U23388 (N_23388,N_22965,N_22781);
and U23389 (N_23389,N_22575,N_22903);
and U23390 (N_23390,N_22763,N_22585);
or U23391 (N_23391,N_22995,N_22781);
xor U23392 (N_23392,N_22823,N_22974);
nand U23393 (N_23393,N_22892,N_22728);
nand U23394 (N_23394,N_22608,N_22880);
xnor U23395 (N_23395,N_22759,N_22961);
xor U23396 (N_23396,N_22548,N_22830);
and U23397 (N_23397,N_22583,N_22772);
nand U23398 (N_23398,N_22904,N_22877);
xor U23399 (N_23399,N_22898,N_22665);
nand U23400 (N_23400,N_22789,N_22513);
xnor U23401 (N_23401,N_22587,N_22672);
or U23402 (N_23402,N_22671,N_22742);
nand U23403 (N_23403,N_22587,N_22934);
xor U23404 (N_23404,N_22508,N_22672);
and U23405 (N_23405,N_22924,N_22861);
xnor U23406 (N_23406,N_22801,N_22593);
or U23407 (N_23407,N_22885,N_22531);
nor U23408 (N_23408,N_22534,N_22704);
xnor U23409 (N_23409,N_22614,N_22995);
nand U23410 (N_23410,N_22595,N_22870);
xnor U23411 (N_23411,N_22939,N_22952);
xor U23412 (N_23412,N_22810,N_22816);
and U23413 (N_23413,N_22507,N_22727);
or U23414 (N_23414,N_22813,N_22957);
or U23415 (N_23415,N_22802,N_22644);
nand U23416 (N_23416,N_22606,N_22856);
and U23417 (N_23417,N_22814,N_22893);
nand U23418 (N_23418,N_22807,N_22687);
and U23419 (N_23419,N_22903,N_22901);
xor U23420 (N_23420,N_22542,N_22722);
nand U23421 (N_23421,N_22750,N_22504);
or U23422 (N_23422,N_22990,N_22624);
nand U23423 (N_23423,N_22850,N_22938);
xnor U23424 (N_23424,N_22628,N_22560);
and U23425 (N_23425,N_22676,N_22654);
or U23426 (N_23426,N_22708,N_22754);
or U23427 (N_23427,N_22517,N_22982);
and U23428 (N_23428,N_22844,N_22829);
nor U23429 (N_23429,N_22642,N_22615);
xnor U23430 (N_23430,N_22697,N_22744);
nand U23431 (N_23431,N_22621,N_22606);
or U23432 (N_23432,N_22883,N_22717);
or U23433 (N_23433,N_22930,N_22844);
nor U23434 (N_23434,N_22575,N_22644);
nand U23435 (N_23435,N_22697,N_22644);
nand U23436 (N_23436,N_22801,N_22617);
xnor U23437 (N_23437,N_22731,N_22866);
nand U23438 (N_23438,N_22574,N_22770);
xor U23439 (N_23439,N_22877,N_22651);
xnor U23440 (N_23440,N_22978,N_22650);
or U23441 (N_23441,N_22550,N_22676);
or U23442 (N_23442,N_22767,N_22644);
xnor U23443 (N_23443,N_22652,N_22900);
nand U23444 (N_23444,N_22605,N_22833);
or U23445 (N_23445,N_22516,N_22696);
nor U23446 (N_23446,N_22654,N_22510);
nand U23447 (N_23447,N_22991,N_22579);
xor U23448 (N_23448,N_22528,N_22630);
or U23449 (N_23449,N_22836,N_22958);
or U23450 (N_23450,N_22500,N_22733);
and U23451 (N_23451,N_22842,N_22783);
or U23452 (N_23452,N_22853,N_22544);
xor U23453 (N_23453,N_22555,N_22945);
xnor U23454 (N_23454,N_22776,N_22732);
nand U23455 (N_23455,N_22856,N_22505);
nor U23456 (N_23456,N_22534,N_22802);
nor U23457 (N_23457,N_22980,N_22529);
nand U23458 (N_23458,N_22897,N_22657);
or U23459 (N_23459,N_22857,N_22822);
and U23460 (N_23460,N_22805,N_22678);
nand U23461 (N_23461,N_22681,N_22695);
nor U23462 (N_23462,N_22834,N_22610);
nand U23463 (N_23463,N_22797,N_22621);
or U23464 (N_23464,N_22694,N_22668);
nand U23465 (N_23465,N_22812,N_22552);
nor U23466 (N_23466,N_22851,N_22715);
and U23467 (N_23467,N_22729,N_22978);
or U23468 (N_23468,N_22827,N_22611);
and U23469 (N_23469,N_22994,N_22766);
xnor U23470 (N_23470,N_22712,N_22810);
nand U23471 (N_23471,N_22783,N_22726);
nor U23472 (N_23472,N_22567,N_22608);
and U23473 (N_23473,N_22629,N_22873);
nand U23474 (N_23474,N_22572,N_22929);
nand U23475 (N_23475,N_22974,N_22656);
nor U23476 (N_23476,N_22650,N_22561);
or U23477 (N_23477,N_22954,N_22838);
nand U23478 (N_23478,N_22880,N_22582);
xnor U23479 (N_23479,N_22930,N_22926);
xor U23480 (N_23480,N_22661,N_22763);
or U23481 (N_23481,N_22922,N_22912);
or U23482 (N_23482,N_22745,N_22970);
xnor U23483 (N_23483,N_22929,N_22774);
nand U23484 (N_23484,N_22994,N_22693);
nand U23485 (N_23485,N_22972,N_22623);
or U23486 (N_23486,N_22561,N_22799);
nor U23487 (N_23487,N_22744,N_22541);
and U23488 (N_23488,N_22760,N_22692);
xnor U23489 (N_23489,N_22532,N_22893);
xnor U23490 (N_23490,N_22813,N_22553);
nand U23491 (N_23491,N_22966,N_22504);
and U23492 (N_23492,N_22870,N_22602);
and U23493 (N_23493,N_22896,N_22779);
or U23494 (N_23494,N_22703,N_22741);
xor U23495 (N_23495,N_22983,N_22825);
and U23496 (N_23496,N_22744,N_22612);
nor U23497 (N_23497,N_22995,N_22826);
nand U23498 (N_23498,N_22703,N_22855);
or U23499 (N_23499,N_22511,N_22962);
nand U23500 (N_23500,N_23105,N_23260);
nand U23501 (N_23501,N_23102,N_23018);
nor U23502 (N_23502,N_23132,N_23366);
nor U23503 (N_23503,N_23093,N_23436);
or U23504 (N_23504,N_23251,N_23185);
nand U23505 (N_23505,N_23006,N_23376);
or U23506 (N_23506,N_23298,N_23430);
nor U23507 (N_23507,N_23320,N_23291);
and U23508 (N_23508,N_23278,N_23177);
nor U23509 (N_23509,N_23374,N_23254);
and U23510 (N_23510,N_23181,N_23394);
nand U23511 (N_23511,N_23170,N_23414);
nand U23512 (N_23512,N_23387,N_23247);
nor U23513 (N_23513,N_23466,N_23079);
and U23514 (N_23514,N_23267,N_23174);
or U23515 (N_23515,N_23144,N_23141);
or U23516 (N_23516,N_23213,N_23187);
and U23517 (N_23517,N_23266,N_23489);
nor U23518 (N_23518,N_23294,N_23463);
nand U23519 (N_23519,N_23021,N_23194);
and U23520 (N_23520,N_23040,N_23250);
xor U23521 (N_23521,N_23146,N_23326);
or U23522 (N_23522,N_23014,N_23403);
xnor U23523 (N_23523,N_23425,N_23171);
and U23524 (N_23524,N_23275,N_23217);
xnor U23525 (N_23525,N_23419,N_23134);
nor U23526 (N_23526,N_23070,N_23051);
nor U23527 (N_23527,N_23169,N_23429);
or U23528 (N_23528,N_23000,N_23451);
nor U23529 (N_23529,N_23321,N_23306);
xnor U23530 (N_23530,N_23381,N_23485);
nand U23531 (N_23531,N_23026,N_23066);
nand U23532 (N_23532,N_23348,N_23074);
and U23533 (N_23533,N_23344,N_23442);
and U23534 (N_23534,N_23044,N_23087);
nand U23535 (N_23535,N_23449,N_23228);
and U23536 (N_23536,N_23071,N_23244);
or U23537 (N_23537,N_23407,N_23452);
and U23538 (N_23538,N_23428,N_23219);
nor U23539 (N_23539,N_23068,N_23384);
or U23540 (N_23540,N_23358,N_23475);
and U23541 (N_23541,N_23098,N_23148);
or U23542 (N_23542,N_23032,N_23340);
or U23543 (N_23543,N_23184,N_23198);
nand U23544 (N_23544,N_23164,N_23193);
nand U23545 (N_23545,N_23375,N_23365);
nand U23546 (N_23546,N_23469,N_23269);
and U23547 (N_23547,N_23318,N_23367);
or U23548 (N_23548,N_23092,N_23031);
nand U23549 (N_23549,N_23133,N_23159);
and U23550 (N_23550,N_23166,N_23048);
xor U23551 (N_23551,N_23362,N_23317);
xor U23552 (N_23552,N_23095,N_23399);
or U23553 (N_23553,N_23036,N_23086);
or U23554 (N_23554,N_23229,N_23163);
or U23555 (N_23555,N_23082,N_23349);
nor U23556 (N_23556,N_23446,N_23025);
nand U23557 (N_23557,N_23136,N_23015);
nand U23558 (N_23558,N_23010,N_23314);
or U23559 (N_23559,N_23024,N_23293);
nand U23560 (N_23560,N_23474,N_23034);
nor U23561 (N_23561,N_23050,N_23478);
nand U23562 (N_23562,N_23303,N_23233);
nand U23563 (N_23563,N_23380,N_23441);
nand U23564 (N_23564,N_23234,N_23307);
nor U23565 (N_23565,N_23055,N_23495);
or U23566 (N_23566,N_23265,N_23395);
xor U23567 (N_23567,N_23491,N_23208);
and U23568 (N_23568,N_23096,N_23085);
or U23569 (N_23569,N_23424,N_23329);
xor U23570 (N_23570,N_23360,N_23322);
or U23571 (N_23571,N_23204,N_23118);
or U23572 (N_23572,N_23196,N_23179);
nand U23573 (N_23573,N_23042,N_23094);
or U23574 (N_23574,N_23284,N_23494);
xor U23575 (N_23575,N_23249,N_23461);
xor U23576 (N_23576,N_23274,N_23112);
xor U23577 (N_23577,N_23155,N_23062);
nand U23578 (N_23578,N_23203,N_23043);
or U23579 (N_23579,N_23296,N_23084);
and U23580 (N_23580,N_23205,N_23427);
nor U23581 (N_23581,N_23346,N_23178);
and U23582 (N_23582,N_23063,N_23336);
or U23583 (N_23583,N_23078,N_23154);
nand U23584 (N_23584,N_23045,N_23257);
nor U23585 (N_23585,N_23361,N_23412);
or U23586 (N_23586,N_23471,N_23191);
xor U23587 (N_23587,N_23328,N_23481);
xor U23588 (N_23588,N_23160,N_23180);
or U23589 (N_23589,N_23280,N_23435);
and U23590 (N_23590,N_23147,N_23281);
nor U23591 (N_23591,N_23288,N_23190);
nand U23592 (N_23592,N_23029,N_23310);
nand U23593 (N_23593,N_23450,N_23099);
or U23594 (N_23594,N_23343,N_23140);
nor U23595 (N_23595,N_23268,N_23312);
or U23596 (N_23596,N_23156,N_23447);
or U23597 (N_23597,N_23316,N_23300);
xor U23598 (N_23598,N_23319,N_23142);
nor U23599 (N_23599,N_23121,N_23245);
or U23600 (N_23600,N_23167,N_23377);
nor U23601 (N_23601,N_23270,N_23123);
xnor U23602 (N_23602,N_23182,N_23420);
xor U23603 (N_23603,N_23347,N_23058);
nor U23604 (N_23604,N_23152,N_23341);
or U23605 (N_23605,N_23331,N_23027);
or U23606 (N_23606,N_23458,N_23139);
xnor U23607 (N_23607,N_23484,N_23223);
xnor U23608 (N_23608,N_23426,N_23324);
nand U23609 (N_23609,N_23261,N_23402);
nand U23610 (N_23610,N_23113,N_23482);
and U23611 (N_23611,N_23172,N_23342);
and U23612 (N_23612,N_23286,N_23235);
xor U23613 (N_23613,N_23097,N_23131);
and U23614 (N_23614,N_23413,N_23090);
xnor U23615 (N_23615,N_23345,N_23214);
nor U23616 (N_23616,N_23248,N_23039);
nand U23617 (N_23617,N_23129,N_23143);
and U23618 (N_23618,N_23239,N_23210);
or U23619 (N_23619,N_23130,N_23415);
or U23620 (N_23620,N_23437,N_23215);
and U23621 (N_23621,N_23041,N_23007);
or U23622 (N_23622,N_23397,N_23005);
xor U23623 (N_23623,N_23158,N_23400);
xor U23624 (N_23624,N_23401,N_23335);
nor U23625 (N_23625,N_23462,N_23243);
nand U23626 (N_23626,N_23404,N_23357);
xnor U23627 (N_23627,N_23101,N_23202);
xnor U23628 (N_23628,N_23313,N_23126);
and U23629 (N_23629,N_23115,N_23081);
or U23630 (N_23630,N_23359,N_23356);
nand U23631 (N_23631,N_23054,N_23282);
or U23632 (N_23632,N_23059,N_23236);
xnor U23633 (N_23633,N_23216,N_23417);
xor U23634 (N_23634,N_23137,N_23109);
or U23635 (N_23635,N_23089,N_23271);
nand U23636 (N_23636,N_23301,N_23150);
nor U23637 (N_23637,N_23393,N_23057);
nor U23638 (N_23638,N_23411,N_23338);
nand U23639 (N_23639,N_23108,N_23127);
nand U23640 (N_23640,N_23408,N_23200);
nor U23641 (N_23641,N_23145,N_23199);
or U23642 (N_23642,N_23297,N_23370);
nor U23643 (N_23643,N_23276,N_23207);
xor U23644 (N_23644,N_23290,N_23398);
nor U23645 (N_23645,N_23176,N_23434);
nor U23646 (N_23646,N_23022,N_23339);
and U23647 (N_23647,N_23444,N_23473);
nor U23648 (N_23648,N_23020,N_23222);
nand U23649 (N_23649,N_23479,N_23038);
xor U23650 (N_23650,N_23119,N_23008);
nor U23651 (N_23651,N_23240,N_23149);
nand U23652 (N_23652,N_23225,N_23459);
nor U23653 (N_23653,N_23226,N_23299);
and U23654 (N_23654,N_23457,N_23383);
nand U23655 (N_23655,N_23390,N_23464);
nor U23656 (N_23656,N_23488,N_23388);
nor U23657 (N_23657,N_23162,N_23253);
and U23658 (N_23658,N_23378,N_23262);
nor U23659 (N_23659,N_23151,N_23332);
and U23660 (N_23660,N_23073,N_23002);
and U23661 (N_23661,N_23497,N_23418);
nand U23662 (N_23662,N_23480,N_23364);
nand U23663 (N_23663,N_23238,N_23256);
and U23664 (N_23664,N_23333,N_23077);
or U23665 (N_23665,N_23135,N_23019);
or U23666 (N_23666,N_23227,N_23075);
and U23667 (N_23667,N_23231,N_23107);
nand U23668 (N_23668,N_23487,N_23277);
and U23669 (N_23669,N_23003,N_23153);
nor U23670 (N_23670,N_23389,N_23432);
xor U23671 (N_23671,N_23258,N_23035);
or U23672 (N_23672,N_23117,N_23354);
and U23673 (N_23673,N_23103,N_23443);
or U23674 (N_23674,N_23211,N_23052);
and U23675 (N_23675,N_23100,N_23065);
and U23676 (N_23676,N_23212,N_23334);
or U23677 (N_23677,N_23421,N_23188);
nand U23678 (N_23678,N_23273,N_23173);
nor U23679 (N_23679,N_23499,N_23009);
and U23680 (N_23680,N_23352,N_23165);
nor U23681 (N_23681,N_23241,N_23279);
xor U23682 (N_23682,N_23138,N_23350);
and U23683 (N_23683,N_23012,N_23124);
and U23684 (N_23684,N_23422,N_23323);
or U23685 (N_23685,N_23295,N_23477);
nand U23686 (N_23686,N_23011,N_23272);
or U23687 (N_23687,N_23056,N_23285);
nand U23688 (N_23688,N_23183,N_23372);
nor U23689 (N_23689,N_23283,N_23302);
and U23690 (N_23690,N_23416,N_23453);
and U23691 (N_23691,N_23385,N_23330);
or U23692 (N_23692,N_23379,N_23033);
nor U23693 (N_23693,N_23083,N_23327);
or U23694 (N_23694,N_23091,N_23391);
xnor U23695 (N_23695,N_23472,N_23197);
and U23696 (N_23696,N_23246,N_23467);
nor U23697 (N_23697,N_23396,N_23221);
xor U23698 (N_23698,N_23433,N_23287);
or U23699 (N_23699,N_23496,N_23493);
or U23700 (N_23700,N_23355,N_23255);
nand U23701 (N_23701,N_23114,N_23309);
nor U23702 (N_23702,N_23168,N_23460);
and U23703 (N_23703,N_23195,N_23064);
nor U23704 (N_23704,N_23382,N_23060);
nor U23705 (N_23705,N_23337,N_23454);
nand U23706 (N_23706,N_23498,N_23049);
and U23707 (N_23707,N_23061,N_23351);
nand U23708 (N_23708,N_23111,N_23106);
nor U23709 (N_23709,N_23023,N_23264);
or U23710 (N_23710,N_23468,N_23325);
nand U23711 (N_23711,N_23311,N_23028);
nand U23712 (N_23712,N_23292,N_23161);
nand U23713 (N_23713,N_23369,N_23186);
or U23714 (N_23714,N_23004,N_23386);
nand U23715 (N_23715,N_23486,N_23069);
and U23716 (N_23716,N_23259,N_23455);
nor U23717 (N_23717,N_23076,N_23465);
and U23718 (N_23718,N_23220,N_23305);
nor U23719 (N_23719,N_23353,N_23067);
nand U23720 (N_23720,N_23209,N_23431);
or U23721 (N_23721,N_23104,N_23122);
nand U23722 (N_23722,N_23047,N_23410);
nor U23723 (N_23723,N_23440,N_23201);
nand U23724 (N_23724,N_23175,N_23189);
or U23725 (N_23725,N_23476,N_23110);
or U23726 (N_23726,N_23406,N_23363);
nor U23727 (N_23727,N_23423,N_23315);
nor U23728 (N_23728,N_23373,N_23289);
xor U23729 (N_23729,N_23120,N_23252);
and U23730 (N_23730,N_23116,N_23013);
or U23731 (N_23731,N_23445,N_23088);
and U23732 (N_23732,N_23371,N_23206);
or U23733 (N_23733,N_23304,N_23368);
nand U23734 (N_23734,N_23224,N_23490);
or U23735 (N_23735,N_23263,N_23218);
xnor U23736 (N_23736,N_23157,N_23470);
nor U23737 (N_23737,N_23405,N_23456);
and U23738 (N_23738,N_23392,N_23125);
or U23739 (N_23739,N_23053,N_23438);
nand U23740 (N_23740,N_23016,N_23037);
or U23741 (N_23741,N_23046,N_23080);
or U23742 (N_23742,N_23230,N_23492);
nand U23743 (N_23743,N_23483,N_23448);
nor U23744 (N_23744,N_23072,N_23030);
and U23745 (N_23745,N_23308,N_23237);
nand U23746 (N_23746,N_23242,N_23017);
nand U23747 (N_23747,N_23439,N_23128);
or U23748 (N_23748,N_23409,N_23192);
nand U23749 (N_23749,N_23232,N_23001);
xnor U23750 (N_23750,N_23426,N_23314);
nand U23751 (N_23751,N_23433,N_23147);
or U23752 (N_23752,N_23479,N_23358);
or U23753 (N_23753,N_23174,N_23090);
xor U23754 (N_23754,N_23463,N_23488);
xnor U23755 (N_23755,N_23080,N_23364);
nand U23756 (N_23756,N_23461,N_23490);
nand U23757 (N_23757,N_23393,N_23301);
xnor U23758 (N_23758,N_23055,N_23484);
and U23759 (N_23759,N_23488,N_23142);
nand U23760 (N_23760,N_23025,N_23035);
or U23761 (N_23761,N_23234,N_23489);
xnor U23762 (N_23762,N_23316,N_23382);
nor U23763 (N_23763,N_23419,N_23477);
nor U23764 (N_23764,N_23193,N_23056);
xnor U23765 (N_23765,N_23125,N_23068);
or U23766 (N_23766,N_23482,N_23148);
nand U23767 (N_23767,N_23197,N_23108);
nand U23768 (N_23768,N_23031,N_23209);
xnor U23769 (N_23769,N_23059,N_23069);
nand U23770 (N_23770,N_23491,N_23133);
xnor U23771 (N_23771,N_23095,N_23128);
and U23772 (N_23772,N_23471,N_23337);
nor U23773 (N_23773,N_23309,N_23203);
or U23774 (N_23774,N_23028,N_23086);
xnor U23775 (N_23775,N_23438,N_23082);
nor U23776 (N_23776,N_23249,N_23003);
xnor U23777 (N_23777,N_23310,N_23429);
xor U23778 (N_23778,N_23094,N_23322);
xor U23779 (N_23779,N_23231,N_23250);
and U23780 (N_23780,N_23111,N_23324);
and U23781 (N_23781,N_23274,N_23439);
or U23782 (N_23782,N_23368,N_23477);
xnor U23783 (N_23783,N_23342,N_23376);
and U23784 (N_23784,N_23036,N_23153);
and U23785 (N_23785,N_23092,N_23320);
nand U23786 (N_23786,N_23040,N_23057);
nor U23787 (N_23787,N_23116,N_23053);
nand U23788 (N_23788,N_23226,N_23430);
or U23789 (N_23789,N_23274,N_23206);
xnor U23790 (N_23790,N_23193,N_23366);
and U23791 (N_23791,N_23285,N_23207);
xnor U23792 (N_23792,N_23157,N_23167);
nand U23793 (N_23793,N_23193,N_23401);
nand U23794 (N_23794,N_23097,N_23444);
nor U23795 (N_23795,N_23382,N_23221);
xor U23796 (N_23796,N_23000,N_23122);
xor U23797 (N_23797,N_23368,N_23498);
nand U23798 (N_23798,N_23450,N_23038);
nor U23799 (N_23799,N_23444,N_23365);
nor U23800 (N_23800,N_23361,N_23033);
and U23801 (N_23801,N_23142,N_23462);
nor U23802 (N_23802,N_23352,N_23215);
nor U23803 (N_23803,N_23239,N_23452);
xnor U23804 (N_23804,N_23297,N_23424);
and U23805 (N_23805,N_23294,N_23201);
and U23806 (N_23806,N_23432,N_23433);
xnor U23807 (N_23807,N_23089,N_23471);
and U23808 (N_23808,N_23175,N_23193);
and U23809 (N_23809,N_23040,N_23287);
and U23810 (N_23810,N_23336,N_23145);
xnor U23811 (N_23811,N_23469,N_23413);
nor U23812 (N_23812,N_23103,N_23486);
xor U23813 (N_23813,N_23020,N_23199);
nor U23814 (N_23814,N_23419,N_23174);
or U23815 (N_23815,N_23087,N_23021);
or U23816 (N_23816,N_23157,N_23378);
xnor U23817 (N_23817,N_23253,N_23093);
nor U23818 (N_23818,N_23388,N_23404);
nor U23819 (N_23819,N_23139,N_23382);
and U23820 (N_23820,N_23220,N_23200);
and U23821 (N_23821,N_23135,N_23065);
or U23822 (N_23822,N_23492,N_23490);
nor U23823 (N_23823,N_23093,N_23255);
or U23824 (N_23824,N_23251,N_23112);
nor U23825 (N_23825,N_23037,N_23353);
xor U23826 (N_23826,N_23366,N_23012);
nand U23827 (N_23827,N_23128,N_23491);
or U23828 (N_23828,N_23070,N_23020);
xnor U23829 (N_23829,N_23002,N_23340);
or U23830 (N_23830,N_23413,N_23099);
nor U23831 (N_23831,N_23025,N_23439);
nand U23832 (N_23832,N_23139,N_23122);
nand U23833 (N_23833,N_23273,N_23108);
nor U23834 (N_23834,N_23471,N_23320);
nand U23835 (N_23835,N_23372,N_23475);
or U23836 (N_23836,N_23481,N_23269);
xor U23837 (N_23837,N_23375,N_23476);
nand U23838 (N_23838,N_23169,N_23127);
nor U23839 (N_23839,N_23272,N_23283);
nand U23840 (N_23840,N_23396,N_23273);
xnor U23841 (N_23841,N_23181,N_23496);
xor U23842 (N_23842,N_23209,N_23032);
or U23843 (N_23843,N_23360,N_23280);
nand U23844 (N_23844,N_23236,N_23028);
and U23845 (N_23845,N_23291,N_23201);
nand U23846 (N_23846,N_23294,N_23381);
xor U23847 (N_23847,N_23327,N_23047);
nand U23848 (N_23848,N_23065,N_23284);
or U23849 (N_23849,N_23246,N_23448);
xor U23850 (N_23850,N_23007,N_23087);
nor U23851 (N_23851,N_23323,N_23450);
nor U23852 (N_23852,N_23312,N_23140);
or U23853 (N_23853,N_23313,N_23328);
xnor U23854 (N_23854,N_23307,N_23346);
xnor U23855 (N_23855,N_23201,N_23322);
nand U23856 (N_23856,N_23400,N_23352);
or U23857 (N_23857,N_23304,N_23398);
nor U23858 (N_23858,N_23418,N_23184);
or U23859 (N_23859,N_23255,N_23472);
xnor U23860 (N_23860,N_23275,N_23186);
nor U23861 (N_23861,N_23421,N_23165);
nor U23862 (N_23862,N_23219,N_23336);
nand U23863 (N_23863,N_23251,N_23442);
or U23864 (N_23864,N_23363,N_23414);
or U23865 (N_23865,N_23279,N_23302);
xor U23866 (N_23866,N_23495,N_23299);
nand U23867 (N_23867,N_23395,N_23075);
nor U23868 (N_23868,N_23105,N_23406);
and U23869 (N_23869,N_23268,N_23332);
xnor U23870 (N_23870,N_23388,N_23155);
and U23871 (N_23871,N_23412,N_23167);
and U23872 (N_23872,N_23255,N_23150);
xnor U23873 (N_23873,N_23164,N_23174);
nand U23874 (N_23874,N_23368,N_23402);
or U23875 (N_23875,N_23296,N_23065);
or U23876 (N_23876,N_23181,N_23409);
nor U23877 (N_23877,N_23284,N_23423);
nand U23878 (N_23878,N_23202,N_23199);
nand U23879 (N_23879,N_23335,N_23019);
nor U23880 (N_23880,N_23134,N_23003);
and U23881 (N_23881,N_23210,N_23265);
xnor U23882 (N_23882,N_23277,N_23044);
and U23883 (N_23883,N_23226,N_23074);
or U23884 (N_23884,N_23458,N_23422);
and U23885 (N_23885,N_23030,N_23249);
nor U23886 (N_23886,N_23018,N_23233);
nor U23887 (N_23887,N_23489,N_23061);
xnor U23888 (N_23888,N_23085,N_23478);
xnor U23889 (N_23889,N_23302,N_23259);
nor U23890 (N_23890,N_23468,N_23057);
nand U23891 (N_23891,N_23246,N_23304);
xnor U23892 (N_23892,N_23432,N_23187);
nand U23893 (N_23893,N_23115,N_23017);
nor U23894 (N_23894,N_23284,N_23294);
and U23895 (N_23895,N_23384,N_23098);
nand U23896 (N_23896,N_23458,N_23185);
nor U23897 (N_23897,N_23116,N_23077);
and U23898 (N_23898,N_23470,N_23068);
nand U23899 (N_23899,N_23037,N_23400);
and U23900 (N_23900,N_23377,N_23271);
and U23901 (N_23901,N_23208,N_23054);
nor U23902 (N_23902,N_23450,N_23427);
nand U23903 (N_23903,N_23085,N_23333);
and U23904 (N_23904,N_23397,N_23372);
nand U23905 (N_23905,N_23281,N_23372);
nor U23906 (N_23906,N_23021,N_23302);
or U23907 (N_23907,N_23451,N_23033);
and U23908 (N_23908,N_23499,N_23260);
nor U23909 (N_23909,N_23217,N_23334);
nand U23910 (N_23910,N_23054,N_23490);
nand U23911 (N_23911,N_23075,N_23107);
nor U23912 (N_23912,N_23314,N_23177);
nand U23913 (N_23913,N_23034,N_23075);
or U23914 (N_23914,N_23268,N_23035);
xnor U23915 (N_23915,N_23378,N_23190);
or U23916 (N_23916,N_23101,N_23042);
and U23917 (N_23917,N_23368,N_23218);
nand U23918 (N_23918,N_23208,N_23092);
or U23919 (N_23919,N_23384,N_23365);
nor U23920 (N_23920,N_23477,N_23053);
or U23921 (N_23921,N_23373,N_23293);
nor U23922 (N_23922,N_23172,N_23488);
nand U23923 (N_23923,N_23218,N_23461);
xnor U23924 (N_23924,N_23356,N_23114);
xor U23925 (N_23925,N_23223,N_23133);
nor U23926 (N_23926,N_23030,N_23479);
nor U23927 (N_23927,N_23494,N_23322);
nor U23928 (N_23928,N_23473,N_23128);
nor U23929 (N_23929,N_23434,N_23276);
nor U23930 (N_23930,N_23283,N_23249);
xor U23931 (N_23931,N_23028,N_23354);
nor U23932 (N_23932,N_23014,N_23341);
or U23933 (N_23933,N_23019,N_23287);
nor U23934 (N_23934,N_23398,N_23148);
nand U23935 (N_23935,N_23393,N_23492);
or U23936 (N_23936,N_23314,N_23027);
and U23937 (N_23937,N_23491,N_23111);
or U23938 (N_23938,N_23199,N_23002);
nand U23939 (N_23939,N_23300,N_23455);
nor U23940 (N_23940,N_23161,N_23382);
and U23941 (N_23941,N_23118,N_23110);
or U23942 (N_23942,N_23484,N_23202);
xnor U23943 (N_23943,N_23428,N_23301);
nand U23944 (N_23944,N_23014,N_23413);
or U23945 (N_23945,N_23192,N_23319);
nand U23946 (N_23946,N_23488,N_23015);
nand U23947 (N_23947,N_23382,N_23368);
and U23948 (N_23948,N_23413,N_23249);
or U23949 (N_23949,N_23017,N_23386);
nor U23950 (N_23950,N_23117,N_23398);
xnor U23951 (N_23951,N_23200,N_23239);
xnor U23952 (N_23952,N_23397,N_23329);
or U23953 (N_23953,N_23146,N_23088);
xnor U23954 (N_23954,N_23416,N_23105);
nand U23955 (N_23955,N_23498,N_23457);
xnor U23956 (N_23956,N_23388,N_23372);
nor U23957 (N_23957,N_23476,N_23388);
nand U23958 (N_23958,N_23315,N_23030);
and U23959 (N_23959,N_23288,N_23401);
xnor U23960 (N_23960,N_23246,N_23013);
and U23961 (N_23961,N_23080,N_23458);
or U23962 (N_23962,N_23182,N_23344);
xor U23963 (N_23963,N_23087,N_23201);
nor U23964 (N_23964,N_23171,N_23043);
or U23965 (N_23965,N_23033,N_23123);
nor U23966 (N_23966,N_23273,N_23453);
nor U23967 (N_23967,N_23187,N_23380);
xor U23968 (N_23968,N_23221,N_23194);
nor U23969 (N_23969,N_23034,N_23403);
or U23970 (N_23970,N_23164,N_23023);
xnor U23971 (N_23971,N_23353,N_23419);
nand U23972 (N_23972,N_23185,N_23296);
and U23973 (N_23973,N_23369,N_23040);
or U23974 (N_23974,N_23103,N_23126);
nor U23975 (N_23975,N_23109,N_23394);
and U23976 (N_23976,N_23197,N_23111);
xnor U23977 (N_23977,N_23429,N_23283);
and U23978 (N_23978,N_23132,N_23352);
nor U23979 (N_23979,N_23104,N_23136);
xnor U23980 (N_23980,N_23159,N_23239);
and U23981 (N_23981,N_23472,N_23215);
nor U23982 (N_23982,N_23384,N_23461);
and U23983 (N_23983,N_23005,N_23142);
nor U23984 (N_23984,N_23157,N_23343);
xnor U23985 (N_23985,N_23403,N_23487);
or U23986 (N_23986,N_23015,N_23347);
xor U23987 (N_23987,N_23342,N_23131);
nand U23988 (N_23988,N_23397,N_23384);
nor U23989 (N_23989,N_23272,N_23030);
nand U23990 (N_23990,N_23327,N_23207);
nor U23991 (N_23991,N_23259,N_23060);
xor U23992 (N_23992,N_23212,N_23096);
or U23993 (N_23993,N_23151,N_23321);
and U23994 (N_23994,N_23338,N_23072);
or U23995 (N_23995,N_23281,N_23363);
nor U23996 (N_23996,N_23090,N_23314);
and U23997 (N_23997,N_23314,N_23358);
nand U23998 (N_23998,N_23143,N_23478);
nor U23999 (N_23999,N_23125,N_23017);
or U24000 (N_24000,N_23734,N_23936);
nor U24001 (N_24001,N_23971,N_23821);
and U24002 (N_24002,N_23602,N_23978);
or U24003 (N_24003,N_23765,N_23860);
xnor U24004 (N_24004,N_23776,N_23916);
nand U24005 (N_24005,N_23729,N_23795);
nand U24006 (N_24006,N_23619,N_23910);
or U24007 (N_24007,N_23719,N_23738);
xor U24008 (N_24008,N_23584,N_23632);
and U24009 (N_24009,N_23702,N_23613);
and U24010 (N_24010,N_23942,N_23786);
nand U24011 (N_24011,N_23504,N_23559);
nor U24012 (N_24012,N_23688,N_23645);
or U24013 (N_24013,N_23778,N_23522);
xnor U24014 (N_24014,N_23984,N_23953);
or U24015 (N_24015,N_23648,N_23892);
xnor U24016 (N_24016,N_23889,N_23770);
nor U24017 (N_24017,N_23638,N_23974);
xor U24018 (N_24018,N_23835,N_23735);
nor U24019 (N_24019,N_23579,N_23580);
nor U24020 (N_24020,N_23950,N_23516);
xnor U24021 (N_24021,N_23962,N_23788);
nand U24022 (N_24022,N_23641,N_23678);
nor U24023 (N_24023,N_23649,N_23654);
and U24024 (N_24024,N_23939,N_23669);
nand U24025 (N_24025,N_23940,N_23752);
nor U24026 (N_24026,N_23699,N_23544);
xnor U24027 (N_24027,N_23691,N_23506);
nor U24028 (N_24028,N_23881,N_23829);
and U24029 (N_24029,N_23594,N_23637);
nand U24030 (N_24030,N_23848,N_23747);
and U24031 (N_24031,N_23710,N_23792);
or U24032 (N_24032,N_23855,N_23592);
xnor U24033 (N_24033,N_23670,N_23650);
or U24034 (N_24034,N_23764,N_23888);
nand U24035 (N_24035,N_23882,N_23864);
or U24036 (N_24036,N_23988,N_23818);
or U24037 (N_24037,N_23926,N_23982);
or U24038 (N_24038,N_23557,N_23871);
or U24039 (N_24039,N_23983,N_23861);
nor U24040 (N_24040,N_23811,N_23514);
nor U24041 (N_24041,N_23798,N_23577);
or U24042 (N_24042,N_23865,N_23543);
or U24043 (N_24043,N_23724,N_23964);
nor U24044 (N_24044,N_23524,N_23558);
xor U24045 (N_24045,N_23695,N_23884);
xor U24046 (N_24046,N_23501,N_23730);
nand U24047 (N_24047,N_23887,N_23685);
nand U24048 (N_24048,N_23521,N_23920);
or U24049 (N_24049,N_23773,N_23938);
nor U24050 (N_24050,N_23966,N_23679);
or U24051 (N_24051,N_23709,N_23624);
nor U24052 (N_24052,N_23947,N_23525);
or U24053 (N_24053,N_23529,N_23631);
or U24054 (N_24054,N_23777,N_23753);
xor U24055 (N_24055,N_23622,N_23697);
or U24056 (N_24056,N_23831,N_23933);
and U24057 (N_24057,N_23652,N_23666);
nand U24058 (N_24058,N_23576,N_23693);
xor U24059 (N_24059,N_23783,N_23875);
xnor U24060 (N_24060,N_23741,N_23689);
xor U24061 (N_24061,N_23834,N_23780);
and U24062 (N_24062,N_23760,N_23690);
nand U24063 (N_24063,N_23832,N_23844);
nand U24064 (N_24064,N_23826,N_23937);
and U24065 (N_24065,N_23841,N_23593);
and U24066 (N_24066,N_23858,N_23909);
nor U24067 (N_24067,N_23737,N_23554);
nor U24068 (N_24068,N_23616,N_23879);
nor U24069 (N_24069,N_23756,N_23902);
xnor U24070 (N_24070,N_23813,N_23930);
or U24071 (N_24071,N_23534,N_23842);
nor U24072 (N_24072,N_23546,N_23564);
nor U24073 (N_24073,N_23548,N_23712);
or U24074 (N_24074,N_23601,N_23809);
nor U24075 (N_24075,N_23611,N_23680);
nor U24076 (N_24076,N_23732,N_23904);
and U24077 (N_24077,N_23701,N_23928);
nand U24078 (N_24078,N_23533,N_23791);
or U24079 (N_24079,N_23977,N_23853);
nor U24080 (N_24080,N_23633,N_23627);
xor U24081 (N_24081,N_23572,N_23567);
xor U24082 (N_24082,N_23790,N_23664);
or U24083 (N_24083,N_23850,N_23614);
or U24084 (N_24084,N_23600,N_23812);
nor U24085 (N_24085,N_23530,N_23932);
or U24086 (N_24086,N_23986,N_23746);
and U24087 (N_24087,N_23662,N_23965);
xnor U24088 (N_24088,N_23757,N_23801);
or U24089 (N_24089,N_23946,N_23672);
nand U24090 (N_24090,N_23763,N_23658);
or U24091 (N_24091,N_23870,N_23714);
nor U24092 (N_24092,N_23895,N_23931);
and U24093 (N_24093,N_23610,N_23976);
nand U24094 (N_24094,N_23805,N_23852);
and U24095 (N_24095,N_23893,N_23868);
nor U24096 (N_24096,N_23731,N_23907);
nor U24097 (N_24097,N_23707,N_23617);
nand U24098 (N_24098,N_23511,N_23566);
or U24099 (N_24099,N_23869,N_23625);
or U24100 (N_24100,N_23924,N_23840);
xnor U24101 (N_24101,N_23628,N_23912);
or U24102 (N_24102,N_23656,N_23908);
nor U24103 (N_24103,N_23991,N_23599);
xnor U24104 (N_24104,N_23513,N_23720);
nor U24105 (N_24105,N_23767,N_23708);
nor U24106 (N_24106,N_23716,N_23794);
nand U24107 (N_24107,N_23929,N_23995);
xor U24108 (N_24108,N_23793,N_23817);
and U24109 (N_24109,N_23553,N_23605);
and U24110 (N_24110,N_23814,N_23917);
or U24111 (N_24111,N_23620,N_23634);
xnor U24112 (N_24112,N_23660,N_23948);
nor U24113 (N_24113,N_23549,N_23980);
or U24114 (N_24114,N_23985,N_23992);
nand U24115 (N_24115,N_23957,N_23918);
or U24116 (N_24116,N_23872,N_23675);
xor U24117 (N_24117,N_23563,N_23545);
and U24118 (N_24118,N_23682,N_23630);
or U24119 (N_24119,N_23542,N_23919);
nor U24120 (N_24120,N_23526,N_23900);
nor U24121 (N_24121,N_23998,N_23540);
nor U24122 (N_24122,N_23573,N_23515);
or U24123 (N_24123,N_23725,N_23717);
nand U24124 (N_24124,N_23990,N_23659);
nor U24125 (N_24125,N_23674,N_23999);
nor U24126 (N_24126,N_23569,N_23843);
and U24127 (N_24127,N_23538,N_23830);
nand U24128 (N_24128,N_23866,N_23694);
nor U24129 (N_24129,N_23596,N_23635);
nand U24130 (N_24130,N_23651,N_23905);
or U24131 (N_24131,N_23973,N_23722);
nor U24132 (N_24132,N_23705,N_23921);
nor U24133 (N_24133,N_23582,N_23657);
or U24134 (N_24134,N_23959,N_23531);
nor U24135 (N_24135,N_23551,N_23598);
nand U24136 (N_24136,N_23517,N_23597);
and U24137 (N_24137,N_23621,N_23862);
and U24138 (N_24138,N_23663,N_23754);
nor U24139 (N_24139,N_23797,N_23804);
and U24140 (N_24140,N_23750,N_23556);
nor U24141 (N_24141,N_23951,N_23822);
nand U24142 (N_24142,N_23775,N_23595);
nor U24143 (N_24143,N_23703,N_23915);
or U24144 (N_24144,N_23827,N_23519);
and U24145 (N_24145,N_23583,N_23771);
nand U24146 (N_24146,N_23736,N_23823);
nand U24147 (N_24147,N_23997,N_23839);
xor U24148 (N_24148,N_23854,N_23768);
nand U24149 (N_24149,N_23743,N_23615);
xor U24150 (N_24150,N_23500,N_23774);
nand U24151 (N_24151,N_23759,N_23537);
nor U24152 (N_24152,N_23568,N_23897);
xor U24153 (N_24153,N_23837,N_23608);
nand U24154 (N_24154,N_23604,N_23640);
xor U24155 (N_24155,N_23914,N_23541);
xnor U24156 (N_24156,N_23518,N_23952);
xor U24157 (N_24157,N_23643,N_23943);
or U24158 (N_24158,N_23913,N_23956);
nor U24159 (N_24159,N_23787,N_23589);
or U24160 (N_24160,N_23681,N_23846);
or U24161 (N_24161,N_23954,N_23536);
nand U24162 (N_24162,N_23588,N_23578);
or U24163 (N_24163,N_23781,N_23935);
and U24164 (N_24164,N_23796,N_23994);
nor U24165 (N_24165,N_23642,N_23883);
xor U24166 (N_24166,N_23603,N_23816);
or U24167 (N_24167,N_23606,N_23799);
and U24168 (N_24168,N_23609,N_23739);
or U24169 (N_24169,N_23721,N_23700);
and U24170 (N_24170,N_23874,N_23993);
xor U24171 (N_24171,N_23876,N_23886);
or U24172 (N_24172,N_23845,N_23510);
nand U24173 (N_24173,N_23550,N_23945);
or U24174 (N_24174,N_23698,N_23981);
nand U24175 (N_24175,N_23728,N_23740);
nand U24176 (N_24176,N_23590,N_23806);
nand U24177 (N_24177,N_23671,N_23639);
xor U24178 (N_24178,N_23989,N_23607);
nor U24179 (N_24179,N_23713,N_23684);
or U24180 (N_24180,N_23523,N_23857);
and U24181 (N_24181,N_23673,N_23968);
and U24182 (N_24182,N_23944,N_23911);
nand U24183 (N_24183,N_23547,N_23979);
nor U24184 (N_24184,N_23923,N_23718);
nor U24185 (N_24185,N_23667,N_23969);
nand U24186 (N_24186,N_23894,N_23512);
xnor U24187 (N_24187,N_23751,N_23655);
or U24188 (N_24188,N_23644,N_23901);
nand U24189 (N_24189,N_23899,N_23555);
nor U24190 (N_24190,N_23769,N_23960);
nand U24191 (N_24191,N_23803,N_23890);
or U24192 (N_24192,N_23665,N_23810);
or U24193 (N_24193,N_23758,N_23742);
xnor U24194 (N_24194,N_23967,N_23898);
xnor U24195 (N_24195,N_23970,N_23727);
nand U24196 (N_24196,N_23527,N_23653);
or U24197 (N_24197,N_23687,N_23851);
and U24198 (N_24198,N_23711,N_23560);
xnor U24199 (N_24199,N_23575,N_23867);
or U24200 (N_24200,N_23683,N_23896);
nor U24201 (N_24201,N_23748,N_23772);
xnor U24202 (N_24202,N_23704,N_23612);
and U24203 (N_24203,N_23880,N_23520);
nor U24204 (N_24204,N_23585,N_23661);
or U24205 (N_24205,N_23996,N_23927);
or U24206 (N_24206,N_23784,N_23581);
or U24207 (N_24207,N_23949,N_23975);
xor U24208 (N_24208,N_23668,N_23779);
nor U24209 (N_24209,N_23903,N_23509);
nand U24210 (N_24210,N_23528,N_23819);
nand U24211 (N_24211,N_23587,N_23696);
xor U24212 (N_24212,N_23877,N_23733);
xnor U24213 (N_24213,N_23802,N_23925);
or U24214 (N_24214,N_23824,N_23987);
or U24215 (N_24215,N_23906,N_23676);
nor U24216 (N_24216,N_23565,N_23873);
and U24217 (N_24217,N_23618,N_23677);
and U24218 (N_24218,N_23539,N_23561);
or U24219 (N_24219,N_23503,N_23508);
nand U24220 (N_24220,N_23552,N_23891);
and U24221 (N_24221,N_23505,N_23825);
xor U24222 (N_24222,N_23847,N_23828);
or U24223 (N_24223,N_23745,N_23726);
and U24224 (N_24224,N_23502,N_23838);
nor U24225 (N_24225,N_23715,N_23692);
and U24226 (N_24226,N_23961,N_23836);
and U24227 (N_24227,N_23972,N_23629);
or U24228 (N_24228,N_23808,N_23766);
and U24229 (N_24229,N_23863,N_23815);
and U24230 (N_24230,N_23623,N_23586);
and U24231 (N_24231,N_23785,N_23749);
nor U24232 (N_24232,N_23646,N_23762);
xor U24233 (N_24233,N_23859,N_23571);
nor U24234 (N_24234,N_23755,N_23570);
nand U24235 (N_24235,N_23507,N_23934);
and U24236 (N_24236,N_23562,N_23833);
or U24237 (N_24237,N_23686,N_23723);
nand U24238 (N_24238,N_23647,N_23574);
nor U24239 (N_24239,N_23744,N_23789);
xnor U24240 (N_24240,N_23955,N_23885);
and U24241 (N_24241,N_23782,N_23941);
xor U24242 (N_24242,N_23922,N_23761);
nand U24243 (N_24243,N_23849,N_23963);
and U24244 (N_24244,N_23636,N_23820);
nand U24245 (N_24245,N_23878,N_23535);
nor U24246 (N_24246,N_23958,N_23591);
nand U24247 (N_24247,N_23800,N_23807);
nor U24248 (N_24248,N_23532,N_23626);
xnor U24249 (N_24249,N_23706,N_23856);
or U24250 (N_24250,N_23938,N_23674);
xor U24251 (N_24251,N_23676,N_23833);
xnor U24252 (N_24252,N_23807,N_23971);
nor U24253 (N_24253,N_23725,N_23654);
nand U24254 (N_24254,N_23661,N_23816);
or U24255 (N_24255,N_23691,N_23965);
nor U24256 (N_24256,N_23734,N_23982);
xnor U24257 (N_24257,N_23689,N_23833);
nor U24258 (N_24258,N_23904,N_23566);
and U24259 (N_24259,N_23979,N_23827);
xor U24260 (N_24260,N_23511,N_23807);
or U24261 (N_24261,N_23767,N_23847);
xor U24262 (N_24262,N_23685,N_23958);
xnor U24263 (N_24263,N_23824,N_23640);
nand U24264 (N_24264,N_23814,N_23668);
xnor U24265 (N_24265,N_23559,N_23612);
or U24266 (N_24266,N_23525,N_23916);
nor U24267 (N_24267,N_23999,N_23960);
xnor U24268 (N_24268,N_23627,N_23523);
nand U24269 (N_24269,N_23991,N_23849);
xor U24270 (N_24270,N_23831,N_23982);
nor U24271 (N_24271,N_23617,N_23772);
xnor U24272 (N_24272,N_23564,N_23827);
nand U24273 (N_24273,N_23548,N_23732);
nand U24274 (N_24274,N_23915,N_23887);
nand U24275 (N_24275,N_23784,N_23734);
or U24276 (N_24276,N_23871,N_23633);
or U24277 (N_24277,N_23783,N_23509);
nor U24278 (N_24278,N_23967,N_23995);
xnor U24279 (N_24279,N_23965,N_23848);
or U24280 (N_24280,N_23778,N_23590);
and U24281 (N_24281,N_23771,N_23887);
nor U24282 (N_24282,N_23733,N_23617);
xnor U24283 (N_24283,N_23610,N_23674);
xor U24284 (N_24284,N_23894,N_23992);
nand U24285 (N_24285,N_23942,N_23882);
or U24286 (N_24286,N_23934,N_23916);
nor U24287 (N_24287,N_23995,N_23615);
nor U24288 (N_24288,N_23760,N_23709);
nand U24289 (N_24289,N_23807,N_23923);
or U24290 (N_24290,N_23540,N_23908);
or U24291 (N_24291,N_23791,N_23746);
nor U24292 (N_24292,N_23510,N_23555);
nand U24293 (N_24293,N_23847,N_23943);
and U24294 (N_24294,N_23912,N_23539);
or U24295 (N_24295,N_23711,N_23983);
and U24296 (N_24296,N_23622,N_23871);
nor U24297 (N_24297,N_23500,N_23971);
xnor U24298 (N_24298,N_23798,N_23983);
nor U24299 (N_24299,N_23626,N_23801);
and U24300 (N_24300,N_23561,N_23845);
or U24301 (N_24301,N_23921,N_23680);
and U24302 (N_24302,N_23519,N_23685);
and U24303 (N_24303,N_23563,N_23704);
xor U24304 (N_24304,N_23819,N_23668);
or U24305 (N_24305,N_23537,N_23603);
xor U24306 (N_24306,N_23850,N_23782);
and U24307 (N_24307,N_23961,N_23959);
or U24308 (N_24308,N_23936,N_23626);
or U24309 (N_24309,N_23555,N_23734);
nand U24310 (N_24310,N_23645,N_23723);
or U24311 (N_24311,N_23901,N_23626);
or U24312 (N_24312,N_23918,N_23660);
nor U24313 (N_24313,N_23702,N_23752);
nor U24314 (N_24314,N_23852,N_23866);
xor U24315 (N_24315,N_23855,N_23681);
xnor U24316 (N_24316,N_23818,N_23914);
and U24317 (N_24317,N_23993,N_23626);
nand U24318 (N_24318,N_23799,N_23662);
nand U24319 (N_24319,N_23532,N_23888);
nand U24320 (N_24320,N_23725,N_23969);
nand U24321 (N_24321,N_23644,N_23715);
or U24322 (N_24322,N_23594,N_23852);
or U24323 (N_24323,N_23522,N_23885);
or U24324 (N_24324,N_23791,N_23939);
xnor U24325 (N_24325,N_23901,N_23874);
xnor U24326 (N_24326,N_23754,N_23766);
xor U24327 (N_24327,N_23781,N_23715);
xnor U24328 (N_24328,N_23804,N_23622);
or U24329 (N_24329,N_23911,N_23893);
nor U24330 (N_24330,N_23609,N_23967);
and U24331 (N_24331,N_23986,N_23635);
or U24332 (N_24332,N_23725,N_23515);
xnor U24333 (N_24333,N_23509,N_23626);
and U24334 (N_24334,N_23885,N_23567);
nand U24335 (N_24335,N_23871,N_23978);
or U24336 (N_24336,N_23588,N_23911);
nor U24337 (N_24337,N_23730,N_23818);
xor U24338 (N_24338,N_23581,N_23529);
nor U24339 (N_24339,N_23525,N_23887);
nor U24340 (N_24340,N_23511,N_23936);
nor U24341 (N_24341,N_23558,N_23553);
and U24342 (N_24342,N_23836,N_23542);
and U24343 (N_24343,N_23577,N_23588);
or U24344 (N_24344,N_23805,N_23722);
or U24345 (N_24345,N_23773,N_23560);
or U24346 (N_24346,N_23929,N_23920);
or U24347 (N_24347,N_23894,N_23631);
or U24348 (N_24348,N_23646,N_23949);
nor U24349 (N_24349,N_23873,N_23697);
nand U24350 (N_24350,N_23749,N_23729);
xnor U24351 (N_24351,N_23939,N_23570);
or U24352 (N_24352,N_23694,N_23885);
nand U24353 (N_24353,N_23798,N_23878);
nand U24354 (N_24354,N_23899,N_23640);
nor U24355 (N_24355,N_23773,N_23890);
or U24356 (N_24356,N_23593,N_23981);
or U24357 (N_24357,N_23697,N_23728);
and U24358 (N_24358,N_23893,N_23690);
and U24359 (N_24359,N_23776,N_23758);
nand U24360 (N_24360,N_23641,N_23539);
or U24361 (N_24361,N_23824,N_23555);
or U24362 (N_24362,N_23610,N_23512);
xnor U24363 (N_24363,N_23881,N_23869);
nand U24364 (N_24364,N_23804,N_23908);
nand U24365 (N_24365,N_23964,N_23908);
nand U24366 (N_24366,N_23563,N_23681);
xor U24367 (N_24367,N_23946,N_23676);
nor U24368 (N_24368,N_23817,N_23684);
xor U24369 (N_24369,N_23591,N_23603);
or U24370 (N_24370,N_23712,N_23906);
or U24371 (N_24371,N_23822,N_23695);
or U24372 (N_24372,N_23743,N_23883);
or U24373 (N_24373,N_23521,N_23931);
and U24374 (N_24374,N_23907,N_23568);
nand U24375 (N_24375,N_23560,N_23782);
and U24376 (N_24376,N_23689,N_23537);
and U24377 (N_24377,N_23820,N_23680);
xnor U24378 (N_24378,N_23869,N_23904);
nor U24379 (N_24379,N_23889,N_23944);
or U24380 (N_24380,N_23885,N_23516);
nor U24381 (N_24381,N_23977,N_23872);
nor U24382 (N_24382,N_23992,N_23811);
or U24383 (N_24383,N_23600,N_23503);
or U24384 (N_24384,N_23915,N_23692);
and U24385 (N_24385,N_23633,N_23679);
xnor U24386 (N_24386,N_23800,N_23702);
and U24387 (N_24387,N_23791,N_23516);
or U24388 (N_24388,N_23759,N_23838);
xnor U24389 (N_24389,N_23712,N_23534);
nand U24390 (N_24390,N_23703,N_23596);
or U24391 (N_24391,N_23766,N_23614);
nor U24392 (N_24392,N_23910,N_23678);
xor U24393 (N_24393,N_23879,N_23602);
or U24394 (N_24394,N_23535,N_23694);
and U24395 (N_24395,N_23587,N_23647);
nor U24396 (N_24396,N_23692,N_23889);
nor U24397 (N_24397,N_23747,N_23938);
nand U24398 (N_24398,N_23967,N_23721);
and U24399 (N_24399,N_23991,N_23525);
nand U24400 (N_24400,N_23564,N_23673);
and U24401 (N_24401,N_23684,N_23884);
or U24402 (N_24402,N_23637,N_23892);
xnor U24403 (N_24403,N_23536,N_23983);
and U24404 (N_24404,N_23639,N_23921);
and U24405 (N_24405,N_23740,N_23630);
and U24406 (N_24406,N_23901,N_23951);
nor U24407 (N_24407,N_23665,N_23979);
nand U24408 (N_24408,N_23883,N_23605);
xor U24409 (N_24409,N_23537,N_23913);
and U24410 (N_24410,N_23596,N_23752);
and U24411 (N_24411,N_23638,N_23772);
nor U24412 (N_24412,N_23637,N_23749);
nor U24413 (N_24413,N_23832,N_23866);
nand U24414 (N_24414,N_23727,N_23845);
nand U24415 (N_24415,N_23736,N_23876);
or U24416 (N_24416,N_23630,N_23915);
and U24417 (N_24417,N_23793,N_23787);
or U24418 (N_24418,N_23742,N_23965);
nor U24419 (N_24419,N_23811,N_23803);
and U24420 (N_24420,N_23847,N_23979);
nand U24421 (N_24421,N_23828,N_23706);
xor U24422 (N_24422,N_23601,N_23776);
nand U24423 (N_24423,N_23988,N_23862);
nor U24424 (N_24424,N_23714,N_23618);
and U24425 (N_24425,N_23826,N_23670);
xnor U24426 (N_24426,N_23911,N_23751);
or U24427 (N_24427,N_23884,N_23740);
and U24428 (N_24428,N_23843,N_23856);
nand U24429 (N_24429,N_23824,N_23734);
nand U24430 (N_24430,N_23953,N_23977);
or U24431 (N_24431,N_23653,N_23897);
xor U24432 (N_24432,N_23716,N_23730);
and U24433 (N_24433,N_23800,N_23904);
nand U24434 (N_24434,N_23990,N_23581);
and U24435 (N_24435,N_23861,N_23880);
and U24436 (N_24436,N_23784,N_23527);
nor U24437 (N_24437,N_23925,N_23727);
and U24438 (N_24438,N_23787,N_23789);
xor U24439 (N_24439,N_23809,N_23661);
nand U24440 (N_24440,N_23957,N_23694);
and U24441 (N_24441,N_23802,N_23744);
or U24442 (N_24442,N_23757,N_23570);
xor U24443 (N_24443,N_23641,N_23596);
nor U24444 (N_24444,N_23545,N_23516);
nor U24445 (N_24445,N_23556,N_23571);
nand U24446 (N_24446,N_23864,N_23559);
nor U24447 (N_24447,N_23719,N_23912);
nor U24448 (N_24448,N_23896,N_23842);
xor U24449 (N_24449,N_23857,N_23755);
or U24450 (N_24450,N_23989,N_23719);
nor U24451 (N_24451,N_23684,N_23986);
xor U24452 (N_24452,N_23674,N_23770);
xor U24453 (N_24453,N_23972,N_23598);
or U24454 (N_24454,N_23701,N_23909);
nand U24455 (N_24455,N_23636,N_23862);
or U24456 (N_24456,N_23820,N_23666);
xor U24457 (N_24457,N_23980,N_23704);
or U24458 (N_24458,N_23985,N_23923);
and U24459 (N_24459,N_23730,N_23869);
and U24460 (N_24460,N_23705,N_23796);
nor U24461 (N_24461,N_23789,N_23823);
nor U24462 (N_24462,N_23960,N_23784);
or U24463 (N_24463,N_23974,N_23577);
nand U24464 (N_24464,N_23995,N_23815);
or U24465 (N_24465,N_23577,N_23657);
xor U24466 (N_24466,N_23750,N_23990);
nand U24467 (N_24467,N_23652,N_23837);
xor U24468 (N_24468,N_23927,N_23801);
or U24469 (N_24469,N_23780,N_23717);
or U24470 (N_24470,N_23991,N_23663);
nand U24471 (N_24471,N_23848,N_23748);
and U24472 (N_24472,N_23868,N_23522);
or U24473 (N_24473,N_23505,N_23524);
xor U24474 (N_24474,N_23925,N_23549);
or U24475 (N_24475,N_23906,N_23650);
nor U24476 (N_24476,N_23543,N_23766);
nor U24477 (N_24477,N_23634,N_23885);
or U24478 (N_24478,N_23916,N_23752);
and U24479 (N_24479,N_23876,N_23828);
or U24480 (N_24480,N_23981,N_23768);
or U24481 (N_24481,N_23516,N_23573);
nor U24482 (N_24482,N_23871,N_23663);
and U24483 (N_24483,N_23887,N_23904);
and U24484 (N_24484,N_23975,N_23577);
xnor U24485 (N_24485,N_23565,N_23663);
and U24486 (N_24486,N_23740,N_23928);
xnor U24487 (N_24487,N_23624,N_23804);
xnor U24488 (N_24488,N_23569,N_23981);
or U24489 (N_24489,N_23693,N_23619);
xnor U24490 (N_24490,N_23991,N_23657);
nand U24491 (N_24491,N_23594,N_23747);
nand U24492 (N_24492,N_23699,N_23739);
and U24493 (N_24493,N_23910,N_23746);
xor U24494 (N_24494,N_23948,N_23877);
or U24495 (N_24495,N_23807,N_23556);
or U24496 (N_24496,N_23868,N_23602);
xnor U24497 (N_24497,N_23681,N_23577);
and U24498 (N_24498,N_23826,N_23838);
and U24499 (N_24499,N_23571,N_23854);
and U24500 (N_24500,N_24443,N_24046);
nor U24501 (N_24501,N_24181,N_24036);
or U24502 (N_24502,N_24496,N_24396);
nand U24503 (N_24503,N_24077,N_24261);
xnor U24504 (N_24504,N_24149,N_24017);
and U24505 (N_24505,N_24198,N_24008);
and U24506 (N_24506,N_24083,N_24402);
nor U24507 (N_24507,N_24400,N_24466);
nand U24508 (N_24508,N_24241,N_24469);
nand U24509 (N_24509,N_24197,N_24015);
or U24510 (N_24510,N_24043,N_24338);
nor U24511 (N_24511,N_24055,N_24356);
xnor U24512 (N_24512,N_24134,N_24244);
or U24513 (N_24513,N_24052,N_24206);
xor U24514 (N_24514,N_24401,N_24139);
nor U24515 (N_24515,N_24119,N_24141);
nand U24516 (N_24516,N_24025,N_24367);
and U24517 (N_24517,N_24259,N_24078);
nor U24518 (N_24518,N_24175,N_24231);
nor U24519 (N_24519,N_24373,N_24242);
xnor U24520 (N_24520,N_24132,N_24263);
or U24521 (N_24521,N_24449,N_24014);
nand U24522 (N_24522,N_24107,N_24344);
xnor U24523 (N_24523,N_24153,N_24359);
xor U24524 (N_24524,N_24349,N_24062);
and U24525 (N_24525,N_24194,N_24346);
and U24526 (N_24526,N_24044,N_24376);
nand U24527 (N_24527,N_24113,N_24184);
nand U24528 (N_24528,N_24022,N_24486);
nor U24529 (N_24529,N_24236,N_24411);
or U24530 (N_24530,N_24410,N_24387);
or U24531 (N_24531,N_24016,N_24092);
and U24532 (N_24532,N_24066,N_24316);
and U24533 (N_24533,N_24024,N_24032);
or U24534 (N_24534,N_24110,N_24326);
or U24535 (N_24535,N_24247,N_24438);
xor U24536 (N_24536,N_24436,N_24164);
nor U24537 (N_24537,N_24255,N_24380);
nand U24538 (N_24538,N_24151,N_24423);
xor U24539 (N_24539,N_24268,N_24461);
nand U24540 (N_24540,N_24470,N_24243);
nand U24541 (N_24541,N_24393,N_24390);
nor U24542 (N_24542,N_24398,N_24005);
and U24543 (N_24543,N_24204,N_24442);
or U24544 (N_24544,N_24127,N_24234);
and U24545 (N_24545,N_24317,N_24130);
nor U24546 (N_24546,N_24477,N_24147);
nand U24547 (N_24547,N_24214,N_24389);
nand U24548 (N_24548,N_24311,N_24002);
nor U24549 (N_24549,N_24099,N_24200);
and U24550 (N_24550,N_24224,N_24122);
nand U24551 (N_24551,N_24416,N_24215);
and U24552 (N_24552,N_24421,N_24383);
xor U24553 (N_24553,N_24456,N_24170);
nand U24554 (N_24554,N_24281,N_24100);
nand U24555 (N_24555,N_24179,N_24125);
nor U24556 (N_24556,N_24260,N_24330);
nand U24557 (N_24557,N_24051,N_24493);
xor U24558 (N_24558,N_24286,N_24165);
and U24559 (N_24559,N_24394,N_24209);
nand U24560 (N_24560,N_24150,N_24483);
nor U24561 (N_24561,N_24156,N_24365);
nand U24562 (N_24562,N_24405,N_24121);
or U24563 (N_24563,N_24427,N_24068);
or U24564 (N_24564,N_24207,N_24135);
xor U24565 (N_24565,N_24013,N_24295);
and U24566 (N_24566,N_24497,N_24377);
nor U24567 (N_24567,N_24293,N_24277);
xor U24568 (N_24568,N_24291,N_24348);
or U24569 (N_24569,N_24126,N_24187);
nand U24570 (N_24570,N_24182,N_24351);
and U24571 (N_24571,N_24391,N_24045);
and U24572 (N_24572,N_24308,N_24345);
nor U24573 (N_24573,N_24482,N_24357);
or U24574 (N_24574,N_24120,N_24418);
and U24575 (N_24575,N_24303,N_24065);
or U24576 (N_24576,N_24446,N_24428);
xor U24577 (N_24577,N_24103,N_24167);
nor U24578 (N_24578,N_24090,N_24142);
or U24579 (N_24579,N_24307,N_24169);
or U24580 (N_24580,N_24274,N_24315);
or U24581 (N_24581,N_24334,N_24434);
nor U24582 (N_24582,N_24350,N_24414);
nand U24583 (N_24583,N_24007,N_24392);
and U24584 (N_24584,N_24484,N_24371);
nand U24585 (N_24585,N_24091,N_24161);
and U24586 (N_24586,N_24035,N_24288);
xnor U24587 (N_24587,N_24202,N_24094);
nor U24588 (N_24588,N_24074,N_24028);
and U24589 (N_24589,N_24180,N_24228);
nor U24590 (N_24590,N_24408,N_24314);
nand U24591 (N_24591,N_24223,N_24254);
xor U24592 (N_24592,N_24395,N_24030);
nand U24593 (N_24593,N_24447,N_24407);
or U24594 (N_24594,N_24148,N_24249);
and U24595 (N_24595,N_24220,N_24088);
xnor U24596 (N_24596,N_24026,N_24257);
xor U24597 (N_24597,N_24105,N_24429);
nor U24598 (N_24598,N_24245,N_24384);
and U24599 (N_24599,N_24431,N_24319);
or U24600 (N_24600,N_24335,N_24041);
xnor U24601 (N_24601,N_24189,N_24485);
and U24602 (N_24602,N_24325,N_24108);
nor U24603 (N_24603,N_24152,N_24409);
nor U24604 (N_24604,N_24232,N_24102);
xnor U24605 (N_24605,N_24454,N_24304);
nand U24606 (N_24606,N_24240,N_24101);
nand U24607 (N_24607,N_24048,N_24208);
and U24608 (N_24608,N_24491,N_24458);
nand U24609 (N_24609,N_24467,N_24494);
or U24610 (N_24610,N_24087,N_24118);
nor U24611 (N_24611,N_24489,N_24333);
nor U24612 (N_24612,N_24219,N_24069);
or U24613 (N_24613,N_24131,N_24355);
and U24614 (N_24614,N_24217,N_24372);
xor U24615 (N_24615,N_24019,N_24027);
nor U24616 (N_24616,N_24448,N_24282);
or U24617 (N_24617,N_24269,N_24265);
nand U24618 (N_24618,N_24321,N_24210);
nand U24619 (N_24619,N_24339,N_24374);
nor U24620 (N_24620,N_24342,N_24138);
xor U24621 (N_24621,N_24341,N_24237);
or U24622 (N_24622,N_24264,N_24067);
xor U24623 (N_24623,N_24085,N_24270);
xnor U24624 (N_24624,N_24424,N_24474);
nand U24625 (N_24625,N_24106,N_24363);
or U24626 (N_24626,N_24413,N_24111);
nor U24627 (N_24627,N_24283,N_24271);
and U24628 (N_24628,N_24299,N_24306);
nor U24629 (N_24629,N_24347,N_24453);
or U24630 (N_24630,N_24001,N_24322);
nand U24631 (N_24631,N_24011,N_24034);
nor U24632 (N_24632,N_24312,N_24188);
and U24633 (N_24633,N_24309,N_24370);
nand U24634 (N_24634,N_24495,N_24163);
nor U24635 (N_24635,N_24463,N_24415);
nand U24636 (N_24636,N_24213,N_24327);
xnor U24637 (N_24637,N_24476,N_24227);
xor U24638 (N_24638,N_24272,N_24487);
nor U24639 (N_24639,N_24058,N_24129);
nor U24640 (N_24640,N_24479,N_24440);
and U24641 (N_24641,N_24352,N_24399);
nor U24642 (N_24642,N_24262,N_24337);
nor U24643 (N_24643,N_24133,N_24221);
and U24644 (N_24644,N_24313,N_24451);
nand U24645 (N_24645,N_24294,N_24042);
xnor U24646 (N_24646,N_24060,N_24287);
and U24647 (N_24647,N_24117,N_24258);
or U24648 (N_24648,N_24097,N_24093);
nand U24649 (N_24649,N_24124,N_24379);
xor U24650 (N_24650,N_24279,N_24137);
and U24651 (N_24651,N_24465,N_24278);
nand U24652 (N_24652,N_24095,N_24292);
xnor U24653 (N_24653,N_24080,N_24144);
nand U24654 (N_24654,N_24166,N_24499);
nor U24655 (N_24655,N_24158,N_24444);
and U24656 (N_24656,N_24201,N_24071);
nor U24657 (N_24657,N_24433,N_24238);
and U24658 (N_24658,N_24039,N_24471);
xor U24659 (N_24659,N_24455,N_24049);
or U24660 (N_24660,N_24381,N_24056);
nor U24661 (N_24661,N_24037,N_24109);
nor U24662 (N_24662,N_24146,N_24353);
nor U24663 (N_24663,N_24432,N_24439);
and U24664 (N_24664,N_24490,N_24004);
or U24665 (N_24665,N_24225,N_24128);
nand U24666 (N_24666,N_24323,N_24403);
nor U24667 (N_24667,N_24155,N_24426);
nand U24668 (N_24668,N_24366,N_24233);
xnor U24669 (N_24669,N_24115,N_24369);
or U24670 (N_24670,N_24360,N_24251);
or U24671 (N_24671,N_24089,N_24159);
xnor U24672 (N_24672,N_24140,N_24437);
and U24673 (N_24673,N_24266,N_24072);
xnor U24674 (N_24674,N_24226,N_24218);
or U24675 (N_24675,N_24445,N_24143);
nor U24676 (N_24676,N_24003,N_24112);
and U24677 (N_24677,N_24116,N_24230);
nand U24678 (N_24678,N_24375,N_24253);
nor U24679 (N_24679,N_24297,N_24123);
xnor U24680 (N_24680,N_24481,N_24450);
nand U24681 (N_24681,N_24000,N_24084);
nand U24682 (N_24682,N_24250,N_24193);
xnor U24683 (N_24683,N_24435,N_24033);
nor U24684 (N_24684,N_24073,N_24050);
and U24685 (N_24685,N_24211,N_24404);
and U24686 (N_24686,N_24229,N_24362);
xnor U24687 (N_24687,N_24192,N_24075);
and U24688 (N_24688,N_24098,N_24488);
nand U24689 (N_24689,N_24205,N_24063);
xnor U24690 (N_24690,N_24320,N_24070);
and U24691 (N_24691,N_24079,N_24328);
and U24692 (N_24692,N_24464,N_24047);
xnor U24693 (N_24693,N_24388,N_24196);
or U24694 (N_24694,N_24441,N_24305);
and U24695 (N_24695,N_24006,N_24267);
xnor U24696 (N_24696,N_24364,N_24290);
nand U24697 (N_24697,N_24023,N_24478);
nor U24698 (N_24698,N_24178,N_24480);
xor U24699 (N_24699,N_24329,N_24252);
nand U24700 (N_24700,N_24324,N_24186);
or U24701 (N_24701,N_24368,N_24385);
nor U24702 (N_24702,N_24457,N_24216);
nor U24703 (N_24703,N_24177,N_24472);
xor U24704 (N_24704,N_24459,N_24212);
or U24705 (N_24705,N_24195,N_24104);
or U24706 (N_24706,N_24061,N_24280);
nand U24707 (N_24707,N_24289,N_24419);
nor U24708 (N_24708,N_24298,N_24029);
and U24709 (N_24709,N_24012,N_24021);
xnor U24710 (N_24710,N_24302,N_24275);
or U24711 (N_24711,N_24276,N_24331);
and U24712 (N_24712,N_24343,N_24336);
and U24713 (N_24713,N_24386,N_24154);
nor U24714 (N_24714,N_24081,N_24301);
nor U24715 (N_24715,N_24422,N_24246);
nor U24716 (N_24716,N_24018,N_24492);
xnor U24717 (N_24717,N_24300,N_24176);
nor U24718 (N_24718,N_24190,N_24114);
or U24719 (N_24719,N_24256,N_24172);
and U24720 (N_24720,N_24010,N_24222);
nor U24721 (N_24721,N_24064,N_24199);
xor U24722 (N_24722,N_24054,N_24358);
nor U24723 (N_24723,N_24168,N_24038);
nand U24724 (N_24724,N_24406,N_24340);
nand U24725 (N_24725,N_24475,N_24473);
xor U24726 (N_24726,N_24318,N_24031);
xnor U24727 (N_24727,N_24332,N_24361);
nor U24728 (N_24728,N_24171,N_24053);
nand U24729 (N_24729,N_24203,N_24160);
or U24730 (N_24730,N_24412,N_24378);
nand U24731 (N_24731,N_24162,N_24183);
xor U24732 (N_24732,N_24076,N_24430);
nor U24733 (N_24733,N_24157,N_24310);
or U24734 (N_24734,N_24452,N_24284);
xor U24735 (N_24735,N_24239,N_24136);
nand U24736 (N_24736,N_24057,N_24460);
nor U24737 (N_24737,N_24354,N_24273);
and U24738 (N_24738,N_24235,N_24173);
nand U24739 (N_24739,N_24382,N_24174);
nor U24740 (N_24740,N_24417,N_24145);
or U24741 (N_24741,N_24397,N_24086);
or U24742 (N_24742,N_24468,N_24248);
xnor U24743 (N_24743,N_24020,N_24191);
and U24744 (N_24744,N_24420,N_24285);
or U24745 (N_24745,N_24462,N_24096);
nand U24746 (N_24746,N_24185,N_24059);
xor U24747 (N_24747,N_24498,N_24296);
xnor U24748 (N_24748,N_24082,N_24040);
or U24749 (N_24749,N_24009,N_24425);
and U24750 (N_24750,N_24165,N_24085);
nand U24751 (N_24751,N_24248,N_24069);
xnor U24752 (N_24752,N_24188,N_24441);
nor U24753 (N_24753,N_24348,N_24083);
nand U24754 (N_24754,N_24187,N_24334);
or U24755 (N_24755,N_24043,N_24082);
xor U24756 (N_24756,N_24402,N_24154);
or U24757 (N_24757,N_24144,N_24150);
or U24758 (N_24758,N_24330,N_24112);
nor U24759 (N_24759,N_24371,N_24494);
xnor U24760 (N_24760,N_24173,N_24063);
or U24761 (N_24761,N_24405,N_24471);
xnor U24762 (N_24762,N_24133,N_24095);
nor U24763 (N_24763,N_24174,N_24403);
nand U24764 (N_24764,N_24357,N_24313);
xnor U24765 (N_24765,N_24383,N_24125);
nor U24766 (N_24766,N_24375,N_24066);
and U24767 (N_24767,N_24053,N_24360);
xnor U24768 (N_24768,N_24126,N_24245);
or U24769 (N_24769,N_24315,N_24097);
nand U24770 (N_24770,N_24368,N_24088);
or U24771 (N_24771,N_24041,N_24000);
or U24772 (N_24772,N_24338,N_24025);
or U24773 (N_24773,N_24207,N_24242);
and U24774 (N_24774,N_24215,N_24347);
or U24775 (N_24775,N_24218,N_24114);
nand U24776 (N_24776,N_24414,N_24145);
or U24777 (N_24777,N_24375,N_24148);
nor U24778 (N_24778,N_24368,N_24242);
nor U24779 (N_24779,N_24166,N_24225);
and U24780 (N_24780,N_24269,N_24225);
and U24781 (N_24781,N_24290,N_24207);
nand U24782 (N_24782,N_24348,N_24020);
or U24783 (N_24783,N_24169,N_24025);
or U24784 (N_24784,N_24223,N_24181);
and U24785 (N_24785,N_24318,N_24491);
and U24786 (N_24786,N_24068,N_24438);
nand U24787 (N_24787,N_24288,N_24475);
and U24788 (N_24788,N_24149,N_24215);
or U24789 (N_24789,N_24478,N_24142);
nor U24790 (N_24790,N_24224,N_24041);
and U24791 (N_24791,N_24296,N_24138);
or U24792 (N_24792,N_24164,N_24016);
xor U24793 (N_24793,N_24001,N_24405);
and U24794 (N_24794,N_24081,N_24487);
nor U24795 (N_24795,N_24118,N_24225);
or U24796 (N_24796,N_24304,N_24413);
or U24797 (N_24797,N_24258,N_24128);
nor U24798 (N_24798,N_24219,N_24195);
or U24799 (N_24799,N_24223,N_24091);
or U24800 (N_24800,N_24349,N_24347);
nor U24801 (N_24801,N_24034,N_24256);
and U24802 (N_24802,N_24334,N_24173);
and U24803 (N_24803,N_24464,N_24059);
xor U24804 (N_24804,N_24001,N_24092);
nor U24805 (N_24805,N_24078,N_24323);
and U24806 (N_24806,N_24086,N_24387);
nand U24807 (N_24807,N_24491,N_24051);
nor U24808 (N_24808,N_24133,N_24245);
nor U24809 (N_24809,N_24011,N_24266);
nand U24810 (N_24810,N_24359,N_24419);
xnor U24811 (N_24811,N_24402,N_24455);
and U24812 (N_24812,N_24359,N_24117);
nand U24813 (N_24813,N_24146,N_24463);
nand U24814 (N_24814,N_24117,N_24003);
nand U24815 (N_24815,N_24436,N_24272);
xor U24816 (N_24816,N_24415,N_24008);
nand U24817 (N_24817,N_24257,N_24478);
or U24818 (N_24818,N_24105,N_24256);
and U24819 (N_24819,N_24117,N_24288);
nand U24820 (N_24820,N_24124,N_24218);
nand U24821 (N_24821,N_24116,N_24292);
nor U24822 (N_24822,N_24334,N_24024);
xnor U24823 (N_24823,N_24171,N_24413);
nand U24824 (N_24824,N_24410,N_24110);
nor U24825 (N_24825,N_24420,N_24111);
nor U24826 (N_24826,N_24142,N_24355);
and U24827 (N_24827,N_24179,N_24134);
and U24828 (N_24828,N_24251,N_24092);
and U24829 (N_24829,N_24234,N_24369);
nand U24830 (N_24830,N_24309,N_24221);
nor U24831 (N_24831,N_24097,N_24106);
or U24832 (N_24832,N_24136,N_24234);
nand U24833 (N_24833,N_24302,N_24444);
xor U24834 (N_24834,N_24441,N_24337);
and U24835 (N_24835,N_24037,N_24366);
and U24836 (N_24836,N_24435,N_24037);
xor U24837 (N_24837,N_24169,N_24045);
xnor U24838 (N_24838,N_24247,N_24415);
and U24839 (N_24839,N_24356,N_24174);
xnor U24840 (N_24840,N_24192,N_24024);
nand U24841 (N_24841,N_24178,N_24186);
nor U24842 (N_24842,N_24416,N_24116);
xor U24843 (N_24843,N_24030,N_24418);
nor U24844 (N_24844,N_24048,N_24113);
and U24845 (N_24845,N_24446,N_24206);
or U24846 (N_24846,N_24268,N_24069);
or U24847 (N_24847,N_24426,N_24238);
or U24848 (N_24848,N_24205,N_24214);
xor U24849 (N_24849,N_24382,N_24485);
and U24850 (N_24850,N_24184,N_24170);
nand U24851 (N_24851,N_24038,N_24232);
nor U24852 (N_24852,N_24479,N_24242);
or U24853 (N_24853,N_24340,N_24320);
or U24854 (N_24854,N_24251,N_24378);
nand U24855 (N_24855,N_24239,N_24280);
nor U24856 (N_24856,N_24343,N_24457);
nor U24857 (N_24857,N_24321,N_24138);
or U24858 (N_24858,N_24049,N_24044);
and U24859 (N_24859,N_24358,N_24012);
nor U24860 (N_24860,N_24169,N_24460);
and U24861 (N_24861,N_24010,N_24143);
nand U24862 (N_24862,N_24136,N_24078);
nand U24863 (N_24863,N_24055,N_24013);
nand U24864 (N_24864,N_24012,N_24476);
xnor U24865 (N_24865,N_24419,N_24163);
and U24866 (N_24866,N_24053,N_24155);
or U24867 (N_24867,N_24355,N_24001);
xnor U24868 (N_24868,N_24406,N_24086);
nor U24869 (N_24869,N_24358,N_24409);
nor U24870 (N_24870,N_24399,N_24284);
or U24871 (N_24871,N_24308,N_24441);
or U24872 (N_24872,N_24419,N_24245);
xnor U24873 (N_24873,N_24402,N_24267);
and U24874 (N_24874,N_24316,N_24030);
xnor U24875 (N_24875,N_24465,N_24195);
nand U24876 (N_24876,N_24144,N_24155);
nand U24877 (N_24877,N_24097,N_24025);
or U24878 (N_24878,N_24211,N_24403);
and U24879 (N_24879,N_24111,N_24406);
nor U24880 (N_24880,N_24484,N_24027);
nor U24881 (N_24881,N_24459,N_24211);
or U24882 (N_24882,N_24086,N_24396);
and U24883 (N_24883,N_24389,N_24051);
or U24884 (N_24884,N_24334,N_24312);
nor U24885 (N_24885,N_24088,N_24038);
or U24886 (N_24886,N_24041,N_24125);
xnor U24887 (N_24887,N_24355,N_24257);
nor U24888 (N_24888,N_24309,N_24231);
nand U24889 (N_24889,N_24270,N_24031);
nand U24890 (N_24890,N_24079,N_24128);
nor U24891 (N_24891,N_24450,N_24471);
nor U24892 (N_24892,N_24138,N_24024);
nand U24893 (N_24893,N_24440,N_24476);
nand U24894 (N_24894,N_24451,N_24256);
and U24895 (N_24895,N_24018,N_24365);
xor U24896 (N_24896,N_24178,N_24499);
nor U24897 (N_24897,N_24150,N_24164);
nand U24898 (N_24898,N_24294,N_24069);
nor U24899 (N_24899,N_24056,N_24284);
and U24900 (N_24900,N_24492,N_24409);
nor U24901 (N_24901,N_24041,N_24143);
or U24902 (N_24902,N_24223,N_24121);
or U24903 (N_24903,N_24275,N_24021);
xnor U24904 (N_24904,N_24026,N_24456);
nor U24905 (N_24905,N_24498,N_24127);
or U24906 (N_24906,N_24071,N_24346);
or U24907 (N_24907,N_24492,N_24060);
nand U24908 (N_24908,N_24218,N_24343);
xor U24909 (N_24909,N_24016,N_24250);
nand U24910 (N_24910,N_24296,N_24408);
and U24911 (N_24911,N_24011,N_24486);
and U24912 (N_24912,N_24343,N_24305);
or U24913 (N_24913,N_24443,N_24052);
xnor U24914 (N_24914,N_24435,N_24041);
nand U24915 (N_24915,N_24338,N_24311);
nor U24916 (N_24916,N_24353,N_24315);
and U24917 (N_24917,N_24336,N_24240);
or U24918 (N_24918,N_24397,N_24054);
nand U24919 (N_24919,N_24198,N_24147);
xnor U24920 (N_24920,N_24481,N_24384);
nor U24921 (N_24921,N_24283,N_24450);
or U24922 (N_24922,N_24372,N_24040);
nor U24923 (N_24923,N_24473,N_24288);
or U24924 (N_24924,N_24034,N_24145);
xnor U24925 (N_24925,N_24104,N_24027);
xnor U24926 (N_24926,N_24276,N_24089);
and U24927 (N_24927,N_24334,N_24333);
and U24928 (N_24928,N_24170,N_24299);
or U24929 (N_24929,N_24360,N_24202);
xnor U24930 (N_24930,N_24242,N_24153);
xnor U24931 (N_24931,N_24353,N_24142);
xnor U24932 (N_24932,N_24311,N_24123);
and U24933 (N_24933,N_24146,N_24297);
nand U24934 (N_24934,N_24498,N_24240);
or U24935 (N_24935,N_24193,N_24212);
nand U24936 (N_24936,N_24094,N_24328);
or U24937 (N_24937,N_24443,N_24317);
and U24938 (N_24938,N_24465,N_24276);
nor U24939 (N_24939,N_24182,N_24337);
xnor U24940 (N_24940,N_24203,N_24251);
nand U24941 (N_24941,N_24403,N_24362);
nor U24942 (N_24942,N_24120,N_24056);
and U24943 (N_24943,N_24048,N_24175);
xnor U24944 (N_24944,N_24180,N_24114);
xnor U24945 (N_24945,N_24348,N_24232);
or U24946 (N_24946,N_24049,N_24432);
xnor U24947 (N_24947,N_24421,N_24304);
and U24948 (N_24948,N_24396,N_24030);
or U24949 (N_24949,N_24439,N_24177);
nand U24950 (N_24950,N_24452,N_24423);
xnor U24951 (N_24951,N_24122,N_24340);
nand U24952 (N_24952,N_24217,N_24367);
nor U24953 (N_24953,N_24255,N_24334);
nand U24954 (N_24954,N_24432,N_24119);
nand U24955 (N_24955,N_24094,N_24009);
or U24956 (N_24956,N_24312,N_24253);
or U24957 (N_24957,N_24159,N_24420);
and U24958 (N_24958,N_24162,N_24225);
or U24959 (N_24959,N_24034,N_24272);
nand U24960 (N_24960,N_24440,N_24135);
nand U24961 (N_24961,N_24197,N_24483);
or U24962 (N_24962,N_24249,N_24158);
xor U24963 (N_24963,N_24002,N_24198);
and U24964 (N_24964,N_24382,N_24436);
and U24965 (N_24965,N_24104,N_24312);
or U24966 (N_24966,N_24395,N_24331);
or U24967 (N_24967,N_24413,N_24057);
nand U24968 (N_24968,N_24129,N_24135);
nor U24969 (N_24969,N_24347,N_24345);
nor U24970 (N_24970,N_24113,N_24213);
or U24971 (N_24971,N_24479,N_24285);
xor U24972 (N_24972,N_24430,N_24497);
nor U24973 (N_24973,N_24446,N_24059);
nor U24974 (N_24974,N_24257,N_24328);
or U24975 (N_24975,N_24153,N_24323);
nor U24976 (N_24976,N_24207,N_24062);
and U24977 (N_24977,N_24438,N_24395);
nor U24978 (N_24978,N_24062,N_24099);
nand U24979 (N_24979,N_24177,N_24470);
and U24980 (N_24980,N_24203,N_24292);
or U24981 (N_24981,N_24474,N_24078);
nor U24982 (N_24982,N_24066,N_24279);
or U24983 (N_24983,N_24275,N_24283);
nand U24984 (N_24984,N_24064,N_24183);
nand U24985 (N_24985,N_24311,N_24406);
or U24986 (N_24986,N_24247,N_24262);
nor U24987 (N_24987,N_24353,N_24272);
nand U24988 (N_24988,N_24410,N_24427);
nor U24989 (N_24989,N_24195,N_24168);
xnor U24990 (N_24990,N_24207,N_24258);
nor U24991 (N_24991,N_24253,N_24453);
nand U24992 (N_24992,N_24219,N_24330);
nand U24993 (N_24993,N_24109,N_24179);
and U24994 (N_24994,N_24375,N_24091);
xor U24995 (N_24995,N_24005,N_24444);
or U24996 (N_24996,N_24299,N_24432);
nor U24997 (N_24997,N_24084,N_24154);
xor U24998 (N_24998,N_24256,N_24234);
nor U24999 (N_24999,N_24209,N_24023);
nand U25000 (N_25000,N_24656,N_24626);
xor U25001 (N_25001,N_24746,N_24562);
nand U25002 (N_25002,N_24581,N_24828);
xor U25003 (N_25003,N_24844,N_24769);
and U25004 (N_25004,N_24613,N_24852);
and U25005 (N_25005,N_24831,N_24723);
nor U25006 (N_25006,N_24735,N_24939);
and U25007 (N_25007,N_24505,N_24582);
or U25008 (N_25008,N_24540,N_24682);
nand U25009 (N_25009,N_24920,N_24619);
xor U25010 (N_25010,N_24830,N_24519);
xor U25011 (N_25011,N_24722,N_24817);
or U25012 (N_25012,N_24821,N_24923);
nor U25013 (N_25013,N_24694,N_24837);
or U25014 (N_25014,N_24739,N_24630);
nand U25015 (N_25015,N_24772,N_24861);
and U25016 (N_25016,N_24760,N_24534);
and U25017 (N_25017,N_24672,N_24584);
nand U25018 (N_25018,N_24840,N_24594);
and U25019 (N_25019,N_24745,N_24781);
or U25020 (N_25020,N_24738,N_24804);
nand U25021 (N_25021,N_24500,N_24707);
and U25022 (N_25022,N_24695,N_24839);
xnor U25023 (N_25023,N_24543,N_24848);
and U25024 (N_25024,N_24554,N_24508);
and U25025 (N_25025,N_24527,N_24668);
or U25026 (N_25026,N_24910,N_24614);
or U25027 (N_25027,N_24846,N_24687);
nor U25028 (N_25028,N_24522,N_24859);
and U25029 (N_25029,N_24531,N_24587);
nor U25030 (N_25030,N_24936,N_24615);
nor U25031 (N_25031,N_24697,N_24811);
nand U25032 (N_25032,N_24711,N_24820);
nand U25033 (N_25033,N_24756,N_24785);
nand U25034 (N_25034,N_24921,N_24970);
and U25035 (N_25035,N_24720,N_24749);
nor U25036 (N_25036,N_24663,N_24965);
or U25037 (N_25037,N_24693,N_24765);
or U25038 (N_25038,N_24547,N_24670);
nand U25039 (N_25039,N_24905,N_24546);
nand U25040 (N_25040,N_24602,N_24768);
xnor U25041 (N_25041,N_24692,N_24911);
and U25042 (N_25042,N_24868,N_24620);
nor U25043 (N_25043,N_24641,N_24872);
and U25044 (N_25044,N_24767,N_24561);
nand U25045 (N_25045,N_24690,N_24995);
nor U25046 (N_25046,N_24925,N_24747);
nand U25047 (N_25047,N_24841,N_24600);
and U25048 (N_25048,N_24887,N_24658);
or U25049 (N_25049,N_24754,N_24704);
nor U25050 (N_25050,N_24855,N_24703);
nor U25051 (N_25051,N_24625,N_24952);
and U25052 (N_25052,N_24974,N_24610);
nor U25053 (N_25053,N_24979,N_24509);
and U25054 (N_25054,N_24971,N_24570);
nor U25055 (N_25055,N_24706,N_24934);
or U25056 (N_25056,N_24753,N_24515);
nor U25057 (N_25057,N_24555,N_24778);
nand U25058 (N_25058,N_24764,N_24699);
xor U25059 (N_25059,N_24601,N_24964);
xor U25060 (N_25060,N_24624,N_24826);
nand U25061 (N_25061,N_24865,N_24973);
nand U25062 (N_25062,N_24871,N_24514);
xor U25063 (N_25063,N_24976,N_24933);
xnor U25064 (N_25064,N_24700,N_24617);
and U25065 (N_25065,N_24943,N_24884);
nand U25066 (N_25066,N_24962,N_24579);
and U25067 (N_25067,N_24511,N_24651);
and U25068 (N_25068,N_24535,N_24931);
xor U25069 (N_25069,N_24966,N_24771);
nand U25070 (N_25070,N_24565,N_24986);
or U25071 (N_25071,N_24633,N_24845);
and U25072 (N_25072,N_24988,N_24686);
or U25073 (N_25073,N_24913,N_24897);
nor U25074 (N_25074,N_24869,N_24850);
xnor U25075 (N_25075,N_24674,N_24843);
or U25076 (N_25076,N_24688,N_24585);
nand U25077 (N_25077,N_24816,N_24621);
and U25078 (N_25078,N_24894,N_24890);
xnor U25079 (N_25079,N_24637,N_24981);
and U25080 (N_25080,N_24542,N_24710);
or U25081 (N_25081,N_24780,N_24895);
nor U25082 (N_25082,N_24683,N_24583);
and U25083 (N_25083,N_24567,N_24676);
or U25084 (N_25084,N_24783,N_24740);
or U25085 (N_25085,N_24712,N_24533);
and U25086 (N_25086,N_24961,N_24792);
xnor U25087 (N_25087,N_24629,N_24824);
and U25088 (N_25088,N_24858,N_24608);
and U25089 (N_25089,N_24953,N_24571);
nor U25090 (N_25090,N_24516,N_24662);
or U25091 (N_25091,N_24959,N_24553);
nand U25092 (N_25092,N_24929,N_24501);
nand U25093 (N_25093,N_24551,N_24664);
nor U25094 (N_25094,N_24681,N_24715);
and U25095 (N_25095,N_24517,N_24597);
nor U25096 (N_25096,N_24901,N_24580);
xor U25097 (N_25097,N_24634,N_24560);
nand U25098 (N_25098,N_24812,N_24870);
and U25099 (N_25099,N_24654,N_24696);
or U25100 (N_25100,N_24725,N_24705);
or U25101 (N_25101,N_24940,N_24607);
nor U25102 (N_25102,N_24805,N_24724);
or U25103 (N_25103,N_24878,N_24822);
or U25104 (N_25104,N_24815,N_24963);
nand U25105 (N_25105,N_24667,N_24666);
and U25106 (N_25106,N_24853,N_24789);
and U25107 (N_25107,N_24829,N_24732);
nor U25108 (N_25108,N_24521,N_24906);
and U25109 (N_25109,N_24566,N_24525);
nand U25110 (N_25110,N_24854,N_24544);
xnor U25111 (N_25111,N_24713,N_24958);
and U25112 (N_25112,N_24969,N_24975);
xor U25113 (N_25113,N_24718,N_24537);
xnor U25114 (N_25114,N_24834,N_24680);
and U25115 (N_25115,N_24794,N_24759);
or U25116 (N_25116,N_24685,N_24838);
nand U25117 (N_25117,N_24532,N_24557);
or U25118 (N_25118,N_24796,N_24742);
nor U25119 (N_25119,N_24642,N_24698);
nand U25120 (N_25120,N_24717,N_24689);
and U25121 (N_25121,N_24653,N_24518);
nand U25122 (N_25122,N_24919,N_24918);
nand U25123 (N_25123,N_24708,N_24507);
or U25124 (N_25124,N_24847,N_24922);
and U25125 (N_25125,N_24675,N_24564);
or U25126 (N_25126,N_24591,N_24833);
or U25127 (N_25127,N_24889,N_24731);
xor U25128 (N_25128,N_24808,N_24504);
nand U25129 (N_25129,N_24892,N_24879);
xnor U25130 (N_25130,N_24999,N_24882);
nor U25131 (N_25131,N_24917,N_24665);
or U25132 (N_25132,N_24596,N_24604);
nand U25133 (N_25133,N_24823,N_24730);
or U25134 (N_25134,N_24590,N_24618);
nand U25135 (N_25135,N_24791,N_24631);
nand U25136 (N_25136,N_24548,N_24948);
or U25137 (N_25137,N_24795,N_24549);
and U25138 (N_25138,N_24636,N_24774);
and U25139 (N_25139,N_24721,N_24782);
xnor U25140 (N_25140,N_24528,N_24652);
xnor U25141 (N_25141,N_24748,N_24599);
and U25142 (N_25142,N_24763,N_24775);
nand U25143 (N_25143,N_24646,N_24661);
or U25144 (N_25144,N_24856,N_24716);
and U25145 (N_25145,N_24813,N_24803);
and U25146 (N_25146,N_24788,N_24526);
or U25147 (N_25147,N_24752,N_24737);
nand U25148 (N_25148,N_24744,N_24896);
xnor U25149 (N_25149,N_24524,N_24766);
or U25150 (N_25150,N_24776,N_24985);
or U25151 (N_25151,N_24891,N_24989);
and U25152 (N_25152,N_24773,N_24992);
nor U25153 (N_25153,N_24714,N_24874);
or U25154 (N_25154,N_24576,N_24678);
nand U25155 (N_25155,N_24942,N_24529);
or U25156 (N_25156,N_24593,N_24867);
nor U25157 (N_25157,N_24757,N_24762);
nand U25158 (N_25158,N_24734,N_24928);
nor U25159 (N_25159,N_24946,N_24603);
nand U25160 (N_25160,N_24941,N_24606);
xnor U25161 (N_25161,N_24914,N_24648);
nand U25162 (N_25162,N_24827,N_24558);
nor U25163 (N_25163,N_24609,N_24937);
nor U25164 (N_25164,N_24881,N_24612);
or U25165 (N_25165,N_24956,N_24876);
xnor U25166 (N_25166,N_24635,N_24523);
nor U25167 (N_25167,N_24954,N_24806);
nand U25168 (N_25168,N_24578,N_24539);
nand U25169 (N_25169,N_24592,N_24586);
nor U25170 (N_25170,N_24967,N_24573);
xor U25171 (N_25171,N_24987,N_24951);
nor U25172 (N_25172,N_24559,N_24947);
xnor U25173 (N_25173,N_24727,N_24673);
or U25174 (N_25174,N_24814,N_24640);
or U25175 (N_25175,N_24807,N_24984);
xnor U25176 (N_25176,N_24893,N_24983);
and U25177 (N_25177,N_24552,N_24860);
nor U25178 (N_25178,N_24647,N_24530);
nand U25179 (N_25179,N_24657,N_24611);
nor U25180 (N_25180,N_24520,N_24944);
xor U25181 (N_25181,N_24902,N_24977);
nor U25182 (N_25182,N_24728,N_24875);
nor U25183 (N_25183,N_24787,N_24729);
and U25184 (N_25184,N_24873,N_24755);
and U25185 (N_25185,N_24563,N_24502);
or U25186 (N_25186,N_24538,N_24972);
or U25187 (N_25187,N_24770,N_24938);
and U25188 (N_25188,N_24643,N_24575);
nor U25189 (N_25189,N_24810,N_24761);
or U25190 (N_25190,N_24733,N_24857);
nor U25191 (N_25191,N_24978,N_24924);
nand U25192 (N_25192,N_24569,N_24842);
nand U25193 (N_25193,N_24702,N_24849);
or U25194 (N_25194,N_24832,N_24750);
or U25195 (N_25195,N_24623,N_24912);
and U25196 (N_25196,N_24510,N_24743);
nor U25197 (N_25197,N_24930,N_24866);
nand U25198 (N_25198,N_24679,N_24957);
or U25199 (N_25199,N_24649,N_24836);
nor U25200 (N_25200,N_24927,N_24800);
xnor U25201 (N_25201,N_24650,N_24536);
or U25202 (N_25202,N_24605,N_24851);
nor U25203 (N_25203,N_24888,N_24994);
and U25204 (N_25204,N_24949,N_24886);
nand U25205 (N_25205,N_24701,N_24777);
nand U25206 (N_25206,N_24932,N_24503);
and U25207 (N_25207,N_24786,N_24598);
xnor U25208 (N_25208,N_24864,N_24751);
nand U25209 (N_25209,N_24877,N_24996);
and U25210 (N_25210,N_24909,N_24628);
and U25211 (N_25211,N_24568,N_24900);
and U25212 (N_25212,N_24574,N_24589);
and U25213 (N_25213,N_24616,N_24935);
or U25214 (N_25214,N_24639,N_24904);
xnor U25215 (N_25215,N_24960,N_24638);
nor U25216 (N_25216,N_24993,N_24885);
xor U25217 (N_25217,N_24990,N_24684);
nor U25218 (N_25218,N_24726,N_24955);
nor U25219 (N_25219,N_24784,N_24916);
and U25220 (N_25220,N_24825,N_24659);
xnor U25221 (N_25221,N_24991,N_24545);
and U25222 (N_25222,N_24719,N_24627);
nor U25223 (N_25223,N_24899,N_24818);
nor U25224 (N_25224,N_24880,N_24798);
nor U25225 (N_25225,N_24982,N_24577);
and U25226 (N_25226,N_24758,N_24588);
or U25227 (N_25227,N_24797,N_24669);
xnor U25228 (N_25228,N_24801,N_24655);
or U25229 (N_25229,N_24709,N_24819);
nand U25230 (N_25230,N_24506,N_24997);
or U25231 (N_25231,N_24926,N_24541);
nor U25232 (N_25232,N_24835,N_24968);
or U25233 (N_25233,N_24907,N_24741);
or U25234 (N_25234,N_24862,N_24632);
xnor U25235 (N_25235,N_24898,N_24677);
nor U25236 (N_25236,N_24945,N_24809);
nor U25237 (N_25237,N_24980,N_24512);
nor U25238 (N_25238,N_24671,N_24799);
or U25239 (N_25239,N_24660,N_24622);
nor U25240 (N_25240,N_24550,N_24998);
and U25241 (N_25241,N_24513,N_24736);
and U25242 (N_25242,N_24644,N_24779);
xnor U25243 (N_25243,N_24556,N_24950);
xor U25244 (N_25244,N_24903,N_24790);
and U25245 (N_25245,N_24595,N_24802);
or U25246 (N_25246,N_24908,N_24691);
and U25247 (N_25247,N_24793,N_24883);
nor U25248 (N_25248,N_24645,N_24863);
nand U25249 (N_25249,N_24915,N_24572);
and U25250 (N_25250,N_24670,N_24565);
and U25251 (N_25251,N_24640,N_24743);
xor U25252 (N_25252,N_24611,N_24927);
xor U25253 (N_25253,N_24568,N_24764);
or U25254 (N_25254,N_24677,N_24878);
nor U25255 (N_25255,N_24504,N_24899);
xnor U25256 (N_25256,N_24980,N_24555);
or U25257 (N_25257,N_24506,N_24782);
nor U25258 (N_25258,N_24627,N_24820);
nand U25259 (N_25259,N_24605,N_24628);
and U25260 (N_25260,N_24844,N_24505);
and U25261 (N_25261,N_24889,N_24972);
nand U25262 (N_25262,N_24538,N_24504);
nand U25263 (N_25263,N_24530,N_24903);
or U25264 (N_25264,N_24528,N_24571);
xor U25265 (N_25265,N_24907,N_24891);
nand U25266 (N_25266,N_24589,N_24873);
and U25267 (N_25267,N_24952,N_24510);
nor U25268 (N_25268,N_24877,N_24523);
nand U25269 (N_25269,N_24868,N_24512);
and U25270 (N_25270,N_24664,N_24778);
and U25271 (N_25271,N_24785,N_24794);
or U25272 (N_25272,N_24715,N_24569);
nor U25273 (N_25273,N_24815,N_24863);
and U25274 (N_25274,N_24889,N_24988);
nor U25275 (N_25275,N_24949,N_24824);
and U25276 (N_25276,N_24949,N_24620);
or U25277 (N_25277,N_24532,N_24970);
nor U25278 (N_25278,N_24777,N_24659);
nor U25279 (N_25279,N_24711,N_24641);
nor U25280 (N_25280,N_24916,N_24849);
and U25281 (N_25281,N_24988,N_24709);
xnor U25282 (N_25282,N_24603,N_24945);
nor U25283 (N_25283,N_24612,N_24624);
nand U25284 (N_25284,N_24867,N_24807);
xnor U25285 (N_25285,N_24671,N_24526);
xnor U25286 (N_25286,N_24775,N_24674);
xnor U25287 (N_25287,N_24936,N_24979);
xor U25288 (N_25288,N_24823,N_24881);
or U25289 (N_25289,N_24748,N_24846);
and U25290 (N_25290,N_24660,N_24531);
and U25291 (N_25291,N_24593,N_24814);
nor U25292 (N_25292,N_24543,N_24999);
xor U25293 (N_25293,N_24622,N_24772);
nor U25294 (N_25294,N_24934,N_24631);
or U25295 (N_25295,N_24822,N_24709);
nor U25296 (N_25296,N_24757,N_24725);
nand U25297 (N_25297,N_24556,N_24645);
nor U25298 (N_25298,N_24573,N_24669);
and U25299 (N_25299,N_24887,N_24967);
xor U25300 (N_25300,N_24604,N_24830);
nor U25301 (N_25301,N_24965,N_24682);
nor U25302 (N_25302,N_24882,N_24582);
nor U25303 (N_25303,N_24988,N_24511);
nand U25304 (N_25304,N_24599,N_24965);
xor U25305 (N_25305,N_24594,N_24648);
nand U25306 (N_25306,N_24983,N_24740);
and U25307 (N_25307,N_24668,N_24871);
and U25308 (N_25308,N_24619,N_24899);
xor U25309 (N_25309,N_24903,N_24743);
and U25310 (N_25310,N_24537,N_24897);
nor U25311 (N_25311,N_24641,N_24988);
or U25312 (N_25312,N_24713,N_24719);
and U25313 (N_25313,N_24607,N_24750);
nor U25314 (N_25314,N_24830,N_24574);
or U25315 (N_25315,N_24672,N_24961);
and U25316 (N_25316,N_24640,N_24724);
nor U25317 (N_25317,N_24929,N_24535);
xnor U25318 (N_25318,N_24638,N_24721);
or U25319 (N_25319,N_24735,N_24695);
and U25320 (N_25320,N_24906,N_24803);
nand U25321 (N_25321,N_24857,N_24784);
or U25322 (N_25322,N_24891,N_24825);
nor U25323 (N_25323,N_24587,N_24930);
nor U25324 (N_25324,N_24977,N_24779);
xnor U25325 (N_25325,N_24737,N_24807);
nor U25326 (N_25326,N_24654,N_24546);
nor U25327 (N_25327,N_24837,N_24550);
nor U25328 (N_25328,N_24529,N_24756);
nand U25329 (N_25329,N_24950,N_24904);
xor U25330 (N_25330,N_24797,N_24739);
and U25331 (N_25331,N_24964,N_24961);
nor U25332 (N_25332,N_24723,N_24717);
nor U25333 (N_25333,N_24976,N_24920);
nor U25334 (N_25334,N_24670,N_24953);
and U25335 (N_25335,N_24881,N_24538);
nor U25336 (N_25336,N_24675,N_24681);
xor U25337 (N_25337,N_24926,N_24889);
xnor U25338 (N_25338,N_24828,N_24868);
or U25339 (N_25339,N_24970,N_24997);
xnor U25340 (N_25340,N_24501,N_24940);
or U25341 (N_25341,N_24829,N_24550);
or U25342 (N_25342,N_24522,N_24917);
nor U25343 (N_25343,N_24829,N_24761);
or U25344 (N_25344,N_24611,N_24676);
and U25345 (N_25345,N_24969,N_24957);
nand U25346 (N_25346,N_24944,N_24797);
nand U25347 (N_25347,N_24514,N_24516);
xnor U25348 (N_25348,N_24629,N_24921);
and U25349 (N_25349,N_24819,N_24714);
and U25350 (N_25350,N_24632,N_24665);
xor U25351 (N_25351,N_24982,N_24876);
nand U25352 (N_25352,N_24635,N_24605);
nor U25353 (N_25353,N_24753,N_24741);
nor U25354 (N_25354,N_24589,N_24923);
and U25355 (N_25355,N_24785,N_24562);
xor U25356 (N_25356,N_24750,N_24735);
xor U25357 (N_25357,N_24761,N_24820);
nor U25358 (N_25358,N_24586,N_24617);
xnor U25359 (N_25359,N_24730,N_24523);
nand U25360 (N_25360,N_24690,N_24899);
and U25361 (N_25361,N_24693,N_24977);
nor U25362 (N_25362,N_24777,N_24844);
nor U25363 (N_25363,N_24572,N_24570);
nand U25364 (N_25364,N_24683,N_24878);
and U25365 (N_25365,N_24736,N_24680);
nand U25366 (N_25366,N_24625,N_24526);
nand U25367 (N_25367,N_24888,N_24839);
nor U25368 (N_25368,N_24607,N_24771);
xnor U25369 (N_25369,N_24595,N_24589);
nor U25370 (N_25370,N_24603,N_24957);
nor U25371 (N_25371,N_24528,N_24702);
or U25372 (N_25372,N_24933,N_24871);
and U25373 (N_25373,N_24649,N_24638);
nand U25374 (N_25374,N_24775,N_24507);
and U25375 (N_25375,N_24661,N_24936);
nand U25376 (N_25376,N_24705,N_24793);
xor U25377 (N_25377,N_24789,N_24767);
nand U25378 (N_25378,N_24766,N_24759);
or U25379 (N_25379,N_24669,N_24636);
and U25380 (N_25380,N_24744,N_24829);
nor U25381 (N_25381,N_24744,N_24738);
xor U25382 (N_25382,N_24826,N_24585);
or U25383 (N_25383,N_24899,N_24987);
and U25384 (N_25384,N_24680,N_24923);
nor U25385 (N_25385,N_24803,N_24684);
or U25386 (N_25386,N_24833,N_24738);
xor U25387 (N_25387,N_24911,N_24672);
and U25388 (N_25388,N_24588,N_24755);
nand U25389 (N_25389,N_24577,N_24639);
or U25390 (N_25390,N_24874,N_24569);
nor U25391 (N_25391,N_24819,N_24912);
xnor U25392 (N_25392,N_24822,N_24946);
and U25393 (N_25393,N_24876,N_24780);
nor U25394 (N_25394,N_24664,N_24925);
nor U25395 (N_25395,N_24712,N_24615);
or U25396 (N_25396,N_24618,N_24609);
or U25397 (N_25397,N_24921,N_24917);
nor U25398 (N_25398,N_24742,N_24610);
or U25399 (N_25399,N_24565,N_24692);
or U25400 (N_25400,N_24948,N_24615);
nor U25401 (N_25401,N_24569,N_24516);
nor U25402 (N_25402,N_24955,N_24528);
xnor U25403 (N_25403,N_24787,N_24519);
xnor U25404 (N_25404,N_24728,N_24523);
nand U25405 (N_25405,N_24650,N_24833);
or U25406 (N_25406,N_24509,N_24731);
nor U25407 (N_25407,N_24715,N_24571);
nor U25408 (N_25408,N_24689,N_24910);
nand U25409 (N_25409,N_24714,N_24587);
or U25410 (N_25410,N_24688,N_24944);
nand U25411 (N_25411,N_24975,N_24952);
or U25412 (N_25412,N_24513,N_24619);
nand U25413 (N_25413,N_24674,N_24677);
nor U25414 (N_25414,N_24751,N_24789);
and U25415 (N_25415,N_24660,N_24596);
nand U25416 (N_25416,N_24976,N_24530);
xnor U25417 (N_25417,N_24556,N_24993);
xor U25418 (N_25418,N_24586,N_24637);
and U25419 (N_25419,N_24546,N_24742);
or U25420 (N_25420,N_24553,N_24592);
or U25421 (N_25421,N_24782,N_24785);
nor U25422 (N_25422,N_24969,N_24927);
and U25423 (N_25423,N_24998,N_24886);
nand U25424 (N_25424,N_24997,N_24942);
nor U25425 (N_25425,N_24975,N_24966);
nand U25426 (N_25426,N_24657,N_24873);
or U25427 (N_25427,N_24692,N_24523);
xor U25428 (N_25428,N_24583,N_24746);
or U25429 (N_25429,N_24519,N_24578);
or U25430 (N_25430,N_24757,N_24709);
and U25431 (N_25431,N_24662,N_24797);
xor U25432 (N_25432,N_24509,N_24589);
nand U25433 (N_25433,N_24950,N_24905);
nand U25434 (N_25434,N_24926,N_24733);
nand U25435 (N_25435,N_24617,N_24610);
and U25436 (N_25436,N_24684,N_24775);
and U25437 (N_25437,N_24524,N_24744);
nand U25438 (N_25438,N_24537,N_24654);
xnor U25439 (N_25439,N_24705,N_24590);
nand U25440 (N_25440,N_24857,N_24697);
and U25441 (N_25441,N_24534,N_24779);
nor U25442 (N_25442,N_24871,N_24818);
and U25443 (N_25443,N_24560,N_24690);
xor U25444 (N_25444,N_24592,N_24963);
xor U25445 (N_25445,N_24656,N_24770);
nand U25446 (N_25446,N_24698,N_24893);
xnor U25447 (N_25447,N_24982,N_24528);
xnor U25448 (N_25448,N_24708,N_24992);
and U25449 (N_25449,N_24961,N_24845);
nor U25450 (N_25450,N_24858,N_24997);
and U25451 (N_25451,N_24949,N_24903);
nor U25452 (N_25452,N_24950,N_24977);
and U25453 (N_25453,N_24610,N_24764);
and U25454 (N_25454,N_24883,N_24544);
xor U25455 (N_25455,N_24605,N_24792);
and U25456 (N_25456,N_24934,N_24791);
or U25457 (N_25457,N_24501,N_24925);
nand U25458 (N_25458,N_24939,N_24799);
nor U25459 (N_25459,N_24521,N_24686);
nand U25460 (N_25460,N_24626,N_24872);
and U25461 (N_25461,N_24588,N_24769);
and U25462 (N_25462,N_24602,N_24776);
nor U25463 (N_25463,N_24649,N_24554);
and U25464 (N_25464,N_24614,N_24951);
xor U25465 (N_25465,N_24967,N_24590);
nand U25466 (N_25466,N_24784,N_24786);
or U25467 (N_25467,N_24502,N_24524);
and U25468 (N_25468,N_24957,N_24972);
and U25469 (N_25469,N_24814,N_24584);
or U25470 (N_25470,N_24936,N_24734);
nand U25471 (N_25471,N_24895,N_24589);
nand U25472 (N_25472,N_24646,N_24689);
nor U25473 (N_25473,N_24505,N_24903);
and U25474 (N_25474,N_24729,N_24802);
xor U25475 (N_25475,N_24723,N_24885);
and U25476 (N_25476,N_24620,N_24935);
nor U25477 (N_25477,N_24788,N_24541);
nor U25478 (N_25478,N_24828,N_24725);
nor U25479 (N_25479,N_24931,N_24710);
and U25480 (N_25480,N_24582,N_24500);
xnor U25481 (N_25481,N_24819,N_24521);
nand U25482 (N_25482,N_24744,N_24818);
and U25483 (N_25483,N_24953,N_24758);
nand U25484 (N_25484,N_24718,N_24643);
nand U25485 (N_25485,N_24706,N_24803);
nor U25486 (N_25486,N_24963,N_24657);
and U25487 (N_25487,N_24921,N_24793);
nand U25488 (N_25488,N_24645,N_24615);
nand U25489 (N_25489,N_24813,N_24721);
or U25490 (N_25490,N_24863,N_24842);
or U25491 (N_25491,N_24940,N_24954);
and U25492 (N_25492,N_24921,N_24868);
and U25493 (N_25493,N_24549,N_24969);
and U25494 (N_25494,N_24796,N_24841);
nor U25495 (N_25495,N_24527,N_24526);
and U25496 (N_25496,N_24676,N_24629);
nand U25497 (N_25497,N_24947,N_24842);
or U25498 (N_25498,N_24758,N_24675);
nand U25499 (N_25499,N_24508,N_24717);
and U25500 (N_25500,N_25226,N_25068);
or U25501 (N_25501,N_25122,N_25279);
nand U25502 (N_25502,N_25019,N_25299);
nor U25503 (N_25503,N_25463,N_25184);
nor U25504 (N_25504,N_25262,N_25159);
nor U25505 (N_25505,N_25442,N_25333);
nor U25506 (N_25506,N_25417,N_25478);
nand U25507 (N_25507,N_25485,N_25462);
and U25508 (N_25508,N_25156,N_25473);
xor U25509 (N_25509,N_25228,N_25407);
nand U25510 (N_25510,N_25298,N_25222);
xor U25511 (N_25511,N_25310,N_25469);
nor U25512 (N_25512,N_25413,N_25346);
xnor U25513 (N_25513,N_25146,N_25321);
or U25514 (N_25514,N_25483,N_25154);
or U25515 (N_25515,N_25108,N_25367);
nor U25516 (N_25516,N_25339,N_25188);
or U25517 (N_25517,N_25396,N_25111);
or U25518 (N_25518,N_25097,N_25081);
nand U25519 (N_25519,N_25471,N_25240);
nor U25520 (N_25520,N_25120,N_25223);
nor U25521 (N_25521,N_25304,N_25128);
nand U25522 (N_25522,N_25351,N_25244);
or U25523 (N_25523,N_25118,N_25271);
or U25524 (N_25524,N_25455,N_25211);
xor U25525 (N_25525,N_25371,N_25054);
or U25526 (N_25526,N_25431,N_25168);
nand U25527 (N_25527,N_25105,N_25134);
or U25528 (N_25528,N_25464,N_25283);
xnor U25529 (N_25529,N_25006,N_25280);
xor U25530 (N_25530,N_25011,N_25058);
or U25531 (N_25531,N_25055,N_25443);
and U25532 (N_25532,N_25123,N_25063);
and U25533 (N_25533,N_25153,N_25099);
or U25534 (N_25534,N_25377,N_25352);
and U25535 (N_25535,N_25340,N_25379);
nor U25536 (N_25536,N_25247,N_25158);
and U25537 (N_25537,N_25130,N_25495);
nor U25538 (N_25538,N_25422,N_25219);
and U25539 (N_25539,N_25014,N_25287);
xor U25540 (N_25540,N_25381,N_25482);
xor U25541 (N_25541,N_25163,N_25364);
and U25542 (N_25542,N_25043,N_25409);
or U25543 (N_25543,N_25079,N_25213);
nand U25544 (N_25544,N_25344,N_25065);
nand U25545 (N_25545,N_25446,N_25424);
nor U25546 (N_25546,N_25400,N_25169);
and U25547 (N_25547,N_25303,N_25257);
or U25548 (N_25548,N_25430,N_25176);
nor U25549 (N_25549,N_25102,N_25467);
nor U25550 (N_25550,N_25235,N_25127);
or U25551 (N_25551,N_25326,N_25353);
and U25552 (N_25552,N_25124,N_25139);
nor U25553 (N_25553,N_25496,N_25293);
nor U25554 (N_25554,N_25217,N_25115);
and U25555 (N_25555,N_25104,N_25276);
and U25556 (N_25556,N_25452,N_25477);
nand U25557 (N_25557,N_25288,N_25461);
or U25558 (N_25558,N_25425,N_25343);
nor U25559 (N_25559,N_25423,N_25162);
xor U25560 (N_25560,N_25465,N_25447);
or U25561 (N_25561,N_25137,N_25218);
xor U25562 (N_25562,N_25200,N_25155);
nand U25563 (N_25563,N_25245,N_25246);
and U25564 (N_25564,N_25183,N_25077);
nand U25565 (N_25565,N_25107,N_25302);
nor U25566 (N_25566,N_25434,N_25345);
xor U25567 (N_25567,N_25480,N_25214);
nand U25568 (N_25568,N_25392,N_25318);
nor U25569 (N_25569,N_25185,N_25349);
and U25570 (N_25570,N_25490,N_25016);
or U25571 (N_25571,N_25397,N_25225);
xnor U25572 (N_25572,N_25263,N_25091);
and U25573 (N_25573,N_25267,N_25207);
and U25574 (N_25574,N_25157,N_25239);
or U25575 (N_25575,N_25451,N_25121);
nand U25576 (N_25576,N_25320,N_25142);
or U25577 (N_25577,N_25062,N_25338);
xnor U25578 (N_25578,N_25281,N_25388);
nor U25579 (N_25579,N_25266,N_25210);
xor U25580 (N_25580,N_25103,N_25275);
xor U25581 (N_25581,N_25323,N_25265);
nor U25582 (N_25582,N_25284,N_25282);
nor U25583 (N_25583,N_25050,N_25256);
and U25584 (N_25584,N_25291,N_25454);
xnor U25585 (N_25585,N_25313,N_25076);
nand U25586 (N_25586,N_25090,N_25309);
or U25587 (N_25587,N_25390,N_25202);
nor U25588 (N_25588,N_25285,N_25190);
and U25589 (N_25589,N_25269,N_25389);
nand U25590 (N_25590,N_25297,N_25393);
nor U25591 (N_25591,N_25368,N_25420);
and U25592 (N_25592,N_25445,N_25365);
nor U25593 (N_25593,N_25316,N_25221);
xnor U25594 (N_25594,N_25067,N_25059);
or U25595 (N_25595,N_25372,N_25060);
xnor U25596 (N_25596,N_25151,N_25023);
nand U25597 (N_25597,N_25362,N_25479);
nor U25598 (N_25598,N_25132,N_25039);
nor U25599 (N_25599,N_25013,N_25319);
or U25600 (N_25600,N_25497,N_25342);
xnor U25601 (N_25601,N_25402,N_25406);
nor U25602 (N_25602,N_25051,N_25233);
nor U25603 (N_25603,N_25251,N_25106);
nand U25604 (N_25604,N_25486,N_25456);
and U25605 (N_25605,N_25459,N_25186);
xnor U25606 (N_25606,N_25037,N_25268);
nand U25607 (N_25607,N_25112,N_25436);
nor U25608 (N_25608,N_25475,N_25029);
nor U25609 (N_25609,N_25189,N_25135);
xnor U25610 (N_25610,N_25136,N_25373);
nand U25611 (N_25611,N_25408,N_25432);
nand U25612 (N_25612,N_25180,N_25195);
and U25613 (N_25613,N_25002,N_25089);
nand U25614 (N_25614,N_25070,N_25057);
or U25615 (N_25615,N_25053,N_25071);
nor U25616 (N_25616,N_25172,N_25378);
nand U25617 (N_25617,N_25131,N_25441);
xnor U25618 (N_25618,N_25008,N_25166);
nor U25619 (N_25619,N_25005,N_25427);
xor U25620 (N_25620,N_25095,N_25332);
nor U25621 (N_25621,N_25040,N_25044);
nand U25622 (N_25622,N_25336,N_25241);
nand U25623 (N_25623,N_25093,N_25492);
and U25624 (N_25624,N_25327,N_25259);
xnor U25625 (N_25625,N_25238,N_25292);
nor U25626 (N_25626,N_25370,N_25468);
xor U25627 (N_25627,N_25253,N_25286);
and U25628 (N_25628,N_25125,N_25003);
nor U25629 (N_25629,N_25160,N_25147);
nand U25630 (N_25630,N_25335,N_25295);
nand U25631 (N_25631,N_25322,N_25341);
xnor U25632 (N_25632,N_25174,N_25260);
or U25633 (N_25633,N_25152,N_25363);
xnor U25634 (N_25634,N_25498,N_25119);
nand U25635 (N_25635,N_25382,N_25435);
nor U25636 (N_25636,N_25359,N_25398);
nor U25637 (N_25637,N_25206,N_25182);
and U25638 (N_25638,N_25272,N_25045);
nor U25639 (N_25639,N_25474,N_25086);
nor U25640 (N_25640,N_25187,N_25437);
xnor U25641 (N_25641,N_25440,N_25024);
nand U25642 (N_25642,N_25041,N_25412);
nor U25643 (N_25643,N_25419,N_25021);
nor U25644 (N_25644,N_25078,N_25109);
nor U25645 (N_25645,N_25209,N_25315);
nand U25646 (N_25646,N_25360,N_25375);
nand U25647 (N_25647,N_25178,N_25227);
nand U25648 (N_25648,N_25012,N_25036);
nand U25649 (N_25649,N_25004,N_25141);
nor U25650 (N_25650,N_25410,N_25411);
and U25651 (N_25651,N_25258,N_25052);
nor U25652 (N_25652,N_25294,N_25224);
nor U25653 (N_25653,N_25374,N_25290);
or U25654 (N_25654,N_25305,N_25049);
xor U25655 (N_25655,N_25032,N_25337);
or U25656 (N_25656,N_25385,N_25025);
xnor U25657 (N_25657,N_25248,N_25350);
nand U25658 (N_25658,N_25354,N_25215);
or U25659 (N_25659,N_25177,N_25080);
nand U25660 (N_25660,N_25236,N_25194);
xnor U25661 (N_25661,N_25018,N_25252);
or U25662 (N_25662,N_25493,N_25391);
or U25663 (N_25663,N_25403,N_25110);
nor U25664 (N_25664,N_25031,N_25317);
xnor U25665 (N_25665,N_25376,N_25231);
nor U25666 (N_25666,N_25444,N_25201);
or U25667 (N_25667,N_25254,N_25237);
xor U25668 (N_25668,N_25173,N_25167);
nor U25669 (N_25669,N_25387,N_25192);
and U25670 (N_25670,N_25384,N_25175);
or U25671 (N_25671,N_25330,N_25191);
or U25672 (N_25672,N_25439,N_25000);
and U25673 (N_25673,N_25449,N_25361);
xor U25674 (N_25674,N_25145,N_25347);
nand U25675 (N_25675,N_25073,N_25116);
or U25676 (N_25676,N_25453,N_25230);
xor U25677 (N_25677,N_25488,N_25399);
nor U25678 (N_25678,N_25092,N_25204);
and U25679 (N_25679,N_25010,N_25181);
nand U25680 (N_25680,N_25289,N_25205);
nor U25681 (N_25681,N_25489,N_25220);
and U25682 (N_25682,N_25007,N_25329);
and U25683 (N_25683,N_25035,N_25415);
nand U25684 (N_25684,N_25296,N_25494);
and U25685 (N_25685,N_25328,N_25426);
and U25686 (N_25686,N_25458,N_25311);
xor U25687 (N_25687,N_25179,N_25331);
nor U25688 (N_25688,N_25307,N_25216);
nand U25689 (N_25689,N_25082,N_25476);
or U25690 (N_25690,N_25033,N_25075);
xor U25691 (N_25691,N_25457,N_25369);
or U25692 (N_25692,N_25056,N_25171);
or U25693 (N_25693,N_25113,N_25199);
or U25694 (N_25694,N_25069,N_25300);
nor U25695 (N_25695,N_25386,N_25366);
or U25696 (N_25696,N_25149,N_25015);
xor U25697 (N_25697,N_25261,N_25416);
nand U25698 (N_25698,N_25487,N_25243);
nand U25699 (N_25699,N_25027,N_25450);
and U25700 (N_25700,N_25394,N_25061);
or U25701 (N_25701,N_25277,N_25026);
nor U25702 (N_25702,N_25255,N_25229);
nor U25703 (N_25703,N_25034,N_25203);
nor U25704 (N_25704,N_25165,N_25356);
nor U25705 (N_25705,N_25481,N_25405);
or U25706 (N_25706,N_25306,N_25499);
nand U25707 (N_25707,N_25438,N_25020);
nand U25708 (N_25708,N_25022,N_25314);
xnor U25709 (N_25709,N_25126,N_25138);
or U25710 (N_25710,N_25148,N_25140);
nor U25711 (N_25711,N_25301,N_25250);
nand U25712 (N_25712,N_25270,N_25421);
xnor U25713 (N_25713,N_25358,N_25466);
xor U25714 (N_25714,N_25150,N_25074);
and U25715 (N_25715,N_25278,N_25087);
or U25716 (N_25716,N_25197,N_25355);
and U25717 (N_25717,N_25009,N_25429);
nor U25718 (N_25718,N_25088,N_25030);
nand U25719 (N_25719,N_25274,N_25418);
or U25720 (N_25720,N_25017,N_25098);
nand U25721 (N_25721,N_25084,N_25083);
nand U25722 (N_25722,N_25273,N_25460);
and U25723 (N_25723,N_25161,N_25348);
nor U25724 (N_25724,N_25001,N_25117);
xor U25725 (N_25725,N_25380,N_25085);
or U25726 (N_25726,N_25170,N_25383);
nand U25727 (N_25727,N_25234,N_25414);
xor U25728 (N_25728,N_25308,N_25094);
and U25729 (N_25729,N_25249,N_25470);
nand U25730 (N_25730,N_25193,N_25028);
nor U25731 (N_25731,N_25048,N_25208);
and U25732 (N_25732,N_25484,N_25472);
xnor U25733 (N_25733,N_25325,N_25491);
and U25734 (N_25734,N_25242,N_25196);
or U25735 (N_25735,N_25143,N_25448);
xor U25736 (N_25736,N_25072,N_25042);
xnor U25737 (N_25737,N_25114,N_25066);
xor U25738 (N_25738,N_25428,N_25395);
nor U25739 (N_25739,N_25198,N_25129);
nand U25740 (N_25740,N_25064,N_25334);
and U25741 (N_25741,N_25404,N_25264);
or U25742 (N_25742,N_25101,N_25357);
xnor U25743 (N_25743,N_25164,N_25232);
nand U25744 (N_25744,N_25212,N_25046);
nor U25745 (N_25745,N_25401,N_25312);
xor U25746 (N_25746,N_25324,N_25144);
nand U25747 (N_25747,N_25433,N_25100);
and U25748 (N_25748,N_25096,N_25133);
nor U25749 (N_25749,N_25038,N_25047);
xor U25750 (N_25750,N_25306,N_25247);
nor U25751 (N_25751,N_25304,N_25161);
or U25752 (N_25752,N_25457,N_25102);
nand U25753 (N_25753,N_25028,N_25017);
nor U25754 (N_25754,N_25110,N_25268);
or U25755 (N_25755,N_25453,N_25391);
and U25756 (N_25756,N_25153,N_25058);
and U25757 (N_25757,N_25279,N_25234);
and U25758 (N_25758,N_25127,N_25460);
or U25759 (N_25759,N_25201,N_25194);
nand U25760 (N_25760,N_25099,N_25363);
xor U25761 (N_25761,N_25433,N_25470);
and U25762 (N_25762,N_25474,N_25159);
and U25763 (N_25763,N_25172,N_25201);
xor U25764 (N_25764,N_25011,N_25068);
or U25765 (N_25765,N_25236,N_25474);
and U25766 (N_25766,N_25187,N_25146);
and U25767 (N_25767,N_25269,N_25159);
nor U25768 (N_25768,N_25067,N_25415);
nor U25769 (N_25769,N_25088,N_25076);
and U25770 (N_25770,N_25450,N_25104);
or U25771 (N_25771,N_25083,N_25109);
or U25772 (N_25772,N_25119,N_25453);
xnor U25773 (N_25773,N_25020,N_25030);
or U25774 (N_25774,N_25267,N_25404);
or U25775 (N_25775,N_25429,N_25337);
and U25776 (N_25776,N_25036,N_25341);
or U25777 (N_25777,N_25048,N_25032);
nand U25778 (N_25778,N_25210,N_25013);
xor U25779 (N_25779,N_25495,N_25246);
and U25780 (N_25780,N_25202,N_25376);
and U25781 (N_25781,N_25436,N_25285);
xor U25782 (N_25782,N_25421,N_25149);
and U25783 (N_25783,N_25148,N_25149);
nor U25784 (N_25784,N_25459,N_25263);
nor U25785 (N_25785,N_25439,N_25104);
nand U25786 (N_25786,N_25479,N_25067);
xor U25787 (N_25787,N_25365,N_25458);
or U25788 (N_25788,N_25266,N_25478);
nand U25789 (N_25789,N_25315,N_25057);
nand U25790 (N_25790,N_25203,N_25207);
xor U25791 (N_25791,N_25361,N_25039);
nand U25792 (N_25792,N_25113,N_25004);
or U25793 (N_25793,N_25161,N_25229);
nand U25794 (N_25794,N_25030,N_25304);
nor U25795 (N_25795,N_25393,N_25110);
xor U25796 (N_25796,N_25178,N_25279);
nor U25797 (N_25797,N_25473,N_25480);
nand U25798 (N_25798,N_25001,N_25436);
and U25799 (N_25799,N_25475,N_25460);
and U25800 (N_25800,N_25268,N_25197);
or U25801 (N_25801,N_25007,N_25463);
and U25802 (N_25802,N_25027,N_25342);
and U25803 (N_25803,N_25363,N_25309);
nor U25804 (N_25804,N_25482,N_25046);
xor U25805 (N_25805,N_25499,N_25490);
and U25806 (N_25806,N_25282,N_25482);
and U25807 (N_25807,N_25016,N_25291);
and U25808 (N_25808,N_25120,N_25421);
xnor U25809 (N_25809,N_25357,N_25041);
nor U25810 (N_25810,N_25374,N_25111);
or U25811 (N_25811,N_25114,N_25102);
and U25812 (N_25812,N_25181,N_25166);
nor U25813 (N_25813,N_25398,N_25246);
nand U25814 (N_25814,N_25027,N_25269);
xnor U25815 (N_25815,N_25270,N_25257);
nor U25816 (N_25816,N_25296,N_25308);
xnor U25817 (N_25817,N_25096,N_25077);
xnor U25818 (N_25818,N_25009,N_25230);
or U25819 (N_25819,N_25089,N_25161);
and U25820 (N_25820,N_25001,N_25014);
nor U25821 (N_25821,N_25239,N_25273);
and U25822 (N_25822,N_25424,N_25452);
xnor U25823 (N_25823,N_25240,N_25224);
or U25824 (N_25824,N_25114,N_25325);
and U25825 (N_25825,N_25087,N_25220);
and U25826 (N_25826,N_25274,N_25293);
xnor U25827 (N_25827,N_25488,N_25087);
and U25828 (N_25828,N_25247,N_25002);
and U25829 (N_25829,N_25219,N_25400);
or U25830 (N_25830,N_25353,N_25380);
nor U25831 (N_25831,N_25357,N_25029);
or U25832 (N_25832,N_25318,N_25045);
or U25833 (N_25833,N_25385,N_25266);
or U25834 (N_25834,N_25471,N_25018);
nand U25835 (N_25835,N_25188,N_25495);
xnor U25836 (N_25836,N_25304,N_25455);
and U25837 (N_25837,N_25088,N_25204);
and U25838 (N_25838,N_25039,N_25417);
nand U25839 (N_25839,N_25145,N_25248);
and U25840 (N_25840,N_25281,N_25049);
nor U25841 (N_25841,N_25017,N_25404);
xnor U25842 (N_25842,N_25320,N_25166);
nand U25843 (N_25843,N_25365,N_25300);
and U25844 (N_25844,N_25097,N_25336);
nor U25845 (N_25845,N_25186,N_25320);
and U25846 (N_25846,N_25325,N_25093);
xor U25847 (N_25847,N_25469,N_25461);
and U25848 (N_25848,N_25384,N_25342);
and U25849 (N_25849,N_25255,N_25321);
nor U25850 (N_25850,N_25026,N_25002);
xnor U25851 (N_25851,N_25387,N_25182);
nand U25852 (N_25852,N_25013,N_25121);
xnor U25853 (N_25853,N_25164,N_25482);
and U25854 (N_25854,N_25410,N_25055);
xnor U25855 (N_25855,N_25427,N_25065);
nand U25856 (N_25856,N_25355,N_25234);
nor U25857 (N_25857,N_25051,N_25439);
and U25858 (N_25858,N_25338,N_25286);
xnor U25859 (N_25859,N_25389,N_25417);
or U25860 (N_25860,N_25250,N_25387);
xor U25861 (N_25861,N_25198,N_25477);
and U25862 (N_25862,N_25208,N_25097);
xor U25863 (N_25863,N_25172,N_25470);
xor U25864 (N_25864,N_25064,N_25411);
nand U25865 (N_25865,N_25272,N_25435);
and U25866 (N_25866,N_25091,N_25195);
or U25867 (N_25867,N_25143,N_25332);
xnor U25868 (N_25868,N_25434,N_25060);
nor U25869 (N_25869,N_25043,N_25304);
xor U25870 (N_25870,N_25031,N_25174);
xnor U25871 (N_25871,N_25089,N_25249);
or U25872 (N_25872,N_25163,N_25387);
or U25873 (N_25873,N_25051,N_25336);
or U25874 (N_25874,N_25288,N_25007);
or U25875 (N_25875,N_25246,N_25364);
or U25876 (N_25876,N_25244,N_25297);
nor U25877 (N_25877,N_25151,N_25170);
or U25878 (N_25878,N_25083,N_25027);
or U25879 (N_25879,N_25188,N_25113);
and U25880 (N_25880,N_25341,N_25167);
or U25881 (N_25881,N_25464,N_25300);
xnor U25882 (N_25882,N_25171,N_25491);
xor U25883 (N_25883,N_25251,N_25389);
and U25884 (N_25884,N_25186,N_25474);
xnor U25885 (N_25885,N_25498,N_25414);
nor U25886 (N_25886,N_25245,N_25052);
or U25887 (N_25887,N_25333,N_25074);
xor U25888 (N_25888,N_25288,N_25313);
nand U25889 (N_25889,N_25463,N_25312);
or U25890 (N_25890,N_25427,N_25306);
xor U25891 (N_25891,N_25465,N_25067);
and U25892 (N_25892,N_25322,N_25118);
xnor U25893 (N_25893,N_25169,N_25239);
xor U25894 (N_25894,N_25162,N_25183);
xor U25895 (N_25895,N_25045,N_25173);
nand U25896 (N_25896,N_25053,N_25185);
nor U25897 (N_25897,N_25268,N_25449);
nor U25898 (N_25898,N_25209,N_25317);
and U25899 (N_25899,N_25167,N_25330);
nor U25900 (N_25900,N_25385,N_25088);
nand U25901 (N_25901,N_25319,N_25378);
nand U25902 (N_25902,N_25264,N_25061);
xnor U25903 (N_25903,N_25019,N_25305);
or U25904 (N_25904,N_25345,N_25291);
or U25905 (N_25905,N_25242,N_25349);
or U25906 (N_25906,N_25442,N_25115);
xnor U25907 (N_25907,N_25198,N_25380);
nand U25908 (N_25908,N_25293,N_25294);
nor U25909 (N_25909,N_25245,N_25042);
nand U25910 (N_25910,N_25284,N_25403);
or U25911 (N_25911,N_25313,N_25391);
or U25912 (N_25912,N_25287,N_25359);
nor U25913 (N_25913,N_25083,N_25368);
or U25914 (N_25914,N_25414,N_25400);
and U25915 (N_25915,N_25245,N_25021);
nand U25916 (N_25916,N_25275,N_25398);
nor U25917 (N_25917,N_25324,N_25290);
and U25918 (N_25918,N_25169,N_25167);
and U25919 (N_25919,N_25374,N_25257);
nand U25920 (N_25920,N_25041,N_25109);
nor U25921 (N_25921,N_25230,N_25329);
nand U25922 (N_25922,N_25346,N_25246);
or U25923 (N_25923,N_25349,N_25271);
and U25924 (N_25924,N_25190,N_25096);
nor U25925 (N_25925,N_25186,N_25342);
and U25926 (N_25926,N_25247,N_25290);
nand U25927 (N_25927,N_25265,N_25162);
nand U25928 (N_25928,N_25090,N_25011);
xor U25929 (N_25929,N_25146,N_25341);
nor U25930 (N_25930,N_25416,N_25104);
and U25931 (N_25931,N_25110,N_25187);
xnor U25932 (N_25932,N_25158,N_25402);
nor U25933 (N_25933,N_25049,N_25343);
or U25934 (N_25934,N_25018,N_25040);
or U25935 (N_25935,N_25116,N_25119);
and U25936 (N_25936,N_25230,N_25043);
or U25937 (N_25937,N_25195,N_25317);
xor U25938 (N_25938,N_25233,N_25199);
nand U25939 (N_25939,N_25363,N_25499);
nand U25940 (N_25940,N_25470,N_25409);
nor U25941 (N_25941,N_25183,N_25407);
nand U25942 (N_25942,N_25276,N_25049);
and U25943 (N_25943,N_25017,N_25198);
nor U25944 (N_25944,N_25014,N_25050);
or U25945 (N_25945,N_25173,N_25197);
and U25946 (N_25946,N_25153,N_25329);
nand U25947 (N_25947,N_25487,N_25421);
nand U25948 (N_25948,N_25181,N_25354);
xor U25949 (N_25949,N_25429,N_25466);
nor U25950 (N_25950,N_25306,N_25180);
xnor U25951 (N_25951,N_25085,N_25192);
nand U25952 (N_25952,N_25057,N_25105);
xnor U25953 (N_25953,N_25219,N_25163);
nand U25954 (N_25954,N_25302,N_25275);
or U25955 (N_25955,N_25346,N_25137);
or U25956 (N_25956,N_25380,N_25028);
nor U25957 (N_25957,N_25241,N_25110);
nor U25958 (N_25958,N_25151,N_25256);
nor U25959 (N_25959,N_25261,N_25002);
or U25960 (N_25960,N_25465,N_25148);
and U25961 (N_25961,N_25355,N_25137);
nand U25962 (N_25962,N_25375,N_25045);
and U25963 (N_25963,N_25295,N_25380);
or U25964 (N_25964,N_25149,N_25243);
or U25965 (N_25965,N_25373,N_25222);
nand U25966 (N_25966,N_25225,N_25443);
or U25967 (N_25967,N_25404,N_25332);
nand U25968 (N_25968,N_25465,N_25419);
nand U25969 (N_25969,N_25052,N_25417);
and U25970 (N_25970,N_25260,N_25247);
and U25971 (N_25971,N_25145,N_25421);
nand U25972 (N_25972,N_25061,N_25474);
or U25973 (N_25973,N_25062,N_25150);
xor U25974 (N_25974,N_25359,N_25014);
and U25975 (N_25975,N_25199,N_25355);
nand U25976 (N_25976,N_25051,N_25407);
nor U25977 (N_25977,N_25164,N_25162);
or U25978 (N_25978,N_25402,N_25177);
nand U25979 (N_25979,N_25274,N_25011);
xor U25980 (N_25980,N_25243,N_25140);
nand U25981 (N_25981,N_25277,N_25096);
xnor U25982 (N_25982,N_25203,N_25083);
or U25983 (N_25983,N_25390,N_25496);
and U25984 (N_25984,N_25407,N_25170);
nand U25985 (N_25985,N_25282,N_25256);
nand U25986 (N_25986,N_25115,N_25334);
and U25987 (N_25987,N_25087,N_25301);
and U25988 (N_25988,N_25414,N_25121);
nand U25989 (N_25989,N_25482,N_25040);
xor U25990 (N_25990,N_25490,N_25157);
and U25991 (N_25991,N_25072,N_25233);
and U25992 (N_25992,N_25373,N_25268);
xor U25993 (N_25993,N_25168,N_25198);
nor U25994 (N_25994,N_25491,N_25162);
nand U25995 (N_25995,N_25349,N_25304);
and U25996 (N_25996,N_25329,N_25060);
nor U25997 (N_25997,N_25065,N_25323);
or U25998 (N_25998,N_25182,N_25032);
xnor U25999 (N_25999,N_25356,N_25270);
and U26000 (N_26000,N_25679,N_25947);
nor U26001 (N_26001,N_25723,N_25642);
xor U26002 (N_26002,N_25885,N_25744);
nand U26003 (N_26003,N_25886,N_25656);
or U26004 (N_26004,N_25576,N_25717);
nand U26005 (N_26005,N_25607,N_25930);
and U26006 (N_26006,N_25553,N_25754);
or U26007 (N_26007,N_25574,N_25884);
xnor U26008 (N_26008,N_25802,N_25568);
xnor U26009 (N_26009,N_25775,N_25640);
nor U26010 (N_26010,N_25601,N_25895);
xnor U26011 (N_26011,N_25936,N_25849);
nor U26012 (N_26012,N_25697,N_25523);
xor U26013 (N_26013,N_25690,N_25643);
xor U26014 (N_26014,N_25801,N_25958);
and U26015 (N_26015,N_25985,N_25605);
and U26016 (N_26016,N_25810,N_25909);
xor U26017 (N_26017,N_25875,N_25862);
or U26018 (N_26018,N_25852,N_25592);
xnor U26019 (N_26019,N_25745,N_25767);
or U26020 (N_26020,N_25560,N_25544);
and U26021 (N_26021,N_25701,N_25575);
xor U26022 (N_26022,N_25880,N_25755);
xnor U26023 (N_26023,N_25883,N_25835);
or U26024 (N_26024,N_25976,N_25861);
nor U26025 (N_26025,N_25736,N_25820);
xnor U26026 (N_26026,N_25946,N_25704);
xor U26027 (N_26027,N_25806,N_25500);
or U26028 (N_26028,N_25757,N_25915);
and U26029 (N_26029,N_25538,N_25663);
or U26030 (N_26030,N_25903,N_25974);
or U26031 (N_26031,N_25808,N_25518);
or U26032 (N_26032,N_25552,N_25831);
or U26033 (N_26033,N_25631,N_25617);
and U26034 (N_26034,N_25562,N_25763);
or U26035 (N_26035,N_25972,N_25781);
and U26036 (N_26036,N_25752,N_25514);
nor U26037 (N_26037,N_25561,N_25776);
nand U26038 (N_26038,N_25864,N_25993);
nand U26039 (N_26039,N_25811,N_25922);
nand U26040 (N_26040,N_25829,N_25839);
xor U26041 (N_26041,N_25652,N_25600);
xor U26042 (N_26042,N_25629,N_25730);
and U26043 (N_26043,N_25804,N_25856);
nand U26044 (N_26044,N_25739,N_25741);
nand U26045 (N_26045,N_25878,N_25869);
and U26046 (N_26046,N_25892,N_25623);
or U26047 (N_26047,N_25522,N_25657);
xor U26048 (N_26048,N_25774,N_25813);
nand U26049 (N_26049,N_25935,N_25511);
nand U26050 (N_26050,N_25727,N_25753);
and U26051 (N_26051,N_25902,N_25718);
or U26052 (N_26052,N_25798,N_25932);
xnor U26053 (N_26053,N_25826,N_25731);
nand U26054 (N_26054,N_25998,N_25703);
and U26055 (N_26055,N_25661,N_25858);
nor U26056 (N_26056,N_25585,N_25799);
and U26057 (N_26057,N_25983,N_25728);
nand U26058 (N_26058,N_25686,N_25664);
nand U26059 (N_26059,N_25773,N_25673);
or U26060 (N_26060,N_25848,N_25805);
and U26061 (N_26061,N_25843,N_25684);
xnor U26062 (N_26062,N_25578,N_25994);
xnor U26063 (N_26063,N_25724,N_25867);
and U26064 (N_26064,N_25768,N_25596);
nand U26065 (N_26065,N_25943,N_25865);
and U26066 (N_26066,N_25857,N_25588);
xor U26067 (N_26067,N_25853,N_25954);
or U26068 (N_26068,N_25982,N_25921);
or U26069 (N_26069,N_25609,N_25780);
or U26070 (N_26070,N_25507,N_25792);
or U26071 (N_26071,N_25997,N_25719);
nand U26072 (N_26072,N_25635,N_25988);
xor U26073 (N_26073,N_25937,N_25658);
xnor U26074 (N_26074,N_25938,N_25554);
xnor U26075 (N_26075,N_25762,N_25659);
xnor U26076 (N_26076,N_25549,N_25868);
nand U26077 (N_26077,N_25587,N_25711);
nor U26078 (N_26078,N_25740,N_25981);
or U26079 (N_26079,N_25772,N_25706);
or U26080 (N_26080,N_25691,N_25709);
nor U26081 (N_26081,N_25577,N_25604);
and U26082 (N_26082,N_25877,N_25590);
nand U26083 (N_26083,N_25565,N_25699);
nand U26084 (N_26084,N_25818,N_25694);
nand U26085 (N_26085,N_25662,N_25509);
or U26086 (N_26086,N_25738,N_25505);
nand U26087 (N_26087,N_25645,N_25615);
and U26088 (N_26088,N_25644,N_25618);
nand U26089 (N_26089,N_25795,N_25622);
nor U26090 (N_26090,N_25546,N_25572);
and U26091 (N_26091,N_25542,N_25681);
xnor U26092 (N_26092,N_25692,N_25667);
xor U26093 (N_26093,N_25608,N_25793);
nand U26094 (N_26094,N_25899,N_25545);
nor U26095 (N_26095,N_25625,N_25917);
nor U26096 (N_26096,N_25566,N_25599);
and U26097 (N_26097,N_25961,N_25732);
xnor U26098 (N_26098,N_25636,N_25823);
xor U26099 (N_26099,N_25606,N_25957);
or U26100 (N_26100,N_25726,N_25879);
xor U26101 (N_26101,N_25713,N_25648);
nor U26102 (N_26102,N_25787,N_25620);
xnor U26103 (N_26103,N_25968,N_25907);
xor U26104 (N_26104,N_25627,N_25613);
and U26105 (N_26105,N_25677,N_25945);
or U26106 (N_26106,N_25626,N_25586);
nor U26107 (N_26107,N_25710,N_25890);
xnor U26108 (N_26108,N_25898,N_25595);
and U26109 (N_26109,N_25926,N_25756);
and U26110 (N_26110,N_25942,N_25859);
nand U26111 (N_26111,N_25678,N_25977);
nor U26112 (N_26112,N_25580,N_25516);
xnor U26113 (N_26113,N_25797,N_25962);
nor U26114 (N_26114,N_25950,N_25929);
nand U26115 (N_26115,N_25573,N_25771);
nand U26116 (N_26116,N_25670,N_25651);
nand U26117 (N_26117,N_25896,N_25931);
and U26118 (N_26118,N_25948,N_25784);
nand U26119 (N_26119,N_25758,N_25668);
nor U26120 (N_26120,N_25525,N_25769);
nand U26121 (N_26121,N_25973,N_25614);
and U26122 (N_26122,N_25876,N_25747);
xor U26123 (N_26123,N_25539,N_25815);
xnor U26124 (N_26124,N_25583,N_25515);
nand U26125 (N_26125,N_25840,N_25814);
nand U26126 (N_26126,N_25888,N_25952);
nand U26127 (N_26127,N_25960,N_25871);
nand U26128 (N_26128,N_25989,N_25912);
nor U26129 (N_26129,N_25838,N_25924);
xnor U26130 (N_26130,N_25581,N_25969);
or U26131 (N_26131,N_25919,N_25688);
nand U26132 (N_26132,N_25743,N_25782);
nand U26133 (N_26133,N_25526,N_25634);
nand U26134 (N_26134,N_25970,N_25923);
nor U26135 (N_26135,N_25870,N_25748);
or U26136 (N_26136,N_25742,N_25847);
or U26137 (N_26137,N_25650,N_25920);
nor U26138 (N_26138,N_25597,N_25939);
or U26139 (N_26139,N_25641,N_25925);
or U26140 (N_26140,N_25543,N_25693);
or U26141 (N_26141,N_25589,N_25638);
xnor U26142 (N_26142,N_25519,N_25541);
and U26143 (N_26143,N_25630,N_25770);
or U26144 (N_26144,N_25729,N_25821);
xnor U26145 (N_26145,N_25517,N_25532);
nand U26146 (N_26146,N_25863,N_25956);
and U26147 (N_26147,N_25512,N_25854);
or U26148 (N_26148,N_25653,N_25944);
xor U26149 (N_26149,N_25833,N_25824);
or U26150 (N_26150,N_25556,N_25905);
and U26151 (N_26151,N_25979,N_25908);
nor U26152 (N_26152,N_25655,N_25819);
or U26153 (N_26153,N_25933,N_25881);
nor U26154 (N_26154,N_25579,N_25911);
or U26155 (N_26155,N_25906,N_25971);
and U26156 (N_26156,N_25708,N_25660);
nand U26157 (N_26157,N_25734,N_25637);
or U26158 (N_26158,N_25715,N_25918);
xnor U26159 (N_26159,N_25674,N_25531);
nor U26160 (N_26160,N_25832,N_25846);
nor U26161 (N_26161,N_25714,N_25809);
or U26162 (N_26162,N_25504,N_25603);
and U26163 (N_26163,N_25891,N_25675);
nand U26164 (N_26164,N_25647,N_25986);
or U26165 (N_26165,N_25992,N_25850);
nand U26166 (N_26166,N_25524,N_25632);
and U26167 (N_26167,N_25963,N_25564);
xor U26168 (N_26168,N_25633,N_25934);
nand U26169 (N_26169,N_25712,N_25967);
nand U26170 (N_26170,N_25803,N_25765);
or U26171 (N_26171,N_25696,N_25991);
and U26172 (N_26172,N_25783,N_25669);
xor U26173 (N_26173,N_25520,N_25766);
or U26174 (N_26174,N_25893,N_25616);
xor U26175 (N_26175,N_25540,N_25513);
nand U26176 (N_26176,N_25707,N_25978);
or U26177 (N_26177,N_25855,N_25700);
nor U26178 (N_26178,N_25800,N_25536);
nor U26179 (N_26179,N_25872,N_25602);
nor U26180 (N_26180,N_25665,N_25502);
nand U26181 (N_26181,N_25702,N_25746);
xnor U26182 (N_26182,N_25949,N_25807);
and U26183 (N_26183,N_25705,N_25558);
or U26184 (N_26184,N_25786,N_25687);
or U26185 (N_26185,N_25582,N_25851);
and U26186 (N_26186,N_25501,N_25980);
nand U26187 (N_26187,N_25698,N_25676);
xnor U26188 (N_26188,N_25759,N_25984);
and U26189 (N_26189,N_25794,N_25913);
nand U26190 (N_26190,N_25951,N_25628);
and U26191 (N_26191,N_25995,N_25928);
and U26192 (N_26192,N_25940,N_25569);
nand U26193 (N_26193,N_25611,N_25591);
xnor U26194 (N_26194,N_25680,N_25844);
or U26195 (N_26195,N_25987,N_25725);
or U26196 (N_26196,N_25535,N_25695);
nand U26197 (N_26197,N_25521,N_25685);
and U26198 (N_26198,N_25735,N_25999);
and U26199 (N_26199,N_25897,N_25889);
and U26200 (N_26200,N_25761,N_25796);
or U26201 (N_26201,N_25764,N_25955);
nand U26202 (N_26202,N_25654,N_25527);
nand U26203 (N_26203,N_25779,N_25845);
nor U26204 (N_26204,N_25567,N_25841);
and U26205 (N_26205,N_25720,N_25594);
and U26206 (N_26206,N_25751,N_25941);
and U26207 (N_26207,N_25975,N_25624);
xor U26208 (N_26208,N_25894,N_25639);
nor U26209 (N_26209,N_25716,N_25812);
xor U26210 (N_26210,N_25836,N_25959);
and U26211 (N_26211,N_25901,N_25721);
nand U26212 (N_26212,N_25619,N_25682);
nor U26213 (N_26213,N_25749,N_25830);
or U26214 (N_26214,N_25816,N_25610);
nand U26215 (N_26215,N_25990,N_25822);
or U26216 (N_26216,N_25666,N_25900);
nand U26217 (N_26217,N_25733,N_25828);
nor U26218 (N_26218,N_25559,N_25672);
nand U26219 (N_26219,N_25827,N_25842);
xor U26220 (N_26220,N_25904,N_25555);
xor U26221 (N_26221,N_25612,N_25530);
nor U26222 (N_26222,N_25533,N_25778);
nand U26223 (N_26223,N_25621,N_25964);
nor U26224 (N_26224,N_25791,N_25563);
xor U26225 (N_26225,N_25550,N_25789);
or U26226 (N_26226,N_25910,N_25966);
or U26227 (N_26227,N_25584,N_25785);
nand U26228 (N_26228,N_25996,N_25873);
or U26229 (N_26229,N_25510,N_25683);
and U26230 (N_26230,N_25866,N_25887);
or U26231 (N_26231,N_25760,N_25529);
nand U26232 (N_26232,N_25570,N_25927);
nor U26233 (N_26233,N_25547,N_25508);
and U26234 (N_26234,N_25503,N_25874);
and U26235 (N_26235,N_25548,N_25817);
and U26236 (N_26236,N_25750,N_25834);
xor U26237 (N_26237,N_25593,N_25534);
nor U26238 (N_26238,N_25825,N_25646);
or U26239 (N_26239,N_25649,N_25737);
or U26240 (N_26240,N_25557,N_25916);
nor U26241 (N_26241,N_25965,N_25528);
nand U26242 (N_26242,N_25790,N_25571);
xor U26243 (N_26243,N_25837,N_25860);
nand U26244 (N_26244,N_25722,N_25914);
nand U26245 (N_26245,N_25689,N_25671);
nand U26246 (N_26246,N_25598,N_25953);
or U26247 (N_26247,N_25506,N_25788);
or U26248 (N_26248,N_25777,N_25551);
nor U26249 (N_26249,N_25537,N_25882);
xnor U26250 (N_26250,N_25757,N_25891);
and U26251 (N_26251,N_25611,N_25692);
nand U26252 (N_26252,N_25636,N_25634);
nand U26253 (N_26253,N_25916,N_25839);
xnor U26254 (N_26254,N_25867,N_25642);
nor U26255 (N_26255,N_25795,N_25784);
or U26256 (N_26256,N_25852,N_25854);
or U26257 (N_26257,N_25764,N_25821);
and U26258 (N_26258,N_25631,N_25853);
and U26259 (N_26259,N_25679,N_25613);
and U26260 (N_26260,N_25563,N_25514);
xnor U26261 (N_26261,N_25528,N_25738);
nand U26262 (N_26262,N_25905,N_25874);
nand U26263 (N_26263,N_25944,N_25584);
nor U26264 (N_26264,N_25775,N_25530);
or U26265 (N_26265,N_25586,N_25644);
nor U26266 (N_26266,N_25858,N_25962);
xnor U26267 (N_26267,N_25752,N_25988);
and U26268 (N_26268,N_25727,N_25698);
nor U26269 (N_26269,N_25680,N_25534);
nor U26270 (N_26270,N_25731,N_25700);
nor U26271 (N_26271,N_25961,N_25929);
nor U26272 (N_26272,N_25728,N_25951);
xor U26273 (N_26273,N_25995,N_25835);
xor U26274 (N_26274,N_25716,N_25534);
nor U26275 (N_26275,N_25650,N_25822);
xnor U26276 (N_26276,N_25583,N_25815);
nor U26277 (N_26277,N_25602,N_25807);
nand U26278 (N_26278,N_25777,N_25840);
nand U26279 (N_26279,N_25511,N_25950);
nand U26280 (N_26280,N_25732,N_25632);
and U26281 (N_26281,N_25940,N_25899);
or U26282 (N_26282,N_25522,N_25691);
or U26283 (N_26283,N_25971,N_25579);
xor U26284 (N_26284,N_25726,N_25806);
and U26285 (N_26285,N_25509,N_25886);
xor U26286 (N_26286,N_25787,N_25845);
nand U26287 (N_26287,N_25565,N_25650);
nor U26288 (N_26288,N_25640,N_25787);
xor U26289 (N_26289,N_25663,N_25759);
xnor U26290 (N_26290,N_25836,N_25710);
and U26291 (N_26291,N_25594,N_25807);
and U26292 (N_26292,N_25798,N_25592);
or U26293 (N_26293,N_25875,N_25541);
xnor U26294 (N_26294,N_25548,N_25932);
nand U26295 (N_26295,N_25820,N_25967);
and U26296 (N_26296,N_25939,N_25908);
xnor U26297 (N_26297,N_25888,N_25911);
and U26298 (N_26298,N_25942,N_25707);
and U26299 (N_26299,N_25967,N_25681);
or U26300 (N_26300,N_25701,N_25960);
xor U26301 (N_26301,N_25926,N_25630);
nand U26302 (N_26302,N_25866,N_25945);
and U26303 (N_26303,N_25834,N_25856);
and U26304 (N_26304,N_25586,N_25562);
nor U26305 (N_26305,N_25663,N_25835);
nor U26306 (N_26306,N_25760,N_25669);
and U26307 (N_26307,N_25703,N_25604);
nand U26308 (N_26308,N_25702,N_25624);
xnor U26309 (N_26309,N_25995,N_25982);
or U26310 (N_26310,N_25712,N_25724);
nor U26311 (N_26311,N_25922,N_25558);
and U26312 (N_26312,N_25599,N_25997);
nand U26313 (N_26313,N_25769,N_25797);
and U26314 (N_26314,N_25972,N_25832);
and U26315 (N_26315,N_25972,N_25913);
or U26316 (N_26316,N_25544,N_25688);
and U26317 (N_26317,N_25692,N_25634);
or U26318 (N_26318,N_25884,N_25602);
nand U26319 (N_26319,N_25581,N_25840);
nor U26320 (N_26320,N_25989,N_25668);
nor U26321 (N_26321,N_25621,N_25532);
and U26322 (N_26322,N_25981,N_25664);
xor U26323 (N_26323,N_25845,N_25663);
nor U26324 (N_26324,N_25791,N_25609);
nand U26325 (N_26325,N_25829,N_25783);
or U26326 (N_26326,N_25896,N_25573);
or U26327 (N_26327,N_25672,N_25752);
xnor U26328 (N_26328,N_25532,N_25555);
xnor U26329 (N_26329,N_25946,N_25582);
or U26330 (N_26330,N_25907,N_25505);
or U26331 (N_26331,N_25674,N_25792);
or U26332 (N_26332,N_25769,N_25682);
and U26333 (N_26333,N_25741,N_25648);
xor U26334 (N_26334,N_25965,N_25620);
or U26335 (N_26335,N_25629,N_25698);
xnor U26336 (N_26336,N_25779,N_25866);
nor U26337 (N_26337,N_25862,N_25930);
xnor U26338 (N_26338,N_25522,N_25952);
xnor U26339 (N_26339,N_25704,N_25562);
xor U26340 (N_26340,N_25900,N_25756);
nor U26341 (N_26341,N_25676,N_25591);
nor U26342 (N_26342,N_25736,N_25561);
or U26343 (N_26343,N_25950,N_25651);
and U26344 (N_26344,N_25954,N_25874);
nor U26345 (N_26345,N_25993,N_25956);
xor U26346 (N_26346,N_25683,N_25663);
nand U26347 (N_26347,N_25556,N_25790);
or U26348 (N_26348,N_25693,N_25765);
and U26349 (N_26349,N_25879,N_25691);
xnor U26350 (N_26350,N_25762,N_25770);
and U26351 (N_26351,N_25918,N_25842);
and U26352 (N_26352,N_25871,N_25675);
or U26353 (N_26353,N_25645,N_25512);
nand U26354 (N_26354,N_25516,N_25601);
and U26355 (N_26355,N_25546,N_25906);
nand U26356 (N_26356,N_25741,N_25540);
and U26357 (N_26357,N_25790,N_25578);
or U26358 (N_26358,N_25639,N_25733);
or U26359 (N_26359,N_25819,N_25770);
or U26360 (N_26360,N_25837,N_25629);
or U26361 (N_26361,N_25515,N_25940);
nand U26362 (N_26362,N_25801,N_25813);
or U26363 (N_26363,N_25726,N_25748);
xor U26364 (N_26364,N_25676,N_25516);
or U26365 (N_26365,N_25811,N_25838);
and U26366 (N_26366,N_25669,N_25520);
nor U26367 (N_26367,N_25572,N_25558);
nand U26368 (N_26368,N_25564,N_25930);
or U26369 (N_26369,N_25983,N_25875);
xnor U26370 (N_26370,N_25610,N_25846);
or U26371 (N_26371,N_25705,N_25858);
nor U26372 (N_26372,N_25679,N_25871);
nor U26373 (N_26373,N_25553,N_25666);
or U26374 (N_26374,N_25862,N_25768);
xnor U26375 (N_26375,N_25788,N_25752);
nand U26376 (N_26376,N_25904,N_25548);
nand U26377 (N_26377,N_25637,N_25756);
or U26378 (N_26378,N_25836,N_25556);
xor U26379 (N_26379,N_25502,N_25925);
or U26380 (N_26380,N_25666,N_25818);
nand U26381 (N_26381,N_25553,N_25911);
nor U26382 (N_26382,N_25885,N_25785);
nor U26383 (N_26383,N_25893,N_25839);
and U26384 (N_26384,N_25816,N_25947);
and U26385 (N_26385,N_25940,N_25523);
or U26386 (N_26386,N_25819,N_25825);
xor U26387 (N_26387,N_25668,N_25602);
xnor U26388 (N_26388,N_25619,N_25627);
nor U26389 (N_26389,N_25713,N_25581);
or U26390 (N_26390,N_25529,N_25710);
nand U26391 (N_26391,N_25508,N_25555);
xor U26392 (N_26392,N_25501,N_25526);
nor U26393 (N_26393,N_25765,N_25997);
nand U26394 (N_26394,N_25663,N_25598);
and U26395 (N_26395,N_25706,N_25540);
and U26396 (N_26396,N_25751,N_25826);
nand U26397 (N_26397,N_25982,N_25726);
and U26398 (N_26398,N_25798,N_25736);
nand U26399 (N_26399,N_25797,N_25662);
nor U26400 (N_26400,N_25587,N_25828);
nor U26401 (N_26401,N_25583,N_25899);
xor U26402 (N_26402,N_25737,N_25844);
nand U26403 (N_26403,N_25823,N_25601);
or U26404 (N_26404,N_25549,N_25841);
xor U26405 (N_26405,N_25742,N_25575);
or U26406 (N_26406,N_25919,N_25680);
or U26407 (N_26407,N_25625,N_25929);
xnor U26408 (N_26408,N_25809,N_25894);
or U26409 (N_26409,N_25811,N_25815);
nand U26410 (N_26410,N_25971,N_25531);
nor U26411 (N_26411,N_25665,N_25725);
or U26412 (N_26412,N_25729,N_25819);
and U26413 (N_26413,N_25561,N_25647);
xnor U26414 (N_26414,N_25926,N_25878);
nand U26415 (N_26415,N_25964,N_25945);
or U26416 (N_26416,N_25751,N_25983);
nor U26417 (N_26417,N_25516,N_25700);
nand U26418 (N_26418,N_25989,N_25830);
xor U26419 (N_26419,N_25573,N_25963);
and U26420 (N_26420,N_25755,N_25793);
xnor U26421 (N_26421,N_25793,N_25865);
or U26422 (N_26422,N_25986,N_25786);
or U26423 (N_26423,N_25904,N_25575);
or U26424 (N_26424,N_25806,N_25977);
nand U26425 (N_26425,N_25933,N_25879);
and U26426 (N_26426,N_25568,N_25523);
xor U26427 (N_26427,N_25786,N_25606);
or U26428 (N_26428,N_25653,N_25586);
nand U26429 (N_26429,N_25530,N_25932);
nand U26430 (N_26430,N_25649,N_25917);
or U26431 (N_26431,N_25798,N_25513);
nor U26432 (N_26432,N_25579,N_25739);
or U26433 (N_26433,N_25992,N_25626);
or U26434 (N_26434,N_25826,N_25892);
or U26435 (N_26435,N_25903,N_25893);
and U26436 (N_26436,N_25627,N_25841);
and U26437 (N_26437,N_25781,N_25834);
nor U26438 (N_26438,N_25557,N_25821);
xnor U26439 (N_26439,N_25697,N_25559);
or U26440 (N_26440,N_25534,N_25607);
and U26441 (N_26441,N_25828,N_25832);
nand U26442 (N_26442,N_25577,N_25754);
or U26443 (N_26443,N_25978,N_25708);
nor U26444 (N_26444,N_25954,N_25603);
nor U26445 (N_26445,N_25737,N_25510);
nor U26446 (N_26446,N_25982,N_25799);
and U26447 (N_26447,N_25550,N_25949);
xor U26448 (N_26448,N_25612,N_25727);
and U26449 (N_26449,N_25560,N_25991);
xnor U26450 (N_26450,N_25647,N_25514);
or U26451 (N_26451,N_25959,N_25879);
and U26452 (N_26452,N_25518,N_25922);
nand U26453 (N_26453,N_25767,N_25686);
xor U26454 (N_26454,N_25972,N_25956);
xnor U26455 (N_26455,N_25987,N_25909);
or U26456 (N_26456,N_25709,N_25974);
nor U26457 (N_26457,N_25806,N_25750);
or U26458 (N_26458,N_25680,N_25784);
nor U26459 (N_26459,N_25562,N_25529);
and U26460 (N_26460,N_25722,N_25807);
nand U26461 (N_26461,N_25941,N_25793);
or U26462 (N_26462,N_25978,N_25692);
and U26463 (N_26463,N_25709,N_25574);
nand U26464 (N_26464,N_25927,N_25818);
or U26465 (N_26465,N_25732,N_25992);
xor U26466 (N_26466,N_25610,N_25699);
nand U26467 (N_26467,N_25946,N_25681);
nor U26468 (N_26468,N_25867,N_25641);
and U26469 (N_26469,N_25800,N_25913);
or U26470 (N_26470,N_25643,N_25854);
xnor U26471 (N_26471,N_25670,N_25792);
and U26472 (N_26472,N_25949,N_25543);
or U26473 (N_26473,N_25528,N_25931);
nand U26474 (N_26474,N_25966,N_25545);
or U26475 (N_26475,N_25651,N_25855);
and U26476 (N_26476,N_25957,N_25714);
xnor U26477 (N_26477,N_25521,N_25893);
and U26478 (N_26478,N_25690,N_25675);
nand U26479 (N_26479,N_25650,N_25849);
nand U26480 (N_26480,N_25938,N_25807);
nor U26481 (N_26481,N_25996,N_25541);
or U26482 (N_26482,N_25867,N_25849);
or U26483 (N_26483,N_25657,N_25752);
nand U26484 (N_26484,N_25569,N_25946);
nand U26485 (N_26485,N_25943,N_25763);
nor U26486 (N_26486,N_25873,N_25777);
nand U26487 (N_26487,N_25675,N_25663);
nor U26488 (N_26488,N_25787,N_25888);
nand U26489 (N_26489,N_25595,N_25707);
nor U26490 (N_26490,N_25647,N_25689);
and U26491 (N_26491,N_25748,N_25555);
nor U26492 (N_26492,N_25657,N_25677);
or U26493 (N_26493,N_25956,N_25597);
nor U26494 (N_26494,N_25544,N_25840);
nor U26495 (N_26495,N_25799,N_25981);
and U26496 (N_26496,N_25647,N_25628);
xnor U26497 (N_26497,N_25623,N_25708);
nor U26498 (N_26498,N_25872,N_25890);
or U26499 (N_26499,N_25813,N_25510);
nand U26500 (N_26500,N_26043,N_26069);
xnor U26501 (N_26501,N_26284,N_26101);
xnor U26502 (N_26502,N_26116,N_26218);
nand U26503 (N_26503,N_26119,N_26251);
nand U26504 (N_26504,N_26370,N_26021);
or U26505 (N_26505,N_26399,N_26011);
or U26506 (N_26506,N_26080,N_26224);
or U26507 (N_26507,N_26219,N_26157);
nor U26508 (N_26508,N_26203,N_26296);
nand U26509 (N_26509,N_26368,N_26003);
or U26510 (N_26510,N_26372,N_26432);
and U26511 (N_26511,N_26105,N_26316);
nand U26512 (N_26512,N_26235,N_26250);
and U26513 (N_26513,N_26115,N_26002);
and U26514 (N_26514,N_26320,N_26163);
xor U26515 (N_26515,N_26268,N_26100);
nand U26516 (N_26516,N_26494,N_26153);
or U26517 (N_26517,N_26177,N_26306);
or U26518 (N_26518,N_26067,N_26242);
nand U26519 (N_26519,N_26089,N_26364);
xnor U26520 (N_26520,N_26376,N_26385);
and U26521 (N_26521,N_26146,N_26197);
and U26522 (N_26522,N_26274,N_26110);
or U26523 (N_26523,N_26038,N_26048);
or U26524 (N_26524,N_26142,N_26132);
or U26525 (N_26525,N_26404,N_26188);
nand U26526 (N_26526,N_26378,N_26304);
and U26527 (N_26527,N_26314,N_26059);
and U26528 (N_26528,N_26046,N_26448);
nand U26529 (N_26529,N_26111,N_26392);
nor U26530 (N_26530,N_26103,N_26033);
or U26531 (N_26531,N_26057,N_26439);
nor U26532 (N_26532,N_26200,N_26366);
or U26533 (N_26533,N_26010,N_26393);
and U26534 (N_26534,N_26354,N_26441);
nor U26535 (N_26535,N_26294,N_26278);
or U26536 (N_26536,N_26211,N_26303);
and U26537 (N_26537,N_26361,N_26324);
xnor U26538 (N_26538,N_26254,N_26359);
nor U26539 (N_26539,N_26257,N_26036);
xnor U26540 (N_26540,N_26126,N_26217);
or U26541 (N_26541,N_26222,N_26071);
nor U26542 (N_26542,N_26493,N_26151);
or U26543 (N_26543,N_26201,N_26076);
nand U26544 (N_26544,N_26438,N_26390);
and U26545 (N_26545,N_26081,N_26206);
xor U26546 (N_26546,N_26476,N_26266);
nand U26547 (N_26547,N_26434,N_26141);
nand U26548 (N_26548,N_26326,N_26283);
nand U26549 (N_26549,N_26156,N_26430);
or U26550 (N_26550,N_26214,N_26220);
nor U26551 (N_26551,N_26459,N_26295);
and U26552 (N_26552,N_26065,N_26144);
nor U26553 (N_26553,N_26102,N_26315);
or U26554 (N_26554,N_26469,N_26427);
and U26555 (N_26555,N_26467,N_26353);
nand U26556 (N_26556,N_26079,N_26092);
nor U26557 (N_26557,N_26025,N_26062);
or U26558 (N_26558,N_26078,N_26009);
or U26559 (N_26559,N_26223,N_26299);
and U26560 (N_26560,N_26475,N_26253);
and U26561 (N_26561,N_26305,N_26377);
nor U26562 (N_26562,N_26258,N_26408);
or U26563 (N_26563,N_26247,N_26014);
nand U26564 (N_26564,N_26168,N_26400);
or U26565 (N_26565,N_26090,N_26122);
and U26566 (N_26566,N_26277,N_26117);
nor U26567 (N_26567,N_26487,N_26174);
nor U26568 (N_26568,N_26421,N_26241);
nand U26569 (N_26569,N_26155,N_26331);
xor U26570 (N_26570,N_26027,N_26125);
xnor U26571 (N_26571,N_26474,N_26281);
xnor U26572 (N_26572,N_26419,N_26016);
and U26573 (N_26573,N_26170,N_26233);
or U26574 (N_26574,N_26489,N_26345);
and U26575 (N_26575,N_26273,N_26275);
nor U26576 (N_26576,N_26171,N_26436);
nor U26577 (N_26577,N_26066,N_26360);
nand U26578 (N_26578,N_26321,N_26135);
xnor U26579 (N_26579,N_26402,N_26019);
xnor U26580 (N_26580,N_26196,N_26232);
and U26581 (N_26581,N_26208,N_26029);
and U26582 (N_26582,N_26347,N_26417);
and U26583 (N_26583,N_26334,N_26446);
nor U26584 (N_26584,N_26030,N_26073);
and U26585 (N_26585,N_26020,N_26215);
nor U26586 (N_26586,N_26087,N_26121);
and U26587 (N_26587,N_26388,N_26428);
and U26588 (N_26588,N_26282,N_26382);
nand U26589 (N_26589,N_26383,N_26271);
and U26590 (N_26590,N_26483,N_26423);
xnor U26591 (N_26591,N_26246,N_26108);
xnor U26592 (N_26592,N_26272,N_26063);
xnor U26593 (N_26593,N_26140,N_26058);
and U26594 (N_26594,N_26128,N_26239);
and U26595 (N_26595,N_26145,N_26228);
or U26596 (N_26596,N_26074,N_26351);
nand U26597 (N_26597,N_26172,N_26431);
or U26598 (N_26598,N_26006,N_26072);
nor U26599 (N_26599,N_26379,N_26084);
and U26600 (N_26600,N_26182,N_26317);
and U26601 (N_26601,N_26449,N_26358);
xor U26602 (N_26602,N_26452,N_26435);
or U26603 (N_26603,N_26056,N_26471);
nand U26604 (N_26604,N_26261,N_26007);
and U26605 (N_26605,N_26028,N_26231);
nand U26606 (N_26606,N_26330,N_26470);
or U26607 (N_26607,N_26210,N_26094);
and U26608 (N_26608,N_26131,N_26134);
or U26609 (N_26609,N_26138,N_26042);
nor U26610 (N_26610,N_26096,N_26327);
or U26611 (N_26611,N_26447,N_26082);
nand U26612 (N_26612,N_26085,N_26098);
nand U26613 (N_26613,N_26004,N_26070);
nand U26614 (N_26614,N_26396,N_26106);
nor U26615 (N_26615,N_26238,N_26161);
nor U26616 (N_26616,N_26104,N_26492);
and U26617 (N_26617,N_26279,N_26124);
or U26618 (N_26618,N_26307,N_26114);
xnor U26619 (N_26619,N_26175,N_26407);
or U26620 (N_26620,N_26276,N_26191);
nor U26621 (N_26621,N_26460,N_26041);
and U26622 (N_26622,N_26367,N_26194);
nand U26623 (N_26623,N_26363,N_26462);
nand U26624 (N_26624,N_26164,N_26183);
nor U26625 (N_26625,N_26213,N_26384);
xnor U26626 (N_26626,N_26323,N_26484);
nor U26627 (N_26627,N_26259,N_26312);
xnor U26628 (N_26628,N_26380,N_26290);
or U26629 (N_26629,N_26234,N_26158);
xor U26630 (N_26630,N_26147,N_26394);
xor U26631 (N_26631,N_26466,N_26237);
nor U26632 (N_26632,N_26189,N_26107);
nor U26633 (N_26633,N_26249,N_26221);
nand U26634 (N_26634,N_26185,N_26022);
nor U26635 (N_26635,N_26485,N_26015);
or U26636 (N_26636,N_26187,N_26287);
and U26637 (N_26637,N_26472,N_26420);
nor U26638 (N_26638,N_26297,N_26288);
or U26639 (N_26639,N_26389,N_26205);
or U26640 (N_26640,N_26301,N_26005);
xnor U26641 (N_26641,N_26053,N_26395);
or U26642 (N_26642,N_26293,N_26473);
nor U26643 (N_26643,N_26083,N_26350);
nor U26644 (N_26644,N_26289,N_26055);
or U26645 (N_26645,N_26349,N_26075);
and U26646 (N_26646,N_26365,N_26403);
nor U26647 (N_26647,N_26012,N_26461);
nor U26648 (N_26648,N_26176,N_26302);
nor U26649 (N_26649,N_26190,N_26456);
nand U26650 (N_26650,N_26442,N_26424);
xor U26651 (N_26651,N_26165,N_26127);
nor U26652 (N_26652,N_26008,N_26341);
xnor U26653 (N_26653,N_26478,N_26267);
nor U26654 (N_26654,N_26137,N_26202);
xor U26655 (N_26655,N_26371,N_26412);
xor U26656 (N_26656,N_26418,N_26387);
and U26657 (N_26657,N_26498,N_26497);
and U26658 (N_26658,N_26488,N_26454);
and U26659 (N_26659,N_26269,N_26047);
nor U26660 (N_26660,N_26225,N_26465);
or U26661 (N_26661,N_26413,N_26313);
and U26662 (N_26662,N_26118,N_26437);
xnor U26663 (N_26663,N_26335,N_26243);
nor U26664 (N_26664,N_26180,N_26166);
xnor U26665 (N_26665,N_26409,N_26322);
xor U26666 (N_26666,N_26130,N_26344);
nor U26667 (N_26667,N_26286,N_26061);
nand U26668 (N_26668,N_26209,N_26248);
nand U26669 (N_26669,N_26255,N_26356);
or U26670 (N_26670,N_26023,N_26049);
nand U26671 (N_26671,N_26481,N_26052);
or U26672 (N_26672,N_26309,N_26149);
nand U26673 (N_26673,N_26308,N_26032);
nor U26674 (N_26674,N_26328,N_26285);
and U26675 (N_26675,N_26491,N_26329);
or U26676 (N_26676,N_26280,N_26026);
and U26677 (N_26677,N_26455,N_26477);
xnor U26678 (N_26678,N_26397,N_26337);
nor U26679 (N_26679,N_26212,N_26216);
nand U26680 (N_26680,N_26192,N_26148);
nand U26681 (N_26681,N_26088,N_26482);
nor U26682 (N_26682,N_26109,N_26339);
or U26683 (N_26683,N_26433,N_26207);
or U26684 (N_26684,N_26486,N_26357);
nor U26685 (N_26685,N_26263,N_26318);
and U26686 (N_26686,N_26369,N_26264);
nand U26687 (N_26687,N_26453,N_26120);
nor U26688 (N_26688,N_26300,N_26480);
nand U26689 (N_26689,N_26373,N_26136);
nand U26690 (N_26690,N_26310,N_26193);
nor U26691 (N_26691,N_26355,N_26195);
or U26692 (N_26692,N_26425,N_26450);
nor U26693 (N_26693,N_26457,N_26252);
or U26694 (N_26694,N_26129,N_26298);
xnor U26695 (N_26695,N_26152,N_26463);
nand U26696 (N_26696,N_26319,N_26181);
xor U26697 (N_26697,N_26143,N_26154);
nand U26698 (N_26698,N_26086,N_26270);
xor U26699 (N_26699,N_26375,N_26338);
and U26700 (N_26700,N_26244,N_26150);
and U26701 (N_26701,N_26227,N_26226);
nor U26702 (N_26702,N_26240,N_26113);
nor U26703 (N_26703,N_26422,N_26311);
xnor U26704 (N_26704,N_26416,N_26405);
and U26705 (N_26705,N_26458,N_26000);
nand U26706 (N_26706,N_26037,N_26346);
nor U26707 (N_26707,N_26068,N_26381);
nor U26708 (N_26708,N_26001,N_26236);
and U26709 (N_26709,N_26013,N_26401);
xor U26710 (N_26710,N_26451,N_26044);
nor U26711 (N_26711,N_26410,N_26179);
and U26712 (N_26712,N_26443,N_26468);
nor U26713 (N_26713,N_26426,N_26045);
nand U26714 (N_26714,N_26095,N_26051);
nand U26715 (N_26715,N_26093,N_26352);
nand U26716 (N_26716,N_26204,N_26265);
nand U26717 (N_26717,N_26050,N_26333);
nand U26718 (N_26718,N_26018,N_26340);
or U26719 (N_26719,N_26374,N_26262);
nor U26720 (N_26720,N_26444,N_26160);
or U26721 (N_26721,N_26325,N_26054);
xor U26722 (N_26722,N_26440,N_26479);
or U26723 (N_26723,N_26167,N_26464);
and U26724 (N_26724,N_26229,N_26411);
or U26725 (N_26725,N_26024,N_26292);
or U26726 (N_26726,N_26332,N_26034);
nor U26727 (N_26727,N_26077,N_26184);
or U26728 (N_26728,N_26245,N_26348);
nand U26729 (N_26729,N_26391,N_26414);
nand U26730 (N_26730,N_26039,N_26260);
nand U26731 (N_26731,N_26031,N_26112);
nand U26732 (N_26732,N_26343,N_26178);
nor U26733 (N_26733,N_26133,N_26199);
nor U26734 (N_26734,N_26035,N_26064);
or U26735 (N_26735,N_26186,N_26099);
nand U26736 (N_26736,N_26060,N_26162);
nand U26737 (N_26737,N_26499,N_26342);
and U26738 (N_26738,N_26198,N_26159);
and U26739 (N_26739,N_26490,N_26291);
nor U26740 (N_26740,N_26398,N_26097);
and U26741 (N_26741,N_26406,N_26123);
nor U26742 (N_26742,N_26415,N_26429);
nand U26743 (N_26743,N_26386,N_26336);
and U26744 (N_26744,N_26169,N_26230);
or U26745 (N_26745,N_26017,N_26445);
nand U26746 (N_26746,N_26173,N_26495);
or U26747 (N_26747,N_26091,N_26139);
nor U26748 (N_26748,N_26040,N_26496);
nand U26749 (N_26749,N_26362,N_26256);
xor U26750 (N_26750,N_26159,N_26167);
xor U26751 (N_26751,N_26181,N_26251);
nand U26752 (N_26752,N_26164,N_26416);
xor U26753 (N_26753,N_26403,N_26374);
xnor U26754 (N_26754,N_26179,N_26347);
and U26755 (N_26755,N_26246,N_26457);
and U26756 (N_26756,N_26339,N_26016);
xnor U26757 (N_26757,N_26243,N_26170);
nand U26758 (N_26758,N_26207,N_26034);
nor U26759 (N_26759,N_26482,N_26473);
or U26760 (N_26760,N_26028,N_26206);
nand U26761 (N_26761,N_26092,N_26326);
or U26762 (N_26762,N_26337,N_26263);
or U26763 (N_26763,N_26048,N_26311);
nor U26764 (N_26764,N_26406,N_26497);
nor U26765 (N_26765,N_26212,N_26456);
nor U26766 (N_26766,N_26451,N_26448);
xnor U26767 (N_26767,N_26409,N_26196);
xnor U26768 (N_26768,N_26260,N_26113);
nand U26769 (N_26769,N_26338,N_26410);
xnor U26770 (N_26770,N_26404,N_26032);
nor U26771 (N_26771,N_26194,N_26027);
nand U26772 (N_26772,N_26332,N_26023);
xnor U26773 (N_26773,N_26350,N_26440);
and U26774 (N_26774,N_26190,N_26243);
xor U26775 (N_26775,N_26158,N_26142);
nand U26776 (N_26776,N_26303,N_26193);
xnor U26777 (N_26777,N_26258,N_26136);
and U26778 (N_26778,N_26288,N_26483);
xnor U26779 (N_26779,N_26327,N_26333);
nand U26780 (N_26780,N_26301,N_26041);
and U26781 (N_26781,N_26480,N_26074);
nor U26782 (N_26782,N_26477,N_26365);
xnor U26783 (N_26783,N_26261,N_26273);
xnor U26784 (N_26784,N_26224,N_26407);
xor U26785 (N_26785,N_26471,N_26014);
nor U26786 (N_26786,N_26266,N_26386);
or U26787 (N_26787,N_26110,N_26237);
and U26788 (N_26788,N_26311,N_26166);
nand U26789 (N_26789,N_26117,N_26054);
and U26790 (N_26790,N_26019,N_26138);
xor U26791 (N_26791,N_26107,N_26024);
and U26792 (N_26792,N_26408,N_26270);
nor U26793 (N_26793,N_26487,N_26057);
nand U26794 (N_26794,N_26283,N_26481);
or U26795 (N_26795,N_26274,N_26212);
xor U26796 (N_26796,N_26433,N_26473);
nand U26797 (N_26797,N_26491,N_26486);
or U26798 (N_26798,N_26116,N_26467);
or U26799 (N_26799,N_26218,N_26226);
nand U26800 (N_26800,N_26227,N_26126);
or U26801 (N_26801,N_26078,N_26093);
nor U26802 (N_26802,N_26244,N_26360);
and U26803 (N_26803,N_26284,N_26129);
and U26804 (N_26804,N_26024,N_26190);
nand U26805 (N_26805,N_26057,N_26355);
xnor U26806 (N_26806,N_26015,N_26055);
or U26807 (N_26807,N_26196,N_26356);
nand U26808 (N_26808,N_26481,N_26450);
and U26809 (N_26809,N_26096,N_26163);
or U26810 (N_26810,N_26048,N_26262);
nor U26811 (N_26811,N_26440,N_26393);
and U26812 (N_26812,N_26117,N_26213);
and U26813 (N_26813,N_26317,N_26309);
or U26814 (N_26814,N_26361,N_26188);
xnor U26815 (N_26815,N_26035,N_26115);
xnor U26816 (N_26816,N_26203,N_26446);
nand U26817 (N_26817,N_26106,N_26214);
or U26818 (N_26818,N_26012,N_26382);
nor U26819 (N_26819,N_26046,N_26341);
xnor U26820 (N_26820,N_26174,N_26331);
nor U26821 (N_26821,N_26362,N_26098);
nand U26822 (N_26822,N_26358,N_26066);
xnor U26823 (N_26823,N_26132,N_26244);
or U26824 (N_26824,N_26470,N_26425);
nand U26825 (N_26825,N_26149,N_26189);
xor U26826 (N_26826,N_26140,N_26097);
nor U26827 (N_26827,N_26408,N_26409);
nor U26828 (N_26828,N_26014,N_26259);
or U26829 (N_26829,N_26444,N_26431);
and U26830 (N_26830,N_26229,N_26371);
nand U26831 (N_26831,N_26207,N_26216);
xnor U26832 (N_26832,N_26145,N_26075);
or U26833 (N_26833,N_26120,N_26104);
xnor U26834 (N_26834,N_26498,N_26222);
nor U26835 (N_26835,N_26164,N_26299);
nor U26836 (N_26836,N_26406,N_26394);
and U26837 (N_26837,N_26013,N_26485);
nand U26838 (N_26838,N_26442,N_26154);
nor U26839 (N_26839,N_26331,N_26323);
nor U26840 (N_26840,N_26153,N_26343);
and U26841 (N_26841,N_26468,N_26052);
xor U26842 (N_26842,N_26408,N_26219);
nand U26843 (N_26843,N_26086,N_26372);
nor U26844 (N_26844,N_26295,N_26155);
or U26845 (N_26845,N_26322,N_26405);
xnor U26846 (N_26846,N_26325,N_26073);
xor U26847 (N_26847,N_26177,N_26125);
and U26848 (N_26848,N_26366,N_26123);
and U26849 (N_26849,N_26483,N_26140);
nand U26850 (N_26850,N_26049,N_26181);
nand U26851 (N_26851,N_26109,N_26091);
or U26852 (N_26852,N_26394,N_26041);
and U26853 (N_26853,N_26406,N_26140);
nand U26854 (N_26854,N_26445,N_26226);
xor U26855 (N_26855,N_26412,N_26447);
or U26856 (N_26856,N_26232,N_26396);
nor U26857 (N_26857,N_26421,N_26180);
xnor U26858 (N_26858,N_26294,N_26450);
nand U26859 (N_26859,N_26359,N_26418);
xor U26860 (N_26860,N_26003,N_26291);
nand U26861 (N_26861,N_26094,N_26267);
nor U26862 (N_26862,N_26298,N_26396);
xnor U26863 (N_26863,N_26106,N_26045);
xnor U26864 (N_26864,N_26088,N_26248);
or U26865 (N_26865,N_26240,N_26049);
and U26866 (N_26866,N_26395,N_26277);
or U26867 (N_26867,N_26053,N_26351);
or U26868 (N_26868,N_26301,N_26275);
nand U26869 (N_26869,N_26247,N_26336);
nand U26870 (N_26870,N_26360,N_26063);
xor U26871 (N_26871,N_26192,N_26228);
xnor U26872 (N_26872,N_26010,N_26066);
nor U26873 (N_26873,N_26393,N_26326);
or U26874 (N_26874,N_26061,N_26295);
and U26875 (N_26875,N_26486,N_26239);
xnor U26876 (N_26876,N_26304,N_26098);
nor U26877 (N_26877,N_26388,N_26475);
xor U26878 (N_26878,N_26053,N_26209);
and U26879 (N_26879,N_26439,N_26344);
xor U26880 (N_26880,N_26292,N_26299);
xnor U26881 (N_26881,N_26280,N_26062);
or U26882 (N_26882,N_26311,N_26324);
or U26883 (N_26883,N_26215,N_26314);
and U26884 (N_26884,N_26149,N_26099);
nor U26885 (N_26885,N_26390,N_26410);
nand U26886 (N_26886,N_26159,N_26356);
and U26887 (N_26887,N_26499,N_26052);
or U26888 (N_26888,N_26339,N_26335);
xor U26889 (N_26889,N_26377,N_26392);
or U26890 (N_26890,N_26451,N_26222);
xnor U26891 (N_26891,N_26242,N_26392);
nor U26892 (N_26892,N_26283,N_26232);
nand U26893 (N_26893,N_26152,N_26131);
and U26894 (N_26894,N_26049,N_26484);
xor U26895 (N_26895,N_26134,N_26492);
nand U26896 (N_26896,N_26353,N_26242);
and U26897 (N_26897,N_26131,N_26284);
nand U26898 (N_26898,N_26382,N_26338);
or U26899 (N_26899,N_26421,N_26258);
and U26900 (N_26900,N_26272,N_26238);
nor U26901 (N_26901,N_26257,N_26327);
xor U26902 (N_26902,N_26086,N_26185);
nor U26903 (N_26903,N_26435,N_26183);
nor U26904 (N_26904,N_26038,N_26133);
and U26905 (N_26905,N_26139,N_26408);
nor U26906 (N_26906,N_26334,N_26231);
and U26907 (N_26907,N_26150,N_26123);
nor U26908 (N_26908,N_26140,N_26380);
or U26909 (N_26909,N_26354,N_26241);
nand U26910 (N_26910,N_26098,N_26252);
and U26911 (N_26911,N_26485,N_26346);
and U26912 (N_26912,N_26367,N_26031);
and U26913 (N_26913,N_26163,N_26150);
nand U26914 (N_26914,N_26006,N_26391);
nand U26915 (N_26915,N_26489,N_26166);
xnor U26916 (N_26916,N_26065,N_26264);
xor U26917 (N_26917,N_26135,N_26482);
xor U26918 (N_26918,N_26154,N_26150);
or U26919 (N_26919,N_26071,N_26096);
nand U26920 (N_26920,N_26177,N_26335);
or U26921 (N_26921,N_26238,N_26460);
or U26922 (N_26922,N_26206,N_26386);
and U26923 (N_26923,N_26384,N_26215);
or U26924 (N_26924,N_26209,N_26074);
or U26925 (N_26925,N_26039,N_26271);
xnor U26926 (N_26926,N_26346,N_26350);
nand U26927 (N_26927,N_26134,N_26405);
or U26928 (N_26928,N_26002,N_26122);
xor U26929 (N_26929,N_26353,N_26083);
xor U26930 (N_26930,N_26161,N_26328);
nor U26931 (N_26931,N_26481,N_26123);
nor U26932 (N_26932,N_26349,N_26388);
nand U26933 (N_26933,N_26495,N_26213);
and U26934 (N_26934,N_26099,N_26176);
nor U26935 (N_26935,N_26453,N_26423);
xnor U26936 (N_26936,N_26144,N_26206);
nor U26937 (N_26937,N_26294,N_26170);
xor U26938 (N_26938,N_26451,N_26275);
and U26939 (N_26939,N_26080,N_26335);
or U26940 (N_26940,N_26331,N_26438);
nor U26941 (N_26941,N_26430,N_26219);
xnor U26942 (N_26942,N_26399,N_26348);
nand U26943 (N_26943,N_26352,N_26126);
nor U26944 (N_26944,N_26330,N_26392);
xor U26945 (N_26945,N_26279,N_26234);
nand U26946 (N_26946,N_26079,N_26364);
and U26947 (N_26947,N_26099,N_26062);
nor U26948 (N_26948,N_26473,N_26043);
and U26949 (N_26949,N_26461,N_26411);
or U26950 (N_26950,N_26004,N_26237);
nor U26951 (N_26951,N_26132,N_26364);
nor U26952 (N_26952,N_26374,N_26008);
nor U26953 (N_26953,N_26190,N_26331);
and U26954 (N_26954,N_26268,N_26176);
xnor U26955 (N_26955,N_26223,N_26077);
and U26956 (N_26956,N_26288,N_26242);
or U26957 (N_26957,N_26364,N_26428);
xnor U26958 (N_26958,N_26008,N_26058);
or U26959 (N_26959,N_26082,N_26103);
and U26960 (N_26960,N_26284,N_26194);
nand U26961 (N_26961,N_26197,N_26263);
or U26962 (N_26962,N_26055,N_26144);
xor U26963 (N_26963,N_26262,N_26178);
nand U26964 (N_26964,N_26123,N_26268);
or U26965 (N_26965,N_26304,N_26478);
or U26966 (N_26966,N_26193,N_26436);
and U26967 (N_26967,N_26438,N_26445);
or U26968 (N_26968,N_26088,N_26004);
and U26969 (N_26969,N_26485,N_26034);
and U26970 (N_26970,N_26120,N_26286);
nor U26971 (N_26971,N_26444,N_26133);
and U26972 (N_26972,N_26171,N_26111);
nor U26973 (N_26973,N_26340,N_26344);
nand U26974 (N_26974,N_26356,N_26304);
xor U26975 (N_26975,N_26461,N_26404);
nand U26976 (N_26976,N_26427,N_26339);
xor U26977 (N_26977,N_26043,N_26187);
nor U26978 (N_26978,N_26331,N_26145);
or U26979 (N_26979,N_26485,N_26345);
nor U26980 (N_26980,N_26241,N_26457);
or U26981 (N_26981,N_26469,N_26265);
nor U26982 (N_26982,N_26023,N_26438);
or U26983 (N_26983,N_26239,N_26428);
and U26984 (N_26984,N_26379,N_26091);
nand U26985 (N_26985,N_26422,N_26308);
or U26986 (N_26986,N_26498,N_26379);
and U26987 (N_26987,N_26456,N_26063);
nand U26988 (N_26988,N_26033,N_26356);
and U26989 (N_26989,N_26097,N_26004);
xor U26990 (N_26990,N_26158,N_26392);
nor U26991 (N_26991,N_26008,N_26451);
or U26992 (N_26992,N_26062,N_26018);
or U26993 (N_26993,N_26379,N_26408);
nor U26994 (N_26994,N_26380,N_26020);
nor U26995 (N_26995,N_26081,N_26142);
or U26996 (N_26996,N_26495,N_26007);
nand U26997 (N_26997,N_26455,N_26303);
nand U26998 (N_26998,N_26046,N_26224);
or U26999 (N_26999,N_26226,N_26132);
xnor U27000 (N_27000,N_26674,N_26863);
xor U27001 (N_27001,N_26635,N_26943);
xor U27002 (N_27002,N_26905,N_26844);
nand U27003 (N_27003,N_26923,N_26697);
xor U27004 (N_27004,N_26717,N_26883);
nand U27005 (N_27005,N_26851,N_26679);
nand U27006 (N_27006,N_26744,N_26505);
and U27007 (N_27007,N_26913,N_26887);
and U27008 (N_27008,N_26530,N_26958);
nand U27009 (N_27009,N_26595,N_26807);
xor U27010 (N_27010,N_26523,N_26539);
xor U27011 (N_27011,N_26654,N_26788);
xor U27012 (N_27012,N_26650,N_26518);
nor U27013 (N_27013,N_26902,N_26980);
nor U27014 (N_27014,N_26576,N_26659);
nor U27015 (N_27015,N_26907,N_26532);
or U27016 (N_27016,N_26831,N_26708);
or U27017 (N_27017,N_26765,N_26737);
nand U27018 (N_27018,N_26810,N_26738);
and U27019 (N_27019,N_26845,N_26553);
or U27020 (N_27020,N_26676,N_26799);
and U27021 (N_27021,N_26824,N_26911);
nor U27022 (N_27022,N_26894,N_26632);
xnor U27023 (N_27023,N_26726,N_26941);
xnor U27024 (N_27024,N_26611,N_26803);
nor U27025 (N_27025,N_26688,N_26874);
nor U27026 (N_27026,N_26939,N_26790);
and U27027 (N_27027,N_26777,N_26964);
or U27028 (N_27028,N_26629,N_26792);
nand U27029 (N_27029,N_26932,N_26565);
or U27030 (N_27030,N_26860,N_26511);
and U27031 (N_27031,N_26948,N_26721);
nor U27032 (N_27032,N_26848,N_26525);
or U27033 (N_27033,N_26936,N_26873);
nand U27034 (N_27034,N_26747,N_26638);
or U27035 (N_27035,N_26605,N_26961);
and U27036 (N_27036,N_26730,N_26742);
nor U27037 (N_27037,N_26935,N_26898);
nand U27038 (N_27038,N_26671,N_26588);
nor U27039 (N_27039,N_26876,N_26604);
xnor U27040 (N_27040,N_26769,N_26597);
and U27041 (N_27041,N_26608,N_26857);
nand U27042 (N_27042,N_26534,N_26673);
nor U27043 (N_27043,N_26925,N_26984);
nor U27044 (N_27044,N_26563,N_26680);
and U27045 (N_27045,N_26692,N_26542);
nand U27046 (N_27046,N_26915,N_26975);
and U27047 (N_27047,N_26933,N_26972);
xor U27048 (N_27048,N_26985,N_26789);
xor U27049 (N_27049,N_26718,N_26685);
nor U27050 (N_27050,N_26806,N_26558);
and U27051 (N_27051,N_26893,N_26849);
and U27052 (N_27052,N_26979,N_26854);
nor U27053 (N_27053,N_26503,N_26639);
or U27054 (N_27054,N_26538,N_26551);
xnor U27055 (N_27055,N_26690,N_26924);
nor U27056 (N_27056,N_26987,N_26776);
nor U27057 (N_27057,N_26770,N_26818);
or U27058 (N_27058,N_26775,N_26591);
nor U27059 (N_27059,N_26645,N_26647);
and U27060 (N_27060,N_26513,N_26837);
and U27061 (N_27061,N_26703,N_26509);
xnor U27062 (N_27062,N_26561,N_26566);
nor U27063 (N_27063,N_26600,N_26570);
nand U27064 (N_27064,N_26559,N_26815);
and U27065 (N_27065,N_26937,N_26914);
nor U27066 (N_27066,N_26821,N_26660);
and U27067 (N_27067,N_26614,N_26990);
and U27068 (N_27068,N_26644,N_26892);
nand U27069 (N_27069,N_26843,N_26675);
nor U27070 (N_27070,N_26541,N_26749);
or U27071 (N_27071,N_26580,N_26965);
and U27072 (N_27072,N_26596,N_26699);
or U27073 (N_27073,N_26947,N_26683);
xor U27074 (N_27074,N_26574,N_26577);
nand U27075 (N_27075,N_26909,N_26521);
nor U27076 (N_27076,N_26888,N_26543);
or U27077 (N_27077,N_26636,N_26507);
nand U27078 (N_27078,N_26537,N_26739);
and U27079 (N_27079,N_26877,N_26613);
xor U27080 (N_27080,N_26899,N_26954);
nor U27081 (N_27081,N_26846,N_26656);
nand U27082 (N_27082,N_26830,N_26750);
or U27083 (N_27083,N_26871,N_26814);
or U27084 (N_27084,N_26993,N_26986);
and U27085 (N_27085,N_26601,N_26631);
nor U27086 (N_27086,N_26897,N_26522);
xnor U27087 (N_27087,N_26524,N_26896);
and U27088 (N_27088,N_26858,N_26784);
and U27089 (N_27089,N_26862,N_26519);
nand U27090 (N_27090,N_26828,N_26516);
and U27091 (N_27091,N_26571,N_26612);
nor U27092 (N_27092,N_26698,N_26569);
xnor U27093 (N_27093,N_26840,N_26763);
and U27094 (N_27094,N_26881,N_26994);
xor U27095 (N_27095,N_26794,N_26998);
xnor U27096 (N_27096,N_26796,N_26700);
xor U27097 (N_27097,N_26785,N_26733);
xnor U27098 (N_27098,N_26872,N_26757);
and U27099 (N_27099,N_26546,N_26836);
and U27100 (N_27100,N_26875,N_26921);
xnor U27101 (N_27101,N_26585,N_26533);
nor U27102 (N_27102,N_26504,N_26602);
nand U27103 (N_27103,N_26802,N_26847);
nor U27104 (N_27104,N_26768,N_26773);
and U27105 (N_27105,N_26946,N_26908);
xor U27106 (N_27106,N_26599,N_26878);
and U27107 (N_27107,N_26633,N_26672);
xnor U27108 (N_27108,N_26512,N_26865);
nand U27109 (N_27109,N_26758,N_26918);
nor U27110 (N_27110,N_26940,N_26801);
nor U27111 (N_27111,N_26514,N_26540);
or U27112 (N_27112,N_26573,N_26651);
nand U27113 (N_27113,N_26842,N_26771);
and U27114 (N_27114,N_26575,N_26767);
nor U27115 (N_27115,N_26832,N_26755);
xnor U27116 (N_27116,N_26916,N_26816);
nand U27117 (N_27117,N_26714,N_26822);
nand U27118 (N_27118,N_26678,N_26502);
nor U27119 (N_27119,N_26564,N_26957);
nor U27120 (N_27120,N_26732,N_26813);
nor U27121 (N_27121,N_26748,N_26616);
or U27122 (N_27122,N_26740,N_26618);
and U27123 (N_27123,N_26751,N_26741);
and U27124 (N_27124,N_26891,N_26760);
or U27125 (N_27125,N_26868,N_26833);
and U27126 (N_27126,N_26969,N_26953);
and U27127 (N_27127,N_26643,N_26900);
and U27128 (N_27128,N_26627,N_26625);
and U27129 (N_27129,N_26962,N_26804);
and U27130 (N_27130,N_26517,N_26641);
nand U27131 (N_27131,N_26753,N_26772);
nand U27132 (N_27132,N_26691,N_26510);
nand U27133 (N_27133,N_26646,N_26999);
nand U27134 (N_27134,N_26855,N_26945);
and U27135 (N_27135,N_26981,N_26684);
and U27136 (N_27136,N_26705,N_26779);
or U27137 (N_27137,N_26694,N_26995);
xnor U27138 (N_27138,N_26707,N_26562);
xnor U27139 (N_27139,N_26929,N_26853);
nor U27140 (N_27140,N_26736,N_26808);
or U27141 (N_27141,N_26992,N_26786);
xor U27142 (N_27142,N_26764,N_26841);
nand U27143 (N_27143,N_26715,N_26560);
nand U27144 (N_27144,N_26956,N_26904);
nand U27145 (N_27145,N_26971,N_26590);
and U27146 (N_27146,N_26531,N_26970);
xnor U27147 (N_27147,N_26890,N_26689);
and U27148 (N_27148,N_26508,N_26670);
nor U27149 (N_27149,N_26548,N_26637);
or U27150 (N_27150,N_26867,N_26687);
xnor U27151 (N_27151,N_26870,N_26834);
and U27152 (N_27152,N_26800,N_26966);
or U27153 (N_27153,N_26527,N_26586);
nor U27154 (N_27154,N_26906,N_26665);
or U27155 (N_27155,N_26667,N_26640);
and U27156 (N_27156,N_26850,N_26617);
nand U27157 (N_27157,N_26649,N_26944);
nor U27158 (N_27158,N_26549,N_26722);
xnor U27159 (N_27159,N_26712,N_26648);
nor U27160 (N_27160,N_26682,N_26653);
and U27161 (N_27161,N_26619,N_26988);
or U27162 (N_27162,N_26880,N_26528);
or U27163 (N_27163,N_26835,N_26989);
nor U27164 (N_27164,N_26955,N_26861);
nor U27165 (N_27165,N_26598,N_26793);
or U27166 (N_27166,N_26746,N_26693);
nor U27167 (N_27167,N_26978,N_26942);
xor U27168 (N_27168,N_26634,N_26663);
nor U27169 (N_27169,N_26568,N_26661);
or U27170 (N_27170,N_26716,N_26728);
nand U27171 (N_27171,N_26938,N_26968);
xor U27172 (N_27172,N_26886,N_26963);
and U27173 (N_27173,N_26838,N_26762);
or U27174 (N_27174,N_26960,N_26529);
and U27175 (N_27175,N_26997,N_26866);
and U27176 (N_27176,N_26535,N_26782);
nor U27177 (N_27177,N_26931,N_26754);
and U27178 (N_27178,N_26713,N_26555);
nor U27179 (N_27179,N_26879,N_26885);
nand U27180 (N_27180,N_26756,N_26526);
xnor U27181 (N_27181,N_26658,N_26922);
or U27182 (N_27182,N_26967,N_26895);
and U27183 (N_27183,N_26928,N_26727);
nand U27184 (N_27184,N_26554,N_26536);
xnor U27185 (N_27185,N_26859,N_26864);
xor U27186 (N_27186,N_26731,N_26583);
xnor U27187 (N_27187,N_26983,N_26884);
nor U27188 (N_27188,N_26766,N_26677);
xnor U27189 (N_27189,N_26706,N_26974);
xor U27190 (N_27190,N_26556,N_26823);
nand U27191 (N_27191,N_26603,N_26709);
or U27192 (N_27192,N_26926,N_26622);
or U27193 (N_27193,N_26630,N_26973);
xor U27194 (N_27194,N_26579,N_26696);
or U27195 (N_27195,N_26686,N_26809);
nand U27196 (N_27196,N_26547,N_26581);
and U27197 (N_27197,N_26780,N_26711);
nor U27198 (N_27198,N_26825,N_26917);
xnor U27199 (N_27199,N_26587,N_26774);
or U27200 (N_27200,N_26695,N_26819);
xor U27201 (N_27201,N_26919,N_26664);
or U27202 (N_27202,N_26621,N_26582);
or U27203 (N_27203,N_26805,N_26552);
and U27204 (N_27204,N_26704,N_26623);
xor U27205 (N_27205,N_26710,N_26642);
nand U27206 (N_27206,N_26949,N_26817);
xor U27207 (N_27207,N_26702,N_26544);
nand U27208 (N_27208,N_26798,N_26500);
or U27209 (N_27209,N_26593,N_26920);
or U27210 (N_27210,N_26669,N_26950);
or U27211 (N_27211,N_26934,N_26506);
nor U27212 (N_27212,N_26820,N_26930);
and U27213 (N_27213,N_26829,N_26620);
nand U27214 (N_27214,N_26951,N_26572);
or U27215 (N_27215,N_26787,N_26578);
xnor U27216 (N_27216,N_26882,N_26557);
xnor U27217 (N_27217,N_26889,N_26996);
and U27218 (N_27218,N_26584,N_26781);
nand U27219 (N_27219,N_26952,N_26912);
and U27220 (N_27220,N_26626,N_26545);
xnor U27221 (N_27221,N_26719,N_26725);
nor U27222 (N_27222,N_26592,N_26991);
and U27223 (N_27223,N_26515,N_26655);
nand U27224 (N_27224,N_26752,N_26657);
and U27225 (N_27225,N_26856,N_26701);
xnor U27226 (N_27226,N_26606,N_26743);
xnor U27227 (N_27227,N_26839,N_26735);
xnor U27228 (N_27228,N_26745,N_26927);
xor U27229 (N_27229,N_26795,N_26826);
or U27230 (N_27230,N_26827,N_26720);
xnor U27231 (N_27231,N_26982,N_26567);
nor U27232 (N_27232,N_26589,N_26783);
or U27233 (N_27233,N_26852,N_26734);
and U27234 (N_27234,N_26610,N_26501);
nor U27235 (N_27235,N_26609,N_26901);
nand U27236 (N_27236,N_26761,N_26666);
nor U27237 (N_27237,N_26724,N_26976);
nand U27238 (N_27238,N_26681,N_26778);
xor U27239 (N_27239,N_26520,N_26662);
nand U27240 (N_27240,N_26668,N_26811);
xnor U27241 (N_27241,N_26812,N_26977);
nand U27242 (N_27242,N_26869,N_26550);
nor U27243 (N_27243,N_26628,N_26759);
or U27244 (N_27244,N_26652,N_26729);
nor U27245 (N_27245,N_26910,N_26607);
nand U27246 (N_27246,N_26797,N_26903);
nor U27247 (N_27247,N_26624,N_26791);
or U27248 (N_27248,N_26959,N_26723);
nor U27249 (N_27249,N_26615,N_26594);
and U27250 (N_27250,N_26591,N_26531);
xor U27251 (N_27251,N_26771,N_26644);
nand U27252 (N_27252,N_26723,N_26729);
or U27253 (N_27253,N_26742,N_26560);
nor U27254 (N_27254,N_26501,N_26581);
nand U27255 (N_27255,N_26816,N_26699);
or U27256 (N_27256,N_26989,N_26943);
nand U27257 (N_27257,N_26749,N_26747);
nor U27258 (N_27258,N_26972,N_26960);
xor U27259 (N_27259,N_26925,N_26735);
or U27260 (N_27260,N_26629,N_26518);
xor U27261 (N_27261,N_26819,N_26903);
xnor U27262 (N_27262,N_26720,N_26973);
xnor U27263 (N_27263,N_26793,N_26735);
nand U27264 (N_27264,N_26917,N_26599);
or U27265 (N_27265,N_26580,N_26949);
or U27266 (N_27266,N_26527,N_26933);
nor U27267 (N_27267,N_26905,N_26522);
nand U27268 (N_27268,N_26881,N_26992);
nand U27269 (N_27269,N_26597,N_26617);
nand U27270 (N_27270,N_26598,N_26539);
or U27271 (N_27271,N_26718,N_26616);
nand U27272 (N_27272,N_26778,N_26535);
xnor U27273 (N_27273,N_26888,N_26995);
nand U27274 (N_27274,N_26956,N_26626);
nand U27275 (N_27275,N_26519,N_26857);
xor U27276 (N_27276,N_26819,N_26933);
or U27277 (N_27277,N_26781,N_26748);
or U27278 (N_27278,N_26844,N_26560);
nor U27279 (N_27279,N_26509,N_26877);
or U27280 (N_27280,N_26554,N_26815);
nand U27281 (N_27281,N_26585,N_26908);
xnor U27282 (N_27282,N_26722,N_26755);
or U27283 (N_27283,N_26549,N_26519);
and U27284 (N_27284,N_26931,N_26974);
or U27285 (N_27285,N_26798,N_26825);
and U27286 (N_27286,N_26594,N_26760);
or U27287 (N_27287,N_26540,N_26922);
nor U27288 (N_27288,N_26998,N_26587);
nor U27289 (N_27289,N_26674,N_26908);
or U27290 (N_27290,N_26747,N_26620);
nor U27291 (N_27291,N_26752,N_26709);
or U27292 (N_27292,N_26569,N_26868);
nand U27293 (N_27293,N_26648,N_26572);
nand U27294 (N_27294,N_26972,N_26921);
nor U27295 (N_27295,N_26523,N_26719);
nor U27296 (N_27296,N_26543,N_26937);
xnor U27297 (N_27297,N_26669,N_26943);
or U27298 (N_27298,N_26754,N_26845);
and U27299 (N_27299,N_26727,N_26807);
or U27300 (N_27300,N_26837,N_26901);
and U27301 (N_27301,N_26828,N_26717);
and U27302 (N_27302,N_26932,N_26645);
or U27303 (N_27303,N_26507,N_26625);
or U27304 (N_27304,N_26877,N_26503);
nor U27305 (N_27305,N_26598,N_26666);
nand U27306 (N_27306,N_26910,N_26900);
nand U27307 (N_27307,N_26935,N_26983);
nor U27308 (N_27308,N_26500,N_26826);
nor U27309 (N_27309,N_26517,N_26610);
xnor U27310 (N_27310,N_26513,N_26526);
and U27311 (N_27311,N_26809,N_26530);
xnor U27312 (N_27312,N_26834,N_26908);
or U27313 (N_27313,N_26895,N_26622);
nor U27314 (N_27314,N_26614,N_26660);
nor U27315 (N_27315,N_26537,N_26982);
or U27316 (N_27316,N_26856,N_26917);
and U27317 (N_27317,N_26584,N_26809);
nand U27318 (N_27318,N_26712,N_26582);
xor U27319 (N_27319,N_26625,N_26701);
nor U27320 (N_27320,N_26924,N_26825);
xor U27321 (N_27321,N_26540,N_26784);
and U27322 (N_27322,N_26528,N_26725);
and U27323 (N_27323,N_26596,N_26756);
or U27324 (N_27324,N_26811,N_26756);
and U27325 (N_27325,N_26761,N_26791);
xor U27326 (N_27326,N_26940,N_26904);
nand U27327 (N_27327,N_26889,N_26852);
nand U27328 (N_27328,N_26981,N_26616);
xnor U27329 (N_27329,N_26864,N_26973);
nor U27330 (N_27330,N_26524,N_26969);
xnor U27331 (N_27331,N_26611,N_26628);
nand U27332 (N_27332,N_26631,N_26521);
or U27333 (N_27333,N_26617,N_26977);
and U27334 (N_27334,N_26737,N_26788);
nor U27335 (N_27335,N_26672,N_26596);
nor U27336 (N_27336,N_26566,N_26901);
and U27337 (N_27337,N_26824,N_26701);
and U27338 (N_27338,N_26779,N_26893);
or U27339 (N_27339,N_26743,N_26894);
or U27340 (N_27340,N_26583,N_26904);
nor U27341 (N_27341,N_26679,N_26888);
xor U27342 (N_27342,N_26569,N_26500);
nor U27343 (N_27343,N_26522,N_26647);
nor U27344 (N_27344,N_26505,N_26686);
or U27345 (N_27345,N_26984,N_26713);
xor U27346 (N_27346,N_26996,N_26972);
nor U27347 (N_27347,N_26592,N_26681);
nor U27348 (N_27348,N_26957,N_26811);
nand U27349 (N_27349,N_26557,N_26591);
xnor U27350 (N_27350,N_26516,N_26648);
and U27351 (N_27351,N_26915,N_26764);
or U27352 (N_27352,N_26887,N_26642);
xnor U27353 (N_27353,N_26862,N_26863);
and U27354 (N_27354,N_26960,N_26628);
nor U27355 (N_27355,N_26568,N_26840);
and U27356 (N_27356,N_26931,N_26753);
and U27357 (N_27357,N_26665,N_26578);
and U27358 (N_27358,N_26805,N_26862);
or U27359 (N_27359,N_26635,N_26810);
nand U27360 (N_27360,N_26568,N_26554);
xnor U27361 (N_27361,N_26699,N_26750);
xor U27362 (N_27362,N_26632,N_26858);
nand U27363 (N_27363,N_26811,N_26582);
and U27364 (N_27364,N_26822,N_26562);
or U27365 (N_27365,N_26697,N_26794);
xnor U27366 (N_27366,N_26988,N_26742);
nor U27367 (N_27367,N_26695,N_26859);
nand U27368 (N_27368,N_26978,N_26506);
and U27369 (N_27369,N_26955,N_26676);
or U27370 (N_27370,N_26757,N_26639);
and U27371 (N_27371,N_26738,N_26965);
nor U27372 (N_27372,N_26873,N_26892);
nor U27373 (N_27373,N_26748,N_26903);
or U27374 (N_27374,N_26676,N_26800);
nor U27375 (N_27375,N_26565,N_26574);
or U27376 (N_27376,N_26833,N_26661);
nand U27377 (N_27377,N_26625,N_26947);
and U27378 (N_27378,N_26868,N_26877);
nor U27379 (N_27379,N_26818,N_26703);
nor U27380 (N_27380,N_26833,N_26866);
nand U27381 (N_27381,N_26562,N_26754);
or U27382 (N_27382,N_26702,N_26815);
and U27383 (N_27383,N_26929,N_26802);
xnor U27384 (N_27384,N_26858,N_26697);
or U27385 (N_27385,N_26648,N_26753);
nand U27386 (N_27386,N_26737,N_26570);
nand U27387 (N_27387,N_26794,N_26986);
nand U27388 (N_27388,N_26828,N_26623);
nand U27389 (N_27389,N_26793,N_26951);
or U27390 (N_27390,N_26932,N_26703);
or U27391 (N_27391,N_26867,N_26724);
nor U27392 (N_27392,N_26511,N_26948);
or U27393 (N_27393,N_26643,N_26667);
and U27394 (N_27394,N_26763,N_26912);
or U27395 (N_27395,N_26898,N_26930);
or U27396 (N_27396,N_26818,N_26702);
nand U27397 (N_27397,N_26625,N_26651);
or U27398 (N_27398,N_26723,N_26754);
xor U27399 (N_27399,N_26804,N_26749);
xor U27400 (N_27400,N_26558,N_26875);
nor U27401 (N_27401,N_26879,N_26938);
and U27402 (N_27402,N_26732,N_26787);
nand U27403 (N_27403,N_26708,N_26844);
nor U27404 (N_27404,N_26642,N_26560);
nand U27405 (N_27405,N_26611,N_26849);
or U27406 (N_27406,N_26589,N_26684);
nand U27407 (N_27407,N_26501,N_26529);
or U27408 (N_27408,N_26702,N_26725);
nor U27409 (N_27409,N_26957,N_26602);
xor U27410 (N_27410,N_26549,N_26643);
xor U27411 (N_27411,N_26706,N_26728);
or U27412 (N_27412,N_26764,N_26799);
xnor U27413 (N_27413,N_26581,N_26871);
nand U27414 (N_27414,N_26735,N_26804);
nor U27415 (N_27415,N_26842,N_26815);
nor U27416 (N_27416,N_26959,N_26870);
and U27417 (N_27417,N_26706,N_26698);
xor U27418 (N_27418,N_26952,N_26537);
nand U27419 (N_27419,N_26988,N_26796);
or U27420 (N_27420,N_26898,N_26957);
or U27421 (N_27421,N_26820,N_26931);
or U27422 (N_27422,N_26899,N_26892);
nor U27423 (N_27423,N_26953,N_26899);
and U27424 (N_27424,N_26768,N_26980);
or U27425 (N_27425,N_26850,N_26687);
xnor U27426 (N_27426,N_26727,N_26840);
nand U27427 (N_27427,N_26763,N_26974);
nor U27428 (N_27428,N_26695,N_26861);
or U27429 (N_27429,N_26647,N_26609);
nand U27430 (N_27430,N_26607,N_26980);
and U27431 (N_27431,N_26765,N_26575);
nand U27432 (N_27432,N_26547,N_26531);
and U27433 (N_27433,N_26524,N_26604);
or U27434 (N_27434,N_26613,N_26879);
nor U27435 (N_27435,N_26697,N_26811);
or U27436 (N_27436,N_26639,N_26505);
and U27437 (N_27437,N_26700,N_26666);
xor U27438 (N_27438,N_26909,N_26686);
or U27439 (N_27439,N_26770,N_26862);
or U27440 (N_27440,N_26632,N_26898);
nor U27441 (N_27441,N_26668,N_26998);
or U27442 (N_27442,N_26693,N_26793);
or U27443 (N_27443,N_26855,N_26829);
or U27444 (N_27444,N_26621,N_26727);
xor U27445 (N_27445,N_26962,N_26932);
or U27446 (N_27446,N_26753,N_26715);
nor U27447 (N_27447,N_26543,N_26929);
or U27448 (N_27448,N_26840,N_26684);
or U27449 (N_27449,N_26661,N_26717);
nand U27450 (N_27450,N_26973,N_26763);
and U27451 (N_27451,N_26621,N_26919);
nand U27452 (N_27452,N_26767,N_26646);
or U27453 (N_27453,N_26988,N_26816);
nor U27454 (N_27454,N_26718,N_26762);
xnor U27455 (N_27455,N_26949,N_26894);
xnor U27456 (N_27456,N_26828,N_26990);
nor U27457 (N_27457,N_26690,N_26573);
nor U27458 (N_27458,N_26664,N_26571);
nand U27459 (N_27459,N_26522,N_26569);
and U27460 (N_27460,N_26583,N_26704);
nor U27461 (N_27461,N_26758,N_26792);
nand U27462 (N_27462,N_26751,N_26820);
and U27463 (N_27463,N_26963,N_26717);
or U27464 (N_27464,N_26966,N_26863);
nand U27465 (N_27465,N_26838,N_26678);
nand U27466 (N_27466,N_26833,N_26916);
nor U27467 (N_27467,N_26515,N_26844);
nor U27468 (N_27468,N_26604,N_26504);
or U27469 (N_27469,N_26974,N_26958);
xnor U27470 (N_27470,N_26940,N_26670);
or U27471 (N_27471,N_26640,N_26930);
nor U27472 (N_27472,N_26692,N_26501);
xnor U27473 (N_27473,N_26601,N_26597);
or U27474 (N_27474,N_26644,N_26987);
xor U27475 (N_27475,N_26679,N_26683);
and U27476 (N_27476,N_26740,N_26718);
nor U27477 (N_27477,N_26601,N_26664);
nor U27478 (N_27478,N_26718,N_26934);
nor U27479 (N_27479,N_26688,N_26681);
or U27480 (N_27480,N_26709,N_26813);
nor U27481 (N_27481,N_26607,N_26888);
xnor U27482 (N_27482,N_26765,N_26983);
nand U27483 (N_27483,N_26661,N_26918);
nand U27484 (N_27484,N_26763,N_26911);
and U27485 (N_27485,N_26849,N_26847);
and U27486 (N_27486,N_26812,N_26983);
and U27487 (N_27487,N_26722,N_26821);
nand U27488 (N_27488,N_26748,N_26669);
and U27489 (N_27489,N_26817,N_26614);
and U27490 (N_27490,N_26880,N_26914);
nor U27491 (N_27491,N_26740,N_26885);
xnor U27492 (N_27492,N_26710,N_26811);
and U27493 (N_27493,N_26995,N_26873);
or U27494 (N_27494,N_26649,N_26777);
xnor U27495 (N_27495,N_26780,N_26879);
or U27496 (N_27496,N_26931,N_26575);
or U27497 (N_27497,N_26572,N_26956);
nand U27498 (N_27498,N_26940,N_26851);
and U27499 (N_27499,N_26904,N_26546);
nand U27500 (N_27500,N_27411,N_27105);
nand U27501 (N_27501,N_27498,N_27388);
nor U27502 (N_27502,N_27390,N_27454);
or U27503 (N_27503,N_27288,N_27141);
nand U27504 (N_27504,N_27004,N_27151);
nand U27505 (N_27505,N_27296,N_27363);
nor U27506 (N_27506,N_27494,N_27387);
or U27507 (N_27507,N_27372,N_27050);
or U27508 (N_27508,N_27384,N_27403);
and U27509 (N_27509,N_27030,N_27070);
xnor U27510 (N_27510,N_27394,N_27412);
xnor U27511 (N_27511,N_27098,N_27063);
nand U27512 (N_27512,N_27162,N_27110);
nor U27513 (N_27513,N_27154,N_27276);
and U27514 (N_27514,N_27464,N_27005);
or U27515 (N_27515,N_27116,N_27294);
and U27516 (N_27516,N_27081,N_27264);
nand U27517 (N_27517,N_27324,N_27139);
nor U27518 (N_27518,N_27121,N_27487);
nand U27519 (N_27519,N_27295,N_27468);
nand U27520 (N_27520,N_27182,N_27416);
nor U27521 (N_27521,N_27404,N_27446);
nor U27522 (N_27522,N_27447,N_27356);
or U27523 (N_27523,N_27473,N_27061);
or U27524 (N_27524,N_27006,N_27339);
and U27525 (N_27525,N_27366,N_27273);
and U27526 (N_27526,N_27223,N_27313);
or U27527 (N_27527,N_27332,N_27108);
nor U27528 (N_27528,N_27365,N_27436);
or U27529 (N_27529,N_27328,N_27274);
or U27530 (N_27530,N_27218,N_27430);
and U27531 (N_27531,N_27143,N_27052);
nor U27532 (N_27532,N_27173,N_27008);
nor U27533 (N_27533,N_27307,N_27248);
and U27534 (N_27534,N_27206,N_27208);
nand U27535 (N_27535,N_27391,N_27376);
nand U27536 (N_27536,N_27240,N_27038);
xnor U27537 (N_27537,N_27286,N_27393);
xor U27538 (N_27538,N_27083,N_27217);
or U27539 (N_27539,N_27456,N_27419);
xor U27540 (N_27540,N_27175,N_27291);
or U27541 (N_27541,N_27170,N_27268);
xnor U27542 (N_27542,N_27104,N_27449);
nor U27543 (N_27543,N_27389,N_27046);
or U27544 (N_27544,N_27212,N_27250);
nand U27545 (N_27545,N_27335,N_27491);
nand U27546 (N_27546,N_27392,N_27087);
xnor U27547 (N_27547,N_27343,N_27044);
nand U27548 (N_27548,N_27001,N_27458);
and U27549 (N_27549,N_27331,N_27074);
nor U27550 (N_27550,N_27041,N_27476);
nor U27551 (N_27551,N_27091,N_27169);
xnor U27552 (N_27552,N_27334,N_27309);
nand U27553 (N_27553,N_27347,N_27472);
nor U27554 (N_27554,N_27002,N_27140);
and U27555 (N_27555,N_27025,N_27158);
and U27556 (N_27556,N_27287,N_27266);
nand U27557 (N_27557,N_27204,N_27306);
or U27558 (N_27558,N_27055,N_27234);
nand U27559 (N_27559,N_27378,N_27144);
nand U27560 (N_27560,N_27118,N_27186);
nand U27561 (N_27561,N_27357,N_27016);
nor U27562 (N_27562,N_27191,N_27370);
nor U27563 (N_27563,N_27202,N_27097);
nor U27564 (N_27564,N_27245,N_27455);
nand U27565 (N_27565,N_27433,N_27445);
xor U27566 (N_27566,N_27318,N_27230);
xnor U27567 (N_27567,N_27185,N_27374);
or U27568 (N_27568,N_27236,N_27222);
nor U27569 (N_27569,N_27113,N_27226);
nor U27570 (N_27570,N_27159,N_27323);
and U27571 (N_27571,N_27137,N_27262);
nor U27572 (N_27572,N_27178,N_27009);
nand U27573 (N_27573,N_27338,N_27232);
nor U27574 (N_27574,N_27478,N_27341);
and U27575 (N_27575,N_27282,N_27233);
and U27576 (N_27576,N_27377,N_27126);
nand U27577 (N_27577,N_27480,N_27012);
xor U27578 (N_27578,N_27125,N_27174);
xnor U27579 (N_27579,N_27089,N_27424);
nor U27580 (N_27580,N_27056,N_27414);
or U27581 (N_27581,N_27285,N_27020);
or U27582 (N_27582,N_27350,N_27453);
xor U27583 (N_27583,N_27405,N_27441);
xor U27584 (N_27584,N_27219,N_27256);
nand U27585 (N_27585,N_27147,N_27239);
nor U27586 (N_27586,N_27259,N_27326);
or U27587 (N_27587,N_27119,N_27431);
nor U27588 (N_27588,N_27459,N_27167);
or U27589 (N_27589,N_27361,N_27073);
or U27590 (N_27590,N_27205,N_27267);
xnor U27591 (N_27591,N_27157,N_27200);
or U27592 (N_27592,N_27255,N_27210);
or U27593 (N_27593,N_27272,N_27235);
nand U27594 (N_27594,N_27409,N_27043);
and U27595 (N_27595,N_27499,N_27152);
and U27596 (N_27596,N_27401,N_27013);
xnor U27597 (N_27597,N_27060,N_27465);
nor U27598 (N_27598,N_27317,N_27461);
or U27599 (N_27599,N_27132,N_27066);
nand U27600 (N_27600,N_27321,N_27155);
nand U27601 (N_27601,N_27349,N_27402);
nor U27602 (N_27602,N_27467,N_27029);
or U27603 (N_27603,N_27076,N_27329);
or U27604 (N_27604,N_27194,N_27034);
xor U27605 (N_27605,N_27327,N_27065);
nor U27606 (N_27606,N_27156,N_27463);
or U27607 (N_27607,N_27054,N_27400);
or U27608 (N_27608,N_27049,N_27123);
nor U27609 (N_27609,N_27423,N_27497);
or U27610 (N_27610,N_27303,N_27386);
nor U27611 (N_27611,N_27358,N_27367);
nand U27612 (N_27612,N_27224,N_27131);
and U27613 (N_27613,N_27422,N_27261);
xor U27614 (N_27614,N_27308,N_27011);
or U27615 (N_27615,N_27086,N_27310);
nand U27616 (N_27616,N_27354,N_27135);
nor U27617 (N_27617,N_27216,N_27382);
nand U27618 (N_27618,N_27022,N_27271);
xnor U27619 (N_27619,N_27032,N_27260);
xnor U27620 (N_27620,N_27100,N_27263);
nor U27621 (N_27621,N_27277,N_27062);
xnor U27622 (N_27622,N_27289,N_27359);
nor U27623 (N_27623,N_27352,N_27312);
and U27624 (N_27624,N_27353,N_27369);
nand U27625 (N_27625,N_27251,N_27021);
and U27626 (N_27626,N_27413,N_27036);
and U27627 (N_27627,N_27068,N_27007);
nand U27628 (N_27628,N_27242,N_27039);
and U27629 (N_27629,N_27283,N_27057);
or U27630 (N_27630,N_27381,N_27138);
and U27631 (N_27631,N_27399,N_27371);
nand U27632 (N_27632,N_27122,N_27124);
xnor U27633 (N_27633,N_27026,N_27168);
nor U27634 (N_27634,N_27019,N_27172);
or U27635 (N_27635,N_27214,N_27102);
or U27636 (N_27636,N_27010,N_27003);
nor U27637 (N_27637,N_27238,N_27257);
xor U27638 (N_27638,N_27336,N_27373);
nor U27639 (N_27639,N_27096,N_27483);
nand U27640 (N_27640,N_27069,N_27333);
or U27641 (N_27641,N_27345,N_27448);
nor U27642 (N_27642,N_27080,N_27213);
and U27643 (N_27643,N_27435,N_27298);
nor U27644 (N_27644,N_27474,N_27244);
nand U27645 (N_27645,N_27439,N_27183);
xor U27646 (N_27646,N_27485,N_27095);
and U27647 (N_27647,N_27093,N_27227);
nor U27648 (N_27648,N_27410,N_27396);
nand U27649 (N_27649,N_27330,N_27107);
or U27650 (N_27650,N_27475,N_27184);
and U27651 (N_27651,N_27228,N_27053);
nand U27652 (N_27652,N_27397,N_27383);
nand U27653 (N_27653,N_27017,N_27425);
or U27654 (N_27654,N_27215,N_27444);
and U27655 (N_27655,N_27302,N_27127);
and U27656 (N_27656,N_27292,N_27112);
nand U27657 (N_27657,N_27406,N_27203);
or U27658 (N_27658,N_27099,N_27495);
nor U27659 (N_27659,N_27418,N_27201);
nor U27660 (N_27660,N_27482,N_27024);
or U27661 (N_27661,N_27432,N_27375);
xnor U27662 (N_27662,N_27166,N_27299);
xnor U27663 (N_27663,N_27164,N_27270);
nand U27664 (N_27664,N_27477,N_27058);
xor U27665 (N_27665,N_27496,N_27189);
and U27666 (N_27666,N_27115,N_27114);
and U27667 (N_27667,N_27325,N_27379);
xnor U27668 (N_27668,N_27160,N_27254);
nand U27669 (N_27669,N_27018,N_27322);
nor U27670 (N_27670,N_27265,N_27094);
nor U27671 (N_27671,N_27171,N_27428);
or U27672 (N_27672,N_27180,N_27243);
nor U27673 (N_27673,N_27072,N_27059);
and U27674 (N_27674,N_27198,N_27351);
nor U27675 (N_27675,N_27035,N_27045);
xnor U27676 (N_27676,N_27101,N_27320);
nor U27677 (N_27677,N_27117,N_27280);
or U27678 (N_27678,N_27197,N_27153);
xnor U27679 (N_27679,N_27490,N_27000);
nor U27680 (N_27680,N_27067,N_27301);
and U27681 (N_27681,N_27231,N_27304);
and U27682 (N_27682,N_27207,N_27048);
nand U27683 (N_27683,N_27315,N_27417);
nand U27684 (N_27684,N_27103,N_27460);
and U27685 (N_27685,N_27293,N_27090);
nand U27686 (N_27686,N_27407,N_27305);
or U27687 (N_27687,N_27470,N_27128);
nor U27688 (N_27688,N_27380,N_27027);
or U27689 (N_27689,N_27130,N_27042);
xnor U27690 (N_27690,N_27385,N_27492);
and U27691 (N_27691,N_27368,N_27275);
or U27692 (N_27692,N_27015,N_27109);
xnor U27693 (N_27693,N_27149,N_27420);
or U27694 (N_27694,N_27342,N_27486);
and U27695 (N_27695,N_27258,N_27075);
nor U27696 (N_27696,N_27340,N_27176);
nor U27697 (N_27697,N_27192,N_27241);
and U27698 (N_27698,N_27079,N_27181);
nor U27699 (N_27699,N_27484,N_27493);
nor U27700 (N_27700,N_27085,N_27023);
nor U27701 (N_27701,N_27082,N_27193);
and U27702 (N_27702,N_27279,N_27408);
xor U27703 (N_27703,N_27092,N_27427);
nand U27704 (N_27704,N_27078,N_27165);
or U27705 (N_27705,N_27064,N_27148);
nand U27706 (N_27706,N_27281,N_27033);
nor U27707 (N_27707,N_27440,N_27084);
nor U27708 (N_27708,N_27037,N_27415);
or U27709 (N_27709,N_27220,N_27188);
nand U27710 (N_27710,N_27450,N_27290);
xor U27711 (N_27711,N_27297,N_27129);
or U27712 (N_27712,N_27161,N_27047);
or U27713 (N_27713,N_27300,N_27150);
nand U27714 (N_27714,N_27195,N_27031);
nand U27715 (N_27715,N_27284,N_27246);
xor U27716 (N_27716,N_27247,N_27221);
and U27717 (N_27717,N_27489,N_27209);
and U27718 (N_27718,N_27443,N_27360);
nor U27719 (N_27719,N_27364,N_27398);
or U27720 (N_27720,N_27196,N_27142);
xor U27721 (N_27721,N_27316,N_27229);
or U27722 (N_27722,N_27253,N_27190);
and U27723 (N_27723,N_27311,N_27438);
nand U27724 (N_27724,N_27362,N_27469);
and U27725 (N_27725,N_27136,N_27337);
nor U27726 (N_27726,N_27479,N_27051);
and U27727 (N_27727,N_27348,N_27481);
xor U27728 (N_27728,N_27225,N_27355);
or U27729 (N_27729,N_27421,N_27462);
xnor U27730 (N_27730,N_27466,N_27249);
xor U27731 (N_27731,N_27040,N_27120);
or U27732 (N_27732,N_27395,N_27426);
xnor U27733 (N_27733,N_27134,N_27451);
nor U27734 (N_27734,N_27088,N_27014);
nor U27735 (N_27735,N_27346,N_27028);
or U27736 (N_27736,N_27199,N_27442);
xor U27737 (N_27737,N_27278,N_27488);
nor U27738 (N_27738,N_27434,N_27187);
and U27739 (N_27739,N_27429,N_27252);
or U27740 (N_27740,N_27344,N_27177);
xor U27741 (N_27741,N_27452,N_27146);
nor U27742 (N_27742,N_27163,N_27269);
or U27743 (N_27743,N_27314,N_27133);
and U27744 (N_27744,N_27179,N_27437);
and U27745 (N_27745,N_27106,N_27211);
and U27746 (N_27746,N_27145,N_27319);
nand U27747 (N_27747,N_27071,N_27111);
nand U27748 (N_27748,N_27471,N_27077);
and U27749 (N_27749,N_27237,N_27457);
or U27750 (N_27750,N_27382,N_27297);
and U27751 (N_27751,N_27289,N_27373);
and U27752 (N_27752,N_27447,N_27027);
and U27753 (N_27753,N_27152,N_27275);
and U27754 (N_27754,N_27002,N_27291);
xor U27755 (N_27755,N_27288,N_27053);
nor U27756 (N_27756,N_27316,N_27490);
xnor U27757 (N_27757,N_27474,N_27269);
xor U27758 (N_27758,N_27134,N_27300);
and U27759 (N_27759,N_27463,N_27138);
nor U27760 (N_27760,N_27094,N_27070);
or U27761 (N_27761,N_27372,N_27235);
or U27762 (N_27762,N_27330,N_27129);
and U27763 (N_27763,N_27446,N_27478);
nor U27764 (N_27764,N_27340,N_27475);
nand U27765 (N_27765,N_27190,N_27252);
xor U27766 (N_27766,N_27058,N_27414);
or U27767 (N_27767,N_27137,N_27219);
or U27768 (N_27768,N_27441,N_27128);
xor U27769 (N_27769,N_27326,N_27363);
nor U27770 (N_27770,N_27456,N_27111);
and U27771 (N_27771,N_27235,N_27331);
or U27772 (N_27772,N_27234,N_27372);
nand U27773 (N_27773,N_27163,N_27015);
nand U27774 (N_27774,N_27227,N_27372);
nor U27775 (N_27775,N_27001,N_27335);
xnor U27776 (N_27776,N_27113,N_27172);
nor U27777 (N_27777,N_27097,N_27451);
and U27778 (N_27778,N_27164,N_27066);
xnor U27779 (N_27779,N_27201,N_27056);
nand U27780 (N_27780,N_27391,N_27400);
nor U27781 (N_27781,N_27391,N_27493);
nand U27782 (N_27782,N_27066,N_27338);
xor U27783 (N_27783,N_27213,N_27196);
and U27784 (N_27784,N_27441,N_27214);
or U27785 (N_27785,N_27261,N_27170);
nor U27786 (N_27786,N_27211,N_27409);
nand U27787 (N_27787,N_27090,N_27487);
nand U27788 (N_27788,N_27300,N_27318);
nor U27789 (N_27789,N_27360,N_27440);
nand U27790 (N_27790,N_27379,N_27465);
or U27791 (N_27791,N_27437,N_27077);
and U27792 (N_27792,N_27430,N_27120);
nand U27793 (N_27793,N_27377,N_27343);
xor U27794 (N_27794,N_27224,N_27197);
nand U27795 (N_27795,N_27486,N_27282);
and U27796 (N_27796,N_27322,N_27338);
or U27797 (N_27797,N_27380,N_27330);
and U27798 (N_27798,N_27447,N_27380);
and U27799 (N_27799,N_27241,N_27218);
or U27800 (N_27800,N_27338,N_27173);
nand U27801 (N_27801,N_27066,N_27385);
nor U27802 (N_27802,N_27105,N_27342);
and U27803 (N_27803,N_27165,N_27262);
nand U27804 (N_27804,N_27118,N_27352);
and U27805 (N_27805,N_27305,N_27278);
nand U27806 (N_27806,N_27350,N_27136);
nand U27807 (N_27807,N_27141,N_27216);
or U27808 (N_27808,N_27478,N_27227);
and U27809 (N_27809,N_27285,N_27337);
nor U27810 (N_27810,N_27409,N_27184);
nor U27811 (N_27811,N_27470,N_27377);
and U27812 (N_27812,N_27416,N_27137);
nor U27813 (N_27813,N_27134,N_27349);
or U27814 (N_27814,N_27177,N_27237);
nand U27815 (N_27815,N_27451,N_27237);
nor U27816 (N_27816,N_27354,N_27104);
and U27817 (N_27817,N_27175,N_27296);
xor U27818 (N_27818,N_27122,N_27019);
and U27819 (N_27819,N_27325,N_27172);
or U27820 (N_27820,N_27351,N_27292);
xnor U27821 (N_27821,N_27425,N_27300);
xor U27822 (N_27822,N_27413,N_27063);
xor U27823 (N_27823,N_27261,N_27443);
nand U27824 (N_27824,N_27289,N_27175);
nor U27825 (N_27825,N_27006,N_27054);
and U27826 (N_27826,N_27442,N_27390);
nor U27827 (N_27827,N_27228,N_27240);
and U27828 (N_27828,N_27385,N_27125);
or U27829 (N_27829,N_27044,N_27484);
and U27830 (N_27830,N_27446,N_27079);
nor U27831 (N_27831,N_27446,N_27106);
xnor U27832 (N_27832,N_27290,N_27057);
nor U27833 (N_27833,N_27182,N_27407);
or U27834 (N_27834,N_27210,N_27027);
nor U27835 (N_27835,N_27494,N_27025);
xor U27836 (N_27836,N_27030,N_27114);
nand U27837 (N_27837,N_27260,N_27248);
nor U27838 (N_27838,N_27438,N_27424);
or U27839 (N_27839,N_27439,N_27374);
and U27840 (N_27840,N_27030,N_27251);
xnor U27841 (N_27841,N_27097,N_27356);
nor U27842 (N_27842,N_27269,N_27305);
nand U27843 (N_27843,N_27487,N_27489);
nor U27844 (N_27844,N_27000,N_27335);
xnor U27845 (N_27845,N_27180,N_27352);
nor U27846 (N_27846,N_27126,N_27223);
xnor U27847 (N_27847,N_27362,N_27081);
xor U27848 (N_27848,N_27035,N_27485);
xnor U27849 (N_27849,N_27062,N_27403);
and U27850 (N_27850,N_27415,N_27090);
xor U27851 (N_27851,N_27057,N_27314);
or U27852 (N_27852,N_27323,N_27199);
nand U27853 (N_27853,N_27121,N_27101);
and U27854 (N_27854,N_27034,N_27339);
nor U27855 (N_27855,N_27108,N_27313);
xnor U27856 (N_27856,N_27111,N_27004);
and U27857 (N_27857,N_27466,N_27204);
or U27858 (N_27858,N_27391,N_27377);
and U27859 (N_27859,N_27282,N_27241);
xnor U27860 (N_27860,N_27301,N_27382);
nor U27861 (N_27861,N_27007,N_27101);
nor U27862 (N_27862,N_27358,N_27488);
xor U27863 (N_27863,N_27031,N_27053);
xor U27864 (N_27864,N_27453,N_27388);
nand U27865 (N_27865,N_27177,N_27076);
nand U27866 (N_27866,N_27317,N_27389);
and U27867 (N_27867,N_27112,N_27066);
and U27868 (N_27868,N_27038,N_27291);
nand U27869 (N_27869,N_27326,N_27064);
and U27870 (N_27870,N_27159,N_27032);
xor U27871 (N_27871,N_27128,N_27453);
xor U27872 (N_27872,N_27410,N_27156);
and U27873 (N_27873,N_27347,N_27235);
and U27874 (N_27874,N_27224,N_27273);
xnor U27875 (N_27875,N_27464,N_27447);
xnor U27876 (N_27876,N_27409,N_27173);
or U27877 (N_27877,N_27457,N_27138);
and U27878 (N_27878,N_27152,N_27061);
nand U27879 (N_27879,N_27425,N_27103);
and U27880 (N_27880,N_27077,N_27478);
or U27881 (N_27881,N_27151,N_27044);
and U27882 (N_27882,N_27022,N_27077);
or U27883 (N_27883,N_27429,N_27446);
nand U27884 (N_27884,N_27084,N_27002);
nand U27885 (N_27885,N_27147,N_27461);
nor U27886 (N_27886,N_27005,N_27010);
xor U27887 (N_27887,N_27408,N_27340);
or U27888 (N_27888,N_27217,N_27004);
nand U27889 (N_27889,N_27074,N_27391);
and U27890 (N_27890,N_27167,N_27126);
nand U27891 (N_27891,N_27164,N_27144);
and U27892 (N_27892,N_27029,N_27436);
nor U27893 (N_27893,N_27033,N_27340);
nand U27894 (N_27894,N_27053,N_27369);
nor U27895 (N_27895,N_27425,N_27167);
or U27896 (N_27896,N_27303,N_27302);
nand U27897 (N_27897,N_27149,N_27165);
or U27898 (N_27898,N_27440,N_27192);
nand U27899 (N_27899,N_27074,N_27055);
or U27900 (N_27900,N_27033,N_27497);
nand U27901 (N_27901,N_27147,N_27039);
and U27902 (N_27902,N_27119,N_27301);
or U27903 (N_27903,N_27442,N_27065);
nand U27904 (N_27904,N_27344,N_27397);
or U27905 (N_27905,N_27163,N_27477);
nor U27906 (N_27906,N_27207,N_27135);
nand U27907 (N_27907,N_27239,N_27097);
or U27908 (N_27908,N_27027,N_27111);
xor U27909 (N_27909,N_27261,N_27412);
nand U27910 (N_27910,N_27068,N_27398);
nor U27911 (N_27911,N_27030,N_27147);
xor U27912 (N_27912,N_27361,N_27227);
nor U27913 (N_27913,N_27412,N_27176);
or U27914 (N_27914,N_27491,N_27259);
xor U27915 (N_27915,N_27060,N_27342);
nor U27916 (N_27916,N_27208,N_27044);
or U27917 (N_27917,N_27281,N_27474);
nand U27918 (N_27918,N_27320,N_27295);
or U27919 (N_27919,N_27383,N_27412);
xnor U27920 (N_27920,N_27390,N_27489);
and U27921 (N_27921,N_27189,N_27216);
and U27922 (N_27922,N_27232,N_27079);
xor U27923 (N_27923,N_27234,N_27162);
or U27924 (N_27924,N_27164,N_27425);
and U27925 (N_27925,N_27272,N_27336);
xor U27926 (N_27926,N_27309,N_27269);
nor U27927 (N_27927,N_27410,N_27306);
xnor U27928 (N_27928,N_27246,N_27343);
nor U27929 (N_27929,N_27476,N_27046);
xnor U27930 (N_27930,N_27365,N_27421);
nor U27931 (N_27931,N_27487,N_27195);
nand U27932 (N_27932,N_27429,N_27389);
and U27933 (N_27933,N_27358,N_27034);
xnor U27934 (N_27934,N_27448,N_27304);
or U27935 (N_27935,N_27147,N_27054);
or U27936 (N_27936,N_27239,N_27000);
xor U27937 (N_27937,N_27059,N_27064);
xor U27938 (N_27938,N_27397,N_27445);
or U27939 (N_27939,N_27205,N_27031);
and U27940 (N_27940,N_27435,N_27471);
xnor U27941 (N_27941,N_27365,N_27134);
and U27942 (N_27942,N_27101,N_27127);
or U27943 (N_27943,N_27068,N_27492);
and U27944 (N_27944,N_27261,N_27265);
nor U27945 (N_27945,N_27393,N_27241);
xor U27946 (N_27946,N_27199,N_27131);
and U27947 (N_27947,N_27393,N_27341);
nor U27948 (N_27948,N_27197,N_27403);
or U27949 (N_27949,N_27233,N_27163);
nand U27950 (N_27950,N_27267,N_27042);
nor U27951 (N_27951,N_27411,N_27468);
or U27952 (N_27952,N_27497,N_27387);
or U27953 (N_27953,N_27080,N_27121);
and U27954 (N_27954,N_27135,N_27063);
nand U27955 (N_27955,N_27430,N_27212);
or U27956 (N_27956,N_27401,N_27212);
or U27957 (N_27957,N_27457,N_27122);
nor U27958 (N_27958,N_27325,N_27341);
or U27959 (N_27959,N_27207,N_27347);
and U27960 (N_27960,N_27231,N_27391);
xnor U27961 (N_27961,N_27064,N_27051);
xnor U27962 (N_27962,N_27068,N_27099);
or U27963 (N_27963,N_27443,N_27075);
or U27964 (N_27964,N_27402,N_27479);
or U27965 (N_27965,N_27002,N_27109);
nor U27966 (N_27966,N_27044,N_27062);
and U27967 (N_27967,N_27022,N_27053);
xnor U27968 (N_27968,N_27027,N_27203);
and U27969 (N_27969,N_27133,N_27173);
or U27970 (N_27970,N_27171,N_27443);
xnor U27971 (N_27971,N_27174,N_27178);
xnor U27972 (N_27972,N_27424,N_27156);
nand U27973 (N_27973,N_27040,N_27011);
or U27974 (N_27974,N_27093,N_27359);
or U27975 (N_27975,N_27366,N_27169);
nand U27976 (N_27976,N_27188,N_27443);
nor U27977 (N_27977,N_27070,N_27154);
and U27978 (N_27978,N_27348,N_27247);
xor U27979 (N_27979,N_27079,N_27323);
xnor U27980 (N_27980,N_27230,N_27114);
and U27981 (N_27981,N_27165,N_27176);
nand U27982 (N_27982,N_27240,N_27168);
nand U27983 (N_27983,N_27311,N_27373);
xnor U27984 (N_27984,N_27227,N_27466);
or U27985 (N_27985,N_27298,N_27061);
xor U27986 (N_27986,N_27319,N_27194);
or U27987 (N_27987,N_27159,N_27367);
and U27988 (N_27988,N_27231,N_27230);
and U27989 (N_27989,N_27316,N_27086);
xor U27990 (N_27990,N_27175,N_27198);
and U27991 (N_27991,N_27340,N_27160);
xnor U27992 (N_27992,N_27331,N_27008);
xnor U27993 (N_27993,N_27036,N_27159);
nand U27994 (N_27994,N_27166,N_27348);
nor U27995 (N_27995,N_27275,N_27160);
nor U27996 (N_27996,N_27270,N_27423);
xnor U27997 (N_27997,N_27119,N_27190);
or U27998 (N_27998,N_27391,N_27042);
xnor U27999 (N_27999,N_27179,N_27447);
and U28000 (N_28000,N_27871,N_27822);
nand U28001 (N_28001,N_27753,N_27733);
xnor U28002 (N_28002,N_27672,N_27521);
and U28003 (N_28003,N_27610,N_27951);
or U28004 (N_28004,N_27855,N_27515);
nor U28005 (N_28005,N_27760,N_27660);
and U28006 (N_28006,N_27970,N_27830);
and U28007 (N_28007,N_27815,N_27783);
and U28008 (N_28008,N_27860,N_27594);
nand U28009 (N_28009,N_27957,N_27514);
xor U28010 (N_28010,N_27982,N_27771);
xnor U28011 (N_28011,N_27625,N_27637);
xnor U28012 (N_28012,N_27881,N_27995);
nor U28013 (N_28013,N_27611,N_27589);
and U28014 (N_28014,N_27757,N_27574);
or U28015 (N_28015,N_27615,N_27917);
nor U28016 (N_28016,N_27973,N_27655);
nor U28017 (N_28017,N_27885,N_27890);
nor U28018 (N_28018,N_27579,N_27682);
and U28019 (N_28019,N_27551,N_27712);
nor U28020 (N_28020,N_27513,N_27724);
nand U28021 (N_28021,N_27522,N_27656);
nand U28022 (N_28022,N_27628,N_27525);
xor U28023 (N_28023,N_27511,N_27889);
nand U28024 (N_28024,N_27820,N_27808);
and U28025 (N_28025,N_27903,N_27623);
and U28026 (N_28026,N_27734,N_27572);
nand U28027 (N_28027,N_27592,N_27802);
and U28028 (N_28028,N_27577,N_27788);
and U28029 (N_28029,N_27789,N_27782);
and U28030 (N_28030,N_27718,N_27784);
xnor U28031 (N_28031,N_27739,N_27750);
and U28032 (N_28032,N_27811,N_27945);
nor U28033 (N_28033,N_27727,N_27692);
and U28034 (N_28034,N_27697,N_27747);
or U28035 (N_28035,N_27532,N_27517);
and U28036 (N_28036,N_27569,N_27967);
xor U28037 (N_28037,N_27715,N_27787);
xor U28038 (N_28038,N_27576,N_27858);
xor U28039 (N_28039,N_27506,N_27662);
nand U28040 (N_28040,N_27813,N_27704);
or U28041 (N_28041,N_27588,N_27863);
nand U28042 (N_28042,N_27875,N_27676);
nand U28043 (N_28043,N_27695,N_27999);
nor U28044 (N_28044,N_27596,N_27763);
nand U28045 (N_28045,N_27601,N_27773);
xnor U28046 (N_28046,N_27657,N_27742);
nand U28047 (N_28047,N_27963,N_27624);
and U28048 (N_28048,N_27717,N_27971);
nor U28049 (N_28049,N_27598,N_27994);
or U28050 (N_28050,N_27914,N_27633);
nor U28051 (N_28051,N_27844,N_27546);
or U28052 (N_28052,N_27866,N_27932);
xor U28053 (N_28053,N_27710,N_27582);
nand U28054 (N_28054,N_27671,N_27986);
and U28055 (N_28055,N_27947,N_27984);
and U28056 (N_28056,N_27836,N_27944);
or U28057 (N_28057,N_27975,N_27520);
and U28058 (N_28058,N_27725,N_27910);
nand U28059 (N_28059,N_27849,N_27749);
and U28060 (N_28060,N_27543,N_27703);
xor U28061 (N_28061,N_27557,N_27814);
nand U28062 (N_28062,N_27711,N_27974);
or U28063 (N_28063,N_27832,N_27681);
or U28064 (N_28064,N_27766,N_27578);
nor U28065 (N_28065,N_27927,N_27678);
and U28066 (N_28066,N_27708,N_27983);
nor U28067 (N_28067,N_27799,N_27874);
nor U28068 (N_28068,N_27533,N_27980);
and U28069 (N_28069,N_27843,N_27921);
xor U28070 (N_28070,N_27738,N_27528);
or U28071 (N_28071,N_27503,N_27892);
xor U28072 (N_28072,N_27857,N_27797);
nand U28073 (N_28073,N_27748,N_27674);
and U28074 (N_28074,N_27758,N_27700);
nand U28075 (N_28075,N_27631,N_27809);
nand U28076 (N_28076,N_27691,N_27790);
and U28077 (N_28077,N_27966,N_27846);
or U28078 (N_28078,N_27764,N_27537);
nor U28079 (N_28079,N_27774,N_27746);
or U28080 (N_28080,N_27828,N_27990);
nand U28081 (N_28081,N_27690,N_27805);
nor U28082 (N_28082,N_27544,N_27934);
and U28083 (N_28083,N_27620,N_27547);
xor U28084 (N_28084,N_27895,N_27972);
nor U28085 (N_28085,N_27619,N_27722);
nand U28086 (N_28086,N_27731,N_27987);
or U28087 (N_28087,N_27922,N_27862);
nor U28088 (N_28088,N_27621,N_27698);
nor U28089 (N_28089,N_27768,N_27998);
or U28090 (N_28090,N_27751,N_27996);
and U28091 (N_28091,N_27694,N_27916);
nand U28092 (N_28092,N_27851,N_27640);
nor U28093 (N_28093,N_27949,N_27599);
and U28094 (N_28094,N_27634,N_27867);
xor U28095 (N_28095,N_27791,N_27852);
xnor U28096 (N_28096,N_27906,N_27679);
or U28097 (N_28097,N_27913,N_27804);
or U28098 (N_28098,N_27912,N_27888);
and U28099 (N_28099,N_27507,N_27549);
or U28100 (N_28100,N_27887,N_27705);
xor U28101 (N_28101,N_27882,N_27516);
nor U28102 (N_28102,N_27677,N_27976);
xor U28103 (N_28103,N_27819,N_27564);
or U28104 (N_28104,N_27649,N_27933);
nand U28105 (N_28105,N_27613,N_27591);
and U28106 (N_28106,N_27683,N_27835);
nand U28107 (N_28107,N_27558,N_27540);
and U28108 (N_28108,N_27873,N_27559);
nor U28109 (N_28109,N_27707,N_27985);
nand U28110 (N_28110,N_27940,N_27955);
or U28111 (N_28111,N_27573,N_27523);
nand U28112 (N_28112,N_27584,N_27833);
nand U28113 (N_28113,N_27817,N_27568);
nand U28114 (N_28114,N_27853,N_27919);
and U28115 (N_28115,N_27652,N_27567);
and U28116 (N_28116,N_27670,N_27969);
xor U28117 (N_28117,N_27684,N_27663);
xnor U28118 (N_28118,N_27512,N_27505);
xnor U28119 (N_28119,N_27566,N_27772);
nor U28120 (N_28120,N_27504,N_27847);
nand U28121 (N_28121,N_27597,N_27648);
or U28122 (N_28122,N_27629,N_27931);
or U28123 (N_28123,N_27950,N_27539);
or U28124 (N_28124,N_27880,N_27571);
nor U28125 (N_28125,N_27778,N_27786);
and U28126 (N_28126,N_27765,N_27541);
nor U28127 (N_28127,N_27879,N_27529);
and U28128 (N_28128,N_27926,N_27812);
or U28129 (N_28129,N_27644,N_27500);
or U28130 (N_28130,N_27713,N_27954);
nand U28131 (N_28131,N_27755,N_27997);
and U28132 (N_28132,N_27626,N_27675);
and U28133 (N_28133,N_27759,N_27581);
or U28134 (N_28134,N_27554,N_27794);
and U28135 (N_28135,N_27925,N_27938);
xnor U28136 (N_28136,N_27904,N_27603);
nor U28137 (N_28137,N_27988,N_27896);
or U28138 (N_28138,N_27714,N_27608);
xnor U28139 (N_28139,N_27767,N_27968);
xor U28140 (N_28140,N_27838,N_27732);
or U28141 (N_28141,N_27865,N_27550);
and U28142 (N_28142,N_27840,N_27769);
nand U28143 (N_28143,N_27908,N_27735);
xnor U28144 (N_28144,N_27891,N_27762);
xor U28145 (N_28145,N_27795,N_27510);
xnor U28146 (N_28146,N_27659,N_27709);
or U28147 (N_28147,N_27870,N_27726);
nand U28148 (N_28148,N_27680,N_27884);
nor U28149 (N_28149,N_27531,N_27518);
and U28150 (N_28150,N_27553,N_27941);
nand U28151 (N_28151,N_27807,N_27614);
nand U28152 (N_28152,N_27555,N_27937);
nand U28153 (N_28153,N_27992,N_27575);
nand U28154 (N_28154,N_27590,N_27991);
nor U28155 (N_28155,N_27989,N_27962);
nor U28156 (N_28156,N_27756,N_27856);
xor U28157 (N_28157,N_27686,N_27861);
xor U28158 (N_28158,N_27607,N_27897);
xor U28159 (N_28159,N_27741,N_27744);
nand U28160 (N_28160,N_27754,N_27622);
nand U28161 (N_28161,N_27929,N_27716);
nand U28162 (N_28162,N_27743,N_27918);
nand U28163 (N_28163,N_27701,N_27570);
nor U28164 (N_28164,N_27580,N_27508);
nor U28165 (N_28165,N_27924,N_27561);
nand U28166 (N_28166,N_27893,N_27850);
xor U28167 (N_28167,N_27779,N_27668);
and U28168 (N_28168,N_27605,N_27770);
and U28169 (N_28169,N_27859,N_27792);
and U28170 (N_28170,N_27501,N_27827);
xnor U28171 (N_28171,N_27693,N_27593);
nor U28172 (N_28172,N_27687,N_27872);
and U28173 (N_28173,N_27689,N_27667);
and U28174 (N_28174,N_27665,N_27720);
nand U28175 (N_28175,N_27796,N_27647);
xnor U28176 (N_28176,N_27978,N_27563);
nand U28177 (N_28177,N_27864,N_27905);
nand U28178 (N_28178,N_27651,N_27638);
xor U28179 (N_28179,N_27509,N_27816);
nand U28180 (N_28180,N_27781,N_27823);
and U28181 (N_28181,N_27834,N_27900);
nor U28182 (N_28182,N_27818,N_27842);
nand U28183 (N_28183,N_27946,N_27630);
nand U28184 (N_28184,N_27752,N_27534);
and U28185 (N_28185,N_27837,N_27587);
or U28186 (N_28186,N_27848,N_27639);
and U28187 (N_28187,N_27723,N_27803);
or U28188 (N_28188,N_27894,N_27761);
and U28189 (N_28189,N_27736,N_27979);
nor U28190 (N_28190,N_27530,N_27923);
xnor U28191 (N_28191,N_27536,N_27737);
nor U28192 (N_28192,N_27775,N_27977);
nand U28193 (N_28193,N_27911,N_27801);
and U28194 (N_28194,N_27653,N_27928);
or U28195 (N_28195,N_27901,N_27777);
or U28196 (N_28196,N_27606,N_27604);
or U28197 (N_28197,N_27959,N_27953);
or U28198 (N_28198,N_27699,N_27961);
xor U28199 (N_28199,N_27646,N_27943);
nand U28200 (N_28200,N_27664,N_27907);
nand U28201 (N_28201,N_27920,N_27616);
nand U28202 (N_28202,N_27658,N_27826);
nand U28203 (N_28203,N_27930,N_27650);
and U28204 (N_28204,N_27902,N_27958);
xnor U28205 (N_28205,N_27627,N_27876);
nor U28206 (N_28206,N_27706,N_27824);
nand U28207 (N_28207,N_27981,N_27810);
xnor U28208 (N_28208,N_27556,N_27585);
and U28209 (N_28209,N_27780,N_27642);
xnor U28210 (N_28210,N_27798,N_27821);
xor U28211 (N_28211,N_27645,N_27730);
and U28212 (N_28212,N_27909,N_27740);
or U28213 (N_28213,N_27854,N_27562);
nor U28214 (N_28214,N_27939,N_27696);
xor U28215 (N_28215,N_27868,N_27524);
nand U28216 (N_28216,N_27538,N_27565);
and U28217 (N_28217,N_27560,N_27719);
nor U28218 (N_28218,N_27702,N_27728);
nor U28219 (N_28219,N_27600,N_27785);
or U28220 (N_28220,N_27643,N_27673);
or U28221 (N_28221,N_27845,N_27898);
xnor U28222 (N_28222,N_27636,N_27877);
nand U28223 (N_28223,N_27685,N_27964);
or U28224 (N_28224,N_27552,N_27502);
xnor U28225 (N_28225,N_27915,N_27899);
nand U28226 (N_28226,N_27806,N_27635);
nand U28227 (N_28227,N_27545,N_27519);
and U28228 (N_28228,N_27793,N_27841);
or U28229 (N_28229,N_27745,N_27542);
or U28230 (N_28230,N_27883,N_27869);
xnor U28231 (N_28231,N_27595,N_27800);
or U28232 (N_28232,N_27831,N_27878);
and U28233 (N_28233,N_27956,N_27993);
nor U28234 (N_28234,N_27632,N_27776);
nor U28235 (N_28235,N_27526,N_27935);
nand U28236 (N_28236,N_27942,N_27948);
nor U28237 (N_28237,N_27548,N_27965);
nor U28238 (N_28238,N_27825,N_27661);
nor U28239 (N_28239,N_27617,N_27535);
or U28240 (N_28240,N_27729,N_27666);
nor U28241 (N_28241,N_27527,N_27721);
xnor U28242 (N_28242,N_27641,N_27936);
xnor U28243 (N_28243,N_27612,N_27886);
xor U28244 (N_28244,N_27654,N_27669);
xor U28245 (N_28245,N_27952,N_27609);
nand U28246 (N_28246,N_27602,N_27586);
xor U28247 (N_28247,N_27583,N_27960);
nor U28248 (N_28248,N_27829,N_27688);
nand U28249 (N_28249,N_27618,N_27839);
or U28250 (N_28250,N_27553,N_27932);
or U28251 (N_28251,N_27579,N_27611);
or U28252 (N_28252,N_27759,N_27534);
nor U28253 (N_28253,N_27666,N_27900);
or U28254 (N_28254,N_27606,N_27999);
xnor U28255 (N_28255,N_27688,N_27963);
nor U28256 (N_28256,N_27878,N_27873);
nor U28257 (N_28257,N_27593,N_27895);
nand U28258 (N_28258,N_27634,N_27560);
and U28259 (N_28259,N_27964,N_27500);
xor U28260 (N_28260,N_27591,N_27521);
xnor U28261 (N_28261,N_27597,N_27509);
nor U28262 (N_28262,N_27518,N_27568);
nor U28263 (N_28263,N_27699,N_27556);
nand U28264 (N_28264,N_27799,N_27770);
nor U28265 (N_28265,N_27640,N_27983);
or U28266 (N_28266,N_27703,N_27580);
nor U28267 (N_28267,N_27774,N_27741);
nand U28268 (N_28268,N_27747,N_27995);
xnor U28269 (N_28269,N_27881,N_27722);
xnor U28270 (N_28270,N_27871,N_27574);
or U28271 (N_28271,N_27934,N_27501);
nand U28272 (N_28272,N_27710,N_27847);
nor U28273 (N_28273,N_27716,N_27813);
xnor U28274 (N_28274,N_27709,N_27830);
nand U28275 (N_28275,N_27951,N_27626);
nand U28276 (N_28276,N_27914,N_27688);
nor U28277 (N_28277,N_27767,N_27913);
or U28278 (N_28278,N_27537,N_27714);
nor U28279 (N_28279,N_27593,N_27833);
and U28280 (N_28280,N_27860,N_27641);
nor U28281 (N_28281,N_27817,N_27933);
and U28282 (N_28282,N_27864,N_27722);
or U28283 (N_28283,N_27967,N_27703);
nand U28284 (N_28284,N_27520,N_27924);
and U28285 (N_28285,N_27741,N_27710);
xor U28286 (N_28286,N_27678,N_27846);
xnor U28287 (N_28287,N_27916,N_27842);
and U28288 (N_28288,N_27754,N_27976);
and U28289 (N_28289,N_27825,N_27915);
nand U28290 (N_28290,N_27979,N_27913);
xor U28291 (N_28291,N_27605,N_27518);
nand U28292 (N_28292,N_27667,N_27634);
and U28293 (N_28293,N_27504,N_27771);
nor U28294 (N_28294,N_27517,N_27743);
nor U28295 (N_28295,N_27625,N_27603);
nor U28296 (N_28296,N_27839,N_27716);
and U28297 (N_28297,N_27723,N_27647);
xnor U28298 (N_28298,N_27876,N_27685);
and U28299 (N_28299,N_27994,N_27799);
nand U28300 (N_28300,N_27556,N_27965);
nand U28301 (N_28301,N_27567,N_27653);
or U28302 (N_28302,N_27590,N_27654);
xnor U28303 (N_28303,N_27522,N_27662);
nand U28304 (N_28304,N_27739,N_27838);
or U28305 (N_28305,N_27617,N_27967);
xor U28306 (N_28306,N_27618,N_27807);
xnor U28307 (N_28307,N_27668,N_27727);
nand U28308 (N_28308,N_27931,N_27994);
xnor U28309 (N_28309,N_27897,N_27638);
or U28310 (N_28310,N_27808,N_27634);
nor U28311 (N_28311,N_27540,N_27615);
or U28312 (N_28312,N_27821,N_27801);
or U28313 (N_28313,N_27668,N_27960);
and U28314 (N_28314,N_27630,N_27515);
nor U28315 (N_28315,N_27930,N_27949);
and U28316 (N_28316,N_27606,N_27536);
nand U28317 (N_28317,N_27724,N_27775);
nand U28318 (N_28318,N_27836,N_27529);
or U28319 (N_28319,N_27889,N_27516);
xor U28320 (N_28320,N_27730,N_27616);
and U28321 (N_28321,N_27637,N_27751);
nand U28322 (N_28322,N_27533,N_27735);
and U28323 (N_28323,N_27917,N_27738);
and U28324 (N_28324,N_27643,N_27698);
and U28325 (N_28325,N_27659,N_27608);
xnor U28326 (N_28326,N_27627,N_27891);
and U28327 (N_28327,N_27760,N_27836);
and U28328 (N_28328,N_27883,N_27916);
or U28329 (N_28329,N_27988,N_27734);
nand U28330 (N_28330,N_27919,N_27623);
or U28331 (N_28331,N_27668,N_27598);
xnor U28332 (N_28332,N_27626,N_27625);
xor U28333 (N_28333,N_27702,N_27932);
nand U28334 (N_28334,N_27862,N_27511);
or U28335 (N_28335,N_27798,N_27571);
nor U28336 (N_28336,N_27754,N_27874);
or U28337 (N_28337,N_27864,N_27757);
nand U28338 (N_28338,N_27984,N_27928);
nand U28339 (N_28339,N_27759,N_27853);
xor U28340 (N_28340,N_27711,N_27575);
or U28341 (N_28341,N_27612,N_27573);
nor U28342 (N_28342,N_27529,N_27898);
or U28343 (N_28343,N_27781,N_27750);
nor U28344 (N_28344,N_27548,N_27560);
or U28345 (N_28345,N_27994,N_27693);
and U28346 (N_28346,N_27658,N_27562);
nor U28347 (N_28347,N_27651,N_27660);
or U28348 (N_28348,N_27709,N_27801);
xor U28349 (N_28349,N_27947,N_27893);
nor U28350 (N_28350,N_27551,N_27875);
or U28351 (N_28351,N_27910,N_27991);
and U28352 (N_28352,N_27536,N_27768);
or U28353 (N_28353,N_27969,N_27757);
and U28354 (N_28354,N_27709,N_27763);
nor U28355 (N_28355,N_27683,N_27976);
or U28356 (N_28356,N_27989,N_27603);
xor U28357 (N_28357,N_27535,N_27732);
nand U28358 (N_28358,N_27853,N_27655);
and U28359 (N_28359,N_27978,N_27709);
and U28360 (N_28360,N_27631,N_27660);
xnor U28361 (N_28361,N_27630,N_27612);
nor U28362 (N_28362,N_27896,N_27692);
nor U28363 (N_28363,N_27506,N_27579);
xnor U28364 (N_28364,N_27909,N_27910);
nor U28365 (N_28365,N_27722,N_27998);
and U28366 (N_28366,N_27898,N_27935);
nor U28367 (N_28367,N_27604,N_27882);
nand U28368 (N_28368,N_27911,N_27523);
nand U28369 (N_28369,N_27857,N_27791);
nand U28370 (N_28370,N_27589,N_27568);
nor U28371 (N_28371,N_27788,N_27850);
xor U28372 (N_28372,N_27663,N_27658);
and U28373 (N_28373,N_27956,N_27725);
or U28374 (N_28374,N_27789,N_27761);
nor U28375 (N_28375,N_27617,N_27705);
nor U28376 (N_28376,N_27757,N_27698);
and U28377 (N_28377,N_27904,N_27755);
xnor U28378 (N_28378,N_27537,N_27884);
nor U28379 (N_28379,N_27935,N_27601);
or U28380 (N_28380,N_27861,N_27715);
nor U28381 (N_28381,N_27783,N_27587);
nor U28382 (N_28382,N_27970,N_27978);
and U28383 (N_28383,N_27795,N_27800);
xnor U28384 (N_28384,N_27949,N_27523);
nor U28385 (N_28385,N_27971,N_27925);
nand U28386 (N_28386,N_27557,N_27794);
xnor U28387 (N_28387,N_27862,N_27949);
nor U28388 (N_28388,N_27975,N_27534);
nand U28389 (N_28389,N_27809,N_27752);
nand U28390 (N_28390,N_27553,N_27827);
nand U28391 (N_28391,N_27752,N_27619);
or U28392 (N_28392,N_27986,N_27944);
xor U28393 (N_28393,N_27567,N_27660);
or U28394 (N_28394,N_27826,N_27987);
nand U28395 (N_28395,N_27868,N_27835);
or U28396 (N_28396,N_27825,N_27500);
xor U28397 (N_28397,N_27959,N_27629);
and U28398 (N_28398,N_27878,N_27949);
and U28399 (N_28399,N_27533,N_27573);
nand U28400 (N_28400,N_27688,N_27955);
xnor U28401 (N_28401,N_27617,N_27979);
and U28402 (N_28402,N_27584,N_27966);
nor U28403 (N_28403,N_27813,N_27602);
nor U28404 (N_28404,N_27808,N_27933);
nor U28405 (N_28405,N_27861,N_27768);
xor U28406 (N_28406,N_27726,N_27722);
nand U28407 (N_28407,N_27969,N_27593);
xnor U28408 (N_28408,N_27873,N_27862);
nor U28409 (N_28409,N_27666,N_27950);
xnor U28410 (N_28410,N_27703,N_27662);
and U28411 (N_28411,N_27552,N_27623);
and U28412 (N_28412,N_27502,N_27808);
nor U28413 (N_28413,N_27545,N_27901);
and U28414 (N_28414,N_27577,N_27872);
xnor U28415 (N_28415,N_27685,N_27887);
or U28416 (N_28416,N_27684,N_27937);
or U28417 (N_28417,N_27801,N_27599);
nor U28418 (N_28418,N_27532,N_27559);
and U28419 (N_28419,N_27615,N_27780);
nor U28420 (N_28420,N_27573,N_27780);
nand U28421 (N_28421,N_27639,N_27511);
and U28422 (N_28422,N_27978,N_27766);
and U28423 (N_28423,N_27781,N_27559);
nand U28424 (N_28424,N_27515,N_27553);
nand U28425 (N_28425,N_27998,N_27640);
nand U28426 (N_28426,N_27576,N_27910);
nand U28427 (N_28427,N_27836,N_27925);
or U28428 (N_28428,N_27505,N_27878);
xnor U28429 (N_28429,N_27881,N_27625);
nand U28430 (N_28430,N_27744,N_27559);
and U28431 (N_28431,N_27842,N_27879);
and U28432 (N_28432,N_27966,N_27704);
and U28433 (N_28433,N_27726,N_27741);
xor U28434 (N_28434,N_27961,N_27685);
nor U28435 (N_28435,N_27842,N_27770);
nand U28436 (N_28436,N_27778,N_27686);
and U28437 (N_28437,N_27841,N_27565);
xnor U28438 (N_28438,N_27560,N_27561);
xor U28439 (N_28439,N_27645,N_27699);
and U28440 (N_28440,N_27541,N_27523);
nor U28441 (N_28441,N_27597,N_27649);
or U28442 (N_28442,N_27685,N_27772);
nand U28443 (N_28443,N_27774,N_27539);
xor U28444 (N_28444,N_27844,N_27566);
and U28445 (N_28445,N_27951,N_27751);
or U28446 (N_28446,N_27847,N_27902);
and U28447 (N_28447,N_27759,N_27821);
or U28448 (N_28448,N_27914,N_27516);
and U28449 (N_28449,N_27742,N_27631);
and U28450 (N_28450,N_27619,N_27706);
nand U28451 (N_28451,N_27784,N_27602);
or U28452 (N_28452,N_27642,N_27814);
or U28453 (N_28453,N_27845,N_27925);
or U28454 (N_28454,N_27911,N_27790);
xor U28455 (N_28455,N_27774,N_27784);
xnor U28456 (N_28456,N_27510,N_27858);
or U28457 (N_28457,N_27850,N_27765);
and U28458 (N_28458,N_27796,N_27523);
xor U28459 (N_28459,N_27606,N_27502);
xor U28460 (N_28460,N_27942,N_27689);
xor U28461 (N_28461,N_27772,N_27719);
nor U28462 (N_28462,N_27813,N_27998);
nand U28463 (N_28463,N_27580,N_27846);
xnor U28464 (N_28464,N_27540,N_27928);
and U28465 (N_28465,N_27562,N_27822);
or U28466 (N_28466,N_27726,N_27599);
nand U28467 (N_28467,N_27794,N_27708);
nand U28468 (N_28468,N_27855,N_27728);
and U28469 (N_28469,N_27801,N_27857);
nand U28470 (N_28470,N_27971,N_27663);
and U28471 (N_28471,N_27954,N_27831);
nand U28472 (N_28472,N_27506,N_27597);
xnor U28473 (N_28473,N_27554,N_27693);
nor U28474 (N_28474,N_27825,N_27806);
and U28475 (N_28475,N_27698,N_27648);
nand U28476 (N_28476,N_27713,N_27700);
nor U28477 (N_28477,N_27531,N_27970);
nor U28478 (N_28478,N_27876,N_27606);
nor U28479 (N_28479,N_27976,N_27634);
or U28480 (N_28480,N_27567,N_27671);
nor U28481 (N_28481,N_27502,N_27644);
or U28482 (N_28482,N_27504,N_27991);
and U28483 (N_28483,N_27562,N_27783);
and U28484 (N_28484,N_27948,N_27969);
nand U28485 (N_28485,N_27612,N_27737);
nand U28486 (N_28486,N_27745,N_27527);
nor U28487 (N_28487,N_27836,N_27993);
and U28488 (N_28488,N_27559,N_27579);
xor U28489 (N_28489,N_27917,N_27976);
or U28490 (N_28490,N_27543,N_27859);
xor U28491 (N_28491,N_27654,N_27989);
nand U28492 (N_28492,N_27827,N_27954);
nand U28493 (N_28493,N_27598,N_27570);
xnor U28494 (N_28494,N_27687,N_27768);
or U28495 (N_28495,N_27884,N_27844);
nor U28496 (N_28496,N_27594,N_27801);
nand U28497 (N_28497,N_27771,N_27646);
and U28498 (N_28498,N_27674,N_27945);
nor U28499 (N_28499,N_27535,N_27638);
or U28500 (N_28500,N_28238,N_28248);
nand U28501 (N_28501,N_28000,N_28343);
nand U28502 (N_28502,N_28329,N_28026);
nand U28503 (N_28503,N_28449,N_28084);
and U28504 (N_28504,N_28482,N_28063);
and U28505 (N_28505,N_28261,N_28221);
or U28506 (N_28506,N_28057,N_28441);
nand U28507 (N_28507,N_28494,N_28283);
and U28508 (N_28508,N_28282,N_28196);
and U28509 (N_28509,N_28170,N_28131);
xor U28510 (N_28510,N_28281,N_28188);
xnor U28511 (N_28511,N_28056,N_28478);
nand U28512 (N_28512,N_28105,N_28124);
or U28513 (N_28513,N_28076,N_28194);
xor U28514 (N_28514,N_28108,N_28390);
nand U28515 (N_28515,N_28177,N_28456);
and U28516 (N_28516,N_28336,N_28290);
nand U28517 (N_28517,N_28444,N_28380);
nor U28518 (N_28518,N_28361,N_28096);
xnor U28519 (N_28519,N_28373,N_28357);
and U28520 (N_28520,N_28067,N_28364);
nand U28521 (N_28521,N_28493,N_28189);
and U28522 (N_28522,N_28034,N_28333);
nor U28523 (N_28523,N_28028,N_28435);
xor U28524 (N_28524,N_28032,N_28351);
nor U28525 (N_28525,N_28392,N_28337);
or U28526 (N_28526,N_28134,N_28440);
or U28527 (N_28527,N_28497,N_28422);
nor U28528 (N_28528,N_28166,N_28182);
nand U28529 (N_28529,N_28437,N_28088);
xor U28530 (N_28530,N_28220,N_28447);
xor U28531 (N_28531,N_28078,N_28402);
nand U28532 (N_28532,N_28274,N_28498);
xnor U28533 (N_28533,N_28383,N_28163);
xor U28534 (N_28534,N_28058,N_28098);
and U28535 (N_28535,N_28403,N_28388);
xnor U28536 (N_28536,N_28037,N_28050);
nand U28537 (N_28537,N_28312,N_28273);
nand U28538 (N_28538,N_28125,N_28384);
nor U28539 (N_28539,N_28216,N_28095);
nor U28540 (N_28540,N_28399,N_28161);
xnor U28541 (N_28541,N_28467,N_28345);
and U28542 (N_28542,N_28442,N_28160);
xor U28543 (N_28543,N_28300,N_28229);
xnor U28544 (N_28544,N_28480,N_28287);
and U28545 (N_28545,N_28374,N_28142);
nand U28546 (N_28546,N_28239,N_28100);
or U28547 (N_28547,N_28330,N_28272);
or U28548 (N_28548,N_28060,N_28307);
nand U28549 (N_28549,N_28308,N_28211);
xor U28550 (N_28550,N_28301,N_28230);
xor U28551 (N_28551,N_28315,N_28214);
nor U28552 (N_28552,N_28020,N_28203);
nor U28553 (N_28553,N_28346,N_28126);
or U28554 (N_28554,N_28303,N_28350);
and U28555 (N_28555,N_28109,N_28049);
nor U28556 (N_28556,N_28231,N_28218);
nor U28557 (N_28557,N_28054,N_28094);
xor U28558 (N_28558,N_28327,N_28097);
nand U28559 (N_28559,N_28082,N_28148);
xor U28560 (N_28560,N_28326,N_28025);
and U28561 (N_28561,N_28270,N_28349);
or U28562 (N_28562,N_28068,N_28314);
and U28563 (N_28563,N_28171,N_28495);
nand U28564 (N_28564,N_28217,N_28065);
or U28565 (N_28565,N_28372,N_28075);
nand U28566 (N_28566,N_28284,N_28450);
nor U28567 (N_28567,N_28199,N_28077);
nand U28568 (N_28568,N_28260,N_28258);
or U28569 (N_28569,N_28409,N_28293);
nor U28570 (N_28570,N_28130,N_28431);
nand U28571 (N_28571,N_28045,N_28458);
nor U28572 (N_28572,N_28310,N_28288);
nand U28573 (N_28573,N_28492,N_28087);
or U28574 (N_28574,N_28061,N_28164);
nor U28575 (N_28575,N_28285,N_28002);
xor U28576 (N_28576,N_28454,N_28240);
xor U28577 (N_28577,N_28404,N_28257);
and U28578 (N_28578,N_28340,N_28022);
nand U28579 (N_28579,N_28151,N_28139);
nor U28580 (N_28580,N_28079,N_28064);
xnor U28581 (N_28581,N_28427,N_28243);
xnor U28582 (N_28582,N_28011,N_28093);
nor U28583 (N_28583,N_28006,N_28407);
xor U28584 (N_28584,N_28292,N_28021);
xnor U28585 (N_28585,N_28081,N_28204);
nor U28586 (N_28586,N_28213,N_28224);
xnor U28587 (N_28587,N_28018,N_28222);
xnor U28588 (N_28588,N_28195,N_28267);
and U28589 (N_28589,N_28236,N_28086);
nand U28590 (N_28590,N_28143,N_28269);
xnor U28591 (N_28591,N_28294,N_28235);
or U28592 (N_28592,N_28119,N_28448);
nor U28593 (N_28593,N_28016,N_28223);
or U28594 (N_28594,N_28190,N_28136);
xor U28595 (N_28595,N_28443,N_28365);
nand U28596 (N_28596,N_28279,N_28362);
and U28597 (N_28597,N_28127,N_28371);
and U28598 (N_28598,N_28378,N_28145);
and U28599 (N_28599,N_28089,N_28162);
and U28600 (N_28600,N_28241,N_28271);
nor U28601 (N_28601,N_28410,N_28138);
nor U28602 (N_28602,N_28265,N_28379);
and U28603 (N_28603,N_28387,N_28040);
xnor U28604 (N_28604,N_28367,N_28348);
xnor U28605 (N_28605,N_28335,N_28116);
and U28606 (N_28606,N_28416,N_28186);
nand U28607 (N_28607,N_28090,N_28484);
xor U28608 (N_28608,N_28320,N_28004);
or U28609 (N_28609,N_28062,N_28318);
nor U28610 (N_28610,N_28313,N_28117);
and U28611 (N_28611,N_28154,N_28152);
nor U28612 (N_28612,N_28246,N_28280);
xnor U28613 (N_28613,N_28092,N_28453);
nand U28614 (N_28614,N_28244,N_28245);
xnor U28615 (N_28615,N_28027,N_28219);
nor U28616 (N_28616,N_28496,N_28368);
nor U28617 (N_28617,N_28069,N_28418);
xnor U28618 (N_28618,N_28356,N_28415);
and U28619 (N_28619,N_28396,N_28306);
nand U28620 (N_28620,N_28200,N_28059);
xor U28621 (N_28621,N_28042,N_28499);
or U28622 (N_28622,N_28311,N_28150);
nand U28623 (N_28623,N_28429,N_28316);
or U28624 (N_28624,N_28250,N_28474);
or U28625 (N_28625,N_28173,N_28375);
nor U28626 (N_28626,N_28408,N_28353);
or U28627 (N_28627,N_28470,N_28234);
xor U28628 (N_28628,N_28401,N_28029);
xnor U28629 (N_28629,N_28339,N_28420);
or U28630 (N_28630,N_28237,N_28263);
xnor U28631 (N_28631,N_28347,N_28299);
or U28632 (N_28632,N_28354,N_28485);
xor U28633 (N_28633,N_28074,N_28111);
xor U28634 (N_28634,N_28465,N_28317);
nor U28635 (N_28635,N_28428,N_28472);
and U28636 (N_28636,N_28191,N_28023);
and U28637 (N_28637,N_28133,N_28319);
and U28638 (N_28638,N_28490,N_28370);
nor U28639 (N_28639,N_28183,N_28035);
nand U28640 (N_28640,N_28338,N_28225);
xnor U28641 (N_28641,N_28102,N_28107);
or U28642 (N_28642,N_28426,N_28406);
xor U28643 (N_28643,N_28491,N_28479);
and U28644 (N_28644,N_28413,N_28425);
or U28645 (N_28645,N_28297,N_28192);
nand U28646 (N_28646,N_28181,N_28039);
xnor U28647 (N_28647,N_28405,N_28120);
and U28648 (N_28648,N_28210,N_28174);
xor U28649 (N_28649,N_28298,N_28206);
xor U28650 (N_28650,N_28172,N_28158);
nand U28651 (N_28651,N_28466,N_28278);
nor U28652 (N_28652,N_28007,N_28106);
and U28653 (N_28653,N_28205,N_28009);
and U28654 (N_28654,N_28460,N_28381);
or U28655 (N_28655,N_28080,N_28430);
and U28656 (N_28656,N_28382,N_28457);
xnor U28657 (N_28657,N_28101,N_28038);
nor U28658 (N_28658,N_28122,N_28424);
nand U28659 (N_28659,N_28099,N_28398);
or U28660 (N_28660,N_28156,N_28411);
nor U28661 (N_28661,N_28013,N_28135);
and U28662 (N_28662,N_28473,N_28085);
nand U28663 (N_28663,N_28197,N_28155);
nor U28664 (N_28664,N_28389,N_28147);
or U28665 (N_28665,N_28209,N_28255);
xor U28666 (N_28666,N_28475,N_28385);
and U28667 (N_28667,N_28008,N_28397);
and U28668 (N_28668,N_28129,N_28024);
nand U28669 (N_28669,N_28198,N_28412);
and U28670 (N_28670,N_28305,N_28140);
or U28671 (N_28671,N_28488,N_28462);
xnor U28672 (N_28672,N_28321,N_28352);
or U28673 (N_28673,N_28187,N_28159);
and U28674 (N_28674,N_28423,N_28463);
nor U28675 (N_28675,N_28328,N_28275);
and U28676 (N_28676,N_28331,N_28110);
nor U28677 (N_28677,N_28168,N_28052);
xor U28678 (N_28678,N_28066,N_28141);
nor U28679 (N_28679,N_28344,N_28010);
nand U28680 (N_28680,N_28358,N_28193);
and U28681 (N_28681,N_28157,N_28451);
xnor U28682 (N_28682,N_28167,N_28091);
or U28683 (N_28683,N_28323,N_28259);
and U28684 (N_28684,N_28048,N_28070);
and U28685 (N_28685,N_28417,N_28366);
and U28686 (N_28686,N_28019,N_28377);
or U28687 (N_28687,N_28446,N_28169);
xnor U28688 (N_28688,N_28264,N_28291);
nand U28689 (N_28689,N_28179,N_28262);
nor U28690 (N_28690,N_28252,N_28268);
nor U28691 (N_28691,N_28289,N_28341);
and U28692 (N_28692,N_28031,N_28251);
nand U28693 (N_28693,N_28360,N_28247);
or U28694 (N_28694,N_28487,N_28342);
nor U28695 (N_28695,N_28051,N_28232);
xor U28696 (N_28696,N_28001,N_28432);
or U28697 (N_28697,N_28137,N_28180);
or U28698 (N_28698,N_28014,N_28419);
nor U28699 (N_28699,N_28445,N_28266);
xnor U28700 (N_28700,N_28144,N_28121);
nand U28701 (N_28701,N_28277,N_28047);
xor U28702 (N_28702,N_28153,N_28322);
or U28703 (N_28703,N_28112,N_28053);
nor U28704 (N_28704,N_28072,N_28477);
and U28705 (N_28705,N_28071,N_28455);
xnor U28706 (N_28706,N_28176,N_28207);
xnor U28707 (N_28707,N_28212,N_28421);
xor U28708 (N_28708,N_28332,N_28483);
nand U28709 (N_28709,N_28215,N_28132);
and U28710 (N_28710,N_28304,N_28175);
and U28711 (N_28711,N_28334,N_28227);
nand U28712 (N_28712,N_28296,N_28184);
nand U28713 (N_28713,N_28471,N_28030);
nand U28714 (N_28714,N_28386,N_28073);
nor U28715 (N_28715,N_28185,N_28489);
or U28716 (N_28716,N_28041,N_28165);
nor U28717 (N_28717,N_28468,N_28146);
nand U28718 (N_28718,N_28395,N_28128);
nor U28719 (N_28719,N_28434,N_28391);
nor U28720 (N_28720,N_28005,N_28043);
nor U28721 (N_28721,N_28439,N_28438);
nor U28722 (N_28722,N_28414,N_28433);
or U28723 (N_28723,N_28233,N_28113);
or U28724 (N_28724,N_28242,N_28461);
xor U28725 (N_28725,N_28118,N_28309);
and U28726 (N_28726,N_28452,N_28149);
nand U28727 (N_28727,N_28178,N_28228);
xnor U28728 (N_28728,N_28201,N_28481);
xor U28729 (N_28729,N_28459,N_28363);
or U28730 (N_28730,N_28104,N_28355);
nand U28731 (N_28731,N_28044,N_28254);
nand U28732 (N_28732,N_28302,N_28055);
nand U28733 (N_28733,N_28015,N_28394);
nand U28734 (N_28734,N_28486,N_28046);
and U28735 (N_28735,N_28017,N_28226);
nor U28736 (N_28736,N_28436,N_28276);
nand U28737 (N_28737,N_28253,N_28295);
and U28738 (N_28738,N_28286,N_28202);
xor U28739 (N_28739,N_28400,N_28476);
nor U28740 (N_28740,N_28115,N_28359);
nand U28741 (N_28741,N_28376,N_28256);
and U28742 (N_28742,N_28393,N_28325);
nand U28743 (N_28743,N_28369,N_28012);
and U28744 (N_28744,N_28036,N_28469);
or U28745 (N_28745,N_28103,N_28464);
and U28746 (N_28746,N_28123,N_28249);
nand U28747 (N_28747,N_28083,N_28324);
and U28748 (N_28748,N_28003,N_28208);
and U28749 (N_28749,N_28114,N_28033);
nor U28750 (N_28750,N_28263,N_28496);
or U28751 (N_28751,N_28482,N_28401);
nand U28752 (N_28752,N_28232,N_28452);
xnor U28753 (N_28753,N_28286,N_28314);
nor U28754 (N_28754,N_28453,N_28233);
or U28755 (N_28755,N_28401,N_28113);
nor U28756 (N_28756,N_28242,N_28067);
or U28757 (N_28757,N_28169,N_28105);
nor U28758 (N_28758,N_28219,N_28328);
or U28759 (N_28759,N_28098,N_28346);
and U28760 (N_28760,N_28276,N_28052);
nor U28761 (N_28761,N_28146,N_28022);
and U28762 (N_28762,N_28226,N_28362);
or U28763 (N_28763,N_28482,N_28466);
xor U28764 (N_28764,N_28332,N_28154);
and U28765 (N_28765,N_28089,N_28473);
xor U28766 (N_28766,N_28148,N_28149);
nand U28767 (N_28767,N_28267,N_28164);
or U28768 (N_28768,N_28125,N_28462);
nor U28769 (N_28769,N_28173,N_28277);
nand U28770 (N_28770,N_28200,N_28006);
xnor U28771 (N_28771,N_28109,N_28081);
or U28772 (N_28772,N_28197,N_28381);
xor U28773 (N_28773,N_28252,N_28178);
nand U28774 (N_28774,N_28417,N_28358);
nand U28775 (N_28775,N_28338,N_28358);
or U28776 (N_28776,N_28433,N_28489);
nor U28777 (N_28777,N_28018,N_28015);
nand U28778 (N_28778,N_28272,N_28110);
xor U28779 (N_28779,N_28408,N_28482);
nor U28780 (N_28780,N_28180,N_28006);
nand U28781 (N_28781,N_28142,N_28402);
or U28782 (N_28782,N_28479,N_28322);
and U28783 (N_28783,N_28438,N_28478);
nor U28784 (N_28784,N_28175,N_28410);
or U28785 (N_28785,N_28120,N_28130);
xor U28786 (N_28786,N_28078,N_28063);
and U28787 (N_28787,N_28328,N_28471);
nand U28788 (N_28788,N_28012,N_28443);
nor U28789 (N_28789,N_28229,N_28186);
nand U28790 (N_28790,N_28054,N_28384);
nand U28791 (N_28791,N_28187,N_28195);
nor U28792 (N_28792,N_28128,N_28093);
or U28793 (N_28793,N_28420,N_28461);
xnor U28794 (N_28794,N_28496,N_28077);
or U28795 (N_28795,N_28411,N_28215);
nor U28796 (N_28796,N_28072,N_28468);
or U28797 (N_28797,N_28136,N_28284);
nor U28798 (N_28798,N_28319,N_28197);
xor U28799 (N_28799,N_28173,N_28314);
nor U28800 (N_28800,N_28428,N_28039);
xor U28801 (N_28801,N_28203,N_28333);
nor U28802 (N_28802,N_28309,N_28472);
nand U28803 (N_28803,N_28386,N_28182);
or U28804 (N_28804,N_28344,N_28499);
nand U28805 (N_28805,N_28059,N_28474);
nor U28806 (N_28806,N_28302,N_28077);
xor U28807 (N_28807,N_28058,N_28191);
nand U28808 (N_28808,N_28073,N_28421);
nand U28809 (N_28809,N_28187,N_28224);
and U28810 (N_28810,N_28423,N_28026);
or U28811 (N_28811,N_28080,N_28349);
or U28812 (N_28812,N_28435,N_28372);
xor U28813 (N_28813,N_28415,N_28009);
and U28814 (N_28814,N_28339,N_28479);
or U28815 (N_28815,N_28387,N_28129);
xnor U28816 (N_28816,N_28359,N_28416);
nand U28817 (N_28817,N_28312,N_28357);
nand U28818 (N_28818,N_28174,N_28102);
and U28819 (N_28819,N_28439,N_28003);
and U28820 (N_28820,N_28159,N_28058);
nor U28821 (N_28821,N_28042,N_28411);
xnor U28822 (N_28822,N_28043,N_28269);
xnor U28823 (N_28823,N_28482,N_28124);
and U28824 (N_28824,N_28309,N_28460);
xnor U28825 (N_28825,N_28334,N_28222);
and U28826 (N_28826,N_28303,N_28022);
or U28827 (N_28827,N_28036,N_28353);
or U28828 (N_28828,N_28150,N_28263);
xor U28829 (N_28829,N_28217,N_28008);
nand U28830 (N_28830,N_28158,N_28062);
xor U28831 (N_28831,N_28052,N_28046);
and U28832 (N_28832,N_28259,N_28005);
and U28833 (N_28833,N_28422,N_28359);
xor U28834 (N_28834,N_28210,N_28037);
nand U28835 (N_28835,N_28049,N_28275);
nor U28836 (N_28836,N_28030,N_28206);
and U28837 (N_28837,N_28429,N_28233);
nor U28838 (N_28838,N_28021,N_28475);
xor U28839 (N_28839,N_28415,N_28110);
nor U28840 (N_28840,N_28215,N_28196);
or U28841 (N_28841,N_28038,N_28162);
nor U28842 (N_28842,N_28466,N_28492);
nand U28843 (N_28843,N_28355,N_28064);
nand U28844 (N_28844,N_28357,N_28475);
and U28845 (N_28845,N_28071,N_28150);
nand U28846 (N_28846,N_28205,N_28270);
or U28847 (N_28847,N_28491,N_28149);
and U28848 (N_28848,N_28116,N_28473);
nor U28849 (N_28849,N_28352,N_28490);
nand U28850 (N_28850,N_28161,N_28071);
xnor U28851 (N_28851,N_28432,N_28479);
xor U28852 (N_28852,N_28187,N_28410);
and U28853 (N_28853,N_28377,N_28078);
and U28854 (N_28854,N_28161,N_28086);
and U28855 (N_28855,N_28236,N_28336);
or U28856 (N_28856,N_28182,N_28167);
or U28857 (N_28857,N_28417,N_28023);
and U28858 (N_28858,N_28331,N_28065);
nor U28859 (N_28859,N_28428,N_28340);
xnor U28860 (N_28860,N_28226,N_28071);
nor U28861 (N_28861,N_28385,N_28454);
or U28862 (N_28862,N_28284,N_28197);
or U28863 (N_28863,N_28236,N_28387);
xnor U28864 (N_28864,N_28128,N_28005);
xor U28865 (N_28865,N_28041,N_28122);
or U28866 (N_28866,N_28221,N_28140);
or U28867 (N_28867,N_28306,N_28381);
and U28868 (N_28868,N_28253,N_28034);
or U28869 (N_28869,N_28234,N_28139);
nand U28870 (N_28870,N_28300,N_28101);
nand U28871 (N_28871,N_28332,N_28238);
nor U28872 (N_28872,N_28471,N_28241);
or U28873 (N_28873,N_28425,N_28086);
xor U28874 (N_28874,N_28123,N_28250);
or U28875 (N_28875,N_28094,N_28162);
and U28876 (N_28876,N_28089,N_28097);
and U28877 (N_28877,N_28176,N_28067);
and U28878 (N_28878,N_28342,N_28234);
xnor U28879 (N_28879,N_28432,N_28325);
and U28880 (N_28880,N_28356,N_28484);
nor U28881 (N_28881,N_28023,N_28077);
xnor U28882 (N_28882,N_28092,N_28433);
nand U28883 (N_28883,N_28438,N_28450);
nand U28884 (N_28884,N_28249,N_28034);
nor U28885 (N_28885,N_28036,N_28481);
nand U28886 (N_28886,N_28271,N_28367);
or U28887 (N_28887,N_28122,N_28351);
or U28888 (N_28888,N_28174,N_28026);
and U28889 (N_28889,N_28108,N_28453);
nand U28890 (N_28890,N_28032,N_28288);
nor U28891 (N_28891,N_28401,N_28149);
nor U28892 (N_28892,N_28268,N_28294);
nand U28893 (N_28893,N_28312,N_28279);
nand U28894 (N_28894,N_28014,N_28301);
nand U28895 (N_28895,N_28494,N_28263);
or U28896 (N_28896,N_28074,N_28310);
nor U28897 (N_28897,N_28315,N_28318);
or U28898 (N_28898,N_28066,N_28076);
xor U28899 (N_28899,N_28340,N_28095);
xor U28900 (N_28900,N_28202,N_28230);
or U28901 (N_28901,N_28396,N_28393);
nand U28902 (N_28902,N_28105,N_28180);
nand U28903 (N_28903,N_28291,N_28266);
nor U28904 (N_28904,N_28486,N_28193);
or U28905 (N_28905,N_28415,N_28278);
and U28906 (N_28906,N_28475,N_28429);
xnor U28907 (N_28907,N_28322,N_28061);
and U28908 (N_28908,N_28320,N_28416);
or U28909 (N_28909,N_28153,N_28309);
xor U28910 (N_28910,N_28322,N_28293);
and U28911 (N_28911,N_28098,N_28131);
and U28912 (N_28912,N_28218,N_28470);
and U28913 (N_28913,N_28235,N_28207);
or U28914 (N_28914,N_28038,N_28266);
nor U28915 (N_28915,N_28060,N_28192);
nor U28916 (N_28916,N_28080,N_28410);
xor U28917 (N_28917,N_28198,N_28208);
nor U28918 (N_28918,N_28182,N_28093);
nand U28919 (N_28919,N_28168,N_28007);
nor U28920 (N_28920,N_28151,N_28242);
and U28921 (N_28921,N_28385,N_28250);
nor U28922 (N_28922,N_28293,N_28207);
nor U28923 (N_28923,N_28127,N_28257);
nand U28924 (N_28924,N_28042,N_28477);
nand U28925 (N_28925,N_28272,N_28440);
nor U28926 (N_28926,N_28101,N_28310);
or U28927 (N_28927,N_28085,N_28468);
nor U28928 (N_28928,N_28448,N_28330);
or U28929 (N_28929,N_28228,N_28361);
nand U28930 (N_28930,N_28043,N_28145);
nand U28931 (N_28931,N_28489,N_28205);
or U28932 (N_28932,N_28032,N_28282);
nand U28933 (N_28933,N_28173,N_28400);
nor U28934 (N_28934,N_28403,N_28367);
or U28935 (N_28935,N_28482,N_28189);
or U28936 (N_28936,N_28057,N_28283);
or U28937 (N_28937,N_28317,N_28336);
nor U28938 (N_28938,N_28054,N_28397);
nor U28939 (N_28939,N_28128,N_28452);
xnor U28940 (N_28940,N_28493,N_28321);
and U28941 (N_28941,N_28111,N_28017);
nand U28942 (N_28942,N_28345,N_28400);
nand U28943 (N_28943,N_28037,N_28051);
and U28944 (N_28944,N_28290,N_28093);
nand U28945 (N_28945,N_28059,N_28031);
nor U28946 (N_28946,N_28220,N_28175);
or U28947 (N_28947,N_28093,N_28221);
xor U28948 (N_28948,N_28234,N_28265);
or U28949 (N_28949,N_28297,N_28097);
or U28950 (N_28950,N_28331,N_28350);
nor U28951 (N_28951,N_28329,N_28362);
xnor U28952 (N_28952,N_28415,N_28144);
or U28953 (N_28953,N_28173,N_28336);
or U28954 (N_28954,N_28180,N_28264);
and U28955 (N_28955,N_28480,N_28323);
or U28956 (N_28956,N_28289,N_28205);
xnor U28957 (N_28957,N_28442,N_28015);
nand U28958 (N_28958,N_28123,N_28274);
xor U28959 (N_28959,N_28002,N_28369);
xor U28960 (N_28960,N_28061,N_28216);
nor U28961 (N_28961,N_28133,N_28405);
nand U28962 (N_28962,N_28232,N_28378);
and U28963 (N_28963,N_28298,N_28234);
nand U28964 (N_28964,N_28424,N_28385);
or U28965 (N_28965,N_28221,N_28429);
nor U28966 (N_28966,N_28249,N_28301);
or U28967 (N_28967,N_28277,N_28213);
nor U28968 (N_28968,N_28079,N_28199);
and U28969 (N_28969,N_28104,N_28173);
xor U28970 (N_28970,N_28457,N_28335);
nor U28971 (N_28971,N_28134,N_28039);
xnor U28972 (N_28972,N_28140,N_28283);
nand U28973 (N_28973,N_28082,N_28290);
or U28974 (N_28974,N_28229,N_28435);
or U28975 (N_28975,N_28252,N_28267);
xnor U28976 (N_28976,N_28326,N_28309);
nand U28977 (N_28977,N_28088,N_28033);
or U28978 (N_28978,N_28063,N_28255);
or U28979 (N_28979,N_28302,N_28035);
xor U28980 (N_28980,N_28372,N_28095);
and U28981 (N_28981,N_28414,N_28271);
xnor U28982 (N_28982,N_28447,N_28034);
and U28983 (N_28983,N_28061,N_28402);
or U28984 (N_28984,N_28373,N_28119);
and U28985 (N_28985,N_28202,N_28200);
and U28986 (N_28986,N_28160,N_28117);
xor U28987 (N_28987,N_28232,N_28450);
nand U28988 (N_28988,N_28121,N_28068);
xnor U28989 (N_28989,N_28030,N_28290);
and U28990 (N_28990,N_28353,N_28395);
and U28991 (N_28991,N_28342,N_28334);
or U28992 (N_28992,N_28151,N_28114);
nor U28993 (N_28993,N_28414,N_28105);
or U28994 (N_28994,N_28154,N_28029);
or U28995 (N_28995,N_28237,N_28298);
or U28996 (N_28996,N_28387,N_28328);
or U28997 (N_28997,N_28277,N_28158);
nand U28998 (N_28998,N_28466,N_28445);
nor U28999 (N_28999,N_28081,N_28310);
and U29000 (N_29000,N_28939,N_28817);
xor U29001 (N_29001,N_28677,N_28639);
nand U29002 (N_29002,N_28622,N_28883);
nor U29003 (N_29003,N_28847,N_28772);
or U29004 (N_29004,N_28995,N_28523);
or U29005 (N_29005,N_28560,N_28660);
nand U29006 (N_29006,N_28513,N_28792);
nor U29007 (N_29007,N_28666,N_28953);
nand U29008 (N_29008,N_28936,N_28575);
or U29009 (N_29009,N_28608,N_28873);
xor U29010 (N_29010,N_28975,N_28797);
and U29011 (N_29011,N_28828,N_28659);
or U29012 (N_29012,N_28816,N_28906);
nand U29013 (N_29013,N_28534,N_28859);
nand U29014 (N_29014,N_28904,N_28796);
or U29015 (N_29015,N_28991,N_28550);
and U29016 (N_29016,N_28500,N_28960);
nand U29017 (N_29017,N_28759,N_28756);
nor U29018 (N_29018,N_28771,N_28985);
xnor U29019 (N_29019,N_28635,N_28658);
and U29020 (N_29020,N_28938,N_28554);
nor U29021 (N_29021,N_28717,N_28800);
nor U29022 (N_29022,N_28624,N_28602);
nand U29023 (N_29023,N_28930,N_28990);
nand U29024 (N_29024,N_28732,N_28885);
xor U29025 (N_29025,N_28768,N_28919);
nand U29026 (N_29026,N_28581,N_28510);
xnor U29027 (N_29027,N_28740,N_28502);
and U29028 (N_29028,N_28853,N_28739);
nand U29029 (N_29029,N_28887,N_28793);
xor U29030 (N_29030,N_28977,N_28537);
nor U29031 (N_29031,N_28863,N_28506);
nor U29032 (N_29032,N_28629,N_28764);
nand U29033 (N_29033,N_28593,N_28869);
xor U29034 (N_29034,N_28905,N_28997);
xor U29035 (N_29035,N_28533,N_28641);
xnor U29036 (N_29036,N_28579,N_28685);
xor U29037 (N_29037,N_28676,N_28778);
xnor U29038 (N_29038,N_28710,N_28516);
and U29039 (N_29039,N_28728,N_28813);
xor U29040 (N_29040,N_28935,N_28942);
nor U29041 (N_29041,N_28802,N_28561);
nor U29042 (N_29042,N_28595,N_28892);
nand U29043 (N_29043,N_28970,N_28804);
xnor U29044 (N_29044,N_28689,N_28881);
and U29045 (N_29045,N_28604,N_28706);
nor U29046 (N_29046,N_28791,N_28774);
xor U29047 (N_29047,N_28803,N_28769);
and U29048 (N_29048,N_28601,N_28786);
and U29049 (N_29049,N_28741,N_28920);
nand U29050 (N_29050,N_28893,N_28807);
xor U29051 (N_29051,N_28866,N_28648);
xor U29052 (N_29052,N_28783,N_28616);
and U29053 (N_29053,N_28614,N_28707);
or U29054 (N_29054,N_28855,N_28746);
xnor U29055 (N_29055,N_28683,N_28765);
or U29056 (N_29056,N_28999,N_28607);
or U29057 (N_29057,N_28580,N_28625);
or U29058 (N_29058,N_28809,N_28574);
and U29059 (N_29059,N_28949,N_28651);
or U29060 (N_29060,N_28891,N_28757);
nor U29061 (N_29061,N_28679,N_28850);
nor U29062 (N_29062,N_28875,N_28958);
and U29063 (N_29063,N_28914,N_28947);
xnor U29064 (N_29064,N_28543,N_28918);
or U29065 (N_29065,N_28584,N_28838);
and U29066 (N_29066,N_28986,N_28650);
and U29067 (N_29067,N_28599,N_28532);
and U29068 (N_29068,N_28656,N_28943);
xnor U29069 (N_29069,N_28664,N_28631);
nand U29070 (N_29070,N_28940,N_28874);
nand U29071 (N_29071,N_28569,N_28860);
xnor U29072 (N_29072,N_28752,N_28929);
nand U29073 (N_29073,N_28567,N_28557);
and U29074 (N_29074,N_28785,N_28609);
or U29075 (N_29075,N_28908,N_28725);
and U29076 (N_29076,N_28723,N_28606);
or U29077 (N_29077,N_28773,N_28505);
nor U29078 (N_29078,N_28552,N_28672);
xor U29079 (N_29079,N_28825,N_28627);
nor U29080 (N_29080,N_28684,N_28907);
and U29081 (N_29081,N_28979,N_28819);
xor U29082 (N_29082,N_28632,N_28527);
or U29083 (N_29083,N_28889,N_28647);
nand U29084 (N_29084,N_28556,N_28509);
xor U29085 (N_29085,N_28511,N_28966);
and U29086 (N_29086,N_28698,N_28541);
or U29087 (N_29087,N_28652,N_28753);
nor U29088 (N_29088,N_28767,N_28718);
or U29089 (N_29089,N_28520,N_28518);
xnor U29090 (N_29090,N_28758,N_28600);
xnor U29091 (N_29091,N_28959,N_28925);
and U29092 (N_29092,N_28750,N_28515);
xor U29093 (N_29093,N_28784,N_28921);
and U29094 (N_29094,N_28680,N_28815);
or U29095 (N_29095,N_28720,N_28603);
and U29096 (N_29096,N_28643,N_28586);
nand U29097 (N_29097,N_28514,N_28909);
nand U29098 (N_29098,N_28738,N_28626);
or U29099 (N_29099,N_28700,N_28628);
nand U29100 (N_29100,N_28981,N_28727);
xor U29101 (N_29101,N_28691,N_28913);
nor U29102 (N_29102,N_28911,N_28983);
nor U29103 (N_29103,N_28834,N_28638);
or U29104 (N_29104,N_28694,N_28782);
and U29105 (N_29105,N_28553,N_28692);
nand U29106 (N_29106,N_28788,N_28988);
or U29107 (N_29107,N_28577,N_28642);
and U29108 (N_29108,N_28634,N_28870);
xnor U29109 (N_29109,N_28596,N_28971);
nor U29110 (N_29110,N_28693,N_28790);
nand U29111 (N_29111,N_28598,N_28766);
xnor U29112 (N_29112,N_28512,N_28877);
nor U29113 (N_29113,N_28799,N_28974);
nand U29114 (N_29114,N_28952,N_28762);
nor U29115 (N_29115,N_28565,N_28617);
nor U29116 (N_29116,N_28779,N_28538);
nor U29117 (N_29117,N_28888,N_28713);
nor U29118 (N_29118,N_28712,N_28775);
nor U29119 (N_29119,N_28879,N_28837);
or U29120 (N_29120,N_28836,N_28835);
or U29121 (N_29121,N_28501,N_28840);
nand U29122 (N_29122,N_28701,N_28528);
or U29123 (N_29123,N_28865,N_28722);
xnor U29124 (N_29124,N_28618,N_28711);
or U29125 (N_29125,N_28503,N_28868);
and U29126 (N_29126,N_28748,N_28856);
or U29127 (N_29127,N_28989,N_28655);
nand U29128 (N_29128,N_28576,N_28962);
and U29129 (N_29129,N_28902,N_28955);
nor U29130 (N_29130,N_28890,N_28956);
nand U29131 (N_29131,N_28849,N_28841);
or U29132 (N_29132,N_28830,N_28927);
and U29133 (N_29133,N_28968,N_28671);
or U29134 (N_29134,N_28716,N_28547);
nor U29135 (N_29135,N_28668,N_28880);
nor U29136 (N_29136,N_28531,N_28726);
or U29137 (N_29137,N_28996,N_28937);
nor U29138 (N_29138,N_28714,N_28854);
xnor U29139 (N_29139,N_28910,N_28594);
xnor U29140 (N_29140,N_28846,N_28839);
or U29141 (N_29141,N_28781,N_28623);
xor U29142 (N_29142,N_28525,N_28969);
and U29143 (N_29143,N_28667,N_28630);
nor U29144 (N_29144,N_28934,N_28964);
and U29145 (N_29145,N_28916,N_28861);
nand U29146 (N_29146,N_28731,N_28946);
or U29147 (N_29147,N_28735,N_28747);
and U29148 (N_29148,N_28578,N_28653);
nor U29149 (N_29149,N_28640,N_28566);
and U29150 (N_29150,N_28944,N_28844);
nand U29151 (N_29151,N_28941,N_28749);
nor U29152 (N_29152,N_28582,N_28917);
or U29153 (N_29153,N_28583,N_28872);
and U29154 (N_29154,N_28744,N_28924);
and U29155 (N_29155,N_28787,N_28862);
nor U29156 (N_29156,N_28669,N_28522);
or U29157 (N_29157,N_28894,N_28549);
nand U29158 (N_29158,N_28504,N_28998);
or U29159 (N_29159,N_28702,N_28670);
xor U29160 (N_29160,N_28857,N_28555);
or U29161 (N_29161,N_28912,N_28573);
xnor U29162 (N_29162,N_28644,N_28688);
nor U29163 (N_29163,N_28585,N_28589);
or U29164 (N_29164,N_28951,N_28649);
nand U29165 (N_29165,N_28780,N_28524);
xor U29166 (N_29166,N_28755,N_28519);
nor U29167 (N_29167,N_28572,N_28903);
xnor U29168 (N_29168,N_28615,N_28987);
or U29169 (N_29169,N_28878,N_28922);
xor U29170 (N_29170,N_28901,N_28950);
xor U29171 (N_29171,N_28590,N_28886);
and U29172 (N_29172,N_28508,N_28657);
and U29173 (N_29173,N_28882,N_28867);
nand U29174 (N_29174,N_28536,N_28611);
and U29175 (N_29175,N_28697,N_28895);
nor U29176 (N_29176,N_28564,N_28754);
nor U29177 (N_29177,N_28984,N_28810);
and U29178 (N_29178,N_28559,N_28967);
nand U29179 (N_29179,N_28829,N_28737);
nand U29180 (N_29180,N_28570,N_28770);
nor U29181 (N_29181,N_28661,N_28805);
xnor U29182 (N_29182,N_28864,N_28963);
or U29183 (N_29183,N_28571,N_28965);
and U29184 (N_29184,N_28546,N_28529);
and U29185 (N_29185,N_28871,N_28690);
nor U29186 (N_29186,N_28826,N_28621);
nor U29187 (N_29187,N_28898,N_28736);
xnor U29188 (N_29188,N_28948,N_28696);
or U29189 (N_29189,N_28897,N_28612);
nor U29190 (N_29190,N_28645,N_28763);
nand U29191 (N_29191,N_28982,N_28708);
nor U29192 (N_29192,N_28721,N_28923);
or U29193 (N_29193,N_28972,N_28823);
and U29194 (N_29194,N_28681,N_28928);
and U29195 (N_29195,N_28932,N_28654);
nor U29196 (N_29196,N_28695,N_28729);
nor U29197 (N_29197,N_28957,N_28831);
nor U29198 (N_29198,N_28709,N_28703);
nor U29199 (N_29199,N_28821,N_28848);
nand U29200 (N_29200,N_28961,N_28926);
xnor U29201 (N_29201,N_28822,N_28761);
xor U29202 (N_29202,N_28814,N_28899);
and U29203 (N_29203,N_28833,N_28827);
xor U29204 (N_29204,N_28539,N_28687);
and U29205 (N_29205,N_28620,N_28592);
nand U29206 (N_29206,N_28665,N_28544);
nor U29207 (N_29207,N_28824,N_28798);
or U29208 (N_29208,N_28795,N_28682);
nor U29209 (N_29209,N_28705,N_28663);
xnor U29210 (N_29210,N_28801,N_28605);
and U29211 (N_29211,N_28587,N_28777);
or U29212 (N_29212,N_28852,N_28733);
nor U29213 (N_29213,N_28588,N_28678);
and U29214 (N_29214,N_28568,N_28530);
xor U29215 (N_29215,N_28931,N_28884);
nand U29216 (N_29216,N_28808,N_28818);
xnor U29217 (N_29217,N_28760,N_28542);
and U29218 (N_29218,N_28820,N_28562);
or U29219 (N_29219,N_28851,N_28633);
xor U29220 (N_29220,N_28673,N_28954);
or U29221 (N_29221,N_28811,N_28719);
nor U29222 (N_29222,N_28558,N_28876);
nand U29223 (N_29223,N_28535,N_28619);
nand U29224 (N_29224,N_28789,N_28858);
and U29225 (N_29225,N_28545,N_28915);
nand U29226 (N_29226,N_28745,N_28591);
and U29227 (N_29227,N_28900,N_28776);
xor U29228 (N_29228,N_28980,N_28507);
and U29229 (N_29229,N_28976,N_28845);
and U29230 (N_29230,N_28662,N_28734);
nand U29231 (N_29231,N_28548,N_28832);
or U29232 (N_29232,N_28521,N_28610);
and U29233 (N_29233,N_28540,N_28704);
nand U29234 (N_29234,N_28794,N_28674);
or U29235 (N_29235,N_28896,N_28637);
and U29236 (N_29236,N_28751,N_28636);
nor U29237 (N_29237,N_28992,N_28743);
nor U29238 (N_29238,N_28699,N_28742);
or U29239 (N_29239,N_28993,N_28724);
nor U29240 (N_29240,N_28613,N_28675);
and U29241 (N_29241,N_28526,N_28686);
or U29242 (N_29242,N_28843,N_28646);
or U29243 (N_29243,N_28563,N_28812);
nand U29244 (N_29244,N_28973,N_28730);
and U29245 (N_29245,N_28806,N_28715);
nand U29246 (N_29246,N_28842,N_28933);
nand U29247 (N_29247,N_28551,N_28978);
and U29248 (N_29248,N_28994,N_28945);
nand U29249 (N_29249,N_28597,N_28517);
nor U29250 (N_29250,N_28957,N_28628);
nor U29251 (N_29251,N_28789,N_28638);
xnor U29252 (N_29252,N_28933,N_28548);
nand U29253 (N_29253,N_28898,N_28744);
nor U29254 (N_29254,N_28573,N_28626);
nand U29255 (N_29255,N_28634,N_28699);
nand U29256 (N_29256,N_28810,N_28887);
or U29257 (N_29257,N_28908,N_28573);
xnor U29258 (N_29258,N_28560,N_28906);
or U29259 (N_29259,N_28875,N_28688);
xnor U29260 (N_29260,N_28791,N_28631);
and U29261 (N_29261,N_28803,N_28666);
xor U29262 (N_29262,N_28721,N_28898);
or U29263 (N_29263,N_28871,N_28874);
or U29264 (N_29264,N_28572,N_28656);
and U29265 (N_29265,N_28517,N_28509);
nor U29266 (N_29266,N_28655,N_28760);
and U29267 (N_29267,N_28857,N_28504);
nand U29268 (N_29268,N_28719,N_28746);
nor U29269 (N_29269,N_28885,N_28653);
xor U29270 (N_29270,N_28534,N_28780);
nor U29271 (N_29271,N_28956,N_28852);
xor U29272 (N_29272,N_28580,N_28960);
and U29273 (N_29273,N_28693,N_28676);
and U29274 (N_29274,N_28658,N_28897);
and U29275 (N_29275,N_28592,N_28735);
and U29276 (N_29276,N_28779,N_28616);
nor U29277 (N_29277,N_28907,N_28671);
nor U29278 (N_29278,N_28818,N_28582);
xor U29279 (N_29279,N_28878,N_28876);
and U29280 (N_29280,N_28601,N_28814);
or U29281 (N_29281,N_28531,N_28785);
nand U29282 (N_29282,N_28995,N_28583);
nand U29283 (N_29283,N_28604,N_28640);
nand U29284 (N_29284,N_28583,N_28856);
nand U29285 (N_29285,N_28784,N_28838);
nand U29286 (N_29286,N_28603,N_28997);
nand U29287 (N_29287,N_28993,N_28542);
nand U29288 (N_29288,N_28511,N_28733);
nand U29289 (N_29289,N_28757,N_28728);
nand U29290 (N_29290,N_28684,N_28788);
xor U29291 (N_29291,N_28858,N_28658);
or U29292 (N_29292,N_28659,N_28916);
xor U29293 (N_29293,N_28638,N_28615);
nand U29294 (N_29294,N_28697,N_28671);
and U29295 (N_29295,N_28719,N_28707);
nand U29296 (N_29296,N_28515,N_28680);
xor U29297 (N_29297,N_28869,N_28846);
xor U29298 (N_29298,N_28781,N_28799);
nand U29299 (N_29299,N_28683,N_28863);
nor U29300 (N_29300,N_28888,N_28777);
or U29301 (N_29301,N_28619,N_28741);
and U29302 (N_29302,N_28779,N_28727);
or U29303 (N_29303,N_28625,N_28683);
and U29304 (N_29304,N_28651,N_28883);
or U29305 (N_29305,N_28806,N_28854);
and U29306 (N_29306,N_28525,N_28751);
nand U29307 (N_29307,N_28818,N_28819);
nor U29308 (N_29308,N_28996,N_28733);
nor U29309 (N_29309,N_28755,N_28751);
xor U29310 (N_29310,N_28705,N_28743);
nor U29311 (N_29311,N_28691,N_28711);
nor U29312 (N_29312,N_28744,N_28822);
nor U29313 (N_29313,N_28913,N_28584);
and U29314 (N_29314,N_28567,N_28704);
nor U29315 (N_29315,N_28956,N_28591);
nand U29316 (N_29316,N_28757,N_28617);
nand U29317 (N_29317,N_28781,N_28529);
xnor U29318 (N_29318,N_28687,N_28985);
and U29319 (N_29319,N_28593,N_28951);
and U29320 (N_29320,N_28583,N_28878);
nor U29321 (N_29321,N_28859,N_28802);
or U29322 (N_29322,N_28567,N_28867);
nor U29323 (N_29323,N_28816,N_28718);
or U29324 (N_29324,N_28709,N_28887);
xor U29325 (N_29325,N_28886,N_28509);
or U29326 (N_29326,N_28690,N_28809);
nor U29327 (N_29327,N_28727,N_28987);
and U29328 (N_29328,N_28540,N_28806);
or U29329 (N_29329,N_28706,N_28753);
nor U29330 (N_29330,N_28513,N_28994);
nor U29331 (N_29331,N_28759,N_28753);
nor U29332 (N_29332,N_28981,N_28700);
or U29333 (N_29333,N_28912,N_28848);
xor U29334 (N_29334,N_28933,N_28705);
nand U29335 (N_29335,N_28662,N_28810);
or U29336 (N_29336,N_28794,N_28541);
or U29337 (N_29337,N_28907,N_28753);
nor U29338 (N_29338,N_28737,N_28551);
or U29339 (N_29339,N_28510,N_28683);
nand U29340 (N_29340,N_28921,N_28802);
nand U29341 (N_29341,N_28909,N_28713);
xor U29342 (N_29342,N_28937,N_28609);
nor U29343 (N_29343,N_28606,N_28622);
and U29344 (N_29344,N_28914,N_28761);
and U29345 (N_29345,N_28967,N_28768);
nand U29346 (N_29346,N_28667,N_28632);
nor U29347 (N_29347,N_28895,N_28955);
xnor U29348 (N_29348,N_28620,N_28845);
xor U29349 (N_29349,N_28619,N_28987);
and U29350 (N_29350,N_28968,N_28879);
nand U29351 (N_29351,N_28698,N_28971);
xor U29352 (N_29352,N_28924,N_28682);
nand U29353 (N_29353,N_28663,N_28642);
and U29354 (N_29354,N_28939,N_28673);
nor U29355 (N_29355,N_28821,N_28669);
nand U29356 (N_29356,N_28785,N_28677);
and U29357 (N_29357,N_28892,N_28739);
xnor U29358 (N_29358,N_28567,N_28814);
or U29359 (N_29359,N_28688,N_28929);
or U29360 (N_29360,N_28506,N_28831);
or U29361 (N_29361,N_28876,N_28858);
nand U29362 (N_29362,N_28721,N_28970);
or U29363 (N_29363,N_28971,N_28741);
and U29364 (N_29364,N_28992,N_28768);
nand U29365 (N_29365,N_28840,N_28698);
or U29366 (N_29366,N_28875,N_28600);
nor U29367 (N_29367,N_28979,N_28647);
nor U29368 (N_29368,N_28845,N_28502);
and U29369 (N_29369,N_28741,N_28702);
nor U29370 (N_29370,N_28817,N_28502);
xnor U29371 (N_29371,N_28954,N_28689);
xor U29372 (N_29372,N_28503,N_28757);
or U29373 (N_29373,N_28967,N_28596);
and U29374 (N_29374,N_28781,N_28633);
nand U29375 (N_29375,N_28871,N_28542);
nor U29376 (N_29376,N_28874,N_28795);
xnor U29377 (N_29377,N_28725,N_28901);
nor U29378 (N_29378,N_28959,N_28625);
or U29379 (N_29379,N_28764,N_28547);
and U29380 (N_29380,N_28932,N_28766);
xnor U29381 (N_29381,N_28779,N_28679);
or U29382 (N_29382,N_28628,N_28540);
nor U29383 (N_29383,N_28964,N_28618);
xnor U29384 (N_29384,N_28577,N_28505);
xor U29385 (N_29385,N_28934,N_28630);
xor U29386 (N_29386,N_28701,N_28713);
xor U29387 (N_29387,N_28524,N_28890);
nand U29388 (N_29388,N_28640,N_28775);
nand U29389 (N_29389,N_28670,N_28858);
nand U29390 (N_29390,N_28836,N_28846);
and U29391 (N_29391,N_28680,N_28647);
or U29392 (N_29392,N_28835,N_28697);
xor U29393 (N_29393,N_28989,N_28516);
xnor U29394 (N_29394,N_28575,N_28635);
nor U29395 (N_29395,N_28757,N_28711);
and U29396 (N_29396,N_28666,N_28508);
xor U29397 (N_29397,N_28643,N_28844);
xnor U29398 (N_29398,N_28890,N_28602);
nor U29399 (N_29399,N_28677,N_28908);
nand U29400 (N_29400,N_28966,N_28845);
nor U29401 (N_29401,N_28869,N_28942);
and U29402 (N_29402,N_28866,N_28707);
nor U29403 (N_29403,N_28592,N_28773);
or U29404 (N_29404,N_28932,N_28572);
and U29405 (N_29405,N_28898,N_28895);
and U29406 (N_29406,N_28784,N_28855);
and U29407 (N_29407,N_28977,N_28708);
nor U29408 (N_29408,N_28513,N_28738);
nor U29409 (N_29409,N_28904,N_28636);
or U29410 (N_29410,N_28942,N_28696);
and U29411 (N_29411,N_28955,N_28711);
or U29412 (N_29412,N_28916,N_28910);
or U29413 (N_29413,N_28875,N_28739);
or U29414 (N_29414,N_28921,N_28929);
or U29415 (N_29415,N_28517,N_28759);
xnor U29416 (N_29416,N_28522,N_28897);
nand U29417 (N_29417,N_28824,N_28595);
xor U29418 (N_29418,N_28582,N_28919);
nand U29419 (N_29419,N_28965,N_28711);
xnor U29420 (N_29420,N_28979,N_28586);
or U29421 (N_29421,N_28948,N_28725);
nand U29422 (N_29422,N_28755,N_28773);
nand U29423 (N_29423,N_28849,N_28884);
nor U29424 (N_29424,N_28630,N_28977);
nand U29425 (N_29425,N_28916,N_28758);
or U29426 (N_29426,N_28948,N_28665);
nor U29427 (N_29427,N_28892,N_28714);
nor U29428 (N_29428,N_28525,N_28581);
or U29429 (N_29429,N_28993,N_28741);
nor U29430 (N_29430,N_28739,N_28763);
nor U29431 (N_29431,N_28770,N_28789);
xor U29432 (N_29432,N_28555,N_28728);
and U29433 (N_29433,N_28534,N_28681);
or U29434 (N_29434,N_28663,N_28926);
xor U29435 (N_29435,N_28689,N_28508);
xor U29436 (N_29436,N_28546,N_28985);
or U29437 (N_29437,N_28852,N_28595);
and U29438 (N_29438,N_28639,N_28534);
nor U29439 (N_29439,N_28837,N_28997);
or U29440 (N_29440,N_28891,N_28614);
nand U29441 (N_29441,N_28782,N_28607);
and U29442 (N_29442,N_28779,N_28656);
nor U29443 (N_29443,N_28556,N_28933);
and U29444 (N_29444,N_28517,N_28827);
and U29445 (N_29445,N_28611,N_28838);
and U29446 (N_29446,N_28993,N_28630);
or U29447 (N_29447,N_28648,N_28616);
nor U29448 (N_29448,N_28519,N_28774);
and U29449 (N_29449,N_28626,N_28846);
or U29450 (N_29450,N_28950,N_28815);
or U29451 (N_29451,N_28553,N_28564);
or U29452 (N_29452,N_28655,N_28778);
xnor U29453 (N_29453,N_28662,N_28908);
nand U29454 (N_29454,N_28934,N_28872);
xor U29455 (N_29455,N_28998,N_28542);
nor U29456 (N_29456,N_28571,N_28778);
nor U29457 (N_29457,N_28974,N_28672);
and U29458 (N_29458,N_28816,N_28934);
nor U29459 (N_29459,N_28743,N_28802);
and U29460 (N_29460,N_28553,N_28945);
or U29461 (N_29461,N_28860,N_28639);
or U29462 (N_29462,N_28884,N_28638);
or U29463 (N_29463,N_28937,N_28781);
nor U29464 (N_29464,N_28613,N_28845);
and U29465 (N_29465,N_28604,N_28611);
or U29466 (N_29466,N_28708,N_28707);
and U29467 (N_29467,N_28631,N_28952);
xnor U29468 (N_29468,N_28862,N_28573);
nand U29469 (N_29469,N_28796,N_28638);
and U29470 (N_29470,N_28637,N_28798);
or U29471 (N_29471,N_28954,N_28577);
nand U29472 (N_29472,N_28615,N_28776);
or U29473 (N_29473,N_28879,N_28806);
or U29474 (N_29474,N_28535,N_28646);
and U29475 (N_29475,N_28600,N_28953);
nor U29476 (N_29476,N_28608,N_28613);
nor U29477 (N_29477,N_28851,N_28998);
xnor U29478 (N_29478,N_28914,N_28529);
nor U29479 (N_29479,N_28914,N_28666);
xnor U29480 (N_29480,N_28957,N_28734);
xor U29481 (N_29481,N_28702,N_28593);
and U29482 (N_29482,N_28970,N_28794);
or U29483 (N_29483,N_28867,N_28538);
nand U29484 (N_29484,N_28738,N_28530);
nand U29485 (N_29485,N_28987,N_28553);
nand U29486 (N_29486,N_28971,N_28813);
and U29487 (N_29487,N_28641,N_28772);
and U29488 (N_29488,N_28841,N_28902);
and U29489 (N_29489,N_28894,N_28763);
nor U29490 (N_29490,N_28613,N_28703);
and U29491 (N_29491,N_28994,N_28596);
xor U29492 (N_29492,N_28605,N_28563);
or U29493 (N_29493,N_28809,N_28661);
and U29494 (N_29494,N_28567,N_28681);
xnor U29495 (N_29495,N_28597,N_28594);
xor U29496 (N_29496,N_28572,N_28813);
and U29497 (N_29497,N_28593,N_28824);
nand U29498 (N_29498,N_28725,N_28605);
nor U29499 (N_29499,N_28633,N_28763);
nor U29500 (N_29500,N_29251,N_29492);
xor U29501 (N_29501,N_29051,N_29041);
nand U29502 (N_29502,N_29203,N_29100);
and U29503 (N_29503,N_29088,N_29068);
xnor U29504 (N_29504,N_29480,N_29071);
nand U29505 (N_29505,N_29336,N_29128);
nor U29506 (N_29506,N_29406,N_29187);
xor U29507 (N_29507,N_29049,N_29377);
and U29508 (N_29508,N_29477,N_29101);
and U29509 (N_29509,N_29345,N_29257);
and U29510 (N_29510,N_29276,N_29390);
xnor U29511 (N_29511,N_29025,N_29389);
xor U29512 (N_29512,N_29288,N_29451);
or U29513 (N_29513,N_29287,N_29226);
nor U29514 (N_29514,N_29077,N_29214);
nand U29515 (N_29515,N_29436,N_29489);
nor U29516 (N_29516,N_29289,N_29125);
nor U29517 (N_29517,N_29338,N_29168);
or U29518 (N_29518,N_29391,N_29471);
xor U29519 (N_29519,N_29475,N_29484);
xnor U29520 (N_29520,N_29096,N_29347);
and U29521 (N_29521,N_29372,N_29178);
xor U29522 (N_29522,N_29173,N_29367);
nand U29523 (N_29523,N_29221,N_29322);
and U29524 (N_29524,N_29274,N_29196);
or U29525 (N_29525,N_29036,N_29004);
nand U29526 (N_29526,N_29405,N_29424);
nand U29527 (N_29527,N_29319,N_29415);
nor U29528 (N_29528,N_29079,N_29121);
nand U29529 (N_29529,N_29120,N_29481);
or U29530 (N_29530,N_29335,N_29235);
nand U29531 (N_29531,N_29151,N_29264);
nand U29532 (N_29532,N_29123,N_29150);
or U29533 (N_29533,N_29225,N_29430);
xnor U29534 (N_29534,N_29198,N_29202);
xor U29535 (N_29535,N_29425,N_29465);
xor U29536 (N_29536,N_29144,N_29247);
xor U29537 (N_29537,N_29158,N_29464);
nor U29538 (N_29538,N_29435,N_29427);
nor U29539 (N_29539,N_29447,N_29473);
or U29540 (N_29540,N_29182,N_29195);
xnor U29541 (N_29541,N_29472,N_29478);
xor U29542 (N_29542,N_29369,N_29012);
or U29543 (N_29543,N_29070,N_29174);
xor U29544 (N_29544,N_29352,N_29163);
and U29545 (N_29545,N_29343,N_29154);
and U29546 (N_29546,N_29236,N_29212);
nand U29547 (N_29547,N_29375,N_29364);
xnor U29548 (N_29548,N_29140,N_29082);
and U29549 (N_29549,N_29024,N_29393);
and U29550 (N_29550,N_29252,N_29362);
xor U29551 (N_29551,N_29126,N_29292);
nor U29552 (N_29552,N_29245,N_29324);
nor U29553 (N_29553,N_29038,N_29043);
nand U29554 (N_29554,N_29035,N_29115);
or U29555 (N_29555,N_29142,N_29205);
xor U29556 (N_29556,N_29180,N_29099);
xor U29557 (N_29557,N_29317,N_29003);
or U29558 (N_29558,N_29186,N_29269);
and U29559 (N_29559,N_29355,N_29404);
xnor U29560 (N_29560,N_29408,N_29055);
and U29561 (N_29561,N_29046,N_29016);
or U29562 (N_29562,N_29417,N_29366);
or U29563 (N_29563,N_29299,N_29078);
or U29564 (N_29564,N_29438,N_29348);
and U29565 (N_29565,N_29179,N_29122);
nor U29566 (N_29566,N_29382,N_29013);
or U29567 (N_29567,N_29111,N_29273);
or U29568 (N_29568,N_29105,N_29048);
xor U29569 (N_29569,N_29431,N_29392);
and U29570 (N_29570,N_29363,N_29297);
and U29571 (N_29571,N_29442,N_29482);
xor U29572 (N_29572,N_29201,N_29228);
or U29573 (N_29573,N_29074,N_29230);
nand U29574 (N_29574,N_29190,N_29107);
xor U29575 (N_29575,N_29119,N_29192);
nor U29576 (N_29576,N_29194,N_29238);
and U29577 (N_29577,N_29490,N_29114);
or U29578 (N_29578,N_29085,N_29279);
nand U29579 (N_29579,N_29374,N_29353);
and U29580 (N_29580,N_29239,N_29081);
xnor U29581 (N_29581,N_29255,N_29161);
xor U29582 (N_29582,N_29327,N_29056);
xor U29583 (N_29583,N_29401,N_29380);
and U29584 (N_29584,N_29095,N_29023);
or U29585 (N_29585,N_29090,N_29193);
and U29586 (N_29586,N_29127,N_29330);
and U29587 (N_29587,N_29429,N_29488);
or U29588 (N_29588,N_29265,N_29331);
or U29589 (N_29589,N_29084,N_29396);
nand U29590 (N_29590,N_29460,N_29141);
nand U29591 (N_29591,N_29479,N_29103);
or U29592 (N_29592,N_29321,N_29307);
nand U29593 (N_29593,N_29493,N_29091);
nand U29594 (N_29594,N_29277,N_29086);
xor U29595 (N_29595,N_29376,N_29446);
or U29596 (N_29596,N_29223,N_29145);
nor U29597 (N_29597,N_29157,N_29263);
xor U29598 (N_29598,N_29188,N_29044);
xnor U29599 (N_29599,N_29286,N_29208);
nor U29600 (N_29600,N_29244,N_29346);
nor U29601 (N_29601,N_29108,N_29116);
nor U29602 (N_29602,N_29132,N_29009);
or U29603 (N_29603,N_29165,N_29207);
nor U29604 (N_29604,N_29309,N_29253);
nand U29605 (N_29605,N_29052,N_29206);
and U29606 (N_29606,N_29155,N_29370);
nor U29607 (N_29607,N_29216,N_29166);
nor U29608 (N_29608,N_29267,N_29323);
nor U29609 (N_29609,N_29296,N_29341);
xor U29610 (N_29610,N_29298,N_29386);
or U29611 (N_29611,N_29177,N_29006);
nand U29612 (N_29612,N_29170,N_29320);
and U29613 (N_29613,N_29470,N_29314);
nor U29614 (N_29614,N_29219,N_29499);
and U29615 (N_29615,N_29448,N_29227);
nand U29616 (N_29616,N_29350,N_29093);
nor U29617 (N_29617,N_29397,N_29066);
nor U29618 (N_29618,N_29444,N_29373);
and U29619 (N_29619,N_29418,N_29266);
nor U29620 (N_29620,N_29129,N_29109);
nand U29621 (N_29621,N_29410,N_29359);
or U29622 (N_29622,N_29017,N_29419);
or U29623 (N_29623,N_29452,N_29434);
or U29624 (N_29624,N_29215,N_29001);
or U29625 (N_29625,N_29342,N_29468);
or U29626 (N_29626,N_29243,N_29304);
nor U29627 (N_29627,N_29360,N_29268);
or U29628 (N_29628,N_29050,N_29047);
nand U29629 (N_29629,N_29199,N_29262);
and U29630 (N_29630,N_29498,N_29291);
xor U29631 (N_29631,N_29010,N_29420);
nand U29632 (N_29632,N_29184,N_29474);
xnor U29633 (N_29633,N_29029,N_29211);
nand U29634 (N_29634,N_29104,N_29260);
or U29635 (N_29635,N_29034,N_29486);
nor U29636 (N_29636,N_29261,N_29285);
or U29637 (N_29637,N_29136,N_29409);
xor U29638 (N_29638,N_29011,N_29306);
or U29639 (N_29639,N_29130,N_29224);
xor U29640 (N_29640,N_29428,N_29463);
nand U29641 (N_29641,N_29258,N_29027);
nor U29642 (N_29642,N_29169,N_29124);
nand U29643 (N_29643,N_29094,N_29149);
and U29644 (N_29644,N_29270,N_29250);
xor U29645 (N_29645,N_29491,N_29313);
nand U29646 (N_29646,N_29028,N_29275);
nor U29647 (N_29647,N_29329,N_29148);
nand U29648 (N_29648,N_29371,N_29057);
nand U29649 (N_29649,N_29040,N_29295);
and U29650 (N_29650,N_29432,N_29459);
xor U29651 (N_29651,N_29118,N_29183);
xnor U29652 (N_29652,N_29272,N_29361);
or U29653 (N_29653,N_29117,N_29171);
nand U29654 (N_29654,N_29018,N_29290);
or U29655 (N_29655,N_29333,N_29349);
nand U29656 (N_29656,N_29421,N_29433);
and U29657 (N_29657,N_29422,N_29497);
nor U29658 (N_29658,N_29368,N_29200);
or U29659 (N_29659,N_29411,N_29053);
nand U29660 (N_29660,N_29007,N_29450);
nand U29661 (N_29661,N_29063,N_29485);
nor U29662 (N_29662,N_29106,N_29426);
nand U29663 (N_29663,N_29249,N_29097);
xnor U29664 (N_29664,N_29339,N_29153);
nor U29665 (N_29665,N_29241,N_29080);
and U29666 (N_29666,N_29256,N_29033);
xnor U29667 (N_29667,N_29072,N_29102);
nor U29668 (N_29668,N_29358,N_29032);
nor U29669 (N_29669,N_29476,N_29354);
and U29670 (N_29670,N_29381,N_29412);
xor U29671 (N_29671,N_29000,N_29437);
nand U29672 (N_29672,N_29454,N_29385);
nand U29673 (N_29673,N_29042,N_29030);
or U29674 (N_29674,N_29164,N_29064);
nor U29675 (N_29675,N_29316,N_29305);
or U29676 (N_29676,N_29445,N_29059);
xor U29677 (N_29677,N_29416,N_29462);
and U29678 (N_29678,N_29020,N_29311);
or U29679 (N_29679,N_29449,N_29162);
or U29680 (N_29680,N_29387,N_29232);
and U29681 (N_29681,N_29443,N_29087);
nor U29682 (N_29682,N_29402,N_29259);
or U29683 (N_29683,N_29334,N_29014);
and U29684 (N_29684,N_29407,N_29423);
and U29685 (N_29685,N_29278,N_29152);
or U29686 (N_29686,N_29282,N_29039);
and U29687 (N_29687,N_29204,N_29133);
or U29688 (N_29688,N_29308,N_29209);
and U29689 (N_29689,N_29318,N_29351);
xor U29690 (N_29690,N_29483,N_29234);
xnor U29691 (N_29691,N_29189,N_29487);
and U29692 (N_29692,N_29167,N_29237);
nand U29693 (N_29693,N_29399,N_29388);
xor U29694 (N_29694,N_29379,N_29015);
nor U29695 (N_29695,N_29332,N_29495);
nor U29696 (N_29696,N_29466,N_29089);
xnor U29697 (N_29697,N_29344,N_29469);
nand U29698 (N_29698,N_29293,N_29312);
or U29699 (N_29699,N_29175,N_29054);
nand U29700 (N_29700,N_29283,N_29340);
and U29701 (N_29701,N_29008,N_29139);
xor U29702 (N_29702,N_29176,N_29172);
or U29703 (N_29703,N_29229,N_29233);
xnor U29704 (N_29704,N_29031,N_29284);
or U29705 (N_29705,N_29138,N_29280);
and U29706 (N_29706,N_29328,N_29067);
nor U29707 (N_29707,N_29400,N_29073);
nand U29708 (N_29708,N_29453,N_29062);
nand U29709 (N_29709,N_29156,N_29456);
or U29710 (N_29710,N_29113,N_29076);
or U29711 (N_29711,N_29461,N_29383);
nor U29712 (N_29712,N_29378,N_29271);
and U29713 (N_29713,N_29137,N_29026);
xor U29714 (N_29714,N_29160,N_29135);
xnor U29715 (N_29715,N_29110,N_29458);
nor U29716 (N_29716,N_29143,N_29315);
or U29717 (N_29717,N_29069,N_29467);
nand U29718 (N_29718,N_29065,N_29414);
nand U29719 (N_29719,N_29440,N_29058);
nand U29720 (N_29720,N_29197,N_29098);
nor U29721 (N_29721,N_29441,N_29356);
nor U29722 (N_29722,N_29002,N_29455);
nor U29723 (N_29723,N_29281,N_29092);
nand U29724 (N_29724,N_29303,N_29384);
or U29725 (N_29725,N_29217,N_29147);
nor U29726 (N_29726,N_29019,N_29301);
and U29727 (N_29727,N_29248,N_29185);
nor U29728 (N_29728,N_29146,N_29398);
nand U29729 (N_29729,N_29496,N_29022);
and U29730 (N_29730,N_29357,N_29310);
nand U29731 (N_29731,N_29045,N_29302);
xnor U29732 (N_29732,N_29365,N_29294);
or U29733 (N_29733,N_29075,N_29326);
and U29734 (N_29734,N_29134,N_29246);
or U29735 (N_29735,N_29325,N_29060);
nor U29736 (N_29736,N_29254,N_29213);
xor U29737 (N_29737,N_29005,N_29112);
nor U29738 (N_29738,N_29403,N_29337);
xor U29739 (N_29739,N_29131,N_29159);
nand U29740 (N_29740,N_29037,N_29181);
xnor U29741 (N_29741,N_29457,N_29191);
nand U29742 (N_29742,N_29300,N_29021);
and U29743 (N_29743,N_29220,N_29395);
nor U29744 (N_29744,N_29210,N_29222);
xnor U29745 (N_29745,N_29242,N_29231);
and U29746 (N_29746,N_29439,N_29494);
xnor U29747 (N_29747,N_29218,N_29061);
nor U29748 (N_29748,N_29413,N_29083);
and U29749 (N_29749,N_29240,N_29394);
and U29750 (N_29750,N_29064,N_29106);
or U29751 (N_29751,N_29372,N_29297);
nor U29752 (N_29752,N_29395,N_29475);
or U29753 (N_29753,N_29071,N_29387);
nor U29754 (N_29754,N_29141,N_29474);
xor U29755 (N_29755,N_29384,N_29213);
nand U29756 (N_29756,N_29448,N_29179);
nor U29757 (N_29757,N_29087,N_29036);
nand U29758 (N_29758,N_29387,N_29441);
or U29759 (N_29759,N_29192,N_29109);
xor U29760 (N_29760,N_29131,N_29312);
xor U29761 (N_29761,N_29072,N_29139);
nand U29762 (N_29762,N_29086,N_29122);
or U29763 (N_29763,N_29091,N_29322);
nor U29764 (N_29764,N_29386,N_29191);
nand U29765 (N_29765,N_29310,N_29359);
or U29766 (N_29766,N_29483,N_29206);
and U29767 (N_29767,N_29147,N_29398);
nor U29768 (N_29768,N_29226,N_29265);
xnor U29769 (N_29769,N_29019,N_29416);
nor U29770 (N_29770,N_29239,N_29187);
or U29771 (N_29771,N_29161,N_29091);
and U29772 (N_29772,N_29252,N_29462);
or U29773 (N_29773,N_29489,N_29367);
and U29774 (N_29774,N_29423,N_29244);
nor U29775 (N_29775,N_29010,N_29474);
nand U29776 (N_29776,N_29484,N_29067);
nand U29777 (N_29777,N_29111,N_29445);
nand U29778 (N_29778,N_29032,N_29282);
nand U29779 (N_29779,N_29163,N_29307);
nor U29780 (N_29780,N_29193,N_29297);
xor U29781 (N_29781,N_29324,N_29096);
nand U29782 (N_29782,N_29408,N_29143);
and U29783 (N_29783,N_29029,N_29254);
xor U29784 (N_29784,N_29162,N_29165);
nand U29785 (N_29785,N_29453,N_29113);
nor U29786 (N_29786,N_29456,N_29179);
xnor U29787 (N_29787,N_29064,N_29444);
nor U29788 (N_29788,N_29077,N_29092);
or U29789 (N_29789,N_29096,N_29184);
nand U29790 (N_29790,N_29276,N_29354);
nor U29791 (N_29791,N_29213,N_29000);
and U29792 (N_29792,N_29478,N_29315);
or U29793 (N_29793,N_29495,N_29473);
or U29794 (N_29794,N_29452,N_29247);
or U29795 (N_29795,N_29118,N_29496);
xnor U29796 (N_29796,N_29280,N_29483);
nor U29797 (N_29797,N_29056,N_29143);
or U29798 (N_29798,N_29390,N_29007);
and U29799 (N_29799,N_29023,N_29370);
and U29800 (N_29800,N_29271,N_29285);
nand U29801 (N_29801,N_29097,N_29054);
xnor U29802 (N_29802,N_29418,N_29389);
or U29803 (N_29803,N_29124,N_29092);
nor U29804 (N_29804,N_29368,N_29242);
and U29805 (N_29805,N_29227,N_29483);
nand U29806 (N_29806,N_29433,N_29427);
or U29807 (N_29807,N_29198,N_29295);
xor U29808 (N_29808,N_29151,N_29387);
nor U29809 (N_29809,N_29423,N_29105);
xnor U29810 (N_29810,N_29427,N_29004);
and U29811 (N_29811,N_29376,N_29410);
xor U29812 (N_29812,N_29102,N_29220);
nor U29813 (N_29813,N_29019,N_29041);
nand U29814 (N_29814,N_29144,N_29255);
and U29815 (N_29815,N_29267,N_29413);
or U29816 (N_29816,N_29193,N_29162);
or U29817 (N_29817,N_29400,N_29150);
nor U29818 (N_29818,N_29035,N_29332);
xnor U29819 (N_29819,N_29251,N_29072);
nand U29820 (N_29820,N_29459,N_29423);
or U29821 (N_29821,N_29126,N_29495);
and U29822 (N_29822,N_29449,N_29098);
and U29823 (N_29823,N_29411,N_29454);
nor U29824 (N_29824,N_29379,N_29169);
xnor U29825 (N_29825,N_29407,N_29042);
and U29826 (N_29826,N_29384,N_29465);
xor U29827 (N_29827,N_29272,N_29336);
or U29828 (N_29828,N_29014,N_29070);
and U29829 (N_29829,N_29305,N_29065);
or U29830 (N_29830,N_29128,N_29117);
xor U29831 (N_29831,N_29106,N_29422);
and U29832 (N_29832,N_29190,N_29365);
nor U29833 (N_29833,N_29209,N_29238);
nor U29834 (N_29834,N_29141,N_29050);
nor U29835 (N_29835,N_29070,N_29065);
xnor U29836 (N_29836,N_29499,N_29238);
nand U29837 (N_29837,N_29239,N_29481);
and U29838 (N_29838,N_29426,N_29018);
xnor U29839 (N_29839,N_29271,N_29477);
and U29840 (N_29840,N_29032,N_29034);
and U29841 (N_29841,N_29238,N_29072);
or U29842 (N_29842,N_29170,N_29487);
and U29843 (N_29843,N_29041,N_29255);
and U29844 (N_29844,N_29423,N_29483);
xor U29845 (N_29845,N_29036,N_29476);
xor U29846 (N_29846,N_29068,N_29428);
nand U29847 (N_29847,N_29102,N_29224);
nand U29848 (N_29848,N_29271,N_29192);
nor U29849 (N_29849,N_29148,N_29386);
and U29850 (N_29850,N_29444,N_29255);
and U29851 (N_29851,N_29490,N_29160);
nor U29852 (N_29852,N_29253,N_29063);
xor U29853 (N_29853,N_29358,N_29397);
xor U29854 (N_29854,N_29146,N_29332);
nand U29855 (N_29855,N_29163,N_29312);
or U29856 (N_29856,N_29385,N_29140);
or U29857 (N_29857,N_29204,N_29107);
nor U29858 (N_29858,N_29405,N_29170);
xnor U29859 (N_29859,N_29111,N_29033);
nand U29860 (N_29860,N_29172,N_29285);
nor U29861 (N_29861,N_29085,N_29282);
nand U29862 (N_29862,N_29439,N_29067);
nor U29863 (N_29863,N_29149,N_29244);
xnor U29864 (N_29864,N_29128,N_29080);
xor U29865 (N_29865,N_29133,N_29028);
nand U29866 (N_29866,N_29139,N_29352);
and U29867 (N_29867,N_29438,N_29089);
nor U29868 (N_29868,N_29331,N_29419);
and U29869 (N_29869,N_29435,N_29279);
nor U29870 (N_29870,N_29164,N_29406);
nand U29871 (N_29871,N_29397,N_29115);
nor U29872 (N_29872,N_29095,N_29477);
or U29873 (N_29873,N_29310,N_29062);
nand U29874 (N_29874,N_29486,N_29050);
nor U29875 (N_29875,N_29444,N_29253);
or U29876 (N_29876,N_29244,N_29402);
nor U29877 (N_29877,N_29098,N_29195);
nor U29878 (N_29878,N_29374,N_29434);
nand U29879 (N_29879,N_29275,N_29235);
or U29880 (N_29880,N_29224,N_29006);
nor U29881 (N_29881,N_29279,N_29370);
nor U29882 (N_29882,N_29241,N_29205);
nor U29883 (N_29883,N_29451,N_29192);
and U29884 (N_29884,N_29488,N_29451);
or U29885 (N_29885,N_29196,N_29024);
nand U29886 (N_29886,N_29147,N_29118);
and U29887 (N_29887,N_29166,N_29014);
or U29888 (N_29888,N_29061,N_29164);
or U29889 (N_29889,N_29350,N_29122);
and U29890 (N_29890,N_29426,N_29458);
nand U29891 (N_29891,N_29382,N_29412);
and U29892 (N_29892,N_29399,N_29319);
nor U29893 (N_29893,N_29170,N_29294);
nor U29894 (N_29894,N_29048,N_29067);
or U29895 (N_29895,N_29425,N_29012);
nand U29896 (N_29896,N_29394,N_29172);
nand U29897 (N_29897,N_29486,N_29247);
or U29898 (N_29898,N_29284,N_29144);
nand U29899 (N_29899,N_29109,N_29173);
nor U29900 (N_29900,N_29276,N_29174);
and U29901 (N_29901,N_29408,N_29037);
xor U29902 (N_29902,N_29477,N_29239);
and U29903 (N_29903,N_29152,N_29331);
or U29904 (N_29904,N_29319,N_29141);
or U29905 (N_29905,N_29129,N_29215);
nand U29906 (N_29906,N_29340,N_29038);
nand U29907 (N_29907,N_29469,N_29225);
xor U29908 (N_29908,N_29442,N_29336);
and U29909 (N_29909,N_29302,N_29125);
nor U29910 (N_29910,N_29288,N_29315);
nand U29911 (N_29911,N_29053,N_29269);
xnor U29912 (N_29912,N_29403,N_29330);
nor U29913 (N_29913,N_29102,N_29355);
xor U29914 (N_29914,N_29475,N_29275);
xor U29915 (N_29915,N_29198,N_29234);
or U29916 (N_29916,N_29172,N_29236);
xor U29917 (N_29917,N_29289,N_29303);
xor U29918 (N_29918,N_29246,N_29236);
or U29919 (N_29919,N_29411,N_29398);
and U29920 (N_29920,N_29068,N_29411);
and U29921 (N_29921,N_29492,N_29143);
or U29922 (N_29922,N_29058,N_29329);
and U29923 (N_29923,N_29213,N_29118);
or U29924 (N_29924,N_29386,N_29235);
xor U29925 (N_29925,N_29456,N_29039);
or U29926 (N_29926,N_29148,N_29433);
nand U29927 (N_29927,N_29357,N_29319);
nor U29928 (N_29928,N_29318,N_29257);
or U29929 (N_29929,N_29113,N_29269);
or U29930 (N_29930,N_29315,N_29312);
nand U29931 (N_29931,N_29195,N_29261);
nor U29932 (N_29932,N_29311,N_29164);
nand U29933 (N_29933,N_29102,N_29426);
or U29934 (N_29934,N_29206,N_29045);
or U29935 (N_29935,N_29451,N_29026);
or U29936 (N_29936,N_29185,N_29246);
xor U29937 (N_29937,N_29186,N_29333);
nor U29938 (N_29938,N_29312,N_29310);
nand U29939 (N_29939,N_29301,N_29322);
xnor U29940 (N_29940,N_29457,N_29158);
and U29941 (N_29941,N_29002,N_29427);
nor U29942 (N_29942,N_29055,N_29223);
or U29943 (N_29943,N_29475,N_29410);
xor U29944 (N_29944,N_29367,N_29172);
xor U29945 (N_29945,N_29210,N_29228);
nand U29946 (N_29946,N_29015,N_29164);
nand U29947 (N_29947,N_29455,N_29103);
xor U29948 (N_29948,N_29343,N_29140);
nand U29949 (N_29949,N_29131,N_29319);
or U29950 (N_29950,N_29338,N_29476);
and U29951 (N_29951,N_29085,N_29419);
nand U29952 (N_29952,N_29419,N_29067);
or U29953 (N_29953,N_29094,N_29402);
xor U29954 (N_29954,N_29246,N_29465);
nor U29955 (N_29955,N_29327,N_29332);
nand U29956 (N_29956,N_29118,N_29294);
and U29957 (N_29957,N_29009,N_29096);
nand U29958 (N_29958,N_29225,N_29331);
nor U29959 (N_29959,N_29384,N_29097);
nand U29960 (N_29960,N_29431,N_29499);
or U29961 (N_29961,N_29369,N_29135);
and U29962 (N_29962,N_29227,N_29482);
nor U29963 (N_29963,N_29301,N_29406);
or U29964 (N_29964,N_29495,N_29068);
or U29965 (N_29965,N_29319,N_29397);
nand U29966 (N_29966,N_29079,N_29133);
nor U29967 (N_29967,N_29081,N_29029);
nand U29968 (N_29968,N_29189,N_29229);
nand U29969 (N_29969,N_29016,N_29410);
or U29970 (N_29970,N_29336,N_29215);
nand U29971 (N_29971,N_29331,N_29376);
or U29972 (N_29972,N_29339,N_29193);
and U29973 (N_29973,N_29009,N_29046);
nor U29974 (N_29974,N_29417,N_29272);
and U29975 (N_29975,N_29056,N_29262);
nand U29976 (N_29976,N_29448,N_29422);
or U29977 (N_29977,N_29492,N_29397);
or U29978 (N_29978,N_29273,N_29253);
xor U29979 (N_29979,N_29468,N_29239);
or U29980 (N_29980,N_29103,N_29373);
or U29981 (N_29981,N_29236,N_29157);
nand U29982 (N_29982,N_29430,N_29285);
xor U29983 (N_29983,N_29358,N_29035);
nor U29984 (N_29984,N_29416,N_29182);
nand U29985 (N_29985,N_29290,N_29082);
xnor U29986 (N_29986,N_29355,N_29493);
nand U29987 (N_29987,N_29172,N_29479);
nor U29988 (N_29988,N_29165,N_29068);
and U29989 (N_29989,N_29036,N_29008);
or U29990 (N_29990,N_29169,N_29421);
or U29991 (N_29991,N_29121,N_29404);
and U29992 (N_29992,N_29493,N_29480);
nand U29993 (N_29993,N_29090,N_29067);
and U29994 (N_29994,N_29280,N_29487);
nor U29995 (N_29995,N_29388,N_29135);
and U29996 (N_29996,N_29292,N_29389);
or U29997 (N_29997,N_29073,N_29372);
xnor U29998 (N_29998,N_29373,N_29475);
or U29999 (N_29999,N_29469,N_29238);
or U30000 (N_30000,N_29987,N_29901);
or U30001 (N_30001,N_29669,N_29518);
or U30002 (N_30002,N_29641,N_29768);
xor U30003 (N_30003,N_29624,N_29652);
nand U30004 (N_30004,N_29918,N_29823);
and U30005 (N_30005,N_29612,N_29658);
and U30006 (N_30006,N_29573,N_29561);
nand U30007 (N_30007,N_29845,N_29967);
nand U30008 (N_30008,N_29826,N_29521);
nor U30009 (N_30009,N_29743,N_29922);
nand U30010 (N_30010,N_29968,N_29530);
and U30011 (N_30011,N_29729,N_29547);
nand U30012 (N_30012,N_29983,N_29992);
nor U30013 (N_30013,N_29995,N_29712);
xor U30014 (N_30014,N_29516,N_29778);
xnor U30015 (N_30015,N_29572,N_29811);
nor U30016 (N_30016,N_29595,N_29731);
and U30017 (N_30017,N_29500,N_29815);
nor U30018 (N_30018,N_29817,N_29505);
nand U30019 (N_30019,N_29606,N_29779);
xor U30020 (N_30020,N_29549,N_29849);
or U30021 (N_30021,N_29524,N_29791);
nand U30022 (N_30022,N_29852,N_29556);
nand U30023 (N_30023,N_29945,N_29875);
or U30024 (N_30024,N_29661,N_29977);
nor U30025 (N_30025,N_29905,N_29858);
nor U30026 (N_30026,N_29944,N_29859);
nor U30027 (N_30027,N_29850,N_29691);
or U30028 (N_30028,N_29884,N_29780);
xor U30029 (N_30029,N_29935,N_29754);
and U30030 (N_30030,N_29949,N_29957);
xor U30031 (N_30031,N_29843,N_29670);
nor U30032 (N_30032,N_29978,N_29896);
xor U30033 (N_30033,N_29985,N_29723);
xor U30034 (N_30034,N_29592,N_29913);
xor U30035 (N_30035,N_29684,N_29876);
and U30036 (N_30036,N_29747,N_29781);
or U30037 (N_30037,N_29761,N_29525);
or U30038 (N_30038,N_29623,N_29711);
nor U30039 (N_30039,N_29839,N_29520);
or U30040 (N_30040,N_29806,N_29504);
and U30041 (N_30041,N_29631,N_29636);
nand U30042 (N_30042,N_29716,N_29900);
nand U30043 (N_30043,N_29677,N_29954);
and U30044 (N_30044,N_29930,N_29535);
nor U30045 (N_30045,N_29756,N_29581);
nand U30046 (N_30046,N_29724,N_29557);
nor U30047 (N_30047,N_29651,N_29663);
nand U30048 (N_30048,N_29979,N_29667);
xor U30049 (N_30049,N_29857,N_29998);
or U30050 (N_30050,N_29709,N_29727);
nand U30051 (N_30051,N_29879,N_29923);
xnor U30052 (N_30052,N_29730,N_29671);
and U30053 (N_30053,N_29751,N_29996);
or U30054 (N_30054,N_29958,N_29868);
nand U30055 (N_30055,N_29862,N_29531);
xor U30056 (N_30056,N_29640,N_29609);
or U30057 (N_30057,N_29655,N_29621);
xor U30058 (N_30058,N_29738,N_29699);
nor U30059 (N_30059,N_29708,N_29582);
xor U30060 (N_30060,N_29537,N_29771);
nand U30061 (N_30061,N_29567,N_29757);
nor U30062 (N_30062,N_29745,N_29578);
or U30063 (N_30063,N_29886,N_29827);
nor U30064 (N_30064,N_29562,N_29566);
and U30065 (N_30065,N_29927,N_29584);
nor U30066 (N_30066,N_29774,N_29969);
nand U30067 (N_30067,N_29994,N_29555);
and U30068 (N_30068,N_29512,N_29855);
xnor U30069 (N_30069,N_29742,N_29615);
or U30070 (N_30070,N_29877,N_29642);
nand U30071 (N_30071,N_29719,N_29825);
nor U30072 (N_30072,N_29588,N_29821);
or U30073 (N_30073,N_29610,N_29763);
nor U30074 (N_30074,N_29540,N_29887);
xnor U30075 (N_30075,N_29666,N_29951);
and U30076 (N_30076,N_29689,N_29888);
xor U30077 (N_30077,N_29790,N_29637);
nor U30078 (N_30078,N_29630,N_29776);
or U30079 (N_30079,N_29902,N_29916);
nand U30080 (N_30080,N_29974,N_29721);
nand U30081 (N_30081,N_29787,N_29828);
and U30082 (N_30082,N_29664,N_29732);
and U30083 (N_30083,N_29596,N_29564);
xor U30084 (N_30084,N_29851,N_29509);
and U30085 (N_30085,N_29894,N_29848);
nor U30086 (N_30086,N_29660,N_29698);
nand U30087 (N_30087,N_29643,N_29799);
or U30088 (N_30088,N_29676,N_29812);
or U30089 (N_30089,N_29937,N_29874);
xnor U30090 (N_30090,N_29854,N_29601);
or U30091 (N_30091,N_29899,N_29717);
or U30092 (N_30092,N_29686,N_29617);
or U30093 (N_30093,N_29869,N_29818);
nand U30094 (N_30094,N_29559,N_29674);
nand U30095 (N_30095,N_29519,N_29841);
nor U30096 (N_30096,N_29837,N_29990);
or U30097 (N_30097,N_29980,N_29824);
nor U30098 (N_30098,N_29737,N_29593);
nand U30099 (N_30099,N_29526,N_29544);
or U30100 (N_30100,N_29972,N_29898);
nand U30101 (N_30101,N_29838,N_29628);
or U30102 (N_30102,N_29836,N_29543);
or U30103 (N_30103,N_29786,N_29539);
and U30104 (N_30104,N_29574,N_29694);
or U30105 (N_30105,N_29625,N_29608);
or U30106 (N_30106,N_29515,N_29668);
xor U30107 (N_30107,N_29613,N_29634);
and U30108 (N_30108,N_29911,N_29976);
xor U30109 (N_30109,N_29897,N_29605);
and U30110 (N_30110,N_29784,N_29679);
or U30111 (N_30111,N_29653,N_29867);
nor U30112 (N_30112,N_29506,N_29554);
and U30113 (N_30113,N_29614,N_29604);
or U30114 (N_30114,N_29750,N_29832);
and U30115 (N_30115,N_29696,N_29794);
nand U30116 (N_30116,N_29587,N_29616);
xor U30117 (N_30117,N_29563,N_29939);
and U30118 (N_30118,N_29864,N_29657);
nand U30119 (N_30119,N_29585,N_29508);
nor U30120 (N_30120,N_29702,N_29758);
nor U30121 (N_30121,N_29597,N_29802);
or U30122 (N_30122,N_29553,N_29770);
nand U30123 (N_30123,N_29704,N_29618);
nor U30124 (N_30124,N_29782,N_29880);
xor U30125 (N_30125,N_29736,N_29991);
or U30126 (N_30126,N_29924,N_29659);
nand U30127 (N_30127,N_29752,N_29589);
nor U30128 (N_30128,N_29932,N_29632);
nand U30129 (N_30129,N_29648,N_29558);
or U30130 (N_30130,N_29946,N_29813);
nor U30131 (N_30131,N_29956,N_29903);
nand U30132 (N_30132,N_29970,N_29542);
nand U30133 (N_30133,N_29649,N_29536);
xnor U30134 (N_30134,N_29744,N_29801);
and U30135 (N_30135,N_29796,N_29760);
nand U30136 (N_30136,N_29997,N_29656);
nand U30137 (N_30137,N_29871,N_29707);
xnor U30138 (N_30138,N_29984,N_29948);
xor U30139 (N_30139,N_29583,N_29591);
and U30140 (N_30140,N_29533,N_29919);
xor U30141 (N_30141,N_29928,N_29749);
nor U30142 (N_30142,N_29775,N_29840);
xnor U30143 (N_30143,N_29912,N_29870);
xnor U30144 (N_30144,N_29988,N_29860);
and U30145 (N_30145,N_29933,N_29940);
nand U30146 (N_30146,N_29726,N_29681);
and U30147 (N_30147,N_29947,N_29693);
nand U30148 (N_30148,N_29810,N_29816);
xor U30149 (N_30149,N_29599,N_29844);
nor U30150 (N_30150,N_29502,N_29690);
nor U30151 (N_30151,N_29622,N_29964);
or U30152 (N_30152,N_29703,N_29685);
nand U30153 (N_30153,N_29741,N_29759);
and U30154 (N_30154,N_29906,N_29706);
and U30155 (N_30155,N_29725,N_29882);
and U30156 (N_30156,N_29907,N_29586);
nand U30157 (N_30157,N_29568,N_29678);
and U30158 (N_30158,N_29603,N_29600);
nand U30159 (N_30159,N_29890,N_29626);
nand U30160 (N_30160,N_29904,N_29769);
or U30161 (N_30161,N_29647,N_29673);
or U30162 (N_30162,N_29680,N_29833);
and U30163 (N_30163,N_29639,N_29739);
and U30164 (N_30164,N_29507,N_29697);
or U30165 (N_30165,N_29962,N_29552);
xor U30166 (N_30166,N_29565,N_29834);
xnor U30167 (N_30167,N_29765,N_29943);
and U30168 (N_30168,N_29773,N_29772);
nor U30169 (N_30169,N_29793,N_29822);
and U30170 (N_30170,N_29528,N_29683);
nand U30171 (N_30171,N_29700,N_29955);
or U30172 (N_30172,N_29797,N_29654);
and U30173 (N_30173,N_29662,N_29701);
nand U30174 (N_30174,N_29873,N_29804);
xor U30175 (N_30175,N_29579,N_29611);
and U30176 (N_30176,N_29534,N_29878);
nand U30177 (N_30177,N_29808,N_29820);
xor U30178 (N_30178,N_29532,N_29783);
xnor U30179 (N_30179,N_29865,N_29513);
nor U30180 (N_30180,N_29715,N_29814);
and U30181 (N_30181,N_29705,N_29510);
and U30182 (N_30182,N_29672,N_29501);
and U30183 (N_30183,N_29594,N_29571);
nand U30184 (N_30184,N_29522,N_29748);
or U30185 (N_30185,N_29925,N_29546);
and U30186 (N_30186,N_29577,N_29527);
and U30187 (N_30187,N_29800,N_29740);
xor U30188 (N_30188,N_29627,N_29926);
nand U30189 (N_30189,N_29830,N_29620);
nor U30190 (N_30190,N_29728,N_29795);
and U30191 (N_30191,N_29819,N_29635);
nor U30192 (N_30192,N_29950,N_29767);
nor U30193 (N_30193,N_29872,N_29942);
xor U30194 (N_30194,N_29598,N_29503);
xor U30195 (N_30195,N_29720,N_29569);
and U30196 (N_30196,N_29785,N_29993);
or U30197 (N_30197,N_29638,N_29682);
and U30198 (N_30198,N_29665,N_29921);
and U30199 (N_30199,N_29734,N_29963);
and U30200 (N_30200,N_29710,N_29910);
or U30201 (N_30201,N_29953,N_29722);
nand U30202 (N_30202,N_29861,N_29931);
nor U30203 (N_30203,N_29803,N_29885);
nand U30204 (N_30204,N_29551,N_29883);
or U30205 (N_30205,N_29908,N_29733);
and U30206 (N_30206,N_29891,N_29692);
and U30207 (N_30207,N_29580,N_29966);
and U30208 (N_30208,N_29941,N_29881);
nand U30209 (N_30209,N_29853,N_29829);
nor U30210 (N_30210,N_29909,N_29619);
and U30211 (N_30211,N_29892,N_29917);
nor U30212 (N_30212,N_29889,N_29753);
or U30213 (N_30213,N_29523,N_29893);
and U30214 (N_30214,N_29576,N_29863);
nand U30215 (N_30215,N_29550,N_29975);
nand U30216 (N_30216,N_29777,N_29529);
nand U30217 (N_30217,N_29755,N_29842);
nand U30218 (N_30218,N_29789,N_29835);
and U30219 (N_30219,N_29590,N_29746);
xor U30220 (N_30220,N_29517,N_29560);
nand U30221 (N_30221,N_29989,N_29645);
or U30222 (N_30222,N_29798,N_29548);
xor U30223 (N_30223,N_29687,N_29846);
nor U30224 (N_30224,N_29809,N_29961);
and U30225 (N_30225,N_29973,N_29982);
nor U30226 (N_30226,N_29807,N_29831);
nor U30227 (N_30227,N_29650,N_29735);
nor U30228 (N_30228,N_29545,N_29538);
and U30229 (N_30229,N_29866,N_29986);
and U30230 (N_30230,N_29514,N_29646);
xor U30231 (N_30231,N_29633,N_29960);
or U30232 (N_30232,N_29570,N_29934);
nor U30233 (N_30233,N_29541,N_29999);
nor U30234 (N_30234,N_29788,N_29607);
and U30235 (N_30235,N_29602,N_29805);
or U30236 (N_30236,N_29644,N_29971);
or U30237 (N_30237,N_29575,N_29952);
or U30238 (N_30238,N_29718,N_29762);
and U30239 (N_30239,N_29675,N_29792);
and U30240 (N_30240,N_29914,N_29981);
xnor U30241 (N_30241,N_29915,N_29965);
or U30242 (N_30242,N_29695,N_29713);
nand U30243 (N_30243,N_29920,N_29938);
or U30244 (N_30244,N_29766,N_29629);
nand U30245 (N_30245,N_29959,N_29936);
nor U30246 (N_30246,N_29764,N_29511);
nand U30247 (N_30247,N_29714,N_29847);
nor U30248 (N_30248,N_29929,N_29856);
and U30249 (N_30249,N_29688,N_29895);
or U30250 (N_30250,N_29981,N_29670);
nor U30251 (N_30251,N_29850,N_29660);
nand U30252 (N_30252,N_29598,N_29711);
or U30253 (N_30253,N_29515,N_29520);
or U30254 (N_30254,N_29832,N_29566);
xnor U30255 (N_30255,N_29664,N_29834);
and U30256 (N_30256,N_29747,N_29993);
and U30257 (N_30257,N_29744,N_29725);
nand U30258 (N_30258,N_29654,N_29927);
xnor U30259 (N_30259,N_29958,N_29651);
or U30260 (N_30260,N_29689,N_29963);
xnor U30261 (N_30261,N_29632,N_29934);
or U30262 (N_30262,N_29931,N_29850);
nand U30263 (N_30263,N_29615,N_29695);
or U30264 (N_30264,N_29917,N_29734);
and U30265 (N_30265,N_29976,N_29522);
nand U30266 (N_30266,N_29537,N_29937);
xnor U30267 (N_30267,N_29740,N_29805);
and U30268 (N_30268,N_29785,N_29639);
or U30269 (N_30269,N_29952,N_29802);
and U30270 (N_30270,N_29885,N_29661);
nand U30271 (N_30271,N_29675,N_29569);
nor U30272 (N_30272,N_29603,N_29588);
and U30273 (N_30273,N_29714,N_29617);
or U30274 (N_30274,N_29784,N_29675);
xor U30275 (N_30275,N_29573,N_29805);
nor U30276 (N_30276,N_29792,N_29506);
and U30277 (N_30277,N_29691,N_29681);
nand U30278 (N_30278,N_29579,N_29887);
nand U30279 (N_30279,N_29859,N_29988);
or U30280 (N_30280,N_29938,N_29812);
and U30281 (N_30281,N_29863,N_29975);
or U30282 (N_30282,N_29751,N_29748);
nor U30283 (N_30283,N_29557,N_29804);
nor U30284 (N_30284,N_29669,N_29608);
xor U30285 (N_30285,N_29525,N_29751);
xnor U30286 (N_30286,N_29848,N_29915);
nand U30287 (N_30287,N_29657,N_29856);
or U30288 (N_30288,N_29942,N_29679);
nor U30289 (N_30289,N_29870,N_29896);
nand U30290 (N_30290,N_29922,N_29624);
nor U30291 (N_30291,N_29950,N_29954);
xnor U30292 (N_30292,N_29946,N_29575);
and U30293 (N_30293,N_29831,N_29778);
nor U30294 (N_30294,N_29529,N_29803);
xor U30295 (N_30295,N_29768,N_29730);
or U30296 (N_30296,N_29686,N_29618);
nand U30297 (N_30297,N_29623,N_29802);
and U30298 (N_30298,N_29711,N_29511);
and U30299 (N_30299,N_29756,N_29747);
nand U30300 (N_30300,N_29595,N_29522);
or U30301 (N_30301,N_29926,N_29670);
nand U30302 (N_30302,N_29614,N_29701);
or U30303 (N_30303,N_29874,N_29691);
or U30304 (N_30304,N_29884,N_29696);
and U30305 (N_30305,N_29535,N_29590);
or U30306 (N_30306,N_29606,N_29926);
nand U30307 (N_30307,N_29687,N_29782);
nand U30308 (N_30308,N_29977,N_29616);
or U30309 (N_30309,N_29949,N_29515);
and U30310 (N_30310,N_29900,N_29813);
nor U30311 (N_30311,N_29862,N_29568);
xnor U30312 (N_30312,N_29703,N_29761);
xor U30313 (N_30313,N_29715,N_29936);
nor U30314 (N_30314,N_29849,N_29721);
and U30315 (N_30315,N_29706,N_29947);
nor U30316 (N_30316,N_29798,N_29783);
or U30317 (N_30317,N_29548,N_29602);
xor U30318 (N_30318,N_29816,N_29869);
nand U30319 (N_30319,N_29643,N_29714);
and U30320 (N_30320,N_29583,N_29973);
or U30321 (N_30321,N_29664,N_29949);
or U30322 (N_30322,N_29879,N_29682);
xnor U30323 (N_30323,N_29571,N_29965);
xnor U30324 (N_30324,N_29727,N_29566);
or U30325 (N_30325,N_29876,N_29633);
and U30326 (N_30326,N_29779,N_29545);
xnor U30327 (N_30327,N_29689,N_29792);
nor U30328 (N_30328,N_29552,N_29752);
nor U30329 (N_30329,N_29716,N_29681);
xor U30330 (N_30330,N_29868,N_29754);
xnor U30331 (N_30331,N_29610,N_29827);
nor U30332 (N_30332,N_29870,N_29660);
and U30333 (N_30333,N_29848,N_29559);
and U30334 (N_30334,N_29910,N_29673);
xnor U30335 (N_30335,N_29532,N_29983);
xor U30336 (N_30336,N_29898,N_29926);
and U30337 (N_30337,N_29676,N_29657);
and U30338 (N_30338,N_29931,N_29666);
and U30339 (N_30339,N_29555,N_29720);
nor U30340 (N_30340,N_29618,N_29709);
or U30341 (N_30341,N_29714,N_29690);
xnor U30342 (N_30342,N_29773,N_29629);
xor U30343 (N_30343,N_29569,N_29845);
nand U30344 (N_30344,N_29592,N_29547);
and U30345 (N_30345,N_29607,N_29659);
nand U30346 (N_30346,N_29585,N_29803);
and U30347 (N_30347,N_29628,N_29923);
xnor U30348 (N_30348,N_29661,N_29997);
nor U30349 (N_30349,N_29953,N_29544);
or U30350 (N_30350,N_29952,N_29759);
or U30351 (N_30351,N_29507,N_29792);
nor U30352 (N_30352,N_29913,N_29946);
nand U30353 (N_30353,N_29677,N_29675);
xnor U30354 (N_30354,N_29554,N_29882);
nand U30355 (N_30355,N_29811,N_29886);
xnor U30356 (N_30356,N_29773,N_29661);
and U30357 (N_30357,N_29996,N_29533);
and U30358 (N_30358,N_29523,N_29549);
nor U30359 (N_30359,N_29721,N_29523);
or U30360 (N_30360,N_29822,N_29575);
xor U30361 (N_30361,N_29660,N_29775);
xnor U30362 (N_30362,N_29983,N_29558);
nand U30363 (N_30363,N_29733,N_29709);
xnor U30364 (N_30364,N_29887,N_29919);
nor U30365 (N_30365,N_29843,N_29605);
or U30366 (N_30366,N_29743,N_29543);
xnor U30367 (N_30367,N_29743,N_29952);
nor U30368 (N_30368,N_29967,N_29690);
and U30369 (N_30369,N_29979,N_29605);
and U30370 (N_30370,N_29584,N_29829);
or U30371 (N_30371,N_29738,N_29603);
nor U30372 (N_30372,N_29563,N_29581);
and U30373 (N_30373,N_29898,N_29515);
xnor U30374 (N_30374,N_29536,N_29611);
xor U30375 (N_30375,N_29892,N_29669);
nand U30376 (N_30376,N_29919,N_29955);
and U30377 (N_30377,N_29653,N_29854);
xor U30378 (N_30378,N_29631,N_29747);
nand U30379 (N_30379,N_29893,N_29736);
or U30380 (N_30380,N_29934,N_29843);
nor U30381 (N_30381,N_29693,N_29851);
nand U30382 (N_30382,N_29726,N_29917);
nor U30383 (N_30383,N_29854,N_29680);
nand U30384 (N_30384,N_29502,N_29561);
nand U30385 (N_30385,N_29581,N_29924);
nand U30386 (N_30386,N_29561,N_29528);
or U30387 (N_30387,N_29657,N_29971);
nand U30388 (N_30388,N_29789,N_29602);
xnor U30389 (N_30389,N_29570,N_29587);
nand U30390 (N_30390,N_29644,N_29681);
nor U30391 (N_30391,N_29963,N_29665);
and U30392 (N_30392,N_29900,N_29809);
nand U30393 (N_30393,N_29543,N_29700);
nand U30394 (N_30394,N_29565,N_29634);
xnor U30395 (N_30395,N_29697,N_29604);
nor U30396 (N_30396,N_29619,N_29745);
nand U30397 (N_30397,N_29973,N_29656);
nand U30398 (N_30398,N_29680,N_29801);
nor U30399 (N_30399,N_29577,N_29851);
or U30400 (N_30400,N_29536,N_29811);
nor U30401 (N_30401,N_29692,N_29621);
or U30402 (N_30402,N_29726,N_29843);
nor U30403 (N_30403,N_29959,N_29604);
or U30404 (N_30404,N_29686,N_29934);
or U30405 (N_30405,N_29852,N_29860);
and U30406 (N_30406,N_29953,N_29504);
nand U30407 (N_30407,N_29752,N_29733);
xnor U30408 (N_30408,N_29788,N_29613);
nand U30409 (N_30409,N_29500,N_29938);
and U30410 (N_30410,N_29934,N_29536);
nor U30411 (N_30411,N_29879,N_29502);
nor U30412 (N_30412,N_29904,N_29556);
and U30413 (N_30413,N_29945,N_29644);
nor U30414 (N_30414,N_29820,N_29959);
and U30415 (N_30415,N_29925,N_29549);
or U30416 (N_30416,N_29954,N_29644);
xnor U30417 (N_30417,N_29863,N_29924);
and U30418 (N_30418,N_29540,N_29780);
and U30419 (N_30419,N_29538,N_29927);
xor U30420 (N_30420,N_29896,N_29988);
and U30421 (N_30421,N_29595,N_29730);
nand U30422 (N_30422,N_29760,N_29882);
nand U30423 (N_30423,N_29672,N_29574);
or U30424 (N_30424,N_29973,N_29711);
nor U30425 (N_30425,N_29957,N_29731);
and U30426 (N_30426,N_29619,N_29891);
nor U30427 (N_30427,N_29763,N_29997);
nor U30428 (N_30428,N_29956,N_29688);
xnor U30429 (N_30429,N_29743,N_29729);
nor U30430 (N_30430,N_29773,N_29711);
nand U30431 (N_30431,N_29727,N_29763);
xor U30432 (N_30432,N_29984,N_29952);
xnor U30433 (N_30433,N_29948,N_29621);
or U30434 (N_30434,N_29711,N_29681);
and U30435 (N_30435,N_29741,N_29969);
xnor U30436 (N_30436,N_29972,N_29985);
or U30437 (N_30437,N_29786,N_29529);
or U30438 (N_30438,N_29743,N_29555);
nor U30439 (N_30439,N_29528,N_29578);
nor U30440 (N_30440,N_29545,N_29853);
nand U30441 (N_30441,N_29969,N_29689);
and U30442 (N_30442,N_29946,N_29795);
nor U30443 (N_30443,N_29650,N_29673);
xnor U30444 (N_30444,N_29686,N_29983);
nand U30445 (N_30445,N_29755,N_29645);
and U30446 (N_30446,N_29716,N_29935);
xor U30447 (N_30447,N_29795,N_29677);
nand U30448 (N_30448,N_29578,N_29842);
xnor U30449 (N_30449,N_29522,N_29580);
and U30450 (N_30450,N_29900,N_29669);
nor U30451 (N_30451,N_29512,N_29505);
nand U30452 (N_30452,N_29591,N_29909);
nor U30453 (N_30453,N_29961,N_29558);
nand U30454 (N_30454,N_29605,N_29917);
and U30455 (N_30455,N_29742,N_29618);
and U30456 (N_30456,N_29559,N_29911);
nand U30457 (N_30457,N_29900,N_29894);
or U30458 (N_30458,N_29850,N_29612);
xnor U30459 (N_30459,N_29857,N_29977);
xor U30460 (N_30460,N_29803,N_29739);
nor U30461 (N_30461,N_29990,N_29983);
xor U30462 (N_30462,N_29873,N_29572);
nor U30463 (N_30463,N_29561,N_29701);
nand U30464 (N_30464,N_29932,N_29693);
xor U30465 (N_30465,N_29547,N_29674);
or U30466 (N_30466,N_29878,N_29852);
or U30467 (N_30467,N_29932,N_29587);
xnor U30468 (N_30468,N_29567,N_29551);
nand U30469 (N_30469,N_29962,N_29571);
nor U30470 (N_30470,N_29699,N_29591);
and U30471 (N_30471,N_29545,N_29947);
or U30472 (N_30472,N_29937,N_29929);
and U30473 (N_30473,N_29978,N_29827);
and U30474 (N_30474,N_29801,N_29718);
and U30475 (N_30475,N_29555,N_29583);
nor U30476 (N_30476,N_29961,N_29548);
xor U30477 (N_30477,N_29926,N_29682);
and U30478 (N_30478,N_29647,N_29812);
xnor U30479 (N_30479,N_29998,N_29858);
xor U30480 (N_30480,N_29930,N_29697);
or U30481 (N_30481,N_29927,N_29576);
nor U30482 (N_30482,N_29512,N_29539);
nor U30483 (N_30483,N_29627,N_29938);
xnor U30484 (N_30484,N_29672,N_29762);
or U30485 (N_30485,N_29713,N_29974);
and U30486 (N_30486,N_29712,N_29728);
or U30487 (N_30487,N_29972,N_29949);
nand U30488 (N_30488,N_29841,N_29861);
nand U30489 (N_30489,N_29876,N_29658);
and U30490 (N_30490,N_29658,N_29619);
nand U30491 (N_30491,N_29954,N_29777);
or U30492 (N_30492,N_29585,N_29786);
and U30493 (N_30493,N_29730,N_29999);
nand U30494 (N_30494,N_29592,N_29713);
xnor U30495 (N_30495,N_29539,N_29791);
nand U30496 (N_30496,N_29676,N_29678);
nor U30497 (N_30497,N_29794,N_29727);
nand U30498 (N_30498,N_29792,N_29618);
and U30499 (N_30499,N_29610,N_29588);
and U30500 (N_30500,N_30485,N_30069);
nor U30501 (N_30501,N_30311,N_30113);
nand U30502 (N_30502,N_30003,N_30443);
xor U30503 (N_30503,N_30248,N_30020);
nand U30504 (N_30504,N_30436,N_30105);
or U30505 (N_30505,N_30049,N_30377);
and U30506 (N_30506,N_30396,N_30175);
xnor U30507 (N_30507,N_30164,N_30432);
xor U30508 (N_30508,N_30180,N_30232);
or U30509 (N_30509,N_30289,N_30317);
and U30510 (N_30510,N_30052,N_30177);
and U30511 (N_30511,N_30440,N_30280);
xor U30512 (N_30512,N_30413,N_30086);
and U30513 (N_30513,N_30424,N_30223);
nor U30514 (N_30514,N_30328,N_30470);
or U30515 (N_30515,N_30045,N_30383);
and U30516 (N_30516,N_30117,N_30406);
xnor U30517 (N_30517,N_30348,N_30015);
nor U30518 (N_30518,N_30090,N_30137);
nor U30519 (N_30519,N_30402,N_30335);
or U30520 (N_30520,N_30420,N_30465);
nand U30521 (N_30521,N_30495,N_30132);
xor U30522 (N_30522,N_30361,N_30190);
xnor U30523 (N_30523,N_30387,N_30059);
nand U30524 (N_30524,N_30179,N_30104);
and U30525 (N_30525,N_30423,N_30374);
or U30526 (N_30526,N_30303,N_30351);
and U30527 (N_30527,N_30360,N_30345);
or U30528 (N_30528,N_30365,N_30134);
nor U30529 (N_30529,N_30314,N_30235);
nor U30530 (N_30530,N_30191,N_30167);
xnor U30531 (N_30531,N_30487,N_30234);
nor U30532 (N_30532,N_30037,N_30123);
and U30533 (N_30533,N_30484,N_30079);
nand U30534 (N_30534,N_30208,N_30039);
xnor U30535 (N_30535,N_30467,N_30353);
or U30536 (N_30536,N_30414,N_30493);
xnor U30537 (N_30537,N_30083,N_30275);
or U30538 (N_30538,N_30033,N_30207);
nor U30539 (N_30539,N_30364,N_30437);
and U30540 (N_30540,N_30333,N_30258);
nand U30541 (N_30541,N_30498,N_30411);
xor U30542 (N_30542,N_30238,N_30142);
xor U30543 (N_30543,N_30141,N_30293);
or U30544 (N_30544,N_30260,N_30252);
nand U30545 (N_30545,N_30272,N_30202);
or U30546 (N_30546,N_30127,N_30192);
and U30547 (N_30547,N_30456,N_30473);
xnor U30548 (N_30548,N_30388,N_30077);
nand U30549 (N_30549,N_30426,N_30261);
nand U30550 (N_30550,N_30425,N_30497);
and U30551 (N_30551,N_30482,N_30469);
nand U30552 (N_30552,N_30165,N_30032);
nor U30553 (N_30553,N_30233,N_30403);
xor U30554 (N_30554,N_30087,N_30370);
and U30555 (N_30555,N_30188,N_30475);
nand U30556 (N_30556,N_30148,N_30285);
and U30557 (N_30557,N_30011,N_30041);
xor U30558 (N_30558,N_30005,N_30267);
nand U30559 (N_30559,N_30031,N_30243);
xor U30560 (N_30560,N_30135,N_30126);
or U30561 (N_30561,N_30189,N_30256);
nand U30562 (N_30562,N_30334,N_30363);
and U30563 (N_30563,N_30093,N_30390);
and U30564 (N_30564,N_30433,N_30157);
and U30565 (N_30565,N_30209,N_30014);
nor U30566 (N_30566,N_30446,N_30292);
or U30567 (N_30567,N_30103,N_30358);
nand U30568 (N_30568,N_30149,N_30236);
nor U30569 (N_30569,N_30125,N_30327);
nor U30570 (N_30570,N_30404,N_30176);
xnor U30571 (N_30571,N_30082,N_30155);
or U30572 (N_30572,N_30376,N_30254);
and U30573 (N_30573,N_30251,N_30009);
nand U30574 (N_30574,N_30051,N_30043);
or U30575 (N_30575,N_30462,N_30483);
nor U30576 (N_30576,N_30464,N_30295);
nor U30577 (N_30577,N_30129,N_30279);
and U30578 (N_30578,N_30128,N_30386);
xnor U30579 (N_30579,N_30085,N_30447);
nor U30580 (N_30580,N_30371,N_30060);
xor U30581 (N_30581,N_30407,N_30118);
nor U30582 (N_30582,N_30222,N_30409);
and U30583 (N_30583,N_30340,N_30078);
nor U30584 (N_30584,N_30047,N_30074);
and U30585 (N_30585,N_30160,N_30455);
xnor U30586 (N_30586,N_30042,N_30186);
and U30587 (N_30587,N_30013,N_30172);
nor U30588 (N_30588,N_30152,N_30076);
nor U30589 (N_30589,N_30318,N_30089);
or U30590 (N_30590,N_30322,N_30324);
and U30591 (N_30591,N_30389,N_30412);
xnor U30592 (N_30592,N_30018,N_30181);
or U30593 (N_30593,N_30193,N_30108);
and U30594 (N_30594,N_30101,N_30169);
nor U30595 (N_30595,N_30491,N_30080);
xnor U30596 (N_30596,N_30326,N_30415);
xnor U30597 (N_30597,N_30022,N_30271);
or U30598 (N_30598,N_30301,N_30174);
nor U30599 (N_30599,N_30244,N_30486);
and U30600 (N_30600,N_30109,N_30283);
and U30601 (N_30601,N_30457,N_30231);
xor U30602 (N_30602,N_30171,N_30441);
nor U30603 (N_30603,N_30266,N_30062);
nor U30604 (N_30604,N_30298,N_30075);
nor U30605 (N_30605,N_30489,N_30217);
nand U30606 (N_30606,N_30354,N_30300);
xnor U30607 (N_30607,N_30056,N_30144);
nand U30608 (N_30608,N_30290,N_30211);
xnor U30609 (N_30609,N_30325,N_30115);
xor U30610 (N_30610,N_30398,N_30268);
nand U30611 (N_30611,N_30000,N_30401);
or U30612 (N_30612,N_30023,N_30431);
or U30613 (N_30613,N_30323,N_30450);
xor U30614 (N_30614,N_30417,N_30378);
xor U30615 (N_30615,N_30224,N_30305);
and U30616 (N_30616,N_30106,N_30245);
xnor U30617 (N_30617,N_30029,N_30346);
nand U30618 (N_30618,N_30499,N_30368);
and U30619 (N_30619,N_30359,N_30435);
nor U30620 (N_30620,N_30269,N_30393);
nor U30621 (N_30621,N_30449,N_30380);
xnor U30622 (N_30622,N_30146,N_30265);
and U30623 (N_30623,N_30057,N_30241);
nor U30624 (N_30624,N_30071,N_30097);
and U30625 (N_30625,N_30344,N_30170);
or U30626 (N_30626,N_30416,N_30028);
and U30627 (N_30627,N_30206,N_30184);
nand U30628 (N_30628,N_30430,N_30130);
nor U30629 (N_30629,N_30400,N_30445);
nand U30630 (N_30630,N_30166,N_30496);
xor U30631 (N_30631,N_30151,N_30147);
nor U30632 (N_30632,N_30477,N_30427);
xor U30633 (N_30633,N_30320,N_30099);
and U30634 (N_30634,N_30024,N_30210);
nor U30635 (N_30635,N_30136,N_30145);
xor U30636 (N_30636,N_30366,N_30395);
nand U30637 (N_30637,N_30220,N_30138);
nor U30638 (N_30638,N_30307,N_30002);
xnor U30639 (N_30639,N_30088,N_30394);
nor U30640 (N_30640,N_30081,N_30439);
or U30641 (N_30641,N_30488,N_30084);
or U30642 (N_30642,N_30038,N_30150);
xnor U30643 (N_30643,N_30237,N_30219);
and U30644 (N_30644,N_30096,N_30228);
or U30645 (N_30645,N_30367,N_30384);
nor U30646 (N_30646,N_30050,N_30299);
and U30647 (N_30647,N_30274,N_30309);
or U30648 (N_30648,N_30214,N_30282);
and U30649 (N_30649,N_30478,N_30458);
xor U30650 (N_30650,N_30040,N_30247);
and U30651 (N_30651,N_30428,N_30154);
or U30652 (N_30652,N_30410,N_30310);
nor U30653 (N_30653,N_30092,N_30156);
and U30654 (N_30654,N_30225,N_30249);
xor U30655 (N_30655,N_30046,N_30054);
nor U30656 (N_30656,N_30195,N_30422);
nand U30657 (N_30657,N_30472,N_30315);
nand U30658 (N_30658,N_30392,N_30369);
xor U30659 (N_30659,N_30494,N_30421);
and U30660 (N_30660,N_30122,N_30007);
nand U30661 (N_30661,N_30316,N_30452);
nand U30662 (N_30662,N_30481,N_30296);
xor U30663 (N_30663,N_30454,N_30466);
and U30664 (N_30664,N_30194,N_30471);
xor U30665 (N_30665,N_30474,N_30408);
nand U30666 (N_30666,N_30330,N_30332);
nor U30667 (N_30667,N_30492,N_30203);
nor U30668 (N_30668,N_30372,N_30100);
nand U30669 (N_30669,N_30444,N_30429);
and U30670 (N_30670,N_30476,N_30215);
and U30671 (N_30671,N_30120,N_30490);
nor U30672 (N_30672,N_30385,N_30264);
xor U30673 (N_30673,N_30338,N_30198);
nand U30674 (N_30674,N_30027,N_30213);
nor U30675 (N_30675,N_30438,N_30112);
nor U30676 (N_30676,N_30331,N_30418);
xnor U30677 (N_30677,N_30070,N_30205);
or U30678 (N_30678,N_30263,N_30111);
or U30679 (N_30679,N_30068,N_30259);
nor U30680 (N_30680,N_30321,N_30017);
and U30681 (N_30681,N_30197,N_30227);
nor U30682 (N_30682,N_30357,N_30201);
and U30683 (N_30683,N_30356,N_30026);
or U30684 (N_30684,N_30319,N_30140);
nor U30685 (N_30685,N_30016,N_30459);
and U30686 (N_30686,N_30161,N_30313);
nor U30687 (N_30687,N_30379,N_30297);
and U30688 (N_30688,N_30284,N_30021);
nor U30689 (N_30689,N_30204,N_30434);
or U30690 (N_30690,N_30012,N_30347);
xor U30691 (N_30691,N_30064,N_30448);
nor U30692 (N_30692,N_30281,N_30067);
nor U30693 (N_30693,N_30162,N_30044);
nor U30694 (N_30694,N_30375,N_30173);
xnor U30695 (N_30695,N_30143,N_30405);
or U30696 (N_30696,N_30278,N_30114);
and U30697 (N_30697,N_30397,N_30006);
nand U30698 (N_30698,N_30183,N_30288);
nor U30699 (N_30699,N_30480,N_30153);
or U30700 (N_30700,N_30262,N_30158);
and U30701 (N_30701,N_30025,N_30312);
xnor U30702 (N_30702,N_30178,N_30239);
xor U30703 (N_30703,N_30066,N_30240);
nand U30704 (N_30704,N_30230,N_30095);
nor U30705 (N_30705,N_30373,N_30063);
xnor U30706 (N_30706,N_30072,N_30362);
or U30707 (N_30707,N_30461,N_30200);
nand U30708 (N_30708,N_30276,N_30419);
nor U30709 (N_30709,N_30034,N_30451);
nand U30710 (N_30710,N_30355,N_30350);
xor U30711 (N_30711,N_30329,N_30229);
xor U30712 (N_30712,N_30302,N_30163);
nand U30713 (N_30713,N_30304,N_30337);
and U30714 (N_30714,N_30286,N_30306);
or U30715 (N_30715,N_30463,N_30107);
or U30716 (N_30716,N_30246,N_30339);
nor U30717 (N_30717,N_30061,N_30212);
xor U30718 (N_30718,N_30159,N_30102);
nor U30719 (N_30719,N_30185,N_30182);
nand U30720 (N_30720,N_30253,N_30294);
and U30721 (N_30721,N_30291,N_30168);
and U30722 (N_30722,N_30255,N_30382);
nor U30723 (N_30723,N_30121,N_30030);
nor U30724 (N_30724,N_30019,N_30065);
nor U30725 (N_30725,N_30352,N_30381);
or U30726 (N_30726,N_30055,N_30391);
xnor U30727 (N_30727,N_30399,N_30308);
nor U30728 (N_30728,N_30035,N_30221);
nand U30729 (N_30729,N_30053,N_30139);
or U30730 (N_30730,N_30270,N_30133);
xnor U30731 (N_30731,N_30287,N_30442);
xnor U30732 (N_30732,N_30342,N_30479);
and U30733 (N_30733,N_30453,N_30001);
nand U30734 (N_30734,N_30091,N_30341);
nand U30735 (N_30735,N_30226,N_30336);
or U30736 (N_30736,N_30343,N_30098);
xnor U30737 (N_30737,N_30187,N_30257);
or U30738 (N_30738,N_30277,N_30460);
xor U30739 (N_30739,N_30110,N_30273);
nand U30740 (N_30740,N_30058,N_30048);
and U30741 (N_30741,N_30131,N_30216);
nand U30742 (N_30742,N_30468,N_30218);
and U30743 (N_30743,N_30242,N_30004);
xnor U30744 (N_30744,N_30250,N_30124);
and U30745 (N_30745,N_30196,N_30199);
or U30746 (N_30746,N_30010,N_30349);
xnor U30747 (N_30747,N_30008,N_30119);
xor U30748 (N_30748,N_30073,N_30094);
or U30749 (N_30749,N_30116,N_30036);
nand U30750 (N_30750,N_30456,N_30011);
or U30751 (N_30751,N_30045,N_30430);
nor U30752 (N_30752,N_30191,N_30100);
xor U30753 (N_30753,N_30256,N_30209);
and U30754 (N_30754,N_30382,N_30398);
and U30755 (N_30755,N_30030,N_30268);
xor U30756 (N_30756,N_30018,N_30138);
or U30757 (N_30757,N_30344,N_30104);
or U30758 (N_30758,N_30277,N_30418);
or U30759 (N_30759,N_30055,N_30245);
nor U30760 (N_30760,N_30324,N_30017);
nand U30761 (N_30761,N_30438,N_30341);
and U30762 (N_30762,N_30465,N_30170);
nor U30763 (N_30763,N_30091,N_30070);
and U30764 (N_30764,N_30270,N_30283);
or U30765 (N_30765,N_30228,N_30378);
nand U30766 (N_30766,N_30372,N_30491);
nand U30767 (N_30767,N_30254,N_30274);
and U30768 (N_30768,N_30402,N_30003);
nand U30769 (N_30769,N_30188,N_30377);
xor U30770 (N_30770,N_30004,N_30352);
nand U30771 (N_30771,N_30052,N_30395);
xnor U30772 (N_30772,N_30302,N_30470);
nand U30773 (N_30773,N_30458,N_30041);
nand U30774 (N_30774,N_30380,N_30240);
nand U30775 (N_30775,N_30179,N_30353);
xnor U30776 (N_30776,N_30417,N_30129);
xor U30777 (N_30777,N_30487,N_30445);
xor U30778 (N_30778,N_30024,N_30102);
or U30779 (N_30779,N_30297,N_30035);
xnor U30780 (N_30780,N_30065,N_30475);
nand U30781 (N_30781,N_30160,N_30432);
nand U30782 (N_30782,N_30485,N_30437);
and U30783 (N_30783,N_30432,N_30330);
nand U30784 (N_30784,N_30279,N_30433);
nand U30785 (N_30785,N_30082,N_30084);
or U30786 (N_30786,N_30171,N_30323);
xnor U30787 (N_30787,N_30457,N_30478);
xor U30788 (N_30788,N_30391,N_30414);
or U30789 (N_30789,N_30159,N_30095);
nand U30790 (N_30790,N_30203,N_30055);
and U30791 (N_30791,N_30373,N_30355);
and U30792 (N_30792,N_30122,N_30274);
nand U30793 (N_30793,N_30497,N_30419);
nand U30794 (N_30794,N_30215,N_30330);
or U30795 (N_30795,N_30188,N_30411);
nand U30796 (N_30796,N_30022,N_30014);
or U30797 (N_30797,N_30110,N_30189);
xnor U30798 (N_30798,N_30390,N_30079);
and U30799 (N_30799,N_30014,N_30206);
and U30800 (N_30800,N_30310,N_30144);
xnor U30801 (N_30801,N_30216,N_30086);
nand U30802 (N_30802,N_30195,N_30378);
and U30803 (N_30803,N_30078,N_30072);
nand U30804 (N_30804,N_30462,N_30166);
and U30805 (N_30805,N_30373,N_30086);
and U30806 (N_30806,N_30137,N_30174);
or U30807 (N_30807,N_30346,N_30363);
and U30808 (N_30808,N_30296,N_30099);
nand U30809 (N_30809,N_30351,N_30144);
or U30810 (N_30810,N_30083,N_30074);
nand U30811 (N_30811,N_30004,N_30347);
and U30812 (N_30812,N_30419,N_30050);
nand U30813 (N_30813,N_30447,N_30351);
nor U30814 (N_30814,N_30188,N_30318);
and U30815 (N_30815,N_30091,N_30134);
nor U30816 (N_30816,N_30290,N_30424);
nor U30817 (N_30817,N_30443,N_30107);
nand U30818 (N_30818,N_30148,N_30032);
nor U30819 (N_30819,N_30443,N_30401);
or U30820 (N_30820,N_30219,N_30032);
xor U30821 (N_30821,N_30094,N_30418);
and U30822 (N_30822,N_30458,N_30204);
and U30823 (N_30823,N_30109,N_30057);
and U30824 (N_30824,N_30074,N_30442);
or U30825 (N_30825,N_30367,N_30119);
nor U30826 (N_30826,N_30432,N_30390);
xor U30827 (N_30827,N_30462,N_30402);
and U30828 (N_30828,N_30270,N_30456);
and U30829 (N_30829,N_30408,N_30350);
nand U30830 (N_30830,N_30023,N_30301);
nand U30831 (N_30831,N_30091,N_30052);
nand U30832 (N_30832,N_30255,N_30484);
nand U30833 (N_30833,N_30492,N_30122);
nand U30834 (N_30834,N_30137,N_30139);
nor U30835 (N_30835,N_30491,N_30063);
nand U30836 (N_30836,N_30360,N_30068);
or U30837 (N_30837,N_30375,N_30481);
or U30838 (N_30838,N_30202,N_30135);
xor U30839 (N_30839,N_30037,N_30433);
or U30840 (N_30840,N_30336,N_30071);
or U30841 (N_30841,N_30377,N_30001);
and U30842 (N_30842,N_30041,N_30261);
nor U30843 (N_30843,N_30292,N_30261);
or U30844 (N_30844,N_30403,N_30335);
and U30845 (N_30845,N_30228,N_30126);
and U30846 (N_30846,N_30375,N_30476);
nand U30847 (N_30847,N_30209,N_30329);
nor U30848 (N_30848,N_30287,N_30049);
and U30849 (N_30849,N_30248,N_30153);
xnor U30850 (N_30850,N_30055,N_30050);
or U30851 (N_30851,N_30025,N_30041);
xnor U30852 (N_30852,N_30381,N_30204);
nor U30853 (N_30853,N_30288,N_30025);
nand U30854 (N_30854,N_30159,N_30139);
or U30855 (N_30855,N_30013,N_30141);
nand U30856 (N_30856,N_30389,N_30473);
nand U30857 (N_30857,N_30391,N_30352);
nor U30858 (N_30858,N_30051,N_30000);
nor U30859 (N_30859,N_30092,N_30102);
nor U30860 (N_30860,N_30127,N_30100);
or U30861 (N_30861,N_30426,N_30366);
xor U30862 (N_30862,N_30397,N_30348);
and U30863 (N_30863,N_30384,N_30401);
xnor U30864 (N_30864,N_30413,N_30096);
or U30865 (N_30865,N_30008,N_30336);
nor U30866 (N_30866,N_30126,N_30372);
and U30867 (N_30867,N_30229,N_30324);
nor U30868 (N_30868,N_30181,N_30036);
or U30869 (N_30869,N_30498,N_30199);
and U30870 (N_30870,N_30070,N_30423);
and U30871 (N_30871,N_30469,N_30095);
and U30872 (N_30872,N_30156,N_30051);
xor U30873 (N_30873,N_30494,N_30341);
nand U30874 (N_30874,N_30107,N_30268);
and U30875 (N_30875,N_30161,N_30058);
and U30876 (N_30876,N_30468,N_30408);
and U30877 (N_30877,N_30354,N_30266);
nand U30878 (N_30878,N_30157,N_30077);
xnor U30879 (N_30879,N_30064,N_30494);
nand U30880 (N_30880,N_30231,N_30210);
nand U30881 (N_30881,N_30432,N_30102);
xor U30882 (N_30882,N_30379,N_30485);
and U30883 (N_30883,N_30379,N_30261);
or U30884 (N_30884,N_30316,N_30088);
nor U30885 (N_30885,N_30257,N_30351);
nand U30886 (N_30886,N_30236,N_30404);
nand U30887 (N_30887,N_30305,N_30090);
nand U30888 (N_30888,N_30261,N_30383);
xor U30889 (N_30889,N_30493,N_30035);
and U30890 (N_30890,N_30404,N_30177);
nand U30891 (N_30891,N_30331,N_30212);
or U30892 (N_30892,N_30462,N_30222);
nand U30893 (N_30893,N_30063,N_30486);
xor U30894 (N_30894,N_30203,N_30054);
nor U30895 (N_30895,N_30107,N_30266);
and U30896 (N_30896,N_30396,N_30373);
or U30897 (N_30897,N_30128,N_30397);
nand U30898 (N_30898,N_30417,N_30242);
nor U30899 (N_30899,N_30237,N_30287);
nor U30900 (N_30900,N_30380,N_30370);
xnor U30901 (N_30901,N_30264,N_30187);
nand U30902 (N_30902,N_30121,N_30394);
xor U30903 (N_30903,N_30045,N_30217);
and U30904 (N_30904,N_30065,N_30080);
and U30905 (N_30905,N_30357,N_30385);
nand U30906 (N_30906,N_30249,N_30478);
xor U30907 (N_30907,N_30206,N_30429);
nand U30908 (N_30908,N_30416,N_30057);
and U30909 (N_30909,N_30357,N_30231);
and U30910 (N_30910,N_30001,N_30338);
nor U30911 (N_30911,N_30085,N_30260);
nand U30912 (N_30912,N_30351,N_30136);
and U30913 (N_30913,N_30385,N_30259);
nor U30914 (N_30914,N_30144,N_30063);
nand U30915 (N_30915,N_30289,N_30383);
nand U30916 (N_30916,N_30208,N_30389);
and U30917 (N_30917,N_30449,N_30043);
or U30918 (N_30918,N_30253,N_30200);
or U30919 (N_30919,N_30219,N_30371);
and U30920 (N_30920,N_30190,N_30188);
nor U30921 (N_30921,N_30073,N_30394);
nor U30922 (N_30922,N_30254,N_30333);
or U30923 (N_30923,N_30041,N_30037);
xnor U30924 (N_30924,N_30255,N_30152);
nand U30925 (N_30925,N_30017,N_30225);
or U30926 (N_30926,N_30004,N_30208);
nand U30927 (N_30927,N_30306,N_30413);
nand U30928 (N_30928,N_30053,N_30410);
nand U30929 (N_30929,N_30129,N_30253);
nor U30930 (N_30930,N_30432,N_30417);
or U30931 (N_30931,N_30090,N_30483);
xor U30932 (N_30932,N_30186,N_30021);
or U30933 (N_30933,N_30257,N_30163);
nor U30934 (N_30934,N_30452,N_30237);
nor U30935 (N_30935,N_30232,N_30306);
or U30936 (N_30936,N_30378,N_30144);
nor U30937 (N_30937,N_30066,N_30315);
xnor U30938 (N_30938,N_30252,N_30102);
nor U30939 (N_30939,N_30087,N_30460);
and U30940 (N_30940,N_30307,N_30276);
or U30941 (N_30941,N_30137,N_30167);
nand U30942 (N_30942,N_30052,N_30495);
and U30943 (N_30943,N_30038,N_30014);
nand U30944 (N_30944,N_30276,N_30131);
nor U30945 (N_30945,N_30459,N_30130);
nor U30946 (N_30946,N_30076,N_30462);
nand U30947 (N_30947,N_30145,N_30387);
or U30948 (N_30948,N_30313,N_30237);
and U30949 (N_30949,N_30230,N_30108);
xor U30950 (N_30950,N_30193,N_30184);
nand U30951 (N_30951,N_30309,N_30063);
nor U30952 (N_30952,N_30097,N_30040);
xor U30953 (N_30953,N_30233,N_30054);
or U30954 (N_30954,N_30044,N_30358);
nand U30955 (N_30955,N_30031,N_30183);
or U30956 (N_30956,N_30399,N_30200);
nor U30957 (N_30957,N_30261,N_30212);
xnor U30958 (N_30958,N_30080,N_30084);
xnor U30959 (N_30959,N_30321,N_30081);
nor U30960 (N_30960,N_30169,N_30482);
nand U30961 (N_30961,N_30190,N_30208);
nor U30962 (N_30962,N_30249,N_30335);
and U30963 (N_30963,N_30269,N_30262);
nand U30964 (N_30964,N_30420,N_30378);
or U30965 (N_30965,N_30097,N_30092);
or U30966 (N_30966,N_30219,N_30124);
xor U30967 (N_30967,N_30248,N_30406);
or U30968 (N_30968,N_30339,N_30283);
xnor U30969 (N_30969,N_30042,N_30005);
or U30970 (N_30970,N_30017,N_30472);
and U30971 (N_30971,N_30062,N_30452);
and U30972 (N_30972,N_30484,N_30296);
nor U30973 (N_30973,N_30375,N_30324);
nand U30974 (N_30974,N_30348,N_30178);
and U30975 (N_30975,N_30262,N_30347);
nor U30976 (N_30976,N_30330,N_30479);
nand U30977 (N_30977,N_30212,N_30389);
nand U30978 (N_30978,N_30353,N_30329);
nand U30979 (N_30979,N_30127,N_30471);
xor U30980 (N_30980,N_30383,N_30194);
nand U30981 (N_30981,N_30120,N_30135);
or U30982 (N_30982,N_30168,N_30147);
nor U30983 (N_30983,N_30224,N_30398);
or U30984 (N_30984,N_30158,N_30334);
xor U30985 (N_30985,N_30462,N_30072);
and U30986 (N_30986,N_30196,N_30314);
or U30987 (N_30987,N_30358,N_30383);
nor U30988 (N_30988,N_30184,N_30372);
or U30989 (N_30989,N_30355,N_30094);
xor U30990 (N_30990,N_30449,N_30255);
xor U30991 (N_30991,N_30015,N_30171);
nor U30992 (N_30992,N_30068,N_30291);
or U30993 (N_30993,N_30246,N_30449);
or U30994 (N_30994,N_30457,N_30495);
nand U30995 (N_30995,N_30491,N_30170);
nor U30996 (N_30996,N_30355,N_30087);
or U30997 (N_30997,N_30123,N_30077);
xor U30998 (N_30998,N_30061,N_30198);
and U30999 (N_30999,N_30376,N_30259);
or U31000 (N_31000,N_30965,N_30975);
and U31001 (N_31001,N_30868,N_30922);
and U31002 (N_31002,N_30822,N_30765);
and U31003 (N_31003,N_30585,N_30886);
nand U31004 (N_31004,N_30783,N_30695);
nand U31005 (N_31005,N_30699,N_30918);
or U31006 (N_31006,N_30731,N_30857);
nor U31007 (N_31007,N_30517,N_30727);
xor U31008 (N_31008,N_30998,N_30656);
and U31009 (N_31009,N_30907,N_30562);
xnor U31010 (N_31010,N_30753,N_30993);
nand U31011 (N_31011,N_30743,N_30528);
and U31012 (N_31012,N_30722,N_30715);
nor U31013 (N_31013,N_30635,N_30609);
and U31014 (N_31014,N_30682,N_30589);
xor U31015 (N_31015,N_30543,N_30734);
or U31016 (N_31016,N_30980,N_30798);
xnor U31017 (N_31017,N_30689,N_30991);
nand U31018 (N_31018,N_30866,N_30782);
nor U31019 (N_31019,N_30844,N_30704);
xor U31020 (N_31020,N_30941,N_30880);
xor U31021 (N_31021,N_30578,N_30651);
or U31022 (N_31022,N_30691,N_30852);
and U31023 (N_31023,N_30505,N_30570);
xor U31024 (N_31024,N_30851,N_30631);
and U31025 (N_31025,N_30660,N_30508);
nand U31026 (N_31026,N_30882,N_30776);
and U31027 (N_31027,N_30772,N_30616);
nand U31028 (N_31028,N_30780,N_30629);
xor U31029 (N_31029,N_30824,N_30919);
nor U31030 (N_31030,N_30754,N_30982);
nor U31031 (N_31031,N_30768,N_30825);
nor U31032 (N_31032,N_30519,N_30739);
nor U31033 (N_31033,N_30846,N_30921);
and U31034 (N_31034,N_30910,N_30775);
nand U31035 (N_31035,N_30872,N_30653);
nand U31036 (N_31036,N_30790,N_30735);
and U31037 (N_31037,N_30569,N_30712);
nor U31038 (N_31038,N_30710,N_30905);
or U31039 (N_31039,N_30697,N_30506);
and U31040 (N_31040,N_30668,N_30586);
or U31041 (N_31041,N_30939,N_30516);
xor U31042 (N_31042,N_30897,N_30583);
xnor U31043 (N_31043,N_30680,N_30549);
and U31044 (N_31044,N_30595,N_30946);
nor U31045 (N_31045,N_30805,N_30658);
xnor U31046 (N_31046,N_30864,N_30796);
nand U31047 (N_31047,N_30748,N_30746);
nor U31048 (N_31048,N_30669,N_30932);
or U31049 (N_31049,N_30675,N_30981);
and U31050 (N_31050,N_30632,N_30779);
or U31051 (N_31051,N_30626,N_30742);
or U31052 (N_31052,N_30771,N_30959);
or U31053 (N_31053,N_30613,N_30802);
and U31054 (N_31054,N_30555,N_30594);
nor U31055 (N_31055,N_30729,N_30944);
xnor U31056 (N_31056,N_30717,N_30719);
xor U31057 (N_31057,N_30614,N_30725);
nand U31058 (N_31058,N_30873,N_30639);
xnor U31059 (N_31059,N_30602,N_30869);
and U31060 (N_31060,N_30707,N_30502);
or U31061 (N_31061,N_30931,N_30924);
nor U31062 (N_31062,N_30995,N_30915);
nor U31063 (N_31063,N_30836,N_30581);
nor U31064 (N_31064,N_30553,N_30877);
or U31065 (N_31065,N_30920,N_30624);
nor U31066 (N_31066,N_30994,N_30795);
or U31067 (N_31067,N_30883,N_30679);
and U31068 (N_31068,N_30789,N_30612);
nand U31069 (N_31069,N_30812,N_30703);
and U31070 (N_31070,N_30533,N_30550);
or U31071 (N_31071,N_30898,N_30503);
xnor U31072 (N_31072,N_30638,N_30966);
nand U31073 (N_31073,N_30800,N_30558);
xnor U31074 (N_31074,N_30590,N_30832);
and U31075 (N_31075,N_30809,N_30620);
and U31076 (N_31076,N_30536,N_30591);
xor U31077 (N_31077,N_30777,N_30509);
nand U31078 (N_31078,N_30955,N_30531);
nand U31079 (N_31079,N_30996,N_30956);
nand U31080 (N_31080,N_30799,N_30925);
and U31081 (N_31081,N_30878,N_30816);
or U31082 (N_31082,N_30997,N_30504);
nand U31083 (N_31083,N_30511,N_30652);
or U31084 (N_31084,N_30523,N_30566);
or U31085 (N_31085,N_30761,N_30501);
nor U31086 (N_31086,N_30810,N_30987);
nor U31087 (N_31087,N_30557,N_30950);
and U31088 (N_31088,N_30870,N_30821);
and U31089 (N_31089,N_30976,N_30530);
and U31090 (N_31090,N_30999,N_30584);
nor U31091 (N_31091,N_30716,N_30657);
nor U31092 (N_31092,N_30641,N_30692);
nor U31093 (N_31093,N_30573,N_30527);
or U31094 (N_31094,N_30636,N_30673);
and U31095 (N_31095,N_30625,N_30733);
and U31096 (N_31096,N_30762,N_30526);
or U31097 (N_31097,N_30760,N_30940);
nand U31098 (N_31098,N_30740,N_30858);
xor U31099 (N_31099,N_30670,N_30726);
nor U31100 (N_31100,N_30512,N_30876);
and U31101 (N_31101,N_30744,N_30930);
or U31102 (N_31102,N_30885,N_30659);
nand U31103 (N_31103,N_30827,N_30648);
xnor U31104 (N_31104,N_30769,N_30745);
or U31105 (N_31105,N_30698,N_30811);
xor U31106 (N_31106,N_30559,N_30714);
nand U31107 (N_31107,N_30646,N_30900);
xor U31108 (N_31108,N_30867,N_30677);
and U31109 (N_31109,N_30603,N_30807);
nor U31110 (N_31110,N_30911,N_30804);
xnor U31111 (N_31111,N_30913,N_30974);
xor U31112 (N_31112,N_30843,N_30791);
and U31113 (N_31113,N_30556,N_30902);
xor U31114 (N_31114,N_30676,N_30899);
or U31115 (N_31115,N_30537,N_30601);
xor U31116 (N_31116,N_30947,N_30784);
nor U31117 (N_31117,N_30606,N_30713);
nand U31118 (N_31118,N_30667,N_30705);
nor U31119 (N_31119,N_30985,N_30644);
or U31120 (N_31120,N_30865,N_30879);
and U31121 (N_31121,N_30835,N_30934);
or U31122 (N_31122,N_30633,N_30935);
xnor U31123 (N_31123,N_30622,N_30514);
nand U31124 (N_31124,N_30888,N_30814);
and U31125 (N_31125,N_30801,N_30618);
xnor U31126 (N_31126,N_30929,N_30671);
nor U31127 (N_31127,N_30515,N_30895);
or U31128 (N_31128,N_30607,N_30684);
nand U31129 (N_31129,N_30926,N_30903);
and U31130 (N_31130,N_30706,N_30828);
and U31131 (N_31131,N_30617,N_30637);
nand U31132 (N_31132,N_30850,N_30649);
nand U31133 (N_31133,N_30535,N_30928);
or U31134 (N_31134,N_30723,N_30741);
nor U31135 (N_31135,N_30938,N_30849);
and U31136 (N_31136,N_30596,N_30778);
xnor U31137 (N_31137,N_30834,N_30874);
nand U31138 (N_31138,N_30972,N_30859);
nand U31139 (N_31139,N_30576,N_30605);
xor U31140 (N_31140,N_30847,N_30848);
and U31141 (N_31141,N_30973,N_30551);
nor U31142 (N_31142,N_30884,N_30520);
xor U31143 (N_31143,N_30964,N_30529);
nor U31144 (N_31144,N_30856,N_30575);
nor U31145 (N_31145,N_30724,N_30957);
or U31146 (N_31146,N_30923,N_30970);
and U31147 (N_31147,N_30540,N_30788);
and U31148 (N_31148,N_30690,N_30665);
nand U31149 (N_31149,N_30702,N_30983);
nand U31150 (N_31150,N_30579,N_30561);
and U31151 (N_31151,N_30942,N_30654);
xnor U31152 (N_31152,N_30841,N_30820);
and U31153 (N_31153,N_30645,N_30563);
or U31154 (N_31154,N_30611,N_30830);
nor U31155 (N_31155,N_30781,N_30989);
nor U31156 (N_31156,N_30554,N_30855);
nor U31157 (N_31157,N_30621,N_30896);
xor U31158 (N_31158,N_30688,N_30891);
or U31159 (N_31159,N_30948,N_30747);
nor U31160 (N_31160,N_30806,N_30518);
and U31161 (N_31161,N_30738,N_30521);
nor U31162 (N_31162,N_30737,N_30541);
and U31163 (N_31163,N_30650,N_30861);
or U31164 (N_31164,N_30732,N_30979);
nor U31165 (N_31165,N_30507,N_30906);
xnor U31166 (N_31166,N_30971,N_30608);
or U31167 (N_31167,N_30890,N_30752);
xnor U31168 (N_31168,N_30937,N_30952);
nor U31169 (N_31169,N_30787,N_30666);
nand U31170 (N_31170,N_30875,N_30615);
or U31171 (N_31171,N_30840,N_30916);
nor U31172 (N_31172,N_30992,N_30962);
or U31173 (N_31173,N_30773,N_30958);
and U31174 (N_31174,N_30592,N_30917);
nand U31175 (N_31175,N_30610,N_30647);
or U31176 (N_31176,N_30571,N_30604);
nand U31177 (N_31177,N_30893,N_30580);
nand U31178 (N_31178,N_30709,N_30863);
nand U31179 (N_31179,N_30845,N_30539);
and U31180 (N_31180,N_30687,N_30547);
or U31181 (N_31181,N_30642,N_30524);
nor U31182 (N_31182,N_30862,N_30853);
and U31183 (N_31183,N_30730,N_30546);
and U31184 (N_31184,N_30661,N_30600);
nor U31185 (N_31185,N_30678,N_30534);
or U31186 (N_31186,N_30860,N_30718);
nor U31187 (N_31187,N_30829,N_30767);
and U31188 (N_31188,N_30587,N_30577);
xor U31189 (N_31189,N_30871,N_30967);
nor U31190 (N_31190,N_30588,N_30751);
or U31191 (N_31191,N_30758,N_30815);
nor U31192 (N_31192,N_30817,N_30977);
nand U31193 (N_31193,N_30525,N_30513);
and U31194 (N_31194,N_30826,N_30510);
nand U31195 (N_31195,N_30623,N_30990);
nor U31196 (N_31196,N_30954,N_30672);
or U31197 (N_31197,N_30969,N_30560);
xnor U31198 (N_31198,N_30598,N_30538);
nand U31199 (N_31199,N_30894,N_30968);
or U31200 (N_31200,N_30839,N_30701);
nand U31201 (N_31201,N_30833,N_30988);
nor U31202 (N_31202,N_30774,N_30755);
xnor U31203 (N_31203,N_30803,N_30818);
or U31204 (N_31204,N_30945,N_30889);
and U31205 (N_31205,N_30770,N_30593);
and U31206 (N_31206,N_30693,N_30854);
nor U31207 (N_31207,N_30663,N_30978);
nand U31208 (N_31208,N_30597,N_30685);
xnor U31209 (N_31209,N_30887,N_30963);
or U31210 (N_31210,N_30912,N_30640);
nand U31211 (N_31211,N_30914,N_30681);
nand U31212 (N_31212,N_30831,N_30548);
or U31213 (N_31213,N_30749,N_30711);
xor U31214 (N_31214,N_30674,N_30881);
or U31215 (N_31215,N_30500,N_30686);
and U31216 (N_31216,N_30764,N_30567);
nor U31217 (N_31217,N_30574,N_30627);
or U31218 (N_31218,N_30984,N_30662);
nor U31219 (N_31219,N_30552,N_30813);
nand U31220 (N_31220,N_30936,N_30757);
or U31221 (N_31221,N_30785,N_30808);
nor U31222 (N_31222,N_30720,N_30927);
nor U31223 (N_31223,N_30700,N_30943);
nor U31224 (N_31224,N_30545,N_30694);
and U31225 (N_31225,N_30683,N_30792);
xnor U31226 (N_31226,N_30901,N_30750);
and U31227 (N_31227,N_30819,N_30763);
nand U31228 (N_31228,N_30634,N_30766);
xor U31229 (N_31229,N_30619,N_30532);
nor U31230 (N_31230,N_30664,N_30542);
or U31231 (N_31231,N_30599,N_30708);
and U31232 (N_31232,N_30961,N_30842);
nor U31233 (N_31233,N_30544,N_30728);
or U31234 (N_31234,N_30630,N_30756);
nand U31235 (N_31235,N_30986,N_30823);
nand U31236 (N_31236,N_30953,N_30572);
nand U31237 (N_31237,N_30522,N_30582);
nand U31238 (N_31238,N_30949,N_30655);
or U31239 (N_31239,N_30908,N_30794);
or U31240 (N_31240,N_30909,N_30797);
xnor U31241 (N_31241,N_30793,N_30759);
and U31242 (N_31242,N_30786,N_30951);
or U31243 (N_31243,N_30564,N_30892);
nor U31244 (N_31244,N_30628,N_30960);
nor U31245 (N_31245,N_30933,N_30565);
xor U31246 (N_31246,N_30721,N_30568);
nor U31247 (N_31247,N_30736,N_30837);
xor U31248 (N_31248,N_30696,N_30904);
nor U31249 (N_31249,N_30838,N_30643);
nand U31250 (N_31250,N_30773,N_30682);
and U31251 (N_31251,N_30702,N_30598);
or U31252 (N_31252,N_30914,N_30802);
nor U31253 (N_31253,N_30796,N_30536);
nand U31254 (N_31254,N_30851,N_30843);
and U31255 (N_31255,N_30978,N_30667);
and U31256 (N_31256,N_30825,N_30544);
and U31257 (N_31257,N_30510,N_30942);
and U31258 (N_31258,N_30708,N_30503);
xor U31259 (N_31259,N_30965,N_30602);
or U31260 (N_31260,N_30941,N_30715);
and U31261 (N_31261,N_30831,N_30676);
or U31262 (N_31262,N_30811,N_30846);
and U31263 (N_31263,N_30928,N_30583);
nor U31264 (N_31264,N_30955,N_30879);
xnor U31265 (N_31265,N_30580,N_30563);
nor U31266 (N_31266,N_30835,N_30771);
and U31267 (N_31267,N_30612,N_30503);
nor U31268 (N_31268,N_30770,N_30677);
xnor U31269 (N_31269,N_30852,N_30571);
and U31270 (N_31270,N_30730,N_30709);
nor U31271 (N_31271,N_30983,N_30753);
nand U31272 (N_31272,N_30840,N_30926);
nor U31273 (N_31273,N_30564,N_30545);
xor U31274 (N_31274,N_30607,N_30803);
xor U31275 (N_31275,N_30610,N_30674);
nor U31276 (N_31276,N_30886,N_30945);
and U31277 (N_31277,N_30925,N_30580);
and U31278 (N_31278,N_30944,N_30806);
nand U31279 (N_31279,N_30660,N_30901);
or U31280 (N_31280,N_30851,N_30609);
nand U31281 (N_31281,N_30599,N_30739);
or U31282 (N_31282,N_30923,N_30973);
nand U31283 (N_31283,N_30707,N_30748);
or U31284 (N_31284,N_30650,N_30924);
and U31285 (N_31285,N_30686,N_30886);
and U31286 (N_31286,N_30621,N_30640);
and U31287 (N_31287,N_30755,N_30677);
nor U31288 (N_31288,N_30928,N_30711);
xor U31289 (N_31289,N_30550,N_30992);
xnor U31290 (N_31290,N_30753,N_30583);
xnor U31291 (N_31291,N_30799,N_30766);
xnor U31292 (N_31292,N_30745,N_30522);
nor U31293 (N_31293,N_30983,N_30813);
or U31294 (N_31294,N_30575,N_30875);
nand U31295 (N_31295,N_30702,N_30504);
nand U31296 (N_31296,N_30665,N_30865);
nor U31297 (N_31297,N_30537,N_30534);
nor U31298 (N_31298,N_30574,N_30537);
nand U31299 (N_31299,N_30858,N_30651);
or U31300 (N_31300,N_30712,N_30610);
nand U31301 (N_31301,N_30947,N_30597);
nand U31302 (N_31302,N_30933,N_30722);
nand U31303 (N_31303,N_30538,N_30809);
nor U31304 (N_31304,N_30548,N_30976);
and U31305 (N_31305,N_30792,N_30594);
nor U31306 (N_31306,N_30741,N_30927);
nor U31307 (N_31307,N_30986,N_30773);
or U31308 (N_31308,N_30772,N_30584);
or U31309 (N_31309,N_30801,N_30853);
or U31310 (N_31310,N_30727,N_30800);
nand U31311 (N_31311,N_30577,N_30573);
and U31312 (N_31312,N_30651,N_30571);
or U31313 (N_31313,N_30778,N_30517);
or U31314 (N_31314,N_30546,N_30903);
or U31315 (N_31315,N_30995,N_30649);
and U31316 (N_31316,N_30972,N_30655);
nand U31317 (N_31317,N_30873,N_30596);
xnor U31318 (N_31318,N_30780,N_30894);
xor U31319 (N_31319,N_30770,N_30766);
nor U31320 (N_31320,N_30679,N_30884);
nand U31321 (N_31321,N_30740,N_30655);
or U31322 (N_31322,N_30540,N_30918);
xnor U31323 (N_31323,N_30911,N_30557);
and U31324 (N_31324,N_30860,N_30533);
or U31325 (N_31325,N_30919,N_30858);
nand U31326 (N_31326,N_30866,N_30923);
or U31327 (N_31327,N_30654,N_30861);
and U31328 (N_31328,N_30707,N_30906);
or U31329 (N_31329,N_30954,N_30878);
xor U31330 (N_31330,N_30533,N_30543);
nand U31331 (N_31331,N_30865,N_30739);
and U31332 (N_31332,N_30598,N_30991);
xnor U31333 (N_31333,N_30685,N_30788);
or U31334 (N_31334,N_30804,N_30739);
nand U31335 (N_31335,N_30957,N_30788);
xor U31336 (N_31336,N_30769,N_30501);
nor U31337 (N_31337,N_30515,N_30533);
or U31338 (N_31338,N_30568,N_30547);
nor U31339 (N_31339,N_30589,N_30942);
nor U31340 (N_31340,N_30708,N_30883);
nand U31341 (N_31341,N_30697,N_30570);
nor U31342 (N_31342,N_30763,N_30595);
nor U31343 (N_31343,N_30705,N_30712);
nor U31344 (N_31344,N_30947,N_30787);
nand U31345 (N_31345,N_30843,N_30935);
nor U31346 (N_31346,N_30828,N_30738);
xnor U31347 (N_31347,N_30993,N_30602);
nor U31348 (N_31348,N_30568,N_30565);
xnor U31349 (N_31349,N_30649,N_30817);
or U31350 (N_31350,N_30549,N_30708);
or U31351 (N_31351,N_30683,N_30736);
or U31352 (N_31352,N_30578,N_30521);
nor U31353 (N_31353,N_30868,N_30699);
and U31354 (N_31354,N_30642,N_30854);
xnor U31355 (N_31355,N_30820,N_30676);
nand U31356 (N_31356,N_30946,N_30516);
xor U31357 (N_31357,N_30969,N_30926);
or U31358 (N_31358,N_30794,N_30927);
nor U31359 (N_31359,N_30672,N_30737);
xnor U31360 (N_31360,N_30561,N_30762);
nor U31361 (N_31361,N_30639,N_30955);
nor U31362 (N_31362,N_30541,N_30911);
nor U31363 (N_31363,N_30874,N_30832);
nand U31364 (N_31364,N_30554,N_30971);
nor U31365 (N_31365,N_30731,N_30890);
nand U31366 (N_31366,N_30700,N_30988);
xnor U31367 (N_31367,N_30632,N_30732);
nand U31368 (N_31368,N_30975,N_30978);
or U31369 (N_31369,N_30727,N_30750);
xor U31370 (N_31370,N_30703,N_30868);
xor U31371 (N_31371,N_30896,N_30529);
nor U31372 (N_31372,N_30603,N_30854);
nor U31373 (N_31373,N_30883,N_30700);
xor U31374 (N_31374,N_30576,N_30526);
xnor U31375 (N_31375,N_30509,N_30714);
nor U31376 (N_31376,N_30862,N_30939);
nor U31377 (N_31377,N_30543,N_30717);
or U31378 (N_31378,N_30997,N_30545);
xor U31379 (N_31379,N_30775,N_30690);
xor U31380 (N_31380,N_30981,N_30560);
nand U31381 (N_31381,N_30520,N_30970);
nand U31382 (N_31382,N_30595,N_30649);
nor U31383 (N_31383,N_30644,N_30957);
nand U31384 (N_31384,N_30872,N_30823);
nand U31385 (N_31385,N_30583,N_30794);
nor U31386 (N_31386,N_30743,N_30566);
and U31387 (N_31387,N_30917,N_30825);
nor U31388 (N_31388,N_30623,N_30951);
nand U31389 (N_31389,N_30958,N_30906);
nor U31390 (N_31390,N_30935,N_30972);
xor U31391 (N_31391,N_30693,N_30757);
xor U31392 (N_31392,N_30877,N_30562);
nand U31393 (N_31393,N_30895,N_30862);
nand U31394 (N_31394,N_30943,N_30591);
xnor U31395 (N_31395,N_30631,N_30538);
nand U31396 (N_31396,N_30927,N_30690);
xor U31397 (N_31397,N_30638,N_30597);
and U31398 (N_31398,N_30940,N_30728);
xor U31399 (N_31399,N_30622,N_30860);
and U31400 (N_31400,N_30546,N_30981);
and U31401 (N_31401,N_30508,N_30949);
nor U31402 (N_31402,N_30673,N_30935);
nand U31403 (N_31403,N_30714,N_30511);
and U31404 (N_31404,N_30741,N_30966);
nand U31405 (N_31405,N_30845,N_30719);
nand U31406 (N_31406,N_30969,N_30674);
xnor U31407 (N_31407,N_30650,N_30806);
nand U31408 (N_31408,N_30878,N_30741);
nand U31409 (N_31409,N_30974,N_30599);
and U31410 (N_31410,N_30663,N_30949);
or U31411 (N_31411,N_30881,N_30919);
nor U31412 (N_31412,N_30891,N_30754);
xnor U31413 (N_31413,N_30857,N_30576);
xnor U31414 (N_31414,N_30887,N_30958);
xnor U31415 (N_31415,N_30745,N_30867);
nand U31416 (N_31416,N_30559,N_30950);
nand U31417 (N_31417,N_30502,N_30728);
xnor U31418 (N_31418,N_30994,N_30928);
nor U31419 (N_31419,N_30866,N_30867);
nand U31420 (N_31420,N_30918,N_30618);
xnor U31421 (N_31421,N_30630,N_30694);
and U31422 (N_31422,N_30762,N_30933);
or U31423 (N_31423,N_30525,N_30721);
and U31424 (N_31424,N_30978,N_30852);
or U31425 (N_31425,N_30737,N_30925);
xnor U31426 (N_31426,N_30648,N_30997);
nand U31427 (N_31427,N_30837,N_30625);
and U31428 (N_31428,N_30943,N_30860);
nor U31429 (N_31429,N_30880,N_30594);
nor U31430 (N_31430,N_30697,N_30512);
or U31431 (N_31431,N_30979,N_30503);
xnor U31432 (N_31432,N_30580,N_30877);
or U31433 (N_31433,N_30766,N_30975);
xnor U31434 (N_31434,N_30547,N_30876);
nor U31435 (N_31435,N_30985,N_30928);
and U31436 (N_31436,N_30573,N_30640);
and U31437 (N_31437,N_30804,N_30802);
or U31438 (N_31438,N_30758,N_30680);
or U31439 (N_31439,N_30847,N_30620);
nand U31440 (N_31440,N_30934,N_30546);
nand U31441 (N_31441,N_30979,N_30664);
or U31442 (N_31442,N_30770,N_30793);
or U31443 (N_31443,N_30914,N_30638);
nand U31444 (N_31444,N_30652,N_30746);
and U31445 (N_31445,N_30994,N_30805);
and U31446 (N_31446,N_30569,N_30544);
xor U31447 (N_31447,N_30969,N_30982);
xor U31448 (N_31448,N_30917,N_30922);
and U31449 (N_31449,N_30913,N_30555);
nor U31450 (N_31450,N_30980,N_30959);
xnor U31451 (N_31451,N_30877,N_30737);
nor U31452 (N_31452,N_30765,N_30838);
and U31453 (N_31453,N_30669,N_30949);
nand U31454 (N_31454,N_30753,N_30929);
or U31455 (N_31455,N_30530,N_30762);
or U31456 (N_31456,N_30575,N_30587);
nor U31457 (N_31457,N_30994,N_30840);
or U31458 (N_31458,N_30904,N_30776);
nand U31459 (N_31459,N_30570,N_30557);
xnor U31460 (N_31460,N_30789,N_30938);
nand U31461 (N_31461,N_30881,N_30945);
and U31462 (N_31462,N_30722,N_30541);
or U31463 (N_31463,N_30500,N_30691);
or U31464 (N_31464,N_30767,N_30950);
xnor U31465 (N_31465,N_30623,N_30997);
nand U31466 (N_31466,N_30835,N_30812);
or U31467 (N_31467,N_30899,N_30838);
nor U31468 (N_31468,N_30801,N_30785);
nand U31469 (N_31469,N_30606,N_30734);
or U31470 (N_31470,N_30638,N_30669);
and U31471 (N_31471,N_30900,N_30521);
xor U31472 (N_31472,N_30782,N_30916);
or U31473 (N_31473,N_30672,N_30973);
or U31474 (N_31474,N_30644,N_30973);
xor U31475 (N_31475,N_30995,N_30648);
nand U31476 (N_31476,N_30693,N_30770);
or U31477 (N_31477,N_30959,N_30721);
nand U31478 (N_31478,N_30762,N_30664);
and U31479 (N_31479,N_30522,N_30804);
or U31480 (N_31480,N_30861,N_30684);
xnor U31481 (N_31481,N_30820,N_30793);
xnor U31482 (N_31482,N_30912,N_30849);
xor U31483 (N_31483,N_30536,N_30520);
and U31484 (N_31484,N_30561,N_30928);
or U31485 (N_31485,N_30605,N_30635);
or U31486 (N_31486,N_30858,N_30789);
nand U31487 (N_31487,N_30753,N_30653);
xnor U31488 (N_31488,N_30756,N_30720);
or U31489 (N_31489,N_30637,N_30741);
xor U31490 (N_31490,N_30570,N_30869);
xnor U31491 (N_31491,N_30917,N_30718);
xnor U31492 (N_31492,N_30770,N_30618);
and U31493 (N_31493,N_30698,N_30927);
or U31494 (N_31494,N_30870,N_30703);
nand U31495 (N_31495,N_30892,N_30928);
xor U31496 (N_31496,N_30794,N_30813);
or U31497 (N_31497,N_30817,N_30568);
or U31498 (N_31498,N_30851,N_30939);
xnor U31499 (N_31499,N_30971,N_30701);
nor U31500 (N_31500,N_31144,N_31497);
nand U31501 (N_31501,N_31450,N_31118);
or U31502 (N_31502,N_31105,N_31174);
and U31503 (N_31503,N_31415,N_31356);
and U31504 (N_31504,N_31158,N_31404);
nand U31505 (N_31505,N_31456,N_31433);
xor U31506 (N_31506,N_31432,N_31452);
nand U31507 (N_31507,N_31303,N_31413);
and U31508 (N_31508,N_31188,N_31051);
nor U31509 (N_31509,N_31238,N_31498);
nand U31510 (N_31510,N_31459,N_31397);
and U31511 (N_31511,N_31420,N_31049);
xnor U31512 (N_31512,N_31067,N_31085);
nor U31513 (N_31513,N_31379,N_31329);
or U31514 (N_31514,N_31249,N_31083);
xnor U31515 (N_31515,N_31493,N_31108);
and U31516 (N_31516,N_31159,N_31279);
xnor U31517 (N_31517,N_31468,N_31295);
xor U31518 (N_31518,N_31489,N_31097);
or U31519 (N_31519,N_31360,N_31488);
xor U31520 (N_31520,N_31322,N_31043);
or U31521 (N_31521,N_31280,N_31338);
nor U31522 (N_31522,N_31168,N_31380);
xor U31523 (N_31523,N_31368,N_31438);
nand U31524 (N_31524,N_31454,N_31487);
and U31525 (N_31525,N_31320,N_31138);
nor U31526 (N_31526,N_31431,N_31022);
nand U31527 (N_31527,N_31445,N_31411);
nor U31528 (N_31528,N_31177,N_31028);
nor U31529 (N_31529,N_31467,N_31142);
xor U31530 (N_31530,N_31209,N_31316);
nand U31531 (N_31531,N_31155,N_31192);
nor U31532 (N_31532,N_31223,N_31275);
nand U31533 (N_31533,N_31392,N_31256);
and U31534 (N_31534,N_31214,N_31100);
nor U31535 (N_31535,N_31492,N_31371);
or U31536 (N_31536,N_31319,N_31171);
or U31537 (N_31537,N_31063,N_31482);
or U31538 (N_31538,N_31311,N_31437);
or U31539 (N_31539,N_31470,N_31023);
nor U31540 (N_31540,N_31087,N_31163);
or U31541 (N_31541,N_31469,N_31326);
nor U31542 (N_31542,N_31427,N_31309);
xnor U31543 (N_31543,N_31170,N_31194);
or U31544 (N_31544,N_31084,N_31211);
xor U31545 (N_31545,N_31354,N_31120);
and U31546 (N_31546,N_31439,N_31068);
and U31547 (N_31547,N_31342,N_31128);
nor U31548 (N_31548,N_31457,N_31201);
and U31549 (N_31549,N_31106,N_31304);
xnor U31550 (N_31550,N_31337,N_31139);
xor U31551 (N_31551,N_31294,N_31341);
and U31552 (N_31552,N_31244,N_31010);
xnor U31553 (N_31553,N_31390,N_31386);
or U31554 (N_31554,N_31261,N_31229);
and U31555 (N_31555,N_31164,N_31013);
xnor U31556 (N_31556,N_31019,N_31025);
or U31557 (N_31557,N_31406,N_31284);
xor U31558 (N_31558,N_31333,N_31388);
and U31559 (N_31559,N_31112,N_31357);
or U31560 (N_31560,N_31160,N_31331);
or U31561 (N_31561,N_31198,N_31286);
or U31562 (N_31562,N_31113,N_31169);
nand U31563 (N_31563,N_31373,N_31074);
nand U31564 (N_31564,N_31178,N_31082);
and U31565 (N_31565,N_31032,N_31024);
and U31566 (N_31566,N_31372,N_31064);
xnor U31567 (N_31567,N_31444,N_31058);
and U31568 (N_31568,N_31091,N_31292);
xnor U31569 (N_31569,N_31047,N_31257);
xnor U31570 (N_31570,N_31347,N_31196);
nor U31571 (N_31571,N_31026,N_31247);
nor U31572 (N_31572,N_31141,N_31015);
or U31573 (N_31573,N_31253,N_31402);
and U31574 (N_31574,N_31018,N_31409);
xnor U31575 (N_31575,N_31167,N_31179);
xor U31576 (N_31576,N_31491,N_31014);
and U31577 (N_31577,N_31393,N_31038);
nand U31578 (N_31578,N_31131,N_31246);
or U31579 (N_31579,N_31375,N_31345);
or U31580 (N_31580,N_31250,N_31274);
and U31581 (N_31581,N_31033,N_31465);
or U31582 (N_31582,N_31396,N_31374);
xnor U31583 (N_31583,N_31208,N_31416);
nand U31584 (N_31584,N_31453,N_31447);
xnor U31585 (N_31585,N_31363,N_31475);
nor U31586 (N_31586,N_31086,N_31003);
xnor U31587 (N_31587,N_31325,N_31387);
nand U31588 (N_31588,N_31340,N_31312);
nor U31589 (N_31589,N_31212,N_31401);
nor U31590 (N_31590,N_31166,N_31195);
nor U31591 (N_31591,N_31417,N_31350);
nand U31592 (N_31592,N_31135,N_31418);
nand U31593 (N_31593,N_31220,N_31059);
nand U31594 (N_31594,N_31185,N_31461);
and U31595 (N_31595,N_31381,N_31385);
xor U31596 (N_31596,N_31412,N_31152);
and U31597 (N_31597,N_31149,N_31148);
or U31598 (N_31598,N_31034,N_31323);
nor U31599 (N_31599,N_31012,N_31232);
xor U31600 (N_31600,N_31234,N_31156);
nor U31601 (N_31601,N_31425,N_31451);
or U31602 (N_31602,N_31165,N_31291);
and U31603 (N_31603,N_31419,N_31109);
nand U31604 (N_31604,N_31040,N_31186);
nand U31605 (N_31605,N_31389,N_31228);
or U31606 (N_31606,N_31313,N_31080);
nor U31607 (N_31607,N_31449,N_31490);
nor U31608 (N_31608,N_31426,N_31035);
xor U31609 (N_31609,N_31362,N_31207);
or U31610 (N_31610,N_31210,N_31036);
nor U31611 (N_31611,N_31495,N_31117);
nor U31612 (N_31612,N_31078,N_31352);
nor U31613 (N_31613,N_31162,N_31069);
nand U31614 (N_31614,N_31219,N_31233);
or U31615 (N_31615,N_31001,N_31030);
or U31616 (N_31616,N_31161,N_31130);
nand U31617 (N_31617,N_31090,N_31218);
nor U31618 (N_31618,N_31006,N_31039);
nand U31619 (N_31619,N_31029,N_31353);
nand U31620 (N_31620,N_31191,N_31182);
nand U31621 (N_31621,N_31187,N_31285);
and U31622 (N_31622,N_31305,N_31296);
and U31623 (N_31623,N_31098,N_31476);
or U31624 (N_31624,N_31369,N_31283);
nor U31625 (N_31625,N_31268,N_31093);
nand U31626 (N_31626,N_31355,N_31440);
xnor U31627 (N_31627,N_31073,N_31403);
xnor U31628 (N_31628,N_31277,N_31344);
and U31629 (N_31629,N_31299,N_31114);
and U31630 (N_31630,N_31293,N_31382);
xor U31631 (N_31631,N_31405,N_31377);
and U31632 (N_31632,N_31494,N_31053);
nand U31633 (N_31633,N_31263,N_31290);
nor U31634 (N_31634,N_31111,N_31222);
nor U31635 (N_31635,N_31298,N_31245);
nand U31636 (N_31636,N_31473,N_31395);
and U31637 (N_31637,N_31157,N_31000);
nand U31638 (N_31638,N_31240,N_31221);
xor U31639 (N_31639,N_31126,N_31251);
nor U31640 (N_31640,N_31276,N_31466);
nand U31641 (N_31641,N_31436,N_31486);
and U31642 (N_31642,N_31496,N_31151);
or U31643 (N_31643,N_31478,N_31349);
and U31644 (N_31644,N_31260,N_31376);
nand U31645 (N_31645,N_31154,N_31480);
and U31646 (N_31646,N_31088,N_31094);
or U31647 (N_31647,N_31455,N_31181);
nor U31648 (N_31648,N_31119,N_31230);
xor U31649 (N_31649,N_31332,N_31180);
or U31650 (N_31650,N_31358,N_31462);
xnor U31651 (N_31651,N_31007,N_31176);
nand U31652 (N_31652,N_31042,N_31242);
nand U31653 (N_31653,N_31122,N_31366);
xor U31654 (N_31654,N_31281,N_31190);
nand U31655 (N_31655,N_31485,N_31458);
and U31656 (N_31656,N_31021,N_31270);
and U31657 (N_31657,N_31370,N_31020);
nand U31658 (N_31658,N_31217,N_31471);
nor U31659 (N_31659,N_31150,N_31205);
or U31660 (N_31660,N_31061,N_31193);
nand U31661 (N_31661,N_31048,N_31173);
xor U31662 (N_31662,N_31045,N_31041);
nor U31663 (N_31663,N_31378,N_31062);
xnor U31664 (N_31664,N_31110,N_31011);
xor U31665 (N_31665,N_31289,N_31060);
xnor U31666 (N_31666,N_31364,N_31384);
xor U31667 (N_31667,N_31282,N_31129);
nor U31668 (N_31668,N_31479,N_31330);
and U31669 (N_31669,N_31423,N_31287);
xor U31670 (N_31670,N_31146,N_31055);
and U31671 (N_31671,N_31300,N_31089);
nor U31672 (N_31672,N_31224,N_31318);
and U31673 (N_31673,N_31079,N_31095);
nor U31674 (N_31674,N_31125,N_31057);
or U31675 (N_31675,N_31199,N_31066);
xnor U31676 (N_31676,N_31474,N_31327);
or U31677 (N_31677,N_31359,N_31065);
nor U31678 (N_31678,N_31351,N_31243);
nor U31679 (N_31679,N_31365,N_31124);
or U31680 (N_31680,N_31434,N_31050);
xor U31681 (N_31681,N_31254,N_31072);
nor U31682 (N_31682,N_31104,N_31056);
nand U31683 (N_31683,N_31203,N_31017);
nand U31684 (N_31684,N_31136,N_31031);
or U31685 (N_31685,N_31346,N_31428);
and U31686 (N_31686,N_31421,N_31481);
and U31687 (N_31687,N_31307,N_31407);
or U31688 (N_31688,N_31009,N_31408);
nand U31689 (N_31689,N_31259,N_31046);
or U31690 (N_31690,N_31202,N_31383);
nand U31691 (N_31691,N_31262,N_31398);
nand U31692 (N_31692,N_31255,N_31092);
or U31693 (N_31693,N_31052,N_31463);
or U31694 (N_31694,N_31241,N_31172);
nand U31695 (N_31695,N_31184,N_31394);
nand U31696 (N_31696,N_31442,N_31410);
nor U31697 (N_31697,N_31215,N_31400);
or U31698 (N_31698,N_31273,N_31239);
nand U31699 (N_31699,N_31483,N_31101);
or U31700 (N_31700,N_31004,N_31127);
nor U31701 (N_31701,N_31143,N_31070);
nor U31702 (N_31702,N_31301,N_31429);
nor U31703 (N_31703,N_31443,N_31140);
or U31704 (N_31704,N_31324,N_31189);
xnor U31705 (N_31705,N_31016,N_31448);
or U31706 (N_31706,N_31071,N_31269);
xor U31707 (N_31707,N_31204,N_31464);
nand U31708 (N_31708,N_31133,N_31308);
nor U31709 (N_31709,N_31484,N_31175);
nor U31710 (N_31710,N_31317,N_31134);
or U31711 (N_31711,N_31315,N_31302);
nand U31712 (N_31712,N_31252,N_31147);
nor U31713 (N_31713,N_31099,N_31226);
and U31714 (N_31714,N_31297,N_31348);
nor U31715 (N_31715,N_31336,N_31446);
nand U31716 (N_31716,N_31361,N_31213);
nor U31717 (N_31717,N_31121,N_31430);
nand U31718 (N_31718,N_31266,N_31096);
xnor U31719 (N_31719,N_31460,N_31328);
or U31720 (N_31720,N_31206,N_31153);
or U31721 (N_31721,N_31435,N_31037);
xnor U31722 (N_31722,N_31391,N_31267);
xor U31723 (N_31723,N_31235,N_31005);
or U31724 (N_31724,N_31216,N_31116);
nor U31725 (N_31725,N_31107,N_31002);
and U31726 (N_31726,N_31008,N_31145);
nor U31727 (N_31727,N_31265,N_31075);
nor U31728 (N_31728,N_31197,N_31103);
xnor U31729 (N_31729,N_31477,N_31472);
nand U31730 (N_31730,N_31422,N_31227);
nand U31731 (N_31731,N_31272,N_31271);
or U31732 (N_31732,N_31076,N_31343);
xnor U31733 (N_31733,N_31236,N_31132);
nor U31734 (N_31734,N_31237,N_31441);
nand U31735 (N_31735,N_31077,N_31027);
nor U31736 (N_31736,N_31044,N_31231);
xnor U31737 (N_31737,N_31310,N_31278);
and U31738 (N_31738,N_31321,N_31248);
and U31739 (N_31739,N_31102,N_31081);
nor U31740 (N_31740,N_31225,N_31054);
and U31741 (N_31741,N_31123,N_31258);
or U31742 (N_31742,N_31424,N_31183);
and U31743 (N_31743,N_31314,N_31115);
nand U31744 (N_31744,N_31137,N_31414);
nand U31745 (N_31745,N_31367,N_31499);
or U31746 (N_31746,N_31288,N_31334);
or U31747 (N_31747,N_31264,N_31399);
and U31748 (N_31748,N_31306,N_31339);
and U31749 (N_31749,N_31200,N_31335);
or U31750 (N_31750,N_31045,N_31419);
xor U31751 (N_31751,N_31295,N_31321);
or U31752 (N_31752,N_31213,N_31006);
and U31753 (N_31753,N_31090,N_31096);
xor U31754 (N_31754,N_31453,N_31049);
or U31755 (N_31755,N_31038,N_31427);
or U31756 (N_31756,N_31101,N_31211);
or U31757 (N_31757,N_31401,N_31448);
xor U31758 (N_31758,N_31340,N_31291);
or U31759 (N_31759,N_31478,N_31335);
nand U31760 (N_31760,N_31411,N_31087);
or U31761 (N_31761,N_31018,N_31187);
or U31762 (N_31762,N_31300,N_31396);
or U31763 (N_31763,N_31285,N_31329);
and U31764 (N_31764,N_31036,N_31426);
xnor U31765 (N_31765,N_31195,N_31432);
nor U31766 (N_31766,N_31450,N_31370);
or U31767 (N_31767,N_31101,N_31384);
xor U31768 (N_31768,N_31380,N_31085);
nand U31769 (N_31769,N_31178,N_31022);
xnor U31770 (N_31770,N_31417,N_31357);
nand U31771 (N_31771,N_31206,N_31158);
nor U31772 (N_31772,N_31048,N_31498);
and U31773 (N_31773,N_31112,N_31018);
nor U31774 (N_31774,N_31018,N_31067);
xnor U31775 (N_31775,N_31309,N_31421);
xnor U31776 (N_31776,N_31004,N_31044);
nor U31777 (N_31777,N_31454,N_31120);
nand U31778 (N_31778,N_31402,N_31026);
nor U31779 (N_31779,N_31465,N_31399);
nand U31780 (N_31780,N_31140,N_31035);
or U31781 (N_31781,N_31315,N_31329);
xnor U31782 (N_31782,N_31329,N_31239);
xnor U31783 (N_31783,N_31489,N_31068);
or U31784 (N_31784,N_31447,N_31470);
or U31785 (N_31785,N_31499,N_31144);
xor U31786 (N_31786,N_31067,N_31013);
or U31787 (N_31787,N_31015,N_31219);
or U31788 (N_31788,N_31415,N_31136);
and U31789 (N_31789,N_31329,N_31479);
or U31790 (N_31790,N_31352,N_31138);
or U31791 (N_31791,N_31494,N_31248);
nand U31792 (N_31792,N_31056,N_31481);
nor U31793 (N_31793,N_31221,N_31401);
and U31794 (N_31794,N_31105,N_31096);
nor U31795 (N_31795,N_31130,N_31008);
nor U31796 (N_31796,N_31019,N_31211);
nand U31797 (N_31797,N_31069,N_31059);
or U31798 (N_31798,N_31460,N_31117);
nand U31799 (N_31799,N_31464,N_31091);
nor U31800 (N_31800,N_31316,N_31360);
or U31801 (N_31801,N_31263,N_31001);
and U31802 (N_31802,N_31334,N_31020);
and U31803 (N_31803,N_31041,N_31039);
xnor U31804 (N_31804,N_31401,N_31022);
nand U31805 (N_31805,N_31012,N_31004);
xor U31806 (N_31806,N_31365,N_31011);
xnor U31807 (N_31807,N_31240,N_31330);
and U31808 (N_31808,N_31380,N_31265);
nand U31809 (N_31809,N_31075,N_31292);
and U31810 (N_31810,N_31374,N_31373);
or U31811 (N_31811,N_31317,N_31048);
and U31812 (N_31812,N_31228,N_31092);
and U31813 (N_31813,N_31351,N_31265);
or U31814 (N_31814,N_31183,N_31102);
nand U31815 (N_31815,N_31044,N_31093);
or U31816 (N_31816,N_31493,N_31013);
and U31817 (N_31817,N_31166,N_31094);
nor U31818 (N_31818,N_31288,N_31251);
xor U31819 (N_31819,N_31110,N_31347);
and U31820 (N_31820,N_31260,N_31168);
xor U31821 (N_31821,N_31108,N_31077);
xor U31822 (N_31822,N_31492,N_31073);
or U31823 (N_31823,N_31184,N_31206);
nand U31824 (N_31824,N_31336,N_31024);
xnor U31825 (N_31825,N_31327,N_31394);
nand U31826 (N_31826,N_31093,N_31454);
or U31827 (N_31827,N_31422,N_31397);
and U31828 (N_31828,N_31061,N_31117);
and U31829 (N_31829,N_31086,N_31315);
and U31830 (N_31830,N_31499,N_31340);
nor U31831 (N_31831,N_31335,N_31132);
and U31832 (N_31832,N_31311,N_31041);
or U31833 (N_31833,N_31060,N_31158);
or U31834 (N_31834,N_31033,N_31000);
xor U31835 (N_31835,N_31144,N_31023);
nor U31836 (N_31836,N_31002,N_31081);
and U31837 (N_31837,N_31026,N_31090);
nand U31838 (N_31838,N_31463,N_31435);
or U31839 (N_31839,N_31412,N_31172);
xor U31840 (N_31840,N_31424,N_31169);
nand U31841 (N_31841,N_31144,N_31435);
xor U31842 (N_31842,N_31403,N_31311);
nor U31843 (N_31843,N_31118,N_31198);
nor U31844 (N_31844,N_31427,N_31464);
and U31845 (N_31845,N_31122,N_31021);
nand U31846 (N_31846,N_31461,N_31102);
nor U31847 (N_31847,N_31286,N_31403);
or U31848 (N_31848,N_31184,N_31237);
nand U31849 (N_31849,N_31148,N_31208);
nor U31850 (N_31850,N_31302,N_31000);
xnor U31851 (N_31851,N_31488,N_31338);
nor U31852 (N_31852,N_31141,N_31264);
nor U31853 (N_31853,N_31182,N_31201);
or U31854 (N_31854,N_31494,N_31263);
xor U31855 (N_31855,N_31142,N_31209);
or U31856 (N_31856,N_31250,N_31103);
and U31857 (N_31857,N_31432,N_31065);
nand U31858 (N_31858,N_31478,N_31402);
nor U31859 (N_31859,N_31051,N_31022);
nand U31860 (N_31860,N_31258,N_31274);
nor U31861 (N_31861,N_31191,N_31188);
nand U31862 (N_31862,N_31332,N_31159);
and U31863 (N_31863,N_31177,N_31291);
and U31864 (N_31864,N_31131,N_31312);
xor U31865 (N_31865,N_31304,N_31208);
or U31866 (N_31866,N_31058,N_31247);
and U31867 (N_31867,N_31350,N_31378);
nand U31868 (N_31868,N_31057,N_31098);
nor U31869 (N_31869,N_31208,N_31158);
and U31870 (N_31870,N_31342,N_31012);
or U31871 (N_31871,N_31313,N_31483);
or U31872 (N_31872,N_31464,N_31169);
nand U31873 (N_31873,N_31165,N_31288);
and U31874 (N_31874,N_31239,N_31248);
or U31875 (N_31875,N_31473,N_31392);
or U31876 (N_31876,N_31424,N_31003);
xor U31877 (N_31877,N_31236,N_31142);
or U31878 (N_31878,N_31318,N_31124);
nor U31879 (N_31879,N_31376,N_31275);
nor U31880 (N_31880,N_31175,N_31070);
nor U31881 (N_31881,N_31422,N_31238);
or U31882 (N_31882,N_31160,N_31380);
or U31883 (N_31883,N_31283,N_31042);
or U31884 (N_31884,N_31207,N_31036);
or U31885 (N_31885,N_31087,N_31332);
nor U31886 (N_31886,N_31356,N_31389);
or U31887 (N_31887,N_31427,N_31416);
nor U31888 (N_31888,N_31270,N_31401);
or U31889 (N_31889,N_31048,N_31362);
nand U31890 (N_31890,N_31467,N_31200);
xnor U31891 (N_31891,N_31225,N_31395);
nor U31892 (N_31892,N_31140,N_31132);
nor U31893 (N_31893,N_31231,N_31043);
nand U31894 (N_31894,N_31090,N_31217);
nor U31895 (N_31895,N_31321,N_31356);
or U31896 (N_31896,N_31099,N_31493);
xnor U31897 (N_31897,N_31093,N_31289);
and U31898 (N_31898,N_31468,N_31480);
nand U31899 (N_31899,N_31430,N_31281);
and U31900 (N_31900,N_31436,N_31214);
xnor U31901 (N_31901,N_31213,N_31048);
xor U31902 (N_31902,N_31183,N_31258);
and U31903 (N_31903,N_31472,N_31442);
nand U31904 (N_31904,N_31109,N_31170);
or U31905 (N_31905,N_31184,N_31411);
and U31906 (N_31906,N_31067,N_31224);
nor U31907 (N_31907,N_31460,N_31355);
xnor U31908 (N_31908,N_31477,N_31359);
nor U31909 (N_31909,N_31363,N_31312);
or U31910 (N_31910,N_31304,N_31214);
nand U31911 (N_31911,N_31091,N_31008);
nand U31912 (N_31912,N_31282,N_31186);
or U31913 (N_31913,N_31138,N_31101);
xnor U31914 (N_31914,N_31256,N_31208);
nor U31915 (N_31915,N_31425,N_31156);
or U31916 (N_31916,N_31289,N_31094);
and U31917 (N_31917,N_31078,N_31458);
xor U31918 (N_31918,N_31494,N_31349);
and U31919 (N_31919,N_31422,N_31073);
nor U31920 (N_31920,N_31328,N_31386);
and U31921 (N_31921,N_31270,N_31476);
nor U31922 (N_31922,N_31362,N_31144);
nand U31923 (N_31923,N_31475,N_31248);
nor U31924 (N_31924,N_31410,N_31394);
nor U31925 (N_31925,N_31340,N_31102);
and U31926 (N_31926,N_31029,N_31022);
or U31927 (N_31927,N_31204,N_31425);
and U31928 (N_31928,N_31466,N_31450);
and U31929 (N_31929,N_31138,N_31076);
xor U31930 (N_31930,N_31181,N_31163);
nand U31931 (N_31931,N_31027,N_31246);
nor U31932 (N_31932,N_31078,N_31361);
nand U31933 (N_31933,N_31081,N_31464);
nor U31934 (N_31934,N_31377,N_31263);
nor U31935 (N_31935,N_31334,N_31265);
xnor U31936 (N_31936,N_31140,N_31052);
and U31937 (N_31937,N_31323,N_31274);
nor U31938 (N_31938,N_31417,N_31328);
nand U31939 (N_31939,N_31030,N_31118);
xnor U31940 (N_31940,N_31429,N_31207);
and U31941 (N_31941,N_31390,N_31041);
nand U31942 (N_31942,N_31263,N_31249);
xnor U31943 (N_31943,N_31147,N_31202);
or U31944 (N_31944,N_31495,N_31199);
and U31945 (N_31945,N_31214,N_31391);
xor U31946 (N_31946,N_31220,N_31029);
nor U31947 (N_31947,N_31111,N_31027);
nor U31948 (N_31948,N_31101,N_31495);
and U31949 (N_31949,N_31352,N_31297);
nor U31950 (N_31950,N_31065,N_31330);
xnor U31951 (N_31951,N_31381,N_31188);
xnor U31952 (N_31952,N_31407,N_31022);
nand U31953 (N_31953,N_31019,N_31307);
xnor U31954 (N_31954,N_31389,N_31272);
and U31955 (N_31955,N_31174,N_31277);
or U31956 (N_31956,N_31489,N_31017);
xor U31957 (N_31957,N_31300,N_31325);
and U31958 (N_31958,N_31160,N_31145);
nor U31959 (N_31959,N_31468,N_31274);
xor U31960 (N_31960,N_31220,N_31126);
or U31961 (N_31961,N_31279,N_31345);
or U31962 (N_31962,N_31125,N_31336);
xor U31963 (N_31963,N_31104,N_31464);
and U31964 (N_31964,N_31361,N_31433);
nor U31965 (N_31965,N_31001,N_31153);
and U31966 (N_31966,N_31294,N_31201);
nor U31967 (N_31967,N_31368,N_31493);
xnor U31968 (N_31968,N_31173,N_31252);
nand U31969 (N_31969,N_31401,N_31452);
nor U31970 (N_31970,N_31401,N_31425);
nand U31971 (N_31971,N_31201,N_31390);
and U31972 (N_31972,N_31075,N_31237);
and U31973 (N_31973,N_31319,N_31143);
nand U31974 (N_31974,N_31105,N_31021);
and U31975 (N_31975,N_31087,N_31043);
nand U31976 (N_31976,N_31050,N_31418);
and U31977 (N_31977,N_31415,N_31194);
nor U31978 (N_31978,N_31157,N_31136);
and U31979 (N_31979,N_31077,N_31356);
nand U31980 (N_31980,N_31392,N_31434);
and U31981 (N_31981,N_31353,N_31471);
nor U31982 (N_31982,N_31161,N_31122);
xor U31983 (N_31983,N_31415,N_31458);
xnor U31984 (N_31984,N_31363,N_31486);
nor U31985 (N_31985,N_31161,N_31181);
xnor U31986 (N_31986,N_31114,N_31307);
and U31987 (N_31987,N_31350,N_31473);
and U31988 (N_31988,N_31235,N_31003);
xor U31989 (N_31989,N_31499,N_31058);
nand U31990 (N_31990,N_31123,N_31214);
xor U31991 (N_31991,N_31072,N_31335);
xor U31992 (N_31992,N_31024,N_31320);
or U31993 (N_31993,N_31213,N_31016);
or U31994 (N_31994,N_31266,N_31083);
xnor U31995 (N_31995,N_31163,N_31462);
nor U31996 (N_31996,N_31435,N_31104);
and U31997 (N_31997,N_31466,N_31067);
and U31998 (N_31998,N_31463,N_31310);
and U31999 (N_31999,N_31188,N_31148);
xnor U32000 (N_32000,N_31806,N_31622);
nor U32001 (N_32001,N_31553,N_31973);
xnor U32002 (N_32002,N_31618,N_31508);
or U32003 (N_32003,N_31886,N_31936);
and U32004 (N_32004,N_31821,N_31650);
nand U32005 (N_32005,N_31891,N_31980);
xnor U32006 (N_32006,N_31981,N_31524);
nor U32007 (N_32007,N_31979,N_31772);
or U32008 (N_32008,N_31518,N_31827);
nand U32009 (N_32009,N_31581,N_31971);
and U32010 (N_32010,N_31710,N_31879);
nor U32011 (N_32011,N_31956,N_31968);
xor U32012 (N_32012,N_31900,N_31636);
and U32013 (N_32013,N_31609,N_31845);
nor U32014 (N_32014,N_31552,N_31637);
and U32015 (N_32015,N_31590,N_31959);
nor U32016 (N_32016,N_31627,N_31632);
or U32017 (N_32017,N_31847,N_31571);
nor U32018 (N_32018,N_31714,N_31987);
nand U32019 (N_32019,N_31967,N_31784);
nor U32020 (N_32020,N_31825,N_31512);
nor U32021 (N_32021,N_31507,N_31584);
nor U32022 (N_32022,N_31708,N_31801);
and U32023 (N_32023,N_31648,N_31659);
xor U32024 (N_32024,N_31942,N_31573);
xor U32025 (N_32025,N_31565,N_31539);
and U32026 (N_32026,N_31780,N_31820);
nand U32027 (N_32027,N_31616,N_31591);
and U32028 (N_32028,N_31997,N_31547);
nand U32029 (N_32029,N_31846,N_31850);
xnor U32030 (N_32030,N_31765,N_31944);
and U32031 (N_32031,N_31652,N_31791);
and U32032 (N_32032,N_31540,N_31705);
nor U32033 (N_32033,N_31727,N_31505);
xnor U32034 (N_32034,N_31937,N_31826);
xor U32035 (N_32035,N_31841,N_31985);
xnor U32036 (N_32036,N_31729,N_31624);
nand U32037 (N_32037,N_31865,N_31773);
or U32038 (N_32038,N_31905,N_31645);
xor U32039 (N_32039,N_31572,N_31833);
nand U32040 (N_32040,N_31692,N_31556);
xnor U32041 (N_32041,N_31520,N_31864);
nand U32042 (N_32042,N_31930,N_31809);
xor U32043 (N_32043,N_31974,N_31764);
nand U32044 (N_32044,N_31906,N_31661);
or U32045 (N_32045,N_31576,N_31603);
and U32046 (N_32046,N_31851,N_31739);
nor U32047 (N_32047,N_31802,N_31824);
nor U32048 (N_32048,N_31588,N_31882);
xor U32049 (N_32049,N_31875,N_31689);
or U32050 (N_32050,N_31907,N_31711);
nor U32051 (N_32051,N_31874,N_31760);
nand U32052 (N_32052,N_31702,N_31940);
nand U32053 (N_32053,N_31790,N_31678);
or U32054 (N_32054,N_31917,N_31545);
nor U32055 (N_32055,N_31675,N_31725);
xnor U32056 (N_32056,N_31561,N_31863);
xor U32057 (N_32057,N_31889,N_31988);
xor U32058 (N_32058,N_31894,N_31876);
or U32059 (N_32059,N_31928,N_31789);
nor U32060 (N_32060,N_31738,N_31862);
or U32061 (N_32061,N_31615,N_31911);
xnor U32062 (N_32062,N_31696,N_31792);
nand U32063 (N_32063,N_31671,N_31803);
nand U32064 (N_32064,N_31502,N_31883);
nor U32065 (N_32065,N_31946,N_31963);
nor U32066 (N_32066,N_31952,N_31606);
and U32067 (N_32067,N_31933,N_31795);
and U32068 (N_32068,N_31690,N_31969);
or U32069 (N_32069,N_31608,N_31643);
and U32070 (N_32070,N_31728,N_31901);
nor U32071 (N_32071,N_31677,N_31631);
nor U32072 (N_32072,N_31517,N_31617);
xnor U32073 (N_32073,N_31630,N_31830);
nand U32074 (N_32074,N_31595,N_31756);
nor U32075 (N_32075,N_31686,N_31994);
nand U32076 (N_32076,N_31807,N_31674);
and U32077 (N_32077,N_31888,N_31966);
and U32078 (N_32078,N_31713,N_31818);
nand U32079 (N_32079,N_31965,N_31817);
and U32080 (N_32080,N_31550,N_31515);
or U32081 (N_32081,N_31812,N_31915);
nor U32082 (N_32082,N_31746,N_31744);
or U32083 (N_32083,N_31724,N_31787);
nor U32084 (N_32084,N_31771,N_31877);
nor U32085 (N_32085,N_31599,N_31899);
nand U32086 (N_32086,N_31623,N_31684);
nor U32087 (N_32087,N_31610,N_31885);
or U32088 (N_32088,N_31737,N_31511);
xor U32089 (N_32089,N_31526,N_31945);
or U32090 (N_32090,N_31558,N_31555);
nand U32091 (N_32091,N_31621,N_31852);
xor U32092 (N_32092,N_31527,N_31763);
or U32093 (N_32093,N_31909,N_31908);
xor U32094 (N_32094,N_31913,N_31996);
or U32095 (N_32095,N_31860,N_31823);
nand U32096 (N_32096,N_31958,N_31878);
or U32097 (N_32097,N_31694,N_31680);
nor U32098 (N_32098,N_31866,N_31718);
and U32099 (N_32099,N_31836,N_31605);
nor U32100 (N_32100,N_31881,N_31897);
and U32101 (N_32101,N_31676,N_31574);
and U32102 (N_32102,N_31948,N_31983);
nor U32103 (N_32103,N_31734,N_31687);
and U32104 (N_32104,N_31612,N_31951);
xor U32105 (N_32105,N_31730,N_31649);
and U32106 (N_32106,N_31736,N_31720);
or U32107 (N_32107,N_31794,N_31740);
xnor U32108 (N_32108,N_31964,N_31761);
nor U32109 (N_32109,N_31577,N_31538);
xor U32110 (N_32110,N_31642,N_31626);
nand U32111 (N_32111,N_31854,N_31837);
and U32112 (N_32112,N_31619,N_31567);
xnor U32113 (N_32113,N_31819,N_31814);
or U32114 (N_32114,N_31660,N_31586);
nor U32115 (N_32115,N_31990,N_31667);
xnor U32116 (N_32116,N_31788,N_31566);
nor U32117 (N_32117,N_31949,N_31564);
or U32118 (N_32118,N_31731,N_31775);
nor U32119 (N_32119,N_31954,N_31717);
xnor U32120 (N_32120,N_31651,N_31604);
nand U32121 (N_32121,N_31976,N_31726);
and U32122 (N_32122,N_31562,N_31848);
nor U32123 (N_32123,N_31554,N_31849);
nor U32124 (N_32124,N_31840,N_31750);
nor U32125 (N_32125,N_31961,N_31892);
nand U32126 (N_32126,N_31743,N_31781);
xor U32127 (N_32127,N_31793,N_31835);
nand U32128 (N_32128,N_31890,N_31665);
nand U32129 (N_32129,N_31931,N_31898);
and U32130 (N_32130,N_31785,N_31646);
and U32131 (N_32131,N_31919,N_31504);
or U32132 (N_32132,N_31842,N_31950);
xor U32133 (N_32133,N_31872,N_31868);
nor U32134 (N_32134,N_31658,N_31767);
and U32135 (N_32135,N_31685,N_31777);
and U32136 (N_32136,N_31568,N_31706);
xor U32137 (N_32137,N_31597,N_31681);
nand U32138 (N_32138,N_31844,N_31559);
nor U32139 (N_32139,N_31880,N_31509);
nand U32140 (N_32140,N_31927,N_31786);
and U32141 (N_32141,N_31815,N_31531);
xnor U32142 (N_32142,N_31633,N_31939);
nor U32143 (N_32143,N_31669,N_31871);
nor U32144 (N_32144,N_31516,N_31867);
or U32145 (N_32145,N_31839,N_31857);
or U32146 (N_32146,N_31923,N_31861);
nor U32147 (N_32147,N_31977,N_31758);
or U32148 (N_32148,N_31639,N_31719);
and U32149 (N_32149,N_31747,N_31647);
and U32150 (N_32150,N_31783,N_31741);
xor U32151 (N_32151,N_31856,N_31598);
nand U32152 (N_32152,N_31592,N_31989);
xnor U32153 (N_32153,N_31766,N_31549);
or U32154 (N_32154,N_31722,N_31723);
nand U32155 (N_32155,N_31672,N_31869);
xnor U32156 (N_32156,N_31635,N_31542);
nor U32157 (N_32157,N_31699,N_31955);
and U32158 (N_32158,N_31528,N_31770);
nor U32159 (N_32159,N_31514,N_31838);
or U32160 (N_32160,N_31829,N_31522);
nand U32161 (N_32161,N_31932,N_31691);
or U32162 (N_32162,N_31887,N_31916);
nand U32163 (N_32163,N_31769,N_31808);
nor U32164 (N_32164,N_31828,N_31593);
nor U32165 (N_32165,N_31701,N_31804);
nor U32166 (N_32166,N_31715,N_31924);
nor U32167 (N_32167,N_31926,N_31503);
xnor U32168 (N_32168,N_31904,N_31798);
nor U32169 (N_32169,N_31557,N_31653);
xor U32170 (N_32170,N_31858,N_31533);
or U32171 (N_32171,N_31682,N_31934);
nand U32172 (N_32172,N_31662,N_31935);
xor U32173 (N_32173,N_31752,N_31683);
xnor U32174 (N_32174,N_31853,N_31941);
nand U32175 (N_32175,N_31673,N_31986);
and U32176 (N_32176,N_31978,N_31800);
or U32177 (N_32177,N_31768,N_31563);
or U32178 (N_32178,N_31938,N_31500);
nand U32179 (N_32179,N_31700,N_31580);
or U32180 (N_32180,N_31628,N_31704);
xnor U32181 (N_32181,N_31991,N_31668);
and U32182 (N_32182,N_31534,N_31745);
nand U32183 (N_32183,N_31543,N_31733);
xor U32184 (N_32184,N_31596,N_31957);
xor U32185 (N_32185,N_31776,N_31920);
nor U32186 (N_32186,N_31697,N_31918);
nand U32187 (N_32187,N_31501,N_31754);
xor U32188 (N_32188,N_31703,N_31896);
xor U32189 (N_32189,N_31510,N_31721);
or U32190 (N_32190,N_31585,N_31583);
xnor U32191 (N_32191,N_31984,N_31893);
or U32192 (N_32192,N_31993,N_31902);
and U32193 (N_32193,N_31587,N_31634);
nor U32194 (N_32194,N_31921,N_31999);
nor U32195 (N_32195,N_31578,N_31855);
or U32196 (N_32196,N_31629,N_31748);
or U32197 (N_32197,N_31607,N_31873);
xnor U32198 (N_32198,N_31625,N_31641);
nor U32199 (N_32199,N_31654,N_31903);
xor U32200 (N_32200,N_31749,N_31506);
and U32201 (N_32201,N_31589,N_31600);
nor U32202 (N_32202,N_31929,N_31755);
nand U32203 (N_32203,N_31666,N_31813);
and U32204 (N_32204,N_31614,N_31947);
or U32205 (N_32205,N_31638,N_31742);
and U32206 (N_32206,N_31620,N_31611);
xnor U32207 (N_32207,N_31799,N_31640);
nand U32208 (N_32208,N_31693,N_31536);
nor U32209 (N_32209,N_31695,N_31805);
or U32210 (N_32210,N_31762,N_31655);
nor U32211 (N_32211,N_31779,N_31822);
xor U32212 (N_32212,N_31521,N_31560);
nand U32213 (N_32213,N_31796,N_31912);
nand U32214 (N_32214,N_31569,N_31656);
and U32215 (N_32215,N_31532,N_31816);
nor U32216 (N_32216,N_31759,N_31782);
nand U32217 (N_32217,N_31753,N_31688);
xor U32218 (N_32218,N_31834,N_31582);
xor U32219 (N_32219,N_31698,N_31757);
and U32220 (N_32220,N_31709,N_31972);
nor U32221 (N_32221,N_31870,N_31519);
xor U32222 (N_32222,N_31679,N_31910);
or U32223 (N_32223,N_31998,N_31570);
nor U32224 (N_32224,N_31975,N_31579);
xor U32225 (N_32225,N_31970,N_31541);
xor U32226 (N_32226,N_31712,N_31523);
xor U32227 (N_32227,N_31657,N_31884);
or U32228 (N_32228,N_31513,N_31962);
or U32229 (N_32229,N_31811,N_31735);
or U32230 (N_32230,N_31832,N_31925);
nand U32231 (N_32231,N_31895,N_31914);
and U32232 (N_32232,N_31774,N_31575);
xnor U32233 (N_32233,N_31732,N_31810);
nor U32234 (N_32234,N_31594,N_31644);
nand U32235 (N_32235,N_31664,N_31544);
xnor U32236 (N_32236,N_31953,N_31663);
nor U32237 (N_32237,N_31602,N_31751);
xor U32238 (N_32238,N_31992,N_31670);
xor U32239 (N_32239,N_31551,N_31982);
xnor U32240 (N_32240,N_31859,N_31546);
nand U32241 (N_32241,N_31548,N_31537);
and U32242 (N_32242,N_31716,N_31797);
nand U32243 (N_32243,N_31530,N_31778);
nand U32244 (N_32244,N_31601,N_31843);
xor U32245 (N_32245,N_31831,N_31529);
xnor U32246 (N_32246,N_31707,N_31960);
and U32247 (N_32247,N_31995,N_31943);
nor U32248 (N_32248,N_31922,N_31613);
nor U32249 (N_32249,N_31525,N_31535);
nor U32250 (N_32250,N_31552,N_31995);
xor U32251 (N_32251,N_31854,N_31610);
and U32252 (N_32252,N_31828,N_31915);
or U32253 (N_32253,N_31735,N_31730);
and U32254 (N_32254,N_31652,N_31750);
xor U32255 (N_32255,N_31832,N_31506);
xnor U32256 (N_32256,N_31908,N_31820);
and U32257 (N_32257,N_31973,N_31546);
or U32258 (N_32258,N_31544,N_31966);
xor U32259 (N_32259,N_31743,N_31653);
nand U32260 (N_32260,N_31598,N_31978);
nor U32261 (N_32261,N_31766,N_31648);
or U32262 (N_32262,N_31864,N_31975);
or U32263 (N_32263,N_31751,N_31515);
nand U32264 (N_32264,N_31871,N_31704);
and U32265 (N_32265,N_31970,N_31514);
or U32266 (N_32266,N_31948,N_31794);
or U32267 (N_32267,N_31951,N_31731);
nand U32268 (N_32268,N_31712,N_31567);
and U32269 (N_32269,N_31921,N_31926);
and U32270 (N_32270,N_31578,N_31651);
nor U32271 (N_32271,N_31933,N_31855);
xor U32272 (N_32272,N_31737,N_31689);
nand U32273 (N_32273,N_31915,N_31738);
or U32274 (N_32274,N_31637,N_31923);
or U32275 (N_32275,N_31954,N_31752);
nor U32276 (N_32276,N_31587,N_31776);
or U32277 (N_32277,N_31878,N_31763);
and U32278 (N_32278,N_31970,N_31911);
nor U32279 (N_32279,N_31838,N_31783);
and U32280 (N_32280,N_31987,N_31717);
and U32281 (N_32281,N_31602,N_31637);
nor U32282 (N_32282,N_31513,N_31656);
or U32283 (N_32283,N_31917,N_31998);
nand U32284 (N_32284,N_31586,N_31644);
and U32285 (N_32285,N_31977,N_31837);
xnor U32286 (N_32286,N_31572,N_31916);
and U32287 (N_32287,N_31657,N_31660);
or U32288 (N_32288,N_31931,N_31663);
nand U32289 (N_32289,N_31555,N_31734);
and U32290 (N_32290,N_31597,N_31972);
xnor U32291 (N_32291,N_31704,N_31817);
xor U32292 (N_32292,N_31570,N_31653);
or U32293 (N_32293,N_31802,N_31768);
and U32294 (N_32294,N_31771,N_31800);
nor U32295 (N_32295,N_31645,N_31644);
nand U32296 (N_32296,N_31561,N_31879);
nand U32297 (N_32297,N_31560,N_31713);
xor U32298 (N_32298,N_31582,N_31669);
xnor U32299 (N_32299,N_31578,N_31588);
xor U32300 (N_32300,N_31994,N_31947);
and U32301 (N_32301,N_31587,N_31757);
nand U32302 (N_32302,N_31722,N_31951);
and U32303 (N_32303,N_31610,N_31946);
nor U32304 (N_32304,N_31897,N_31777);
nor U32305 (N_32305,N_31931,N_31583);
xnor U32306 (N_32306,N_31765,N_31561);
nor U32307 (N_32307,N_31764,N_31852);
nor U32308 (N_32308,N_31691,N_31870);
xnor U32309 (N_32309,N_31963,N_31596);
xnor U32310 (N_32310,N_31817,N_31520);
xnor U32311 (N_32311,N_31590,N_31628);
or U32312 (N_32312,N_31881,N_31723);
nor U32313 (N_32313,N_31747,N_31653);
xnor U32314 (N_32314,N_31580,N_31639);
xor U32315 (N_32315,N_31552,N_31660);
and U32316 (N_32316,N_31736,N_31768);
nand U32317 (N_32317,N_31932,N_31950);
xnor U32318 (N_32318,N_31973,N_31997);
nand U32319 (N_32319,N_31970,N_31609);
and U32320 (N_32320,N_31849,N_31698);
nor U32321 (N_32321,N_31689,N_31987);
xnor U32322 (N_32322,N_31641,N_31972);
xnor U32323 (N_32323,N_31986,N_31744);
and U32324 (N_32324,N_31759,N_31676);
and U32325 (N_32325,N_31557,N_31715);
nand U32326 (N_32326,N_31559,N_31823);
nand U32327 (N_32327,N_31772,N_31904);
nor U32328 (N_32328,N_31863,N_31737);
xnor U32329 (N_32329,N_31967,N_31746);
nor U32330 (N_32330,N_31996,N_31786);
or U32331 (N_32331,N_31608,N_31509);
nor U32332 (N_32332,N_31984,N_31785);
or U32333 (N_32333,N_31557,N_31624);
nor U32334 (N_32334,N_31562,N_31940);
nand U32335 (N_32335,N_31502,N_31578);
and U32336 (N_32336,N_31939,N_31881);
and U32337 (N_32337,N_31519,N_31840);
or U32338 (N_32338,N_31612,N_31565);
xnor U32339 (N_32339,N_31655,N_31787);
xor U32340 (N_32340,N_31964,N_31898);
or U32341 (N_32341,N_31741,N_31975);
xor U32342 (N_32342,N_31886,N_31856);
and U32343 (N_32343,N_31954,N_31730);
nor U32344 (N_32344,N_31923,N_31992);
xnor U32345 (N_32345,N_31584,N_31649);
and U32346 (N_32346,N_31553,N_31763);
nor U32347 (N_32347,N_31997,N_31819);
xor U32348 (N_32348,N_31774,N_31615);
nor U32349 (N_32349,N_31841,N_31612);
nand U32350 (N_32350,N_31684,N_31993);
nand U32351 (N_32351,N_31875,N_31572);
and U32352 (N_32352,N_31694,N_31544);
nor U32353 (N_32353,N_31734,N_31851);
and U32354 (N_32354,N_31645,N_31565);
nand U32355 (N_32355,N_31887,N_31818);
and U32356 (N_32356,N_31835,N_31758);
nor U32357 (N_32357,N_31664,N_31578);
xor U32358 (N_32358,N_31782,N_31554);
nor U32359 (N_32359,N_31536,N_31576);
xnor U32360 (N_32360,N_31571,N_31827);
nand U32361 (N_32361,N_31652,N_31816);
nor U32362 (N_32362,N_31955,N_31618);
nand U32363 (N_32363,N_31741,N_31757);
nor U32364 (N_32364,N_31736,N_31729);
or U32365 (N_32365,N_31735,N_31867);
xor U32366 (N_32366,N_31922,N_31818);
xor U32367 (N_32367,N_31891,N_31976);
and U32368 (N_32368,N_31827,N_31778);
and U32369 (N_32369,N_31731,N_31844);
xnor U32370 (N_32370,N_31535,N_31898);
xnor U32371 (N_32371,N_31899,N_31762);
and U32372 (N_32372,N_31595,N_31893);
or U32373 (N_32373,N_31741,N_31920);
nand U32374 (N_32374,N_31603,N_31524);
or U32375 (N_32375,N_31668,N_31815);
or U32376 (N_32376,N_31652,N_31899);
and U32377 (N_32377,N_31987,N_31544);
xnor U32378 (N_32378,N_31640,N_31688);
xnor U32379 (N_32379,N_31919,N_31865);
nor U32380 (N_32380,N_31711,N_31637);
and U32381 (N_32381,N_31912,N_31576);
or U32382 (N_32382,N_31718,N_31902);
xor U32383 (N_32383,N_31887,N_31695);
and U32384 (N_32384,N_31769,N_31552);
nor U32385 (N_32385,N_31873,N_31535);
or U32386 (N_32386,N_31786,N_31504);
nand U32387 (N_32387,N_31691,N_31911);
and U32388 (N_32388,N_31968,N_31630);
nand U32389 (N_32389,N_31505,N_31938);
nor U32390 (N_32390,N_31560,N_31755);
and U32391 (N_32391,N_31679,N_31531);
or U32392 (N_32392,N_31991,N_31861);
nor U32393 (N_32393,N_31568,N_31842);
nor U32394 (N_32394,N_31646,N_31922);
nand U32395 (N_32395,N_31706,N_31729);
nor U32396 (N_32396,N_31676,N_31598);
and U32397 (N_32397,N_31940,N_31861);
and U32398 (N_32398,N_31598,N_31666);
xor U32399 (N_32399,N_31608,N_31826);
nand U32400 (N_32400,N_31863,N_31703);
nor U32401 (N_32401,N_31576,N_31881);
or U32402 (N_32402,N_31614,N_31595);
nor U32403 (N_32403,N_31813,N_31762);
and U32404 (N_32404,N_31547,N_31813);
xnor U32405 (N_32405,N_31949,N_31838);
xor U32406 (N_32406,N_31553,N_31953);
nor U32407 (N_32407,N_31822,N_31920);
and U32408 (N_32408,N_31993,N_31700);
or U32409 (N_32409,N_31917,N_31506);
nand U32410 (N_32410,N_31820,N_31815);
and U32411 (N_32411,N_31769,N_31560);
nand U32412 (N_32412,N_31879,N_31698);
or U32413 (N_32413,N_31664,N_31629);
xor U32414 (N_32414,N_31556,N_31736);
and U32415 (N_32415,N_31760,N_31664);
nand U32416 (N_32416,N_31569,N_31787);
nor U32417 (N_32417,N_31797,N_31859);
nor U32418 (N_32418,N_31516,N_31529);
nor U32419 (N_32419,N_31861,N_31794);
nor U32420 (N_32420,N_31551,N_31552);
nand U32421 (N_32421,N_31655,N_31952);
nand U32422 (N_32422,N_31756,N_31729);
nand U32423 (N_32423,N_31503,N_31999);
or U32424 (N_32424,N_31550,N_31990);
or U32425 (N_32425,N_31804,N_31875);
xnor U32426 (N_32426,N_31712,N_31667);
xor U32427 (N_32427,N_31909,N_31638);
xnor U32428 (N_32428,N_31874,N_31957);
nor U32429 (N_32429,N_31882,N_31608);
or U32430 (N_32430,N_31664,N_31654);
nor U32431 (N_32431,N_31796,N_31819);
nand U32432 (N_32432,N_31750,N_31751);
nor U32433 (N_32433,N_31500,N_31954);
xor U32434 (N_32434,N_31508,N_31806);
nand U32435 (N_32435,N_31857,N_31736);
nor U32436 (N_32436,N_31900,N_31901);
nand U32437 (N_32437,N_31526,N_31620);
nand U32438 (N_32438,N_31783,N_31563);
or U32439 (N_32439,N_31813,N_31968);
and U32440 (N_32440,N_31818,N_31522);
and U32441 (N_32441,N_31709,N_31813);
and U32442 (N_32442,N_31902,N_31517);
nand U32443 (N_32443,N_31897,N_31820);
xnor U32444 (N_32444,N_31907,N_31686);
xnor U32445 (N_32445,N_31835,N_31964);
and U32446 (N_32446,N_31950,N_31891);
nor U32447 (N_32447,N_31585,N_31824);
xnor U32448 (N_32448,N_31876,N_31968);
and U32449 (N_32449,N_31789,N_31755);
or U32450 (N_32450,N_31809,N_31925);
and U32451 (N_32451,N_31983,N_31708);
and U32452 (N_32452,N_31762,N_31722);
or U32453 (N_32453,N_31595,N_31655);
nand U32454 (N_32454,N_31770,N_31821);
nor U32455 (N_32455,N_31955,N_31646);
nor U32456 (N_32456,N_31939,N_31522);
nand U32457 (N_32457,N_31893,N_31754);
or U32458 (N_32458,N_31713,N_31619);
and U32459 (N_32459,N_31865,N_31530);
or U32460 (N_32460,N_31795,N_31861);
or U32461 (N_32461,N_31799,N_31829);
nor U32462 (N_32462,N_31615,N_31866);
nor U32463 (N_32463,N_31698,N_31960);
or U32464 (N_32464,N_31812,N_31767);
nand U32465 (N_32465,N_31999,N_31559);
nand U32466 (N_32466,N_31574,N_31628);
or U32467 (N_32467,N_31583,N_31521);
and U32468 (N_32468,N_31972,N_31998);
or U32469 (N_32469,N_31629,N_31997);
nor U32470 (N_32470,N_31789,N_31997);
or U32471 (N_32471,N_31966,N_31501);
and U32472 (N_32472,N_31595,N_31994);
or U32473 (N_32473,N_31507,N_31655);
xor U32474 (N_32474,N_31872,N_31751);
and U32475 (N_32475,N_31767,N_31648);
xnor U32476 (N_32476,N_31992,N_31772);
xnor U32477 (N_32477,N_31549,N_31914);
nor U32478 (N_32478,N_31926,N_31502);
nand U32479 (N_32479,N_31692,N_31539);
nand U32480 (N_32480,N_31838,N_31773);
nor U32481 (N_32481,N_31538,N_31788);
nor U32482 (N_32482,N_31788,N_31526);
or U32483 (N_32483,N_31737,N_31566);
nand U32484 (N_32484,N_31715,N_31587);
xnor U32485 (N_32485,N_31729,N_31950);
nor U32486 (N_32486,N_31960,N_31920);
xor U32487 (N_32487,N_31667,N_31593);
nor U32488 (N_32488,N_31798,N_31899);
xor U32489 (N_32489,N_31634,N_31531);
and U32490 (N_32490,N_31580,N_31584);
nand U32491 (N_32491,N_31644,N_31895);
and U32492 (N_32492,N_31989,N_31605);
xor U32493 (N_32493,N_31807,N_31683);
nor U32494 (N_32494,N_31556,N_31715);
and U32495 (N_32495,N_31897,N_31602);
nand U32496 (N_32496,N_31653,N_31962);
nor U32497 (N_32497,N_31844,N_31993);
or U32498 (N_32498,N_31989,N_31688);
nor U32499 (N_32499,N_31827,N_31710);
nand U32500 (N_32500,N_32065,N_32230);
nand U32501 (N_32501,N_32344,N_32140);
nor U32502 (N_32502,N_32089,N_32010);
and U32503 (N_32503,N_32396,N_32057);
nand U32504 (N_32504,N_32478,N_32496);
nand U32505 (N_32505,N_32136,N_32406);
nor U32506 (N_32506,N_32076,N_32143);
and U32507 (N_32507,N_32146,N_32129);
nand U32508 (N_32508,N_32167,N_32159);
and U32509 (N_32509,N_32062,N_32055);
and U32510 (N_32510,N_32228,N_32108);
xnor U32511 (N_32511,N_32234,N_32451);
and U32512 (N_32512,N_32053,N_32186);
nor U32513 (N_32513,N_32027,N_32215);
xor U32514 (N_32514,N_32123,N_32029);
or U32515 (N_32515,N_32270,N_32105);
nor U32516 (N_32516,N_32034,N_32403);
nor U32517 (N_32517,N_32154,N_32480);
or U32518 (N_32518,N_32364,N_32144);
nand U32519 (N_32519,N_32350,N_32329);
nor U32520 (N_32520,N_32286,N_32210);
xnor U32521 (N_32521,N_32173,N_32223);
or U32522 (N_32522,N_32420,N_32443);
and U32523 (N_32523,N_32033,N_32337);
nor U32524 (N_32524,N_32224,N_32128);
nor U32525 (N_32525,N_32067,N_32229);
nor U32526 (N_32526,N_32479,N_32375);
nor U32527 (N_32527,N_32149,N_32362);
xnor U32528 (N_32528,N_32139,N_32115);
and U32529 (N_32529,N_32411,N_32259);
xor U32530 (N_32530,N_32104,N_32485);
nand U32531 (N_32531,N_32384,N_32371);
or U32532 (N_32532,N_32110,N_32388);
and U32533 (N_32533,N_32390,N_32241);
xor U32534 (N_32534,N_32491,N_32473);
nand U32535 (N_32535,N_32386,N_32111);
or U32536 (N_32536,N_32185,N_32310);
or U32537 (N_32537,N_32077,N_32037);
and U32538 (N_32538,N_32025,N_32194);
nor U32539 (N_32539,N_32081,N_32145);
and U32540 (N_32540,N_32488,N_32410);
xnor U32541 (N_32541,N_32045,N_32263);
xor U32542 (N_32542,N_32351,N_32097);
nand U32543 (N_32543,N_32002,N_32465);
xor U32544 (N_32544,N_32417,N_32486);
nor U32545 (N_32545,N_32213,N_32178);
xor U32546 (N_32546,N_32214,N_32013);
xor U32547 (N_32547,N_32205,N_32005);
nand U32548 (N_32548,N_32138,N_32031);
and U32549 (N_32549,N_32369,N_32078);
nor U32550 (N_32550,N_32352,N_32211);
and U32551 (N_32551,N_32304,N_32357);
and U32552 (N_32552,N_32152,N_32343);
nand U32553 (N_32553,N_32012,N_32462);
or U32554 (N_32554,N_32428,N_32006);
or U32555 (N_32555,N_32358,N_32481);
nand U32556 (N_32556,N_32319,N_32269);
nand U32557 (N_32557,N_32107,N_32294);
nand U32558 (N_32558,N_32445,N_32400);
nor U32559 (N_32559,N_32436,N_32249);
nor U32560 (N_32560,N_32376,N_32256);
or U32561 (N_32561,N_32096,N_32168);
nand U32562 (N_32562,N_32426,N_32166);
nor U32563 (N_32563,N_32233,N_32477);
nand U32564 (N_32564,N_32268,N_32074);
nor U32565 (N_32565,N_32300,N_32433);
nand U32566 (N_32566,N_32121,N_32299);
and U32567 (N_32567,N_32165,N_32289);
xor U32568 (N_32568,N_32274,N_32177);
xnor U32569 (N_32569,N_32209,N_32278);
nand U32570 (N_32570,N_32212,N_32174);
nand U32571 (N_32571,N_32306,N_32463);
nor U32572 (N_32572,N_32418,N_32322);
nor U32573 (N_32573,N_32125,N_32349);
and U32574 (N_32574,N_32252,N_32320);
nand U32575 (N_32575,N_32079,N_32151);
nor U32576 (N_32576,N_32179,N_32456);
nor U32577 (N_32577,N_32007,N_32216);
nor U32578 (N_32578,N_32372,N_32338);
nand U32579 (N_32579,N_32469,N_32137);
xor U32580 (N_32580,N_32244,N_32100);
nor U32581 (N_32581,N_32356,N_32460);
and U32582 (N_32582,N_32226,N_32247);
and U32583 (N_32583,N_32328,N_32448);
nor U32584 (N_32584,N_32391,N_32271);
nor U32585 (N_32585,N_32492,N_32172);
and U32586 (N_32586,N_32240,N_32370);
xnor U32587 (N_32587,N_32109,N_32028);
or U32588 (N_32588,N_32208,N_32225);
nand U32589 (N_32589,N_32093,N_32133);
xor U32590 (N_32590,N_32346,N_32302);
nor U32591 (N_32591,N_32219,N_32325);
nor U32592 (N_32592,N_32001,N_32222);
nand U32593 (N_32593,N_32412,N_32307);
or U32594 (N_32594,N_32316,N_32251);
nor U32595 (N_32595,N_32475,N_32071);
nand U32596 (N_32596,N_32347,N_32373);
nand U32597 (N_32597,N_32085,N_32378);
nor U32598 (N_32598,N_32311,N_32439);
nor U32599 (N_32599,N_32336,N_32155);
nand U32600 (N_32600,N_32361,N_32287);
or U32601 (N_32601,N_32455,N_32339);
or U32602 (N_32602,N_32308,N_32374);
xor U32603 (N_32603,N_32392,N_32323);
nor U32604 (N_32604,N_32267,N_32070);
nor U32605 (N_32605,N_32206,N_32314);
or U32606 (N_32606,N_32203,N_32243);
nand U32607 (N_32607,N_32056,N_32345);
and U32608 (N_32608,N_32068,N_32430);
and U32609 (N_32609,N_32359,N_32353);
nand U32610 (N_32610,N_32472,N_32080);
and U32611 (N_32611,N_32232,N_32094);
nor U32612 (N_32612,N_32360,N_32072);
nor U32613 (N_32613,N_32116,N_32134);
and U32614 (N_32614,N_32266,N_32497);
or U32615 (N_32615,N_32444,N_32262);
nand U32616 (N_32616,N_32471,N_32021);
nand U32617 (N_32617,N_32091,N_32237);
or U32618 (N_32618,N_32126,N_32181);
xnor U32619 (N_32619,N_32342,N_32389);
xnor U32620 (N_32620,N_32161,N_32184);
xor U32621 (N_32621,N_32408,N_32318);
nor U32622 (N_32622,N_32331,N_32162);
nand U32623 (N_32623,N_32498,N_32246);
or U32624 (N_32624,N_32402,N_32164);
nand U32625 (N_32625,N_32175,N_32404);
xnor U32626 (N_32626,N_32313,N_32365);
nand U32627 (N_32627,N_32039,N_32321);
nor U32628 (N_32628,N_32422,N_32051);
or U32629 (N_32629,N_32153,N_32054);
or U32630 (N_32630,N_32221,N_32409);
or U32631 (N_32631,N_32305,N_32442);
nor U32632 (N_32632,N_32207,N_32122);
nand U32633 (N_32633,N_32189,N_32459);
nor U32634 (N_32634,N_32324,N_32193);
nor U32635 (N_32635,N_32484,N_32394);
nor U32636 (N_32636,N_32038,N_32483);
and U32637 (N_32637,N_32292,N_32330);
xor U32638 (N_32638,N_32106,N_32204);
or U32639 (N_32639,N_32022,N_32495);
xnor U32640 (N_32640,N_32197,N_32272);
nand U32641 (N_32641,N_32066,N_32295);
nor U32642 (N_32642,N_32141,N_32470);
nor U32643 (N_32643,N_32385,N_32253);
and U32644 (N_32644,N_32147,N_32291);
nor U32645 (N_32645,N_32103,N_32142);
nand U32646 (N_32646,N_32060,N_32160);
or U32647 (N_32647,N_32298,N_32405);
and U32648 (N_32648,N_32303,N_32014);
or U32649 (N_32649,N_32296,N_32335);
xnor U32650 (N_32650,N_32148,N_32490);
or U32651 (N_32651,N_32383,N_32461);
xnor U32652 (N_32652,N_32341,N_32285);
nand U32653 (N_32653,N_32042,N_32407);
nor U32654 (N_32654,N_32132,N_32059);
xor U32655 (N_32655,N_32450,N_32395);
and U32656 (N_32656,N_32124,N_32366);
nand U32657 (N_32657,N_32258,N_32454);
nand U32658 (N_32658,N_32414,N_32280);
nor U32659 (N_32659,N_32277,N_32087);
or U32660 (N_32660,N_32281,N_32023);
nand U32661 (N_32661,N_32158,N_32419);
and U32662 (N_32662,N_32000,N_32457);
nand U32663 (N_32663,N_32061,N_32282);
xor U32664 (N_32664,N_32196,N_32199);
xnor U32665 (N_32665,N_32327,N_32261);
xnor U32666 (N_32666,N_32003,N_32192);
nor U32667 (N_32667,N_32309,N_32381);
nand U32668 (N_32668,N_32447,N_32086);
xnor U32669 (N_32669,N_32088,N_32018);
nand U32670 (N_32670,N_32424,N_32084);
and U32671 (N_32671,N_32058,N_32217);
nor U32672 (N_32672,N_32064,N_32393);
and U32673 (N_32673,N_32069,N_32044);
nor U32674 (N_32674,N_32101,N_32052);
and U32675 (N_32675,N_32260,N_32113);
or U32676 (N_32676,N_32004,N_32255);
and U32677 (N_32677,N_32170,N_32202);
nand U32678 (N_32678,N_32176,N_32432);
nand U32679 (N_32679,N_32333,N_32095);
nand U32680 (N_32680,N_32015,N_32188);
or U32681 (N_32681,N_32187,N_32427);
xnor U32682 (N_32682,N_32248,N_32182);
and U32683 (N_32683,N_32279,N_32464);
and U32684 (N_32684,N_32401,N_32127);
nor U32685 (N_32685,N_32191,N_32200);
xnor U32686 (N_32686,N_32030,N_32367);
nand U32687 (N_32687,N_32046,N_32040);
and U32688 (N_32688,N_32231,N_32315);
nor U32689 (N_32689,N_32008,N_32284);
nor U32690 (N_32690,N_32032,N_32135);
nand U32691 (N_32691,N_32446,N_32254);
nand U32692 (N_32692,N_32382,N_32399);
xnor U32693 (N_32693,N_32397,N_32063);
xnor U32694 (N_32694,N_32326,N_32201);
nor U32695 (N_32695,N_32379,N_32340);
nor U32696 (N_32696,N_32016,N_32082);
nor U32697 (N_32697,N_32236,N_32494);
or U32698 (N_32698,N_32163,N_32437);
or U32699 (N_32699,N_32434,N_32043);
and U32700 (N_32700,N_32238,N_32312);
nand U32701 (N_32701,N_32265,N_32301);
and U32702 (N_32702,N_32245,N_32435);
xor U32703 (N_32703,N_32227,N_32334);
xor U32704 (N_32704,N_32425,N_32467);
nor U32705 (N_32705,N_32499,N_32348);
nand U32706 (N_32706,N_32190,N_32120);
xor U32707 (N_32707,N_32102,N_32119);
nor U32708 (N_32708,N_32288,N_32368);
and U32709 (N_32709,N_32180,N_32041);
nor U32710 (N_32710,N_32156,N_32297);
xor U32711 (N_32711,N_32114,N_32011);
nor U32712 (N_32712,N_32449,N_32235);
or U32713 (N_32713,N_32489,N_32466);
and U32714 (N_32714,N_32283,N_32090);
and U32715 (N_32715,N_32257,N_32264);
nand U32716 (N_32716,N_32276,N_32474);
nor U32717 (N_32717,N_32387,N_32441);
and U32718 (N_32718,N_32009,N_32150);
and U32719 (N_32719,N_32354,N_32493);
nor U32720 (N_32720,N_32423,N_32429);
nand U32721 (N_32721,N_32118,N_32024);
nor U32722 (N_32722,N_32083,N_32112);
and U32723 (N_32723,N_32036,N_32092);
nand U32724 (N_32724,N_32075,N_32413);
and U32725 (N_32725,N_32380,N_32130);
and U32726 (N_32726,N_32273,N_32431);
nor U32727 (N_32727,N_32421,N_32035);
nand U32728 (N_32728,N_32017,N_32476);
or U32729 (N_32729,N_32117,N_32098);
xor U32730 (N_32730,N_32099,N_32440);
xor U32731 (N_32731,N_32050,N_32218);
or U32732 (N_32732,N_32073,N_32171);
nand U32733 (N_32733,N_32398,N_32049);
and U32734 (N_32734,N_32250,N_32377);
and U32735 (N_32735,N_32332,N_32047);
xor U32736 (N_32736,N_32293,N_32453);
nand U32737 (N_32737,N_32019,N_32020);
nand U32738 (N_32738,N_32198,N_32183);
and U32739 (N_32739,N_32317,N_32468);
nand U32740 (N_32740,N_32438,N_32290);
or U32741 (N_32741,N_32242,N_32482);
and U32742 (N_32742,N_32131,N_32458);
xnor U32743 (N_32743,N_32452,N_32157);
nor U32744 (N_32744,N_32195,N_32355);
nor U32745 (N_32745,N_32220,N_32487);
nand U32746 (N_32746,N_32048,N_32416);
nand U32747 (N_32747,N_32239,N_32169);
nand U32748 (N_32748,N_32026,N_32415);
or U32749 (N_32749,N_32275,N_32363);
xor U32750 (N_32750,N_32212,N_32095);
xnor U32751 (N_32751,N_32348,N_32209);
nor U32752 (N_32752,N_32406,N_32212);
nand U32753 (N_32753,N_32272,N_32274);
and U32754 (N_32754,N_32020,N_32426);
nor U32755 (N_32755,N_32182,N_32429);
or U32756 (N_32756,N_32409,N_32111);
nor U32757 (N_32757,N_32386,N_32254);
or U32758 (N_32758,N_32034,N_32077);
nor U32759 (N_32759,N_32077,N_32241);
and U32760 (N_32760,N_32201,N_32086);
or U32761 (N_32761,N_32307,N_32468);
and U32762 (N_32762,N_32270,N_32487);
xnor U32763 (N_32763,N_32251,N_32108);
nor U32764 (N_32764,N_32493,N_32344);
or U32765 (N_32765,N_32280,N_32411);
xnor U32766 (N_32766,N_32169,N_32317);
xor U32767 (N_32767,N_32433,N_32331);
and U32768 (N_32768,N_32086,N_32175);
nor U32769 (N_32769,N_32295,N_32396);
and U32770 (N_32770,N_32106,N_32079);
or U32771 (N_32771,N_32094,N_32237);
xor U32772 (N_32772,N_32365,N_32355);
nand U32773 (N_32773,N_32231,N_32110);
xnor U32774 (N_32774,N_32038,N_32439);
xor U32775 (N_32775,N_32325,N_32364);
xor U32776 (N_32776,N_32327,N_32360);
nor U32777 (N_32777,N_32458,N_32332);
and U32778 (N_32778,N_32313,N_32268);
nor U32779 (N_32779,N_32432,N_32471);
nand U32780 (N_32780,N_32080,N_32097);
or U32781 (N_32781,N_32421,N_32288);
and U32782 (N_32782,N_32349,N_32225);
xor U32783 (N_32783,N_32262,N_32196);
nand U32784 (N_32784,N_32176,N_32243);
xnor U32785 (N_32785,N_32308,N_32288);
and U32786 (N_32786,N_32133,N_32493);
xor U32787 (N_32787,N_32173,N_32150);
and U32788 (N_32788,N_32282,N_32491);
nand U32789 (N_32789,N_32202,N_32281);
nor U32790 (N_32790,N_32181,N_32045);
nand U32791 (N_32791,N_32434,N_32000);
xor U32792 (N_32792,N_32004,N_32362);
or U32793 (N_32793,N_32365,N_32155);
or U32794 (N_32794,N_32263,N_32270);
nor U32795 (N_32795,N_32297,N_32117);
and U32796 (N_32796,N_32363,N_32278);
and U32797 (N_32797,N_32345,N_32120);
or U32798 (N_32798,N_32002,N_32069);
xor U32799 (N_32799,N_32476,N_32307);
or U32800 (N_32800,N_32439,N_32420);
or U32801 (N_32801,N_32196,N_32393);
and U32802 (N_32802,N_32230,N_32124);
xor U32803 (N_32803,N_32114,N_32194);
and U32804 (N_32804,N_32107,N_32400);
nor U32805 (N_32805,N_32437,N_32027);
xnor U32806 (N_32806,N_32054,N_32247);
or U32807 (N_32807,N_32018,N_32201);
nor U32808 (N_32808,N_32100,N_32175);
xor U32809 (N_32809,N_32208,N_32246);
nor U32810 (N_32810,N_32100,N_32042);
xnor U32811 (N_32811,N_32441,N_32186);
and U32812 (N_32812,N_32152,N_32099);
and U32813 (N_32813,N_32265,N_32388);
xor U32814 (N_32814,N_32115,N_32140);
and U32815 (N_32815,N_32025,N_32224);
xnor U32816 (N_32816,N_32442,N_32402);
xnor U32817 (N_32817,N_32001,N_32214);
nor U32818 (N_32818,N_32154,N_32204);
nand U32819 (N_32819,N_32137,N_32408);
xor U32820 (N_32820,N_32251,N_32044);
or U32821 (N_32821,N_32491,N_32072);
and U32822 (N_32822,N_32487,N_32138);
xor U32823 (N_32823,N_32134,N_32182);
and U32824 (N_32824,N_32214,N_32345);
nor U32825 (N_32825,N_32326,N_32001);
or U32826 (N_32826,N_32271,N_32036);
xor U32827 (N_32827,N_32235,N_32423);
xnor U32828 (N_32828,N_32293,N_32284);
nand U32829 (N_32829,N_32091,N_32082);
nand U32830 (N_32830,N_32339,N_32407);
and U32831 (N_32831,N_32153,N_32477);
nand U32832 (N_32832,N_32196,N_32135);
xor U32833 (N_32833,N_32246,N_32347);
or U32834 (N_32834,N_32453,N_32189);
nand U32835 (N_32835,N_32122,N_32447);
xnor U32836 (N_32836,N_32120,N_32140);
nand U32837 (N_32837,N_32103,N_32081);
nor U32838 (N_32838,N_32307,N_32482);
nor U32839 (N_32839,N_32236,N_32206);
or U32840 (N_32840,N_32260,N_32100);
xor U32841 (N_32841,N_32233,N_32316);
xnor U32842 (N_32842,N_32191,N_32197);
nand U32843 (N_32843,N_32307,N_32236);
and U32844 (N_32844,N_32454,N_32449);
nor U32845 (N_32845,N_32229,N_32276);
nor U32846 (N_32846,N_32221,N_32052);
xnor U32847 (N_32847,N_32260,N_32005);
or U32848 (N_32848,N_32017,N_32068);
nand U32849 (N_32849,N_32224,N_32003);
and U32850 (N_32850,N_32358,N_32016);
xnor U32851 (N_32851,N_32158,N_32013);
xor U32852 (N_32852,N_32374,N_32159);
xnor U32853 (N_32853,N_32452,N_32306);
and U32854 (N_32854,N_32146,N_32400);
nor U32855 (N_32855,N_32009,N_32121);
xnor U32856 (N_32856,N_32372,N_32297);
xor U32857 (N_32857,N_32027,N_32116);
nand U32858 (N_32858,N_32175,N_32177);
xor U32859 (N_32859,N_32223,N_32265);
nor U32860 (N_32860,N_32282,N_32404);
xor U32861 (N_32861,N_32414,N_32229);
nor U32862 (N_32862,N_32305,N_32070);
nand U32863 (N_32863,N_32383,N_32200);
nor U32864 (N_32864,N_32467,N_32166);
and U32865 (N_32865,N_32427,N_32182);
nor U32866 (N_32866,N_32366,N_32051);
nor U32867 (N_32867,N_32067,N_32025);
or U32868 (N_32868,N_32190,N_32024);
and U32869 (N_32869,N_32437,N_32356);
and U32870 (N_32870,N_32056,N_32098);
and U32871 (N_32871,N_32000,N_32375);
xnor U32872 (N_32872,N_32473,N_32194);
nand U32873 (N_32873,N_32161,N_32175);
nand U32874 (N_32874,N_32436,N_32427);
nor U32875 (N_32875,N_32373,N_32315);
or U32876 (N_32876,N_32245,N_32432);
or U32877 (N_32877,N_32137,N_32332);
nand U32878 (N_32878,N_32096,N_32035);
or U32879 (N_32879,N_32469,N_32406);
nor U32880 (N_32880,N_32483,N_32441);
and U32881 (N_32881,N_32249,N_32093);
xnor U32882 (N_32882,N_32125,N_32123);
nor U32883 (N_32883,N_32001,N_32155);
nor U32884 (N_32884,N_32046,N_32402);
nor U32885 (N_32885,N_32341,N_32491);
nand U32886 (N_32886,N_32489,N_32458);
xnor U32887 (N_32887,N_32440,N_32454);
or U32888 (N_32888,N_32351,N_32244);
nand U32889 (N_32889,N_32217,N_32498);
nor U32890 (N_32890,N_32338,N_32038);
and U32891 (N_32891,N_32462,N_32418);
xnor U32892 (N_32892,N_32010,N_32302);
and U32893 (N_32893,N_32177,N_32188);
xnor U32894 (N_32894,N_32321,N_32460);
nand U32895 (N_32895,N_32488,N_32083);
or U32896 (N_32896,N_32123,N_32461);
xor U32897 (N_32897,N_32228,N_32321);
and U32898 (N_32898,N_32347,N_32213);
xnor U32899 (N_32899,N_32460,N_32342);
and U32900 (N_32900,N_32107,N_32040);
and U32901 (N_32901,N_32181,N_32473);
nor U32902 (N_32902,N_32097,N_32488);
or U32903 (N_32903,N_32206,N_32127);
or U32904 (N_32904,N_32332,N_32190);
xor U32905 (N_32905,N_32170,N_32234);
nand U32906 (N_32906,N_32348,N_32188);
or U32907 (N_32907,N_32152,N_32400);
nand U32908 (N_32908,N_32147,N_32167);
nor U32909 (N_32909,N_32235,N_32043);
or U32910 (N_32910,N_32251,N_32320);
and U32911 (N_32911,N_32154,N_32285);
xnor U32912 (N_32912,N_32034,N_32489);
and U32913 (N_32913,N_32320,N_32285);
nor U32914 (N_32914,N_32060,N_32157);
nand U32915 (N_32915,N_32325,N_32051);
nand U32916 (N_32916,N_32457,N_32462);
or U32917 (N_32917,N_32261,N_32316);
nor U32918 (N_32918,N_32243,N_32385);
or U32919 (N_32919,N_32465,N_32237);
nand U32920 (N_32920,N_32041,N_32123);
xnor U32921 (N_32921,N_32069,N_32032);
or U32922 (N_32922,N_32441,N_32237);
nor U32923 (N_32923,N_32298,N_32157);
xor U32924 (N_32924,N_32303,N_32293);
xor U32925 (N_32925,N_32014,N_32163);
or U32926 (N_32926,N_32236,N_32303);
and U32927 (N_32927,N_32213,N_32040);
xor U32928 (N_32928,N_32473,N_32224);
nor U32929 (N_32929,N_32336,N_32427);
or U32930 (N_32930,N_32291,N_32461);
nand U32931 (N_32931,N_32415,N_32471);
nor U32932 (N_32932,N_32408,N_32391);
nand U32933 (N_32933,N_32083,N_32024);
nor U32934 (N_32934,N_32199,N_32435);
and U32935 (N_32935,N_32392,N_32391);
nor U32936 (N_32936,N_32138,N_32002);
or U32937 (N_32937,N_32270,N_32033);
xor U32938 (N_32938,N_32135,N_32112);
xnor U32939 (N_32939,N_32205,N_32090);
or U32940 (N_32940,N_32357,N_32434);
xor U32941 (N_32941,N_32070,N_32093);
xor U32942 (N_32942,N_32001,N_32019);
nand U32943 (N_32943,N_32119,N_32065);
nor U32944 (N_32944,N_32399,N_32200);
xor U32945 (N_32945,N_32291,N_32132);
or U32946 (N_32946,N_32194,N_32370);
xnor U32947 (N_32947,N_32033,N_32182);
and U32948 (N_32948,N_32393,N_32136);
and U32949 (N_32949,N_32105,N_32067);
nand U32950 (N_32950,N_32457,N_32256);
or U32951 (N_32951,N_32218,N_32390);
and U32952 (N_32952,N_32143,N_32334);
xor U32953 (N_32953,N_32026,N_32003);
or U32954 (N_32954,N_32232,N_32100);
and U32955 (N_32955,N_32385,N_32103);
and U32956 (N_32956,N_32374,N_32455);
xor U32957 (N_32957,N_32205,N_32270);
xnor U32958 (N_32958,N_32498,N_32499);
xor U32959 (N_32959,N_32078,N_32119);
nor U32960 (N_32960,N_32118,N_32496);
nor U32961 (N_32961,N_32406,N_32113);
nor U32962 (N_32962,N_32361,N_32007);
and U32963 (N_32963,N_32074,N_32225);
and U32964 (N_32964,N_32427,N_32282);
nor U32965 (N_32965,N_32154,N_32256);
and U32966 (N_32966,N_32109,N_32419);
nor U32967 (N_32967,N_32478,N_32231);
and U32968 (N_32968,N_32325,N_32392);
xor U32969 (N_32969,N_32401,N_32214);
and U32970 (N_32970,N_32217,N_32473);
nand U32971 (N_32971,N_32087,N_32048);
and U32972 (N_32972,N_32449,N_32437);
nor U32973 (N_32973,N_32471,N_32468);
nand U32974 (N_32974,N_32302,N_32126);
nor U32975 (N_32975,N_32236,N_32258);
nand U32976 (N_32976,N_32198,N_32216);
xor U32977 (N_32977,N_32156,N_32382);
xnor U32978 (N_32978,N_32190,N_32425);
nand U32979 (N_32979,N_32347,N_32221);
xor U32980 (N_32980,N_32496,N_32391);
nand U32981 (N_32981,N_32358,N_32461);
nand U32982 (N_32982,N_32040,N_32456);
xor U32983 (N_32983,N_32498,N_32473);
xor U32984 (N_32984,N_32037,N_32313);
nor U32985 (N_32985,N_32070,N_32454);
and U32986 (N_32986,N_32282,N_32246);
nor U32987 (N_32987,N_32395,N_32300);
nand U32988 (N_32988,N_32125,N_32171);
and U32989 (N_32989,N_32266,N_32293);
nand U32990 (N_32990,N_32471,N_32357);
nand U32991 (N_32991,N_32202,N_32235);
nand U32992 (N_32992,N_32415,N_32115);
and U32993 (N_32993,N_32138,N_32193);
xnor U32994 (N_32994,N_32166,N_32044);
or U32995 (N_32995,N_32251,N_32400);
nor U32996 (N_32996,N_32014,N_32074);
xnor U32997 (N_32997,N_32165,N_32392);
nand U32998 (N_32998,N_32301,N_32444);
nand U32999 (N_32999,N_32317,N_32388);
xor U33000 (N_33000,N_32768,N_32789);
and U33001 (N_33001,N_32791,N_32525);
or U33002 (N_33002,N_32905,N_32573);
and U33003 (N_33003,N_32839,N_32888);
nand U33004 (N_33004,N_32620,N_32769);
nand U33005 (N_33005,N_32536,N_32503);
nor U33006 (N_33006,N_32514,N_32603);
or U33007 (N_33007,N_32925,N_32749);
and U33008 (N_33008,N_32940,N_32647);
or U33009 (N_33009,N_32733,N_32863);
or U33010 (N_33010,N_32630,N_32838);
and U33011 (N_33011,N_32668,N_32785);
nor U33012 (N_33012,N_32725,N_32656);
nor U33013 (N_33013,N_32866,N_32677);
xor U33014 (N_33014,N_32640,N_32822);
nand U33015 (N_33015,N_32897,N_32505);
xor U33016 (N_33016,N_32534,N_32676);
xor U33017 (N_33017,N_32535,N_32641);
xor U33018 (N_33018,N_32973,N_32986);
xnor U33019 (N_33019,N_32841,N_32758);
xor U33020 (N_33020,N_32735,N_32646);
or U33021 (N_33021,N_32670,N_32949);
xor U33022 (N_33022,N_32806,N_32605);
and U33023 (N_33023,N_32844,N_32974);
and U33024 (N_33024,N_32527,N_32858);
nor U33025 (N_33025,N_32734,N_32522);
nand U33026 (N_33026,N_32941,N_32853);
nand U33027 (N_33027,N_32955,N_32933);
nor U33028 (N_33028,N_32642,N_32880);
and U33029 (N_33029,N_32786,N_32626);
or U33030 (N_33030,N_32851,N_32645);
nor U33031 (N_33031,N_32512,N_32988);
or U33032 (N_33032,N_32910,N_32728);
or U33033 (N_33033,N_32837,N_32588);
or U33034 (N_33034,N_32765,N_32520);
xor U33035 (N_33035,N_32766,N_32629);
nand U33036 (N_33036,N_32756,N_32750);
xor U33037 (N_33037,N_32873,N_32554);
and U33038 (N_33038,N_32990,N_32589);
nand U33039 (N_33039,N_32587,N_32875);
or U33040 (N_33040,N_32767,N_32681);
or U33041 (N_33041,N_32693,N_32740);
nand U33042 (N_33042,N_32931,N_32657);
nand U33043 (N_33043,N_32964,N_32994);
xnor U33044 (N_33044,N_32682,N_32528);
xnor U33045 (N_33045,N_32703,N_32590);
nand U33046 (N_33046,N_32654,N_32576);
xnor U33047 (N_33047,N_32529,N_32661);
and U33048 (N_33048,N_32914,N_32803);
nor U33049 (N_33049,N_32978,N_32778);
nand U33050 (N_33050,N_32755,N_32730);
nand U33051 (N_33051,N_32606,N_32736);
and U33052 (N_33052,N_32784,N_32928);
nand U33053 (N_33053,N_32510,N_32989);
nor U33054 (N_33054,N_32917,N_32753);
xor U33055 (N_33055,N_32698,N_32560);
or U33056 (N_33056,N_32744,N_32660);
and U33057 (N_33057,N_32859,N_32961);
or U33058 (N_33058,N_32846,N_32594);
and U33059 (N_33059,N_32591,N_32686);
xnor U33060 (N_33060,N_32948,N_32570);
and U33061 (N_33061,N_32991,N_32622);
nand U33062 (N_33062,N_32516,N_32965);
xnor U33063 (N_33063,N_32501,N_32831);
nand U33064 (N_33064,N_32855,N_32679);
or U33065 (N_33065,N_32892,N_32739);
or U33066 (N_33066,N_32705,N_32809);
xor U33067 (N_33067,N_32638,N_32530);
and U33068 (N_33068,N_32615,N_32883);
nor U33069 (N_33069,N_32884,N_32559);
or U33070 (N_33070,N_32712,N_32509);
and U33071 (N_33071,N_32592,N_32548);
nand U33072 (N_33072,N_32816,N_32850);
xnor U33073 (N_33073,N_32960,N_32600);
xor U33074 (N_33074,N_32671,N_32760);
nand U33075 (N_33075,N_32796,N_32781);
and U33076 (N_33076,N_32823,N_32927);
or U33077 (N_33077,N_32867,N_32821);
nand U33078 (N_33078,N_32618,N_32631);
or U33079 (N_33079,N_32721,N_32602);
nand U33080 (N_33080,N_32956,N_32757);
or U33081 (N_33081,N_32706,N_32819);
nor U33082 (N_33082,N_32727,N_32979);
nand U33083 (N_33083,N_32957,N_32623);
xnor U33084 (N_33084,N_32718,N_32687);
and U33085 (N_33085,N_32524,N_32691);
or U33086 (N_33086,N_32665,N_32737);
nand U33087 (N_33087,N_32860,N_32754);
nand U33088 (N_33088,N_32871,N_32540);
xnor U33089 (N_33089,N_32586,N_32865);
nand U33090 (N_33090,N_32616,N_32729);
nand U33091 (N_33091,N_32827,N_32982);
nand U33092 (N_33092,N_32663,N_32811);
nor U33093 (N_33093,N_32523,N_32843);
and U33094 (N_33094,N_32929,N_32558);
or U33095 (N_33095,N_32993,N_32842);
nor U33096 (N_33096,N_32526,N_32511);
xnor U33097 (N_33097,N_32607,N_32696);
xor U33098 (N_33098,N_32984,N_32814);
and U33099 (N_33099,N_32908,N_32857);
xor U33100 (N_33100,N_32713,N_32909);
or U33101 (N_33101,N_32655,N_32751);
xnor U33102 (N_33102,N_32748,N_32566);
nand U33103 (N_33103,N_32920,N_32787);
nor U33104 (N_33104,N_32674,N_32967);
nand U33105 (N_33105,N_32584,N_32653);
and U33106 (N_33106,N_32862,N_32543);
or U33107 (N_33107,N_32808,N_32724);
and U33108 (N_33108,N_32697,N_32699);
and U33109 (N_33109,N_32627,N_32969);
nand U33110 (N_33110,N_32612,N_32864);
nor U33111 (N_33111,N_32707,N_32692);
nand U33112 (N_33112,N_32572,N_32950);
xor U33113 (N_33113,N_32804,N_32644);
or U33114 (N_33114,N_32911,N_32714);
nand U33115 (N_33115,N_32711,N_32595);
or U33116 (N_33116,N_32719,N_32889);
nand U33117 (N_33117,N_32829,N_32688);
and U33118 (N_33118,N_32885,N_32856);
nand U33119 (N_33119,N_32980,N_32907);
or U33120 (N_33120,N_32801,N_32893);
and U33121 (N_33121,N_32683,N_32938);
or U33122 (N_33122,N_32992,N_32828);
nor U33123 (N_33123,N_32678,N_32902);
and U33124 (N_33124,N_32848,N_32834);
or U33125 (N_33125,N_32762,N_32886);
xor U33126 (N_33126,N_32771,N_32502);
nand U33127 (N_33127,N_32847,N_32568);
and U33128 (N_33128,N_32652,N_32635);
nor U33129 (N_33129,N_32557,N_32545);
nand U33130 (N_33130,N_32575,N_32983);
nor U33131 (N_33131,N_32799,N_32539);
and U33132 (N_33132,N_32824,N_32672);
nor U33133 (N_33133,N_32924,N_32872);
and U33134 (N_33134,N_32611,N_32985);
nand U33135 (N_33135,N_32722,N_32604);
and U33136 (N_33136,N_32977,N_32966);
or U33137 (N_33137,N_32997,N_32664);
nor U33138 (N_33138,N_32541,N_32946);
and U33139 (N_33139,N_32794,N_32521);
and U33140 (N_33140,N_32962,N_32564);
nand U33141 (N_33141,N_32628,N_32579);
xnor U33142 (N_33142,N_32710,N_32731);
and U33143 (N_33143,N_32770,N_32639);
nand U33144 (N_33144,N_32807,N_32658);
or U33145 (N_33145,N_32613,N_32648);
and U33146 (N_33146,N_32608,N_32596);
nor U33147 (N_33147,N_32832,N_32849);
xor U33148 (N_33148,N_32976,N_32783);
nand U33149 (N_33149,N_32836,N_32773);
or U33150 (N_33150,N_32567,N_32798);
xnor U33151 (N_33151,N_32553,N_32634);
or U33152 (N_33152,N_32578,N_32542);
and U33153 (N_33153,N_32732,N_32702);
xnor U33154 (N_33154,N_32632,N_32593);
or U33155 (N_33155,N_32825,N_32515);
xnor U33156 (N_33156,N_32562,N_32550);
and U33157 (N_33157,N_32854,N_32812);
nand U33158 (N_33158,N_32574,N_32695);
xor U33159 (N_33159,N_32936,N_32921);
nand U33160 (N_33160,N_32890,N_32903);
xnor U33161 (N_33161,N_32970,N_32617);
nor U33162 (N_33162,N_32585,N_32926);
nand U33163 (N_33163,N_32565,N_32820);
and U33164 (N_33164,N_32896,N_32598);
nor U33165 (N_33165,N_32552,N_32555);
nand U33166 (N_33166,N_32556,N_32915);
or U33167 (N_33167,N_32882,N_32998);
or U33168 (N_33168,N_32899,N_32852);
or U33169 (N_33169,N_32944,N_32715);
or U33170 (N_33170,N_32700,N_32636);
and U33171 (N_33171,N_32869,N_32800);
nand U33172 (N_33172,N_32795,N_32504);
nor U33173 (N_33173,N_32930,N_32959);
nor U33174 (N_33174,N_32895,N_32942);
and U33175 (N_33175,N_32995,N_32935);
xnor U33176 (N_33176,N_32513,N_32934);
or U33177 (N_33177,N_32675,N_32782);
nor U33178 (N_33178,N_32532,N_32651);
nand U33179 (N_33179,N_32500,N_32738);
and U33180 (N_33180,N_32887,N_32996);
nand U33181 (N_33181,N_32601,N_32761);
xor U33182 (N_33182,N_32818,N_32861);
or U33183 (N_33183,N_32610,N_32519);
or U33184 (N_33184,N_32544,N_32830);
or U33185 (N_33185,N_32810,N_32793);
and U33186 (N_33186,N_32547,N_32746);
and U33187 (N_33187,N_32833,N_32900);
nor U33188 (N_33188,N_32981,N_32633);
nand U33189 (N_33189,N_32840,N_32792);
and U33190 (N_33190,N_32788,N_32741);
and U33191 (N_33191,N_32747,N_32764);
or U33192 (N_33192,N_32694,N_32987);
or U33193 (N_33193,N_32943,N_32802);
and U33194 (N_33194,N_32922,N_32621);
xor U33195 (N_33195,N_32720,N_32813);
nand U33196 (N_33196,N_32582,N_32906);
nor U33197 (N_33197,N_32625,N_32951);
or U33198 (N_33198,N_32901,N_32637);
nor U33199 (N_33199,N_32680,N_32538);
xor U33200 (N_33200,N_32561,N_32999);
or U33201 (N_33201,N_32937,N_32916);
nand U33202 (N_33202,N_32904,N_32614);
nor U33203 (N_33203,N_32772,N_32546);
and U33204 (N_33204,N_32790,N_32963);
nor U33205 (N_33205,N_32918,N_32742);
nand U33206 (N_33206,N_32780,N_32533);
xnor U33207 (N_33207,N_32569,N_32577);
and U33208 (N_33208,N_32506,N_32701);
or U33209 (N_33209,N_32953,N_32975);
and U33210 (N_33210,N_32537,N_32779);
nand U33211 (N_33211,N_32716,N_32923);
nor U33212 (N_33212,N_32549,N_32583);
or U33213 (N_33213,N_32717,N_32891);
xor U33214 (N_33214,N_32726,N_32815);
and U33215 (N_33215,N_32759,N_32684);
or U33216 (N_33216,N_32894,N_32878);
xor U33217 (N_33217,N_32835,N_32580);
xor U33218 (N_33218,N_32939,N_32919);
or U33219 (N_33219,N_32752,N_32667);
nand U33220 (N_33220,N_32673,N_32805);
nor U33221 (N_33221,N_32704,N_32507);
nor U33222 (N_33222,N_32968,N_32581);
and U33223 (N_33223,N_32972,N_32649);
nand U33224 (N_33224,N_32709,N_32826);
or U33225 (N_33225,N_32912,N_32817);
and U33226 (N_33226,N_32874,N_32690);
nor U33227 (N_33227,N_32774,N_32597);
nor U33228 (N_33228,N_32551,N_32881);
and U33229 (N_33229,N_32877,N_32954);
nand U33230 (N_33230,N_32743,N_32650);
or U33231 (N_33231,N_32763,N_32518);
or U33232 (N_33232,N_32845,N_32666);
xnor U33233 (N_33233,N_32870,N_32508);
nand U33234 (N_33234,N_32971,N_32952);
nand U33235 (N_33235,N_32745,N_32723);
and U33236 (N_33236,N_32876,N_32947);
and U33237 (N_33237,N_32689,N_32913);
or U33238 (N_33238,N_32517,N_32563);
and U33239 (N_33239,N_32599,N_32643);
nor U33240 (N_33240,N_32945,N_32932);
xnor U33241 (N_33241,N_32797,N_32868);
and U33242 (N_33242,N_32685,N_32662);
nor U33243 (N_33243,N_32708,N_32531);
nand U33244 (N_33244,N_32958,N_32609);
or U33245 (N_33245,N_32777,N_32669);
xnor U33246 (N_33246,N_32879,N_32659);
xnor U33247 (N_33247,N_32775,N_32624);
nand U33248 (N_33248,N_32776,N_32571);
xor U33249 (N_33249,N_32619,N_32898);
or U33250 (N_33250,N_32915,N_32672);
nand U33251 (N_33251,N_32792,N_32559);
or U33252 (N_33252,N_32759,N_32566);
or U33253 (N_33253,N_32923,N_32611);
xor U33254 (N_33254,N_32909,N_32785);
nand U33255 (N_33255,N_32651,N_32881);
xor U33256 (N_33256,N_32546,N_32536);
xor U33257 (N_33257,N_32864,N_32921);
nand U33258 (N_33258,N_32625,N_32838);
xnor U33259 (N_33259,N_32835,N_32851);
nor U33260 (N_33260,N_32624,N_32618);
nand U33261 (N_33261,N_32843,N_32741);
nand U33262 (N_33262,N_32674,N_32953);
xnor U33263 (N_33263,N_32818,N_32722);
xor U33264 (N_33264,N_32656,N_32869);
nand U33265 (N_33265,N_32665,N_32899);
xnor U33266 (N_33266,N_32653,N_32919);
xnor U33267 (N_33267,N_32564,N_32511);
nor U33268 (N_33268,N_32832,N_32536);
and U33269 (N_33269,N_32669,N_32774);
and U33270 (N_33270,N_32801,N_32683);
nand U33271 (N_33271,N_32930,N_32911);
or U33272 (N_33272,N_32764,N_32791);
xor U33273 (N_33273,N_32823,N_32577);
and U33274 (N_33274,N_32571,N_32560);
nand U33275 (N_33275,N_32862,N_32789);
and U33276 (N_33276,N_32865,N_32678);
nand U33277 (N_33277,N_32840,N_32850);
nor U33278 (N_33278,N_32749,N_32563);
xnor U33279 (N_33279,N_32589,N_32936);
or U33280 (N_33280,N_32652,N_32583);
or U33281 (N_33281,N_32591,N_32876);
or U33282 (N_33282,N_32530,N_32549);
or U33283 (N_33283,N_32724,N_32929);
and U33284 (N_33284,N_32704,N_32703);
and U33285 (N_33285,N_32535,N_32649);
and U33286 (N_33286,N_32925,N_32683);
nand U33287 (N_33287,N_32544,N_32547);
xor U33288 (N_33288,N_32521,N_32745);
xnor U33289 (N_33289,N_32881,N_32610);
or U33290 (N_33290,N_32718,N_32770);
nor U33291 (N_33291,N_32574,N_32597);
or U33292 (N_33292,N_32850,N_32670);
or U33293 (N_33293,N_32550,N_32532);
and U33294 (N_33294,N_32666,N_32797);
and U33295 (N_33295,N_32566,N_32928);
nor U33296 (N_33296,N_32884,N_32808);
xnor U33297 (N_33297,N_32971,N_32745);
nand U33298 (N_33298,N_32674,N_32808);
and U33299 (N_33299,N_32714,N_32881);
nand U33300 (N_33300,N_32884,N_32502);
and U33301 (N_33301,N_32883,N_32610);
nor U33302 (N_33302,N_32856,N_32881);
and U33303 (N_33303,N_32762,N_32985);
or U33304 (N_33304,N_32935,N_32733);
nand U33305 (N_33305,N_32633,N_32653);
or U33306 (N_33306,N_32907,N_32669);
and U33307 (N_33307,N_32697,N_32505);
nor U33308 (N_33308,N_32712,N_32861);
xnor U33309 (N_33309,N_32953,N_32834);
nand U33310 (N_33310,N_32929,N_32541);
xnor U33311 (N_33311,N_32710,N_32667);
nor U33312 (N_33312,N_32938,N_32652);
nor U33313 (N_33313,N_32595,N_32527);
nor U33314 (N_33314,N_32906,N_32634);
xnor U33315 (N_33315,N_32706,N_32544);
nor U33316 (N_33316,N_32545,N_32806);
nor U33317 (N_33317,N_32622,N_32718);
nor U33318 (N_33318,N_32782,N_32707);
and U33319 (N_33319,N_32564,N_32964);
xor U33320 (N_33320,N_32835,N_32895);
or U33321 (N_33321,N_32801,N_32676);
nor U33322 (N_33322,N_32986,N_32795);
and U33323 (N_33323,N_32740,N_32699);
nand U33324 (N_33324,N_32795,N_32990);
nor U33325 (N_33325,N_32844,N_32675);
and U33326 (N_33326,N_32514,N_32986);
nand U33327 (N_33327,N_32998,N_32846);
xor U33328 (N_33328,N_32649,N_32898);
and U33329 (N_33329,N_32825,N_32672);
nor U33330 (N_33330,N_32541,N_32745);
and U33331 (N_33331,N_32836,N_32720);
and U33332 (N_33332,N_32547,N_32736);
nor U33333 (N_33333,N_32918,N_32636);
nor U33334 (N_33334,N_32901,N_32930);
or U33335 (N_33335,N_32942,N_32731);
nand U33336 (N_33336,N_32737,N_32958);
nor U33337 (N_33337,N_32758,N_32543);
xor U33338 (N_33338,N_32961,N_32607);
nand U33339 (N_33339,N_32542,N_32931);
or U33340 (N_33340,N_32672,N_32868);
and U33341 (N_33341,N_32839,N_32953);
or U33342 (N_33342,N_32852,N_32700);
or U33343 (N_33343,N_32502,N_32706);
nand U33344 (N_33344,N_32866,N_32971);
nand U33345 (N_33345,N_32640,N_32771);
nand U33346 (N_33346,N_32667,N_32884);
xnor U33347 (N_33347,N_32862,N_32812);
and U33348 (N_33348,N_32765,N_32782);
and U33349 (N_33349,N_32593,N_32773);
and U33350 (N_33350,N_32724,N_32591);
xnor U33351 (N_33351,N_32913,N_32703);
or U33352 (N_33352,N_32966,N_32752);
nand U33353 (N_33353,N_32928,N_32586);
and U33354 (N_33354,N_32561,N_32676);
or U33355 (N_33355,N_32721,N_32563);
or U33356 (N_33356,N_32919,N_32813);
and U33357 (N_33357,N_32720,N_32770);
and U33358 (N_33358,N_32666,N_32603);
or U33359 (N_33359,N_32876,N_32882);
or U33360 (N_33360,N_32733,N_32713);
nand U33361 (N_33361,N_32858,N_32622);
nor U33362 (N_33362,N_32534,N_32725);
or U33363 (N_33363,N_32696,N_32687);
xor U33364 (N_33364,N_32837,N_32655);
and U33365 (N_33365,N_32861,N_32650);
and U33366 (N_33366,N_32776,N_32825);
nand U33367 (N_33367,N_32780,N_32952);
nand U33368 (N_33368,N_32685,N_32935);
nand U33369 (N_33369,N_32792,N_32872);
or U33370 (N_33370,N_32961,N_32786);
and U33371 (N_33371,N_32502,N_32653);
and U33372 (N_33372,N_32781,N_32754);
and U33373 (N_33373,N_32868,N_32758);
and U33374 (N_33374,N_32848,N_32699);
xnor U33375 (N_33375,N_32516,N_32903);
nand U33376 (N_33376,N_32872,N_32734);
and U33377 (N_33377,N_32797,N_32634);
or U33378 (N_33378,N_32509,N_32603);
nor U33379 (N_33379,N_32826,N_32896);
nand U33380 (N_33380,N_32819,N_32500);
nor U33381 (N_33381,N_32673,N_32760);
nor U33382 (N_33382,N_32577,N_32952);
or U33383 (N_33383,N_32879,N_32962);
and U33384 (N_33384,N_32500,N_32896);
nand U33385 (N_33385,N_32524,N_32532);
xor U33386 (N_33386,N_32816,N_32544);
xnor U33387 (N_33387,N_32611,N_32519);
nand U33388 (N_33388,N_32893,N_32803);
and U33389 (N_33389,N_32642,N_32945);
nand U33390 (N_33390,N_32685,N_32630);
xor U33391 (N_33391,N_32633,N_32743);
and U33392 (N_33392,N_32801,N_32871);
xnor U33393 (N_33393,N_32780,N_32801);
xnor U33394 (N_33394,N_32586,N_32862);
and U33395 (N_33395,N_32783,N_32862);
xnor U33396 (N_33396,N_32520,N_32954);
nor U33397 (N_33397,N_32651,N_32742);
nand U33398 (N_33398,N_32934,N_32638);
nor U33399 (N_33399,N_32521,N_32917);
and U33400 (N_33400,N_32867,N_32875);
xor U33401 (N_33401,N_32738,N_32771);
xor U33402 (N_33402,N_32620,N_32716);
nand U33403 (N_33403,N_32559,N_32669);
xor U33404 (N_33404,N_32529,N_32857);
nor U33405 (N_33405,N_32656,N_32950);
and U33406 (N_33406,N_32573,N_32931);
xor U33407 (N_33407,N_32732,N_32743);
xor U33408 (N_33408,N_32626,N_32971);
and U33409 (N_33409,N_32739,N_32539);
nor U33410 (N_33410,N_32580,N_32940);
xor U33411 (N_33411,N_32942,N_32558);
nand U33412 (N_33412,N_32619,N_32752);
nand U33413 (N_33413,N_32862,N_32805);
xnor U33414 (N_33414,N_32810,N_32708);
or U33415 (N_33415,N_32834,N_32726);
xnor U33416 (N_33416,N_32545,N_32514);
and U33417 (N_33417,N_32825,N_32621);
xnor U33418 (N_33418,N_32690,N_32562);
and U33419 (N_33419,N_32740,N_32585);
nor U33420 (N_33420,N_32921,N_32536);
nor U33421 (N_33421,N_32628,N_32553);
and U33422 (N_33422,N_32582,N_32878);
or U33423 (N_33423,N_32526,N_32822);
nor U33424 (N_33424,N_32874,N_32657);
xnor U33425 (N_33425,N_32740,N_32914);
and U33426 (N_33426,N_32724,N_32805);
and U33427 (N_33427,N_32759,N_32540);
or U33428 (N_33428,N_32691,N_32523);
nand U33429 (N_33429,N_32745,N_32651);
and U33430 (N_33430,N_32933,N_32861);
xnor U33431 (N_33431,N_32935,N_32818);
or U33432 (N_33432,N_32548,N_32935);
or U33433 (N_33433,N_32703,N_32513);
and U33434 (N_33434,N_32661,N_32957);
and U33435 (N_33435,N_32747,N_32873);
xor U33436 (N_33436,N_32706,N_32809);
or U33437 (N_33437,N_32703,N_32648);
xnor U33438 (N_33438,N_32657,N_32786);
nand U33439 (N_33439,N_32958,N_32519);
xor U33440 (N_33440,N_32640,N_32926);
and U33441 (N_33441,N_32764,N_32565);
xor U33442 (N_33442,N_32848,N_32969);
and U33443 (N_33443,N_32908,N_32903);
and U33444 (N_33444,N_32634,N_32917);
nand U33445 (N_33445,N_32822,N_32787);
nor U33446 (N_33446,N_32842,N_32571);
xnor U33447 (N_33447,N_32672,N_32934);
and U33448 (N_33448,N_32889,N_32780);
and U33449 (N_33449,N_32733,N_32592);
or U33450 (N_33450,N_32773,N_32609);
nor U33451 (N_33451,N_32558,N_32595);
nor U33452 (N_33452,N_32790,N_32763);
nor U33453 (N_33453,N_32952,N_32801);
or U33454 (N_33454,N_32854,N_32856);
nor U33455 (N_33455,N_32918,N_32623);
or U33456 (N_33456,N_32721,N_32850);
nand U33457 (N_33457,N_32504,N_32735);
nor U33458 (N_33458,N_32980,N_32552);
and U33459 (N_33459,N_32881,N_32926);
nand U33460 (N_33460,N_32677,N_32734);
or U33461 (N_33461,N_32929,N_32658);
nor U33462 (N_33462,N_32583,N_32968);
or U33463 (N_33463,N_32757,N_32955);
or U33464 (N_33464,N_32999,N_32789);
or U33465 (N_33465,N_32598,N_32811);
or U33466 (N_33466,N_32672,N_32998);
nand U33467 (N_33467,N_32745,N_32571);
or U33468 (N_33468,N_32770,N_32936);
xor U33469 (N_33469,N_32951,N_32789);
nand U33470 (N_33470,N_32617,N_32949);
xnor U33471 (N_33471,N_32823,N_32854);
nand U33472 (N_33472,N_32981,N_32606);
or U33473 (N_33473,N_32941,N_32559);
nand U33474 (N_33474,N_32937,N_32948);
xnor U33475 (N_33475,N_32743,N_32680);
xor U33476 (N_33476,N_32608,N_32619);
and U33477 (N_33477,N_32788,N_32569);
nor U33478 (N_33478,N_32938,N_32986);
xnor U33479 (N_33479,N_32919,N_32771);
and U33480 (N_33480,N_32957,N_32684);
and U33481 (N_33481,N_32526,N_32962);
or U33482 (N_33482,N_32566,N_32965);
xnor U33483 (N_33483,N_32881,N_32940);
xnor U33484 (N_33484,N_32992,N_32631);
xnor U33485 (N_33485,N_32528,N_32691);
xnor U33486 (N_33486,N_32905,N_32750);
and U33487 (N_33487,N_32731,N_32879);
nand U33488 (N_33488,N_32720,N_32643);
or U33489 (N_33489,N_32893,N_32796);
nand U33490 (N_33490,N_32970,N_32753);
and U33491 (N_33491,N_32551,N_32696);
and U33492 (N_33492,N_32917,N_32500);
nand U33493 (N_33493,N_32884,N_32970);
and U33494 (N_33494,N_32859,N_32928);
xor U33495 (N_33495,N_32639,N_32504);
or U33496 (N_33496,N_32506,N_32915);
and U33497 (N_33497,N_32723,N_32581);
and U33498 (N_33498,N_32881,N_32704);
xor U33499 (N_33499,N_32521,N_32696);
or U33500 (N_33500,N_33007,N_33452);
and U33501 (N_33501,N_33337,N_33454);
nor U33502 (N_33502,N_33060,N_33308);
and U33503 (N_33503,N_33176,N_33320);
nor U33504 (N_33504,N_33338,N_33271);
or U33505 (N_33505,N_33158,N_33098);
xor U33506 (N_33506,N_33016,N_33023);
or U33507 (N_33507,N_33254,N_33185);
or U33508 (N_33508,N_33301,N_33475);
nor U33509 (N_33509,N_33384,N_33289);
xnor U33510 (N_33510,N_33377,N_33027);
or U33511 (N_33511,N_33412,N_33022);
or U33512 (N_33512,N_33472,N_33351);
or U33513 (N_33513,N_33370,N_33123);
and U33514 (N_33514,N_33434,N_33249);
or U33515 (N_33515,N_33133,N_33479);
and U33516 (N_33516,N_33122,N_33362);
or U33517 (N_33517,N_33152,N_33182);
nor U33518 (N_33518,N_33471,N_33113);
xor U33519 (N_33519,N_33183,N_33467);
xnor U33520 (N_33520,N_33488,N_33364);
and U33521 (N_33521,N_33495,N_33489);
xnor U33522 (N_33522,N_33455,N_33059);
or U33523 (N_33523,N_33040,N_33269);
and U33524 (N_33524,N_33336,N_33312);
and U33525 (N_33525,N_33103,N_33304);
xnor U33526 (N_33526,N_33109,N_33196);
and U33527 (N_33527,N_33374,N_33490);
and U33528 (N_33528,N_33086,N_33418);
xnor U33529 (N_33529,N_33139,N_33095);
nor U33530 (N_33530,N_33356,N_33118);
and U33531 (N_33531,N_33012,N_33339);
nor U33532 (N_33532,N_33078,N_33470);
and U33533 (N_33533,N_33244,N_33033);
xnor U33534 (N_33534,N_33295,N_33409);
or U33535 (N_33535,N_33100,N_33415);
xor U33536 (N_33536,N_33447,N_33230);
and U33537 (N_33537,N_33225,N_33258);
nor U33538 (N_33538,N_33208,N_33314);
xnor U33539 (N_33539,N_33330,N_33044);
or U33540 (N_33540,N_33285,N_33465);
xnor U33541 (N_33541,N_33408,N_33069);
or U33542 (N_33542,N_33353,N_33316);
or U33543 (N_33543,N_33202,N_33063);
xnor U33544 (N_33544,N_33228,N_33165);
xor U33545 (N_33545,N_33021,N_33420);
nand U33546 (N_33546,N_33147,N_33431);
xor U33547 (N_33547,N_33065,N_33270);
nor U33548 (N_33548,N_33449,N_33221);
xnor U33549 (N_33549,N_33045,N_33264);
and U33550 (N_33550,N_33077,N_33001);
or U33551 (N_33551,N_33284,N_33425);
nor U33552 (N_33552,N_33240,N_33138);
and U33553 (N_33553,N_33052,N_33400);
or U33554 (N_33554,N_33127,N_33150);
nand U33555 (N_33555,N_33290,N_33085);
nor U33556 (N_33556,N_33166,N_33019);
or U33557 (N_33557,N_33143,N_33395);
and U33558 (N_33558,N_33005,N_33126);
or U33559 (N_33559,N_33499,N_33256);
xor U33560 (N_33560,N_33392,N_33481);
nor U33561 (N_33561,N_33232,N_33004);
xor U33562 (N_33562,N_33432,N_33048);
or U33563 (N_33563,N_33288,N_33000);
xor U33564 (N_33564,N_33198,N_33410);
and U33565 (N_33565,N_33051,N_33006);
xnor U33566 (N_33566,N_33421,N_33298);
or U33567 (N_33567,N_33383,N_33056);
or U33568 (N_33568,N_33154,N_33193);
and U33569 (N_33569,N_33219,N_33419);
nand U33570 (N_33570,N_33307,N_33076);
xnor U33571 (N_33571,N_33414,N_33087);
xnor U33572 (N_33572,N_33486,N_33061);
nand U33573 (N_33573,N_33120,N_33387);
nor U33574 (N_33574,N_33020,N_33363);
nor U33575 (N_33575,N_33009,N_33468);
nand U33576 (N_33576,N_33313,N_33318);
or U33577 (N_33577,N_33135,N_33112);
nor U33578 (N_33578,N_33426,N_33071);
xnor U33579 (N_33579,N_33132,N_33178);
or U33580 (N_33580,N_33203,N_33277);
xnor U33581 (N_33581,N_33382,N_33391);
or U33582 (N_33582,N_33393,N_33360);
nand U33583 (N_33583,N_33204,N_33278);
nor U33584 (N_33584,N_33101,N_33119);
xnor U33585 (N_33585,N_33011,N_33276);
or U33586 (N_33586,N_33218,N_33429);
xor U33587 (N_33587,N_33014,N_33174);
nand U33588 (N_33588,N_33042,N_33032);
or U33589 (N_33589,N_33261,N_33124);
xnor U33590 (N_33590,N_33036,N_33046);
nand U33591 (N_33591,N_33246,N_33188);
xnor U33592 (N_33592,N_33145,N_33441);
or U33593 (N_33593,N_33149,N_33229);
and U33594 (N_33594,N_33241,N_33070);
nand U33595 (N_33595,N_33283,N_33030);
and U33596 (N_33596,N_33235,N_33025);
nor U33597 (N_33597,N_33247,N_33398);
nand U33598 (N_33598,N_33034,N_33309);
nor U33599 (N_33599,N_33265,N_33252);
xor U33600 (N_33600,N_33068,N_33179);
nand U33601 (N_33601,N_33168,N_33137);
xnor U33602 (N_33602,N_33177,N_33315);
xor U33603 (N_33603,N_33136,N_33456);
and U33604 (N_33604,N_33194,N_33236);
and U33605 (N_33605,N_33024,N_33453);
nor U33606 (N_33606,N_33080,N_33195);
nand U33607 (N_33607,N_33368,N_33379);
and U33608 (N_33608,N_33212,N_33376);
and U33609 (N_33609,N_33233,N_33496);
and U33610 (N_33610,N_33107,N_33057);
or U33611 (N_33611,N_33237,N_33348);
xor U33612 (N_33612,N_33028,N_33116);
and U33613 (N_33613,N_33220,N_33280);
or U33614 (N_33614,N_33227,N_33350);
and U33615 (N_33615,N_33342,N_33155);
or U33616 (N_33616,N_33494,N_33401);
and U33617 (N_33617,N_33172,N_33018);
and U33618 (N_33618,N_33164,N_33192);
nor U33619 (N_33619,N_33482,N_33319);
or U33620 (N_33620,N_33389,N_33476);
nand U33621 (N_33621,N_33074,N_33037);
nand U33622 (N_33622,N_33157,N_33324);
xnor U33623 (N_33623,N_33451,N_33303);
or U33624 (N_33624,N_33413,N_33416);
or U33625 (N_33625,N_33015,N_33201);
nor U33626 (N_33626,N_33478,N_33210);
nor U33627 (N_33627,N_33458,N_33366);
or U33628 (N_33628,N_33187,N_33491);
nor U33629 (N_33629,N_33073,N_33444);
or U33630 (N_33630,N_33081,N_33106);
or U33631 (N_33631,N_33373,N_33343);
xnor U33632 (N_33632,N_33231,N_33438);
nand U33633 (N_33633,N_33114,N_33224);
or U33634 (N_33634,N_33072,N_33128);
and U33635 (N_33635,N_33485,N_33251);
nor U33636 (N_33636,N_33422,N_33492);
or U33637 (N_33637,N_33305,N_33245);
and U33638 (N_33638,N_33053,N_33323);
xnor U33639 (N_33639,N_33129,N_33347);
nor U33640 (N_33640,N_33222,N_33099);
and U33641 (N_33641,N_33215,N_33281);
or U33642 (N_33642,N_33002,N_33105);
and U33643 (N_33643,N_33260,N_33175);
and U33644 (N_33644,N_33206,N_33255);
and U33645 (N_33645,N_33423,N_33017);
nor U33646 (N_33646,N_33405,N_33144);
nor U33647 (N_33647,N_33250,N_33010);
xor U33648 (N_33648,N_33248,N_33075);
xnor U33649 (N_33649,N_33321,N_33142);
or U33650 (N_33650,N_33067,N_33209);
xnor U33651 (N_33651,N_33365,N_33029);
xor U33652 (N_33652,N_33197,N_33153);
and U33653 (N_33653,N_33117,N_33160);
and U33654 (N_33654,N_33013,N_33386);
nor U33655 (N_33655,N_33341,N_33424);
nand U33656 (N_33656,N_33167,N_33340);
xor U33657 (N_33657,N_33151,N_33043);
and U33658 (N_33658,N_33125,N_33039);
or U33659 (N_33659,N_33066,N_33131);
or U33660 (N_33660,N_33058,N_33403);
nor U33661 (N_33661,N_33399,N_33311);
nand U33662 (N_33662,N_33190,N_33189);
nand U33663 (N_33663,N_33430,N_33367);
or U33664 (N_33664,N_33170,N_33091);
nand U33665 (N_33665,N_33273,N_33439);
or U33666 (N_33666,N_33262,N_33450);
nand U33667 (N_33667,N_33322,N_33388);
nand U33668 (N_33668,N_33079,N_33031);
and U33669 (N_33669,N_33358,N_33442);
and U33670 (N_33670,N_33417,N_33146);
or U33671 (N_33671,N_33180,N_33089);
xnor U33672 (N_33672,N_33286,N_33361);
or U33673 (N_33673,N_33092,N_33480);
or U33674 (N_33674,N_33159,N_33497);
xnor U33675 (N_33675,N_33243,N_33108);
or U33676 (N_33676,N_33104,N_33349);
nor U33677 (N_33677,N_33448,N_33357);
or U33678 (N_33678,N_33083,N_33205);
nand U33679 (N_33679,N_33428,N_33390);
or U33680 (N_33680,N_33272,N_33263);
nand U33681 (N_33681,N_33207,N_33473);
and U33682 (N_33682,N_33211,N_33162);
and U33683 (N_33683,N_33064,N_33306);
nand U33684 (N_33684,N_33084,N_33437);
xor U33685 (N_33685,N_33186,N_33094);
nand U33686 (N_33686,N_33385,N_33234);
xor U33687 (N_33687,N_33433,N_33474);
and U33688 (N_33688,N_33460,N_33082);
or U33689 (N_33689,N_33394,N_33381);
nand U33690 (N_33690,N_33161,N_33335);
nand U33691 (N_33691,N_33375,N_33354);
xnor U33692 (N_33692,N_33242,N_33140);
nand U33693 (N_33693,N_33477,N_33445);
xor U33694 (N_33694,N_33096,N_33008);
or U33695 (N_33695,N_33191,N_33291);
or U33696 (N_33696,N_33169,N_33216);
xnor U33697 (N_33697,N_33110,N_33466);
xor U33698 (N_33698,N_33292,N_33090);
or U33699 (N_33699,N_33371,N_33333);
nor U33700 (N_33700,N_33464,N_33498);
xnor U33701 (N_33701,N_33047,N_33493);
xnor U33702 (N_33702,N_33462,N_33440);
nand U33703 (N_33703,N_33300,N_33130);
and U33704 (N_33704,N_33093,N_33055);
nand U33705 (N_33705,N_33487,N_33334);
and U33706 (N_33706,N_33436,N_33181);
or U33707 (N_33707,N_33253,N_33310);
nor U33708 (N_33708,N_33279,N_33294);
or U33709 (N_33709,N_33331,N_33097);
or U33710 (N_33710,N_33378,N_33049);
nor U33711 (N_33711,N_33050,N_33443);
and U33712 (N_33712,N_33184,N_33275);
and U33713 (N_33713,N_33327,N_33459);
nand U33714 (N_33714,N_33111,N_33346);
xor U33715 (N_33715,N_33328,N_33163);
or U33716 (N_33716,N_33293,N_33282);
and U33717 (N_33717,N_33266,N_33239);
nor U33718 (N_33718,N_33088,N_33296);
and U33719 (N_33719,N_33062,N_33317);
or U33720 (N_33720,N_33287,N_33380);
and U33721 (N_33721,N_33035,N_33121);
nor U33722 (N_33722,N_33226,N_33329);
xor U33723 (N_33723,N_33435,N_33446);
nor U33724 (N_33724,N_33268,N_33171);
or U33725 (N_33725,N_33404,N_33427);
nand U33726 (N_33726,N_33359,N_33483);
xnor U33727 (N_33727,N_33259,N_33214);
nor U33728 (N_33728,N_33200,N_33134);
xor U33729 (N_33729,N_33325,N_33297);
and U33730 (N_33730,N_33173,N_33397);
xor U33731 (N_33731,N_33461,N_33355);
or U33732 (N_33732,N_33332,N_33156);
and U33733 (N_33733,N_33463,N_33148);
and U33734 (N_33734,N_33238,N_33369);
and U33735 (N_33735,N_33326,N_33102);
and U33736 (N_33736,N_33257,N_33223);
nor U33737 (N_33737,N_33299,N_33026);
nand U33738 (N_33738,N_33141,N_33344);
or U33739 (N_33739,N_33038,N_33457);
nor U33740 (N_33740,N_33003,N_33054);
or U33741 (N_33741,N_33345,N_33217);
or U33742 (N_33742,N_33274,N_33199);
nor U33743 (N_33743,N_33469,N_33402);
nand U33744 (N_33744,N_33396,N_33406);
nor U33745 (N_33745,N_33411,N_33484);
or U33746 (N_33746,N_33352,N_33302);
and U33747 (N_33747,N_33041,N_33115);
or U33748 (N_33748,N_33407,N_33372);
nor U33749 (N_33749,N_33213,N_33267);
xor U33750 (N_33750,N_33472,N_33371);
nand U33751 (N_33751,N_33330,N_33218);
or U33752 (N_33752,N_33168,N_33199);
and U33753 (N_33753,N_33485,N_33093);
or U33754 (N_33754,N_33078,N_33135);
nand U33755 (N_33755,N_33438,N_33420);
xnor U33756 (N_33756,N_33155,N_33244);
nand U33757 (N_33757,N_33422,N_33318);
nor U33758 (N_33758,N_33261,N_33324);
and U33759 (N_33759,N_33186,N_33001);
xor U33760 (N_33760,N_33286,N_33292);
nand U33761 (N_33761,N_33196,N_33375);
nand U33762 (N_33762,N_33448,N_33350);
or U33763 (N_33763,N_33464,N_33495);
and U33764 (N_33764,N_33471,N_33332);
xnor U33765 (N_33765,N_33257,N_33339);
or U33766 (N_33766,N_33013,N_33463);
and U33767 (N_33767,N_33330,N_33216);
or U33768 (N_33768,N_33275,N_33201);
or U33769 (N_33769,N_33378,N_33201);
nand U33770 (N_33770,N_33016,N_33203);
or U33771 (N_33771,N_33488,N_33391);
nand U33772 (N_33772,N_33301,N_33227);
or U33773 (N_33773,N_33491,N_33478);
xor U33774 (N_33774,N_33220,N_33338);
nand U33775 (N_33775,N_33337,N_33134);
and U33776 (N_33776,N_33213,N_33042);
nor U33777 (N_33777,N_33437,N_33021);
nor U33778 (N_33778,N_33237,N_33477);
or U33779 (N_33779,N_33070,N_33198);
or U33780 (N_33780,N_33265,N_33248);
or U33781 (N_33781,N_33245,N_33499);
or U33782 (N_33782,N_33043,N_33192);
nor U33783 (N_33783,N_33037,N_33423);
or U33784 (N_33784,N_33051,N_33275);
or U33785 (N_33785,N_33411,N_33425);
nor U33786 (N_33786,N_33417,N_33032);
nand U33787 (N_33787,N_33413,N_33155);
nor U33788 (N_33788,N_33030,N_33160);
xnor U33789 (N_33789,N_33177,N_33450);
or U33790 (N_33790,N_33226,N_33413);
and U33791 (N_33791,N_33132,N_33186);
or U33792 (N_33792,N_33059,N_33122);
nand U33793 (N_33793,N_33264,N_33100);
and U33794 (N_33794,N_33273,N_33031);
and U33795 (N_33795,N_33395,N_33026);
nor U33796 (N_33796,N_33484,N_33078);
nand U33797 (N_33797,N_33375,N_33194);
nand U33798 (N_33798,N_33047,N_33058);
nand U33799 (N_33799,N_33433,N_33260);
and U33800 (N_33800,N_33152,N_33431);
xnor U33801 (N_33801,N_33489,N_33115);
or U33802 (N_33802,N_33478,N_33017);
nor U33803 (N_33803,N_33233,N_33161);
or U33804 (N_33804,N_33333,N_33109);
xor U33805 (N_33805,N_33079,N_33278);
or U33806 (N_33806,N_33387,N_33213);
or U33807 (N_33807,N_33428,N_33484);
nand U33808 (N_33808,N_33432,N_33382);
or U33809 (N_33809,N_33160,N_33340);
or U33810 (N_33810,N_33454,N_33370);
xor U33811 (N_33811,N_33055,N_33048);
or U33812 (N_33812,N_33385,N_33213);
xnor U33813 (N_33813,N_33342,N_33273);
nand U33814 (N_33814,N_33440,N_33452);
and U33815 (N_33815,N_33108,N_33087);
nor U33816 (N_33816,N_33483,N_33097);
nor U33817 (N_33817,N_33311,N_33268);
nand U33818 (N_33818,N_33218,N_33179);
xor U33819 (N_33819,N_33193,N_33129);
or U33820 (N_33820,N_33499,N_33298);
nor U33821 (N_33821,N_33329,N_33089);
and U33822 (N_33822,N_33046,N_33396);
and U33823 (N_33823,N_33060,N_33429);
and U33824 (N_33824,N_33435,N_33470);
nor U33825 (N_33825,N_33040,N_33071);
nor U33826 (N_33826,N_33060,N_33049);
xor U33827 (N_33827,N_33249,N_33107);
or U33828 (N_33828,N_33451,N_33350);
and U33829 (N_33829,N_33206,N_33389);
or U33830 (N_33830,N_33285,N_33165);
or U33831 (N_33831,N_33131,N_33332);
nor U33832 (N_33832,N_33184,N_33042);
xnor U33833 (N_33833,N_33372,N_33086);
nand U33834 (N_33834,N_33398,N_33269);
xor U33835 (N_33835,N_33245,N_33274);
nand U33836 (N_33836,N_33492,N_33221);
nand U33837 (N_33837,N_33141,N_33130);
nor U33838 (N_33838,N_33409,N_33269);
and U33839 (N_33839,N_33054,N_33462);
nand U33840 (N_33840,N_33453,N_33311);
xor U33841 (N_33841,N_33326,N_33172);
or U33842 (N_33842,N_33131,N_33027);
and U33843 (N_33843,N_33130,N_33489);
and U33844 (N_33844,N_33224,N_33380);
nor U33845 (N_33845,N_33084,N_33367);
and U33846 (N_33846,N_33342,N_33071);
nand U33847 (N_33847,N_33137,N_33355);
and U33848 (N_33848,N_33127,N_33489);
or U33849 (N_33849,N_33069,N_33260);
nor U33850 (N_33850,N_33339,N_33165);
xnor U33851 (N_33851,N_33237,N_33281);
nor U33852 (N_33852,N_33335,N_33397);
and U33853 (N_33853,N_33422,N_33379);
or U33854 (N_33854,N_33159,N_33113);
nor U33855 (N_33855,N_33028,N_33354);
and U33856 (N_33856,N_33039,N_33095);
and U33857 (N_33857,N_33104,N_33249);
nand U33858 (N_33858,N_33495,N_33398);
and U33859 (N_33859,N_33225,N_33008);
or U33860 (N_33860,N_33381,N_33031);
nor U33861 (N_33861,N_33435,N_33099);
nor U33862 (N_33862,N_33294,N_33333);
or U33863 (N_33863,N_33046,N_33062);
nand U33864 (N_33864,N_33226,N_33440);
nand U33865 (N_33865,N_33475,N_33356);
and U33866 (N_33866,N_33398,N_33365);
and U33867 (N_33867,N_33097,N_33366);
nor U33868 (N_33868,N_33242,N_33361);
or U33869 (N_33869,N_33435,N_33052);
nor U33870 (N_33870,N_33253,N_33395);
or U33871 (N_33871,N_33286,N_33109);
xor U33872 (N_33872,N_33389,N_33180);
or U33873 (N_33873,N_33408,N_33033);
and U33874 (N_33874,N_33046,N_33001);
xor U33875 (N_33875,N_33027,N_33040);
or U33876 (N_33876,N_33031,N_33255);
nor U33877 (N_33877,N_33409,N_33177);
or U33878 (N_33878,N_33495,N_33272);
and U33879 (N_33879,N_33381,N_33342);
or U33880 (N_33880,N_33373,N_33160);
nor U33881 (N_33881,N_33381,N_33372);
and U33882 (N_33882,N_33005,N_33475);
and U33883 (N_33883,N_33351,N_33439);
and U33884 (N_33884,N_33003,N_33427);
and U33885 (N_33885,N_33054,N_33129);
and U33886 (N_33886,N_33092,N_33071);
or U33887 (N_33887,N_33300,N_33295);
nand U33888 (N_33888,N_33497,N_33444);
nor U33889 (N_33889,N_33266,N_33218);
nor U33890 (N_33890,N_33019,N_33012);
and U33891 (N_33891,N_33296,N_33389);
nand U33892 (N_33892,N_33452,N_33160);
xor U33893 (N_33893,N_33138,N_33401);
nor U33894 (N_33894,N_33128,N_33376);
nor U33895 (N_33895,N_33089,N_33319);
or U33896 (N_33896,N_33303,N_33289);
nand U33897 (N_33897,N_33168,N_33447);
nand U33898 (N_33898,N_33052,N_33151);
nand U33899 (N_33899,N_33442,N_33031);
nand U33900 (N_33900,N_33464,N_33410);
nor U33901 (N_33901,N_33032,N_33153);
nor U33902 (N_33902,N_33388,N_33420);
and U33903 (N_33903,N_33403,N_33148);
nor U33904 (N_33904,N_33313,N_33029);
xor U33905 (N_33905,N_33482,N_33405);
and U33906 (N_33906,N_33104,N_33256);
xnor U33907 (N_33907,N_33378,N_33306);
nand U33908 (N_33908,N_33013,N_33475);
or U33909 (N_33909,N_33047,N_33260);
xor U33910 (N_33910,N_33191,N_33345);
and U33911 (N_33911,N_33370,N_33263);
xnor U33912 (N_33912,N_33263,N_33492);
nand U33913 (N_33913,N_33288,N_33001);
nor U33914 (N_33914,N_33073,N_33478);
nor U33915 (N_33915,N_33498,N_33034);
and U33916 (N_33916,N_33414,N_33170);
nor U33917 (N_33917,N_33095,N_33356);
nand U33918 (N_33918,N_33311,N_33022);
nor U33919 (N_33919,N_33295,N_33123);
or U33920 (N_33920,N_33167,N_33126);
xor U33921 (N_33921,N_33485,N_33078);
and U33922 (N_33922,N_33327,N_33360);
or U33923 (N_33923,N_33358,N_33207);
xor U33924 (N_33924,N_33084,N_33486);
xor U33925 (N_33925,N_33198,N_33008);
nand U33926 (N_33926,N_33099,N_33389);
and U33927 (N_33927,N_33174,N_33111);
nor U33928 (N_33928,N_33149,N_33021);
or U33929 (N_33929,N_33491,N_33318);
and U33930 (N_33930,N_33489,N_33128);
nand U33931 (N_33931,N_33335,N_33015);
xor U33932 (N_33932,N_33173,N_33408);
and U33933 (N_33933,N_33080,N_33424);
nand U33934 (N_33934,N_33444,N_33155);
nor U33935 (N_33935,N_33495,N_33271);
or U33936 (N_33936,N_33485,N_33358);
xor U33937 (N_33937,N_33339,N_33390);
or U33938 (N_33938,N_33262,N_33313);
nor U33939 (N_33939,N_33111,N_33007);
and U33940 (N_33940,N_33020,N_33287);
nand U33941 (N_33941,N_33148,N_33032);
and U33942 (N_33942,N_33313,N_33423);
xor U33943 (N_33943,N_33469,N_33388);
or U33944 (N_33944,N_33192,N_33140);
or U33945 (N_33945,N_33200,N_33102);
nand U33946 (N_33946,N_33335,N_33251);
and U33947 (N_33947,N_33450,N_33364);
nor U33948 (N_33948,N_33155,N_33069);
nand U33949 (N_33949,N_33444,N_33076);
xor U33950 (N_33950,N_33070,N_33416);
and U33951 (N_33951,N_33440,N_33359);
nor U33952 (N_33952,N_33379,N_33011);
and U33953 (N_33953,N_33477,N_33102);
or U33954 (N_33954,N_33153,N_33250);
xor U33955 (N_33955,N_33299,N_33129);
nor U33956 (N_33956,N_33369,N_33116);
and U33957 (N_33957,N_33442,N_33409);
and U33958 (N_33958,N_33427,N_33341);
and U33959 (N_33959,N_33267,N_33367);
and U33960 (N_33960,N_33106,N_33444);
nor U33961 (N_33961,N_33100,N_33228);
xnor U33962 (N_33962,N_33161,N_33239);
xor U33963 (N_33963,N_33106,N_33434);
xnor U33964 (N_33964,N_33347,N_33379);
and U33965 (N_33965,N_33154,N_33161);
nand U33966 (N_33966,N_33058,N_33445);
nor U33967 (N_33967,N_33201,N_33029);
nand U33968 (N_33968,N_33389,N_33041);
nor U33969 (N_33969,N_33258,N_33161);
nand U33970 (N_33970,N_33361,N_33439);
nor U33971 (N_33971,N_33116,N_33038);
nand U33972 (N_33972,N_33431,N_33397);
xor U33973 (N_33973,N_33442,N_33494);
nand U33974 (N_33974,N_33236,N_33260);
xnor U33975 (N_33975,N_33492,N_33319);
nor U33976 (N_33976,N_33469,N_33206);
nor U33977 (N_33977,N_33180,N_33499);
and U33978 (N_33978,N_33011,N_33279);
and U33979 (N_33979,N_33156,N_33430);
and U33980 (N_33980,N_33480,N_33161);
nor U33981 (N_33981,N_33261,N_33327);
and U33982 (N_33982,N_33158,N_33264);
or U33983 (N_33983,N_33046,N_33415);
and U33984 (N_33984,N_33166,N_33076);
nor U33985 (N_33985,N_33448,N_33020);
nor U33986 (N_33986,N_33257,N_33146);
nand U33987 (N_33987,N_33165,N_33061);
and U33988 (N_33988,N_33367,N_33369);
nor U33989 (N_33989,N_33117,N_33019);
nand U33990 (N_33990,N_33404,N_33441);
xor U33991 (N_33991,N_33046,N_33312);
nand U33992 (N_33992,N_33108,N_33133);
nor U33993 (N_33993,N_33219,N_33467);
or U33994 (N_33994,N_33261,N_33464);
and U33995 (N_33995,N_33146,N_33345);
nor U33996 (N_33996,N_33443,N_33453);
xnor U33997 (N_33997,N_33400,N_33219);
or U33998 (N_33998,N_33349,N_33160);
nand U33999 (N_33999,N_33116,N_33196);
and U34000 (N_34000,N_33705,N_33893);
and U34001 (N_34001,N_33833,N_33726);
xor U34002 (N_34002,N_33891,N_33764);
nor U34003 (N_34003,N_33921,N_33791);
nor U34004 (N_34004,N_33771,N_33665);
or U34005 (N_34005,N_33751,N_33901);
or U34006 (N_34006,N_33863,N_33699);
xnor U34007 (N_34007,N_33508,N_33558);
and U34008 (N_34008,N_33523,N_33760);
and U34009 (N_34009,N_33567,N_33814);
xnor U34010 (N_34010,N_33526,N_33533);
nand U34011 (N_34011,N_33664,N_33974);
or U34012 (N_34012,N_33953,N_33715);
nand U34013 (N_34013,N_33511,N_33939);
or U34014 (N_34014,N_33542,N_33720);
nor U34015 (N_34015,N_33604,N_33871);
xnor U34016 (N_34016,N_33972,N_33849);
nand U34017 (N_34017,N_33827,N_33842);
xor U34018 (N_34018,N_33870,N_33808);
nand U34019 (N_34019,N_33589,N_33765);
nor U34020 (N_34020,N_33584,N_33860);
nor U34021 (N_34021,N_33884,N_33971);
xor U34022 (N_34022,N_33718,N_33634);
and U34023 (N_34023,N_33928,N_33988);
xnor U34024 (N_34024,N_33740,N_33596);
and U34025 (N_34025,N_33835,N_33630);
nor U34026 (N_34026,N_33735,N_33894);
nor U34027 (N_34027,N_33976,N_33631);
xor U34028 (N_34028,N_33609,N_33600);
and U34029 (N_34029,N_33668,N_33745);
nor U34030 (N_34030,N_33557,N_33970);
nor U34031 (N_34031,N_33637,N_33982);
xnor U34032 (N_34032,N_33969,N_33963);
nand U34033 (N_34033,N_33981,N_33749);
and U34034 (N_34034,N_33859,N_33626);
nor U34035 (N_34035,N_33978,N_33979);
nand U34036 (N_34036,N_33962,N_33758);
nor U34037 (N_34037,N_33714,N_33992);
or U34038 (N_34038,N_33582,N_33638);
xor U34039 (N_34039,N_33537,N_33704);
nand U34040 (N_34040,N_33728,N_33941);
xor U34041 (N_34041,N_33580,N_33995);
and U34042 (N_34042,N_33551,N_33524);
nand U34043 (N_34043,N_33673,N_33856);
xnor U34044 (N_34044,N_33964,N_33581);
nor U34045 (N_34045,N_33539,N_33920);
and U34046 (N_34046,N_33651,N_33773);
nand U34047 (N_34047,N_33563,N_33815);
xnor U34048 (N_34048,N_33877,N_33913);
nor U34049 (N_34049,N_33676,N_33989);
and U34050 (N_34050,N_33555,N_33876);
nand U34051 (N_34051,N_33807,N_33883);
nor U34052 (N_34052,N_33938,N_33624);
xnor U34053 (N_34053,N_33927,N_33690);
or U34054 (N_34054,N_33657,N_33691);
nand U34055 (N_34055,N_33506,N_33512);
nand U34056 (N_34056,N_33597,N_33510);
or U34057 (N_34057,N_33959,N_33850);
nand U34058 (N_34058,N_33552,N_33578);
nor U34059 (N_34059,N_33830,N_33899);
and U34060 (N_34060,N_33944,N_33812);
nor U34061 (N_34061,N_33940,N_33906);
nand U34062 (N_34062,N_33579,N_33562);
nand U34063 (N_34063,N_33924,N_33824);
and U34064 (N_34064,N_33618,N_33683);
xor U34065 (N_34065,N_33732,N_33711);
xor U34066 (N_34066,N_33783,N_33559);
nand U34067 (N_34067,N_33753,N_33900);
xnor U34068 (N_34068,N_33525,N_33514);
or U34069 (N_34069,N_33937,N_33646);
and U34070 (N_34070,N_33809,N_33892);
xnor U34071 (N_34071,N_33547,N_33535);
nand U34072 (N_34072,N_33606,N_33887);
and U34073 (N_34073,N_33810,N_33687);
nand U34074 (N_34074,N_33566,N_33724);
and U34075 (N_34075,N_33952,N_33702);
nand U34076 (N_34076,N_33588,N_33549);
nor U34077 (N_34077,N_33583,N_33922);
nor U34078 (N_34078,N_33832,N_33528);
nand U34079 (N_34079,N_33518,N_33957);
xor U34080 (N_34080,N_33793,N_33532);
and U34081 (N_34081,N_33569,N_33980);
nand U34082 (N_34082,N_33727,N_33917);
and U34083 (N_34083,N_33990,N_33916);
or U34084 (N_34084,N_33688,N_33722);
nand U34085 (N_34085,N_33905,N_33909);
or U34086 (N_34086,N_33674,N_33775);
and U34087 (N_34087,N_33541,N_33954);
and U34088 (N_34088,N_33741,N_33858);
and U34089 (N_34089,N_33534,N_33520);
nor U34090 (N_34090,N_33748,N_33947);
and U34091 (N_34091,N_33786,N_33666);
or U34092 (N_34092,N_33650,N_33544);
and U34093 (N_34093,N_33521,N_33930);
nand U34094 (N_34094,N_33986,N_33813);
nor U34095 (N_34095,N_33966,N_33782);
or U34096 (N_34096,N_33693,N_33914);
and U34097 (N_34097,N_33878,N_33872);
xnor U34098 (N_34098,N_33627,N_33737);
xor U34099 (N_34099,N_33647,N_33632);
nand U34100 (N_34100,N_33703,N_33854);
and U34101 (N_34101,N_33586,N_33902);
and U34102 (N_34102,N_33507,N_33848);
or U34103 (N_34103,N_33671,N_33866);
and U34104 (N_34104,N_33656,N_33910);
xor U34105 (N_34105,N_33698,N_33785);
xor U34106 (N_34106,N_33923,N_33948);
nor U34107 (N_34107,N_33649,N_33853);
nand U34108 (N_34108,N_33912,N_33999);
or U34109 (N_34109,N_33955,N_33795);
xor U34110 (N_34110,N_33843,N_33709);
nand U34111 (N_34111,N_33767,N_33847);
and U34112 (N_34112,N_33502,N_33756);
nor U34113 (N_34113,N_33961,N_33678);
nand U34114 (N_34114,N_33874,N_33540);
xor U34115 (N_34115,N_33769,N_33820);
and U34116 (N_34116,N_33716,N_33772);
nand U34117 (N_34117,N_33529,N_33774);
xnor U34118 (N_34118,N_33919,N_33811);
and U34119 (N_34119,N_33790,N_33846);
nand U34120 (N_34120,N_33652,N_33680);
and U34121 (N_34121,N_33573,N_33743);
xor U34122 (N_34122,N_33513,N_33757);
or U34123 (N_34123,N_33956,N_33677);
nand U34124 (N_34124,N_33763,N_33788);
or U34125 (N_34125,N_33958,N_33752);
and U34126 (N_34126,N_33733,N_33951);
xor U34127 (N_34127,N_33610,N_33779);
or U34128 (N_34128,N_33991,N_33550);
xnor U34129 (N_34129,N_33519,N_33780);
and U34130 (N_34130,N_33831,N_33682);
nor U34131 (N_34131,N_33985,N_33868);
nand U34132 (N_34132,N_33837,N_33929);
or U34133 (N_34133,N_33516,N_33725);
and U34134 (N_34134,N_33554,N_33823);
nand U34135 (N_34135,N_33770,N_33864);
or U34136 (N_34136,N_33967,N_33857);
or U34137 (N_34137,N_33568,N_33731);
xnor U34138 (N_34138,N_33911,N_33655);
xor U34139 (N_34139,N_33661,N_33706);
nor U34140 (N_34140,N_33625,N_33907);
or U34141 (N_34141,N_33590,N_33708);
nand U34142 (N_34142,N_33645,N_33926);
nor U34143 (N_34143,N_33681,N_33816);
xnor U34144 (N_34144,N_33710,N_33766);
or U34145 (N_34145,N_33908,N_33641);
xor U34146 (N_34146,N_33619,N_33796);
nor U34147 (N_34147,N_33603,N_33792);
and U34148 (N_34148,N_33505,N_33742);
or U34149 (N_34149,N_33615,N_33977);
nand U34150 (N_34150,N_33997,N_33915);
nor U34151 (N_34151,N_33623,N_33897);
nand U34152 (N_34152,N_33801,N_33660);
nor U34153 (N_34153,N_33889,N_33784);
or U34154 (N_34154,N_33851,N_33781);
nand U34155 (N_34155,N_33755,N_33594);
nor U34156 (N_34156,N_33895,N_33515);
or U34157 (N_34157,N_33548,N_33746);
or U34158 (N_34158,N_33778,N_33734);
or U34159 (N_34159,N_33888,N_33598);
or U34160 (N_34160,N_33662,N_33822);
nand U34161 (N_34161,N_33730,N_33806);
or U34162 (N_34162,N_33560,N_33684);
nand U34163 (N_34163,N_33918,N_33570);
and U34164 (N_34164,N_33576,N_33669);
nand U34165 (N_34165,N_33949,N_33828);
nor U34166 (N_34166,N_33933,N_33836);
and U34167 (N_34167,N_33636,N_33564);
nand U34168 (N_34168,N_33865,N_33571);
xnor U34169 (N_34169,N_33546,N_33601);
or U34170 (N_34170,N_33613,N_33696);
and U34171 (N_34171,N_33761,N_33852);
xnor U34172 (N_34172,N_33768,N_33993);
nand U34173 (N_34173,N_33943,N_33736);
xor U34174 (N_34174,N_33595,N_33607);
nor U34175 (N_34175,N_33994,N_33719);
nor U34176 (N_34176,N_33592,N_33577);
nand U34177 (N_34177,N_33501,N_33983);
nand U34178 (N_34178,N_33574,N_33500);
xnor U34179 (N_34179,N_33886,N_33712);
or U34180 (N_34180,N_33739,N_33531);
and U34181 (N_34181,N_33617,N_33628);
xor U34182 (N_34182,N_33804,N_33965);
nor U34183 (N_34183,N_33679,N_33862);
or U34184 (N_34184,N_33925,N_33935);
xnor U34185 (N_34185,N_33629,N_33565);
and U34186 (N_34186,N_33762,N_33984);
or U34187 (N_34187,N_33729,N_33553);
nor U34188 (N_34188,N_33975,N_33701);
nor U34189 (N_34189,N_33840,N_33643);
nor U34190 (N_34190,N_33844,N_33898);
xor U34191 (N_34191,N_33838,N_33819);
nor U34192 (N_34192,N_33659,N_33721);
or U34193 (N_34193,N_33572,N_33616);
nand U34194 (N_34194,N_33653,N_33517);
nand U34195 (N_34195,N_33799,N_33834);
xnor U34196 (N_34196,N_33612,N_33882);
or U34197 (N_34197,N_33587,N_33904);
or U34198 (N_34198,N_33973,N_33996);
nand U34199 (N_34199,N_33880,N_33946);
xnor U34200 (N_34200,N_33538,N_33585);
or U34201 (N_34201,N_33504,N_33713);
nor U34202 (N_34202,N_33803,N_33556);
or U34203 (N_34203,N_33707,N_33530);
and U34204 (N_34204,N_33670,N_33658);
or U34205 (N_34205,N_33942,N_33503);
nand U34206 (N_34206,N_33509,N_33821);
nor U34207 (N_34207,N_33692,N_33945);
nor U34208 (N_34208,N_33861,N_33817);
and U34209 (N_34209,N_33675,N_33960);
xnor U34210 (N_34210,N_33744,N_33561);
nor U34211 (N_34211,N_33841,N_33931);
xor U34212 (N_34212,N_33845,N_33934);
nand U34213 (N_34213,N_33695,N_33620);
or U34214 (N_34214,N_33777,N_33903);
or U34215 (N_34215,N_33789,N_33672);
xnor U34216 (N_34216,N_33611,N_33802);
and U34217 (N_34217,N_33717,N_33593);
nor U34218 (N_34218,N_33879,N_33527);
nor U34219 (N_34219,N_33968,N_33543);
nand U34220 (N_34220,N_33747,N_33787);
and U34221 (N_34221,N_33738,N_33697);
nor U34222 (N_34222,N_33633,N_33798);
nor U34223 (N_34223,N_33826,N_33754);
nand U34224 (N_34224,N_33855,N_33750);
nand U34225 (N_34225,N_33950,N_33591);
nor U34226 (N_34226,N_33522,N_33885);
xor U34227 (N_34227,N_33686,N_33622);
or U34228 (N_34228,N_33881,N_33869);
or U34229 (N_34229,N_33536,N_33896);
and U34230 (N_34230,N_33700,N_33575);
nor U34231 (N_34231,N_33602,N_33605);
and U34232 (N_34232,N_33776,N_33797);
and U34233 (N_34233,N_33621,N_33599);
and U34234 (N_34234,N_33818,N_33873);
nor U34235 (N_34235,N_33829,N_33936);
nor U34236 (N_34236,N_33998,N_33663);
or U34237 (N_34237,N_33825,N_33689);
nor U34238 (N_34238,N_33639,N_33685);
or U34239 (N_34239,N_33987,N_33759);
xnor U34240 (N_34240,N_33635,N_33839);
and U34241 (N_34241,N_33667,N_33694);
or U34242 (N_34242,N_33794,N_33723);
nand U34243 (N_34243,N_33654,N_33640);
xnor U34244 (N_34244,N_33644,N_33867);
or U34245 (N_34245,N_33800,N_33875);
and U34246 (N_34246,N_33642,N_33932);
nor U34247 (N_34247,N_33545,N_33890);
or U34248 (N_34248,N_33805,N_33648);
nor U34249 (N_34249,N_33614,N_33608);
and U34250 (N_34250,N_33554,N_33879);
and U34251 (N_34251,N_33733,N_33727);
nand U34252 (N_34252,N_33838,N_33783);
and U34253 (N_34253,N_33765,N_33777);
and U34254 (N_34254,N_33577,N_33622);
nand U34255 (N_34255,N_33960,N_33774);
xnor U34256 (N_34256,N_33959,N_33799);
nand U34257 (N_34257,N_33968,N_33823);
nor U34258 (N_34258,N_33850,N_33563);
and U34259 (N_34259,N_33723,N_33562);
nand U34260 (N_34260,N_33658,N_33798);
nor U34261 (N_34261,N_33705,N_33730);
xnor U34262 (N_34262,N_33940,N_33686);
nor U34263 (N_34263,N_33871,N_33516);
nor U34264 (N_34264,N_33505,N_33645);
and U34265 (N_34265,N_33856,N_33926);
and U34266 (N_34266,N_33740,N_33530);
xnor U34267 (N_34267,N_33621,N_33951);
xnor U34268 (N_34268,N_33665,N_33842);
and U34269 (N_34269,N_33932,N_33608);
or U34270 (N_34270,N_33526,N_33865);
nor U34271 (N_34271,N_33837,N_33984);
and U34272 (N_34272,N_33567,N_33786);
or U34273 (N_34273,N_33689,N_33557);
or U34274 (N_34274,N_33817,N_33666);
nor U34275 (N_34275,N_33582,N_33865);
nor U34276 (N_34276,N_33738,N_33623);
xnor U34277 (N_34277,N_33615,N_33879);
and U34278 (N_34278,N_33580,N_33831);
and U34279 (N_34279,N_33537,N_33593);
or U34280 (N_34280,N_33612,N_33641);
and U34281 (N_34281,N_33792,N_33540);
or U34282 (N_34282,N_33745,N_33637);
nand U34283 (N_34283,N_33564,N_33671);
nand U34284 (N_34284,N_33586,N_33974);
xor U34285 (N_34285,N_33817,N_33903);
nor U34286 (N_34286,N_33940,N_33993);
or U34287 (N_34287,N_33858,N_33930);
nand U34288 (N_34288,N_33588,N_33971);
and U34289 (N_34289,N_33924,N_33521);
xor U34290 (N_34290,N_33851,N_33630);
or U34291 (N_34291,N_33688,N_33733);
xnor U34292 (N_34292,N_33919,N_33843);
and U34293 (N_34293,N_33610,N_33505);
or U34294 (N_34294,N_33857,N_33606);
nor U34295 (N_34295,N_33564,N_33589);
nor U34296 (N_34296,N_33969,N_33977);
and U34297 (N_34297,N_33646,N_33830);
nor U34298 (N_34298,N_33998,N_33713);
nand U34299 (N_34299,N_33510,N_33734);
xnor U34300 (N_34300,N_33730,N_33891);
nand U34301 (N_34301,N_33565,N_33502);
or U34302 (N_34302,N_33718,N_33806);
nor U34303 (N_34303,N_33558,N_33520);
nand U34304 (N_34304,N_33595,N_33936);
and U34305 (N_34305,N_33796,N_33975);
nand U34306 (N_34306,N_33961,N_33668);
nor U34307 (N_34307,N_33719,N_33681);
and U34308 (N_34308,N_33685,N_33660);
xor U34309 (N_34309,N_33647,N_33510);
nor U34310 (N_34310,N_33684,N_33670);
or U34311 (N_34311,N_33554,N_33870);
and U34312 (N_34312,N_33702,N_33955);
or U34313 (N_34313,N_33868,N_33926);
nor U34314 (N_34314,N_33810,N_33840);
nor U34315 (N_34315,N_33518,N_33873);
or U34316 (N_34316,N_33644,N_33643);
and U34317 (N_34317,N_33951,N_33732);
xnor U34318 (N_34318,N_33918,N_33767);
nor U34319 (N_34319,N_33525,N_33907);
or U34320 (N_34320,N_33613,N_33919);
and U34321 (N_34321,N_33609,N_33836);
or U34322 (N_34322,N_33829,N_33588);
or U34323 (N_34323,N_33871,N_33780);
or U34324 (N_34324,N_33606,N_33797);
nor U34325 (N_34325,N_33703,N_33691);
nor U34326 (N_34326,N_33714,N_33970);
nand U34327 (N_34327,N_33873,N_33667);
nor U34328 (N_34328,N_33752,N_33956);
nand U34329 (N_34329,N_33641,N_33836);
and U34330 (N_34330,N_33683,N_33903);
nand U34331 (N_34331,N_33539,N_33547);
xnor U34332 (N_34332,N_33703,N_33968);
xnor U34333 (N_34333,N_33639,N_33831);
or U34334 (N_34334,N_33679,N_33808);
nand U34335 (N_34335,N_33759,N_33669);
nand U34336 (N_34336,N_33844,N_33777);
xor U34337 (N_34337,N_33705,N_33623);
nor U34338 (N_34338,N_33706,N_33821);
nand U34339 (N_34339,N_33711,N_33757);
and U34340 (N_34340,N_33961,N_33626);
nor U34341 (N_34341,N_33933,N_33851);
nand U34342 (N_34342,N_33912,N_33717);
nor U34343 (N_34343,N_33815,N_33734);
or U34344 (N_34344,N_33929,N_33644);
nor U34345 (N_34345,N_33562,N_33857);
nor U34346 (N_34346,N_33724,N_33887);
xor U34347 (N_34347,N_33923,N_33687);
nand U34348 (N_34348,N_33842,N_33997);
or U34349 (N_34349,N_33640,N_33541);
nand U34350 (N_34350,N_33673,N_33946);
and U34351 (N_34351,N_33861,N_33583);
nand U34352 (N_34352,N_33619,N_33667);
or U34353 (N_34353,N_33922,N_33793);
nand U34354 (N_34354,N_33627,N_33885);
or U34355 (N_34355,N_33706,N_33961);
xnor U34356 (N_34356,N_33884,N_33632);
or U34357 (N_34357,N_33551,N_33892);
and U34358 (N_34358,N_33848,N_33960);
nand U34359 (N_34359,N_33756,N_33985);
or U34360 (N_34360,N_33993,N_33567);
xnor U34361 (N_34361,N_33572,N_33978);
nor U34362 (N_34362,N_33748,N_33901);
nor U34363 (N_34363,N_33552,N_33929);
nand U34364 (N_34364,N_33889,N_33635);
or U34365 (N_34365,N_33506,N_33732);
nand U34366 (N_34366,N_33609,N_33841);
nand U34367 (N_34367,N_33975,N_33962);
and U34368 (N_34368,N_33878,N_33577);
nand U34369 (N_34369,N_33786,N_33823);
xnor U34370 (N_34370,N_33825,N_33587);
xnor U34371 (N_34371,N_33557,N_33839);
xnor U34372 (N_34372,N_33855,N_33639);
nand U34373 (N_34373,N_33813,N_33599);
xor U34374 (N_34374,N_33861,N_33714);
or U34375 (N_34375,N_33650,N_33793);
nand U34376 (N_34376,N_33738,N_33813);
nand U34377 (N_34377,N_33878,N_33933);
and U34378 (N_34378,N_33975,N_33948);
and U34379 (N_34379,N_33765,N_33965);
xnor U34380 (N_34380,N_33801,N_33735);
and U34381 (N_34381,N_33710,N_33825);
nor U34382 (N_34382,N_33935,N_33768);
nand U34383 (N_34383,N_33720,N_33512);
nand U34384 (N_34384,N_33921,N_33674);
or U34385 (N_34385,N_33516,N_33577);
nand U34386 (N_34386,N_33960,N_33680);
nand U34387 (N_34387,N_33684,N_33766);
xor U34388 (N_34388,N_33507,N_33824);
and U34389 (N_34389,N_33891,N_33731);
nand U34390 (N_34390,N_33827,N_33600);
nor U34391 (N_34391,N_33624,N_33886);
and U34392 (N_34392,N_33802,N_33645);
or U34393 (N_34393,N_33866,N_33751);
nor U34394 (N_34394,N_33692,N_33633);
nand U34395 (N_34395,N_33760,N_33848);
or U34396 (N_34396,N_33746,N_33897);
xnor U34397 (N_34397,N_33650,N_33571);
nor U34398 (N_34398,N_33673,N_33936);
or U34399 (N_34399,N_33850,N_33796);
nor U34400 (N_34400,N_33726,N_33531);
or U34401 (N_34401,N_33602,N_33575);
xor U34402 (N_34402,N_33696,N_33645);
xor U34403 (N_34403,N_33896,N_33872);
and U34404 (N_34404,N_33767,N_33732);
nand U34405 (N_34405,N_33967,N_33926);
or U34406 (N_34406,N_33687,N_33641);
and U34407 (N_34407,N_33990,N_33738);
nand U34408 (N_34408,N_33597,N_33694);
nor U34409 (N_34409,N_33552,N_33902);
xnor U34410 (N_34410,N_33602,N_33979);
xor U34411 (N_34411,N_33672,N_33502);
xnor U34412 (N_34412,N_33583,N_33774);
nor U34413 (N_34413,N_33918,N_33945);
xnor U34414 (N_34414,N_33677,N_33513);
nor U34415 (N_34415,N_33960,N_33642);
nand U34416 (N_34416,N_33814,N_33944);
nor U34417 (N_34417,N_33967,N_33599);
xnor U34418 (N_34418,N_33932,N_33839);
nand U34419 (N_34419,N_33934,N_33921);
nand U34420 (N_34420,N_33539,N_33968);
nor U34421 (N_34421,N_33553,N_33738);
nand U34422 (N_34422,N_33685,N_33719);
nand U34423 (N_34423,N_33738,N_33537);
nand U34424 (N_34424,N_33539,N_33572);
xor U34425 (N_34425,N_33627,N_33500);
and U34426 (N_34426,N_33666,N_33777);
nand U34427 (N_34427,N_33584,N_33578);
and U34428 (N_34428,N_33951,N_33762);
nand U34429 (N_34429,N_33710,N_33959);
nor U34430 (N_34430,N_33585,N_33985);
nor U34431 (N_34431,N_33531,N_33688);
or U34432 (N_34432,N_33971,N_33791);
nor U34433 (N_34433,N_33888,N_33965);
and U34434 (N_34434,N_33984,N_33796);
nor U34435 (N_34435,N_33681,N_33705);
or U34436 (N_34436,N_33772,N_33840);
nand U34437 (N_34437,N_33927,N_33589);
nand U34438 (N_34438,N_33662,N_33555);
or U34439 (N_34439,N_33957,N_33722);
nor U34440 (N_34440,N_33671,N_33740);
xor U34441 (N_34441,N_33831,N_33573);
or U34442 (N_34442,N_33797,N_33876);
xnor U34443 (N_34443,N_33804,N_33582);
nand U34444 (N_34444,N_33940,N_33887);
or U34445 (N_34445,N_33921,N_33773);
and U34446 (N_34446,N_33743,N_33732);
and U34447 (N_34447,N_33527,N_33517);
or U34448 (N_34448,N_33514,N_33829);
nor U34449 (N_34449,N_33735,N_33725);
xnor U34450 (N_34450,N_33956,N_33639);
nand U34451 (N_34451,N_33696,N_33518);
nor U34452 (N_34452,N_33816,N_33915);
xnor U34453 (N_34453,N_33715,N_33876);
or U34454 (N_34454,N_33765,N_33830);
nor U34455 (N_34455,N_33661,N_33539);
or U34456 (N_34456,N_33681,N_33992);
or U34457 (N_34457,N_33554,N_33665);
or U34458 (N_34458,N_33522,N_33706);
xnor U34459 (N_34459,N_33757,N_33510);
nand U34460 (N_34460,N_33837,N_33935);
or U34461 (N_34461,N_33735,N_33767);
nor U34462 (N_34462,N_33544,N_33667);
or U34463 (N_34463,N_33673,N_33587);
xor U34464 (N_34464,N_33885,N_33743);
nor U34465 (N_34465,N_33501,N_33986);
nor U34466 (N_34466,N_33907,N_33939);
and U34467 (N_34467,N_33777,N_33672);
nor U34468 (N_34468,N_33838,N_33534);
xnor U34469 (N_34469,N_33677,N_33543);
or U34470 (N_34470,N_33863,N_33547);
or U34471 (N_34471,N_33579,N_33715);
or U34472 (N_34472,N_33820,N_33512);
xor U34473 (N_34473,N_33894,N_33729);
nor U34474 (N_34474,N_33501,N_33605);
or U34475 (N_34475,N_33600,N_33714);
and U34476 (N_34476,N_33818,N_33550);
and U34477 (N_34477,N_33607,N_33873);
and U34478 (N_34478,N_33835,N_33708);
xnor U34479 (N_34479,N_33810,N_33835);
nand U34480 (N_34480,N_33721,N_33554);
xor U34481 (N_34481,N_33582,N_33752);
xor U34482 (N_34482,N_33907,N_33880);
and U34483 (N_34483,N_33706,N_33959);
nor U34484 (N_34484,N_33799,N_33501);
nor U34485 (N_34485,N_33823,N_33569);
nor U34486 (N_34486,N_33711,N_33870);
nand U34487 (N_34487,N_33641,N_33615);
and U34488 (N_34488,N_33852,N_33727);
nand U34489 (N_34489,N_33525,N_33716);
xnor U34490 (N_34490,N_33632,N_33613);
and U34491 (N_34491,N_33628,N_33793);
nor U34492 (N_34492,N_33538,N_33626);
xor U34493 (N_34493,N_33593,N_33745);
xnor U34494 (N_34494,N_33895,N_33773);
or U34495 (N_34495,N_33815,N_33616);
xnor U34496 (N_34496,N_33690,N_33618);
or U34497 (N_34497,N_33502,N_33683);
nor U34498 (N_34498,N_33844,N_33917);
or U34499 (N_34499,N_33874,N_33868);
or U34500 (N_34500,N_34035,N_34123);
xor U34501 (N_34501,N_34292,N_34331);
nor U34502 (N_34502,N_34218,N_34055);
nor U34503 (N_34503,N_34401,N_34230);
or U34504 (N_34504,N_34485,N_34117);
nor U34505 (N_34505,N_34071,N_34447);
nand U34506 (N_34506,N_34153,N_34466);
nor U34507 (N_34507,N_34087,N_34224);
nor U34508 (N_34508,N_34255,N_34263);
nor U34509 (N_34509,N_34484,N_34237);
nand U34510 (N_34510,N_34465,N_34273);
xor U34511 (N_34511,N_34046,N_34079);
nand U34512 (N_34512,N_34043,N_34160);
nor U34513 (N_34513,N_34450,N_34262);
or U34514 (N_34514,N_34487,N_34395);
nor U34515 (N_34515,N_34392,N_34282);
nand U34516 (N_34516,N_34471,N_34173);
nand U34517 (N_34517,N_34125,N_34396);
nor U34518 (N_34518,N_34380,N_34095);
or U34519 (N_34519,N_34072,N_34184);
and U34520 (N_34520,N_34427,N_34330);
and U34521 (N_34521,N_34214,N_34412);
and U34522 (N_34522,N_34496,N_34404);
or U34523 (N_34523,N_34171,N_34200);
xnor U34524 (N_34524,N_34267,N_34403);
or U34525 (N_34525,N_34062,N_34113);
nor U34526 (N_34526,N_34144,N_34418);
xnor U34527 (N_34527,N_34190,N_34299);
nor U34528 (N_34528,N_34383,N_34446);
nand U34529 (N_34529,N_34333,N_34287);
nand U34530 (N_34530,N_34008,N_34378);
xnor U34531 (N_34531,N_34139,N_34470);
nor U34532 (N_34532,N_34250,N_34460);
nand U34533 (N_34533,N_34099,N_34235);
nand U34534 (N_34534,N_34059,N_34488);
nor U34535 (N_34535,N_34397,N_34207);
xor U34536 (N_34536,N_34416,N_34133);
xnor U34537 (N_34537,N_34238,N_34081);
or U34538 (N_34538,N_34111,N_34351);
nand U34539 (N_34539,N_34122,N_34024);
nand U34540 (N_34540,N_34166,N_34402);
nand U34541 (N_34541,N_34345,N_34121);
or U34542 (N_34542,N_34258,N_34246);
and U34543 (N_34543,N_34359,N_34411);
xor U34544 (N_34544,N_34228,N_34256);
and U34545 (N_34545,N_34169,N_34322);
nand U34546 (N_34546,N_34315,N_34325);
nand U34547 (N_34547,N_34353,N_34432);
nand U34548 (N_34548,N_34134,N_34327);
or U34549 (N_34549,N_34157,N_34464);
nand U34550 (N_34550,N_34083,N_34451);
or U34551 (N_34551,N_34461,N_34372);
or U34552 (N_34552,N_34023,N_34311);
and U34553 (N_34553,N_34280,N_34149);
and U34554 (N_34554,N_34114,N_34268);
or U34555 (N_34555,N_34360,N_34198);
nor U34556 (N_34556,N_34456,N_34305);
or U34557 (N_34557,N_34017,N_34349);
nand U34558 (N_34558,N_34105,N_34068);
nor U34559 (N_34559,N_34319,N_34410);
or U34560 (N_34560,N_34009,N_34208);
xnor U34561 (N_34561,N_34340,N_34152);
nor U34562 (N_34562,N_34381,N_34039);
or U34563 (N_34563,N_34475,N_34300);
or U34564 (N_34564,N_34251,N_34119);
or U34565 (N_34565,N_34002,N_34006);
or U34566 (N_34566,N_34248,N_34356);
nand U34567 (N_34567,N_34400,N_34457);
nor U34568 (N_34568,N_34147,N_34220);
xnor U34569 (N_34569,N_34435,N_34141);
xnor U34570 (N_34570,N_34474,N_34350);
nand U34571 (N_34571,N_34309,N_34495);
or U34572 (N_34572,N_34061,N_34329);
xor U34573 (N_34573,N_34472,N_34398);
nor U34574 (N_34574,N_34366,N_34388);
nor U34575 (N_34575,N_34056,N_34005);
nand U34576 (N_34576,N_34037,N_34490);
or U34577 (N_34577,N_34227,N_34084);
and U34578 (N_34578,N_34212,N_34272);
nor U34579 (N_34579,N_34162,N_34003);
nand U34580 (N_34580,N_34449,N_34343);
xnor U34581 (N_34581,N_34029,N_34074);
or U34582 (N_34582,N_34129,N_34321);
nor U34583 (N_34583,N_34478,N_34086);
nor U34584 (N_34584,N_34463,N_34399);
xor U34585 (N_34585,N_34443,N_34430);
and U34586 (N_34586,N_34177,N_34124);
nor U34587 (N_34587,N_34453,N_34483);
and U34588 (N_34588,N_34452,N_34182);
xor U34589 (N_34589,N_34000,N_34091);
nor U34590 (N_34590,N_34110,N_34140);
or U34591 (N_34591,N_34192,N_34339);
and U34592 (N_34592,N_34025,N_34323);
xnor U34593 (N_34593,N_34243,N_34232);
or U34594 (N_34594,N_34441,N_34486);
or U34595 (N_34595,N_34259,N_34172);
nand U34596 (N_34596,N_34201,N_34298);
nand U34597 (N_34597,N_34328,N_34165);
nand U34598 (N_34598,N_34245,N_34194);
nor U34599 (N_34599,N_34438,N_34363);
or U34600 (N_34600,N_34247,N_34209);
or U34601 (N_34601,N_34436,N_34310);
xnor U34602 (N_34602,N_34468,N_34219);
or U34603 (N_34603,N_34415,N_34320);
nor U34604 (N_34604,N_34163,N_34313);
or U34605 (N_34605,N_34308,N_34082);
nand U34606 (N_34606,N_34269,N_34052);
nand U34607 (N_34607,N_34021,N_34264);
or U34608 (N_34608,N_34492,N_34130);
nor U34609 (N_34609,N_34189,N_34389);
and U34610 (N_34610,N_34088,N_34317);
nand U34611 (N_34611,N_34040,N_34181);
or U34612 (N_34612,N_34249,N_34213);
or U34613 (N_34613,N_34342,N_34090);
nor U34614 (N_34614,N_34065,N_34234);
nand U34615 (N_34615,N_34151,N_34284);
or U34616 (N_34616,N_34275,N_34473);
and U34617 (N_34617,N_34354,N_34004);
or U34618 (N_34618,N_34096,N_34112);
and U34619 (N_34619,N_34188,N_34116);
xnor U34620 (N_34620,N_34390,N_34285);
and U34621 (N_34621,N_34047,N_34393);
and U34622 (N_34622,N_34196,N_34186);
nand U34623 (N_34623,N_34027,N_34304);
and U34624 (N_34624,N_34306,N_34458);
or U34625 (N_34625,N_34482,N_34455);
and U34626 (N_34626,N_34085,N_34377);
nand U34627 (N_34627,N_34075,N_34289);
nand U34628 (N_34628,N_34375,N_34089);
or U34629 (N_34629,N_34373,N_34332);
nand U34630 (N_34630,N_34143,N_34481);
nand U34631 (N_34631,N_34498,N_34344);
or U34632 (N_34632,N_34296,N_34467);
nand U34633 (N_34633,N_34421,N_34108);
nor U34634 (N_34634,N_34261,N_34109);
and U34635 (N_34635,N_34358,N_34476);
nor U34636 (N_34636,N_34431,N_34058);
nor U34637 (N_34637,N_34131,N_34494);
xnor U34638 (N_34638,N_34033,N_34026);
or U34639 (N_34639,N_34491,N_34374);
and U34640 (N_34640,N_34078,N_34369);
nand U34641 (N_34641,N_34428,N_34176);
nor U34642 (N_34642,N_34288,N_34417);
xnor U34643 (N_34643,N_34080,N_34132);
and U34644 (N_34644,N_34335,N_34077);
and U34645 (N_34645,N_34422,N_34437);
xor U34646 (N_34646,N_34120,N_34225);
nor U34647 (N_34647,N_34093,N_34053);
and U34648 (N_34648,N_34352,N_34100);
nor U34649 (N_34649,N_34146,N_34312);
or U34650 (N_34650,N_34307,N_34054);
xor U34651 (N_34651,N_34303,N_34019);
nand U34652 (N_34652,N_34101,N_34076);
nand U34653 (N_34653,N_34098,N_34191);
xor U34654 (N_34654,N_34297,N_34367);
or U34655 (N_34655,N_34391,N_34217);
xor U34656 (N_34656,N_34407,N_34286);
nand U34657 (N_34657,N_34066,N_34038);
and U34658 (N_34658,N_34185,N_34069);
or U34659 (N_34659,N_34326,N_34257);
nor U34660 (N_34660,N_34142,N_34097);
or U34661 (N_34661,N_34167,N_34223);
nor U34662 (N_34662,N_34362,N_34007);
xor U34663 (N_34663,N_34278,N_34150);
nor U34664 (N_34664,N_34324,N_34197);
xnor U34665 (N_34665,N_34244,N_34252);
and U34666 (N_34666,N_34161,N_34229);
and U34667 (N_34667,N_34063,N_34290);
and U34668 (N_34668,N_34341,N_34445);
or U34669 (N_34669,N_34064,N_34092);
and U34670 (N_34670,N_34001,N_34126);
and U34671 (N_34671,N_34148,N_34236);
and U34672 (N_34672,N_34420,N_34294);
nand U34673 (N_34673,N_34239,N_34060);
and U34674 (N_34674,N_34204,N_34115);
xor U34675 (N_34675,N_34454,N_34222);
xor U34676 (N_34676,N_34419,N_34336);
and U34677 (N_34677,N_34202,N_34364);
nand U34678 (N_34678,N_34205,N_34357);
and U34679 (N_34679,N_34011,N_34382);
xor U34680 (N_34680,N_34102,N_34216);
or U34681 (N_34681,N_34107,N_34044);
nand U34682 (N_34682,N_34276,N_34241);
nand U34683 (N_34683,N_34018,N_34016);
and U34684 (N_34684,N_34265,N_34106);
xnor U34685 (N_34685,N_34070,N_34210);
xor U34686 (N_34686,N_34370,N_34379);
or U34687 (N_34687,N_34424,N_34045);
nand U34688 (N_34688,N_34409,N_34423);
or U34689 (N_34689,N_34159,N_34015);
nor U34690 (N_34690,N_34477,N_34187);
nand U34691 (N_34691,N_34179,N_34057);
or U34692 (N_34692,N_34281,N_34155);
nand U34693 (N_34693,N_34014,N_34406);
nor U34694 (N_34694,N_34041,N_34413);
and U34695 (N_34695,N_34469,N_34429);
xnor U34696 (N_34696,N_34387,N_34012);
nand U34697 (N_34697,N_34384,N_34073);
nand U34698 (N_34698,N_34355,N_34137);
and U34699 (N_34699,N_34371,N_34094);
nand U34700 (N_34700,N_34361,N_34158);
xor U34701 (N_34701,N_34376,N_34254);
or U34702 (N_34702,N_34348,N_34104);
nand U34703 (N_34703,N_34433,N_34013);
or U34704 (N_34704,N_34180,N_34283);
nand U34705 (N_34705,N_34240,N_34439);
nor U34706 (N_34706,N_34291,N_34170);
or U34707 (N_34707,N_34405,N_34260);
nand U34708 (N_34708,N_34028,N_34316);
or U34709 (N_34709,N_34030,N_34215);
xnor U34710 (N_34710,N_34231,N_34489);
or U34711 (N_34711,N_34274,N_34242);
or U34712 (N_34712,N_34293,N_34385);
nor U34713 (N_34713,N_34497,N_34199);
xnor U34714 (N_34714,N_34270,N_34118);
nor U34715 (N_34715,N_34206,N_34459);
or U34716 (N_34716,N_34386,N_34164);
nand U34717 (N_34717,N_34042,N_34499);
nand U34718 (N_34718,N_34020,N_34347);
xnor U34719 (N_34719,N_34338,N_34434);
nor U34720 (N_34720,N_34211,N_34048);
or U34721 (N_34721,N_34195,N_34156);
xor U34722 (N_34722,N_34136,N_34138);
and U34723 (N_34723,N_34425,N_34334);
nor U34724 (N_34724,N_34031,N_34168);
and U34725 (N_34725,N_34032,N_34444);
and U34726 (N_34726,N_34414,N_34034);
nand U34727 (N_34727,N_34036,N_34426);
xor U34728 (N_34728,N_34301,N_34337);
xnor U34729 (N_34729,N_34295,N_34050);
and U34730 (N_34730,N_34314,N_34493);
nor U34731 (N_34731,N_34178,N_34408);
nor U34732 (N_34732,N_34440,N_34051);
or U34733 (N_34733,N_34479,N_34226);
and U34734 (N_34734,N_34221,N_34175);
xor U34735 (N_34735,N_34154,N_34480);
or U34736 (N_34736,N_34022,N_34233);
nor U34737 (N_34737,N_34203,N_34442);
and U34738 (N_34738,N_34253,N_34103);
or U34739 (N_34739,N_34049,N_34302);
nor U34740 (N_34740,N_34135,N_34145);
nand U34741 (N_34741,N_34346,N_34448);
and U34742 (N_34742,N_34174,N_34368);
and U34743 (N_34743,N_34271,N_34318);
nand U34744 (N_34744,N_34128,N_34277);
nor U34745 (N_34745,N_34127,N_34183);
or U34746 (N_34746,N_34365,N_34010);
nor U34747 (N_34747,N_34279,N_34067);
or U34748 (N_34748,N_34462,N_34266);
and U34749 (N_34749,N_34394,N_34193);
and U34750 (N_34750,N_34003,N_34111);
or U34751 (N_34751,N_34102,N_34435);
or U34752 (N_34752,N_34495,N_34453);
xor U34753 (N_34753,N_34027,N_34408);
xor U34754 (N_34754,N_34224,N_34359);
xor U34755 (N_34755,N_34432,N_34490);
nand U34756 (N_34756,N_34414,N_34190);
nand U34757 (N_34757,N_34076,N_34350);
nand U34758 (N_34758,N_34017,N_34431);
and U34759 (N_34759,N_34355,N_34008);
nand U34760 (N_34760,N_34198,N_34278);
xnor U34761 (N_34761,N_34313,N_34035);
xnor U34762 (N_34762,N_34365,N_34055);
and U34763 (N_34763,N_34344,N_34384);
or U34764 (N_34764,N_34357,N_34424);
xor U34765 (N_34765,N_34216,N_34343);
and U34766 (N_34766,N_34167,N_34453);
nand U34767 (N_34767,N_34114,N_34214);
or U34768 (N_34768,N_34477,N_34161);
xnor U34769 (N_34769,N_34387,N_34441);
nand U34770 (N_34770,N_34090,N_34467);
nor U34771 (N_34771,N_34039,N_34105);
or U34772 (N_34772,N_34409,N_34107);
nor U34773 (N_34773,N_34328,N_34038);
nor U34774 (N_34774,N_34142,N_34433);
or U34775 (N_34775,N_34059,N_34347);
nand U34776 (N_34776,N_34480,N_34149);
or U34777 (N_34777,N_34213,N_34229);
xnor U34778 (N_34778,N_34001,N_34495);
or U34779 (N_34779,N_34216,N_34001);
nor U34780 (N_34780,N_34174,N_34425);
xor U34781 (N_34781,N_34004,N_34455);
nand U34782 (N_34782,N_34181,N_34282);
nor U34783 (N_34783,N_34109,N_34259);
and U34784 (N_34784,N_34102,N_34423);
nor U34785 (N_34785,N_34238,N_34023);
nor U34786 (N_34786,N_34297,N_34298);
xnor U34787 (N_34787,N_34122,N_34365);
or U34788 (N_34788,N_34122,N_34447);
nand U34789 (N_34789,N_34034,N_34381);
nand U34790 (N_34790,N_34373,N_34497);
or U34791 (N_34791,N_34439,N_34374);
and U34792 (N_34792,N_34000,N_34119);
nor U34793 (N_34793,N_34428,N_34036);
xor U34794 (N_34794,N_34161,N_34492);
xnor U34795 (N_34795,N_34420,N_34231);
nor U34796 (N_34796,N_34079,N_34315);
xor U34797 (N_34797,N_34119,N_34088);
nor U34798 (N_34798,N_34284,N_34132);
xor U34799 (N_34799,N_34168,N_34101);
and U34800 (N_34800,N_34132,N_34212);
or U34801 (N_34801,N_34368,N_34232);
nor U34802 (N_34802,N_34102,N_34326);
and U34803 (N_34803,N_34433,N_34363);
or U34804 (N_34804,N_34078,N_34102);
and U34805 (N_34805,N_34374,N_34100);
and U34806 (N_34806,N_34493,N_34020);
xnor U34807 (N_34807,N_34161,N_34213);
nor U34808 (N_34808,N_34460,N_34313);
and U34809 (N_34809,N_34392,N_34424);
xor U34810 (N_34810,N_34395,N_34294);
nand U34811 (N_34811,N_34274,N_34281);
nand U34812 (N_34812,N_34212,N_34267);
xor U34813 (N_34813,N_34202,N_34042);
or U34814 (N_34814,N_34334,N_34187);
or U34815 (N_34815,N_34450,N_34111);
nand U34816 (N_34816,N_34390,N_34082);
nor U34817 (N_34817,N_34081,N_34358);
and U34818 (N_34818,N_34099,N_34180);
or U34819 (N_34819,N_34042,N_34391);
nor U34820 (N_34820,N_34238,N_34163);
nor U34821 (N_34821,N_34110,N_34366);
nand U34822 (N_34822,N_34388,N_34141);
nor U34823 (N_34823,N_34009,N_34426);
nor U34824 (N_34824,N_34127,N_34336);
xor U34825 (N_34825,N_34303,N_34393);
nor U34826 (N_34826,N_34107,N_34230);
or U34827 (N_34827,N_34129,N_34447);
nand U34828 (N_34828,N_34416,N_34056);
or U34829 (N_34829,N_34447,N_34294);
nand U34830 (N_34830,N_34119,N_34393);
nor U34831 (N_34831,N_34027,N_34294);
and U34832 (N_34832,N_34137,N_34354);
xor U34833 (N_34833,N_34248,N_34082);
xnor U34834 (N_34834,N_34197,N_34496);
or U34835 (N_34835,N_34024,N_34097);
and U34836 (N_34836,N_34041,N_34175);
nor U34837 (N_34837,N_34493,N_34355);
nor U34838 (N_34838,N_34104,N_34000);
nor U34839 (N_34839,N_34159,N_34465);
or U34840 (N_34840,N_34235,N_34349);
xnor U34841 (N_34841,N_34294,N_34290);
nor U34842 (N_34842,N_34201,N_34053);
nor U34843 (N_34843,N_34218,N_34265);
or U34844 (N_34844,N_34283,N_34486);
and U34845 (N_34845,N_34432,N_34264);
nand U34846 (N_34846,N_34301,N_34332);
xor U34847 (N_34847,N_34110,N_34156);
nor U34848 (N_34848,N_34184,N_34364);
or U34849 (N_34849,N_34021,N_34051);
and U34850 (N_34850,N_34076,N_34306);
or U34851 (N_34851,N_34141,N_34465);
or U34852 (N_34852,N_34312,N_34168);
nand U34853 (N_34853,N_34284,N_34190);
and U34854 (N_34854,N_34059,N_34410);
and U34855 (N_34855,N_34187,N_34243);
or U34856 (N_34856,N_34389,N_34099);
and U34857 (N_34857,N_34337,N_34259);
and U34858 (N_34858,N_34383,N_34166);
nor U34859 (N_34859,N_34276,N_34289);
and U34860 (N_34860,N_34366,N_34416);
xor U34861 (N_34861,N_34389,N_34091);
xor U34862 (N_34862,N_34023,N_34012);
xnor U34863 (N_34863,N_34473,N_34261);
nand U34864 (N_34864,N_34264,N_34373);
and U34865 (N_34865,N_34360,N_34105);
nor U34866 (N_34866,N_34148,N_34019);
nor U34867 (N_34867,N_34494,N_34068);
nand U34868 (N_34868,N_34196,N_34135);
or U34869 (N_34869,N_34452,N_34255);
and U34870 (N_34870,N_34262,N_34402);
nor U34871 (N_34871,N_34064,N_34160);
xnor U34872 (N_34872,N_34119,N_34114);
xor U34873 (N_34873,N_34439,N_34157);
nand U34874 (N_34874,N_34057,N_34293);
nor U34875 (N_34875,N_34186,N_34341);
xor U34876 (N_34876,N_34267,N_34448);
or U34877 (N_34877,N_34260,N_34468);
nand U34878 (N_34878,N_34477,N_34213);
xnor U34879 (N_34879,N_34226,N_34495);
xnor U34880 (N_34880,N_34326,N_34096);
nand U34881 (N_34881,N_34236,N_34037);
nand U34882 (N_34882,N_34214,N_34246);
nand U34883 (N_34883,N_34186,N_34393);
xnor U34884 (N_34884,N_34112,N_34034);
xor U34885 (N_34885,N_34251,N_34415);
nor U34886 (N_34886,N_34297,N_34410);
or U34887 (N_34887,N_34492,N_34410);
and U34888 (N_34888,N_34480,N_34062);
nand U34889 (N_34889,N_34020,N_34044);
and U34890 (N_34890,N_34336,N_34334);
or U34891 (N_34891,N_34175,N_34268);
nor U34892 (N_34892,N_34373,N_34406);
or U34893 (N_34893,N_34449,N_34000);
nor U34894 (N_34894,N_34282,N_34407);
and U34895 (N_34895,N_34211,N_34346);
and U34896 (N_34896,N_34053,N_34153);
or U34897 (N_34897,N_34428,N_34235);
or U34898 (N_34898,N_34136,N_34282);
nor U34899 (N_34899,N_34126,N_34066);
xor U34900 (N_34900,N_34279,N_34325);
nand U34901 (N_34901,N_34499,N_34066);
nand U34902 (N_34902,N_34213,N_34185);
and U34903 (N_34903,N_34368,N_34273);
xnor U34904 (N_34904,N_34136,N_34007);
xor U34905 (N_34905,N_34056,N_34403);
nor U34906 (N_34906,N_34274,N_34110);
nor U34907 (N_34907,N_34068,N_34030);
xor U34908 (N_34908,N_34047,N_34193);
xor U34909 (N_34909,N_34267,N_34278);
nand U34910 (N_34910,N_34141,N_34361);
or U34911 (N_34911,N_34144,N_34342);
xor U34912 (N_34912,N_34170,N_34387);
or U34913 (N_34913,N_34369,N_34210);
nand U34914 (N_34914,N_34427,N_34300);
and U34915 (N_34915,N_34434,N_34033);
nor U34916 (N_34916,N_34289,N_34390);
xor U34917 (N_34917,N_34256,N_34040);
nor U34918 (N_34918,N_34066,N_34441);
xor U34919 (N_34919,N_34492,N_34244);
or U34920 (N_34920,N_34278,N_34013);
nand U34921 (N_34921,N_34163,N_34368);
and U34922 (N_34922,N_34386,N_34103);
nand U34923 (N_34923,N_34105,N_34448);
nand U34924 (N_34924,N_34264,N_34314);
nor U34925 (N_34925,N_34113,N_34216);
nand U34926 (N_34926,N_34369,N_34070);
nor U34927 (N_34927,N_34355,N_34174);
xnor U34928 (N_34928,N_34427,N_34011);
nor U34929 (N_34929,N_34277,N_34036);
xor U34930 (N_34930,N_34492,N_34432);
or U34931 (N_34931,N_34250,N_34414);
and U34932 (N_34932,N_34297,N_34369);
nor U34933 (N_34933,N_34046,N_34492);
or U34934 (N_34934,N_34425,N_34368);
nand U34935 (N_34935,N_34275,N_34351);
xnor U34936 (N_34936,N_34087,N_34356);
or U34937 (N_34937,N_34356,N_34088);
nand U34938 (N_34938,N_34071,N_34146);
or U34939 (N_34939,N_34007,N_34471);
nor U34940 (N_34940,N_34382,N_34368);
or U34941 (N_34941,N_34349,N_34019);
xor U34942 (N_34942,N_34032,N_34030);
and U34943 (N_34943,N_34150,N_34258);
nor U34944 (N_34944,N_34202,N_34326);
or U34945 (N_34945,N_34370,N_34189);
nor U34946 (N_34946,N_34296,N_34478);
nor U34947 (N_34947,N_34130,N_34419);
nor U34948 (N_34948,N_34411,N_34050);
nor U34949 (N_34949,N_34287,N_34350);
nand U34950 (N_34950,N_34079,N_34231);
xnor U34951 (N_34951,N_34359,N_34384);
xor U34952 (N_34952,N_34271,N_34051);
nor U34953 (N_34953,N_34185,N_34361);
or U34954 (N_34954,N_34327,N_34363);
xor U34955 (N_34955,N_34245,N_34140);
or U34956 (N_34956,N_34366,N_34303);
nor U34957 (N_34957,N_34134,N_34038);
nand U34958 (N_34958,N_34114,N_34053);
nand U34959 (N_34959,N_34124,N_34224);
or U34960 (N_34960,N_34443,N_34386);
nand U34961 (N_34961,N_34181,N_34073);
and U34962 (N_34962,N_34089,N_34270);
nand U34963 (N_34963,N_34154,N_34178);
or U34964 (N_34964,N_34166,N_34485);
nand U34965 (N_34965,N_34313,N_34042);
nor U34966 (N_34966,N_34364,N_34326);
or U34967 (N_34967,N_34332,N_34034);
or U34968 (N_34968,N_34183,N_34061);
nand U34969 (N_34969,N_34068,N_34312);
and U34970 (N_34970,N_34047,N_34324);
nand U34971 (N_34971,N_34376,N_34469);
nor U34972 (N_34972,N_34162,N_34282);
nand U34973 (N_34973,N_34264,N_34254);
nor U34974 (N_34974,N_34033,N_34042);
or U34975 (N_34975,N_34378,N_34486);
and U34976 (N_34976,N_34447,N_34349);
nor U34977 (N_34977,N_34420,N_34151);
nand U34978 (N_34978,N_34496,N_34182);
or U34979 (N_34979,N_34142,N_34324);
nand U34980 (N_34980,N_34418,N_34051);
nor U34981 (N_34981,N_34428,N_34373);
nor U34982 (N_34982,N_34354,N_34279);
nor U34983 (N_34983,N_34183,N_34217);
nor U34984 (N_34984,N_34396,N_34218);
xor U34985 (N_34985,N_34450,N_34285);
or U34986 (N_34986,N_34035,N_34307);
or U34987 (N_34987,N_34020,N_34312);
and U34988 (N_34988,N_34212,N_34372);
nor U34989 (N_34989,N_34394,N_34176);
nor U34990 (N_34990,N_34270,N_34104);
nand U34991 (N_34991,N_34175,N_34083);
nor U34992 (N_34992,N_34069,N_34456);
nand U34993 (N_34993,N_34246,N_34077);
xor U34994 (N_34994,N_34061,N_34132);
or U34995 (N_34995,N_34061,N_34346);
xnor U34996 (N_34996,N_34498,N_34104);
xor U34997 (N_34997,N_34082,N_34362);
and U34998 (N_34998,N_34423,N_34295);
nor U34999 (N_34999,N_34203,N_34120);
and U35000 (N_35000,N_34660,N_34609);
xnor U35001 (N_35001,N_34669,N_34711);
nand U35002 (N_35002,N_34570,N_34507);
nor U35003 (N_35003,N_34792,N_34807);
or U35004 (N_35004,N_34813,N_34758);
nor U35005 (N_35005,N_34786,N_34699);
xor U35006 (N_35006,N_34635,N_34793);
xnor U35007 (N_35007,N_34958,N_34674);
or U35008 (N_35008,N_34659,N_34845);
xor U35009 (N_35009,N_34504,N_34578);
xor U35010 (N_35010,N_34521,N_34545);
and U35011 (N_35011,N_34831,N_34735);
nor U35012 (N_35012,N_34751,N_34827);
xnor U35013 (N_35013,N_34910,N_34867);
xor U35014 (N_35014,N_34940,N_34528);
and U35015 (N_35015,N_34936,N_34708);
nor U35016 (N_35016,N_34869,N_34858);
or U35017 (N_35017,N_34822,N_34789);
or U35018 (N_35018,N_34951,N_34955);
nor U35019 (N_35019,N_34879,N_34995);
and U35020 (N_35020,N_34830,N_34608);
xnor U35021 (N_35021,N_34833,N_34851);
xnor U35022 (N_35022,N_34641,N_34969);
and U35023 (N_35023,N_34954,N_34871);
or U35024 (N_35024,N_34706,N_34580);
nor U35025 (N_35025,N_34853,N_34559);
nor U35026 (N_35026,N_34664,N_34791);
nor U35027 (N_35027,N_34882,N_34992);
and U35028 (N_35028,N_34614,N_34774);
nor U35029 (N_35029,N_34937,N_34957);
nand U35030 (N_35030,N_34982,N_34811);
or U35031 (N_35031,N_34935,N_34551);
or U35032 (N_35032,N_34956,N_34908);
and U35033 (N_35033,N_34546,N_34556);
xor U35034 (N_35034,N_34779,N_34803);
nor U35035 (N_35035,N_34874,N_34634);
xor U35036 (N_35036,N_34595,N_34610);
nor U35037 (N_35037,N_34650,N_34941);
nor U35038 (N_35038,N_34772,N_34938);
and U35039 (N_35039,N_34619,N_34698);
and U35040 (N_35040,N_34922,N_34932);
and U35041 (N_35041,N_34880,N_34892);
and U35042 (N_35042,N_34796,N_34859);
or U35043 (N_35043,N_34978,N_34657);
or U35044 (N_35044,N_34946,N_34763);
nand U35045 (N_35045,N_34638,N_34847);
nor U35046 (N_35046,N_34555,N_34678);
nand U35047 (N_35047,N_34615,N_34891);
xnor U35048 (N_35048,N_34719,N_34677);
nand U35049 (N_35049,N_34740,N_34966);
or U35050 (N_35050,N_34945,N_34596);
nand U35051 (N_35051,N_34761,N_34987);
nor U35052 (N_35052,N_34921,N_34737);
and U35053 (N_35053,N_34848,N_34990);
and U35054 (N_35054,N_34630,N_34773);
nand U35055 (N_35055,N_34997,N_34994);
and U35056 (N_35056,N_34632,N_34971);
or U35057 (N_35057,N_34839,N_34778);
nand U35058 (N_35058,N_34523,N_34804);
or U35059 (N_35059,N_34747,N_34574);
and U35060 (N_35060,N_34693,N_34538);
xnor U35061 (N_35061,N_34524,N_34587);
xnor U35062 (N_35062,N_34968,N_34513);
nor U35063 (N_35063,N_34679,N_34683);
xnor U35064 (N_35064,N_34734,N_34633);
nor U35065 (N_35065,N_34733,N_34864);
xor U35066 (N_35066,N_34857,N_34602);
and U35067 (N_35067,N_34808,N_34739);
and U35068 (N_35068,N_34999,N_34500);
nand U35069 (N_35069,N_34564,N_34710);
or U35070 (N_35070,N_34919,N_34600);
xor U35071 (N_35071,N_34884,N_34964);
xnor U35072 (N_35072,N_34947,N_34703);
or U35073 (N_35073,N_34742,N_34985);
or U35074 (N_35074,N_34736,N_34729);
nand U35075 (N_35075,N_34877,N_34939);
xnor U35076 (N_35076,N_34592,N_34581);
xor U35077 (N_35077,N_34780,N_34821);
nor U35078 (N_35078,N_34759,N_34642);
or U35079 (N_35079,N_34636,N_34585);
or U35080 (N_35080,N_34561,N_34510);
nor U35081 (N_35081,N_34897,N_34640);
or U35082 (N_35082,N_34658,N_34505);
xnor U35083 (N_35083,N_34888,N_34989);
nand U35084 (N_35084,N_34746,N_34894);
nand U35085 (N_35085,N_34601,N_34981);
and U35086 (N_35086,N_34668,N_34893);
nor U35087 (N_35087,N_34986,N_34644);
or U35088 (N_35088,N_34547,N_34661);
nor U35089 (N_35089,N_34576,N_34916);
nor U35090 (N_35090,N_34506,N_34797);
nand U35091 (N_35091,N_34973,N_34842);
xor U35092 (N_35092,N_34700,N_34933);
nand U35093 (N_35093,N_34996,N_34714);
xor U35094 (N_35094,N_34537,N_34655);
xnor U35095 (N_35095,N_34536,N_34828);
nand U35096 (N_35096,N_34691,N_34667);
or U35097 (N_35097,N_34611,N_34784);
or U35098 (N_35098,N_34550,N_34928);
and U35099 (N_35099,N_34573,N_34509);
nand U35100 (N_35100,N_34627,N_34695);
and U35101 (N_35101,N_34905,N_34866);
nor U35102 (N_35102,N_34944,N_34948);
xor U35103 (N_35103,N_34631,N_34790);
nand U35104 (N_35104,N_34984,N_34666);
nand U35105 (N_35105,N_34967,N_34868);
or U35106 (N_35106,N_34885,N_34569);
nand U35107 (N_35107,N_34852,N_34607);
nand U35108 (N_35108,N_34593,N_34620);
or U35109 (N_35109,N_34770,N_34533);
or U35110 (N_35110,N_34654,N_34701);
and U35111 (N_35111,N_34961,N_34902);
xor U35112 (N_35112,N_34512,N_34820);
or U35113 (N_35113,N_34907,N_34777);
nand U35114 (N_35114,N_34625,N_34579);
and U35115 (N_35115,N_34577,N_34924);
xnor U35116 (N_35116,N_34818,N_34860);
nand U35117 (N_35117,N_34878,N_34741);
nand U35118 (N_35118,N_34671,N_34713);
nor U35119 (N_35119,N_34656,N_34899);
or U35120 (N_35120,N_34890,N_34844);
nor U35121 (N_35121,N_34623,N_34534);
or U35122 (N_35122,N_34525,N_34603);
and U35123 (N_35123,N_34898,N_34697);
nor U35124 (N_35124,N_34516,N_34687);
xor U35125 (N_35125,N_34979,N_34988);
nor U35126 (N_35126,N_34583,N_34680);
and U35127 (N_35127,N_34911,N_34712);
xor U35128 (N_35128,N_34834,N_34819);
nand U35129 (N_35129,N_34785,N_34681);
nor U35130 (N_35130,N_34977,N_34552);
and U35131 (N_35131,N_34753,N_34624);
xnor U35132 (N_35132,N_34738,N_34931);
nand U35133 (N_35133,N_34673,N_34704);
xor U35134 (N_35134,N_34835,N_34917);
nand U35135 (N_35135,N_34915,N_34855);
nor U35136 (N_35136,N_34745,N_34717);
nor U35137 (N_35137,N_34544,N_34563);
xnor U35138 (N_35138,N_34970,N_34870);
xor U35139 (N_35139,N_34618,N_34775);
xor U35140 (N_35140,N_34501,N_34653);
or U35141 (N_35141,N_34548,N_34726);
nor U35142 (N_35142,N_34912,N_34502);
nand U35143 (N_35143,N_34511,N_34663);
or U35144 (N_35144,N_34597,N_34974);
and U35145 (N_35145,N_34766,N_34722);
and U35146 (N_35146,N_34856,N_34575);
and U35147 (N_35147,N_34508,N_34562);
or U35148 (N_35148,N_34826,N_34814);
xnor U35149 (N_35149,N_34702,N_34960);
xor U35150 (N_35150,N_34598,N_34727);
nor U35151 (N_35151,N_34621,N_34926);
nand U35152 (N_35152,N_34557,N_34558);
xor U35153 (N_35153,N_34591,N_34589);
nor U35154 (N_35154,N_34617,N_34705);
xor U35155 (N_35155,N_34901,N_34983);
or U35156 (N_35156,N_34628,N_34676);
nor U35157 (N_35157,N_34684,N_34637);
nor U35158 (N_35158,N_34692,N_34754);
or U35159 (N_35159,N_34724,N_34689);
nand U35160 (N_35160,N_34530,N_34943);
xnor U35161 (N_35161,N_34837,N_34825);
nand U35162 (N_35162,N_34812,N_34795);
and U35163 (N_35163,N_34662,N_34686);
xnor U35164 (N_35164,N_34881,N_34760);
nor U35165 (N_35165,N_34709,N_34622);
and U35166 (N_35166,N_34720,N_34975);
or U35167 (N_35167,N_34909,N_34648);
and U35168 (N_35168,N_34883,N_34762);
nor U35169 (N_35169,N_34612,N_34675);
and U35170 (N_35170,N_34872,N_34800);
xnor U35171 (N_35171,N_34651,N_34571);
or U35172 (N_35172,N_34694,N_34672);
xnor U35173 (N_35173,N_34887,N_34904);
or U35174 (N_35174,N_34913,N_34590);
nor U35175 (N_35175,N_34929,N_34554);
nand U35176 (N_35176,N_34542,N_34755);
nand U35177 (N_35177,N_34549,N_34876);
xnor U35178 (N_35178,N_34519,N_34993);
nor U35179 (N_35179,N_34716,N_34854);
nor U35180 (N_35180,N_34965,N_34604);
nand U35181 (N_35181,N_34923,N_34731);
or U35182 (N_35182,N_34721,N_34862);
nand U35183 (N_35183,N_34688,N_34748);
and U35184 (N_35184,N_34873,N_34567);
and U35185 (N_35185,N_34998,N_34788);
nor U35186 (N_35186,N_34730,N_34950);
nor U35187 (N_35187,N_34843,N_34906);
and U35188 (N_35188,N_34942,N_34850);
or U35189 (N_35189,N_34782,N_34514);
nor U35190 (N_35190,N_34526,N_34809);
and U35191 (N_35191,N_34531,N_34728);
nand U35192 (N_35192,N_34920,N_34841);
nand U35193 (N_35193,N_34914,N_34517);
nor U35194 (N_35194,N_34723,N_34553);
nor U35195 (N_35195,N_34865,N_34582);
or U35196 (N_35196,N_34832,N_34535);
xnor U35197 (N_35197,N_34749,N_34903);
and U35198 (N_35198,N_34829,N_34817);
nand U35199 (N_35199,N_34769,N_34849);
or U35200 (N_35200,N_34586,N_34838);
nor U35201 (N_35201,N_34836,N_34799);
xor U35202 (N_35202,N_34765,N_34918);
and U35203 (N_35203,N_34639,N_34645);
or U35204 (N_35204,N_34520,N_34889);
xnor U35205 (N_35205,N_34715,N_34696);
and U35206 (N_35206,N_34626,N_34802);
and U35207 (N_35207,N_34806,N_34794);
or U35208 (N_35208,N_34568,N_34540);
and U35209 (N_35209,N_34652,N_34805);
or U35210 (N_35210,N_34665,N_34588);
xnor U35211 (N_35211,N_34605,N_34962);
or U35212 (N_35212,N_34752,N_34781);
and U35213 (N_35213,N_34798,N_34801);
xnor U35214 (N_35214,N_34646,N_34863);
nor U35215 (N_35215,N_34670,N_34750);
nor U35216 (N_35216,N_34565,N_34522);
nor U35217 (N_35217,N_34543,N_34599);
xnor U35218 (N_35218,N_34518,N_34810);
nand U35219 (N_35219,N_34566,N_34616);
nand U35220 (N_35220,N_34732,N_34815);
nand U35221 (N_35221,N_34744,N_34976);
nor U35222 (N_35222,N_34952,N_34725);
and U35223 (N_35223,N_34953,N_34900);
nor U35224 (N_35224,N_34886,N_34823);
and U35225 (N_35225,N_34606,N_34682);
nand U35226 (N_35226,N_34594,N_34718);
and U35227 (N_35227,N_34572,N_34963);
or U35228 (N_35228,N_34690,N_34560);
and U35229 (N_35229,N_34515,N_34707);
nand U35230 (N_35230,N_34629,N_34816);
or U35231 (N_35231,N_34768,N_34927);
or U35232 (N_35232,N_34743,N_34934);
nor U35233 (N_35233,N_34613,N_34756);
or U35234 (N_35234,N_34840,N_34972);
xor U35235 (N_35235,N_34527,N_34764);
and U35236 (N_35236,N_34861,N_34771);
nand U35237 (N_35237,N_34541,N_34529);
and U35238 (N_35238,N_34930,N_34783);
and U35239 (N_35239,N_34875,N_34649);
or U35240 (N_35240,N_34767,N_34647);
nand U35241 (N_35241,N_34503,N_34949);
nand U35242 (N_35242,N_34757,N_34959);
and U35243 (N_35243,N_34532,N_34776);
and U35244 (N_35244,N_34896,N_34895);
nand U35245 (N_35245,N_34685,N_34980);
and U35246 (N_35246,N_34846,N_34643);
nor U35247 (N_35247,N_34991,N_34584);
nor U35248 (N_35248,N_34539,N_34787);
or U35249 (N_35249,N_34925,N_34824);
xnor U35250 (N_35250,N_34704,N_34866);
xor U35251 (N_35251,N_34552,N_34502);
nor U35252 (N_35252,N_34782,N_34510);
and U35253 (N_35253,N_34580,N_34838);
nand U35254 (N_35254,N_34560,N_34534);
and U35255 (N_35255,N_34966,N_34521);
or U35256 (N_35256,N_34552,N_34911);
nand U35257 (N_35257,N_34557,N_34924);
xnor U35258 (N_35258,N_34831,N_34579);
xor U35259 (N_35259,N_34585,N_34763);
nand U35260 (N_35260,N_34719,N_34752);
or U35261 (N_35261,N_34548,N_34773);
or U35262 (N_35262,N_34634,N_34984);
nor U35263 (N_35263,N_34918,N_34704);
xnor U35264 (N_35264,N_34976,N_34876);
xor U35265 (N_35265,N_34681,N_34884);
or U35266 (N_35266,N_34560,N_34967);
xor U35267 (N_35267,N_34592,N_34764);
xnor U35268 (N_35268,N_34532,N_34896);
nor U35269 (N_35269,N_34609,N_34839);
or U35270 (N_35270,N_34585,N_34809);
xnor U35271 (N_35271,N_34892,N_34856);
xor U35272 (N_35272,N_34931,N_34982);
or U35273 (N_35273,N_34532,N_34849);
and U35274 (N_35274,N_34915,N_34731);
or U35275 (N_35275,N_34727,N_34630);
nor U35276 (N_35276,N_34778,N_34922);
nor U35277 (N_35277,N_34723,N_34685);
or U35278 (N_35278,N_34564,N_34744);
and U35279 (N_35279,N_34795,N_34939);
or U35280 (N_35280,N_34631,N_34659);
or U35281 (N_35281,N_34943,N_34783);
xor U35282 (N_35282,N_34987,N_34603);
nor U35283 (N_35283,N_34987,N_34797);
nor U35284 (N_35284,N_34980,N_34779);
nor U35285 (N_35285,N_34693,N_34682);
or U35286 (N_35286,N_34716,N_34897);
and U35287 (N_35287,N_34876,N_34800);
and U35288 (N_35288,N_34940,N_34653);
nand U35289 (N_35289,N_34963,N_34704);
nand U35290 (N_35290,N_34864,N_34541);
nand U35291 (N_35291,N_34786,N_34980);
or U35292 (N_35292,N_34800,N_34887);
or U35293 (N_35293,N_34591,N_34944);
nor U35294 (N_35294,N_34634,N_34672);
and U35295 (N_35295,N_34526,N_34578);
nand U35296 (N_35296,N_34771,N_34602);
and U35297 (N_35297,N_34935,N_34894);
and U35298 (N_35298,N_34945,N_34830);
or U35299 (N_35299,N_34929,N_34548);
or U35300 (N_35300,N_34768,N_34952);
or U35301 (N_35301,N_34581,N_34562);
and U35302 (N_35302,N_34843,N_34534);
xor U35303 (N_35303,N_34815,N_34871);
nor U35304 (N_35304,N_34617,N_34936);
nor U35305 (N_35305,N_34627,N_34643);
and U35306 (N_35306,N_34552,N_34571);
nor U35307 (N_35307,N_34830,N_34844);
and U35308 (N_35308,N_34518,N_34641);
or U35309 (N_35309,N_34581,N_34549);
xor U35310 (N_35310,N_34743,N_34878);
and U35311 (N_35311,N_34663,N_34887);
or U35312 (N_35312,N_34871,N_34804);
or U35313 (N_35313,N_34942,N_34597);
nand U35314 (N_35314,N_34900,N_34709);
or U35315 (N_35315,N_34582,N_34670);
or U35316 (N_35316,N_34640,N_34851);
xnor U35317 (N_35317,N_34542,N_34974);
or U35318 (N_35318,N_34504,N_34585);
nor U35319 (N_35319,N_34692,N_34673);
nor U35320 (N_35320,N_34875,N_34571);
and U35321 (N_35321,N_34940,N_34869);
or U35322 (N_35322,N_34619,N_34854);
nor U35323 (N_35323,N_34641,N_34563);
xnor U35324 (N_35324,N_34853,N_34574);
nand U35325 (N_35325,N_34966,N_34698);
nor U35326 (N_35326,N_34881,N_34580);
and U35327 (N_35327,N_34760,N_34633);
or U35328 (N_35328,N_34719,N_34872);
or U35329 (N_35329,N_34718,N_34516);
or U35330 (N_35330,N_34857,N_34643);
xor U35331 (N_35331,N_34628,N_34587);
or U35332 (N_35332,N_34580,N_34991);
xor U35333 (N_35333,N_34660,N_34581);
nor U35334 (N_35334,N_34711,N_34572);
and U35335 (N_35335,N_34552,N_34605);
nand U35336 (N_35336,N_34989,N_34907);
xnor U35337 (N_35337,N_34901,N_34660);
and U35338 (N_35338,N_34573,N_34992);
xnor U35339 (N_35339,N_34605,N_34902);
or U35340 (N_35340,N_34550,N_34622);
nand U35341 (N_35341,N_34968,N_34817);
xor U35342 (N_35342,N_34585,N_34818);
or U35343 (N_35343,N_34668,N_34920);
nor U35344 (N_35344,N_34593,N_34591);
nand U35345 (N_35345,N_34695,N_34966);
xnor U35346 (N_35346,N_34843,N_34688);
nand U35347 (N_35347,N_34834,N_34690);
nand U35348 (N_35348,N_34636,N_34538);
or U35349 (N_35349,N_34773,N_34686);
xor U35350 (N_35350,N_34517,N_34577);
xnor U35351 (N_35351,N_34938,N_34642);
nor U35352 (N_35352,N_34641,N_34997);
and U35353 (N_35353,N_34707,N_34840);
nand U35354 (N_35354,N_34995,N_34936);
xor U35355 (N_35355,N_34953,N_34740);
nor U35356 (N_35356,N_34503,N_34701);
or U35357 (N_35357,N_34664,N_34626);
or U35358 (N_35358,N_34546,N_34630);
xnor U35359 (N_35359,N_34826,N_34675);
nand U35360 (N_35360,N_34980,N_34546);
nor U35361 (N_35361,N_34773,N_34762);
nor U35362 (N_35362,N_34951,N_34677);
or U35363 (N_35363,N_34525,N_34503);
or U35364 (N_35364,N_34640,N_34580);
xor U35365 (N_35365,N_34955,N_34606);
and U35366 (N_35366,N_34737,N_34976);
and U35367 (N_35367,N_34883,N_34864);
or U35368 (N_35368,N_34610,N_34772);
and U35369 (N_35369,N_34968,N_34800);
xnor U35370 (N_35370,N_34827,N_34978);
xnor U35371 (N_35371,N_34554,N_34634);
xnor U35372 (N_35372,N_34637,N_34619);
nor U35373 (N_35373,N_34579,N_34646);
nor U35374 (N_35374,N_34738,N_34537);
xnor U35375 (N_35375,N_34927,N_34921);
or U35376 (N_35376,N_34895,N_34583);
and U35377 (N_35377,N_34513,N_34719);
xnor U35378 (N_35378,N_34728,N_34753);
nand U35379 (N_35379,N_34810,N_34935);
nand U35380 (N_35380,N_34839,N_34990);
or U35381 (N_35381,N_34822,N_34511);
nand U35382 (N_35382,N_34616,N_34503);
xor U35383 (N_35383,N_34906,N_34509);
or U35384 (N_35384,N_34567,N_34760);
or U35385 (N_35385,N_34995,N_34637);
nor U35386 (N_35386,N_34504,N_34861);
or U35387 (N_35387,N_34985,N_34960);
xnor U35388 (N_35388,N_34795,N_34643);
xor U35389 (N_35389,N_34780,N_34946);
or U35390 (N_35390,N_34930,N_34834);
nand U35391 (N_35391,N_34701,N_34941);
nand U35392 (N_35392,N_34774,N_34517);
nand U35393 (N_35393,N_34955,N_34795);
nand U35394 (N_35394,N_34884,N_34987);
nor U35395 (N_35395,N_34748,N_34860);
xor U35396 (N_35396,N_34650,N_34765);
nor U35397 (N_35397,N_34829,N_34836);
nand U35398 (N_35398,N_34847,N_34694);
nor U35399 (N_35399,N_34832,N_34971);
and U35400 (N_35400,N_34920,N_34674);
or U35401 (N_35401,N_34980,N_34678);
nor U35402 (N_35402,N_34816,N_34897);
nor U35403 (N_35403,N_34991,N_34575);
nor U35404 (N_35404,N_34876,N_34641);
or U35405 (N_35405,N_34544,N_34714);
or U35406 (N_35406,N_34978,N_34739);
and U35407 (N_35407,N_34501,N_34699);
nand U35408 (N_35408,N_34857,N_34595);
xor U35409 (N_35409,N_34634,N_34944);
nand U35410 (N_35410,N_34930,N_34765);
xnor U35411 (N_35411,N_34622,N_34819);
and U35412 (N_35412,N_34778,N_34881);
nor U35413 (N_35413,N_34512,N_34954);
nand U35414 (N_35414,N_34751,N_34643);
xor U35415 (N_35415,N_34842,N_34805);
nor U35416 (N_35416,N_34841,N_34766);
and U35417 (N_35417,N_34938,N_34730);
xnor U35418 (N_35418,N_34977,N_34608);
and U35419 (N_35419,N_34660,N_34568);
nand U35420 (N_35420,N_34909,N_34546);
and U35421 (N_35421,N_34974,N_34547);
or U35422 (N_35422,N_34758,N_34531);
or U35423 (N_35423,N_34882,N_34952);
xor U35424 (N_35424,N_34693,N_34651);
and U35425 (N_35425,N_34627,N_34789);
and U35426 (N_35426,N_34539,N_34650);
nand U35427 (N_35427,N_34780,N_34661);
nor U35428 (N_35428,N_34979,N_34794);
nor U35429 (N_35429,N_34986,N_34903);
or U35430 (N_35430,N_34510,N_34590);
or U35431 (N_35431,N_34679,N_34759);
or U35432 (N_35432,N_34533,N_34602);
nor U35433 (N_35433,N_34856,N_34823);
nor U35434 (N_35434,N_34607,N_34664);
nor U35435 (N_35435,N_34595,N_34848);
and U35436 (N_35436,N_34783,N_34923);
and U35437 (N_35437,N_34972,N_34604);
xor U35438 (N_35438,N_34560,N_34929);
and U35439 (N_35439,N_34779,N_34901);
and U35440 (N_35440,N_34830,N_34921);
nor U35441 (N_35441,N_34720,N_34967);
or U35442 (N_35442,N_34655,N_34878);
nand U35443 (N_35443,N_34648,N_34951);
nor U35444 (N_35444,N_34569,N_34690);
nand U35445 (N_35445,N_34769,N_34818);
xnor U35446 (N_35446,N_34879,N_34697);
nor U35447 (N_35447,N_34802,N_34850);
or U35448 (N_35448,N_34914,N_34942);
or U35449 (N_35449,N_34567,N_34540);
nor U35450 (N_35450,N_34891,N_34763);
and U35451 (N_35451,N_34777,N_34953);
nand U35452 (N_35452,N_34969,N_34723);
nand U35453 (N_35453,N_34872,N_34704);
xnor U35454 (N_35454,N_34586,N_34991);
xnor U35455 (N_35455,N_34760,N_34697);
xnor U35456 (N_35456,N_34940,N_34688);
or U35457 (N_35457,N_34554,N_34638);
nand U35458 (N_35458,N_34613,N_34964);
xor U35459 (N_35459,N_34584,N_34536);
and U35460 (N_35460,N_34873,N_34509);
xor U35461 (N_35461,N_34879,N_34736);
or U35462 (N_35462,N_34779,N_34929);
xor U35463 (N_35463,N_34795,N_34953);
and U35464 (N_35464,N_34694,N_34783);
or U35465 (N_35465,N_34936,N_34830);
nand U35466 (N_35466,N_34638,N_34848);
xnor U35467 (N_35467,N_34934,N_34667);
nor U35468 (N_35468,N_34966,N_34948);
nand U35469 (N_35469,N_34551,N_34863);
or U35470 (N_35470,N_34727,N_34954);
xnor U35471 (N_35471,N_34934,N_34853);
xnor U35472 (N_35472,N_34686,N_34971);
or U35473 (N_35473,N_34966,N_34836);
and U35474 (N_35474,N_34582,N_34604);
nor U35475 (N_35475,N_34664,N_34501);
nand U35476 (N_35476,N_34671,N_34871);
nand U35477 (N_35477,N_34993,N_34522);
or U35478 (N_35478,N_34758,N_34704);
xnor U35479 (N_35479,N_34790,N_34883);
nand U35480 (N_35480,N_34819,N_34541);
or U35481 (N_35481,N_34768,N_34790);
and U35482 (N_35482,N_34993,N_34960);
nor U35483 (N_35483,N_34675,N_34904);
nor U35484 (N_35484,N_34905,N_34618);
xor U35485 (N_35485,N_34687,N_34736);
nor U35486 (N_35486,N_34980,N_34718);
nor U35487 (N_35487,N_34527,N_34884);
and U35488 (N_35488,N_34543,N_34683);
nor U35489 (N_35489,N_34578,N_34556);
nor U35490 (N_35490,N_34578,N_34854);
xor U35491 (N_35491,N_34796,N_34795);
nand U35492 (N_35492,N_34890,N_34684);
or U35493 (N_35493,N_34703,N_34694);
nor U35494 (N_35494,N_34845,N_34824);
and U35495 (N_35495,N_34941,N_34518);
and U35496 (N_35496,N_34747,N_34790);
xnor U35497 (N_35497,N_34507,N_34724);
or U35498 (N_35498,N_34678,N_34908);
nand U35499 (N_35499,N_34898,N_34825);
nor U35500 (N_35500,N_35127,N_35217);
nor U35501 (N_35501,N_35357,N_35448);
nor U35502 (N_35502,N_35422,N_35071);
xnor U35503 (N_35503,N_35451,N_35339);
nor U35504 (N_35504,N_35157,N_35183);
and U35505 (N_35505,N_35450,N_35314);
nor U35506 (N_35506,N_35259,N_35193);
or U35507 (N_35507,N_35036,N_35185);
xor U35508 (N_35508,N_35198,N_35149);
xor U35509 (N_35509,N_35081,N_35122);
nand U35510 (N_35510,N_35444,N_35344);
or U35511 (N_35511,N_35272,N_35351);
nand U35512 (N_35512,N_35225,N_35123);
or U35513 (N_35513,N_35263,N_35464);
xnor U35514 (N_35514,N_35423,N_35385);
or U35515 (N_35515,N_35163,N_35166);
xnor U35516 (N_35516,N_35206,N_35102);
xor U35517 (N_35517,N_35126,N_35396);
nand U35518 (N_35518,N_35147,N_35281);
or U35519 (N_35519,N_35354,N_35466);
nor U35520 (N_35520,N_35400,N_35214);
xor U35521 (N_35521,N_35329,N_35181);
nor U35522 (N_35522,N_35031,N_35349);
nor U35523 (N_35523,N_35401,N_35285);
and U35524 (N_35524,N_35200,N_35276);
nor U35525 (N_35525,N_35017,N_35201);
nand U35526 (N_35526,N_35374,N_35029);
nand U35527 (N_35527,N_35160,N_35256);
nor U35528 (N_35528,N_35076,N_35038);
and U35529 (N_35529,N_35377,N_35268);
nor U35530 (N_35530,N_35155,N_35330);
nand U35531 (N_35531,N_35059,N_35037);
nor U35532 (N_35532,N_35371,N_35194);
nand U35533 (N_35533,N_35300,N_35104);
nand U35534 (N_35534,N_35299,N_35261);
xor U35535 (N_35535,N_35061,N_35048);
or U35536 (N_35536,N_35139,N_35082);
nand U35537 (N_35537,N_35458,N_35387);
and U35538 (N_35538,N_35294,N_35467);
nand U35539 (N_35539,N_35136,N_35121);
xor U35540 (N_35540,N_35493,N_35487);
xor U35541 (N_35541,N_35169,N_35283);
nand U35542 (N_35542,N_35132,N_35352);
and U35543 (N_35543,N_35110,N_35485);
xnor U35544 (N_35544,N_35045,N_35087);
xnor U35545 (N_35545,N_35465,N_35421);
xor U35546 (N_35546,N_35446,N_35328);
nand U35547 (N_35547,N_35057,N_35364);
xor U35548 (N_35548,N_35360,N_35321);
xnor U35549 (N_35549,N_35088,N_35186);
and U35550 (N_35550,N_35437,N_35179);
xnor U35551 (N_35551,N_35405,N_35411);
or U35552 (N_35552,N_35098,N_35095);
or U35553 (N_35553,N_35338,N_35266);
xnor U35554 (N_35554,N_35035,N_35289);
or U35555 (N_35555,N_35106,N_35178);
nand U35556 (N_35556,N_35473,N_35431);
and U35557 (N_35557,N_35222,N_35074);
nor U35558 (N_35558,N_35042,N_35243);
nor U35559 (N_35559,N_35273,N_35288);
or U35560 (N_35560,N_35153,N_35317);
nor U35561 (N_35561,N_35051,N_35196);
or U35562 (N_35562,N_35447,N_35008);
nor U35563 (N_35563,N_35054,N_35184);
xor U35564 (N_35564,N_35327,N_35402);
xor U35565 (N_35565,N_35489,N_35118);
or U35566 (N_35566,N_35303,N_35032);
nand U35567 (N_35567,N_35305,N_35286);
xnor U35568 (N_35568,N_35469,N_35232);
and U35569 (N_35569,N_35372,N_35470);
or U35570 (N_35570,N_35192,N_35416);
nor U35571 (N_35571,N_35237,N_35128);
or U35572 (N_35572,N_35379,N_35412);
nor U35573 (N_35573,N_35430,N_35455);
and U35574 (N_35574,N_35320,N_35226);
xnor U35575 (N_35575,N_35311,N_35063);
nand U35576 (N_35576,N_35207,N_35340);
nor U35577 (N_35577,N_35108,N_35271);
and U35578 (N_35578,N_35066,N_35148);
and U35579 (N_35579,N_35367,N_35420);
xor U35580 (N_35580,N_35060,N_35248);
or U35581 (N_35581,N_35174,N_35004);
xor U35582 (N_35582,N_35393,N_35432);
and U35583 (N_35583,N_35254,N_35052);
or U35584 (N_35584,N_35488,N_35348);
nand U35585 (N_35585,N_35406,N_35041);
xnor U35586 (N_35586,N_35144,N_35424);
or U35587 (N_35587,N_35366,N_35233);
nand U35588 (N_35588,N_35204,N_35274);
nor U35589 (N_35589,N_35199,N_35064);
xnor U35590 (N_35590,N_35461,N_35165);
nand U35591 (N_35591,N_35113,N_35275);
nand U35592 (N_35592,N_35495,N_35075);
xor U35593 (N_35593,N_35101,N_35494);
and U35594 (N_35594,N_35111,N_35456);
nand U35595 (N_35595,N_35449,N_35191);
nor U35596 (N_35596,N_35492,N_35409);
and U35597 (N_35597,N_35323,N_35397);
or U35598 (N_35598,N_35212,N_35152);
or U35599 (N_35599,N_35359,N_35480);
nor U35600 (N_35600,N_35413,N_35429);
or U35601 (N_35601,N_35202,N_35011);
or U35602 (N_35602,N_35114,N_35287);
nor U35603 (N_35603,N_35089,N_35255);
nand U35604 (N_35604,N_35253,N_35053);
nand U35605 (N_35605,N_35213,N_35484);
xnor U35606 (N_35606,N_35270,N_35188);
nor U35607 (N_35607,N_35441,N_35296);
xnor U35608 (N_35608,N_35290,N_35067);
and U35609 (N_35609,N_35389,N_35230);
and U35610 (N_35610,N_35224,N_35369);
xor U35611 (N_35611,N_35282,N_35242);
or U35612 (N_35612,N_35040,N_35180);
nor U35613 (N_35613,N_35249,N_35109);
nor U35614 (N_35614,N_35319,N_35235);
and U35615 (N_35615,N_35105,N_35209);
nor U35616 (N_35616,N_35332,N_35002);
and U35617 (N_35617,N_35361,N_35151);
nand U35618 (N_35618,N_35131,N_35190);
nand U35619 (N_35619,N_35070,N_35245);
or U35620 (N_35620,N_35014,N_35195);
and U35621 (N_35621,N_35310,N_35291);
or U35622 (N_35622,N_35125,N_35384);
or U35623 (N_35623,N_35459,N_35418);
nand U35624 (N_35624,N_35221,N_35069);
xnor U35625 (N_35625,N_35471,N_35313);
nor U35626 (N_35626,N_35007,N_35425);
nand U35627 (N_35627,N_35141,N_35231);
xnor U35628 (N_35628,N_35143,N_35028);
nor U35629 (N_35629,N_35244,N_35238);
and U35630 (N_35630,N_35358,N_35398);
and U35631 (N_35631,N_35050,N_35073);
nand U35632 (N_35632,N_35015,N_35370);
and U35633 (N_35633,N_35172,N_35077);
or U35634 (N_35634,N_35026,N_35262);
xnor U35635 (N_35635,N_35220,N_35043);
nand U35636 (N_35636,N_35468,N_35463);
nand U35637 (N_35637,N_35390,N_35403);
or U35638 (N_35638,N_35404,N_35365);
nand U35639 (N_35639,N_35162,N_35499);
xnor U35640 (N_35640,N_35001,N_35010);
and U35641 (N_35641,N_35307,N_35295);
nand U35642 (N_35642,N_35435,N_35427);
or U35643 (N_35643,N_35177,N_35000);
and U35644 (N_35644,N_35170,N_35216);
nand U35645 (N_35645,N_35247,N_35033);
or U35646 (N_35646,N_35013,N_35312);
xor U35647 (N_35647,N_35280,N_35129);
xnor U35648 (N_35648,N_35150,N_35453);
or U35649 (N_35649,N_35267,N_35086);
or U35650 (N_35650,N_35410,N_35208);
nand U35651 (N_35651,N_35146,N_35161);
nand U35652 (N_35652,N_35115,N_35293);
nand U35653 (N_35653,N_35134,N_35454);
and U35654 (N_35654,N_35100,N_35058);
or U35655 (N_35655,N_35251,N_35333);
nand U35656 (N_35656,N_35353,N_35407);
nor U35657 (N_35657,N_35240,N_35167);
xor U35658 (N_35658,N_35119,N_35419);
xnor U35659 (N_35659,N_35097,N_35414);
and U35660 (N_35660,N_35335,N_35065);
nand U35661 (N_35661,N_35342,N_35496);
or U35662 (N_35662,N_35223,N_35093);
and U35663 (N_35663,N_35391,N_35072);
or U35664 (N_35664,N_35378,N_35439);
nand U35665 (N_35665,N_35080,N_35219);
or U35666 (N_35666,N_35016,N_35375);
nand U35667 (N_35667,N_35306,N_35138);
xor U35668 (N_35668,N_35145,N_35482);
xnor U35669 (N_35669,N_35490,N_35137);
or U35670 (N_35670,N_35443,N_35355);
and U35671 (N_35671,N_35175,N_35047);
and U35672 (N_35672,N_35227,N_35085);
or U35673 (N_35673,N_35373,N_35498);
nor U35674 (N_35674,N_35395,N_35362);
nand U35675 (N_35675,N_35479,N_35483);
nand U35676 (N_35676,N_35246,N_35241);
or U35677 (N_35677,N_35257,N_35331);
xor U35678 (N_35678,N_35046,N_35279);
and U35679 (N_35679,N_35452,N_35383);
and U35680 (N_35680,N_35034,N_35039);
xor U35681 (N_35681,N_35210,N_35445);
nand U35682 (N_35682,N_35229,N_35239);
xor U35683 (N_35683,N_35068,N_35368);
or U35684 (N_35684,N_35124,N_35345);
nor U35685 (N_35685,N_35044,N_35326);
nor U35686 (N_35686,N_35434,N_35252);
and U35687 (N_35687,N_35301,N_35099);
nor U35688 (N_35688,N_35159,N_35096);
xor U35689 (N_35689,N_35158,N_35460);
nor U35690 (N_35690,N_35382,N_35135);
or U35691 (N_35691,N_35055,N_35341);
nor U35692 (N_35692,N_35024,N_35474);
or U35693 (N_35693,N_35325,N_35250);
or U35694 (N_35694,N_35260,N_35302);
xor U35695 (N_35695,N_35164,N_35472);
nand U35696 (N_35696,N_35203,N_35012);
nor U35697 (N_35697,N_35297,N_35103);
and U35698 (N_35698,N_35003,N_35337);
and U35699 (N_35699,N_35117,N_35477);
xor U35700 (N_35700,N_35090,N_35284);
xnor U35701 (N_35701,N_35417,N_35133);
and U35702 (N_35702,N_35234,N_35049);
and U35703 (N_35703,N_35215,N_35324);
nor U35704 (N_35704,N_35176,N_35107);
xnor U35705 (N_35705,N_35020,N_35091);
or U35706 (N_35706,N_35316,N_35497);
nand U35707 (N_35707,N_35092,N_35298);
and U35708 (N_35708,N_35462,N_35440);
or U35709 (N_35709,N_35236,N_35415);
nor U35710 (N_35710,N_35386,N_35350);
nand U35711 (N_35711,N_35381,N_35392);
and U35712 (N_35712,N_35264,N_35171);
nand U35713 (N_35713,N_35187,N_35478);
xor U35714 (N_35714,N_35292,N_35309);
or U35715 (N_35715,N_35457,N_35142);
or U35716 (N_35716,N_35491,N_35258);
nand U35717 (N_35717,N_35356,N_35140);
or U35718 (N_35718,N_35426,N_35376);
and U35719 (N_35719,N_35343,N_35428);
or U35720 (N_35720,N_35436,N_35442);
nand U35721 (N_35721,N_35380,N_35218);
or U35722 (N_35722,N_35308,N_35009);
nand U35723 (N_35723,N_35278,N_35346);
nor U35724 (N_35724,N_35006,N_35363);
xor U35725 (N_35725,N_35168,N_35475);
xnor U35726 (N_35726,N_35336,N_35394);
or U35727 (N_35727,N_35438,N_35022);
nand U35728 (N_35728,N_35156,N_35304);
or U35729 (N_35729,N_35205,N_35120);
xor U35730 (N_35730,N_35189,N_35173);
nand U35731 (N_35731,N_35027,N_35078);
and U35732 (N_35732,N_35269,N_35322);
nand U35733 (N_35733,N_35116,N_35265);
nand U35734 (N_35734,N_35079,N_35023);
nand U35735 (N_35735,N_35228,N_35018);
nor U35736 (N_35736,N_35084,N_35154);
and U35737 (N_35737,N_35025,N_35211);
xor U35738 (N_35738,N_35005,N_35334);
or U35739 (N_35739,N_35486,N_35315);
nand U35740 (N_35740,N_35277,N_35182);
and U35741 (N_35741,N_35094,N_35056);
nor U35742 (N_35742,N_35062,N_35481);
and U35743 (N_35743,N_35433,N_35021);
xnor U35744 (N_35744,N_35318,N_35130);
nor U35745 (N_35745,N_35347,N_35388);
xor U35746 (N_35746,N_35399,N_35197);
and U35747 (N_35747,N_35083,N_35408);
or U35748 (N_35748,N_35112,N_35019);
xnor U35749 (N_35749,N_35030,N_35476);
xnor U35750 (N_35750,N_35080,N_35047);
and U35751 (N_35751,N_35278,N_35368);
or U35752 (N_35752,N_35133,N_35072);
or U35753 (N_35753,N_35093,N_35091);
nand U35754 (N_35754,N_35266,N_35064);
xnor U35755 (N_35755,N_35146,N_35183);
xor U35756 (N_35756,N_35425,N_35185);
nor U35757 (N_35757,N_35293,N_35022);
xor U35758 (N_35758,N_35479,N_35156);
and U35759 (N_35759,N_35126,N_35312);
xor U35760 (N_35760,N_35048,N_35089);
xor U35761 (N_35761,N_35168,N_35253);
nand U35762 (N_35762,N_35403,N_35302);
nor U35763 (N_35763,N_35236,N_35393);
or U35764 (N_35764,N_35300,N_35461);
nor U35765 (N_35765,N_35383,N_35091);
nor U35766 (N_35766,N_35112,N_35447);
nand U35767 (N_35767,N_35393,N_35238);
xnor U35768 (N_35768,N_35255,N_35297);
or U35769 (N_35769,N_35076,N_35374);
and U35770 (N_35770,N_35395,N_35477);
nor U35771 (N_35771,N_35143,N_35099);
nand U35772 (N_35772,N_35017,N_35019);
and U35773 (N_35773,N_35236,N_35460);
and U35774 (N_35774,N_35392,N_35323);
xor U35775 (N_35775,N_35477,N_35424);
nand U35776 (N_35776,N_35487,N_35015);
or U35777 (N_35777,N_35334,N_35312);
xor U35778 (N_35778,N_35322,N_35217);
xor U35779 (N_35779,N_35137,N_35076);
nor U35780 (N_35780,N_35094,N_35191);
nor U35781 (N_35781,N_35276,N_35258);
and U35782 (N_35782,N_35312,N_35350);
nand U35783 (N_35783,N_35206,N_35182);
xor U35784 (N_35784,N_35363,N_35001);
or U35785 (N_35785,N_35124,N_35013);
xor U35786 (N_35786,N_35318,N_35431);
nand U35787 (N_35787,N_35036,N_35104);
xnor U35788 (N_35788,N_35412,N_35021);
xnor U35789 (N_35789,N_35273,N_35080);
xor U35790 (N_35790,N_35202,N_35349);
nor U35791 (N_35791,N_35483,N_35317);
nand U35792 (N_35792,N_35451,N_35187);
nor U35793 (N_35793,N_35137,N_35090);
and U35794 (N_35794,N_35235,N_35064);
or U35795 (N_35795,N_35110,N_35255);
xor U35796 (N_35796,N_35056,N_35015);
nor U35797 (N_35797,N_35222,N_35316);
or U35798 (N_35798,N_35416,N_35490);
xor U35799 (N_35799,N_35463,N_35088);
nand U35800 (N_35800,N_35056,N_35370);
nor U35801 (N_35801,N_35257,N_35384);
nor U35802 (N_35802,N_35253,N_35121);
nand U35803 (N_35803,N_35121,N_35015);
nand U35804 (N_35804,N_35140,N_35423);
xor U35805 (N_35805,N_35170,N_35058);
xor U35806 (N_35806,N_35073,N_35072);
and U35807 (N_35807,N_35396,N_35203);
nor U35808 (N_35808,N_35398,N_35161);
nor U35809 (N_35809,N_35080,N_35381);
and U35810 (N_35810,N_35148,N_35442);
and U35811 (N_35811,N_35295,N_35242);
nand U35812 (N_35812,N_35026,N_35401);
nor U35813 (N_35813,N_35074,N_35087);
xor U35814 (N_35814,N_35036,N_35351);
xnor U35815 (N_35815,N_35023,N_35437);
xor U35816 (N_35816,N_35212,N_35390);
and U35817 (N_35817,N_35181,N_35157);
or U35818 (N_35818,N_35117,N_35431);
xnor U35819 (N_35819,N_35268,N_35396);
or U35820 (N_35820,N_35375,N_35157);
nand U35821 (N_35821,N_35151,N_35492);
nand U35822 (N_35822,N_35055,N_35439);
or U35823 (N_35823,N_35240,N_35489);
nand U35824 (N_35824,N_35442,N_35486);
xnor U35825 (N_35825,N_35070,N_35198);
or U35826 (N_35826,N_35195,N_35006);
and U35827 (N_35827,N_35158,N_35134);
xnor U35828 (N_35828,N_35021,N_35056);
or U35829 (N_35829,N_35057,N_35173);
and U35830 (N_35830,N_35120,N_35458);
nor U35831 (N_35831,N_35441,N_35113);
or U35832 (N_35832,N_35084,N_35168);
or U35833 (N_35833,N_35059,N_35114);
and U35834 (N_35834,N_35017,N_35038);
or U35835 (N_35835,N_35222,N_35077);
nor U35836 (N_35836,N_35214,N_35234);
nand U35837 (N_35837,N_35471,N_35368);
and U35838 (N_35838,N_35316,N_35305);
or U35839 (N_35839,N_35125,N_35119);
nand U35840 (N_35840,N_35425,N_35472);
nor U35841 (N_35841,N_35079,N_35204);
nor U35842 (N_35842,N_35337,N_35234);
xnor U35843 (N_35843,N_35265,N_35367);
nand U35844 (N_35844,N_35330,N_35345);
and U35845 (N_35845,N_35017,N_35334);
and U35846 (N_35846,N_35476,N_35114);
xor U35847 (N_35847,N_35102,N_35243);
and U35848 (N_35848,N_35312,N_35356);
nor U35849 (N_35849,N_35409,N_35226);
and U35850 (N_35850,N_35257,N_35056);
xnor U35851 (N_35851,N_35151,N_35199);
nor U35852 (N_35852,N_35439,N_35193);
and U35853 (N_35853,N_35087,N_35016);
xnor U35854 (N_35854,N_35131,N_35184);
xor U35855 (N_35855,N_35029,N_35270);
xor U35856 (N_35856,N_35199,N_35351);
xor U35857 (N_35857,N_35240,N_35077);
nand U35858 (N_35858,N_35303,N_35292);
xnor U35859 (N_35859,N_35043,N_35103);
nand U35860 (N_35860,N_35120,N_35116);
nor U35861 (N_35861,N_35440,N_35272);
nor U35862 (N_35862,N_35456,N_35156);
xnor U35863 (N_35863,N_35302,N_35418);
xor U35864 (N_35864,N_35055,N_35476);
nor U35865 (N_35865,N_35128,N_35416);
nand U35866 (N_35866,N_35264,N_35026);
nor U35867 (N_35867,N_35258,N_35355);
nor U35868 (N_35868,N_35310,N_35272);
nor U35869 (N_35869,N_35010,N_35365);
nand U35870 (N_35870,N_35275,N_35289);
xor U35871 (N_35871,N_35364,N_35359);
and U35872 (N_35872,N_35125,N_35314);
nor U35873 (N_35873,N_35313,N_35058);
nor U35874 (N_35874,N_35377,N_35114);
and U35875 (N_35875,N_35072,N_35225);
or U35876 (N_35876,N_35286,N_35219);
and U35877 (N_35877,N_35215,N_35162);
and U35878 (N_35878,N_35344,N_35109);
nor U35879 (N_35879,N_35394,N_35314);
nor U35880 (N_35880,N_35362,N_35044);
xor U35881 (N_35881,N_35193,N_35376);
nand U35882 (N_35882,N_35150,N_35357);
nand U35883 (N_35883,N_35221,N_35419);
and U35884 (N_35884,N_35336,N_35391);
nand U35885 (N_35885,N_35227,N_35280);
nor U35886 (N_35886,N_35037,N_35441);
nor U35887 (N_35887,N_35064,N_35355);
nand U35888 (N_35888,N_35049,N_35486);
xor U35889 (N_35889,N_35286,N_35137);
nand U35890 (N_35890,N_35092,N_35055);
and U35891 (N_35891,N_35288,N_35295);
and U35892 (N_35892,N_35303,N_35397);
and U35893 (N_35893,N_35468,N_35296);
or U35894 (N_35894,N_35017,N_35138);
or U35895 (N_35895,N_35391,N_35367);
and U35896 (N_35896,N_35358,N_35207);
nor U35897 (N_35897,N_35111,N_35038);
nand U35898 (N_35898,N_35381,N_35181);
nand U35899 (N_35899,N_35148,N_35450);
xor U35900 (N_35900,N_35398,N_35061);
or U35901 (N_35901,N_35424,N_35247);
nand U35902 (N_35902,N_35386,N_35055);
nor U35903 (N_35903,N_35219,N_35481);
nor U35904 (N_35904,N_35290,N_35422);
nand U35905 (N_35905,N_35206,N_35459);
nand U35906 (N_35906,N_35485,N_35129);
xor U35907 (N_35907,N_35215,N_35278);
nor U35908 (N_35908,N_35400,N_35365);
or U35909 (N_35909,N_35000,N_35251);
or U35910 (N_35910,N_35347,N_35192);
or U35911 (N_35911,N_35119,N_35176);
nand U35912 (N_35912,N_35489,N_35197);
nand U35913 (N_35913,N_35327,N_35105);
or U35914 (N_35914,N_35144,N_35017);
or U35915 (N_35915,N_35248,N_35244);
nor U35916 (N_35916,N_35035,N_35084);
xnor U35917 (N_35917,N_35438,N_35133);
nor U35918 (N_35918,N_35117,N_35179);
and U35919 (N_35919,N_35414,N_35092);
and U35920 (N_35920,N_35358,N_35085);
and U35921 (N_35921,N_35070,N_35307);
and U35922 (N_35922,N_35354,N_35029);
nor U35923 (N_35923,N_35061,N_35325);
or U35924 (N_35924,N_35069,N_35295);
xor U35925 (N_35925,N_35168,N_35211);
xor U35926 (N_35926,N_35394,N_35046);
nor U35927 (N_35927,N_35286,N_35214);
and U35928 (N_35928,N_35030,N_35036);
and U35929 (N_35929,N_35075,N_35285);
or U35930 (N_35930,N_35383,N_35242);
nand U35931 (N_35931,N_35427,N_35446);
xnor U35932 (N_35932,N_35222,N_35408);
and U35933 (N_35933,N_35373,N_35473);
xor U35934 (N_35934,N_35070,N_35452);
nand U35935 (N_35935,N_35125,N_35482);
and U35936 (N_35936,N_35361,N_35341);
or U35937 (N_35937,N_35432,N_35476);
or U35938 (N_35938,N_35247,N_35047);
nand U35939 (N_35939,N_35086,N_35095);
nand U35940 (N_35940,N_35469,N_35138);
nand U35941 (N_35941,N_35146,N_35378);
nor U35942 (N_35942,N_35326,N_35237);
or U35943 (N_35943,N_35376,N_35317);
or U35944 (N_35944,N_35434,N_35076);
xnor U35945 (N_35945,N_35332,N_35328);
and U35946 (N_35946,N_35337,N_35484);
nor U35947 (N_35947,N_35428,N_35019);
nand U35948 (N_35948,N_35154,N_35447);
nor U35949 (N_35949,N_35478,N_35349);
and U35950 (N_35950,N_35263,N_35463);
xor U35951 (N_35951,N_35234,N_35487);
and U35952 (N_35952,N_35173,N_35077);
and U35953 (N_35953,N_35235,N_35304);
nand U35954 (N_35954,N_35499,N_35079);
and U35955 (N_35955,N_35215,N_35160);
or U35956 (N_35956,N_35071,N_35365);
nor U35957 (N_35957,N_35126,N_35149);
and U35958 (N_35958,N_35030,N_35071);
xor U35959 (N_35959,N_35388,N_35431);
nand U35960 (N_35960,N_35237,N_35221);
nand U35961 (N_35961,N_35290,N_35295);
nand U35962 (N_35962,N_35305,N_35462);
and U35963 (N_35963,N_35485,N_35036);
nor U35964 (N_35964,N_35422,N_35001);
xnor U35965 (N_35965,N_35414,N_35218);
or U35966 (N_35966,N_35172,N_35042);
xor U35967 (N_35967,N_35012,N_35417);
nand U35968 (N_35968,N_35400,N_35294);
or U35969 (N_35969,N_35079,N_35349);
nor U35970 (N_35970,N_35176,N_35040);
or U35971 (N_35971,N_35287,N_35112);
and U35972 (N_35972,N_35303,N_35496);
or U35973 (N_35973,N_35357,N_35443);
xnor U35974 (N_35974,N_35033,N_35430);
and U35975 (N_35975,N_35435,N_35499);
nor U35976 (N_35976,N_35228,N_35114);
or U35977 (N_35977,N_35043,N_35260);
xor U35978 (N_35978,N_35245,N_35279);
xnor U35979 (N_35979,N_35484,N_35184);
xnor U35980 (N_35980,N_35094,N_35060);
nor U35981 (N_35981,N_35077,N_35323);
xor U35982 (N_35982,N_35003,N_35482);
nor U35983 (N_35983,N_35072,N_35167);
or U35984 (N_35984,N_35487,N_35454);
xnor U35985 (N_35985,N_35041,N_35471);
nor U35986 (N_35986,N_35007,N_35015);
nand U35987 (N_35987,N_35368,N_35153);
and U35988 (N_35988,N_35257,N_35118);
nand U35989 (N_35989,N_35265,N_35436);
xnor U35990 (N_35990,N_35294,N_35166);
and U35991 (N_35991,N_35458,N_35071);
nor U35992 (N_35992,N_35332,N_35434);
nand U35993 (N_35993,N_35223,N_35389);
nand U35994 (N_35994,N_35212,N_35322);
and U35995 (N_35995,N_35297,N_35139);
nor U35996 (N_35996,N_35122,N_35079);
nor U35997 (N_35997,N_35242,N_35272);
nand U35998 (N_35998,N_35314,N_35239);
and U35999 (N_35999,N_35110,N_35312);
nor U36000 (N_36000,N_35880,N_35649);
nand U36001 (N_36001,N_35692,N_35665);
xnor U36002 (N_36002,N_35801,N_35504);
and U36003 (N_36003,N_35948,N_35572);
and U36004 (N_36004,N_35652,N_35549);
and U36005 (N_36005,N_35562,N_35538);
and U36006 (N_36006,N_35621,N_35785);
and U36007 (N_36007,N_35802,N_35755);
nand U36008 (N_36008,N_35635,N_35990);
nor U36009 (N_36009,N_35569,N_35727);
xor U36010 (N_36010,N_35546,N_35899);
or U36011 (N_36011,N_35852,N_35557);
xor U36012 (N_36012,N_35505,N_35595);
or U36013 (N_36013,N_35689,N_35747);
and U36014 (N_36014,N_35873,N_35932);
xnor U36015 (N_36015,N_35623,N_35981);
or U36016 (N_36016,N_35742,N_35817);
nand U36017 (N_36017,N_35591,N_35667);
xnor U36018 (N_36018,N_35530,N_35512);
nor U36019 (N_36019,N_35641,N_35904);
and U36020 (N_36020,N_35729,N_35881);
xor U36021 (N_36021,N_35977,N_35625);
xnor U36022 (N_36022,N_35638,N_35675);
or U36023 (N_36023,N_35999,N_35519);
and U36024 (N_36024,N_35806,N_35671);
and U36025 (N_36025,N_35712,N_35531);
nor U36026 (N_36026,N_35517,N_35986);
and U36027 (N_36027,N_35878,N_35887);
and U36028 (N_36028,N_35861,N_35753);
nand U36029 (N_36029,N_35745,N_35971);
and U36030 (N_36030,N_35846,N_35944);
nor U36031 (N_36031,N_35574,N_35915);
or U36032 (N_36032,N_35776,N_35658);
xnor U36033 (N_36033,N_35919,N_35643);
nor U36034 (N_36034,N_35525,N_35906);
or U36035 (N_36035,N_35927,N_35735);
xnor U36036 (N_36036,N_35866,N_35763);
nor U36037 (N_36037,N_35653,N_35767);
nor U36038 (N_36038,N_35898,N_35637);
and U36039 (N_36039,N_35679,N_35894);
or U36040 (N_36040,N_35891,N_35993);
nand U36041 (N_36041,N_35811,N_35760);
nand U36042 (N_36042,N_35998,N_35945);
nor U36043 (N_36043,N_35959,N_35740);
xnor U36044 (N_36044,N_35573,N_35568);
and U36045 (N_36045,N_35644,N_35983);
xnor U36046 (N_36046,N_35940,N_35500);
and U36047 (N_36047,N_35989,N_35600);
nand U36048 (N_36048,N_35654,N_35870);
xor U36049 (N_36049,N_35553,N_35547);
nor U36050 (N_36050,N_35624,N_35699);
or U36051 (N_36051,N_35849,N_35963);
nand U36052 (N_36052,N_35586,N_35656);
xnor U36053 (N_36053,N_35892,N_35579);
nor U36054 (N_36054,N_35765,N_35929);
xnor U36055 (N_36055,N_35795,N_35863);
nor U36056 (N_36056,N_35506,N_35746);
and U36057 (N_36057,N_35698,N_35736);
or U36058 (N_36058,N_35916,N_35961);
xnor U36059 (N_36059,N_35908,N_35951);
nor U36060 (N_36060,N_35516,N_35994);
nand U36061 (N_36061,N_35859,N_35783);
and U36062 (N_36062,N_35770,N_35888);
nand U36063 (N_36063,N_35613,N_35634);
xor U36064 (N_36064,N_35732,N_35616);
or U36065 (N_36065,N_35905,N_35956);
xor U36066 (N_36066,N_35840,N_35851);
nor U36067 (N_36067,N_35936,N_35758);
or U36068 (N_36068,N_35798,N_35545);
or U36069 (N_36069,N_35576,N_35722);
nand U36070 (N_36070,N_35787,N_35819);
xor U36071 (N_36071,N_35800,N_35781);
or U36072 (N_36072,N_35918,N_35604);
nor U36073 (N_36073,N_35877,N_35669);
or U36074 (N_36074,N_35743,N_35921);
or U36075 (N_36075,N_35911,N_35885);
nor U36076 (N_36076,N_35879,N_35782);
and U36077 (N_36077,N_35681,N_35741);
nor U36078 (N_36078,N_35552,N_35672);
nand U36079 (N_36079,N_35833,N_35984);
and U36080 (N_36080,N_35587,N_35633);
nand U36081 (N_36081,N_35701,N_35839);
or U36082 (N_36082,N_35834,N_35578);
nor U36083 (N_36083,N_35555,N_35780);
nand U36084 (N_36084,N_35651,N_35571);
or U36085 (N_36085,N_35813,N_35541);
or U36086 (N_36086,N_35510,N_35966);
nand U36087 (N_36087,N_35594,N_35793);
nand U36088 (N_36088,N_35581,N_35855);
nand U36089 (N_36089,N_35975,N_35639);
or U36090 (N_36090,N_35985,N_35559);
nor U36091 (N_36091,N_35827,N_35872);
nor U36092 (N_36092,N_35564,N_35799);
or U36093 (N_36093,N_35874,N_35942);
nand U36094 (N_36094,N_35841,N_35536);
xor U36095 (N_36095,N_35982,N_35717);
and U36096 (N_36096,N_35901,N_35766);
and U36097 (N_36097,N_35968,N_35540);
xnor U36098 (N_36098,N_35853,N_35821);
nor U36099 (N_36099,N_35589,N_35804);
nor U36100 (N_36100,N_35752,N_35797);
nand U36101 (N_36101,N_35835,N_35693);
nand U36102 (N_36102,N_35764,N_35514);
and U36103 (N_36103,N_35721,N_35734);
nor U36104 (N_36104,N_35532,N_35503);
nand U36105 (N_36105,N_35596,N_35744);
nand U36106 (N_36106,N_35969,N_35580);
nor U36107 (N_36107,N_35836,N_35809);
xor U36108 (N_36108,N_35676,N_35978);
nand U36109 (N_36109,N_35768,N_35593);
nand U36110 (N_36110,N_35778,N_35823);
nand U36111 (N_36111,N_35537,N_35920);
nor U36112 (N_36112,N_35958,N_35794);
nor U36113 (N_36113,N_35903,N_35749);
xor U36114 (N_36114,N_35726,N_35640);
or U36115 (N_36115,N_35524,N_35756);
nor U36116 (N_36116,N_35627,N_35923);
xnor U36117 (N_36117,N_35738,N_35997);
or U36118 (N_36118,N_35703,N_35714);
and U36119 (N_36119,N_35868,N_35584);
nand U36120 (N_36120,N_35660,N_35677);
or U36121 (N_36121,N_35526,N_35709);
xor U36122 (N_36122,N_35612,N_35825);
nor U36123 (N_36123,N_35535,N_35928);
or U36124 (N_36124,N_35611,N_35558);
nand U36125 (N_36125,N_35934,N_35523);
and U36126 (N_36126,N_35790,N_35869);
xor U36127 (N_36127,N_35702,N_35824);
xor U36128 (N_36128,N_35585,N_35583);
xor U36129 (N_36129,N_35931,N_35862);
xnor U36130 (N_36130,N_35622,N_35960);
or U36131 (N_36131,N_35707,N_35691);
and U36132 (N_36132,N_35647,N_35886);
nand U36133 (N_36133,N_35914,N_35694);
xnor U36134 (N_36134,N_35501,N_35715);
or U36135 (N_36135,N_35737,N_35664);
nand U36136 (N_36136,N_35803,N_35662);
xor U36137 (N_36137,N_35987,N_35631);
or U36138 (N_36138,N_35848,N_35561);
xnor U36139 (N_36139,N_35609,N_35567);
nor U36140 (N_36140,N_35954,N_35864);
xor U36141 (N_36141,N_35871,N_35507);
xor U36142 (N_36142,N_35674,N_35509);
or U36143 (N_36143,N_35724,N_35808);
nor U36144 (N_36144,N_35970,N_35617);
and U36145 (N_36145,N_35713,N_35615);
xnor U36146 (N_36146,N_35935,N_35543);
nor U36147 (N_36147,N_35511,N_35807);
xor U36148 (N_36148,N_35889,N_35947);
or U36149 (N_36149,N_35720,N_35774);
and U36150 (N_36150,N_35614,N_35933);
xor U36151 (N_36151,N_35599,N_35648);
and U36152 (N_36152,N_35771,N_35937);
and U36153 (N_36153,N_35542,N_35534);
or U36154 (N_36154,N_35645,N_35812);
or U36155 (N_36155,N_35815,N_35902);
or U36156 (N_36156,N_35603,N_35730);
nand U36157 (N_36157,N_35816,N_35706);
and U36158 (N_36158,N_35518,N_35792);
and U36159 (N_36159,N_35759,N_35551);
and U36160 (N_36160,N_35723,N_35943);
or U36161 (N_36161,N_35605,N_35661);
nor U36162 (N_36162,N_35688,N_35831);
nand U36163 (N_36163,N_35708,N_35527);
and U36164 (N_36164,N_35704,N_35773);
and U36165 (N_36165,N_35907,N_35655);
nor U36166 (N_36166,N_35750,N_35754);
nand U36167 (N_36167,N_35762,N_35979);
nor U36168 (N_36168,N_35590,N_35913);
nand U36169 (N_36169,N_35965,N_35520);
nand U36170 (N_36170,N_35521,N_35854);
and U36171 (N_36171,N_35618,N_35900);
or U36172 (N_36172,N_35897,N_35533);
or U36173 (N_36173,N_35739,N_35528);
or U36174 (N_36174,N_35857,N_35974);
nor U36175 (N_36175,N_35620,N_35629);
and U36176 (N_36176,N_35630,N_35563);
xnor U36177 (N_36177,N_35619,N_35560);
or U36178 (N_36178,N_35964,N_35922);
nand U36179 (N_36179,N_35992,N_35515);
nand U36180 (N_36180,N_35912,N_35976);
or U36181 (N_36181,N_35626,N_35601);
and U36182 (N_36182,N_35941,N_35716);
and U36183 (N_36183,N_35733,N_35867);
xor U36184 (N_36184,N_35950,N_35845);
nand U36185 (N_36185,N_35632,N_35847);
or U36186 (N_36186,N_35683,N_35636);
or U36187 (N_36187,N_35842,N_35577);
and U36188 (N_36188,N_35829,N_35876);
xor U36189 (N_36189,N_35769,N_35687);
nand U36190 (N_36190,N_35598,N_35554);
and U36191 (N_36191,N_35610,N_35988);
xnor U36192 (N_36192,N_35882,N_35991);
and U36193 (N_36193,N_35678,N_35796);
nor U36194 (N_36194,N_35779,N_35939);
and U36195 (N_36195,N_35843,N_35711);
nand U36196 (N_36196,N_35957,N_35751);
and U36197 (N_36197,N_35772,N_35895);
nor U36198 (N_36198,N_35684,N_35725);
nor U36199 (N_36199,N_35565,N_35513);
nand U36200 (N_36200,N_35522,N_35502);
and U36201 (N_36201,N_35659,N_35850);
nand U36202 (N_36202,N_35777,N_35710);
or U36203 (N_36203,N_35925,N_35628);
nor U36204 (N_36204,N_35875,N_35731);
xnor U36205 (N_36205,N_35909,N_35728);
or U36206 (N_36206,N_35930,N_35910);
nor U36207 (N_36207,N_35607,N_35953);
and U36208 (N_36208,N_35663,N_35697);
xor U36209 (N_36209,N_35818,N_35860);
or U36210 (N_36210,N_35788,N_35972);
xor U36211 (N_36211,N_35666,N_35805);
nand U36212 (N_36212,N_35826,N_35686);
nor U36213 (N_36213,N_35592,N_35890);
nand U36214 (N_36214,N_35784,N_35883);
xnor U36215 (N_36215,N_35865,N_35657);
xnor U36216 (N_36216,N_35757,N_35996);
nand U36217 (N_36217,N_35588,N_35838);
or U36218 (N_36218,N_35575,N_35582);
xnor U36219 (N_36219,N_35837,N_35539);
and U36220 (N_36220,N_35566,N_35967);
nor U36221 (N_36221,N_35608,N_35844);
or U36222 (N_36222,N_35810,N_35650);
and U36223 (N_36223,N_35670,N_35548);
and U36224 (N_36224,N_35938,N_35775);
nor U36225 (N_36225,N_35700,N_35789);
nor U36226 (N_36226,N_35508,N_35761);
xor U36227 (N_36227,N_35544,N_35597);
and U36228 (N_36228,N_35832,N_35550);
nor U36229 (N_36229,N_35926,N_35748);
or U36230 (N_36230,N_35696,N_35830);
xnor U36231 (N_36231,N_35680,N_35642);
nand U36232 (N_36232,N_35952,N_35690);
and U36233 (N_36233,N_35858,N_35822);
nand U36234 (N_36234,N_35570,N_35820);
nor U36235 (N_36235,N_35529,N_35718);
nand U36236 (N_36236,N_35856,N_35646);
or U36237 (N_36237,N_35917,N_35682);
or U36238 (N_36238,N_35995,N_35668);
nand U36239 (N_36239,N_35828,N_35719);
nor U36240 (N_36240,N_35602,N_35896);
nand U36241 (N_36241,N_35786,N_35673);
xnor U36242 (N_36242,N_35962,N_35606);
and U36243 (N_36243,N_35946,N_35924);
nand U36244 (N_36244,N_35695,N_35556);
nand U36245 (N_36245,N_35973,N_35980);
and U36246 (N_36246,N_35893,N_35949);
xnor U36247 (N_36247,N_35791,N_35685);
nor U36248 (N_36248,N_35884,N_35955);
xor U36249 (N_36249,N_35705,N_35814);
and U36250 (N_36250,N_35907,N_35814);
nor U36251 (N_36251,N_35612,N_35962);
nand U36252 (N_36252,N_35876,N_35550);
nor U36253 (N_36253,N_35522,N_35720);
or U36254 (N_36254,N_35693,N_35639);
nand U36255 (N_36255,N_35811,N_35974);
xnor U36256 (N_36256,N_35934,N_35863);
and U36257 (N_36257,N_35525,N_35915);
or U36258 (N_36258,N_35770,N_35979);
or U36259 (N_36259,N_35797,N_35600);
nor U36260 (N_36260,N_35843,N_35898);
and U36261 (N_36261,N_35770,N_35576);
or U36262 (N_36262,N_35587,N_35562);
nand U36263 (N_36263,N_35962,N_35989);
xnor U36264 (N_36264,N_35685,N_35985);
nand U36265 (N_36265,N_35679,N_35887);
or U36266 (N_36266,N_35765,N_35819);
and U36267 (N_36267,N_35703,N_35768);
nand U36268 (N_36268,N_35669,N_35959);
or U36269 (N_36269,N_35569,N_35539);
nand U36270 (N_36270,N_35891,N_35506);
nor U36271 (N_36271,N_35734,N_35749);
or U36272 (N_36272,N_35907,N_35988);
or U36273 (N_36273,N_35859,N_35928);
nand U36274 (N_36274,N_35988,N_35715);
xor U36275 (N_36275,N_35961,N_35588);
nand U36276 (N_36276,N_35545,N_35674);
or U36277 (N_36277,N_35802,N_35915);
nor U36278 (N_36278,N_35959,N_35883);
xnor U36279 (N_36279,N_35921,N_35556);
nand U36280 (N_36280,N_35647,N_35594);
xnor U36281 (N_36281,N_35703,N_35622);
and U36282 (N_36282,N_35843,N_35871);
xnor U36283 (N_36283,N_35989,N_35725);
and U36284 (N_36284,N_35626,N_35851);
and U36285 (N_36285,N_35785,N_35522);
nand U36286 (N_36286,N_35750,N_35541);
and U36287 (N_36287,N_35804,N_35741);
xnor U36288 (N_36288,N_35864,N_35698);
nor U36289 (N_36289,N_35770,N_35715);
xor U36290 (N_36290,N_35601,N_35680);
or U36291 (N_36291,N_35887,N_35721);
and U36292 (N_36292,N_35997,N_35902);
nor U36293 (N_36293,N_35857,N_35530);
nand U36294 (N_36294,N_35875,N_35911);
and U36295 (N_36295,N_35772,N_35873);
or U36296 (N_36296,N_35931,N_35653);
xnor U36297 (N_36297,N_35704,N_35929);
xnor U36298 (N_36298,N_35883,N_35774);
and U36299 (N_36299,N_35987,N_35843);
or U36300 (N_36300,N_35961,N_35930);
nand U36301 (N_36301,N_35930,N_35781);
or U36302 (N_36302,N_35966,N_35722);
and U36303 (N_36303,N_35946,N_35822);
xnor U36304 (N_36304,N_35746,N_35861);
nor U36305 (N_36305,N_35738,N_35628);
nand U36306 (N_36306,N_35564,N_35973);
nor U36307 (N_36307,N_35782,N_35590);
and U36308 (N_36308,N_35985,N_35933);
xor U36309 (N_36309,N_35916,N_35662);
and U36310 (N_36310,N_35641,N_35682);
or U36311 (N_36311,N_35983,N_35674);
or U36312 (N_36312,N_35504,N_35532);
nand U36313 (N_36313,N_35710,N_35561);
nand U36314 (N_36314,N_35502,N_35757);
nand U36315 (N_36315,N_35688,N_35524);
and U36316 (N_36316,N_35535,N_35657);
xor U36317 (N_36317,N_35725,N_35552);
and U36318 (N_36318,N_35958,N_35851);
nand U36319 (N_36319,N_35765,N_35789);
and U36320 (N_36320,N_35976,N_35806);
nor U36321 (N_36321,N_35790,N_35548);
nor U36322 (N_36322,N_35677,N_35663);
or U36323 (N_36323,N_35640,N_35831);
nand U36324 (N_36324,N_35811,N_35666);
or U36325 (N_36325,N_35968,N_35975);
nor U36326 (N_36326,N_35833,N_35707);
nand U36327 (N_36327,N_35727,N_35647);
nand U36328 (N_36328,N_35564,N_35914);
nor U36329 (N_36329,N_35769,N_35907);
xnor U36330 (N_36330,N_35810,N_35687);
or U36331 (N_36331,N_35552,N_35948);
nand U36332 (N_36332,N_35783,N_35979);
and U36333 (N_36333,N_35623,N_35854);
nor U36334 (N_36334,N_35980,N_35721);
nand U36335 (N_36335,N_35692,N_35627);
nor U36336 (N_36336,N_35853,N_35678);
or U36337 (N_36337,N_35520,N_35833);
or U36338 (N_36338,N_35784,N_35625);
nor U36339 (N_36339,N_35573,N_35720);
xnor U36340 (N_36340,N_35823,N_35721);
or U36341 (N_36341,N_35712,N_35544);
nand U36342 (N_36342,N_35783,N_35693);
xor U36343 (N_36343,N_35798,N_35775);
nand U36344 (N_36344,N_35813,N_35978);
nand U36345 (N_36345,N_35618,N_35571);
nor U36346 (N_36346,N_35753,N_35582);
and U36347 (N_36347,N_35595,N_35840);
and U36348 (N_36348,N_35946,N_35768);
nand U36349 (N_36349,N_35647,N_35692);
nor U36350 (N_36350,N_35696,N_35624);
xor U36351 (N_36351,N_35629,N_35564);
nand U36352 (N_36352,N_35858,N_35553);
nor U36353 (N_36353,N_35520,N_35793);
and U36354 (N_36354,N_35586,N_35879);
and U36355 (N_36355,N_35858,N_35991);
nand U36356 (N_36356,N_35842,N_35555);
and U36357 (N_36357,N_35650,N_35787);
nor U36358 (N_36358,N_35764,N_35719);
nand U36359 (N_36359,N_35806,N_35784);
xor U36360 (N_36360,N_35712,N_35599);
xor U36361 (N_36361,N_35977,N_35887);
or U36362 (N_36362,N_35575,N_35754);
nand U36363 (N_36363,N_35833,N_35788);
and U36364 (N_36364,N_35530,N_35709);
and U36365 (N_36365,N_35714,N_35887);
nor U36366 (N_36366,N_35680,N_35827);
or U36367 (N_36367,N_35751,N_35583);
nand U36368 (N_36368,N_35776,N_35636);
xor U36369 (N_36369,N_35930,N_35582);
nand U36370 (N_36370,N_35885,N_35720);
and U36371 (N_36371,N_35719,N_35555);
and U36372 (N_36372,N_35879,N_35893);
and U36373 (N_36373,N_35941,N_35569);
or U36374 (N_36374,N_35959,N_35676);
and U36375 (N_36375,N_35695,N_35991);
nand U36376 (N_36376,N_35928,N_35826);
or U36377 (N_36377,N_35965,N_35973);
nor U36378 (N_36378,N_35751,N_35550);
and U36379 (N_36379,N_35768,N_35595);
nor U36380 (N_36380,N_35584,N_35537);
and U36381 (N_36381,N_35947,N_35958);
or U36382 (N_36382,N_35875,N_35812);
nor U36383 (N_36383,N_35678,N_35858);
nor U36384 (N_36384,N_35995,N_35823);
xnor U36385 (N_36385,N_35690,N_35848);
or U36386 (N_36386,N_35809,N_35806);
xor U36387 (N_36387,N_35952,N_35541);
or U36388 (N_36388,N_35722,N_35907);
nand U36389 (N_36389,N_35864,N_35953);
or U36390 (N_36390,N_35841,N_35769);
or U36391 (N_36391,N_35538,N_35605);
or U36392 (N_36392,N_35751,N_35625);
nor U36393 (N_36393,N_35757,N_35930);
nor U36394 (N_36394,N_35613,N_35715);
nand U36395 (N_36395,N_35937,N_35787);
nand U36396 (N_36396,N_35997,N_35797);
nor U36397 (N_36397,N_35656,N_35867);
nor U36398 (N_36398,N_35629,N_35945);
and U36399 (N_36399,N_35923,N_35859);
nand U36400 (N_36400,N_35781,N_35981);
or U36401 (N_36401,N_35879,N_35788);
and U36402 (N_36402,N_35651,N_35827);
xnor U36403 (N_36403,N_35510,N_35533);
nor U36404 (N_36404,N_35539,N_35662);
or U36405 (N_36405,N_35995,N_35986);
and U36406 (N_36406,N_35960,N_35615);
nand U36407 (N_36407,N_35795,N_35942);
or U36408 (N_36408,N_35885,N_35656);
or U36409 (N_36409,N_35829,N_35619);
and U36410 (N_36410,N_35564,N_35501);
xnor U36411 (N_36411,N_35711,N_35615);
nand U36412 (N_36412,N_35910,N_35800);
or U36413 (N_36413,N_35540,N_35934);
and U36414 (N_36414,N_35855,N_35794);
nor U36415 (N_36415,N_35738,N_35817);
nor U36416 (N_36416,N_35548,N_35515);
xor U36417 (N_36417,N_35762,N_35750);
or U36418 (N_36418,N_35943,N_35578);
nor U36419 (N_36419,N_35833,N_35559);
or U36420 (N_36420,N_35852,N_35664);
or U36421 (N_36421,N_35898,N_35784);
xnor U36422 (N_36422,N_35535,N_35914);
nand U36423 (N_36423,N_35624,N_35898);
nor U36424 (N_36424,N_35986,N_35748);
or U36425 (N_36425,N_35983,N_35595);
nand U36426 (N_36426,N_35614,N_35779);
nand U36427 (N_36427,N_35922,N_35832);
and U36428 (N_36428,N_35582,N_35838);
or U36429 (N_36429,N_35829,N_35786);
nor U36430 (N_36430,N_35623,N_35837);
xnor U36431 (N_36431,N_35765,N_35541);
or U36432 (N_36432,N_35684,N_35938);
or U36433 (N_36433,N_35527,N_35998);
or U36434 (N_36434,N_35790,N_35998);
or U36435 (N_36435,N_35531,N_35882);
nand U36436 (N_36436,N_35698,N_35687);
nand U36437 (N_36437,N_35890,N_35833);
nand U36438 (N_36438,N_35599,N_35878);
nand U36439 (N_36439,N_35531,N_35811);
or U36440 (N_36440,N_35892,N_35621);
nand U36441 (N_36441,N_35639,N_35544);
nand U36442 (N_36442,N_35911,N_35871);
or U36443 (N_36443,N_35672,N_35521);
or U36444 (N_36444,N_35975,N_35905);
or U36445 (N_36445,N_35635,N_35629);
xor U36446 (N_36446,N_35679,N_35959);
xnor U36447 (N_36447,N_35536,N_35605);
and U36448 (N_36448,N_35664,N_35756);
or U36449 (N_36449,N_35812,N_35746);
xor U36450 (N_36450,N_35590,N_35920);
or U36451 (N_36451,N_35752,N_35584);
and U36452 (N_36452,N_35539,N_35744);
and U36453 (N_36453,N_35943,N_35818);
nor U36454 (N_36454,N_35726,N_35504);
nor U36455 (N_36455,N_35964,N_35965);
nor U36456 (N_36456,N_35995,N_35831);
xor U36457 (N_36457,N_35965,N_35621);
or U36458 (N_36458,N_35868,N_35778);
or U36459 (N_36459,N_35895,N_35744);
or U36460 (N_36460,N_35544,N_35966);
and U36461 (N_36461,N_35939,N_35787);
nor U36462 (N_36462,N_35862,N_35740);
nand U36463 (N_36463,N_35784,N_35677);
nor U36464 (N_36464,N_35893,N_35578);
and U36465 (N_36465,N_35706,N_35741);
nor U36466 (N_36466,N_35576,N_35679);
or U36467 (N_36467,N_35570,N_35733);
and U36468 (N_36468,N_35980,N_35794);
xor U36469 (N_36469,N_35892,N_35842);
nor U36470 (N_36470,N_35938,N_35589);
and U36471 (N_36471,N_35929,N_35991);
and U36472 (N_36472,N_35508,N_35824);
nor U36473 (N_36473,N_35536,N_35521);
nand U36474 (N_36474,N_35716,N_35538);
or U36475 (N_36475,N_35871,N_35673);
and U36476 (N_36476,N_35605,N_35737);
nand U36477 (N_36477,N_35840,N_35985);
nor U36478 (N_36478,N_35537,N_35905);
nor U36479 (N_36479,N_35616,N_35922);
nand U36480 (N_36480,N_35607,N_35633);
xor U36481 (N_36481,N_35848,N_35621);
or U36482 (N_36482,N_35955,N_35574);
or U36483 (N_36483,N_35644,N_35906);
nor U36484 (N_36484,N_35773,N_35836);
nor U36485 (N_36485,N_35635,N_35589);
nor U36486 (N_36486,N_35665,N_35546);
nor U36487 (N_36487,N_35561,N_35999);
xor U36488 (N_36488,N_35947,N_35653);
nand U36489 (N_36489,N_35612,N_35696);
and U36490 (N_36490,N_35628,N_35870);
nor U36491 (N_36491,N_35681,N_35533);
nand U36492 (N_36492,N_35544,N_35696);
nor U36493 (N_36493,N_35504,N_35581);
and U36494 (N_36494,N_35762,N_35902);
nor U36495 (N_36495,N_35944,N_35697);
and U36496 (N_36496,N_35922,N_35662);
xor U36497 (N_36497,N_35609,N_35848);
or U36498 (N_36498,N_35662,N_35959);
nand U36499 (N_36499,N_35551,N_35994);
or U36500 (N_36500,N_36042,N_36077);
or U36501 (N_36501,N_36204,N_36103);
or U36502 (N_36502,N_36378,N_36478);
nand U36503 (N_36503,N_36376,N_36245);
and U36504 (N_36504,N_36238,N_36106);
and U36505 (N_36505,N_36421,N_36315);
or U36506 (N_36506,N_36325,N_36097);
nand U36507 (N_36507,N_36021,N_36467);
xnor U36508 (N_36508,N_36131,N_36236);
nand U36509 (N_36509,N_36076,N_36407);
and U36510 (N_36510,N_36203,N_36200);
nor U36511 (N_36511,N_36011,N_36473);
and U36512 (N_36512,N_36453,N_36486);
and U36513 (N_36513,N_36319,N_36424);
nor U36514 (N_36514,N_36208,N_36457);
and U36515 (N_36515,N_36195,N_36252);
or U36516 (N_36516,N_36328,N_36210);
nor U36517 (N_36517,N_36072,N_36334);
nor U36518 (N_36518,N_36257,N_36029);
nand U36519 (N_36519,N_36189,N_36154);
xor U36520 (N_36520,N_36332,N_36417);
nand U36521 (N_36521,N_36192,N_36469);
and U36522 (N_36522,N_36498,N_36307);
nand U36523 (N_36523,N_36085,N_36070);
and U36524 (N_36524,N_36089,N_36460);
nand U36525 (N_36525,N_36401,N_36005);
and U36526 (N_36526,N_36282,N_36000);
xnor U36527 (N_36527,N_36162,N_36350);
nor U36528 (N_36528,N_36436,N_36003);
or U36529 (N_36529,N_36080,N_36191);
nor U36530 (N_36530,N_36057,N_36043);
nor U36531 (N_36531,N_36355,N_36234);
and U36532 (N_36532,N_36260,N_36075);
xnor U36533 (N_36533,N_36489,N_36354);
nor U36534 (N_36534,N_36285,N_36212);
nand U36535 (N_36535,N_36109,N_36296);
xnor U36536 (N_36536,N_36441,N_36083);
nor U36537 (N_36537,N_36311,N_36430);
xnor U36538 (N_36538,N_36400,N_36199);
and U36539 (N_36539,N_36037,N_36278);
nand U36540 (N_36540,N_36362,N_36277);
nand U36541 (N_36541,N_36027,N_36004);
nor U36542 (N_36542,N_36348,N_36454);
or U36543 (N_36543,N_36187,N_36279);
xor U36544 (N_36544,N_36286,N_36496);
or U36545 (N_36545,N_36410,N_36019);
xor U36546 (N_36546,N_36049,N_36024);
xor U36547 (N_36547,N_36048,N_36265);
and U36548 (N_36548,N_36146,N_36062);
nor U36549 (N_36549,N_36125,N_36082);
and U36550 (N_36550,N_36133,N_36312);
nand U36551 (N_36551,N_36117,N_36433);
or U36552 (N_36552,N_36351,N_36113);
xnor U36553 (N_36553,N_36287,N_36389);
or U36554 (N_36554,N_36377,N_36026);
nand U36555 (N_36555,N_36206,N_36357);
xor U36556 (N_36556,N_36263,N_36463);
nor U36557 (N_36557,N_36405,N_36333);
and U36558 (N_36558,N_36120,N_36174);
and U36559 (N_36559,N_36258,N_36472);
xnor U36560 (N_36560,N_36305,N_36214);
and U36561 (N_36561,N_36318,N_36339);
nor U36562 (N_36562,N_36336,N_36255);
or U36563 (N_36563,N_36313,N_36271);
xor U36564 (N_36564,N_36017,N_36155);
nor U36565 (N_36565,N_36274,N_36012);
xnor U36566 (N_36566,N_36244,N_36101);
xnor U36567 (N_36567,N_36159,N_36451);
xnor U36568 (N_36568,N_36253,N_36338);
and U36569 (N_36569,N_36134,N_36020);
nor U36570 (N_36570,N_36414,N_36492);
nor U36571 (N_36571,N_36322,N_36055);
or U36572 (N_36572,N_36434,N_36108);
nor U36573 (N_36573,N_36280,N_36440);
xor U36574 (N_36574,N_36297,N_36471);
nor U36575 (N_36575,N_36122,N_36152);
nor U36576 (N_36576,N_36160,N_36474);
or U36577 (N_36577,N_36481,N_36235);
and U36578 (N_36578,N_36476,N_36197);
xnor U36579 (N_36579,N_36078,N_36010);
or U36580 (N_36580,N_36015,N_36326);
xnor U36581 (N_36581,N_36262,N_36217);
and U36582 (N_36582,N_36161,N_36237);
nor U36583 (N_36583,N_36053,N_36371);
or U36584 (N_36584,N_36395,N_36304);
nor U36585 (N_36585,N_36095,N_36446);
xor U36586 (N_36586,N_36393,N_36046);
xnor U36587 (N_36587,N_36018,N_36028);
xnor U36588 (N_36588,N_36182,N_36099);
nand U36589 (N_36589,N_36294,N_36135);
nand U36590 (N_36590,N_36115,N_36231);
and U36591 (N_36591,N_36107,N_36181);
xnor U36592 (N_36592,N_36205,N_36466);
and U36593 (N_36593,N_36419,N_36216);
or U36594 (N_36594,N_36295,N_36105);
xor U36595 (N_36595,N_36386,N_36458);
nor U36596 (N_36596,N_36063,N_36060);
xor U36597 (N_36597,N_36058,N_36227);
nand U36598 (N_36598,N_36173,N_36218);
or U36599 (N_36599,N_36284,N_36143);
or U36600 (N_36600,N_36270,N_36121);
nand U36601 (N_36601,N_36165,N_36225);
or U36602 (N_36602,N_36438,N_36369);
and U36603 (N_36603,N_36385,N_36242);
xor U36604 (N_36604,N_36324,N_36314);
xnor U36605 (N_36605,N_36413,N_36123);
nor U36606 (N_36606,N_36249,N_36394);
and U36607 (N_36607,N_36002,N_36136);
nand U36608 (N_36608,N_36390,N_36047);
or U36609 (N_36609,N_36248,N_36347);
nand U36610 (N_36610,N_36493,N_36186);
or U36611 (N_36611,N_36241,N_36480);
or U36612 (N_36612,N_36128,N_36180);
nor U36613 (N_36613,N_36246,N_36110);
nand U36614 (N_36614,N_36071,N_36375);
and U36615 (N_36615,N_36422,N_36129);
and U36616 (N_36616,N_36153,N_36172);
xnor U36617 (N_36617,N_36138,N_36426);
or U36618 (N_36618,N_36444,N_36151);
nand U36619 (N_36619,N_36084,N_36013);
nand U36620 (N_36620,N_36088,N_36292);
nand U36621 (N_36621,N_36465,N_36485);
or U36622 (N_36622,N_36345,N_36140);
and U36623 (N_36623,N_36014,N_36384);
and U36624 (N_36624,N_36251,N_36127);
nand U36625 (N_36625,N_36183,N_36156);
or U36626 (N_36626,N_36034,N_36300);
xor U36627 (N_36627,N_36420,N_36202);
and U36628 (N_36628,N_36423,N_36118);
nor U36629 (N_36629,N_36171,N_36170);
xnor U36630 (N_36630,N_36494,N_36056);
or U36631 (N_36631,N_36448,N_36461);
nand U36632 (N_36632,N_36051,N_36289);
or U36633 (N_36633,N_36147,N_36100);
nor U36634 (N_36634,N_36373,N_36228);
xor U36635 (N_36635,N_36068,N_36041);
xnor U36636 (N_36636,N_36209,N_36178);
or U36637 (N_36637,N_36233,N_36185);
nand U36638 (N_36638,N_36213,N_36343);
nor U36639 (N_36639,N_36353,N_36222);
nand U36640 (N_36640,N_36379,N_36179);
or U36641 (N_36641,N_36139,N_36247);
nor U36642 (N_36642,N_36243,N_36256);
nand U36643 (N_36643,N_36148,N_36207);
nor U36644 (N_36644,N_36090,N_36340);
nand U36645 (N_36645,N_36094,N_36337);
nor U36646 (N_36646,N_36442,N_36308);
or U36647 (N_36647,N_36499,N_36276);
and U36648 (N_36648,N_36468,N_36363);
nand U36649 (N_36649,N_36387,N_36086);
nor U36650 (N_36650,N_36215,N_36261);
nor U36651 (N_36651,N_36408,N_36416);
or U36652 (N_36652,N_36437,N_36272);
or U36653 (N_36653,N_36145,N_36367);
or U36654 (N_36654,N_36490,N_36327);
nor U36655 (N_36655,N_36035,N_36365);
or U36656 (N_36656,N_36001,N_36358);
and U36657 (N_36657,N_36016,N_36445);
and U36658 (N_36658,N_36310,N_36045);
nand U36659 (N_36659,N_36427,N_36303);
xnor U36660 (N_36660,N_36226,N_36198);
nor U36661 (N_36661,N_36025,N_36491);
xor U36662 (N_36662,N_36023,N_36190);
and U36663 (N_36663,N_36061,N_36392);
nand U36664 (N_36664,N_36477,N_36240);
nor U36665 (N_36665,N_36119,N_36224);
nand U36666 (N_36666,N_36330,N_36092);
nor U36667 (N_36667,N_36239,N_36067);
or U36668 (N_36668,N_36130,N_36044);
and U36669 (N_36669,N_36415,N_36223);
or U36670 (N_36670,N_36169,N_36428);
xnor U36671 (N_36671,N_36273,N_36383);
xnor U36672 (N_36672,N_36009,N_36031);
xor U36673 (N_36673,N_36142,N_36033);
xnor U36674 (N_36674,N_36066,N_36264);
nor U36675 (N_36675,N_36331,N_36150);
nor U36676 (N_36676,N_36281,N_36299);
and U36677 (N_36677,N_36488,N_36201);
and U36678 (N_36678,N_36032,N_36073);
nand U36679 (N_36679,N_36450,N_36137);
nor U36680 (N_36680,N_36196,N_36435);
nor U36681 (N_36681,N_36036,N_36194);
nand U36682 (N_36682,N_36316,N_36403);
nor U36683 (N_36683,N_36166,N_36176);
and U36684 (N_36684,N_36470,N_36069);
or U36685 (N_36685,N_36102,N_36341);
nor U36686 (N_36686,N_36402,N_36329);
nor U36687 (N_36687,N_36008,N_36364);
nor U36688 (N_36688,N_36431,N_36432);
or U36689 (N_36689,N_36309,N_36374);
nor U36690 (N_36690,N_36346,N_36291);
xnor U36691 (N_36691,N_36269,N_36093);
nand U36692 (N_36692,N_36081,N_36456);
nor U36693 (N_36693,N_36360,N_36497);
and U36694 (N_36694,N_36323,N_36211);
xor U36695 (N_36695,N_36104,N_36030);
nor U36696 (N_36696,N_36164,N_36158);
and U36697 (N_36697,N_36114,N_36418);
or U36698 (N_36698,N_36290,N_36361);
nand U36699 (N_36699,N_36391,N_36482);
and U36700 (N_36700,N_36396,N_36429);
nor U36701 (N_36701,N_36479,N_36059);
and U36702 (N_36702,N_36232,N_36447);
xor U36703 (N_36703,N_36098,N_36177);
or U36704 (N_36704,N_36399,N_36259);
and U36705 (N_36705,N_36050,N_36254);
or U36706 (N_36706,N_36320,N_36054);
nand U36707 (N_36707,N_36483,N_36382);
nor U36708 (N_36708,N_36184,N_36266);
nand U36709 (N_36709,N_36381,N_36188);
xnor U36710 (N_36710,N_36275,N_36288);
xor U36711 (N_36711,N_36168,N_36149);
nor U36712 (N_36712,N_36301,N_36366);
nor U36713 (N_36713,N_36144,N_36359);
or U36714 (N_36714,N_36038,N_36409);
xnor U36715 (N_36715,N_36349,N_36335);
or U36716 (N_36716,N_36157,N_36380);
xor U36717 (N_36717,N_36007,N_36230);
xor U36718 (N_36718,N_36462,N_36368);
xnor U36719 (N_36719,N_36406,N_36495);
or U36720 (N_36720,N_36302,N_36124);
and U36721 (N_36721,N_36175,N_36283);
nand U36722 (N_36722,N_36221,N_36111);
and U36723 (N_36723,N_36163,N_36317);
or U36724 (N_36724,N_36219,N_36132);
or U36725 (N_36725,N_36372,N_36052);
nor U36726 (N_36726,N_36321,N_36370);
xor U36727 (N_36727,N_36344,N_36464);
xor U36728 (N_36728,N_36397,N_36268);
nor U36729 (N_36729,N_36306,N_36443);
and U36730 (N_36730,N_36411,N_36229);
nor U36731 (N_36731,N_36452,N_36074);
and U36732 (N_36732,N_36250,N_36455);
nor U36733 (N_36733,N_36220,N_36298);
xor U36734 (N_36734,N_36193,N_36022);
and U36735 (N_36735,N_36352,N_36167);
nand U36736 (N_36736,N_36096,N_36065);
or U36737 (N_36737,N_36006,N_36388);
nand U36738 (N_36738,N_36449,N_36484);
xor U36739 (N_36739,N_36293,N_36039);
xor U36740 (N_36740,N_36267,N_36475);
and U36741 (N_36741,N_36091,N_36079);
xor U36742 (N_36742,N_36404,N_36487);
xor U36743 (N_36743,N_36356,N_36412);
nor U36744 (N_36744,N_36398,N_36459);
nand U36745 (N_36745,N_36116,N_36064);
xor U36746 (N_36746,N_36040,N_36425);
nor U36747 (N_36747,N_36087,N_36141);
nand U36748 (N_36748,N_36126,N_36112);
xor U36749 (N_36749,N_36342,N_36439);
nor U36750 (N_36750,N_36470,N_36084);
and U36751 (N_36751,N_36103,N_36331);
nor U36752 (N_36752,N_36271,N_36475);
nand U36753 (N_36753,N_36065,N_36165);
nor U36754 (N_36754,N_36316,N_36232);
xor U36755 (N_36755,N_36219,N_36225);
xor U36756 (N_36756,N_36031,N_36348);
or U36757 (N_36757,N_36361,N_36019);
nand U36758 (N_36758,N_36445,N_36414);
nor U36759 (N_36759,N_36158,N_36233);
xor U36760 (N_36760,N_36039,N_36281);
or U36761 (N_36761,N_36365,N_36106);
and U36762 (N_36762,N_36274,N_36396);
or U36763 (N_36763,N_36292,N_36426);
nand U36764 (N_36764,N_36419,N_36095);
nor U36765 (N_36765,N_36306,N_36039);
or U36766 (N_36766,N_36412,N_36477);
and U36767 (N_36767,N_36228,N_36244);
nor U36768 (N_36768,N_36491,N_36133);
nor U36769 (N_36769,N_36305,N_36257);
and U36770 (N_36770,N_36289,N_36094);
nand U36771 (N_36771,N_36012,N_36489);
nand U36772 (N_36772,N_36495,N_36197);
nand U36773 (N_36773,N_36027,N_36254);
xor U36774 (N_36774,N_36315,N_36097);
or U36775 (N_36775,N_36273,N_36398);
nand U36776 (N_36776,N_36301,N_36189);
nor U36777 (N_36777,N_36033,N_36046);
nand U36778 (N_36778,N_36112,N_36343);
xnor U36779 (N_36779,N_36353,N_36474);
and U36780 (N_36780,N_36157,N_36365);
nand U36781 (N_36781,N_36479,N_36001);
nor U36782 (N_36782,N_36078,N_36271);
nand U36783 (N_36783,N_36185,N_36333);
xor U36784 (N_36784,N_36310,N_36419);
nor U36785 (N_36785,N_36354,N_36088);
or U36786 (N_36786,N_36417,N_36226);
nor U36787 (N_36787,N_36498,N_36382);
or U36788 (N_36788,N_36351,N_36129);
xnor U36789 (N_36789,N_36439,N_36100);
xnor U36790 (N_36790,N_36414,N_36191);
or U36791 (N_36791,N_36171,N_36463);
xor U36792 (N_36792,N_36044,N_36068);
nor U36793 (N_36793,N_36026,N_36359);
nand U36794 (N_36794,N_36214,N_36289);
and U36795 (N_36795,N_36153,N_36133);
or U36796 (N_36796,N_36121,N_36367);
nand U36797 (N_36797,N_36213,N_36397);
nor U36798 (N_36798,N_36086,N_36039);
xor U36799 (N_36799,N_36425,N_36448);
and U36800 (N_36800,N_36148,N_36257);
or U36801 (N_36801,N_36464,N_36019);
nor U36802 (N_36802,N_36402,N_36290);
xnor U36803 (N_36803,N_36101,N_36421);
and U36804 (N_36804,N_36022,N_36249);
nand U36805 (N_36805,N_36065,N_36240);
nor U36806 (N_36806,N_36324,N_36166);
or U36807 (N_36807,N_36078,N_36087);
or U36808 (N_36808,N_36324,N_36136);
and U36809 (N_36809,N_36279,N_36126);
xor U36810 (N_36810,N_36062,N_36491);
nor U36811 (N_36811,N_36172,N_36495);
or U36812 (N_36812,N_36029,N_36464);
xor U36813 (N_36813,N_36299,N_36013);
or U36814 (N_36814,N_36043,N_36310);
or U36815 (N_36815,N_36267,N_36463);
nor U36816 (N_36816,N_36151,N_36481);
or U36817 (N_36817,N_36214,N_36456);
nor U36818 (N_36818,N_36261,N_36222);
xor U36819 (N_36819,N_36058,N_36421);
and U36820 (N_36820,N_36242,N_36201);
nor U36821 (N_36821,N_36092,N_36222);
nor U36822 (N_36822,N_36162,N_36201);
or U36823 (N_36823,N_36320,N_36064);
xnor U36824 (N_36824,N_36132,N_36201);
nand U36825 (N_36825,N_36460,N_36212);
nand U36826 (N_36826,N_36109,N_36431);
xor U36827 (N_36827,N_36420,N_36282);
or U36828 (N_36828,N_36492,N_36084);
and U36829 (N_36829,N_36185,N_36136);
xnor U36830 (N_36830,N_36279,N_36034);
or U36831 (N_36831,N_36235,N_36031);
xor U36832 (N_36832,N_36403,N_36176);
nor U36833 (N_36833,N_36305,N_36190);
or U36834 (N_36834,N_36441,N_36162);
or U36835 (N_36835,N_36186,N_36371);
nand U36836 (N_36836,N_36322,N_36272);
and U36837 (N_36837,N_36265,N_36156);
nand U36838 (N_36838,N_36269,N_36221);
or U36839 (N_36839,N_36303,N_36286);
or U36840 (N_36840,N_36395,N_36255);
xor U36841 (N_36841,N_36211,N_36308);
xnor U36842 (N_36842,N_36186,N_36112);
or U36843 (N_36843,N_36419,N_36022);
or U36844 (N_36844,N_36411,N_36255);
or U36845 (N_36845,N_36085,N_36380);
nand U36846 (N_36846,N_36372,N_36351);
and U36847 (N_36847,N_36378,N_36273);
xnor U36848 (N_36848,N_36182,N_36166);
nand U36849 (N_36849,N_36213,N_36281);
or U36850 (N_36850,N_36161,N_36019);
xor U36851 (N_36851,N_36062,N_36294);
xor U36852 (N_36852,N_36024,N_36125);
and U36853 (N_36853,N_36297,N_36146);
or U36854 (N_36854,N_36233,N_36425);
xnor U36855 (N_36855,N_36043,N_36100);
and U36856 (N_36856,N_36418,N_36485);
nor U36857 (N_36857,N_36062,N_36097);
or U36858 (N_36858,N_36468,N_36427);
and U36859 (N_36859,N_36183,N_36150);
xor U36860 (N_36860,N_36457,N_36182);
nand U36861 (N_36861,N_36352,N_36488);
and U36862 (N_36862,N_36280,N_36324);
xnor U36863 (N_36863,N_36157,N_36432);
or U36864 (N_36864,N_36241,N_36471);
xor U36865 (N_36865,N_36282,N_36077);
and U36866 (N_36866,N_36399,N_36030);
xnor U36867 (N_36867,N_36372,N_36195);
or U36868 (N_36868,N_36340,N_36302);
and U36869 (N_36869,N_36121,N_36105);
xnor U36870 (N_36870,N_36005,N_36327);
and U36871 (N_36871,N_36103,N_36199);
xor U36872 (N_36872,N_36269,N_36480);
or U36873 (N_36873,N_36069,N_36111);
and U36874 (N_36874,N_36353,N_36074);
and U36875 (N_36875,N_36154,N_36396);
nand U36876 (N_36876,N_36068,N_36470);
and U36877 (N_36877,N_36456,N_36391);
nand U36878 (N_36878,N_36055,N_36390);
xor U36879 (N_36879,N_36110,N_36477);
or U36880 (N_36880,N_36139,N_36459);
or U36881 (N_36881,N_36200,N_36452);
or U36882 (N_36882,N_36479,N_36237);
xor U36883 (N_36883,N_36175,N_36059);
xnor U36884 (N_36884,N_36238,N_36372);
xnor U36885 (N_36885,N_36180,N_36131);
or U36886 (N_36886,N_36317,N_36172);
or U36887 (N_36887,N_36183,N_36284);
nor U36888 (N_36888,N_36132,N_36074);
nor U36889 (N_36889,N_36030,N_36273);
xor U36890 (N_36890,N_36267,N_36033);
xnor U36891 (N_36891,N_36071,N_36274);
xnor U36892 (N_36892,N_36239,N_36417);
or U36893 (N_36893,N_36264,N_36278);
xnor U36894 (N_36894,N_36114,N_36166);
xor U36895 (N_36895,N_36379,N_36017);
or U36896 (N_36896,N_36029,N_36241);
nor U36897 (N_36897,N_36135,N_36180);
xnor U36898 (N_36898,N_36145,N_36237);
nand U36899 (N_36899,N_36323,N_36271);
nand U36900 (N_36900,N_36117,N_36295);
xor U36901 (N_36901,N_36162,N_36231);
nand U36902 (N_36902,N_36330,N_36471);
or U36903 (N_36903,N_36191,N_36466);
nor U36904 (N_36904,N_36085,N_36347);
xnor U36905 (N_36905,N_36060,N_36110);
and U36906 (N_36906,N_36145,N_36230);
xor U36907 (N_36907,N_36447,N_36472);
nor U36908 (N_36908,N_36363,N_36465);
nand U36909 (N_36909,N_36458,N_36394);
and U36910 (N_36910,N_36447,N_36322);
xnor U36911 (N_36911,N_36033,N_36293);
or U36912 (N_36912,N_36227,N_36014);
nor U36913 (N_36913,N_36073,N_36221);
and U36914 (N_36914,N_36009,N_36318);
or U36915 (N_36915,N_36467,N_36228);
nor U36916 (N_36916,N_36226,N_36235);
xnor U36917 (N_36917,N_36213,N_36435);
and U36918 (N_36918,N_36064,N_36207);
nand U36919 (N_36919,N_36106,N_36399);
nor U36920 (N_36920,N_36266,N_36005);
nor U36921 (N_36921,N_36037,N_36028);
nor U36922 (N_36922,N_36452,N_36175);
or U36923 (N_36923,N_36155,N_36396);
and U36924 (N_36924,N_36241,N_36197);
or U36925 (N_36925,N_36321,N_36145);
nand U36926 (N_36926,N_36365,N_36303);
nor U36927 (N_36927,N_36067,N_36478);
nand U36928 (N_36928,N_36431,N_36294);
xor U36929 (N_36929,N_36055,N_36168);
and U36930 (N_36930,N_36334,N_36313);
nand U36931 (N_36931,N_36460,N_36488);
or U36932 (N_36932,N_36029,N_36112);
nand U36933 (N_36933,N_36374,N_36288);
or U36934 (N_36934,N_36059,N_36060);
and U36935 (N_36935,N_36187,N_36444);
and U36936 (N_36936,N_36140,N_36273);
nor U36937 (N_36937,N_36315,N_36159);
and U36938 (N_36938,N_36165,N_36069);
and U36939 (N_36939,N_36328,N_36499);
nand U36940 (N_36940,N_36365,N_36165);
nand U36941 (N_36941,N_36329,N_36056);
or U36942 (N_36942,N_36258,N_36257);
xor U36943 (N_36943,N_36320,N_36175);
xnor U36944 (N_36944,N_36024,N_36078);
nor U36945 (N_36945,N_36185,N_36246);
nand U36946 (N_36946,N_36291,N_36161);
nand U36947 (N_36947,N_36189,N_36429);
xnor U36948 (N_36948,N_36379,N_36370);
and U36949 (N_36949,N_36224,N_36188);
xnor U36950 (N_36950,N_36073,N_36351);
nand U36951 (N_36951,N_36303,N_36426);
or U36952 (N_36952,N_36006,N_36437);
or U36953 (N_36953,N_36101,N_36118);
or U36954 (N_36954,N_36134,N_36391);
nand U36955 (N_36955,N_36440,N_36406);
nor U36956 (N_36956,N_36195,N_36384);
xnor U36957 (N_36957,N_36273,N_36040);
and U36958 (N_36958,N_36201,N_36204);
xnor U36959 (N_36959,N_36279,N_36256);
xnor U36960 (N_36960,N_36251,N_36030);
nor U36961 (N_36961,N_36096,N_36215);
nor U36962 (N_36962,N_36083,N_36303);
nor U36963 (N_36963,N_36108,N_36347);
xnor U36964 (N_36964,N_36327,N_36359);
and U36965 (N_36965,N_36084,N_36160);
nand U36966 (N_36966,N_36090,N_36101);
or U36967 (N_36967,N_36292,N_36224);
xor U36968 (N_36968,N_36283,N_36275);
nand U36969 (N_36969,N_36096,N_36418);
and U36970 (N_36970,N_36075,N_36370);
or U36971 (N_36971,N_36185,N_36224);
xor U36972 (N_36972,N_36363,N_36117);
nor U36973 (N_36973,N_36485,N_36232);
nand U36974 (N_36974,N_36106,N_36104);
and U36975 (N_36975,N_36104,N_36374);
and U36976 (N_36976,N_36132,N_36003);
and U36977 (N_36977,N_36441,N_36187);
xor U36978 (N_36978,N_36356,N_36424);
or U36979 (N_36979,N_36125,N_36149);
nand U36980 (N_36980,N_36105,N_36064);
nand U36981 (N_36981,N_36165,N_36242);
or U36982 (N_36982,N_36435,N_36296);
nand U36983 (N_36983,N_36127,N_36401);
nand U36984 (N_36984,N_36205,N_36260);
nor U36985 (N_36985,N_36413,N_36498);
xor U36986 (N_36986,N_36283,N_36263);
xor U36987 (N_36987,N_36311,N_36035);
or U36988 (N_36988,N_36216,N_36427);
or U36989 (N_36989,N_36279,N_36107);
nor U36990 (N_36990,N_36258,N_36218);
and U36991 (N_36991,N_36305,N_36081);
xnor U36992 (N_36992,N_36073,N_36141);
or U36993 (N_36993,N_36199,N_36105);
nor U36994 (N_36994,N_36434,N_36318);
or U36995 (N_36995,N_36282,N_36424);
or U36996 (N_36996,N_36305,N_36064);
nor U36997 (N_36997,N_36218,N_36487);
xor U36998 (N_36998,N_36305,N_36037);
xnor U36999 (N_36999,N_36187,N_36213);
nor U37000 (N_37000,N_36783,N_36623);
xnor U37001 (N_37001,N_36670,N_36822);
nor U37002 (N_37002,N_36744,N_36504);
or U37003 (N_37003,N_36694,N_36799);
nor U37004 (N_37004,N_36802,N_36530);
nand U37005 (N_37005,N_36642,N_36551);
nand U37006 (N_37006,N_36829,N_36650);
xor U37007 (N_37007,N_36858,N_36658);
nand U37008 (N_37008,N_36663,N_36500);
xnor U37009 (N_37009,N_36748,N_36685);
nor U37010 (N_37010,N_36548,N_36973);
nor U37011 (N_37011,N_36654,N_36794);
and U37012 (N_37012,N_36765,N_36553);
nand U37013 (N_37013,N_36933,N_36746);
nor U37014 (N_37014,N_36714,N_36993);
nand U37015 (N_37015,N_36664,N_36651);
nor U37016 (N_37016,N_36624,N_36760);
and U37017 (N_37017,N_36903,N_36560);
or U37018 (N_37018,N_36841,N_36740);
or U37019 (N_37019,N_36676,N_36606);
or U37020 (N_37020,N_36649,N_36696);
nand U37021 (N_37021,N_36784,N_36666);
nor U37022 (N_37022,N_36808,N_36835);
nor U37023 (N_37023,N_36597,N_36859);
nand U37024 (N_37024,N_36743,N_36704);
or U37025 (N_37025,N_36892,N_36894);
nor U37026 (N_37026,N_36758,N_36752);
nand U37027 (N_37027,N_36939,N_36628);
nor U37028 (N_37028,N_36620,N_36819);
xor U37029 (N_37029,N_36821,N_36526);
or U37030 (N_37030,N_36779,N_36812);
nand U37031 (N_37031,N_36803,N_36713);
nand U37032 (N_37032,N_36898,N_36976);
or U37033 (N_37033,N_36766,N_36961);
and U37034 (N_37034,N_36964,N_36817);
or U37035 (N_37035,N_36706,N_36691);
nand U37036 (N_37036,N_36680,N_36907);
xnor U37037 (N_37037,N_36512,N_36615);
nor U37038 (N_37038,N_36791,N_36667);
or U37039 (N_37039,N_36991,N_36850);
xor U37040 (N_37040,N_36879,N_36724);
nor U37041 (N_37041,N_36816,N_36878);
nor U37042 (N_37042,N_36872,N_36904);
xnor U37043 (N_37043,N_36517,N_36775);
nand U37044 (N_37044,N_36644,N_36999);
and U37045 (N_37045,N_36736,N_36842);
nor U37046 (N_37046,N_36622,N_36897);
nor U37047 (N_37047,N_36837,N_36936);
and U37048 (N_37048,N_36908,N_36870);
nand U37049 (N_37049,N_36956,N_36574);
and U37050 (N_37050,N_36727,N_36967);
and U37051 (N_37051,N_36506,N_36739);
and U37052 (N_37052,N_36928,N_36601);
xor U37053 (N_37053,N_36968,N_36987);
nor U37054 (N_37054,N_36954,N_36661);
nand U37055 (N_37055,N_36519,N_36798);
and U37056 (N_37056,N_36565,N_36756);
nand U37057 (N_37057,N_36877,N_36679);
or U37058 (N_37058,N_36825,N_36625);
and U37059 (N_37059,N_36689,N_36762);
nand U37060 (N_37060,N_36545,N_36922);
nor U37061 (N_37061,N_36638,N_36722);
nor U37062 (N_37062,N_36533,N_36735);
and U37063 (N_37063,N_36693,N_36719);
or U37064 (N_37064,N_36721,N_36801);
nor U37065 (N_37065,N_36789,N_36909);
xor U37066 (N_37066,N_36866,N_36600);
and U37067 (N_37067,N_36602,N_36945);
nand U37068 (N_37068,N_36927,N_36848);
and U37069 (N_37069,N_36709,N_36668);
and U37070 (N_37070,N_36838,N_36675);
and U37071 (N_37071,N_36505,N_36930);
nor U37072 (N_37072,N_36828,N_36959);
and U37073 (N_37073,N_36516,N_36585);
and U37074 (N_37074,N_36809,N_36570);
xor U37075 (N_37075,N_36528,N_36645);
nand U37076 (N_37076,N_36787,N_36546);
xnor U37077 (N_37077,N_36906,N_36705);
or U37078 (N_37078,N_36941,N_36750);
nand U37079 (N_37079,N_36647,N_36678);
and U37080 (N_37080,N_36896,N_36582);
xnor U37081 (N_37081,N_36648,N_36734);
nor U37082 (N_37082,N_36621,N_36699);
nor U37083 (N_37083,N_36926,N_36915);
or U37084 (N_37084,N_36711,N_36981);
or U37085 (N_37085,N_36852,N_36772);
nor U37086 (N_37086,N_36700,N_36770);
or U37087 (N_37087,N_36525,N_36588);
nand U37088 (N_37088,N_36882,N_36938);
and U37089 (N_37089,N_36832,N_36531);
nand U37090 (N_37090,N_36815,N_36916);
and U37091 (N_37091,N_36830,N_36539);
xnor U37092 (N_37092,N_36738,N_36501);
nand U37093 (N_37093,N_36745,N_36535);
or U37094 (N_37094,N_36509,N_36918);
and U37095 (N_37095,N_36611,N_36807);
nor U37096 (N_37096,N_36614,N_36590);
nor U37097 (N_37097,N_36749,N_36782);
nand U37098 (N_37098,N_36952,N_36890);
nand U37099 (N_37099,N_36834,N_36855);
nand U37100 (N_37100,N_36559,N_36811);
or U37101 (N_37101,N_36681,N_36598);
and U37102 (N_37102,N_36912,N_36786);
nand U37103 (N_37103,N_36547,N_36527);
xor U37104 (N_37104,N_36901,N_36864);
and U37105 (N_37105,N_36989,N_36780);
and U37106 (N_37106,N_36845,N_36684);
nand U37107 (N_37107,N_36975,N_36979);
and U37108 (N_37108,N_36751,N_36990);
xor U37109 (N_37109,N_36919,N_36594);
nand U37110 (N_37110,N_36905,N_36960);
nand U37111 (N_37111,N_36708,N_36637);
or U37112 (N_37112,N_36683,N_36659);
xnor U37113 (N_37113,N_36576,N_36994);
or U37114 (N_37114,N_36558,N_36702);
xor U37115 (N_37115,N_36963,N_36677);
nand U37116 (N_37116,N_36520,N_36716);
or U37117 (N_37117,N_36703,N_36549);
and U37118 (N_37118,N_36513,N_36853);
nor U37119 (N_37119,N_36865,N_36537);
or U37120 (N_37120,N_36595,N_36523);
xor U37121 (N_37121,N_36715,N_36730);
nor U37122 (N_37122,N_36998,N_36910);
nor U37123 (N_37123,N_36885,N_36793);
nor U37124 (N_37124,N_36717,N_36640);
and U37125 (N_37125,N_36764,N_36902);
or U37126 (N_37126,N_36969,N_36682);
nor U37127 (N_37127,N_36965,N_36889);
nand U37128 (N_37128,N_36995,N_36688);
nand U37129 (N_37129,N_36771,N_36507);
or U37130 (N_37130,N_36543,N_36583);
and U37131 (N_37131,N_36951,N_36591);
xnor U37132 (N_37132,N_36725,N_36788);
and U37133 (N_37133,N_36985,N_36592);
or U37134 (N_37134,N_36753,N_36626);
and U37135 (N_37135,N_36818,N_36660);
nand U37136 (N_37136,N_36851,N_36880);
xor U37137 (N_37137,N_36564,N_36757);
nor U37138 (N_37138,N_36742,N_36871);
nor U37139 (N_37139,N_36631,N_36921);
or U37140 (N_37140,N_36502,N_36982);
xor U37141 (N_37141,N_36643,N_36729);
or U37142 (N_37142,N_36737,N_36728);
xor U37143 (N_37143,N_36632,N_36712);
and U37144 (N_37144,N_36781,N_36607);
xnor U37145 (N_37145,N_36687,N_36934);
and U37146 (N_37146,N_36813,N_36862);
and U37147 (N_37147,N_36785,N_36810);
nand U37148 (N_37148,N_36718,N_36731);
or U37149 (N_37149,N_36804,N_36863);
nand U37150 (N_37150,N_36575,N_36867);
nor U37151 (N_37151,N_36795,N_36581);
nor U37152 (N_37152,N_36827,N_36972);
and U37153 (N_37153,N_36697,N_36920);
xnor U37154 (N_37154,N_36673,N_36943);
nand U37155 (N_37155,N_36536,N_36833);
or U37156 (N_37156,N_36980,N_36511);
or U37157 (N_37157,N_36763,N_36883);
nor U37158 (N_37158,N_36733,N_36541);
and U37159 (N_37159,N_36847,N_36978);
xor U37160 (N_37160,N_36630,N_36657);
or U37161 (N_37161,N_36875,N_36768);
xnor U37162 (N_37162,N_36792,N_36773);
or U37163 (N_37163,N_36844,N_36970);
or U37164 (N_37164,N_36568,N_36924);
or U37165 (N_37165,N_36633,N_36698);
xor U37166 (N_37166,N_36911,N_36937);
nand U37167 (N_37167,N_36997,N_36947);
xor U37168 (N_37168,N_36988,N_36518);
or U37169 (N_37169,N_36655,N_36949);
nor U37170 (N_37170,N_36653,N_36707);
or U37171 (N_37171,N_36514,N_36613);
or U37172 (N_37172,N_36935,N_36586);
and U37173 (N_37173,N_36710,N_36610);
and U37174 (N_37174,N_36669,N_36836);
nand U37175 (N_37175,N_36895,N_36604);
xnor U37176 (N_37176,N_36508,N_36522);
nand U37177 (N_37177,N_36652,N_36876);
nor U37178 (N_37178,N_36831,N_36596);
xnor U37179 (N_37179,N_36942,N_36857);
or U37180 (N_37180,N_36977,N_36843);
or U37181 (N_37181,N_36948,N_36776);
nor U37182 (N_37182,N_36955,N_36913);
xor U37183 (N_37183,N_36550,N_36665);
nor U37184 (N_37184,N_36566,N_36887);
nor U37185 (N_37185,N_36608,N_36805);
xnor U37186 (N_37186,N_36777,N_36953);
or U37187 (N_37187,N_36720,N_36839);
nor U37188 (N_37188,N_36940,N_36577);
nor U37189 (N_37189,N_36755,N_36524);
xor U37190 (N_37190,N_36567,N_36619);
nor U37191 (N_37191,N_36754,N_36603);
nor U37192 (N_37192,N_36983,N_36886);
nor U37193 (N_37193,N_36569,N_36534);
and U37194 (N_37194,N_36899,N_36846);
nand U37195 (N_37195,N_36767,N_36557);
nor U37196 (N_37196,N_36891,N_36609);
or U37197 (N_37197,N_36695,N_36860);
nand U37198 (N_37198,N_36823,N_36634);
or U37199 (N_37199,N_36931,N_36554);
and U37200 (N_37200,N_36820,N_36900);
nand U37201 (N_37201,N_36540,N_36572);
nor U37202 (N_37202,N_36556,N_36605);
and U37203 (N_37203,N_36573,N_36946);
xor U37204 (N_37204,N_36814,N_36962);
nor U37205 (N_37205,N_36996,N_36555);
nand U37206 (N_37206,N_36761,N_36701);
and U37207 (N_37207,N_36984,N_36587);
and U37208 (N_37208,N_36690,N_36542);
and U37209 (N_37209,N_36723,N_36790);
nor U37210 (N_37210,N_36616,N_36593);
nand U37211 (N_37211,N_36974,N_36639);
nand U37212 (N_37212,N_36824,N_36503);
xnor U37213 (N_37213,N_36726,N_36579);
nand U37214 (N_37214,N_36923,N_36914);
xor U37215 (N_37215,N_36800,N_36646);
nor U37216 (N_37216,N_36774,N_36874);
nand U37217 (N_37217,N_36884,N_36563);
and U37218 (N_37218,N_36641,N_36769);
and U37219 (N_37219,N_36747,N_36856);
or U37220 (N_37220,N_36966,N_36741);
and U37221 (N_37221,N_36635,N_36562);
nand U37222 (N_37222,N_36932,N_36636);
nor U37223 (N_37223,N_36840,N_36854);
and U37224 (N_37224,N_36629,N_36552);
nor U37225 (N_37225,N_36797,N_36950);
nor U37226 (N_37226,N_36662,N_36580);
xor U37227 (N_37227,N_36612,N_36671);
or U37228 (N_37228,N_36599,N_36849);
or U37229 (N_37229,N_36627,N_36617);
xor U37230 (N_37230,N_36861,N_36971);
nor U37231 (N_37231,N_36868,N_36618);
nand U37232 (N_37232,N_36826,N_36515);
nand U37233 (N_37233,N_36917,N_36888);
nand U37234 (N_37234,N_36584,N_36925);
nor U37235 (N_37235,N_36686,N_36571);
and U37236 (N_37236,N_36778,N_36521);
xnor U37237 (N_37237,N_36692,N_36561);
nand U37238 (N_37238,N_36589,N_36893);
nand U37239 (N_37239,N_36869,N_36958);
and U37240 (N_37240,N_36986,N_36957);
nor U37241 (N_37241,N_36578,N_36944);
nor U37242 (N_37242,N_36929,N_36674);
and U37243 (N_37243,N_36873,N_36732);
nor U37244 (N_37244,N_36796,N_36532);
nor U37245 (N_37245,N_36806,N_36759);
or U37246 (N_37246,N_36672,N_36544);
or U37247 (N_37247,N_36510,N_36881);
and U37248 (N_37248,N_36992,N_36538);
or U37249 (N_37249,N_36529,N_36656);
nor U37250 (N_37250,N_36644,N_36983);
and U37251 (N_37251,N_36915,N_36966);
xor U37252 (N_37252,N_36980,N_36576);
or U37253 (N_37253,N_36722,N_36523);
or U37254 (N_37254,N_36874,N_36887);
and U37255 (N_37255,N_36529,N_36701);
xnor U37256 (N_37256,N_36793,N_36606);
nor U37257 (N_37257,N_36958,N_36792);
and U37258 (N_37258,N_36675,N_36659);
nand U37259 (N_37259,N_36784,N_36906);
or U37260 (N_37260,N_36553,N_36999);
or U37261 (N_37261,N_36561,N_36773);
or U37262 (N_37262,N_36640,N_36669);
or U37263 (N_37263,N_36752,N_36692);
or U37264 (N_37264,N_36610,N_36883);
xnor U37265 (N_37265,N_36985,N_36925);
or U37266 (N_37266,N_36558,N_36827);
xnor U37267 (N_37267,N_36951,N_36542);
nor U37268 (N_37268,N_36605,N_36773);
xor U37269 (N_37269,N_36685,N_36725);
nor U37270 (N_37270,N_36505,N_36676);
nor U37271 (N_37271,N_36906,N_36795);
nor U37272 (N_37272,N_36671,N_36740);
xnor U37273 (N_37273,N_36621,N_36595);
nand U37274 (N_37274,N_36775,N_36840);
nor U37275 (N_37275,N_36734,N_36544);
xor U37276 (N_37276,N_36904,N_36893);
nand U37277 (N_37277,N_36976,N_36733);
and U37278 (N_37278,N_36960,N_36569);
xor U37279 (N_37279,N_36685,N_36691);
xnor U37280 (N_37280,N_36817,N_36560);
nor U37281 (N_37281,N_36848,N_36668);
and U37282 (N_37282,N_36898,N_36721);
nand U37283 (N_37283,N_36738,N_36685);
xnor U37284 (N_37284,N_36677,N_36885);
nor U37285 (N_37285,N_36598,N_36529);
xnor U37286 (N_37286,N_36602,N_36756);
nor U37287 (N_37287,N_36779,N_36985);
and U37288 (N_37288,N_36927,N_36978);
nor U37289 (N_37289,N_36814,N_36808);
and U37290 (N_37290,N_36716,N_36978);
or U37291 (N_37291,N_36707,N_36987);
and U37292 (N_37292,N_36828,N_36569);
and U37293 (N_37293,N_36820,N_36809);
nor U37294 (N_37294,N_36779,N_36548);
nor U37295 (N_37295,N_36921,N_36649);
xor U37296 (N_37296,N_36923,N_36624);
nand U37297 (N_37297,N_36957,N_36930);
xnor U37298 (N_37298,N_36920,N_36908);
nor U37299 (N_37299,N_36698,N_36613);
and U37300 (N_37300,N_36649,N_36905);
nand U37301 (N_37301,N_36623,N_36634);
and U37302 (N_37302,N_36593,N_36559);
and U37303 (N_37303,N_36908,N_36970);
nand U37304 (N_37304,N_36564,N_36848);
or U37305 (N_37305,N_36866,N_36686);
xor U37306 (N_37306,N_36695,N_36827);
and U37307 (N_37307,N_36647,N_36812);
xor U37308 (N_37308,N_36584,N_36714);
or U37309 (N_37309,N_36923,N_36900);
nor U37310 (N_37310,N_36827,N_36867);
nor U37311 (N_37311,N_36874,N_36744);
nor U37312 (N_37312,N_36697,N_36527);
xnor U37313 (N_37313,N_36977,N_36765);
nor U37314 (N_37314,N_36761,N_36743);
xnor U37315 (N_37315,N_36905,N_36846);
nor U37316 (N_37316,N_36923,N_36657);
or U37317 (N_37317,N_36965,N_36941);
and U37318 (N_37318,N_36632,N_36792);
or U37319 (N_37319,N_36613,N_36648);
nand U37320 (N_37320,N_36945,N_36696);
nor U37321 (N_37321,N_36629,N_36852);
or U37322 (N_37322,N_36514,N_36857);
nor U37323 (N_37323,N_36504,N_36627);
xor U37324 (N_37324,N_36875,N_36989);
and U37325 (N_37325,N_36803,N_36898);
nor U37326 (N_37326,N_36521,N_36556);
or U37327 (N_37327,N_36804,N_36868);
nor U37328 (N_37328,N_36982,N_36753);
xnor U37329 (N_37329,N_36914,N_36576);
and U37330 (N_37330,N_36768,N_36977);
nand U37331 (N_37331,N_36541,N_36518);
nor U37332 (N_37332,N_36854,N_36620);
or U37333 (N_37333,N_36752,N_36532);
or U37334 (N_37334,N_36774,N_36625);
nor U37335 (N_37335,N_36878,N_36546);
nand U37336 (N_37336,N_36767,N_36519);
or U37337 (N_37337,N_36576,N_36653);
and U37338 (N_37338,N_36853,N_36820);
nor U37339 (N_37339,N_36805,N_36865);
nand U37340 (N_37340,N_36939,N_36814);
nand U37341 (N_37341,N_36784,N_36915);
nor U37342 (N_37342,N_36934,N_36583);
or U37343 (N_37343,N_36777,N_36547);
nand U37344 (N_37344,N_36957,N_36610);
nand U37345 (N_37345,N_36601,N_36857);
xnor U37346 (N_37346,N_36761,N_36546);
nand U37347 (N_37347,N_36604,N_36743);
xnor U37348 (N_37348,N_36808,N_36575);
xor U37349 (N_37349,N_36647,N_36602);
and U37350 (N_37350,N_36794,N_36622);
xnor U37351 (N_37351,N_36717,N_36786);
nor U37352 (N_37352,N_36825,N_36506);
nand U37353 (N_37353,N_36789,N_36764);
nand U37354 (N_37354,N_36519,N_36788);
or U37355 (N_37355,N_36513,N_36772);
nor U37356 (N_37356,N_36769,N_36692);
xnor U37357 (N_37357,N_36953,N_36827);
nor U37358 (N_37358,N_36936,N_36974);
nand U37359 (N_37359,N_36946,N_36529);
and U37360 (N_37360,N_36563,N_36622);
or U37361 (N_37361,N_36990,N_36764);
nand U37362 (N_37362,N_36545,N_36742);
xnor U37363 (N_37363,N_36674,N_36707);
and U37364 (N_37364,N_36653,N_36638);
nor U37365 (N_37365,N_36540,N_36985);
xnor U37366 (N_37366,N_36551,N_36750);
nand U37367 (N_37367,N_36857,N_36627);
or U37368 (N_37368,N_36929,N_36849);
xor U37369 (N_37369,N_36822,N_36918);
and U37370 (N_37370,N_36687,N_36850);
and U37371 (N_37371,N_36899,N_36940);
nor U37372 (N_37372,N_36766,N_36555);
or U37373 (N_37373,N_36761,N_36776);
nand U37374 (N_37374,N_36555,N_36979);
xor U37375 (N_37375,N_36947,N_36624);
nor U37376 (N_37376,N_36613,N_36840);
nand U37377 (N_37377,N_36692,N_36530);
xnor U37378 (N_37378,N_36638,N_36831);
nand U37379 (N_37379,N_36685,N_36838);
nand U37380 (N_37380,N_36778,N_36838);
or U37381 (N_37381,N_36974,N_36645);
nand U37382 (N_37382,N_36710,N_36832);
or U37383 (N_37383,N_36840,N_36895);
xnor U37384 (N_37384,N_36582,N_36650);
nor U37385 (N_37385,N_36897,N_36844);
and U37386 (N_37386,N_36670,N_36957);
nor U37387 (N_37387,N_36751,N_36899);
xnor U37388 (N_37388,N_36955,N_36967);
nand U37389 (N_37389,N_36721,N_36749);
or U37390 (N_37390,N_36541,N_36727);
and U37391 (N_37391,N_36766,N_36739);
xor U37392 (N_37392,N_36565,N_36672);
nor U37393 (N_37393,N_36528,N_36705);
nor U37394 (N_37394,N_36981,N_36902);
or U37395 (N_37395,N_36649,N_36999);
and U37396 (N_37396,N_36926,N_36957);
xor U37397 (N_37397,N_36946,N_36647);
nor U37398 (N_37398,N_36508,N_36775);
nand U37399 (N_37399,N_36875,N_36991);
nand U37400 (N_37400,N_36966,N_36563);
xnor U37401 (N_37401,N_36767,N_36534);
xor U37402 (N_37402,N_36796,N_36943);
nand U37403 (N_37403,N_36568,N_36929);
or U37404 (N_37404,N_36976,N_36528);
xor U37405 (N_37405,N_36951,N_36911);
xor U37406 (N_37406,N_36502,N_36707);
and U37407 (N_37407,N_36504,N_36512);
nor U37408 (N_37408,N_36718,N_36639);
and U37409 (N_37409,N_36731,N_36958);
xnor U37410 (N_37410,N_36576,N_36668);
xor U37411 (N_37411,N_36622,N_36667);
nor U37412 (N_37412,N_36506,N_36683);
nand U37413 (N_37413,N_36803,N_36815);
or U37414 (N_37414,N_36628,N_36933);
xor U37415 (N_37415,N_36538,N_36745);
and U37416 (N_37416,N_36569,N_36613);
or U37417 (N_37417,N_36989,N_36960);
and U37418 (N_37418,N_36825,N_36615);
nand U37419 (N_37419,N_36709,N_36653);
nor U37420 (N_37420,N_36760,N_36596);
nand U37421 (N_37421,N_36797,N_36622);
or U37422 (N_37422,N_36888,N_36523);
nand U37423 (N_37423,N_36639,N_36992);
and U37424 (N_37424,N_36596,N_36819);
nor U37425 (N_37425,N_36693,N_36868);
or U37426 (N_37426,N_36752,N_36647);
nand U37427 (N_37427,N_36896,N_36863);
nor U37428 (N_37428,N_36900,N_36951);
nand U37429 (N_37429,N_36775,N_36969);
xnor U37430 (N_37430,N_36608,N_36638);
and U37431 (N_37431,N_36603,N_36779);
or U37432 (N_37432,N_36863,N_36607);
or U37433 (N_37433,N_36903,N_36548);
nor U37434 (N_37434,N_36575,N_36703);
nand U37435 (N_37435,N_36811,N_36703);
and U37436 (N_37436,N_36749,N_36909);
nand U37437 (N_37437,N_36625,N_36781);
nand U37438 (N_37438,N_36598,N_36829);
nor U37439 (N_37439,N_36877,N_36736);
and U37440 (N_37440,N_36769,N_36673);
nand U37441 (N_37441,N_36519,N_36502);
nand U37442 (N_37442,N_36778,N_36705);
xnor U37443 (N_37443,N_36807,N_36508);
xor U37444 (N_37444,N_36985,N_36922);
or U37445 (N_37445,N_36629,N_36521);
nand U37446 (N_37446,N_36990,N_36962);
nand U37447 (N_37447,N_36967,N_36609);
nand U37448 (N_37448,N_36865,N_36765);
xor U37449 (N_37449,N_36701,N_36979);
and U37450 (N_37450,N_36783,N_36932);
nor U37451 (N_37451,N_36892,N_36879);
nand U37452 (N_37452,N_36979,N_36583);
nor U37453 (N_37453,N_36924,N_36521);
and U37454 (N_37454,N_36692,N_36528);
and U37455 (N_37455,N_36687,N_36924);
nor U37456 (N_37456,N_36745,N_36966);
xor U37457 (N_37457,N_36875,N_36911);
xnor U37458 (N_37458,N_36543,N_36520);
nand U37459 (N_37459,N_36759,N_36833);
and U37460 (N_37460,N_36741,N_36792);
nor U37461 (N_37461,N_36574,N_36820);
and U37462 (N_37462,N_36559,N_36581);
xnor U37463 (N_37463,N_36814,N_36662);
or U37464 (N_37464,N_36987,N_36509);
or U37465 (N_37465,N_36889,N_36860);
nor U37466 (N_37466,N_36545,N_36586);
nand U37467 (N_37467,N_36969,N_36638);
nor U37468 (N_37468,N_36735,N_36540);
and U37469 (N_37469,N_36548,N_36526);
nor U37470 (N_37470,N_36917,N_36501);
and U37471 (N_37471,N_36526,N_36641);
xnor U37472 (N_37472,N_36572,N_36897);
or U37473 (N_37473,N_36950,N_36927);
and U37474 (N_37474,N_36548,N_36758);
xor U37475 (N_37475,N_36620,N_36617);
or U37476 (N_37476,N_36530,N_36721);
nor U37477 (N_37477,N_36832,N_36702);
and U37478 (N_37478,N_36939,N_36786);
or U37479 (N_37479,N_36516,N_36683);
and U37480 (N_37480,N_36878,N_36885);
xor U37481 (N_37481,N_36501,N_36594);
nor U37482 (N_37482,N_36775,N_36987);
or U37483 (N_37483,N_36584,N_36842);
or U37484 (N_37484,N_36891,N_36588);
nand U37485 (N_37485,N_36913,N_36954);
xnor U37486 (N_37486,N_36778,N_36815);
nor U37487 (N_37487,N_36659,N_36604);
nor U37488 (N_37488,N_36744,N_36640);
xor U37489 (N_37489,N_36502,N_36816);
nor U37490 (N_37490,N_36657,N_36548);
or U37491 (N_37491,N_36722,N_36945);
or U37492 (N_37492,N_36966,N_36747);
or U37493 (N_37493,N_36750,N_36971);
or U37494 (N_37494,N_36636,N_36868);
xnor U37495 (N_37495,N_36739,N_36897);
xnor U37496 (N_37496,N_36569,N_36683);
nand U37497 (N_37497,N_36831,N_36609);
nand U37498 (N_37498,N_36792,N_36533);
xnor U37499 (N_37499,N_36589,N_36536);
or U37500 (N_37500,N_37257,N_37285);
or U37501 (N_37501,N_37065,N_37218);
nand U37502 (N_37502,N_37015,N_37389);
nor U37503 (N_37503,N_37379,N_37106);
or U37504 (N_37504,N_37442,N_37225);
and U37505 (N_37505,N_37358,N_37027);
nand U37506 (N_37506,N_37055,N_37247);
nor U37507 (N_37507,N_37166,N_37046);
nor U37508 (N_37508,N_37264,N_37428);
nor U37509 (N_37509,N_37460,N_37110);
nor U37510 (N_37510,N_37012,N_37359);
or U37511 (N_37511,N_37413,N_37215);
and U37512 (N_37512,N_37439,N_37382);
nor U37513 (N_37513,N_37350,N_37420);
nor U37514 (N_37514,N_37151,N_37498);
nor U37515 (N_37515,N_37083,N_37422);
and U37516 (N_37516,N_37292,N_37430);
nand U37517 (N_37517,N_37071,N_37037);
nor U37518 (N_37518,N_37353,N_37066);
xnor U37519 (N_37519,N_37217,N_37371);
and U37520 (N_37520,N_37143,N_37079);
and U37521 (N_37521,N_37078,N_37149);
and U37522 (N_37522,N_37458,N_37276);
and U37523 (N_37523,N_37459,N_37440);
nand U37524 (N_37524,N_37323,N_37213);
xor U37525 (N_37525,N_37049,N_37118);
or U37526 (N_37526,N_37408,N_37111);
nor U37527 (N_37527,N_37416,N_37096);
nand U37528 (N_37528,N_37004,N_37122);
or U37529 (N_37529,N_37080,N_37329);
nand U37530 (N_37530,N_37465,N_37219);
xnor U37531 (N_37531,N_37008,N_37221);
nand U37532 (N_37532,N_37053,N_37333);
or U37533 (N_37533,N_37157,N_37284);
nor U37534 (N_37534,N_37128,N_37487);
nor U37535 (N_37535,N_37330,N_37355);
nor U37536 (N_37536,N_37261,N_37423);
or U37537 (N_37537,N_37373,N_37170);
nor U37538 (N_37538,N_37271,N_37057);
nor U37539 (N_37539,N_37473,N_37274);
nor U37540 (N_37540,N_37448,N_37287);
nor U37541 (N_37541,N_37165,N_37265);
and U37542 (N_37542,N_37259,N_37002);
xor U37543 (N_37543,N_37331,N_37208);
nand U37544 (N_37544,N_37435,N_37246);
nand U37545 (N_37545,N_37385,N_37212);
xor U37546 (N_37546,N_37061,N_37025);
or U37547 (N_37547,N_37150,N_37456);
nand U37548 (N_37548,N_37005,N_37467);
xor U37549 (N_37549,N_37494,N_37245);
nor U37550 (N_37550,N_37437,N_37471);
and U37551 (N_37551,N_37202,N_37235);
or U37552 (N_37552,N_37132,N_37103);
nand U37553 (N_37553,N_37200,N_37068);
and U37554 (N_37554,N_37444,N_37431);
nor U37555 (N_37555,N_37306,N_37196);
and U37556 (N_37556,N_37238,N_37023);
nor U37557 (N_37557,N_37433,N_37039);
or U37558 (N_37558,N_37030,N_37268);
and U37559 (N_37559,N_37227,N_37364);
nand U37560 (N_37560,N_37045,N_37484);
nor U37561 (N_37561,N_37229,N_37336);
xor U37562 (N_37562,N_37088,N_37014);
nand U37563 (N_37563,N_37480,N_37470);
xnor U37564 (N_37564,N_37197,N_37130);
or U37565 (N_37565,N_37137,N_37022);
nor U37566 (N_37566,N_37171,N_37239);
xor U37567 (N_37567,N_37376,N_37499);
or U37568 (N_37568,N_37497,N_37328);
or U37569 (N_37569,N_37119,N_37206);
or U37570 (N_37570,N_37266,N_37293);
nor U37571 (N_37571,N_37421,N_37135);
and U37572 (N_37572,N_37181,N_37131);
nand U37573 (N_37573,N_37378,N_37192);
or U37574 (N_37574,N_37154,N_37018);
xnor U37575 (N_37575,N_37267,N_37064);
nor U37576 (N_37576,N_37094,N_37205);
and U37577 (N_37577,N_37496,N_37273);
nand U37578 (N_37578,N_37492,N_37199);
nor U37579 (N_37579,N_37003,N_37256);
or U37580 (N_37580,N_37072,N_37436);
nor U37581 (N_37581,N_37427,N_37400);
nor U37582 (N_37582,N_37322,N_37134);
nand U37583 (N_37583,N_37425,N_37429);
or U37584 (N_37584,N_37317,N_37334);
or U37585 (N_37585,N_37097,N_37186);
nor U37586 (N_37586,N_37320,N_37013);
and U37587 (N_37587,N_37146,N_37370);
and U37588 (N_37588,N_37249,N_37415);
and U37589 (N_37589,N_37188,N_37391);
xor U37590 (N_37590,N_37356,N_37193);
xor U37591 (N_37591,N_37207,N_37381);
and U37592 (N_37592,N_37228,N_37033);
or U37593 (N_37593,N_37093,N_37189);
nand U37594 (N_37594,N_37384,N_37307);
xnor U37595 (N_37595,N_37269,N_37432);
nor U37596 (N_37596,N_37403,N_37315);
and U37597 (N_37597,N_37383,N_37401);
and U37598 (N_37598,N_37301,N_37407);
and U37599 (N_37599,N_37342,N_37153);
nand U37600 (N_37600,N_37295,N_37234);
nor U37601 (N_37601,N_37214,N_37100);
nor U37602 (N_37602,N_37184,N_37062);
or U37603 (N_37603,N_37481,N_37105);
nor U37604 (N_37604,N_37424,N_37489);
or U37605 (N_37605,N_37127,N_37253);
xnor U37606 (N_37606,N_37280,N_37028);
and U37607 (N_37607,N_37325,N_37191);
xor U37608 (N_37608,N_37445,N_37449);
xor U37609 (N_37609,N_37164,N_37176);
or U37610 (N_37610,N_37405,N_37337);
or U37611 (N_37611,N_37126,N_37162);
nand U37612 (N_37612,N_37161,N_37495);
nor U37613 (N_37613,N_37201,N_37412);
nand U37614 (N_37614,N_37308,N_37124);
xor U37615 (N_37615,N_37224,N_37374);
and U37616 (N_37616,N_37419,N_37446);
nand U37617 (N_37617,N_37402,N_37275);
nand U37618 (N_37618,N_37279,N_37115);
and U37619 (N_37619,N_37313,N_37380);
xnor U37620 (N_37620,N_37177,N_37011);
nand U37621 (N_37621,N_37318,N_37410);
or U37622 (N_37622,N_37411,N_37038);
nor U37623 (N_37623,N_37372,N_37314);
nand U37624 (N_37624,N_37145,N_37368);
and U37625 (N_37625,N_37147,N_37406);
nor U37626 (N_37626,N_37136,N_37469);
or U37627 (N_37627,N_37485,N_37144);
nand U37628 (N_37628,N_37462,N_37148);
and U37629 (N_37629,N_37360,N_37168);
or U37630 (N_37630,N_37354,N_37232);
xor U37631 (N_37631,N_37296,N_37248);
nor U37632 (N_37632,N_37390,N_37043);
nor U37633 (N_37633,N_37133,N_37347);
xnor U37634 (N_37634,N_37466,N_37309);
nand U37635 (N_37635,N_37475,N_37396);
and U37636 (N_37636,N_37050,N_37319);
xor U37637 (N_37637,N_37107,N_37036);
or U37638 (N_37638,N_37051,N_37081);
nor U37639 (N_37639,N_37090,N_37117);
nand U37640 (N_37640,N_37101,N_37476);
or U37641 (N_37641,N_37087,N_37159);
nor U37642 (N_37642,N_37116,N_37048);
nand U37643 (N_37643,N_37233,N_37299);
nand U37644 (N_37644,N_37175,N_37388);
nand U37645 (N_37645,N_37204,N_37001);
and U37646 (N_37646,N_37254,N_37182);
and U37647 (N_37647,N_37085,N_37277);
xnor U37648 (N_37648,N_37298,N_37345);
nor U37649 (N_37649,N_37488,N_37349);
nand U37650 (N_37650,N_37016,N_37138);
nor U37651 (N_37651,N_37341,N_37351);
xor U37652 (N_37652,N_37102,N_37029);
nor U37653 (N_37653,N_37092,N_37316);
nand U37654 (N_37654,N_37392,N_37231);
and U37655 (N_37655,N_37252,N_37026);
and U37656 (N_37656,N_37443,N_37386);
or U37657 (N_37657,N_37357,N_37417);
nor U37658 (N_37658,N_37461,N_37312);
or U37659 (N_37659,N_37352,N_37291);
nand U37660 (N_37660,N_37441,N_37335);
and U37661 (N_37661,N_37009,N_37398);
or U37662 (N_37662,N_37032,N_37361);
xnor U37663 (N_37663,N_37024,N_37251);
nand U37664 (N_37664,N_37198,N_37450);
xor U37665 (N_37665,N_37099,N_37075);
nand U37666 (N_37666,N_37108,N_37222);
nand U37667 (N_37667,N_37120,N_37211);
nor U37668 (N_37668,N_37304,N_37305);
xnor U37669 (N_37669,N_37019,N_37243);
nor U37670 (N_37670,N_37183,N_37490);
nor U37671 (N_37671,N_37453,N_37086);
nor U37672 (N_37672,N_37223,N_37399);
xnor U37673 (N_37673,N_37226,N_37302);
or U37674 (N_37674,N_37190,N_37452);
nor U37675 (N_37675,N_37338,N_37123);
nand U37676 (N_37676,N_37455,N_37158);
and U37677 (N_37677,N_37114,N_37010);
nor U37678 (N_37678,N_37270,N_37472);
nor U37679 (N_37679,N_37281,N_37040);
nand U37680 (N_37680,N_37426,N_37017);
or U37681 (N_37681,N_37031,N_37262);
nand U37682 (N_37682,N_37109,N_37167);
nand U37683 (N_37683,N_37067,N_37365);
and U37684 (N_37684,N_37203,N_37104);
xor U37685 (N_37685,N_37082,N_37242);
or U37686 (N_37686,N_37076,N_37058);
and U37687 (N_37687,N_37451,N_37327);
nor U37688 (N_37688,N_37035,N_37041);
or U37689 (N_37689,N_37283,N_37187);
and U37690 (N_37690,N_37139,N_37464);
or U37691 (N_37691,N_37121,N_37363);
or U37692 (N_37692,N_37178,N_37369);
nor U37693 (N_37693,N_37260,N_37077);
or U37694 (N_37694,N_37324,N_37414);
nand U37695 (N_37695,N_37244,N_37060);
or U37696 (N_37696,N_37377,N_37367);
xor U37697 (N_37697,N_37089,N_37052);
nor U37698 (N_37698,N_37073,N_37042);
and U37699 (N_37699,N_37095,N_37034);
xor U37700 (N_37700,N_37290,N_37155);
nor U37701 (N_37701,N_37393,N_37258);
nor U37702 (N_37702,N_37179,N_37418);
xor U37703 (N_37703,N_37348,N_37434);
or U37704 (N_37704,N_37021,N_37288);
xnor U37705 (N_37705,N_37209,N_37152);
nor U37706 (N_37706,N_37395,N_37069);
and U37707 (N_37707,N_37479,N_37091);
or U37708 (N_37708,N_37272,N_37054);
xor U37709 (N_37709,N_37438,N_37230);
xor U37710 (N_37710,N_37063,N_37474);
nor U37711 (N_37711,N_37263,N_37156);
xnor U37712 (N_37712,N_37163,N_37056);
and U37713 (N_37713,N_37236,N_37482);
nor U37714 (N_37714,N_37397,N_37074);
nor U37715 (N_37715,N_37174,N_37404);
and U37716 (N_37716,N_37084,N_37326);
xnor U37717 (N_37717,N_37220,N_37006);
or U37718 (N_37718,N_37297,N_37409);
or U37719 (N_37719,N_37394,N_37194);
nand U37720 (N_37720,N_37059,N_37493);
or U37721 (N_37721,N_37240,N_37255);
nand U37722 (N_37722,N_37020,N_37483);
nor U37723 (N_37723,N_37160,N_37344);
nor U37724 (N_37724,N_37346,N_37294);
or U37725 (N_37725,N_37142,N_37447);
or U37726 (N_37726,N_37180,N_37007);
nand U37727 (N_37727,N_37310,N_37286);
nor U37728 (N_37728,N_37486,N_37343);
nand U37729 (N_37729,N_37454,N_37303);
nor U37730 (N_37730,N_37468,N_37321);
nand U37731 (N_37731,N_37300,N_37457);
and U37732 (N_37732,N_37125,N_37311);
nand U37733 (N_37733,N_37241,N_37129);
xor U37734 (N_37734,N_37478,N_37173);
nor U37735 (N_37735,N_37387,N_37375);
or U37736 (N_37736,N_37332,N_37000);
and U37737 (N_37737,N_37491,N_37362);
xnor U37738 (N_37738,N_37113,N_37463);
xnor U37739 (N_37739,N_37282,N_37047);
or U37740 (N_37740,N_37185,N_37044);
nand U37741 (N_37741,N_37169,N_37210);
xnor U37742 (N_37742,N_37172,N_37140);
and U37743 (N_37743,N_37070,N_37340);
and U37744 (N_37744,N_37278,N_37195);
xor U37745 (N_37745,N_37339,N_37477);
nand U37746 (N_37746,N_37289,N_37141);
and U37747 (N_37747,N_37098,N_37366);
or U37748 (N_37748,N_37250,N_37237);
xor U37749 (N_37749,N_37112,N_37216);
nor U37750 (N_37750,N_37072,N_37318);
xnor U37751 (N_37751,N_37464,N_37302);
nand U37752 (N_37752,N_37253,N_37463);
nand U37753 (N_37753,N_37000,N_37046);
and U37754 (N_37754,N_37121,N_37454);
xnor U37755 (N_37755,N_37353,N_37084);
or U37756 (N_37756,N_37069,N_37315);
and U37757 (N_37757,N_37279,N_37219);
nand U37758 (N_37758,N_37336,N_37055);
xor U37759 (N_37759,N_37105,N_37097);
or U37760 (N_37760,N_37350,N_37182);
or U37761 (N_37761,N_37198,N_37322);
nor U37762 (N_37762,N_37203,N_37043);
xnor U37763 (N_37763,N_37111,N_37495);
xor U37764 (N_37764,N_37262,N_37238);
and U37765 (N_37765,N_37356,N_37010);
or U37766 (N_37766,N_37433,N_37401);
nor U37767 (N_37767,N_37321,N_37255);
and U37768 (N_37768,N_37352,N_37162);
nand U37769 (N_37769,N_37057,N_37263);
nand U37770 (N_37770,N_37426,N_37235);
or U37771 (N_37771,N_37374,N_37447);
and U37772 (N_37772,N_37081,N_37230);
or U37773 (N_37773,N_37160,N_37472);
or U37774 (N_37774,N_37415,N_37435);
nand U37775 (N_37775,N_37434,N_37325);
and U37776 (N_37776,N_37025,N_37423);
nand U37777 (N_37777,N_37377,N_37445);
nor U37778 (N_37778,N_37494,N_37344);
and U37779 (N_37779,N_37280,N_37427);
xnor U37780 (N_37780,N_37398,N_37015);
nor U37781 (N_37781,N_37153,N_37148);
nand U37782 (N_37782,N_37010,N_37166);
nor U37783 (N_37783,N_37479,N_37146);
or U37784 (N_37784,N_37404,N_37421);
and U37785 (N_37785,N_37108,N_37256);
xnor U37786 (N_37786,N_37022,N_37044);
xnor U37787 (N_37787,N_37159,N_37337);
nand U37788 (N_37788,N_37085,N_37118);
nor U37789 (N_37789,N_37474,N_37292);
and U37790 (N_37790,N_37064,N_37435);
nor U37791 (N_37791,N_37097,N_37004);
nand U37792 (N_37792,N_37299,N_37234);
or U37793 (N_37793,N_37359,N_37340);
xnor U37794 (N_37794,N_37020,N_37280);
or U37795 (N_37795,N_37378,N_37193);
nor U37796 (N_37796,N_37424,N_37168);
nand U37797 (N_37797,N_37305,N_37084);
nand U37798 (N_37798,N_37159,N_37361);
nand U37799 (N_37799,N_37171,N_37205);
or U37800 (N_37800,N_37291,N_37209);
and U37801 (N_37801,N_37381,N_37152);
nand U37802 (N_37802,N_37254,N_37255);
xnor U37803 (N_37803,N_37174,N_37323);
xnor U37804 (N_37804,N_37471,N_37452);
nand U37805 (N_37805,N_37274,N_37013);
or U37806 (N_37806,N_37274,N_37021);
nor U37807 (N_37807,N_37453,N_37315);
or U37808 (N_37808,N_37326,N_37175);
xor U37809 (N_37809,N_37420,N_37435);
nor U37810 (N_37810,N_37021,N_37360);
nor U37811 (N_37811,N_37278,N_37120);
and U37812 (N_37812,N_37398,N_37062);
and U37813 (N_37813,N_37267,N_37261);
or U37814 (N_37814,N_37196,N_37167);
xor U37815 (N_37815,N_37261,N_37428);
nand U37816 (N_37816,N_37161,N_37037);
and U37817 (N_37817,N_37223,N_37332);
nor U37818 (N_37818,N_37403,N_37239);
nor U37819 (N_37819,N_37032,N_37328);
nand U37820 (N_37820,N_37122,N_37154);
or U37821 (N_37821,N_37473,N_37143);
nor U37822 (N_37822,N_37467,N_37036);
xnor U37823 (N_37823,N_37463,N_37182);
xor U37824 (N_37824,N_37408,N_37134);
xor U37825 (N_37825,N_37214,N_37057);
and U37826 (N_37826,N_37004,N_37149);
and U37827 (N_37827,N_37239,N_37137);
or U37828 (N_37828,N_37117,N_37498);
nor U37829 (N_37829,N_37453,N_37478);
nor U37830 (N_37830,N_37158,N_37493);
xnor U37831 (N_37831,N_37368,N_37137);
nand U37832 (N_37832,N_37071,N_37096);
or U37833 (N_37833,N_37182,N_37013);
or U37834 (N_37834,N_37408,N_37074);
nor U37835 (N_37835,N_37300,N_37333);
xor U37836 (N_37836,N_37227,N_37061);
nand U37837 (N_37837,N_37141,N_37421);
and U37838 (N_37838,N_37210,N_37404);
nor U37839 (N_37839,N_37016,N_37141);
or U37840 (N_37840,N_37191,N_37300);
or U37841 (N_37841,N_37303,N_37294);
and U37842 (N_37842,N_37206,N_37229);
xnor U37843 (N_37843,N_37064,N_37364);
xor U37844 (N_37844,N_37313,N_37316);
or U37845 (N_37845,N_37249,N_37486);
or U37846 (N_37846,N_37078,N_37493);
nor U37847 (N_37847,N_37126,N_37244);
and U37848 (N_37848,N_37345,N_37409);
nor U37849 (N_37849,N_37050,N_37217);
nor U37850 (N_37850,N_37113,N_37334);
or U37851 (N_37851,N_37071,N_37384);
and U37852 (N_37852,N_37459,N_37227);
nor U37853 (N_37853,N_37435,N_37402);
and U37854 (N_37854,N_37356,N_37073);
nand U37855 (N_37855,N_37100,N_37108);
nor U37856 (N_37856,N_37162,N_37302);
or U37857 (N_37857,N_37139,N_37400);
nor U37858 (N_37858,N_37058,N_37112);
nor U37859 (N_37859,N_37222,N_37374);
xnor U37860 (N_37860,N_37165,N_37082);
nand U37861 (N_37861,N_37366,N_37016);
xnor U37862 (N_37862,N_37310,N_37422);
nor U37863 (N_37863,N_37360,N_37321);
or U37864 (N_37864,N_37153,N_37042);
nand U37865 (N_37865,N_37370,N_37337);
nor U37866 (N_37866,N_37362,N_37466);
nand U37867 (N_37867,N_37020,N_37055);
nor U37868 (N_37868,N_37387,N_37061);
xnor U37869 (N_37869,N_37082,N_37087);
nor U37870 (N_37870,N_37120,N_37070);
nand U37871 (N_37871,N_37295,N_37322);
or U37872 (N_37872,N_37461,N_37147);
nor U37873 (N_37873,N_37453,N_37246);
nor U37874 (N_37874,N_37292,N_37145);
nand U37875 (N_37875,N_37285,N_37059);
and U37876 (N_37876,N_37297,N_37085);
nand U37877 (N_37877,N_37466,N_37054);
or U37878 (N_37878,N_37232,N_37008);
xor U37879 (N_37879,N_37114,N_37273);
or U37880 (N_37880,N_37239,N_37260);
nor U37881 (N_37881,N_37475,N_37472);
xnor U37882 (N_37882,N_37407,N_37057);
xnor U37883 (N_37883,N_37366,N_37108);
nand U37884 (N_37884,N_37055,N_37398);
xor U37885 (N_37885,N_37459,N_37034);
xnor U37886 (N_37886,N_37242,N_37094);
or U37887 (N_37887,N_37457,N_37021);
nand U37888 (N_37888,N_37038,N_37109);
nor U37889 (N_37889,N_37205,N_37466);
and U37890 (N_37890,N_37118,N_37371);
and U37891 (N_37891,N_37091,N_37466);
xnor U37892 (N_37892,N_37433,N_37192);
and U37893 (N_37893,N_37068,N_37060);
or U37894 (N_37894,N_37156,N_37237);
and U37895 (N_37895,N_37041,N_37208);
xnor U37896 (N_37896,N_37232,N_37054);
nor U37897 (N_37897,N_37094,N_37210);
and U37898 (N_37898,N_37186,N_37315);
nand U37899 (N_37899,N_37177,N_37344);
xnor U37900 (N_37900,N_37345,N_37210);
xor U37901 (N_37901,N_37181,N_37218);
nand U37902 (N_37902,N_37497,N_37111);
xnor U37903 (N_37903,N_37190,N_37175);
nand U37904 (N_37904,N_37461,N_37283);
xnor U37905 (N_37905,N_37244,N_37270);
or U37906 (N_37906,N_37478,N_37196);
nor U37907 (N_37907,N_37492,N_37411);
nand U37908 (N_37908,N_37425,N_37073);
nor U37909 (N_37909,N_37122,N_37227);
xor U37910 (N_37910,N_37144,N_37027);
and U37911 (N_37911,N_37414,N_37309);
nor U37912 (N_37912,N_37060,N_37079);
or U37913 (N_37913,N_37067,N_37481);
nor U37914 (N_37914,N_37253,N_37306);
or U37915 (N_37915,N_37059,N_37074);
nor U37916 (N_37916,N_37212,N_37271);
nand U37917 (N_37917,N_37134,N_37297);
nand U37918 (N_37918,N_37030,N_37120);
or U37919 (N_37919,N_37153,N_37177);
nor U37920 (N_37920,N_37358,N_37353);
xnor U37921 (N_37921,N_37442,N_37046);
xnor U37922 (N_37922,N_37368,N_37148);
or U37923 (N_37923,N_37449,N_37429);
or U37924 (N_37924,N_37350,N_37039);
nand U37925 (N_37925,N_37236,N_37309);
or U37926 (N_37926,N_37247,N_37114);
xnor U37927 (N_37927,N_37204,N_37194);
nand U37928 (N_37928,N_37390,N_37102);
nor U37929 (N_37929,N_37235,N_37090);
xor U37930 (N_37930,N_37241,N_37326);
nand U37931 (N_37931,N_37313,N_37038);
xor U37932 (N_37932,N_37188,N_37133);
nor U37933 (N_37933,N_37192,N_37481);
or U37934 (N_37934,N_37243,N_37306);
and U37935 (N_37935,N_37106,N_37358);
nor U37936 (N_37936,N_37191,N_37042);
nand U37937 (N_37937,N_37436,N_37336);
nand U37938 (N_37938,N_37396,N_37054);
and U37939 (N_37939,N_37331,N_37435);
nand U37940 (N_37940,N_37216,N_37007);
nor U37941 (N_37941,N_37119,N_37379);
or U37942 (N_37942,N_37173,N_37409);
and U37943 (N_37943,N_37092,N_37019);
nand U37944 (N_37944,N_37300,N_37183);
nand U37945 (N_37945,N_37281,N_37193);
nand U37946 (N_37946,N_37464,N_37305);
nor U37947 (N_37947,N_37228,N_37304);
xnor U37948 (N_37948,N_37326,N_37400);
nor U37949 (N_37949,N_37086,N_37267);
xor U37950 (N_37950,N_37307,N_37103);
nor U37951 (N_37951,N_37212,N_37433);
and U37952 (N_37952,N_37411,N_37101);
or U37953 (N_37953,N_37233,N_37153);
or U37954 (N_37954,N_37301,N_37447);
nor U37955 (N_37955,N_37363,N_37186);
or U37956 (N_37956,N_37042,N_37410);
nor U37957 (N_37957,N_37368,N_37027);
nand U37958 (N_37958,N_37091,N_37279);
nor U37959 (N_37959,N_37356,N_37125);
nand U37960 (N_37960,N_37001,N_37495);
nand U37961 (N_37961,N_37392,N_37394);
and U37962 (N_37962,N_37263,N_37085);
or U37963 (N_37963,N_37168,N_37103);
nand U37964 (N_37964,N_37098,N_37471);
xnor U37965 (N_37965,N_37180,N_37484);
xnor U37966 (N_37966,N_37412,N_37379);
or U37967 (N_37967,N_37109,N_37148);
xnor U37968 (N_37968,N_37306,N_37166);
xnor U37969 (N_37969,N_37002,N_37445);
or U37970 (N_37970,N_37427,N_37380);
nand U37971 (N_37971,N_37335,N_37019);
or U37972 (N_37972,N_37447,N_37288);
xor U37973 (N_37973,N_37440,N_37191);
xnor U37974 (N_37974,N_37388,N_37223);
xnor U37975 (N_37975,N_37096,N_37145);
and U37976 (N_37976,N_37018,N_37255);
nand U37977 (N_37977,N_37371,N_37143);
and U37978 (N_37978,N_37090,N_37251);
nor U37979 (N_37979,N_37416,N_37050);
nor U37980 (N_37980,N_37349,N_37247);
nor U37981 (N_37981,N_37160,N_37019);
nand U37982 (N_37982,N_37075,N_37357);
or U37983 (N_37983,N_37353,N_37345);
or U37984 (N_37984,N_37072,N_37181);
nand U37985 (N_37985,N_37366,N_37352);
nor U37986 (N_37986,N_37057,N_37346);
nor U37987 (N_37987,N_37072,N_37345);
and U37988 (N_37988,N_37450,N_37150);
xor U37989 (N_37989,N_37319,N_37188);
nand U37990 (N_37990,N_37170,N_37126);
nor U37991 (N_37991,N_37153,N_37330);
or U37992 (N_37992,N_37404,N_37060);
and U37993 (N_37993,N_37006,N_37120);
and U37994 (N_37994,N_37251,N_37369);
or U37995 (N_37995,N_37344,N_37307);
or U37996 (N_37996,N_37267,N_37236);
nand U37997 (N_37997,N_37473,N_37141);
and U37998 (N_37998,N_37178,N_37185);
xor U37999 (N_37999,N_37302,N_37378);
and U38000 (N_38000,N_37980,N_37616);
and U38001 (N_38001,N_37706,N_37632);
nor U38002 (N_38002,N_37537,N_37508);
xor U38003 (N_38003,N_37802,N_37822);
or U38004 (N_38004,N_37887,N_37660);
nor U38005 (N_38005,N_37920,N_37948);
nor U38006 (N_38006,N_37534,N_37964);
or U38007 (N_38007,N_37691,N_37925);
nand U38008 (N_38008,N_37649,N_37690);
xnor U38009 (N_38009,N_37525,N_37772);
nand U38010 (N_38010,N_37864,N_37747);
nor U38011 (N_38011,N_37638,N_37795);
nand U38012 (N_38012,N_37698,N_37914);
and U38013 (N_38013,N_37781,N_37613);
or U38014 (N_38014,N_37503,N_37778);
or U38015 (N_38015,N_37930,N_37669);
nor U38016 (N_38016,N_37788,N_37833);
and U38017 (N_38017,N_37528,N_37770);
nand U38018 (N_38018,N_37851,N_37883);
nor U38019 (N_38019,N_37659,N_37861);
or U38020 (N_38020,N_37652,N_37745);
nand U38021 (N_38021,N_37868,N_37843);
or U38022 (N_38022,N_37714,N_37985);
or U38023 (N_38023,N_37908,N_37927);
and U38024 (N_38024,N_37876,N_37682);
nand U38025 (N_38025,N_37517,N_37607);
or U38026 (N_38026,N_37898,N_37764);
and U38027 (N_38027,N_37553,N_37824);
or U38028 (N_38028,N_37611,N_37685);
or U38029 (N_38029,N_37830,N_37974);
nand U38030 (N_38030,N_37521,N_37842);
nand U38031 (N_38031,N_37501,N_37535);
or U38032 (N_38032,N_37711,N_37606);
xor U38033 (N_38033,N_37641,N_37979);
xor U38034 (N_38034,N_37716,N_37936);
and U38035 (N_38035,N_37813,N_37857);
nand U38036 (N_38036,N_37963,N_37730);
and U38037 (N_38037,N_37972,N_37539);
nor U38038 (N_38038,N_37831,N_37579);
and U38039 (N_38039,N_37926,N_37633);
nand U38040 (N_38040,N_37951,N_37835);
nor U38041 (N_38041,N_37882,N_37961);
or U38042 (N_38042,N_37913,N_37618);
and U38043 (N_38043,N_37810,N_37792);
and U38044 (N_38044,N_37688,N_37605);
xor U38045 (N_38045,N_37811,N_37976);
or U38046 (N_38046,N_37960,N_37958);
nand U38047 (N_38047,N_37574,N_37837);
nor U38048 (N_38048,N_37860,N_37939);
and U38049 (N_38049,N_37738,N_37526);
and U38050 (N_38050,N_37762,N_37694);
nor U38051 (N_38051,N_37749,N_37756);
nand U38052 (N_38052,N_37829,N_37905);
xnor U38053 (N_38053,N_37916,N_37752);
nand U38054 (N_38054,N_37945,N_37547);
nor U38055 (N_38055,N_37946,N_37949);
nor U38056 (N_38056,N_37911,N_37844);
nand U38057 (N_38057,N_37877,N_37990);
nand U38058 (N_38058,N_37769,N_37594);
and U38059 (N_38059,N_37970,N_37982);
xor U38060 (N_38060,N_37922,N_37999);
xor U38061 (N_38061,N_37603,N_37773);
and U38062 (N_38062,N_37771,N_37591);
nand U38063 (N_38063,N_37507,N_37689);
nand U38064 (N_38064,N_37601,N_37997);
or U38065 (N_38065,N_37696,N_37944);
nand U38066 (N_38066,N_37973,N_37677);
nor U38067 (N_38067,N_37675,N_37597);
xnor U38068 (N_38068,N_37702,N_37672);
and U38069 (N_38069,N_37955,N_37619);
nor U38070 (N_38070,N_37583,N_37518);
nor U38071 (N_38071,N_37741,N_37943);
or U38072 (N_38072,N_37530,N_37524);
and U38073 (N_38073,N_37719,N_37701);
or U38074 (N_38074,N_37707,N_37840);
nand U38075 (N_38075,N_37823,N_37753);
or U38076 (N_38076,N_37971,N_37984);
and U38077 (N_38077,N_37871,N_37846);
and U38078 (N_38078,N_37581,N_37998);
xor U38079 (N_38079,N_37504,N_37636);
or U38080 (N_38080,N_37931,N_37630);
or U38081 (N_38081,N_37673,N_37902);
nor U38082 (N_38082,N_37895,N_37721);
and U38083 (N_38083,N_37536,N_37687);
nor U38084 (N_38084,N_37584,N_37548);
or U38085 (N_38085,N_37748,N_37661);
and U38086 (N_38086,N_37765,N_37897);
and U38087 (N_38087,N_37845,N_37903);
and U38088 (N_38088,N_37968,N_37639);
or U38089 (N_38089,N_37545,N_37587);
nand U38090 (N_38090,N_37866,N_37839);
or U38091 (N_38091,N_37523,N_37855);
xnor U38092 (N_38092,N_37777,N_37870);
or U38093 (N_38093,N_37667,N_37774);
nand U38094 (N_38094,N_37737,N_37631);
and U38095 (N_38095,N_37890,N_37541);
nand U38096 (N_38096,N_37783,N_37733);
or U38097 (N_38097,N_37695,N_37699);
nand U38098 (N_38098,N_37917,N_37867);
nand U38099 (N_38099,N_37912,N_37683);
nor U38100 (N_38100,N_37801,N_37635);
and U38101 (N_38101,N_37856,N_37620);
nand U38102 (N_38102,N_37686,N_37546);
nor U38103 (N_38103,N_37891,N_37570);
nor U38104 (N_38104,N_37848,N_37836);
and U38105 (N_38105,N_37894,N_37726);
xnor U38106 (N_38106,N_37780,N_37556);
nor U38107 (N_38107,N_37700,N_37983);
nand U38108 (N_38108,N_37892,N_37743);
or U38109 (N_38109,N_37826,N_37657);
and U38110 (N_38110,N_37977,N_37820);
and U38111 (N_38111,N_37703,N_37608);
xor U38112 (N_38112,N_37676,N_37531);
nor U38113 (N_38113,N_37713,N_37874);
nand U38114 (N_38114,N_37992,N_37950);
nor U38115 (N_38115,N_37626,N_37612);
or U38116 (N_38116,N_37940,N_37670);
or U38117 (N_38117,N_37858,N_37907);
nand U38118 (N_38118,N_37995,N_37589);
nand U38119 (N_38119,N_37881,N_37763);
nand U38120 (N_38120,N_37720,N_37712);
xnor U38121 (N_38121,N_37991,N_37827);
and U38122 (N_38122,N_37599,N_37760);
or U38123 (N_38123,N_37723,N_37566);
nor U38124 (N_38124,N_37662,N_37684);
nor U38125 (N_38125,N_37564,N_37527);
xnor U38126 (N_38126,N_37989,N_37893);
nand U38127 (N_38127,N_37679,N_37511);
and U38128 (N_38128,N_37933,N_37932);
nand U38129 (N_38129,N_37655,N_37622);
and U38130 (N_38130,N_37568,N_37896);
and U38131 (N_38131,N_37578,N_37617);
nand U38132 (N_38132,N_37596,N_37966);
xor U38133 (N_38133,N_37766,N_37804);
xor U38134 (N_38134,N_37602,N_37551);
and U38135 (N_38135,N_37558,N_37921);
nand U38136 (N_38136,N_37656,N_37625);
xor U38137 (N_38137,N_37799,N_37888);
nor U38138 (N_38138,N_37915,N_37767);
xor U38139 (N_38139,N_37965,N_37592);
xnor U38140 (N_38140,N_37538,N_37665);
nand U38141 (N_38141,N_37994,N_37727);
xor U38142 (N_38142,N_37807,N_37668);
xor U38143 (N_38143,N_37585,N_37614);
nand U38144 (N_38144,N_37953,N_37704);
xnor U38145 (N_38145,N_37885,N_37873);
or U38146 (N_38146,N_37814,N_37658);
and U38147 (N_38147,N_37934,N_37506);
and U38148 (N_38148,N_37593,N_37549);
and U38149 (N_38149,N_37697,N_37879);
nor U38150 (N_38150,N_37821,N_37825);
and U38151 (N_38151,N_37654,N_37938);
nor U38152 (N_38152,N_37988,N_37828);
xnor U38153 (N_38153,N_37775,N_37906);
nand U38154 (N_38154,N_37648,N_37862);
or U38155 (N_38155,N_37744,N_37941);
xor U38156 (N_38156,N_37650,N_37812);
and U38157 (N_38157,N_37852,N_37803);
xnor U38158 (N_38158,N_37975,N_37645);
or U38159 (N_38159,N_37863,N_37969);
nand U38160 (N_38160,N_37954,N_37731);
xor U38161 (N_38161,N_37751,N_37609);
xnor U38162 (N_38162,N_37981,N_37865);
nand U38163 (N_38163,N_37816,N_37629);
and U38164 (N_38164,N_37937,N_37910);
and U38165 (N_38165,N_37554,N_37878);
and U38166 (N_38166,N_37834,N_37758);
and U38167 (N_38167,N_37595,N_37776);
and U38168 (N_38168,N_37790,N_37952);
or U38169 (N_38169,N_37853,N_37901);
and U38170 (N_38170,N_37663,N_37886);
xnor U38171 (N_38171,N_37520,N_37815);
xnor U38172 (N_38172,N_37653,N_37900);
or U38173 (N_38173,N_37563,N_37582);
nor U38174 (N_38174,N_37782,N_37515);
nor U38175 (N_38175,N_37957,N_37859);
xnor U38176 (N_38176,N_37544,N_37550);
nor U38177 (N_38177,N_37516,N_37509);
xnor U38178 (N_38178,N_37746,N_37722);
nor U38179 (N_38179,N_37791,N_37996);
and U38180 (N_38180,N_37789,N_37604);
or U38181 (N_38181,N_37987,N_37797);
or U38182 (N_38182,N_37959,N_37728);
xor U38183 (N_38183,N_37500,N_37598);
nor U38184 (N_38184,N_37717,N_37875);
xor U38185 (N_38185,N_37519,N_37784);
or U38186 (N_38186,N_37757,N_37787);
nand U38187 (N_38187,N_37838,N_37580);
nand U38188 (N_38188,N_37678,N_37889);
or U38189 (N_38189,N_37725,N_37627);
nand U38190 (N_38190,N_37806,N_37674);
and U38191 (N_38191,N_37572,N_37805);
or U38192 (N_38192,N_37935,N_37732);
nor U38193 (N_38193,N_37904,N_37586);
nand U38194 (N_38194,N_37588,N_37565);
nand U38195 (N_38195,N_37628,N_37739);
and U38196 (N_38196,N_37512,N_37647);
or U38197 (N_38197,N_37542,N_37567);
or U38198 (N_38198,N_37850,N_37754);
nand U38199 (N_38199,N_37817,N_37575);
nor U38200 (N_38200,N_37557,N_37561);
and U38201 (N_38201,N_37899,N_37569);
nand U38202 (N_38202,N_37522,N_37734);
nor U38203 (N_38203,N_37590,N_37967);
nand U38204 (N_38204,N_37786,N_37540);
and U38205 (N_38205,N_37841,N_37798);
or U38206 (N_38206,N_37750,N_37708);
nand U38207 (N_38207,N_37529,N_37884);
or U38208 (N_38208,N_37642,N_37793);
and U38209 (N_38209,N_37615,N_37577);
nand U38210 (N_38210,N_37552,N_37768);
xor U38211 (N_38211,N_37740,N_37718);
or U38212 (N_38212,N_37571,N_37923);
and U38213 (N_38213,N_37929,N_37819);
nand U38214 (N_38214,N_37724,N_37710);
nand U38215 (N_38215,N_37505,N_37735);
xnor U38216 (N_38216,N_37736,N_37555);
or U38217 (N_38217,N_37681,N_37779);
xnor U38218 (N_38218,N_37854,N_37847);
xnor U38219 (N_38219,N_37705,N_37514);
and U38220 (N_38220,N_37947,N_37956);
xnor U38221 (N_38221,N_37573,N_37794);
or U38222 (N_38222,N_37513,N_37576);
or U38223 (N_38223,N_37909,N_37640);
nor U38224 (N_38224,N_37624,N_37942);
nor U38225 (N_38225,N_37621,N_37644);
nor U38226 (N_38226,N_37962,N_37869);
xor U38227 (N_38227,N_37634,N_37533);
or U38228 (N_38228,N_37510,N_37643);
nand U38229 (N_38229,N_37872,N_37693);
nand U38230 (N_38230,N_37919,N_37715);
or U38231 (N_38231,N_37646,N_37832);
or U38232 (N_38232,N_37560,N_37543);
xnor U38233 (N_38233,N_37924,N_37651);
nor U38234 (N_38234,N_37800,N_37502);
or U38235 (N_38235,N_37671,N_37709);
and U38236 (N_38236,N_37637,N_37680);
and U38237 (N_38237,N_37532,N_37559);
nand U38238 (N_38238,N_37755,N_37666);
xor U38239 (N_38239,N_37759,N_37610);
xnor U38240 (N_38240,N_37978,N_37809);
or U38241 (N_38241,N_37761,N_37729);
and U38242 (N_38242,N_37993,N_37785);
nand U38243 (N_38243,N_37796,N_37562);
or U38244 (N_38244,N_37623,N_37818);
and U38245 (N_38245,N_37692,N_37742);
or U38246 (N_38246,N_37664,N_37880);
and U38247 (N_38247,N_37928,N_37986);
nand U38248 (N_38248,N_37918,N_37600);
nand U38249 (N_38249,N_37808,N_37849);
nand U38250 (N_38250,N_37633,N_37796);
or U38251 (N_38251,N_37976,N_37824);
nand U38252 (N_38252,N_37735,N_37828);
nor U38253 (N_38253,N_37651,N_37585);
and U38254 (N_38254,N_37892,N_37905);
nor U38255 (N_38255,N_37789,N_37560);
xor U38256 (N_38256,N_37745,N_37697);
and U38257 (N_38257,N_37786,N_37604);
nand U38258 (N_38258,N_37917,N_37630);
xnor U38259 (N_38259,N_37763,N_37670);
nand U38260 (N_38260,N_37864,N_37587);
or U38261 (N_38261,N_37554,N_37635);
nand U38262 (N_38262,N_37555,N_37717);
and U38263 (N_38263,N_37784,N_37779);
nor U38264 (N_38264,N_37818,N_37639);
nor U38265 (N_38265,N_37795,N_37888);
or U38266 (N_38266,N_37574,N_37704);
or U38267 (N_38267,N_37761,N_37733);
nand U38268 (N_38268,N_37619,N_37920);
nand U38269 (N_38269,N_37846,N_37617);
or U38270 (N_38270,N_37923,N_37699);
xnor U38271 (N_38271,N_37534,N_37624);
xor U38272 (N_38272,N_37979,N_37902);
and U38273 (N_38273,N_37936,N_37759);
and U38274 (N_38274,N_37806,N_37926);
or U38275 (N_38275,N_37573,N_37868);
xnor U38276 (N_38276,N_37991,N_37714);
and U38277 (N_38277,N_37985,N_37704);
or U38278 (N_38278,N_37902,N_37840);
or U38279 (N_38279,N_37666,N_37779);
xor U38280 (N_38280,N_37725,N_37641);
nand U38281 (N_38281,N_37709,N_37933);
xor U38282 (N_38282,N_37810,N_37643);
and U38283 (N_38283,N_37862,N_37735);
nor U38284 (N_38284,N_37891,N_37533);
nor U38285 (N_38285,N_37647,N_37604);
nand U38286 (N_38286,N_37758,N_37860);
and U38287 (N_38287,N_37500,N_37816);
and U38288 (N_38288,N_37649,N_37985);
nor U38289 (N_38289,N_37898,N_37552);
nand U38290 (N_38290,N_37533,N_37541);
nor U38291 (N_38291,N_37633,N_37592);
nor U38292 (N_38292,N_37761,N_37714);
nand U38293 (N_38293,N_37565,N_37655);
and U38294 (N_38294,N_37518,N_37978);
and U38295 (N_38295,N_37799,N_37871);
and U38296 (N_38296,N_37865,N_37987);
or U38297 (N_38297,N_37943,N_37957);
nor U38298 (N_38298,N_37611,N_37533);
and U38299 (N_38299,N_37529,N_37574);
and U38300 (N_38300,N_37877,N_37814);
nand U38301 (N_38301,N_37843,N_37650);
xnor U38302 (N_38302,N_37632,N_37502);
and U38303 (N_38303,N_37844,N_37971);
or U38304 (N_38304,N_37683,N_37761);
and U38305 (N_38305,N_37914,N_37907);
or U38306 (N_38306,N_37854,N_37512);
xnor U38307 (N_38307,N_37515,N_37899);
nand U38308 (N_38308,N_37719,N_37864);
xor U38309 (N_38309,N_37558,N_37923);
or U38310 (N_38310,N_37859,N_37927);
nor U38311 (N_38311,N_37518,N_37513);
xor U38312 (N_38312,N_37734,N_37609);
nor U38313 (N_38313,N_37927,N_37697);
and U38314 (N_38314,N_37962,N_37578);
and U38315 (N_38315,N_37617,N_37969);
or U38316 (N_38316,N_37609,N_37855);
nand U38317 (N_38317,N_37549,N_37819);
nor U38318 (N_38318,N_37837,N_37880);
nor U38319 (N_38319,N_37866,N_37674);
or U38320 (N_38320,N_37803,N_37711);
nand U38321 (N_38321,N_37809,N_37705);
and U38322 (N_38322,N_37998,N_37858);
xor U38323 (N_38323,N_37656,N_37710);
and U38324 (N_38324,N_37742,N_37582);
xnor U38325 (N_38325,N_37907,N_37670);
or U38326 (N_38326,N_37598,N_37518);
nand U38327 (N_38327,N_37646,N_37971);
nand U38328 (N_38328,N_37551,N_37577);
nand U38329 (N_38329,N_37744,N_37545);
nand U38330 (N_38330,N_37625,N_37875);
xnor U38331 (N_38331,N_37698,N_37797);
and U38332 (N_38332,N_37737,N_37521);
or U38333 (N_38333,N_37643,N_37752);
and U38334 (N_38334,N_37945,N_37664);
nor U38335 (N_38335,N_37871,N_37889);
nand U38336 (N_38336,N_37852,N_37779);
xnor U38337 (N_38337,N_37654,N_37648);
or U38338 (N_38338,N_37632,N_37789);
nor U38339 (N_38339,N_37567,N_37766);
nor U38340 (N_38340,N_37597,N_37566);
xnor U38341 (N_38341,N_37853,N_37662);
and U38342 (N_38342,N_37840,N_37920);
nor U38343 (N_38343,N_37650,N_37747);
nor U38344 (N_38344,N_37833,N_37618);
xnor U38345 (N_38345,N_37738,N_37941);
nor U38346 (N_38346,N_37893,N_37915);
nand U38347 (N_38347,N_37676,N_37580);
or U38348 (N_38348,N_37934,N_37852);
nor U38349 (N_38349,N_37538,N_37518);
nand U38350 (N_38350,N_37948,N_37507);
nand U38351 (N_38351,N_37629,N_37951);
nor U38352 (N_38352,N_37701,N_37512);
or U38353 (N_38353,N_37814,N_37899);
or U38354 (N_38354,N_37522,N_37861);
xnor U38355 (N_38355,N_37921,N_37507);
or U38356 (N_38356,N_37747,N_37927);
or U38357 (N_38357,N_37815,N_37792);
xnor U38358 (N_38358,N_37812,N_37607);
or U38359 (N_38359,N_37984,N_37654);
nand U38360 (N_38360,N_37685,N_37794);
nor U38361 (N_38361,N_37973,N_37975);
or U38362 (N_38362,N_37897,N_37577);
and U38363 (N_38363,N_37855,N_37893);
nor U38364 (N_38364,N_37778,N_37968);
or U38365 (N_38365,N_37607,N_37879);
nor U38366 (N_38366,N_37745,N_37783);
and U38367 (N_38367,N_37795,N_37966);
nor U38368 (N_38368,N_37777,N_37802);
or U38369 (N_38369,N_37648,N_37744);
and U38370 (N_38370,N_37988,N_37997);
or U38371 (N_38371,N_37882,N_37604);
or U38372 (N_38372,N_37897,N_37754);
xor U38373 (N_38373,N_37910,N_37880);
xor U38374 (N_38374,N_37681,N_37978);
nand U38375 (N_38375,N_37991,N_37962);
xor U38376 (N_38376,N_37810,N_37743);
or U38377 (N_38377,N_37586,N_37920);
xnor U38378 (N_38378,N_37618,N_37950);
nor U38379 (N_38379,N_37936,N_37628);
or U38380 (N_38380,N_37934,N_37660);
and U38381 (N_38381,N_37731,N_37712);
xnor U38382 (N_38382,N_37710,N_37944);
nand U38383 (N_38383,N_37872,N_37882);
and U38384 (N_38384,N_37994,N_37971);
nor U38385 (N_38385,N_37735,N_37646);
xnor U38386 (N_38386,N_37941,N_37948);
or U38387 (N_38387,N_37524,N_37878);
xnor U38388 (N_38388,N_37742,N_37768);
xor U38389 (N_38389,N_37821,N_37976);
nand U38390 (N_38390,N_37712,N_37634);
and U38391 (N_38391,N_37643,N_37964);
nor U38392 (N_38392,N_37634,N_37836);
or U38393 (N_38393,N_37999,N_37994);
and U38394 (N_38394,N_37761,N_37700);
or U38395 (N_38395,N_37861,N_37725);
or U38396 (N_38396,N_37731,N_37601);
xnor U38397 (N_38397,N_37588,N_37608);
nor U38398 (N_38398,N_37758,N_37631);
nor U38399 (N_38399,N_37972,N_37571);
nand U38400 (N_38400,N_37719,N_37882);
and U38401 (N_38401,N_37705,N_37791);
nor U38402 (N_38402,N_37531,N_37601);
nand U38403 (N_38403,N_37593,N_37967);
nand U38404 (N_38404,N_37698,N_37912);
xor U38405 (N_38405,N_37608,N_37809);
or U38406 (N_38406,N_37608,N_37636);
nand U38407 (N_38407,N_37981,N_37971);
xor U38408 (N_38408,N_37846,N_37633);
or U38409 (N_38409,N_37562,N_37983);
or U38410 (N_38410,N_37586,N_37984);
nor U38411 (N_38411,N_37985,N_37505);
nor U38412 (N_38412,N_37535,N_37732);
nand U38413 (N_38413,N_37866,N_37947);
xor U38414 (N_38414,N_37541,N_37732);
xor U38415 (N_38415,N_37501,N_37651);
and U38416 (N_38416,N_37508,N_37768);
and U38417 (N_38417,N_37839,N_37653);
and U38418 (N_38418,N_37786,N_37545);
nand U38419 (N_38419,N_37710,N_37894);
nand U38420 (N_38420,N_37911,N_37806);
or U38421 (N_38421,N_37905,N_37620);
nor U38422 (N_38422,N_37966,N_37601);
xnor U38423 (N_38423,N_37701,N_37965);
or U38424 (N_38424,N_37814,N_37862);
or U38425 (N_38425,N_37516,N_37543);
nor U38426 (N_38426,N_37719,N_37692);
xor U38427 (N_38427,N_37994,N_37767);
nand U38428 (N_38428,N_37742,N_37887);
xor U38429 (N_38429,N_37960,N_37567);
or U38430 (N_38430,N_37534,N_37794);
and U38431 (N_38431,N_37794,N_37780);
xor U38432 (N_38432,N_37528,N_37794);
and U38433 (N_38433,N_37532,N_37796);
or U38434 (N_38434,N_37568,N_37614);
or U38435 (N_38435,N_37947,N_37558);
nand U38436 (N_38436,N_37665,N_37995);
nor U38437 (N_38437,N_37670,N_37617);
and U38438 (N_38438,N_37570,N_37987);
and U38439 (N_38439,N_37570,N_37772);
or U38440 (N_38440,N_37907,N_37984);
nand U38441 (N_38441,N_37808,N_37935);
and U38442 (N_38442,N_37983,N_37705);
or U38443 (N_38443,N_37720,N_37651);
nor U38444 (N_38444,N_37701,N_37996);
xor U38445 (N_38445,N_37915,N_37838);
xnor U38446 (N_38446,N_37590,N_37690);
and U38447 (N_38447,N_37630,N_37670);
nand U38448 (N_38448,N_37658,N_37535);
nand U38449 (N_38449,N_37659,N_37576);
and U38450 (N_38450,N_37964,N_37576);
or U38451 (N_38451,N_37889,N_37938);
nand U38452 (N_38452,N_37677,N_37946);
and U38453 (N_38453,N_37862,N_37971);
and U38454 (N_38454,N_37629,N_37560);
xor U38455 (N_38455,N_37978,N_37659);
or U38456 (N_38456,N_37748,N_37796);
nand U38457 (N_38457,N_37517,N_37870);
nand U38458 (N_38458,N_37511,N_37829);
nor U38459 (N_38459,N_37791,N_37752);
xor U38460 (N_38460,N_37868,N_37810);
or U38461 (N_38461,N_37534,N_37753);
nand U38462 (N_38462,N_37850,N_37642);
xnor U38463 (N_38463,N_37618,N_37911);
or U38464 (N_38464,N_37897,N_37996);
or U38465 (N_38465,N_37703,N_37580);
nor U38466 (N_38466,N_37638,N_37966);
nand U38467 (N_38467,N_37889,N_37562);
nor U38468 (N_38468,N_37572,N_37742);
nor U38469 (N_38469,N_37826,N_37896);
nor U38470 (N_38470,N_37604,N_37837);
nor U38471 (N_38471,N_37591,N_37540);
or U38472 (N_38472,N_37866,N_37772);
nor U38473 (N_38473,N_37919,N_37762);
nor U38474 (N_38474,N_37929,N_37741);
nor U38475 (N_38475,N_37852,N_37652);
and U38476 (N_38476,N_37817,N_37729);
nand U38477 (N_38477,N_37760,N_37509);
and U38478 (N_38478,N_37548,N_37606);
xnor U38479 (N_38479,N_37842,N_37740);
xor U38480 (N_38480,N_37562,N_37585);
and U38481 (N_38481,N_37557,N_37618);
xor U38482 (N_38482,N_37605,N_37864);
nand U38483 (N_38483,N_37997,N_37667);
xor U38484 (N_38484,N_37796,N_37746);
nor U38485 (N_38485,N_37964,N_37876);
or U38486 (N_38486,N_37603,N_37870);
nand U38487 (N_38487,N_37549,N_37542);
xnor U38488 (N_38488,N_37967,N_37739);
nand U38489 (N_38489,N_37679,N_37541);
and U38490 (N_38490,N_37542,N_37675);
or U38491 (N_38491,N_37977,N_37674);
nand U38492 (N_38492,N_37822,N_37675);
and U38493 (N_38493,N_37968,N_37719);
nand U38494 (N_38494,N_37658,N_37561);
xor U38495 (N_38495,N_37645,N_37736);
or U38496 (N_38496,N_37891,N_37791);
and U38497 (N_38497,N_37925,N_37693);
or U38498 (N_38498,N_37976,N_37777);
nor U38499 (N_38499,N_37842,N_37917);
xor U38500 (N_38500,N_38111,N_38125);
nand U38501 (N_38501,N_38102,N_38114);
nor U38502 (N_38502,N_38479,N_38216);
and U38503 (N_38503,N_38331,N_38217);
nor U38504 (N_38504,N_38134,N_38237);
nor U38505 (N_38505,N_38087,N_38082);
nand U38506 (N_38506,N_38289,N_38170);
nand U38507 (N_38507,N_38232,N_38422);
and U38508 (N_38508,N_38341,N_38010);
or U38509 (N_38509,N_38024,N_38033);
nor U38510 (N_38510,N_38107,N_38393);
nor U38511 (N_38511,N_38363,N_38303);
xor U38512 (N_38512,N_38262,N_38366);
nor U38513 (N_38513,N_38357,N_38060);
nand U38514 (N_38514,N_38345,N_38263);
and U38515 (N_38515,N_38412,N_38239);
xor U38516 (N_38516,N_38273,N_38380);
or U38517 (N_38517,N_38004,N_38038);
or U38518 (N_38518,N_38052,N_38280);
nand U38519 (N_38519,N_38208,N_38297);
xor U38520 (N_38520,N_38238,N_38181);
and U38521 (N_38521,N_38295,N_38453);
or U38522 (N_38522,N_38104,N_38118);
xnor U38523 (N_38523,N_38196,N_38356);
and U38524 (N_38524,N_38046,N_38346);
nor U38525 (N_38525,N_38340,N_38031);
xor U38526 (N_38526,N_38386,N_38016);
nor U38527 (N_38527,N_38207,N_38351);
or U38528 (N_38528,N_38235,N_38186);
nand U38529 (N_38529,N_38395,N_38091);
xnor U38530 (N_38530,N_38197,N_38265);
nor U38531 (N_38531,N_38483,N_38308);
and U38532 (N_38532,N_38244,N_38193);
and U38533 (N_38533,N_38309,N_38173);
xnor U38534 (N_38534,N_38218,N_38471);
nor U38535 (N_38535,N_38079,N_38122);
nand U38536 (N_38536,N_38204,N_38490);
and U38537 (N_38537,N_38360,N_38361);
and U38538 (N_38538,N_38246,N_38319);
nor U38539 (N_38539,N_38450,N_38150);
nand U38540 (N_38540,N_38165,N_38278);
xor U38541 (N_38541,N_38113,N_38228);
nor U38542 (N_38542,N_38005,N_38473);
nand U38543 (N_38543,N_38027,N_38013);
nor U38544 (N_38544,N_38375,N_38063);
or U38545 (N_38545,N_38410,N_38190);
xnor U38546 (N_38546,N_38030,N_38347);
and U38547 (N_38547,N_38466,N_38406);
or U38548 (N_38548,N_38183,N_38401);
and U38549 (N_38549,N_38432,N_38390);
nor U38550 (N_38550,N_38428,N_38469);
nor U38551 (N_38551,N_38408,N_38126);
and U38552 (N_38552,N_38459,N_38311);
nor U38553 (N_38553,N_38089,N_38068);
or U38554 (N_38554,N_38270,N_38279);
nand U38555 (N_38555,N_38103,N_38168);
nor U38556 (N_38556,N_38298,N_38236);
or U38557 (N_38557,N_38369,N_38499);
nand U38558 (N_38558,N_38172,N_38336);
xor U38559 (N_38559,N_38189,N_38036);
xor U38560 (N_38560,N_38026,N_38137);
or U38561 (N_38561,N_38159,N_38350);
or U38562 (N_38562,N_38066,N_38166);
xnor U38563 (N_38563,N_38081,N_38040);
xor U38564 (N_38564,N_38313,N_38498);
nor U38565 (N_38565,N_38439,N_38489);
xnor U38566 (N_38566,N_38225,N_38250);
nand U38567 (N_38567,N_38149,N_38438);
and U38568 (N_38568,N_38025,N_38153);
nand U38569 (N_38569,N_38458,N_38203);
xnor U38570 (N_38570,N_38051,N_38397);
and U38571 (N_38571,N_38230,N_38160);
xnor U38572 (N_38572,N_38413,N_38171);
or U38573 (N_38573,N_38185,N_38077);
or U38574 (N_38574,N_38292,N_38272);
and U38575 (N_38575,N_38404,N_38222);
and U38576 (N_38576,N_38106,N_38449);
or U38577 (N_38577,N_38461,N_38074);
xor U38578 (N_38578,N_38129,N_38318);
xnor U38579 (N_38579,N_38055,N_38426);
and U38580 (N_38580,N_38001,N_38493);
nor U38581 (N_38581,N_38117,N_38101);
or U38582 (N_38582,N_38241,N_38049);
or U38583 (N_38583,N_38056,N_38044);
xor U38584 (N_38584,N_38067,N_38156);
or U38585 (N_38585,N_38492,N_38215);
xnor U38586 (N_38586,N_38097,N_38271);
nand U38587 (N_38587,N_38000,N_38023);
and U38588 (N_38588,N_38353,N_38269);
nand U38589 (N_38589,N_38274,N_38064);
nand U38590 (N_38590,N_38403,N_38096);
xnor U38591 (N_38591,N_38478,N_38317);
nand U38592 (N_38592,N_38048,N_38304);
and U38593 (N_38593,N_38121,N_38420);
or U38594 (N_38594,N_38099,N_38179);
xor U38595 (N_38595,N_38291,N_38212);
nor U38596 (N_38596,N_38021,N_38437);
xor U38597 (N_38597,N_38327,N_38145);
nor U38598 (N_38598,N_38136,N_38042);
or U38599 (N_38599,N_38022,N_38451);
xor U38600 (N_38600,N_38391,N_38251);
or U38601 (N_38601,N_38180,N_38339);
nand U38602 (N_38602,N_38491,N_38258);
nand U38603 (N_38603,N_38110,N_38431);
nand U38604 (N_38604,N_38465,N_38226);
nor U38605 (N_38605,N_38070,N_38047);
nor U38606 (N_38606,N_38164,N_38039);
and U38607 (N_38607,N_38456,N_38028);
xor U38608 (N_38608,N_38383,N_38482);
xnor U38609 (N_38609,N_38050,N_38109);
xnor U38610 (N_38610,N_38470,N_38384);
nor U38611 (N_38611,N_38205,N_38201);
or U38612 (N_38612,N_38371,N_38299);
or U38613 (N_38613,N_38264,N_38300);
nand U38614 (N_38614,N_38368,N_38276);
and U38615 (N_38615,N_38476,N_38133);
nand U38616 (N_38616,N_38095,N_38090);
and U38617 (N_38617,N_38256,N_38116);
xnor U38618 (N_38618,N_38169,N_38301);
nor U38619 (N_38619,N_38058,N_38310);
and U38620 (N_38620,N_38488,N_38455);
nor U38621 (N_38621,N_38247,N_38381);
nand U38622 (N_38622,N_38061,N_38322);
or U38623 (N_38623,N_38143,N_38198);
nor U38624 (N_38624,N_38321,N_38480);
and U38625 (N_38625,N_38253,N_38192);
xor U38626 (N_38626,N_38372,N_38359);
nor U38627 (N_38627,N_38120,N_38324);
xor U38628 (N_38628,N_38379,N_38259);
nand U38629 (N_38629,N_38337,N_38487);
or U38630 (N_38630,N_38037,N_38243);
nor U38631 (N_38631,N_38154,N_38175);
xnor U38632 (N_38632,N_38072,N_38484);
or U38633 (N_38633,N_38364,N_38481);
and U38634 (N_38634,N_38157,N_38220);
or U38635 (N_38635,N_38445,N_38349);
nand U38636 (N_38636,N_38421,N_38396);
or U38637 (N_38637,N_38325,N_38088);
nor U38638 (N_38638,N_38436,N_38108);
nand U38639 (N_38639,N_38221,N_38261);
xnor U38640 (N_38640,N_38152,N_38094);
nor U38641 (N_38641,N_38442,N_38315);
nand U38642 (N_38642,N_38003,N_38281);
nor U38643 (N_38643,N_38015,N_38440);
nor U38644 (N_38644,N_38184,N_38139);
xnor U38645 (N_38645,N_38370,N_38302);
xor U38646 (N_38646,N_38448,N_38352);
nor U38647 (N_38647,N_38494,N_38080);
and U38648 (N_38648,N_38135,N_38332);
nor U38649 (N_38649,N_38376,N_38115);
and U38650 (N_38650,N_38290,N_38100);
nand U38651 (N_38651,N_38255,N_38213);
xnor U38652 (N_38652,N_38326,N_38233);
xor U38653 (N_38653,N_38377,N_38177);
or U38654 (N_38654,N_38444,N_38284);
nor U38655 (N_38655,N_38374,N_38307);
and U38656 (N_38656,N_38083,N_38141);
nor U38657 (N_38657,N_38035,N_38405);
xnor U38658 (N_38658,N_38214,N_38424);
nor U38659 (N_38659,N_38306,N_38282);
nand U38660 (N_38660,N_38275,N_38447);
and U38661 (N_38661,N_38441,N_38389);
or U38662 (N_38662,N_38019,N_38124);
nor U38663 (N_38663,N_38132,N_38178);
or U38664 (N_38664,N_38210,N_38316);
xnor U38665 (N_38665,N_38425,N_38417);
nor U38666 (N_38666,N_38314,N_38069);
nand U38667 (N_38667,N_38227,N_38358);
nor U38668 (N_38668,N_38486,N_38495);
nand U38669 (N_38669,N_38194,N_38078);
nand U38670 (N_38670,N_38443,N_38224);
xnor U38671 (N_38671,N_38076,N_38248);
nor U38672 (N_38672,N_38474,N_38329);
nor U38673 (N_38673,N_38053,N_38423);
nand U38674 (N_38674,N_38388,N_38131);
nand U38675 (N_38675,N_38142,N_38007);
nor U38676 (N_38676,N_38464,N_38286);
xor U38677 (N_38677,N_38161,N_38254);
xnor U38678 (N_38678,N_38174,N_38249);
nand U38679 (N_38679,N_38231,N_38006);
xor U38680 (N_38680,N_38446,N_38362);
nor U38681 (N_38681,N_38054,N_38029);
and U38682 (N_38682,N_38268,N_38385);
xor U38683 (N_38683,N_38407,N_38415);
xnor U38684 (N_38684,N_38387,N_38293);
nand U38685 (N_38685,N_38211,N_38206);
xnor U38686 (N_38686,N_38034,N_38127);
or U38687 (N_38687,N_38373,N_38285);
nand U38688 (N_38688,N_38092,N_38199);
and U38689 (N_38689,N_38163,N_38367);
and U38690 (N_38690,N_38002,N_38496);
and U38691 (N_38691,N_38342,N_38283);
and U38692 (N_38692,N_38017,N_38200);
or U38693 (N_38693,N_38382,N_38123);
nand U38694 (N_38694,N_38202,N_38485);
nor U38695 (N_38695,N_38457,N_38119);
xnor U38696 (N_38696,N_38075,N_38093);
and U38697 (N_38697,N_38312,N_38155);
nand U38698 (N_38698,N_38062,N_38140);
nor U38699 (N_38699,N_38433,N_38071);
nand U38700 (N_38700,N_38151,N_38234);
xor U38701 (N_38701,N_38338,N_38260);
or U38702 (N_38702,N_38158,N_38398);
xor U38703 (N_38703,N_38012,N_38330);
xnor U38704 (N_38704,N_38147,N_38288);
xor U38705 (N_38705,N_38065,N_38245);
nand U38706 (N_38706,N_38348,N_38320);
xor U38707 (N_38707,N_38223,N_38112);
nor U38708 (N_38708,N_38414,N_38355);
or U38709 (N_38709,N_38411,N_38419);
or U38710 (N_38710,N_38009,N_38468);
or U38711 (N_38711,N_38462,N_38188);
nand U38712 (N_38712,N_38335,N_38430);
or U38713 (N_38713,N_38242,N_38267);
or U38714 (N_38714,N_38463,N_38323);
nor U38715 (N_38715,N_38287,N_38365);
or U38716 (N_38716,N_38146,N_38333);
xor U38717 (N_38717,N_38475,N_38187);
nand U38718 (N_38718,N_38014,N_38343);
or U38719 (N_38719,N_38257,N_38328);
or U38720 (N_38720,N_38252,N_38045);
and U38721 (N_38721,N_38148,N_38138);
xnor U38722 (N_38722,N_38167,N_38057);
nor U38723 (N_38723,N_38305,N_38427);
nand U38724 (N_38724,N_38409,N_38105);
or U38725 (N_38725,N_38195,N_38394);
xnor U38726 (N_38726,N_38086,N_38059);
and U38727 (N_38727,N_38008,N_38032);
nor U38728 (N_38728,N_38402,N_38229);
nor U38729 (N_38729,N_38429,N_38277);
xor U38730 (N_38730,N_38294,N_38144);
xor U38731 (N_38731,N_38191,N_38454);
and U38732 (N_38732,N_38098,N_38085);
and U38733 (N_38733,N_38011,N_38435);
xor U38734 (N_38734,N_38497,N_38334);
nor U38735 (N_38735,N_38219,N_38452);
nand U38736 (N_38736,N_38018,N_38209);
nand U38737 (N_38737,N_38354,N_38073);
and U38738 (N_38738,N_38020,N_38434);
nor U38739 (N_38739,N_38162,N_38392);
nor U38740 (N_38740,N_38472,N_38043);
and U38741 (N_38741,N_38344,N_38400);
and U38742 (N_38742,N_38084,N_38416);
nor U38743 (N_38743,N_38399,N_38041);
and U38744 (N_38744,N_38418,N_38182);
nand U38745 (N_38745,N_38460,N_38240);
or U38746 (N_38746,N_38378,N_38296);
nor U38747 (N_38747,N_38128,N_38477);
or U38748 (N_38748,N_38130,N_38176);
nor U38749 (N_38749,N_38467,N_38266);
or U38750 (N_38750,N_38282,N_38255);
nand U38751 (N_38751,N_38260,N_38226);
and U38752 (N_38752,N_38205,N_38211);
and U38753 (N_38753,N_38017,N_38280);
nand U38754 (N_38754,N_38358,N_38271);
nor U38755 (N_38755,N_38404,N_38240);
and U38756 (N_38756,N_38447,N_38026);
and U38757 (N_38757,N_38417,N_38381);
nor U38758 (N_38758,N_38033,N_38356);
and U38759 (N_38759,N_38486,N_38150);
or U38760 (N_38760,N_38325,N_38214);
and U38761 (N_38761,N_38363,N_38095);
or U38762 (N_38762,N_38391,N_38263);
or U38763 (N_38763,N_38241,N_38122);
or U38764 (N_38764,N_38291,N_38220);
nand U38765 (N_38765,N_38262,N_38078);
and U38766 (N_38766,N_38221,N_38488);
and U38767 (N_38767,N_38269,N_38394);
nand U38768 (N_38768,N_38354,N_38389);
nor U38769 (N_38769,N_38023,N_38242);
nor U38770 (N_38770,N_38109,N_38348);
xor U38771 (N_38771,N_38412,N_38217);
and U38772 (N_38772,N_38431,N_38078);
or U38773 (N_38773,N_38410,N_38066);
xor U38774 (N_38774,N_38128,N_38243);
nand U38775 (N_38775,N_38094,N_38403);
or U38776 (N_38776,N_38330,N_38167);
nand U38777 (N_38777,N_38064,N_38282);
nand U38778 (N_38778,N_38420,N_38406);
xnor U38779 (N_38779,N_38051,N_38304);
nand U38780 (N_38780,N_38340,N_38488);
xor U38781 (N_38781,N_38187,N_38319);
and U38782 (N_38782,N_38267,N_38442);
or U38783 (N_38783,N_38154,N_38342);
nor U38784 (N_38784,N_38099,N_38172);
nor U38785 (N_38785,N_38011,N_38236);
xnor U38786 (N_38786,N_38068,N_38337);
nand U38787 (N_38787,N_38177,N_38151);
and U38788 (N_38788,N_38031,N_38025);
or U38789 (N_38789,N_38151,N_38436);
xnor U38790 (N_38790,N_38070,N_38443);
nor U38791 (N_38791,N_38311,N_38467);
nand U38792 (N_38792,N_38059,N_38301);
or U38793 (N_38793,N_38064,N_38115);
nand U38794 (N_38794,N_38147,N_38353);
or U38795 (N_38795,N_38311,N_38438);
xor U38796 (N_38796,N_38447,N_38346);
nor U38797 (N_38797,N_38269,N_38315);
nor U38798 (N_38798,N_38111,N_38424);
nor U38799 (N_38799,N_38174,N_38025);
nand U38800 (N_38800,N_38161,N_38166);
or U38801 (N_38801,N_38054,N_38124);
nor U38802 (N_38802,N_38067,N_38476);
nand U38803 (N_38803,N_38073,N_38246);
and U38804 (N_38804,N_38131,N_38096);
nor U38805 (N_38805,N_38431,N_38185);
nand U38806 (N_38806,N_38043,N_38079);
and U38807 (N_38807,N_38415,N_38014);
or U38808 (N_38808,N_38472,N_38019);
xnor U38809 (N_38809,N_38073,N_38142);
or U38810 (N_38810,N_38190,N_38273);
nand U38811 (N_38811,N_38416,N_38370);
xnor U38812 (N_38812,N_38314,N_38343);
xnor U38813 (N_38813,N_38225,N_38397);
nand U38814 (N_38814,N_38100,N_38484);
xnor U38815 (N_38815,N_38266,N_38267);
or U38816 (N_38816,N_38130,N_38269);
nor U38817 (N_38817,N_38237,N_38135);
nand U38818 (N_38818,N_38006,N_38137);
nand U38819 (N_38819,N_38170,N_38234);
nand U38820 (N_38820,N_38442,N_38271);
nand U38821 (N_38821,N_38454,N_38486);
nor U38822 (N_38822,N_38438,N_38312);
xnor U38823 (N_38823,N_38478,N_38323);
and U38824 (N_38824,N_38427,N_38413);
xor U38825 (N_38825,N_38408,N_38463);
nor U38826 (N_38826,N_38348,N_38138);
nor U38827 (N_38827,N_38394,N_38084);
nand U38828 (N_38828,N_38314,N_38392);
nand U38829 (N_38829,N_38498,N_38074);
nand U38830 (N_38830,N_38080,N_38432);
nand U38831 (N_38831,N_38497,N_38441);
nor U38832 (N_38832,N_38420,N_38339);
nand U38833 (N_38833,N_38160,N_38373);
nand U38834 (N_38834,N_38493,N_38306);
nand U38835 (N_38835,N_38131,N_38260);
xnor U38836 (N_38836,N_38099,N_38058);
xor U38837 (N_38837,N_38193,N_38369);
xnor U38838 (N_38838,N_38196,N_38274);
xor U38839 (N_38839,N_38330,N_38290);
xnor U38840 (N_38840,N_38194,N_38026);
and U38841 (N_38841,N_38017,N_38178);
or U38842 (N_38842,N_38271,N_38284);
and U38843 (N_38843,N_38290,N_38303);
or U38844 (N_38844,N_38072,N_38143);
xor U38845 (N_38845,N_38050,N_38360);
and U38846 (N_38846,N_38344,N_38014);
xnor U38847 (N_38847,N_38373,N_38191);
nand U38848 (N_38848,N_38331,N_38426);
nand U38849 (N_38849,N_38312,N_38102);
or U38850 (N_38850,N_38284,N_38069);
nand U38851 (N_38851,N_38435,N_38419);
and U38852 (N_38852,N_38470,N_38467);
nor U38853 (N_38853,N_38269,N_38461);
or U38854 (N_38854,N_38045,N_38234);
and U38855 (N_38855,N_38345,N_38282);
nand U38856 (N_38856,N_38491,N_38339);
or U38857 (N_38857,N_38480,N_38000);
xnor U38858 (N_38858,N_38161,N_38018);
and U38859 (N_38859,N_38195,N_38162);
nand U38860 (N_38860,N_38496,N_38489);
or U38861 (N_38861,N_38356,N_38283);
and U38862 (N_38862,N_38170,N_38220);
xnor U38863 (N_38863,N_38139,N_38460);
nor U38864 (N_38864,N_38202,N_38326);
nor U38865 (N_38865,N_38199,N_38336);
nor U38866 (N_38866,N_38428,N_38411);
xnor U38867 (N_38867,N_38424,N_38227);
or U38868 (N_38868,N_38382,N_38268);
xnor U38869 (N_38869,N_38127,N_38185);
nand U38870 (N_38870,N_38113,N_38348);
xor U38871 (N_38871,N_38372,N_38039);
or U38872 (N_38872,N_38437,N_38444);
and U38873 (N_38873,N_38271,N_38376);
nor U38874 (N_38874,N_38324,N_38139);
nand U38875 (N_38875,N_38366,N_38478);
xnor U38876 (N_38876,N_38155,N_38006);
and U38877 (N_38877,N_38009,N_38459);
xor U38878 (N_38878,N_38272,N_38488);
and U38879 (N_38879,N_38348,N_38099);
and U38880 (N_38880,N_38082,N_38287);
or U38881 (N_38881,N_38126,N_38235);
or U38882 (N_38882,N_38068,N_38165);
and U38883 (N_38883,N_38427,N_38139);
xor U38884 (N_38884,N_38323,N_38394);
nand U38885 (N_38885,N_38257,N_38393);
nor U38886 (N_38886,N_38129,N_38409);
xor U38887 (N_38887,N_38423,N_38001);
xnor U38888 (N_38888,N_38350,N_38130);
nor U38889 (N_38889,N_38380,N_38215);
or U38890 (N_38890,N_38274,N_38388);
nand U38891 (N_38891,N_38096,N_38057);
nand U38892 (N_38892,N_38384,N_38097);
nand U38893 (N_38893,N_38040,N_38488);
and U38894 (N_38894,N_38040,N_38478);
nor U38895 (N_38895,N_38045,N_38321);
nand U38896 (N_38896,N_38032,N_38058);
nand U38897 (N_38897,N_38440,N_38095);
and U38898 (N_38898,N_38423,N_38429);
xnor U38899 (N_38899,N_38289,N_38460);
and U38900 (N_38900,N_38120,N_38425);
nor U38901 (N_38901,N_38171,N_38291);
and U38902 (N_38902,N_38360,N_38284);
nor U38903 (N_38903,N_38431,N_38229);
xor U38904 (N_38904,N_38110,N_38236);
and U38905 (N_38905,N_38020,N_38116);
nand U38906 (N_38906,N_38356,N_38277);
nand U38907 (N_38907,N_38429,N_38192);
and U38908 (N_38908,N_38423,N_38183);
or U38909 (N_38909,N_38000,N_38234);
xor U38910 (N_38910,N_38327,N_38207);
or U38911 (N_38911,N_38323,N_38245);
and U38912 (N_38912,N_38114,N_38317);
nand U38913 (N_38913,N_38244,N_38284);
nor U38914 (N_38914,N_38086,N_38327);
nand U38915 (N_38915,N_38282,N_38081);
nor U38916 (N_38916,N_38159,N_38345);
nor U38917 (N_38917,N_38313,N_38124);
nand U38918 (N_38918,N_38493,N_38011);
and U38919 (N_38919,N_38486,N_38140);
and U38920 (N_38920,N_38447,N_38271);
nor U38921 (N_38921,N_38347,N_38339);
nor U38922 (N_38922,N_38477,N_38311);
nand U38923 (N_38923,N_38435,N_38045);
and U38924 (N_38924,N_38495,N_38422);
xor U38925 (N_38925,N_38261,N_38406);
xor U38926 (N_38926,N_38053,N_38076);
nand U38927 (N_38927,N_38167,N_38149);
or U38928 (N_38928,N_38450,N_38055);
nor U38929 (N_38929,N_38487,N_38436);
or U38930 (N_38930,N_38328,N_38467);
and U38931 (N_38931,N_38199,N_38061);
nand U38932 (N_38932,N_38451,N_38476);
nand U38933 (N_38933,N_38092,N_38164);
nand U38934 (N_38934,N_38458,N_38082);
or U38935 (N_38935,N_38043,N_38236);
nor U38936 (N_38936,N_38065,N_38016);
nor U38937 (N_38937,N_38013,N_38108);
nand U38938 (N_38938,N_38243,N_38265);
xnor U38939 (N_38939,N_38475,N_38416);
and U38940 (N_38940,N_38382,N_38338);
or U38941 (N_38941,N_38060,N_38351);
nor U38942 (N_38942,N_38291,N_38215);
xor U38943 (N_38943,N_38072,N_38032);
nor U38944 (N_38944,N_38120,N_38220);
xnor U38945 (N_38945,N_38190,N_38453);
and U38946 (N_38946,N_38227,N_38152);
nor U38947 (N_38947,N_38080,N_38004);
or U38948 (N_38948,N_38055,N_38194);
nand U38949 (N_38949,N_38197,N_38450);
or U38950 (N_38950,N_38289,N_38028);
and U38951 (N_38951,N_38062,N_38197);
and U38952 (N_38952,N_38132,N_38006);
or U38953 (N_38953,N_38093,N_38066);
nor U38954 (N_38954,N_38154,N_38262);
xor U38955 (N_38955,N_38252,N_38231);
nand U38956 (N_38956,N_38485,N_38473);
nand U38957 (N_38957,N_38031,N_38466);
nand U38958 (N_38958,N_38390,N_38064);
nor U38959 (N_38959,N_38241,N_38032);
xnor U38960 (N_38960,N_38396,N_38321);
or U38961 (N_38961,N_38167,N_38267);
and U38962 (N_38962,N_38029,N_38270);
and U38963 (N_38963,N_38297,N_38042);
nand U38964 (N_38964,N_38193,N_38491);
xor U38965 (N_38965,N_38007,N_38392);
nand U38966 (N_38966,N_38252,N_38369);
nor U38967 (N_38967,N_38248,N_38305);
or U38968 (N_38968,N_38270,N_38430);
nand U38969 (N_38969,N_38130,N_38160);
nor U38970 (N_38970,N_38386,N_38276);
nor U38971 (N_38971,N_38446,N_38074);
xor U38972 (N_38972,N_38071,N_38044);
nor U38973 (N_38973,N_38270,N_38378);
xnor U38974 (N_38974,N_38098,N_38040);
or U38975 (N_38975,N_38457,N_38239);
or U38976 (N_38976,N_38260,N_38386);
xor U38977 (N_38977,N_38332,N_38251);
or U38978 (N_38978,N_38457,N_38070);
or U38979 (N_38979,N_38375,N_38199);
nor U38980 (N_38980,N_38247,N_38313);
and U38981 (N_38981,N_38130,N_38236);
and U38982 (N_38982,N_38002,N_38058);
or U38983 (N_38983,N_38488,N_38381);
and U38984 (N_38984,N_38026,N_38369);
nand U38985 (N_38985,N_38383,N_38014);
and U38986 (N_38986,N_38287,N_38065);
or U38987 (N_38987,N_38182,N_38453);
nor U38988 (N_38988,N_38167,N_38415);
xor U38989 (N_38989,N_38002,N_38484);
xor U38990 (N_38990,N_38112,N_38113);
or U38991 (N_38991,N_38330,N_38259);
and U38992 (N_38992,N_38140,N_38135);
and U38993 (N_38993,N_38074,N_38492);
nor U38994 (N_38994,N_38446,N_38042);
or U38995 (N_38995,N_38072,N_38144);
nand U38996 (N_38996,N_38291,N_38032);
nor U38997 (N_38997,N_38431,N_38158);
and U38998 (N_38998,N_38053,N_38253);
or U38999 (N_38999,N_38359,N_38084);
and U39000 (N_39000,N_38886,N_38595);
or U39001 (N_39001,N_38537,N_38619);
nand U39002 (N_39002,N_38572,N_38573);
xnor U39003 (N_39003,N_38753,N_38790);
xor U39004 (N_39004,N_38629,N_38877);
or U39005 (N_39005,N_38838,N_38749);
nor U39006 (N_39006,N_38531,N_38785);
and U39007 (N_39007,N_38897,N_38824);
nand U39008 (N_39008,N_38518,N_38647);
nand U39009 (N_39009,N_38942,N_38501);
nor U39010 (N_39010,N_38937,N_38664);
xnor U39011 (N_39011,N_38624,N_38744);
or U39012 (N_39012,N_38894,N_38740);
and U39013 (N_39013,N_38934,N_38657);
nor U39014 (N_39014,N_38812,N_38507);
nand U39015 (N_39015,N_38515,N_38636);
nand U39016 (N_39016,N_38644,N_38728);
and U39017 (N_39017,N_38993,N_38530);
or U39018 (N_39018,N_38848,N_38618);
and U39019 (N_39019,N_38841,N_38856);
nand U39020 (N_39020,N_38820,N_38589);
nor U39021 (N_39021,N_38638,N_38954);
or U39022 (N_39022,N_38566,N_38750);
xnor U39023 (N_39023,N_38581,N_38852);
xor U39024 (N_39024,N_38959,N_38569);
or U39025 (N_39025,N_38722,N_38688);
and U39026 (N_39026,N_38985,N_38796);
nor U39027 (N_39027,N_38522,N_38693);
or U39028 (N_39028,N_38694,N_38761);
nor U39029 (N_39029,N_38822,N_38900);
or U39030 (N_39030,N_38653,N_38945);
or U39031 (N_39031,N_38803,N_38818);
and U39032 (N_39032,N_38873,N_38550);
nand U39033 (N_39033,N_38703,N_38777);
nand U39034 (N_39034,N_38545,N_38743);
xnor U39035 (N_39035,N_38633,N_38971);
xnor U39036 (N_39036,N_38964,N_38516);
or U39037 (N_39037,N_38755,N_38650);
or U39038 (N_39038,N_38720,N_38963);
and U39039 (N_39039,N_38560,N_38599);
xor U39040 (N_39040,N_38865,N_38682);
xnor U39041 (N_39041,N_38733,N_38787);
or U39042 (N_39042,N_38527,N_38604);
or U39043 (N_39043,N_38860,N_38536);
or U39044 (N_39044,N_38692,N_38977);
nand U39045 (N_39045,N_38605,N_38730);
xnor U39046 (N_39046,N_38882,N_38980);
or U39047 (N_39047,N_38649,N_38794);
nor U39048 (N_39048,N_38994,N_38760);
nor U39049 (N_39049,N_38738,N_38764);
and U39050 (N_39050,N_38811,N_38885);
and U39051 (N_39051,N_38817,N_38890);
xnor U39052 (N_39052,N_38992,N_38702);
nand U39053 (N_39053,N_38867,N_38783);
nand U39054 (N_39054,N_38815,N_38514);
xnor U39055 (N_39055,N_38806,N_38565);
and U39056 (N_39056,N_38614,N_38928);
nand U39057 (N_39057,N_38758,N_38641);
or U39058 (N_39058,N_38902,N_38616);
and U39059 (N_39059,N_38621,N_38791);
or U39060 (N_39060,N_38823,N_38912);
or U39061 (N_39061,N_38906,N_38691);
xor U39062 (N_39062,N_38668,N_38947);
and U39063 (N_39063,N_38524,N_38962);
nor U39064 (N_39064,N_38667,N_38996);
nand U39065 (N_39065,N_38632,N_38951);
or U39066 (N_39066,N_38930,N_38591);
or U39067 (N_39067,N_38800,N_38946);
and U39068 (N_39068,N_38982,N_38975);
nand U39069 (N_39069,N_38613,N_38686);
xor U39070 (N_39070,N_38768,N_38935);
nor U39071 (N_39071,N_38568,N_38779);
xnor U39072 (N_39072,N_38874,N_38825);
nand U39073 (N_39073,N_38797,N_38799);
nand U39074 (N_39074,N_38503,N_38917);
nand U39075 (N_39075,N_38948,N_38695);
nor U39076 (N_39076,N_38655,N_38725);
xnor U39077 (N_39077,N_38802,N_38956);
xnor U39078 (N_39078,N_38659,N_38561);
or U39079 (N_39079,N_38711,N_38924);
nand U39080 (N_39080,N_38795,N_38741);
or U39081 (N_39081,N_38871,N_38850);
and U39082 (N_39082,N_38685,N_38634);
xor U39083 (N_39083,N_38875,N_38615);
nor U39084 (N_39084,N_38533,N_38859);
nand U39085 (N_39085,N_38835,N_38723);
nand U39086 (N_39086,N_38721,N_38814);
nor U39087 (N_39087,N_38757,N_38654);
and U39088 (N_39088,N_38774,N_38969);
nand U39089 (N_39089,N_38767,N_38889);
and U39090 (N_39090,N_38652,N_38562);
nor U39091 (N_39091,N_38517,N_38829);
or U39092 (N_39092,N_38913,N_38832);
xnor U39093 (N_39093,N_38710,N_38775);
xor U39094 (N_39094,N_38953,N_38706);
nor U39095 (N_39095,N_38771,N_38549);
and U39096 (N_39096,N_38714,N_38669);
nor U39097 (N_39097,N_38580,N_38929);
nor U39098 (N_39098,N_38781,N_38736);
or U39099 (N_39099,N_38923,N_38862);
xor U39100 (N_39100,N_38888,N_38986);
and U39101 (N_39101,N_38567,N_38610);
nor U39102 (N_39102,N_38950,N_38826);
nand U39103 (N_39103,N_38600,N_38601);
and U39104 (N_39104,N_38520,N_38548);
xnor U39105 (N_39105,N_38833,N_38784);
nor U39106 (N_39106,N_38509,N_38671);
xor U39107 (N_39107,N_38938,N_38602);
xor U39108 (N_39108,N_38708,N_38645);
or U39109 (N_39109,N_38675,N_38915);
or U39110 (N_39110,N_38626,N_38592);
or U39111 (N_39111,N_38680,N_38981);
nand U39112 (N_39112,N_38635,N_38926);
nor U39113 (N_39113,N_38907,N_38807);
or U39114 (N_39114,N_38553,N_38842);
nand U39115 (N_39115,N_38958,N_38961);
nor U39116 (N_39116,N_38861,N_38909);
or U39117 (N_39117,N_38539,N_38792);
or U39118 (N_39118,N_38870,N_38968);
and U39119 (N_39119,N_38662,N_38831);
xnor U39120 (N_39120,N_38704,N_38908);
and U39121 (N_39121,N_38979,N_38991);
nand U39122 (N_39122,N_38804,N_38925);
nand U39123 (N_39123,N_38656,N_38574);
and U39124 (N_39124,N_38513,N_38866);
and U39125 (N_39125,N_38511,N_38701);
or U39126 (N_39126,N_38663,N_38816);
xnor U39127 (N_39127,N_38544,N_38739);
xor U39128 (N_39128,N_38960,N_38727);
and U39129 (N_39129,N_38555,N_38878);
and U39130 (N_39130,N_38830,N_38696);
and U39131 (N_39131,N_38598,N_38504);
nand U39132 (N_39132,N_38640,N_38508);
or U39133 (N_39133,N_38526,N_38851);
and U39134 (N_39134,N_38809,N_38563);
and U39135 (N_39135,N_38987,N_38998);
nand U39136 (N_39136,N_38609,N_38919);
and U39137 (N_39137,N_38528,N_38944);
and U39138 (N_39138,N_38612,N_38939);
nor U39139 (N_39139,N_38898,N_38678);
xor U39140 (N_39140,N_38868,N_38745);
nand U39141 (N_39141,N_38596,N_38690);
xnor U39142 (N_39142,N_38782,N_38765);
or U39143 (N_39143,N_38952,N_38810);
nor U39144 (N_39144,N_38903,N_38532);
or U39145 (N_39145,N_38525,N_38546);
nor U39146 (N_39146,N_38697,N_38978);
nor U39147 (N_39147,N_38763,N_38506);
nand U39148 (N_39148,N_38715,N_38689);
or U39149 (N_39149,N_38941,N_38705);
nor U39150 (N_39150,N_38995,N_38554);
nor U39151 (N_39151,N_38651,N_38769);
nand U39152 (N_39152,N_38583,N_38737);
xnor U39153 (N_39153,N_38735,N_38780);
and U39154 (N_39154,N_38786,N_38731);
nor U39155 (N_39155,N_38707,N_38932);
xnor U39156 (N_39156,N_38990,N_38788);
nor U39157 (N_39157,N_38857,N_38827);
nand U39158 (N_39158,N_38687,N_38872);
nand U39159 (N_39159,N_38716,N_38772);
xor U39160 (N_39160,N_38608,N_38603);
nand U39161 (N_39161,N_38869,N_38793);
xnor U39162 (N_39162,N_38754,N_38984);
or U39163 (N_39163,N_38564,N_38893);
nor U39164 (N_39164,N_38502,N_38684);
nand U39165 (N_39165,N_38983,N_38557);
and U39166 (N_39166,N_38660,N_38798);
nand U39167 (N_39167,N_38597,N_38551);
or U39168 (N_39168,N_38679,N_38789);
or U39169 (N_39169,N_38940,N_38931);
nand U39170 (N_39170,N_38673,N_38805);
or U39171 (N_39171,N_38876,N_38746);
nor U39172 (N_39172,N_38523,N_38911);
or U39173 (N_39173,N_38665,N_38698);
or U39174 (N_39174,N_38813,N_38547);
xor U39175 (N_39175,N_38594,N_38582);
and U39176 (N_39176,N_38970,N_38578);
nor U39177 (N_39177,N_38751,N_38719);
nand U39178 (N_39178,N_38521,N_38834);
or U39179 (N_39179,N_38606,N_38748);
or U39180 (N_39180,N_38623,N_38855);
and U39181 (N_39181,N_38974,N_38639);
xor U39182 (N_39182,N_38839,N_38895);
xnor U39183 (N_39183,N_38646,N_38726);
xor U39184 (N_39184,N_38770,N_38622);
nand U39185 (N_39185,N_38676,N_38534);
and U39186 (N_39186,N_38905,N_38590);
xor U39187 (N_39187,N_38752,N_38529);
nor U39188 (N_39188,N_38700,N_38593);
nor U39189 (N_39189,N_38880,N_38648);
or U39190 (N_39190,N_38577,N_38864);
and U39191 (N_39191,N_38519,N_38899);
nand U39192 (N_39192,N_38819,N_38840);
xor U39193 (N_39193,N_38677,N_38747);
nand U39194 (N_39194,N_38957,N_38742);
nand U39195 (N_39195,N_38879,N_38642);
nand U39196 (N_39196,N_38965,N_38828);
or U39197 (N_39197,N_38637,N_38910);
nand U39198 (N_39198,N_38718,N_38922);
and U39199 (N_39199,N_38611,N_38836);
xor U39200 (N_39200,N_38936,N_38584);
or U39201 (N_39201,N_38571,N_38713);
and U39202 (N_39202,N_38552,N_38661);
and U39203 (N_39203,N_38724,N_38844);
or U39204 (N_39204,N_38778,N_38989);
xor U39205 (N_39205,N_38541,N_38588);
nand U39206 (N_39206,N_38625,N_38628);
xor U39207 (N_39207,N_38999,N_38843);
nand U39208 (N_39208,N_38921,N_38955);
nand U39209 (N_39209,N_38883,N_38631);
nor U39210 (N_39210,N_38881,N_38837);
nor U39211 (N_39211,N_38846,N_38556);
xnor U39212 (N_39212,N_38863,N_38579);
and U39213 (N_39213,N_38683,N_38674);
nor U39214 (N_39214,N_38587,N_38933);
nor U39215 (N_39215,N_38808,N_38887);
nor U39216 (N_39216,N_38916,N_38847);
or U39217 (N_39217,N_38670,N_38821);
nor U39218 (N_39218,N_38709,N_38559);
nand U39219 (N_39219,N_38884,N_38505);
nand U39220 (N_39220,N_38801,N_38943);
nand U39221 (N_39221,N_38976,N_38672);
nand U39222 (N_39222,N_38967,N_38845);
nand U39223 (N_39223,N_38949,N_38756);
nor U39224 (N_39224,N_38892,N_38658);
nand U39225 (N_39225,N_38712,N_38558);
nand U39226 (N_39226,N_38627,N_38666);
and U39227 (N_39227,N_38510,N_38540);
xnor U39228 (N_39228,N_38729,N_38500);
xnor U39229 (N_39229,N_38542,N_38585);
and U39230 (N_39230,N_38914,N_38576);
or U39231 (N_39231,N_38891,N_38918);
nand U39232 (N_39232,N_38732,N_38586);
nand U39233 (N_39233,N_38570,N_38988);
xnor U39234 (N_39234,N_38997,N_38901);
or U39235 (N_39235,N_38630,N_38512);
or U39236 (N_39236,N_38973,N_38896);
and U39237 (N_39237,N_38543,N_38762);
and U39238 (N_39238,N_38699,N_38904);
nor U39239 (N_39239,N_38643,N_38966);
and U39240 (N_39240,N_38776,N_38858);
xor U39241 (N_39241,N_38849,N_38617);
nand U39242 (N_39242,N_38972,N_38681);
nor U39243 (N_39243,N_38620,N_38759);
and U39244 (N_39244,N_38766,N_38535);
or U39245 (N_39245,N_38853,N_38854);
or U39246 (N_39246,N_38717,N_38927);
nor U39247 (N_39247,N_38607,N_38538);
xnor U39248 (N_39248,N_38734,N_38575);
or U39249 (N_39249,N_38920,N_38773);
nand U39250 (N_39250,N_38736,N_38858);
xor U39251 (N_39251,N_38801,N_38550);
xnor U39252 (N_39252,N_38671,N_38632);
nor U39253 (N_39253,N_38823,N_38900);
and U39254 (N_39254,N_38911,N_38991);
and U39255 (N_39255,N_38863,N_38733);
nand U39256 (N_39256,N_38556,N_38607);
nor U39257 (N_39257,N_38601,N_38695);
nor U39258 (N_39258,N_38534,N_38998);
and U39259 (N_39259,N_38932,N_38523);
xor U39260 (N_39260,N_38762,N_38779);
and U39261 (N_39261,N_38885,N_38791);
nor U39262 (N_39262,N_38521,N_38684);
or U39263 (N_39263,N_38658,N_38946);
or U39264 (N_39264,N_38970,N_38816);
xnor U39265 (N_39265,N_38787,N_38849);
or U39266 (N_39266,N_38714,N_38757);
nand U39267 (N_39267,N_38715,N_38792);
nor U39268 (N_39268,N_38851,N_38911);
or U39269 (N_39269,N_38699,N_38885);
or U39270 (N_39270,N_38665,N_38626);
xnor U39271 (N_39271,N_38851,N_38828);
or U39272 (N_39272,N_38936,N_38958);
nand U39273 (N_39273,N_38957,N_38741);
xnor U39274 (N_39274,N_38703,N_38636);
or U39275 (N_39275,N_38936,N_38727);
and U39276 (N_39276,N_38684,N_38600);
xnor U39277 (N_39277,N_38530,N_38501);
and U39278 (N_39278,N_38685,N_38713);
or U39279 (N_39279,N_38748,N_38820);
and U39280 (N_39280,N_38676,N_38526);
nor U39281 (N_39281,N_38954,N_38844);
xor U39282 (N_39282,N_38954,N_38947);
nand U39283 (N_39283,N_38632,N_38551);
nor U39284 (N_39284,N_38953,N_38514);
nand U39285 (N_39285,N_38623,N_38578);
and U39286 (N_39286,N_38781,N_38843);
nor U39287 (N_39287,N_38843,N_38857);
or U39288 (N_39288,N_38760,N_38960);
or U39289 (N_39289,N_38753,N_38539);
nand U39290 (N_39290,N_38941,N_38590);
nor U39291 (N_39291,N_38878,N_38743);
nor U39292 (N_39292,N_38874,N_38901);
xnor U39293 (N_39293,N_38503,N_38951);
and U39294 (N_39294,N_38547,N_38722);
and U39295 (N_39295,N_38746,N_38629);
and U39296 (N_39296,N_38895,N_38945);
nand U39297 (N_39297,N_38937,N_38533);
nor U39298 (N_39298,N_38914,N_38730);
nand U39299 (N_39299,N_38504,N_38858);
or U39300 (N_39300,N_38868,N_38727);
and U39301 (N_39301,N_38612,N_38655);
nor U39302 (N_39302,N_38763,N_38942);
or U39303 (N_39303,N_38999,N_38735);
nor U39304 (N_39304,N_38729,N_38872);
nor U39305 (N_39305,N_38914,N_38503);
nand U39306 (N_39306,N_38757,N_38517);
nor U39307 (N_39307,N_38570,N_38620);
and U39308 (N_39308,N_38840,N_38805);
xor U39309 (N_39309,N_38989,N_38654);
xor U39310 (N_39310,N_38647,N_38795);
nor U39311 (N_39311,N_38906,N_38773);
nor U39312 (N_39312,N_38519,N_38997);
and U39313 (N_39313,N_38942,N_38776);
nand U39314 (N_39314,N_38807,N_38646);
and U39315 (N_39315,N_38863,N_38768);
nor U39316 (N_39316,N_38930,N_38949);
xor U39317 (N_39317,N_38512,N_38876);
and U39318 (N_39318,N_38995,N_38613);
xor U39319 (N_39319,N_38732,N_38607);
nor U39320 (N_39320,N_38550,N_38551);
nand U39321 (N_39321,N_38574,N_38772);
nor U39322 (N_39322,N_38896,N_38670);
nand U39323 (N_39323,N_38688,N_38842);
and U39324 (N_39324,N_38892,N_38765);
nand U39325 (N_39325,N_38804,N_38769);
and U39326 (N_39326,N_38866,N_38771);
nor U39327 (N_39327,N_38604,N_38747);
and U39328 (N_39328,N_38834,N_38542);
or U39329 (N_39329,N_38846,N_38850);
or U39330 (N_39330,N_38904,N_38738);
xor U39331 (N_39331,N_38700,N_38694);
xor U39332 (N_39332,N_38960,N_38612);
or U39333 (N_39333,N_38763,N_38730);
and U39334 (N_39334,N_38692,N_38956);
nor U39335 (N_39335,N_38630,N_38559);
xor U39336 (N_39336,N_38981,N_38716);
and U39337 (N_39337,N_38987,N_38548);
xnor U39338 (N_39338,N_38925,N_38791);
xor U39339 (N_39339,N_38868,N_38592);
nand U39340 (N_39340,N_38679,N_38585);
or U39341 (N_39341,N_38688,N_38726);
or U39342 (N_39342,N_38572,N_38773);
nor U39343 (N_39343,N_38681,N_38651);
or U39344 (N_39344,N_38603,N_38657);
xor U39345 (N_39345,N_38846,N_38920);
or U39346 (N_39346,N_38629,N_38884);
nor U39347 (N_39347,N_38989,N_38824);
xnor U39348 (N_39348,N_38827,N_38734);
xor U39349 (N_39349,N_38999,N_38827);
xor U39350 (N_39350,N_38862,N_38652);
nor U39351 (N_39351,N_38659,N_38600);
nor U39352 (N_39352,N_38558,N_38665);
or U39353 (N_39353,N_38695,N_38815);
nor U39354 (N_39354,N_38835,N_38952);
and U39355 (N_39355,N_38856,N_38975);
nor U39356 (N_39356,N_38732,N_38780);
xnor U39357 (N_39357,N_38645,N_38846);
xnor U39358 (N_39358,N_38955,N_38956);
nor U39359 (N_39359,N_38811,N_38845);
or U39360 (N_39360,N_38590,N_38942);
nand U39361 (N_39361,N_38869,N_38687);
nor U39362 (N_39362,N_38722,N_38701);
xor U39363 (N_39363,N_38763,N_38529);
nor U39364 (N_39364,N_38646,N_38937);
or U39365 (N_39365,N_38735,N_38917);
and U39366 (N_39366,N_38755,N_38524);
nand U39367 (N_39367,N_38558,N_38836);
nor U39368 (N_39368,N_38720,N_38681);
nand U39369 (N_39369,N_38703,N_38591);
or U39370 (N_39370,N_38673,N_38501);
xnor U39371 (N_39371,N_38521,N_38851);
xnor U39372 (N_39372,N_38549,N_38812);
nand U39373 (N_39373,N_38507,N_38895);
nor U39374 (N_39374,N_38755,N_38672);
or U39375 (N_39375,N_38636,N_38586);
nor U39376 (N_39376,N_38910,N_38911);
nor U39377 (N_39377,N_38891,N_38781);
or U39378 (N_39378,N_38722,N_38609);
and U39379 (N_39379,N_38578,N_38850);
and U39380 (N_39380,N_38800,N_38735);
xor U39381 (N_39381,N_38621,N_38961);
or U39382 (N_39382,N_38975,N_38685);
or U39383 (N_39383,N_38738,N_38907);
nor U39384 (N_39384,N_38679,N_38966);
nor U39385 (N_39385,N_38636,N_38540);
nor U39386 (N_39386,N_38531,N_38993);
or U39387 (N_39387,N_38584,N_38689);
xor U39388 (N_39388,N_38826,N_38668);
and U39389 (N_39389,N_38621,N_38510);
nor U39390 (N_39390,N_38760,N_38920);
or U39391 (N_39391,N_38835,N_38895);
and U39392 (N_39392,N_38852,N_38834);
or U39393 (N_39393,N_38875,N_38541);
nor U39394 (N_39394,N_38878,N_38762);
and U39395 (N_39395,N_38945,N_38536);
xnor U39396 (N_39396,N_38983,N_38665);
nor U39397 (N_39397,N_38741,N_38667);
or U39398 (N_39398,N_38903,N_38881);
xnor U39399 (N_39399,N_38908,N_38675);
nand U39400 (N_39400,N_38765,N_38589);
and U39401 (N_39401,N_38645,N_38600);
xnor U39402 (N_39402,N_38531,N_38708);
nor U39403 (N_39403,N_38822,N_38885);
xnor U39404 (N_39404,N_38557,N_38944);
and U39405 (N_39405,N_38528,N_38523);
nand U39406 (N_39406,N_38511,N_38871);
nand U39407 (N_39407,N_38709,N_38554);
and U39408 (N_39408,N_38587,N_38871);
nand U39409 (N_39409,N_38520,N_38806);
xor U39410 (N_39410,N_38536,N_38818);
or U39411 (N_39411,N_38760,N_38692);
nor U39412 (N_39412,N_38657,N_38621);
and U39413 (N_39413,N_38772,N_38691);
or U39414 (N_39414,N_38545,N_38672);
nand U39415 (N_39415,N_38511,N_38866);
nand U39416 (N_39416,N_38842,N_38871);
nor U39417 (N_39417,N_38604,N_38739);
or U39418 (N_39418,N_38573,N_38509);
and U39419 (N_39419,N_38645,N_38781);
nor U39420 (N_39420,N_38738,N_38888);
xnor U39421 (N_39421,N_38940,N_38509);
nor U39422 (N_39422,N_38749,N_38616);
nor U39423 (N_39423,N_38607,N_38736);
or U39424 (N_39424,N_38804,N_38533);
nand U39425 (N_39425,N_38795,N_38826);
nor U39426 (N_39426,N_38645,N_38881);
and U39427 (N_39427,N_38591,N_38543);
nand U39428 (N_39428,N_38555,N_38723);
and U39429 (N_39429,N_38830,N_38621);
and U39430 (N_39430,N_38848,N_38786);
nand U39431 (N_39431,N_38642,N_38651);
and U39432 (N_39432,N_38855,N_38688);
and U39433 (N_39433,N_38958,N_38752);
and U39434 (N_39434,N_38608,N_38634);
nor U39435 (N_39435,N_38999,N_38769);
or U39436 (N_39436,N_38806,N_38992);
and U39437 (N_39437,N_38695,N_38609);
xor U39438 (N_39438,N_38624,N_38534);
xor U39439 (N_39439,N_38672,N_38701);
and U39440 (N_39440,N_38588,N_38900);
or U39441 (N_39441,N_38667,N_38901);
and U39442 (N_39442,N_38970,N_38811);
xnor U39443 (N_39443,N_38965,N_38652);
and U39444 (N_39444,N_38817,N_38819);
or U39445 (N_39445,N_38903,N_38748);
or U39446 (N_39446,N_38823,N_38643);
nor U39447 (N_39447,N_38784,N_38510);
or U39448 (N_39448,N_38959,N_38934);
xor U39449 (N_39449,N_38511,N_38897);
nand U39450 (N_39450,N_38683,N_38699);
and U39451 (N_39451,N_38733,N_38565);
or U39452 (N_39452,N_38923,N_38560);
nor U39453 (N_39453,N_38978,N_38928);
or U39454 (N_39454,N_38661,N_38651);
nor U39455 (N_39455,N_38720,N_38621);
and U39456 (N_39456,N_38904,N_38824);
or U39457 (N_39457,N_38984,N_38911);
xnor U39458 (N_39458,N_38666,N_38543);
nand U39459 (N_39459,N_38850,N_38986);
nand U39460 (N_39460,N_38872,N_38785);
and U39461 (N_39461,N_38563,N_38602);
or U39462 (N_39462,N_38642,N_38571);
xor U39463 (N_39463,N_38658,N_38617);
nand U39464 (N_39464,N_38842,N_38641);
or U39465 (N_39465,N_38832,N_38678);
or U39466 (N_39466,N_38617,N_38521);
and U39467 (N_39467,N_38948,N_38613);
or U39468 (N_39468,N_38970,N_38953);
nand U39469 (N_39469,N_38656,N_38728);
and U39470 (N_39470,N_38551,N_38978);
nor U39471 (N_39471,N_38644,N_38661);
nand U39472 (N_39472,N_38654,N_38501);
and U39473 (N_39473,N_38629,N_38873);
nor U39474 (N_39474,N_38500,N_38856);
nand U39475 (N_39475,N_38997,N_38618);
nand U39476 (N_39476,N_38845,N_38771);
nor U39477 (N_39477,N_38552,N_38731);
and U39478 (N_39478,N_38683,N_38681);
and U39479 (N_39479,N_38539,N_38736);
xnor U39480 (N_39480,N_38690,N_38559);
nor U39481 (N_39481,N_38547,N_38581);
nor U39482 (N_39482,N_38960,N_38773);
or U39483 (N_39483,N_38696,N_38788);
xnor U39484 (N_39484,N_38748,N_38847);
or U39485 (N_39485,N_38839,N_38717);
or U39486 (N_39486,N_38657,N_38748);
xor U39487 (N_39487,N_38843,N_38777);
xor U39488 (N_39488,N_38792,N_38998);
and U39489 (N_39489,N_38811,N_38936);
nand U39490 (N_39490,N_38628,N_38794);
xnor U39491 (N_39491,N_38831,N_38541);
or U39492 (N_39492,N_38936,N_38734);
and U39493 (N_39493,N_38885,N_38819);
and U39494 (N_39494,N_38577,N_38876);
and U39495 (N_39495,N_38823,N_38893);
xor U39496 (N_39496,N_38755,N_38506);
and U39497 (N_39497,N_38784,N_38700);
nor U39498 (N_39498,N_38883,N_38687);
and U39499 (N_39499,N_38904,N_38668);
or U39500 (N_39500,N_39327,N_39252);
xnor U39501 (N_39501,N_39111,N_39463);
or U39502 (N_39502,N_39088,N_39203);
xnor U39503 (N_39503,N_39403,N_39116);
nor U39504 (N_39504,N_39165,N_39396);
and U39505 (N_39505,N_39235,N_39376);
nand U39506 (N_39506,N_39166,N_39206);
and U39507 (N_39507,N_39259,N_39004);
nor U39508 (N_39508,N_39388,N_39082);
or U39509 (N_39509,N_39216,N_39227);
and U39510 (N_39510,N_39373,N_39352);
and U39511 (N_39511,N_39257,N_39431);
and U39512 (N_39512,N_39309,N_39341);
and U39513 (N_39513,N_39021,N_39129);
and U39514 (N_39514,N_39126,N_39127);
nand U39515 (N_39515,N_39387,N_39400);
xor U39516 (N_39516,N_39321,N_39398);
nand U39517 (N_39517,N_39414,N_39083);
and U39518 (N_39518,N_39303,N_39152);
or U39519 (N_39519,N_39307,N_39212);
and U39520 (N_39520,N_39174,N_39093);
nand U39521 (N_39521,N_39356,N_39042);
and U39522 (N_39522,N_39035,N_39416);
nor U39523 (N_39523,N_39099,N_39329);
nand U39524 (N_39524,N_39214,N_39061);
and U39525 (N_39525,N_39399,N_39304);
and U39526 (N_39526,N_39480,N_39181);
and U39527 (N_39527,N_39000,N_39449);
and U39528 (N_39528,N_39448,N_39168);
xor U39529 (N_39529,N_39405,N_39494);
nand U39530 (N_39530,N_39009,N_39043);
nand U39531 (N_39531,N_39192,N_39084);
or U39532 (N_39532,N_39158,N_39490);
nand U39533 (N_39533,N_39051,N_39308);
nor U39534 (N_39534,N_39339,N_39143);
or U39535 (N_39535,N_39036,N_39180);
nor U39536 (N_39536,N_39495,N_39306);
or U39537 (N_39537,N_39250,N_39401);
nand U39538 (N_39538,N_39328,N_39315);
or U39539 (N_39539,N_39270,N_39022);
and U39540 (N_39540,N_39187,N_39440);
nor U39541 (N_39541,N_39207,N_39200);
and U39542 (N_39542,N_39362,N_39185);
nand U39543 (N_39543,N_39027,N_39374);
nand U39544 (N_39544,N_39001,N_39481);
or U39545 (N_39545,N_39242,N_39363);
xor U39546 (N_39546,N_39156,N_39075);
nand U39547 (N_39547,N_39170,N_39380);
or U39548 (N_39548,N_39425,N_39101);
nand U39549 (N_39549,N_39205,N_39058);
and U39550 (N_39550,N_39169,N_39371);
xnor U39551 (N_39551,N_39256,N_39057);
or U39552 (N_39552,N_39369,N_39472);
nand U39553 (N_39553,N_39432,N_39012);
nor U39554 (N_39554,N_39092,N_39062);
and U39555 (N_39555,N_39109,N_39177);
nand U39556 (N_39556,N_39439,N_39367);
nor U39557 (N_39557,N_39199,N_39159);
xnor U39558 (N_39558,N_39137,N_39391);
or U39559 (N_39559,N_39343,N_39118);
and U39560 (N_39560,N_39110,N_39372);
xnor U39561 (N_39561,N_39468,N_39120);
nor U39562 (N_39562,N_39311,N_39213);
or U39563 (N_39563,N_39124,N_39183);
and U39564 (N_39564,N_39247,N_39474);
and U39565 (N_39565,N_39114,N_39332);
nor U39566 (N_39566,N_39263,N_39154);
nor U39567 (N_39567,N_39121,N_39103);
nor U39568 (N_39568,N_39450,N_39473);
nand U39569 (N_39569,N_39335,N_39288);
or U39570 (N_39570,N_39079,N_39067);
nand U39571 (N_39571,N_39316,N_39095);
and U39572 (N_39572,N_39003,N_39064);
and U39573 (N_39573,N_39090,N_39323);
or U39574 (N_39574,N_39423,N_39385);
xor U39575 (N_39575,N_39264,N_39390);
nor U39576 (N_39576,N_39318,N_39469);
and U39577 (N_39577,N_39106,N_39486);
or U39578 (N_39578,N_39119,N_39364);
and U39579 (N_39579,N_39085,N_39146);
or U39580 (N_39580,N_39040,N_39254);
or U39581 (N_39581,N_39453,N_39145);
nand U39582 (N_39582,N_39208,N_39418);
nor U39583 (N_39583,N_39476,N_39066);
nor U39584 (N_39584,N_39383,N_39055);
and U39585 (N_39585,N_39394,N_39324);
nand U39586 (N_39586,N_39457,N_39375);
and U39587 (N_39587,N_39191,N_39193);
nand U39588 (N_39588,N_39301,N_39445);
nand U39589 (N_39589,N_39462,N_39345);
nand U39590 (N_39590,N_39104,N_39144);
nor U39591 (N_39591,N_39413,N_39248);
nor U39592 (N_39592,N_39015,N_39164);
nand U39593 (N_39593,N_39455,N_39297);
or U39594 (N_39594,N_39482,N_39293);
or U39595 (N_39595,N_39132,N_39330);
or U39596 (N_39596,N_39096,N_39005);
xnor U39597 (N_39597,N_39049,N_39081);
or U39598 (N_39598,N_39140,N_39386);
nor U39599 (N_39599,N_39354,N_39342);
and U39600 (N_39600,N_39044,N_39219);
or U39601 (N_39601,N_39404,N_39148);
and U39602 (N_39602,N_39268,N_39086);
or U39603 (N_39603,N_39428,N_39437);
nand U39604 (N_39604,N_39435,N_39115);
nor U39605 (N_39605,N_39267,N_39430);
nand U39606 (N_39606,N_39131,N_39338);
nor U39607 (N_39607,N_39029,N_39229);
or U39608 (N_39608,N_39026,N_39477);
or U39609 (N_39609,N_39278,N_39161);
or U39610 (N_39610,N_39353,N_39417);
nand U39611 (N_39611,N_39107,N_39023);
xnor U39612 (N_39612,N_39382,N_39359);
or U39613 (N_39613,N_39046,N_39179);
or U39614 (N_39614,N_39461,N_39025);
xnor U39615 (N_39615,N_39325,N_39243);
and U39616 (N_39616,N_39237,N_39296);
xnor U39617 (N_39617,N_39034,N_39031);
xor U39618 (N_39618,N_39442,N_39011);
and U39619 (N_39619,N_39077,N_39291);
xnor U39620 (N_39620,N_39286,N_39196);
xor U39621 (N_39621,N_39033,N_39497);
xnor U39622 (N_39622,N_39313,N_39108);
or U39623 (N_39623,N_39251,N_39141);
or U39624 (N_39624,N_39334,N_39253);
xor U39625 (N_39625,N_39028,N_39408);
or U39626 (N_39626,N_39467,N_39456);
and U39627 (N_39627,N_39298,N_39422);
xnor U39628 (N_39628,N_39190,N_39002);
nor U39629 (N_39629,N_39194,N_39326);
nor U39630 (N_39630,N_39420,N_39249);
xor U39631 (N_39631,N_39128,N_39491);
and U39632 (N_39632,N_39117,N_39483);
xnor U39633 (N_39633,N_39322,N_39098);
or U39634 (N_39634,N_39211,N_39138);
nand U39635 (N_39635,N_39224,N_39195);
or U39636 (N_39636,N_39300,N_39451);
nand U39637 (N_39637,N_39393,N_39238);
nand U39638 (N_39638,N_39045,N_39355);
xor U39639 (N_39639,N_39290,N_39361);
nor U39640 (N_39640,N_39007,N_39246);
nor U39641 (N_39641,N_39239,N_39014);
and U39642 (N_39642,N_39032,N_39037);
and U39643 (N_39643,N_39030,N_39410);
nand U39644 (N_39644,N_39424,N_39493);
and U39645 (N_39645,N_39272,N_39038);
and U39646 (N_39646,N_39188,N_39167);
and U39647 (N_39647,N_39094,N_39498);
or U39648 (N_39648,N_39478,N_39142);
nor U39649 (N_39649,N_39366,N_39344);
nand U39650 (N_39650,N_39070,N_39225);
or U39651 (N_39651,N_39265,N_39283);
nor U39652 (N_39652,N_39245,N_39310);
or U39653 (N_39653,N_39172,N_39230);
nor U39654 (N_39654,N_39226,N_39319);
nor U39655 (N_39655,N_39091,N_39411);
and U39656 (N_39656,N_39269,N_39349);
and U39657 (N_39657,N_39302,N_39487);
and U39658 (N_39658,N_39273,N_39184);
or U39659 (N_39659,N_39289,N_39133);
xnor U39660 (N_39660,N_39006,N_39295);
or U39661 (N_39661,N_39065,N_39294);
and U39662 (N_39662,N_39008,N_39053);
xnor U39663 (N_39663,N_39488,N_39266);
xnor U39664 (N_39664,N_39357,N_39047);
xor U39665 (N_39665,N_39470,N_39071);
and U39666 (N_39666,N_39402,N_39360);
or U39667 (N_39667,N_39136,N_39333);
or U39668 (N_39668,N_39466,N_39039);
nand U39669 (N_39669,N_39279,N_39378);
nand U39670 (N_39670,N_39492,N_39441);
xor U39671 (N_39671,N_39056,N_39340);
and U39672 (N_39672,N_39160,N_39073);
xor U39673 (N_39673,N_39351,N_39052);
nand U39674 (N_39674,N_39346,N_39010);
and U39675 (N_39675,N_39149,N_39087);
or U39676 (N_39676,N_39175,N_39421);
or U39677 (N_39677,N_39444,N_39134);
and U39678 (N_39678,N_39178,N_39072);
nand U39679 (N_39679,N_39409,N_39163);
and U39680 (N_39680,N_39048,N_39189);
nand U39681 (N_39681,N_39234,N_39348);
nand U39682 (N_39682,N_39429,N_39013);
nand U39683 (N_39683,N_39292,N_39475);
nand U39684 (N_39684,N_39223,N_39460);
xnor U39685 (N_39685,N_39201,N_39240);
or U39686 (N_39686,N_39016,N_39122);
nand U39687 (N_39687,N_39496,N_39068);
xor U39688 (N_39688,N_39438,N_39317);
xnor U39689 (N_39689,N_39381,N_39287);
or U39690 (N_39690,N_39210,N_39434);
nand U39691 (N_39691,N_39260,N_39222);
xnor U39692 (N_39692,N_39426,N_39060);
and U39693 (N_39693,N_39337,N_39130);
xor U39694 (N_39694,N_39280,N_39489);
and U39695 (N_39695,N_39209,N_39089);
nor U39696 (N_39696,N_39097,N_39078);
or U39697 (N_39697,N_39105,N_39314);
and U39698 (N_39698,N_39282,N_39019);
and U39699 (N_39699,N_39215,N_39198);
xnor U39700 (N_39700,N_39231,N_39244);
xor U39701 (N_39701,N_39471,N_39024);
xnor U39702 (N_39702,N_39059,N_39112);
and U39703 (N_39703,N_39419,N_39299);
nor U39704 (N_39704,N_39074,N_39336);
and U39705 (N_39705,N_39102,N_39312);
nand U39706 (N_39706,N_39204,N_39162);
and U39707 (N_39707,N_39433,N_39135);
and U39708 (N_39708,N_39485,N_39350);
or U39709 (N_39709,N_39173,N_39446);
or U39710 (N_39710,N_39018,N_39241);
nor U39711 (N_39711,N_39465,N_39275);
or U39712 (N_39712,N_39017,N_39384);
nand U39713 (N_39713,N_39202,N_39365);
or U39714 (N_39714,N_39284,N_39368);
or U39715 (N_39715,N_39370,N_39281);
xnor U39716 (N_39716,N_39020,N_39377);
nand U39717 (N_39717,N_39125,N_39186);
nand U39718 (N_39718,N_39262,N_39147);
and U39719 (N_39719,N_39151,N_39320);
and U39720 (N_39720,N_39150,N_39054);
or U39721 (N_39721,N_39447,N_39255);
and U39722 (N_39722,N_39197,N_39080);
or U39723 (N_39723,N_39220,N_39407);
nand U39724 (N_39724,N_39155,N_39221);
nor U39725 (N_39725,N_39258,N_39076);
and U39726 (N_39726,N_39123,N_39458);
nand U39727 (N_39727,N_39443,N_39499);
and U39728 (N_39728,N_39452,N_39415);
nor U39729 (N_39729,N_39397,N_39063);
and U39730 (N_39730,N_39484,N_39276);
and U39731 (N_39731,N_39347,N_39232);
nand U39732 (N_39732,N_39050,N_39412);
nor U39733 (N_39733,N_39285,N_39389);
or U39734 (N_39734,N_39218,N_39113);
or U39735 (N_39735,N_39464,N_39459);
nor U39736 (N_39736,N_39395,N_39331);
or U39737 (N_39737,N_39182,N_39236);
and U39738 (N_39738,N_39406,N_39436);
nor U39739 (N_39739,N_39358,N_39157);
xor U39740 (N_39740,N_39100,N_39153);
nand U39741 (N_39741,N_39479,N_39427);
nor U39742 (N_39742,N_39217,N_39305);
nand U39743 (N_39743,N_39277,N_39392);
and U39744 (N_39744,N_39069,N_39041);
xnor U39745 (N_39745,N_39261,N_39171);
xor U39746 (N_39746,N_39271,N_39274);
or U39747 (N_39747,N_39139,N_39228);
nand U39748 (N_39748,N_39233,N_39176);
or U39749 (N_39749,N_39379,N_39454);
nand U39750 (N_39750,N_39167,N_39001);
nand U39751 (N_39751,N_39035,N_39179);
nor U39752 (N_39752,N_39468,N_39154);
or U39753 (N_39753,N_39426,N_39491);
xor U39754 (N_39754,N_39050,N_39395);
and U39755 (N_39755,N_39413,N_39021);
xor U39756 (N_39756,N_39400,N_39055);
xnor U39757 (N_39757,N_39252,N_39100);
and U39758 (N_39758,N_39416,N_39195);
or U39759 (N_39759,N_39060,N_39281);
or U39760 (N_39760,N_39432,N_39296);
and U39761 (N_39761,N_39192,N_39183);
nand U39762 (N_39762,N_39210,N_39242);
or U39763 (N_39763,N_39215,N_39034);
nor U39764 (N_39764,N_39083,N_39340);
xnor U39765 (N_39765,N_39409,N_39207);
and U39766 (N_39766,N_39229,N_39154);
and U39767 (N_39767,N_39227,N_39071);
or U39768 (N_39768,N_39470,N_39115);
xor U39769 (N_39769,N_39191,N_39079);
xor U39770 (N_39770,N_39027,N_39201);
nor U39771 (N_39771,N_39199,N_39176);
nand U39772 (N_39772,N_39181,N_39458);
and U39773 (N_39773,N_39490,N_39450);
or U39774 (N_39774,N_39010,N_39353);
nand U39775 (N_39775,N_39436,N_39489);
nor U39776 (N_39776,N_39267,N_39367);
nor U39777 (N_39777,N_39476,N_39150);
xnor U39778 (N_39778,N_39415,N_39257);
or U39779 (N_39779,N_39422,N_39451);
nor U39780 (N_39780,N_39459,N_39399);
and U39781 (N_39781,N_39125,N_39141);
nand U39782 (N_39782,N_39372,N_39470);
and U39783 (N_39783,N_39121,N_39288);
or U39784 (N_39784,N_39420,N_39204);
nor U39785 (N_39785,N_39093,N_39314);
xnor U39786 (N_39786,N_39336,N_39474);
and U39787 (N_39787,N_39144,N_39219);
or U39788 (N_39788,N_39288,N_39086);
or U39789 (N_39789,N_39438,N_39307);
or U39790 (N_39790,N_39400,N_39039);
and U39791 (N_39791,N_39305,N_39477);
nand U39792 (N_39792,N_39288,N_39245);
nor U39793 (N_39793,N_39068,N_39091);
and U39794 (N_39794,N_39166,N_39384);
xnor U39795 (N_39795,N_39294,N_39315);
nor U39796 (N_39796,N_39074,N_39211);
or U39797 (N_39797,N_39450,N_39391);
or U39798 (N_39798,N_39035,N_39082);
or U39799 (N_39799,N_39411,N_39180);
nor U39800 (N_39800,N_39228,N_39097);
nand U39801 (N_39801,N_39180,N_39067);
and U39802 (N_39802,N_39274,N_39343);
xor U39803 (N_39803,N_39202,N_39024);
or U39804 (N_39804,N_39215,N_39137);
or U39805 (N_39805,N_39161,N_39483);
and U39806 (N_39806,N_39346,N_39309);
xnor U39807 (N_39807,N_39273,N_39333);
nor U39808 (N_39808,N_39322,N_39077);
xor U39809 (N_39809,N_39075,N_39446);
nor U39810 (N_39810,N_39313,N_39061);
xnor U39811 (N_39811,N_39026,N_39408);
xnor U39812 (N_39812,N_39283,N_39325);
xnor U39813 (N_39813,N_39401,N_39039);
or U39814 (N_39814,N_39311,N_39103);
or U39815 (N_39815,N_39435,N_39464);
nor U39816 (N_39816,N_39249,N_39436);
xnor U39817 (N_39817,N_39170,N_39315);
nand U39818 (N_39818,N_39487,N_39440);
nand U39819 (N_39819,N_39185,N_39108);
xnor U39820 (N_39820,N_39301,N_39087);
or U39821 (N_39821,N_39034,N_39194);
xnor U39822 (N_39822,N_39208,N_39252);
and U39823 (N_39823,N_39281,N_39007);
and U39824 (N_39824,N_39351,N_39213);
xnor U39825 (N_39825,N_39067,N_39281);
nand U39826 (N_39826,N_39345,N_39112);
nand U39827 (N_39827,N_39370,N_39196);
or U39828 (N_39828,N_39030,N_39000);
nor U39829 (N_39829,N_39435,N_39305);
nand U39830 (N_39830,N_39177,N_39348);
or U39831 (N_39831,N_39250,N_39354);
nor U39832 (N_39832,N_39298,N_39181);
xnor U39833 (N_39833,N_39166,N_39138);
nand U39834 (N_39834,N_39360,N_39310);
nand U39835 (N_39835,N_39290,N_39386);
nor U39836 (N_39836,N_39310,N_39492);
and U39837 (N_39837,N_39378,N_39397);
and U39838 (N_39838,N_39402,N_39485);
nand U39839 (N_39839,N_39102,N_39071);
or U39840 (N_39840,N_39085,N_39361);
xor U39841 (N_39841,N_39084,N_39351);
xnor U39842 (N_39842,N_39469,N_39373);
and U39843 (N_39843,N_39148,N_39081);
xnor U39844 (N_39844,N_39435,N_39353);
nand U39845 (N_39845,N_39102,N_39251);
or U39846 (N_39846,N_39296,N_39411);
nor U39847 (N_39847,N_39330,N_39352);
xnor U39848 (N_39848,N_39456,N_39263);
xnor U39849 (N_39849,N_39485,N_39036);
nor U39850 (N_39850,N_39044,N_39002);
nor U39851 (N_39851,N_39439,N_39496);
or U39852 (N_39852,N_39481,N_39310);
nor U39853 (N_39853,N_39037,N_39024);
nor U39854 (N_39854,N_39440,N_39485);
nor U39855 (N_39855,N_39174,N_39249);
nand U39856 (N_39856,N_39342,N_39280);
nand U39857 (N_39857,N_39205,N_39060);
or U39858 (N_39858,N_39207,N_39233);
xnor U39859 (N_39859,N_39444,N_39360);
and U39860 (N_39860,N_39201,N_39207);
nor U39861 (N_39861,N_39308,N_39179);
nand U39862 (N_39862,N_39294,N_39362);
and U39863 (N_39863,N_39083,N_39133);
nor U39864 (N_39864,N_39399,N_39298);
nand U39865 (N_39865,N_39137,N_39418);
nand U39866 (N_39866,N_39050,N_39306);
and U39867 (N_39867,N_39338,N_39170);
xnor U39868 (N_39868,N_39011,N_39203);
nand U39869 (N_39869,N_39326,N_39086);
nor U39870 (N_39870,N_39112,N_39070);
xnor U39871 (N_39871,N_39058,N_39221);
nor U39872 (N_39872,N_39074,N_39394);
or U39873 (N_39873,N_39318,N_39271);
and U39874 (N_39874,N_39401,N_39481);
or U39875 (N_39875,N_39499,N_39270);
and U39876 (N_39876,N_39432,N_39053);
nor U39877 (N_39877,N_39211,N_39392);
nand U39878 (N_39878,N_39372,N_39156);
nor U39879 (N_39879,N_39480,N_39417);
xor U39880 (N_39880,N_39167,N_39198);
xnor U39881 (N_39881,N_39120,N_39351);
nor U39882 (N_39882,N_39399,N_39385);
or U39883 (N_39883,N_39224,N_39316);
nor U39884 (N_39884,N_39429,N_39012);
and U39885 (N_39885,N_39353,N_39364);
xnor U39886 (N_39886,N_39001,N_39248);
or U39887 (N_39887,N_39151,N_39340);
nand U39888 (N_39888,N_39060,N_39497);
and U39889 (N_39889,N_39302,N_39070);
or U39890 (N_39890,N_39129,N_39088);
or U39891 (N_39891,N_39123,N_39174);
nor U39892 (N_39892,N_39248,N_39198);
xor U39893 (N_39893,N_39355,N_39275);
xnor U39894 (N_39894,N_39377,N_39287);
xor U39895 (N_39895,N_39467,N_39108);
and U39896 (N_39896,N_39409,N_39406);
nand U39897 (N_39897,N_39302,N_39079);
and U39898 (N_39898,N_39095,N_39113);
and U39899 (N_39899,N_39230,N_39244);
or U39900 (N_39900,N_39383,N_39398);
xnor U39901 (N_39901,N_39288,N_39116);
or U39902 (N_39902,N_39203,N_39041);
xnor U39903 (N_39903,N_39380,N_39333);
and U39904 (N_39904,N_39290,N_39101);
and U39905 (N_39905,N_39354,N_39353);
nor U39906 (N_39906,N_39489,N_39391);
nand U39907 (N_39907,N_39486,N_39362);
xor U39908 (N_39908,N_39073,N_39168);
nand U39909 (N_39909,N_39259,N_39118);
or U39910 (N_39910,N_39121,N_39184);
nand U39911 (N_39911,N_39043,N_39242);
nor U39912 (N_39912,N_39048,N_39154);
nor U39913 (N_39913,N_39151,N_39044);
and U39914 (N_39914,N_39059,N_39003);
xnor U39915 (N_39915,N_39091,N_39080);
xor U39916 (N_39916,N_39334,N_39054);
or U39917 (N_39917,N_39059,N_39122);
nor U39918 (N_39918,N_39156,N_39460);
nand U39919 (N_39919,N_39441,N_39229);
xor U39920 (N_39920,N_39052,N_39055);
and U39921 (N_39921,N_39439,N_39295);
nor U39922 (N_39922,N_39283,N_39151);
xor U39923 (N_39923,N_39484,N_39178);
or U39924 (N_39924,N_39041,N_39321);
nor U39925 (N_39925,N_39223,N_39054);
xor U39926 (N_39926,N_39472,N_39067);
nor U39927 (N_39927,N_39026,N_39440);
or U39928 (N_39928,N_39297,N_39029);
nand U39929 (N_39929,N_39212,N_39495);
and U39930 (N_39930,N_39007,N_39311);
and U39931 (N_39931,N_39129,N_39119);
xnor U39932 (N_39932,N_39306,N_39342);
or U39933 (N_39933,N_39108,N_39437);
xor U39934 (N_39934,N_39325,N_39299);
or U39935 (N_39935,N_39233,N_39287);
nor U39936 (N_39936,N_39061,N_39324);
or U39937 (N_39937,N_39281,N_39136);
nand U39938 (N_39938,N_39252,N_39398);
and U39939 (N_39939,N_39217,N_39007);
nand U39940 (N_39940,N_39300,N_39145);
xor U39941 (N_39941,N_39390,N_39086);
or U39942 (N_39942,N_39008,N_39188);
nand U39943 (N_39943,N_39113,N_39240);
xnor U39944 (N_39944,N_39284,N_39386);
nand U39945 (N_39945,N_39135,N_39352);
nand U39946 (N_39946,N_39066,N_39482);
nand U39947 (N_39947,N_39374,N_39496);
nand U39948 (N_39948,N_39260,N_39279);
nor U39949 (N_39949,N_39029,N_39232);
and U39950 (N_39950,N_39015,N_39474);
nor U39951 (N_39951,N_39158,N_39171);
or U39952 (N_39952,N_39445,N_39032);
and U39953 (N_39953,N_39064,N_39436);
nor U39954 (N_39954,N_39252,N_39454);
or U39955 (N_39955,N_39249,N_39467);
and U39956 (N_39956,N_39462,N_39472);
nand U39957 (N_39957,N_39280,N_39185);
nor U39958 (N_39958,N_39365,N_39401);
nand U39959 (N_39959,N_39024,N_39237);
nand U39960 (N_39960,N_39171,N_39358);
nor U39961 (N_39961,N_39303,N_39397);
xnor U39962 (N_39962,N_39364,N_39233);
xnor U39963 (N_39963,N_39468,N_39435);
nor U39964 (N_39964,N_39265,N_39100);
xnor U39965 (N_39965,N_39012,N_39252);
nand U39966 (N_39966,N_39433,N_39374);
xor U39967 (N_39967,N_39077,N_39369);
nor U39968 (N_39968,N_39323,N_39334);
and U39969 (N_39969,N_39189,N_39245);
or U39970 (N_39970,N_39373,N_39035);
xor U39971 (N_39971,N_39309,N_39289);
and U39972 (N_39972,N_39394,N_39109);
or U39973 (N_39973,N_39400,N_39215);
or U39974 (N_39974,N_39166,N_39055);
xor U39975 (N_39975,N_39174,N_39225);
xor U39976 (N_39976,N_39454,N_39310);
nand U39977 (N_39977,N_39459,N_39486);
nand U39978 (N_39978,N_39282,N_39126);
xnor U39979 (N_39979,N_39469,N_39499);
xnor U39980 (N_39980,N_39317,N_39382);
nor U39981 (N_39981,N_39213,N_39053);
or U39982 (N_39982,N_39246,N_39338);
or U39983 (N_39983,N_39494,N_39158);
nand U39984 (N_39984,N_39227,N_39341);
nor U39985 (N_39985,N_39140,N_39262);
nor U39986 (N_39986,N_39315,N_39228);
nor U39987 (N_39987,N_39014,N_39034);
nor U39988 (N_39988,N_39372,N_39290);
or U39989 (N_39989,N_39136,N_39300);
or U39990 (N_39990,N_39450,N_39121);
nand U39991 (N_39991,N_39287,N_39013);
nand U39992 (N_39992,N_39006,N_39177);
xnor U39993 (N_39993,N_39306,N_39104);
or U39994 (N_39994,N_39498,N_39317);
nand U39995 (N_39995,N_39294,N_39372);
nor U39996 (N_39996,N_39007,N_39312);
nand U39997 (N_39997,N_39325,N_39270);
or U39998 (N_39998,N_39339,N_39053);
or U39999 (N_39999,N_39412,N_39144);
nand U40000 (N_40000,N_39899,N_39716);
nand U40001 (N_40001,N_39526,N_39965);
nand U40002 (N_40002,N_39536,N_39921);
or U40003 (N_40003,N_39616,N_39868);
xor U40004 (N_40004,N_39556,N_39508);
nand U40005 (N_40005,N_39957,N_39988);
nand U40006 (N_40006,N_39719,N_39749);
or U40007 (N_40007,N_39960,N_39664);
nand U40008 (N_40008,N_39581,N_39561);
or U40009 (N_40009,N_39961,N_39819);
or U40010 (N_40010,N_39609,N_39946);
or U40011 (N_40011,N_39678,N_39850);
xnor U40012 (N_40012,N_39816,N_39714);
nand U40013 (N_40013,N_39847,N_39689);
and U40014 (N_40014,N_39766,N_39785);
nor U40015 (N_40015,N_39618,N_39895);
or U40016 (N_40016,N_39948,N_39559);
nor U40017 (N_40017,N_39791,N_39949);
xor U40018 (N_40018,N_39625,N_39748);
and U40019 (N_40019,N_39881,N_39637);
xnor U40020 (N_40020,N_39548,N_39509);
or U40021 (N_40021,N_39677,N_39597);
nand U40022 (N_40022,N_39913,N_39639);
xor U40023 (N_40023,N_39926,N_39553);
nand U40024 (N_40024,N_39586,N_39519);
xnor U40025 (N_40025,N_39826,N_39722);
nor U40026 (N_40026,N_39825,N_39588);
nand U40027 (N_40027,N_39869,N_39872);
nand U40028 (N_40028,N_39940,N_39514);
nand U40029 (N_40029,N_39699,N_39930);
or U40030 (N_40030,N_39773,N_39587);
or U40031 (N_40031,N_39684,N_39758);
or U40032 (N_40032,N_39855,N_39551);
nand U40033 (N_40033,N_39840,N_39734);
and U40034 (N_40034,N_39835,N_39781);
nand U40035 (N_40035,N_39518,N_39631);
xor U40036 (N_40036,N_39828,N_39800);
nand U40037 (N_40037,N_39848,N_39761);
nor U40038 (N_40038,N_39894,N_39697);
xnor U40039 (N_40039,N_39995,N_39602);
xnor U40040 (N_40040,N_39670,N_39683);
xnor U40041 (N_40041,N_39686,N_39552);
nor U40042 (N_40042,N_39731,N_39896);
nand U40043 (N_40043,N_39992,N_39768);
or U40044 (N_40044,N_39964,N_39577);
or U40045 (N_40045,N_39517,N_39541);
and U40046 (N_40046,N_39971,N_39891);
and U40047 (N_40047,N_39568,N_39929);
and U40048 (N_40048,N_39582,N_39524);
xor U40049 (N_40049,N_39626,N_39762);
nor U40050 (N_40050,N_39744,N_39500);
or U40051 (N_40051,N_39924,N_39994);
and U40052 (N_40052,N_39707,N_39943);
nor U40053 (N_40053,N_39874,N_39736);
xor U40054 (N_40054,N_39877,N_39737);
xor U40055 (N_40055,N_39706,N_39538);
nand U40056 (N_40056,N_39607,N_39531);
nand U40057 (N_40057,N_39764,N_39563);
nor U40058 (N_40058,N_39991,N_39735);
and U40059 (N_40059,N_39729,N_39910);
and U40060 (N_40060,N_39693,N_39922);
and U40061 (N_40061,N_39525,N_39657);
or U40062 (N_40062,N_39507,N_39520);
or U40063 (N_40063,N_39919,N_39644);
nor U40064 (N_40064,N_39743,N_39837);
nor U40065 (N_40065,N_39622,N_39888);
nor U40066 (N_40066,N_39557,N_39634);
xnor U40067 (N_40067,N_39599,N_39604);
nor U40068 (N_40068,N_39688,N_39522);
xnor U40069 (N_40069,N_39720,N_39628);
nor U40070 (N_40070,N_39777,N_39590);
and U40071 (N_40071,N_39844,N_39876);
nor U40072 (N_40072,N_39680,N_39763);
nand U40073 (N_40073,N_39663,N_39516);
xor U40074 (N_40074,N_39882,N_39562);
or U40075 (N_40075,N_39851,N_39667);
xnor U40076 (N_40076,N_39576,N_39886);
xor U40077 (N_40077,N_39713,N_39540);
and U40078 (N_40078,N_39905,N_39727);
and U40079 (N_40079,N_39972,N_39760);
and U40080 (N_40080,N_39928,N_39963);
or U40081 (N_40081,N_39787,N_39594);
xnor U40082 (N_40082,N_39936,N_39528);
nor U40083 (N_40083,N_39813,N_39756);
nand U40084 (N_40084,N_39726,N_39580);
xnor U40085 (N_40085,N_39887,N_39932);
nand U40086 (N_40086,N_39914,N_39671);
or U40087 (N_40087,N_39504,N_39752);
nor U40088 (N_40088,N_39765,N_39695);
nor U40089 (N_40089,N_39739,N_39814);
nand U40090 (N_40090,N_39705,N_39614);
nor U40091 (N_40091,N_39902,N_39821);
nand U40092 (N_40092,N_39794,N_39619);
nor U40093 (N_40093,N_39983,N_39757);
and U40094 (N_40094,N_39672,N_39854);
nor U40095 (N_40095,N_39550,N_39792);
nand U40096 (N_40096,N_39673,N_39645);
xor U40097 (N_40097,N_39786,N_39998);
xor U40098 (N_40098,N_39530,N_39805);
or U40099 (N_40099,N_39651,N_39674);
xor U40100 (N_40100,N_39574,N_39901);
nor U40101 (N_40101,N_39897,N_39935);
nor U40102 (N_40102,N_39579,N_39687);
and U40103 (N_40103,N_39993,N_39560);
or U40104 (N_40104,N_39630,N_39959);
xor U40105 (N_40105,N_39798,N_39648);
and U40106 (N_40106,N_39621,N_39989);
nor U40107 (N_40107,N_39823,N_39656);
and U40108 (N_40108,N_39985,N_39937);
nor U40109 (N_40109,N_39849,N_39542);
xnor U40110 (N_40110,N_39703,N_39808);
or U40111 (N_40111,N_39506,N_39543);
nor U40112 (N_40112,N_39832,N_39523);
nor U40113 (N_40113,N_39638,N_39810);
xnor U40114 (N_40114,N_39567,N_39533);
or U40115 (N_40115,N_39903,N_39747);
or U40116 (N_40116,N_39841,N_39941);
nand U40117 (N_40117,N_39564,N_39584);
xor U40118 (N_40118,N_39733,N_39605);
nor U40119 (N_40119,N_39806,N_39973);
nor U40120 (N_40120,N_39596,N_39569);
nand U40121 (N_40121,N_39640,N_39724);
nor U40122 (N_40122,N_39575,N_39978);
xor U40123 (N_40123,N_39950,N_39570);
xor U40124 (N_40124,N_39898,N_39804);
xnor U40125 (N_40125,N_39939,N_39968);
or U40126 (N_40126,N_39999,N_39878);
or U40127 (N_40127,N_39947,N_39955);
or U40128 (N_40128,N_39967,N_39982);
nor U40129 (N_40129,N_39970,N_39865);
xor U40130 (N_40130,N_39740,N_39641);
and U40131 (N_40131,N_39723,N_39836);
xor U40132 (N_40132,N_39775,N_39824);
nor U40133 (N_40133,N_39751,N_39502);
nand U40134 (N_40134,N_39938,N_39698);
nor U40135 (N_40135,N_39613,N_39709);
nand U40136 (N_40136,N_39984,N_39746);
nor U40137 (N_40137,N_39815,N_39701);
or U40138 (N_40138,N_39554,N_39573);
and U40139 (N_40139,N_39863,N_39803);
xnor U40140 (N_40140,N_39704,N_39527);
and U40141 (N_40141,N_39708,N_39510);
and U40142 (N_40142,N_39535,N_39655);
and U40143 (N_40143,N_39976,N_39750);
nand U40144 (N_40144,N_39931,N_39916);
xnor U40145 (N_40145,N_39732,N_39912);
nor U40146 (N_40146,N_39608,N_39691);
and U40147 (N_40147,N_39846,N_39990);
xor U40148 (N_40148,N_39742,N_39893);
nor U40149 (N_40149,N_39512,N_39890);
and U40150 (N_40150,N_39532,N_39521);
nand U40151 (N_40151,N_39856,N_39546);
or U40152 (N_40152,N_39710,N_39636);
and U40153 (N_40153,N_39754,N_39859);
nor U40154 (N_40154,N_39980,N_39996);
nor U40155 (N_40155,N_39873,N_39771);
nor U40156 (N_40156,N_39629,N_39730);
nand U40157 (N_40157,N_39981,N_39759);
and U40158 (N_40158,N_39889,N_39774);
xor U40159 (N_40159,N_39880,N_39820);
and U40160 (N_40160,N_39601,N_39962);
or U40161 (N_40161,N_39852,N_39652);
and U40162 (N_40162,N_39627,N_39923);
xor U40163 (N_40163,N_39862,N_39665);
and U40164 (N_40164,N_39864,N_39918);
nand U40165 (N_40165,N_39915,N_39911);
or U40166 (N_40166,N_39501,N_39958);
or U40167 (N_40167,N_39845,N_39544);
xnor U40168 (N_40168,N_39945,N_39583);
or U40169 (N_40169,N_39843,N_39585);
nand U40170 (N_40170,N_39809,N_39801);
and U40171 (N_40171,N_39690,N_39666);
or U40172 (N_40172,N_39593,N_39831);
nand U40173 (N_40173,N_39977,N_39812);
xor U40174 (N_40174,N_39830,N_39660);
xor U40175 (N_40175,N_39776,N_39646);
nand U40176 (N_40176,N_39696,N_39642);
or U40177 (N_40177,N_39956,N_39503);
nand U40178 (N_40178,N_39592,N_39974);
and U40179 (N_40179,N_39649,N_39871);
and U40180 (N_40180,N_39661,N_39537);
and U40181 (N_40181,N_39987,N_39595);
or U40182 (N_40182,N_39909,N_39860);
xnor U40183 (N_40183,N_39857,N_39838);
or U40184 (N_40184,N_39591,N_39834);
xor U40185 (N_40185,N_39904,N_39600);
nand U40186 (N_40186,N_39545,N_39799);
xor U40187 (N_40187,N_39505,N_39782);
and U40188 (N_40188,N_39951,N_39753);
nor U40189 (N_40189,N_39632,N_39668);
xnor U40190 (N_40190,N_39702,N_39685);
nand U40191 (N_40191,N_39817,N_39927);
xnor U40192 (N_40192,N_39783,N_39717);
and U40193 (N_40193,N_39784,N_39885);
or U40194 (N_40194,N_39529,N_39884);
or U40195 (N_40195,N_39953,N_39615);
xnor U40196 (N_40196,N_39802,N_39853);
and U40197 (N_40197,N_39547,N_39997);
xnor U40198 (N_40198,N_39767,N_39606);
xor U40199 (N_40199,N_39611,N_39807);
and U40200 (N_40200,N_39669,N_39907);
or U40201 (N_40201,N_39659,N_39900);
nor U40202 (N_40202,N_39979,N_39738);
or U40203 (N_40203,N_39650,N_39858);
or U40204 (N_40204,N_39692,N_39610);
nor U40205 (N_40205,N_39612,N_39966);
nand U40206 (N_40206,N_39513,N_39617);
xor U40207 (N_40207,N_39906,N_39558);
nand U40208 (N_40208,N_39623,N_39725);
and U40209 (N_40209,N_39788,N_39839);
and U40210 (N_40210,N_39694,N_39633);
nor U40211 (N_40211,N_39549,N_39986);
or U40212 (N_40212,N_39675,N_39866);
nand U40213 (N_40213,N_39578,N_39620);
nand U40214 (N_40214,N_39572,N_39511);
xor U40215 (N_40215,N_39954,N_39711);
or U40216 (N_40216,N_39875,N_39712);
nor U40217 (N_40217,N_39565,N_39755);
nor U40218 (N_40218,N_39975,N_39571);
or U40219 (N_40219,N_39793,N_39917);
nand U40220 (N_40220,N_39870,N_39778);
and U40221 (N_40221,N_39933,N_39741);
xor U40222 (N_40222,N_39908,N_39879);
xnor U40223 (N_40223,N_39676,N_39654);
nand U40224 (N_40224,N_39624,N_39681);
or U40225 (N_40225,N_39944,N_39925);
nor U40226 (N_40226,N_39643,N_39934);
and U40227 (N_40227,N_39833,N_39769);
and U40228 (N_40228,N_39790,N_39653);
xor U40229 (N_40229,N_39779,N_39797);
nor U40230 (N_40230,N_39796,N_39682);
nand U40231 (N_40231,N_39883,N_39811);
nand U40232 (N_40232,N_39969,N_39728);
xor U40233 (N_40233,N_39721,N_39555);
and U40234 (N_40234,N_39679,N_39598);
xnor U40235 (N_40235,N_39867,N_39795);
and U40236 (N_40236,N_39647,N_39861);
nand U40237 (N_40237,N_39818,N_39515);
or U40238 (N_40238,N_39700,N_39603);
xor U40239 (N_40239,N_39772,N_39780);
and U40240 (N_40240,N_39745,N_39715);
nor U40241 (N_40241,N_39789,N_39942);
xnor U40242 (N_40242,N_39662,N_39635);
nor U40243 (N_40243,N_39892,N_39952);
nor U40244 (N_40244,N_39829,N_39822);
xor U40245 (N_40245,N_39827,N_39566);
nand U40246 (N_40246,N_39718,N_39658);
nor U40247 (N_40247,N_39534,N_39589);
and U40248 (N_40248,N_39842,N_39539);
nor U40249 (N_40249,N_39920,N_39770);
nor U40250 (N_40250,N_39579,N_39945);
xnor U40251 (N_40251,N_39513,N_39658);
or U40252 (N_40252,N_39994,N_39917);
or U40253 (N_40253,N_39911,N_39684);
or U40254 (N_40254,N_39959,N_39537);
nand U40255 (N_40255,N_39598,N_39526);
nand U40256 (N_40256,N_39912,N_39859);
or U40257 (N_40257,N_39612,N_39598);
nand U40258 (N_40258,N_39849,N_39665);
nor U40259 (N_40259,N_39946,N_39854);
or U40260 (N_40260,N_39651,N_39689);
and U40261 (N_40261,N_39726,N_39755);
nand U40262 (N_40262,N_39762,N_39573);
xnor U40263 (N_40263,N_39663,N_39565);
and U40264 (N_40264,N_39697,N_39787);
or U40265 (N_40265,N_39843,N_39874);
and U40266 (N_40266,N_39889,N_39758);
and U40267 (N_40267,N_39693,N_39602);
xnor U40268 (N_40268,N_39507,N_39826);
or U40269 (N_40269,N_39726,N_39538);
xnor U40270 (N_40270,N_39554,N_39540);
or U40271 (N_40271,N_39853,N_39630);
xor U40272 (N_40272,N_39823,N_39508);
and U40273 (N_40273,N_39507,N_39714);
nand U40274 (N_40274,N_39741,N_39573);
nand U40275 (N_40275,N_39923,N_39571);
xor U40276 (N_40276,N_39834,N_39997);
nand U40277 (N_40277,N_39816,N_39845);
or U40278 (N_40278,N_39848,N_39591);
or U40279 (N_40279,N_39874,N_39705);
nor U40280 (N_40280,N_39801,N_39883);
nand U40281 (N_40281,N_39513,N_39533);
or U40282 (N_40282,N_39604,N_39649);
and U40283 (N_40283,N_39853,N_39859);
nor U40284 (N_40284,N_39557,N_39931);
or U40285 (N_40285,N_39715,N_39992);
nand U40286 (N_40286,N_39776,N_39541);
xor U40287 (N_40287,N_39609,N_39809);
xor U40288 (N_40288,N_39669,N_39528);
and U40289 (N_40289,N_39986,N_39802);
and U40290 (N_40290,N_39698,N_39621);
and U40291 (N_40291,N_39704,N_39779);
nand U40292 (N_40292,N_39579,N_39582);
xnor U40293 (N_40293,N_39514,N_39836);
nor U40294 (N_40294,N_39886,N_39637);
nand U40295 (N_40295,N_39942,N_39979);
nand U40296 (N_40296,N_39869,N_39645);
nor U40297 (N_40297,N_39922,N_39890);
nand U40298 (N_40298,N_39922,N_39799);
nand U40299 (N_40299,N_39742,N_39852);
or U40300 (N_40300,N_39623,N_39795);
nor U40301 (N_40301,N_39547,N_39912);
and U40302 (N_40302,N_39682,N_39527);
or U40303 (N_40303,N_39993,N_39812);
xnor U40304 (N_40304,N_39686,N_39981);
and U40305 (N_40305,N_39940,N_39595);
xor U40306 (N_40306,N_39832,N_39794);
nor U40307 (N_40307,N_39644,N_39528);
nor U40308 (N_40308,N_39634,N_39987);
nor U40309 (N_40309,N_39972,N_39532);
and U40310 (N_40310,N_39810,N_39997);
or U40311 (N_40311,N_39590,N_39537);
nor U40312 (N_40312,N_39826,N_39624);
nand U40313 (N_40313,N_39694,N_39887);
or U40314 (N_40314,N_39537,N_39513);
xor U40315 (N_40315,N_39660,N_39737);
xnor U40316 (N_40316,N_39564,N_39946);
and U40317 (N_40317,N_39958,N_39631);
and U40318 (N_40318,N_39752,N_39753);
and U40319 (N_40319,N_39586,N_39576);
xor U40320 (N_40320,N_39674,N_39731);
nor U40321 (N_40321,N_39787,N_39786);
xnor U40322 (N_40322,N_39812,N_39704);
nand U40323 (N_40323,N_39503,N_39677);
or U40324 (N_40324,N_39958,N_39632);
and U40325 (N_40325,N_39844,N_39864);
and U40326 (N_40326,N_39768,N_39552);
xor U40327 (N_40327,N_39876,N_39764);
nor U40328 (N_40328,N_39847,N_39650);
or U40329 (N_40329,N_39604,N_39841);
nor U40330 (N_40330,N_39897,N_39705);
and U40331 (N_40331,N_39984,N_39848);
or U40332 (N_40332,N_39638,N_39924);
nor U40333 (N_40333,N_39506,N_39797);
or U40334 (N_40334,N_39710,N_39976);
nor U40335 (N_40335,N_39829,N_39805);
nor U40336 (N_40336,N_39825,N_39670);
nand U40337 (N_40337,N_39781,N_39606);
nor U40338 (N_40338,N_39619,N_39940);
xor U40339 (N_40339,N_39933,N_39879);
and U40340 (N_40340,N_39933,N_39526);
xnor U40341 (N_40341,N_39665,N_39712);
nand U40342 (N_40342,N_39805,N_39674);
nor U40343 (N_40343,N_39742,N_39914);
nand U40344 (N_40344,N_39599,N_39719);
or U40345 (N_40345,N_39810,N_39512);
and U40346 (N_40346,N_39714,N_39842);
nor U40347 (N_40347,N_39789,N_39947);
nand U40348 (N_40348,N_39609,N_39937);
nand U40349 (N_40349,N_39632,N_39782);
nor U40350 (N_40350,N_39761,N_39945);
or U40351 (N_40351,N_39829,N_39738);
or U40352 (N_40352,N_39919,N_39799);
or U40353 (N_40353,N_39954,N_39533);
nand U40354 (N_40354,N_39893,N_39556);
or U40355 (N_40355,N_39875,N_39684);
nor U40356 (N_40356,N_39956,N_39963);
nor U40357 (N_40357,N_39592,N_39867);
nand U40358 (N_40358,N_39504,N_39634);
nand U40359 (N_40359,N_39539,N_39578);
nand U40360 (N_40360,N_39820,N_39861);
or U40361 (N_40361,N_39823,N_39728);
nand U40362 (N_40362,N_39855,N_39543);
xor U40363 (N_40363,N_39709,N_39937);
nand U40364 (N_40364,N_39618,N_39913);
or U40365 (N_40365,N_39723,N_39631);
xnor U40366 (N_40366,N_39592,N_39791);
xnor U40367 (N_40367,N_39926,N_39923);
xor U40368 (N_40368,N_39746,N_39819);
and U40369 (N_40369,N_39542,N_39645);
nor U40370 (N_40370,N_39695,N_39587);
or U40371 (N_40371,N_39954,N_39740);
and U40372 (N_40372,N_39717,N_39590);
nor U40373 (N_40373,N_39695,N_39747);
or U40374 (N_40374,N_39528,N_39944);
and U40375 (N_40375,N_39797,N_39545);
nor U40376 (N_40376,N_39853,N_39664);
or U40377 (N_40377,N_39827,N_39765);
or U40378 (N_40378,N_39996,N_39864);
or U40379 (N_40379,N_39510,N_39862);
or U40380 (N_40380,N_39714,N_39707);
and U40381 (N_40381,N_39753,N_39982);
and U40382 (N_40382,N_39707,N_39586);
nand U40383 (N_40383,N_39876,N_39596);
or U40384 (N_40384,N_39646,N_39536);
and U40385 (N_40385,N_39953,N_39613);
nand U40386 (N_40386,N_39582,N_39986);
and U40387 (N_40387,N_39548,N_39713);
and U40388 (N_40388,N_39549,N_39932);
and U40389 (N_40389,N_39523,N_39818);
nor U40390 (N_40390,N_39533,N_39782);
nand U40391 (N_40391,N_39716,N_39715);
nand U40392 (N_40392,N_39755,N_39974);
nor U40393 (N_40393,N_39733,N_39881);
or U40394 (N_40394,N_39913,N_39548);
or U40395 (N_40395,N_39836,N_39721);
nand U40396 (N_40396,N_39954,N_39952);
xor U40397 (N_40397,N_39505,N_39718);
xor U40398 (N_40398,N_39561,N_39766);
nand U40399 (N_40399,N_39591,N_39762);
nand U40400 (N_40400,N_39845,N_39947);
xor U40401 (N_40401,N_39858,N_39986);
and U40402 (N_40402,N_39639,N_39769);
nand U40403 (N_40403,N_39712,N_39623);
xor U40404 (N_40404,N_39814,N_39713);
nand U40405 (N_40405,N_39961,N_39798);
or U40406 (N_40406,N_39689,N_39569);
xor U40407 (N_40407,N_39604,N_39808);
nor U40408 (N_40408,N_39931,N_39583);
and U40409 (N_40409,N_39622,N_39808);
or U40410 (N_40410,N_39501,N_39570);
and U40411 (N_40411,N_39811,N_39553);
or U40412 (N_40412,N_39918,N_39838);
and U40413 (N_40413,N_39811,N_39818);
nand U40414 (N_40414,N_39718,N_39829);
and U40415 (N_40415,N_39734,N_39790);
or U40416 (N_40416,N_39518,N_39625);
nor U40417 (N_40417,N_39912,N_39806);
and U40418 (N_40418,N_39726,N_39614);
nand U40419 (N_40419,N_39961,N_39831);
and U40420 (N_40420,N_39890,N_39541);
xnor U40421 (N_40421,N_39947,N_39666);
or U40422 (N_40422,N_39829,N_39672);
or U40423 (N_40423,N_39732,N_39987);
or U40424 (N_40424,N_39563,N_39594);
or U40425 (N_40425,N_39608,N_39699);
nor U40426 (N_40426,N_39722,N_39674);
xnor U40427 (N_40427,N_39678,N_39916);
and U40428 (N_40428,N_39615,N_39507);
nor U40429 (N_40429,N_39883,N_39755);
and U40430 (N_40430,N_39605,N_39962);
nor U40431 (N_40431,N_39750,N_39978);
xor U40432 (N_40432,N_39858,N_39881);
xor U40433 (N_40433,N_39501,N_39545);
and U40434 (N_40434,N_39887,N_39689);
nand U40435 (N_40435,N_39723,N_39588);
nand U40436 (N_40436,N_39527,N_39877);
nand U40437 (N_40437,N_39549,N_39758);
nand U40438 (N_40438,N_39502,N_39971);
xor U40439 (N_40439,N_39910,N_39710);
or U40440 (N_40440,N_39821,N_39783);
nand U40441 (N_40441,N_39726,N_39842);
nor U40442 (N_40442,N_39877,N_39576);
xnor U40443 (N_40443,N_39741,N_39655);
nor U40444 (N_40444,N_39553,N_39747);
and U40445 (N_40445,N_39827,N_39558);
or U40446 (N_40446,N_39703,N_39586);
xnor U40447 (N_40447,N_39993,N_39586);
nor U40448 (N_40448,N_39903,N_39765);
xor U40449 (N_40449,N_39816,N_39643);
nor U40450 (N_40450,N_39562,N_39692);
nor U40451 (N_40451,N_39504,N_39944);
or U40452 (N_40452,N_39890,N_39838);
nor U40453 (N_40453,N_39669,N_39663);
xor U40454 (N_40454,N_39834,N_39833);
or U40455 (N_40455,N_39581,N_39752);
nor U40456 (N_40456,N_39897,N_39750);
or U40457 (N_40457,N_39687,N_39965);
nor U40458 (N_40458,N_39670,N_39631);
nor U40459 (N_40459,N_39980,N_39567);
or U40460 (N_40460,N_39654,N_39609);
nand U40461 (N_40461,N_39666,N_39855);
nand U40462 (N_40462,N_39883,N_39614);
xor U40463 (N_40463,N_39623,N_39590);
and U40464 (N_40464,N_39716,N_39543);
and U40465 (N_40465,N_39787,N_39810);
and U40466 (N_40466,N_39847,N_39893);
nor U40467 (N_40467,N_39565,N_39527);
nand U40468 (N_40468,N_39501,N_39518);
nor U40469 (N_40469,N_39552,N_39527);
xor U40470 (N_40470,N_39531,N_39588);
and U40471 (N_40471,N_39622,N_39527);
nor U40472 (N_40472,N_39839,N_39977);
nand U40473 (N_40473,N_39778,N_39502);
and U40474 (N_40474,N_39584,N_39599);
nand U40475 (N_40475,N_39527,N_39647);
nor U40476 (N_40476,N_39986,N_39646);
xor U40477 (N_40477,N_39940,N_39548);
and U40478 (N_40478,N_39788,N_39581);
xnor U40479 (N_40479,N_39513,N_39918);
nand U40480 (N_40480,N_39624,N_39667);
or U40481 (N_40481,N_39600,N_39724);
xnor U40482 (N_40482,N_39500,N_39548);
nand U40483 (N_40483,N_39602,N_39541);
nand U40484 (N_40484,N_39506,N_39672);
nand U40485 (N_40485,N_39576,N_39787);
nor U40486 (N_40486,N_39999,N_39719);
and U40487 (N_40487,N_39647,N_39999);
xor U40488 (N_40488,N_39710,N_39600);
nor U40489 (N_40489,N_39637,N_39669);
nand U40490 (N_40490,N_39565,N_39939);
and U40491 (N_40491,N_39793,N_39995);
or U40492 (N_40492,N_39800,N_39554);
or U40493 (N_40493,N_39720,N_39890);
nor U40494 (N_40494,N_39640,N_39966);
nand U40495 (N_40495,N_39802,N_39877);
and U40496 (N_40496,N_39598,N_39537);
nand U40497 (N_40497,N_39591,N_39622);
nand U40498 (N_40498,N_39870,N_39942);
nand U40499 (N_40499,N_39519,N_39520);
nor U40500 (N_40500,N_40264,N_40380);
nand U40501 (N_40501,N_40113,N_40315);
or U40502 (N_40502,N_40388,N_40486);
nand U40503 (N_40503,N_40228,N_40194);
nand U40504 (N_40504,N_40133,N_40102);
or U40505 (N_40505,N_40387,N_40129);
xor U40506 (N_40506,N_40067,N_40345);
nand U40507 (N_40507,N_40358,N_40327);
nand U40508 (N_40508,N_40151,N_40470);
xor U40509 (N_40509,N_40082,N_40379);
xor U40510 (N_40510,N_40302,N_40354);
xnor U40511 (N_40511,N_40017,N_40420);
nor U40512 (N_40512,N_40161,N_40022);
nor U40513 (N_40513,N_40477,N_40197);
nand U40514 (N_40514,N_40040,N_40253);
or U40515 (N_40515,N_40414,N_40394);
and U40516 (N_40516,N_40474,N_40135);
nand U40517 (N_40517,N_40426,N_40066);
nor U40518 (N_40518,N_40064,N_40236);
nor U40519 (N_40519,N_40068,N_40196);
xor U40520 (N_40520,N_40273,N_40294);
or U40521 (N_40521,N_40001,N_40329);
and U40522 (N_40522,N_40124,N_40347);
or U40523 (N_40523,N_40257,N_40226);
nand U40524 (N_40524,N_40446,N_40229);
nor U40525 (N_40525,N_40363,N_40009);
nor U40526 (N_40526,N_40353,N_40167);
and U40527 (N_40527,N_40313,N_40378);
or U40528 (N_40528,N_40030,N_40391);
nand U40529 (N_40529,N_40037,N_40206);
and U40530 (N_40530,N_40381,N_40403);
and U40531 (N_40531,N_40393,N_40475);
or U40532 (N_40532,N_40468,N_40193);
nor U40533 (N_40533,N_40424,N_40232);
and U40534 (N_40534,N_40285,N_40110);
nor U40535 (N_40535,N_40341,N_40283);
and U40536 (N_40536,N_40377,N_40158);
xor U40537 (N_40537,N_40091,N_40335);
nand U40538 (N_40538,N_40138,N_40152);
nor U40539 (N_40539,N_40044,N_40428);
nand U40540 (N_40540,N_40280,N_40328);
nand U40541 (N_40541,N_40089,N_40410);
nand U40542 (N_40542,N_40142,N_40185);
or U40543 (N_40543,N_40062,N_40427);
nand U40544 (N_40544,N_40339,N_40056);
xnor U40545 (N_40545,N_40049,N_40259);
nand U40546 (N_40546,N_40060,N_40351);
nor U40547 (N_40547,N_40467,N_40035);
xor U40548 (N_40548,N_40465,N_40237);
nor U40549 (N_40549,N_40348,N_40119);
and U40550 (N_40550,N_40238,N_40332);
nor U40551 (N_40551,N_40079,N_40286);
nor U40552 (N_40552,N_40109,N_40442);
and U40553 (N_40553,N_40092,N_40163);
nand U40554 (N_40554,N_40183,N_40104);
or U40555 (N_40555,N_40343,N_40225);
nor U40556 (N_40556,N_40490,N_40365);
or U40557 (N_40557,N_40148,N_40246);
or U40558 (N_40558,N_40195,N_40330);
nor U40559 (N_40559,N_40240,N_40205);
nand U40560 (N_40560,N_40250,N_40033);
xnor U40561 (N_40561,N_40170,N_40473);
nor U40562 (N_40562,N_40412,N_40457);
nand U40563 (N_40563,N_40310,N_40362);
nor U40564 (N_40564,N_40212,N_40112);
xor U40565 (N_40565,N_40449,N_40289);
and U40566 (N_40566,N_40032,N_40139);
and U40567 (N_40567,N_40231,N_40123);
nor U40568 (N_40568,N_40070,N_40439);
or U40569 (N_40569,N_40488,N_40479);
xnor U40570 (N_40570,N_40413,N_40118);
nor U40571 (N_40571,N_40371,N_40029);
and U40572 (N_40572,N_40171,N_40207);
nor U40573 (N_40573,N_40301,N_40012);
nor U40574 (N_40574,N_40369,N_40011);
xnor U40575 (N_40575,N_40499,N_40077);
nor U40576 (N_40576,N_40080,N_40149);
or U40577 (N_40577,N_40491,N_40088);
xor U40578 (N_40578,N_40191,N_40466);
nand U40579 (N_40579,N_40284,N_40462);
or U40580 (N_40580,N_40046,N_40014);
xor U40581 (N_40581,N_40188,N_40279);
nand U40582 (N_40582,N_40293,N_40125);
nand U40583 (N_40583,N_40209,N_40199);
or U40584 (N_40584,N_40055,N_40447);
or U40585 (N_40585,N_40227,N_40311);
nor U40586 (N_40586,N_40108,N_40053);
or U40587 (N_40587,N_40431,N_40287);
or U40588 (N_40588,N_40083,N_40141);
nor U40589 (N_40589,N_40072,N_40370);
nor U40590 (N_40590,N_40150,N_40024);
or U40591 (N_40591,N_40090,N_40432);
and U40592 (N_40592,N_40127,N_40058);
nor U40593 (N_40593,N_40305,N_40215);
and U40594 (N_40594,N_40153,N_40027);
nand U40595 (N_40595,N_40342,N_40034);
nand U40596 (N_40596,N_40320,N_40270);
xor U40597 (N_40597,N_40374,N_40364);
nand U40598 (N_40598,N_40013,N_40298);
and U40599 (N_40599,N_40344,N_40415);
and U40600 (N_40600,N_40075,N_40251);
nor U40601 (N_40601,N_40047,N_40222);
or U40602 (N_40602,N_40140,N_40101);
nor U40603 (N_40603,N_40445,N_40248);
nor U40604 (N_40604,N_40247,N_40172);
or U40605 (N_40605,N_40454,N_40453);
nor U40606 (N_40606,N_40189,N_40389);
xor U40607 (N_40607,N_40476,N_40418);
xor U40608 (N_40608,N_40334,N_40355);
nand U40609 (N_40609,N_40276,N_40312);
nand U40610 (N_40610,N_40041,N_40460);
nor U40611 (N_40611,N_40282,N_40448);
nand U40612 (N_40612,N_40210,N_40103);
xnor U40613 (N_40613,N_40039,N_40241);
nor U40614 (N_40614,N_40292,N_40021);
nand U40615 (N_40615,N_40242,N_40459);
nand U40616 (N_40616,N_40106,N_40233);
nor U40617 (N_40617,N_40409,N_40425);
or U40618 (N_40618,N_40497,N_40169);
or U40619 (N_40619,N_40063,N_40376);
xnor U40620 (N_40620,N_40494,N_40239);
or U40621 (N_40621,N_40417,N_40213);
and U40622 (N_40622,N_40146,N_40249);
xor U40623 (N_40623,N_40097,N_40020);
nand U40624 (N_40624,N_40093,N_40084);
nor U40625 (N_40625,N_40086,N_40190);
or U40626 (N_40626,N_40223,N_40166);
and U40627 (N_40627,N_40290,N_40438);
nor U40628 (N_40628,N_40321,N_40078);
nor U40629 (N_40629,N_40122,N_40407);
nand U40630 (N_40630,N_40252,N_40304);
and U40631 (N_40631,N_40297,N_40202);
xnor U40632 (N_40632,N_40179,N_40015);
nand U40633 (N_40633,N_40054,N_40385);
and U40634 (N_40634,N_40450,N_40340);
or U40635 (N_40635,N_40137,N_40042);
nor U40636 (N_40636,N_40319,N_40099);
nor U40637 (N_40637,N_40255,N_40131);
nor U40638 (N_40638,N_40398,N_40208);
nor U40639 (N_40639,N_40436,N_40472);
nor U40640 (N_40640,N_40366,N_40295);
nor U40641 (N_40641,N_40437,N_40395);
xor U40642 (N_40642,N_40201,N_40368);
nor U40643 (N_40643,N_40372,N_40274);
nand U40644 (N_40644,N_40105,N_40263);
and U40645 (N_40645,N_40361,N_40406);
nand U40646 (N_40646,N_40235,N_40128);
xor U40647 (N_40647,N_40126,N_40258);
or U40648 (N_40648,N_40052,N_40117);
xnor U40649 (N_40649,N_40455,N_40224);
and U40650 (N_40650,N_40057,N_40308);
nand U40651 (N_40651,N_40478,N_40303);
or U40652 (N_40652,N_40186,N_40456);
and U40653 (N_40653,N_40234,N_40217);
nand U40654 (N_40654,N_40177,N_40367);
xnor U40655 (N_40655,N_40458,N_40159);
and U40656 (N_40656,N_40045,N_40480);
and U40657 (N_40657,N_40346,N_40154);
or U40658 (N_40658,N_40300,N_40408);
xor U40659 (N_40659,N_40493,N_40435);
and U40660 (N_40660,N_40107,N_40271);
and U40661 (N_40661,N_40400,N_40096);
nor U40662 (N_40662,N_40182,N_40336);
nand U40663 (N_40663,N_40005,N_40357);
xor U40664 (N_40664,N_40007,N_40350);
nand U40665 (N_40665,N_40115,N_40178);
nand U40666 (N_40666,N_40405,N_40245);
xnor U40667 (N_40667,N_40069,N_40430);
or U40668 (N_40668,N_40114,N_40173);
nor U40669 (N_40669,N_40485,N_40204);
nand U40670 (N_40670,N_40421,N_40397);
nand U40671 (N_40671,N_40065,N_40331);
nor U40672 (N_40672,N_40230,N_40051);
and U40673 (N_40673,N_40322,N_40416);
nand U40674 (N_40674,N_40098,N_40309);
and U40675 (N_40675,N_40306,N_40451);
or U40676 (N_40676,N_40198,N_40071);
nor U40677 (N_40677,N_40471,N_40487);
nor U40678 (N_40678,N_40275,N_40121);
and U40679 (N_40679,N_40073,N_40337);
nor U40680 (N_40680,N_40254,N_40087);
or U40681 (N_40681,N_40323,N_40267);
nand U40682 (N_40682,N_40489,N_40419);
and U40683 (N_40683,N_40076,N_40243);
or U40684 (N_40684,N_40116,N_40324);
and U40685 (N_40685,N_40220,N_40100);
and U40686 (N_40686,N_40061,N_40299);
xnor U40687 (N_40687,N_40461,N_40440);
nand U40688 (N_40688,N_40010,N_40085);
xnor U40689 (N_40689,N_40018,N_40281);
nor U40690 (N_40690,N_40296,N_40145);
nand U40691 (N_40691,N_40349,N_40175);
nor U40692 (N_40692,N_40482,N_40025);
or U40693 (N_40693,N_40433,N_40260);
or U40694 (N_40694,N_40000,N_40404);
and U40695 (N_40695,N_40006,N_40272);
xor U40696 (N_40696,N_40483,N_40036);
or U40697 (N_40697,N_40307,N_40143);
nand U40698 (N_40698,N_40095,N_40402);
xnor U40699 (N_40699,N_40481,N_40288);
xor U40700 (N_40700,N_40023,N_40390);
nor U40701 (N_40701,N_40168,N_40333);
or U40702 (N_40702,N_40094,N_40463);
xor U40703 (N_40703,N_40180,N_40192);
or U40704 (N_40704,N_40050,N_40269);
and U40705 (N_40705,N_40160,N_40016);
or U40706 (N_40706,N_40261,N_40136);
xnor U40707 (N_40707,N_40003,N_40111);
xor U40708 (N_40708,N_40059,N_40434);
nand U40709 (N_40709,N_40375,N_40081);
nand U40710 (N_40710,N_40422,N_40469);
and U40711 (N_40711,N_40028,N_40443);
nand U40712 (N_40712,N_40317,N_40155);
or U40713 (N_40713,N_40256,N_40384);
or U40714 (N_40714,N_40266,N_40074);
or U40715 (N_40715,N_40268,N_40164);
and U40716 (N_40716,N_40120,N_40211);
or U40717 (N_40717,N_40382,N_40026);
xnor U40718 (N_40718,N_40399,N_40359);
or U40719 (N_40719,N_40356,N_40214);
xor U40720 (N_40720,N_40495,N_40498);
or U40721 (N_40721,N_40244,N_40444);
nand U40722 (N_40722,N_40144,N_40203);
nor U40723 (N_40723,N_40219,N_40130);
xor U40724 (N_40724,N_40165,N_40265);
or U40725 (N_40725,N_40360,N_40277);
and U40726 (N_40726,N_40134,N_40314);
or U40727 (N_40727,N_40019,N_40423);
or U40728 (N_40728,N_40156,N_40386);
xnor U40729 (N_40729,N_40200,N_40218);
nor U40730 (N_40730,N_40338,N_40325);
and U40731 (N_40731,N_40484,N_40043);
nor U40732 (N_40732,N_40132,N_40401);
xor U40733 (N_40733,N_40216,N_40429);
xnor U40734 (N_40734,N_40031,N_40174);
nor U40735 (N_40735,N_40278,N_40352);
xor U40736 (N_40736,N_40373,N_40048);
and U40737 (N_40737,N_40038,N_40008);
xor U40738 (N_40738,N_40392,N_40187);
and U40739 (N_40739,N_40318,N_40184);
or U40740 (N_40740,N_40411,N_40383);
nor U40741 (N_40741,N_40004,N_40492);
and U40742 (N_40742,N_40162,N_40181);
nand U40743 (N_40743,N_40221,N_40326);
and U40744 (N_40744,N_40002,N_40316);
or U40745 (N_40745,N_40441,N_40496);
and U40746 (N_40746,N_40157,N_40452);
or U40747 (N_40747,N_40176,N_40147);
and U40748 (N_40748,N_40291,N_40262);
nor U40749 (N_40749,N_40396,N_40464);
and U40750 (N_40750,N_40013,N_40293);
nor U40751 (N_40751,N_40145,N_40030);
and U40752 (N_40752,N_40178,N_40176);
or U40753 (N_40753,N_40392,N_40307);
or U40754 (N_40754,N_40200,N_40157);
xnor U40755 (N_40755,N_40460,N_40470);
nor U40756 (N_40756,N_40105,N_40063);
or U40757 (N_40757,N_40029,N_40337);
nor U40758 (N_40758,N_40358,N_40086);
and U40759 (N_40759,N_40409,N_40086);
xor U40760 (N_40760,N_40074,N_40035);
nor U40761 (N_40761,N_40118,N_40108);
xnor U40762 (N_40762,N_40407,N_40268);
nand U40763 (N_40763,N_40247,N_40192);
or U40764 (N_40764,N_40255,N_40121);
xnor U40765 (N_40765,N_40099,N_40221);
or U40766 (N_40766,N_40346,N_40212);
nand U40767 (N_40767,N_40048,N_40238);
nand U40768 (N_40768,N_40037,N_40217);
and U40769 (N_40769,N_40389,N_40076);
xor U40770 (N_40770,N_40006,N_40412);
xnor U40771 (N_40771,N_40180,N_40476);
xnor U40772 (N_40772,N_40210,N_40290);
nor U40773 (N_40773,N_40450,N_40082);
nor U40774 (N_40774,N_40213,N_40339);
nand U40775 (N_40775,N_40431,N_40145);
and U40776 (N_40776,N_40268,N_40450);
or U40777 (N_40777,N_40449,N_40070);
or U40778 (N_40778,N_40064,N_40286);
and U40779 (N_40779,N_40425,N_40395);
xor U40780 (N_40780,N_40349,N_40029);
or U40781 (N_40781,N_40007,N_40364);
and U40782 (N_40782,N_40022,N_40422);
nor U40783 (N_40783,N_40421,N_40426);
and U40784 (N_40784,N_40128,N_40402);
nand U40785 (N_40785,N_40163,N_40284);
or U40786 (N_40786,N_40075,N_40116);
nor U40787 (N_40787,N_40486,N_40215);
xor U40788 (N_40788,N_40345,N_40169);
nor U40789 (N_40789,N_40153,N_40479);
nor U40790 (N_40790,N_40078,N_40403);
nor U40791 (N_40791,N_40180,N_40168);
xnor U40792 (N_40792,N_40048,N_40323);
nor U40793 (N_40793,N_40482,N_40109);
xor U40794 (N_40794,N_40053,N_40064);
nor U40795 (N_40795,N_40377,N_40239);
nor U40796 (N_40796,N_40184,N_40362);
and U40797 (N_40797,N_40359,N_40232);
nor U40798 (N_40798,N_40350,N_40214);
nor U40799 (N_40799,N_40375,N_40135);
xor U40800 (N_40800,N_40198,N_40455);
xnor U40801 (N_40801,N_40131,N_40206);
nor U40802 (N_40802,N_40177,N_40095);
and U40803 (N_40803,N_40208,N_40094);
nor U40804 (N_40804,N_40227,N_40065);
and U40805 (N_40805,N_40054,N_40106);
and U40806 (N_40806,N_40276,N_40057);
nand U40807 (N_40807,N_40080,N_40379);
nand U40808 (N_40808,N_40317,N_40082);
nand U40809 (N_40809,N_40036,N_40380);
nor U40810 (N_40810,N_40452,N_40305);
and U40811 (N_40811,N_40244,N_40073);
nor U40812 (N_40812,N_40410,N_40394);
or U40813 (N_40813,N_40105,N_40362);
or U40814 (N_40814,N_40143,N_40196);
nor U40815 (N_40815,N_40190,N_40234);
nor U40816 (N_40816,N_40106,N_40180);
and U40817 (N_40817,N_40087,N_40031);
xor U40818 (N_40818,N_40469,N_40095);
nand U40819 (N_40819,N_40393,N_40216);
nor U40820 (N_40820,N_40182,N_40226);
or U40821 (N_40821,N_40161,N_40117);
or U40822 (N_40822,N_40406,N_40467);
xnor U40823 (N_40823,N_40272,N_40046);
or U40824 (N_40824,N_40163,N_40468);
xnor U40825 (N_40825,N_40435,N_40229);
nor U40826 (N_40826,N_40174,N_40378);
nor U40827 (N_40827,N_40282,N_40161);
nor U40828 (N_40828,N_40220,N_40137);
nor U40829 (N_40829,N_40280,N_40467);
and U40830 (N_40830,N_40393,N_40177);
nand U40831 (N_40831,N_40217,N_40163);
or U40832 (N_40832,N_40477,N_40069);
and U40833 (N_40833,N_40454,N_40307);
and U40834 (N_40834,N_40355,N_40369);
nor U40835 (N_40835,N_40144,N_40278);
xor U40836 (N_40836,N_40121,N_40093);
or U40837 (N_40837,N_40282,N_40027);
xnor U40838 (N_40838,N_40059,N_40116);
and U40839 (N_40839,N_40398,N_40236);
nand U40840 (N_40840,N_40299,N_40023);
nor U40841 (N_40841,N_40252,N_40211);
and U40842 (N_40842,N_40189,N_40331);
nor U40843 (N_40843,N_40226,N_40365);
nand U40844 (N_40844,N_40142,N_40235);
xor U40845 (N_40845,N_40101,N_40342);
xor U40846 (N_40846,N_40251,N_40253);
or U40847 (N_40847,N_40077,N_40130);
xor U40848 (N_40848,N_40169,N_40178);
or U40849 (N_40849,N_40288,N_40398);
nor U40850 (N_40850,N_40089,N_40206);
and U40851 (N_40851,N_40060,N_40376);
nor U40852 (N_40852,N_40333,N_40478);
nor U40853 (N_40853,N_40286,N_40451);
xnor U40854 (N_40854,N_40145,N_40146);
xor U40855 (N_40855,N_40264,N_40012);
nor U40856 (N_40856,N_40112,N_40142);
xnor U40857 (N_40857,N_40434,N_40155);
xnor U40858 (N_40858,N_40404,N_40128);
xor U40859 (N_40859,N_40105,N_40314);
nand U40860 (N_40860,N_40432,N_40022);
xor U40861 (N_40861,N_40331,N_40045);
and U40862 (N_40862,N_40111,N_40378);
nor U40863 (N_40863,N_40107,N_40335);
xnor U40864 (N_40864,N_40090,N_40026);
xor U40865 (N_40865,N_40457,N_40496);
or U40866 (N_40866,N_40403,N_40171);
or U40867 (N_40867,N_40358,N_40423);
and U40868 (N_40868,N_40398,N_40439);
nor U40869 (N_40869,N_40013,N_40035);
nor U40870 (N_40870,N_40094,N_40465);
and U40871 (N_40871,N_40250,N_40028);
xor U40872 (N_40872,N_40422,N_40307);
or U40873 (N_40873,N_40143,N_40193);
or U40874 (N_40874,N_40338,N_40055);
nand U40875 (N_40875,N_40469,N_40434);
xnor U40876 (N_40876,N_40370,N_40242);
nor U40877 (N_40877,N_40268,N_40317);
xor U40878 (N_40878,N_40231,N_40388);
nand U40879 (N_40879,N_40310,N_40238);
or U40880 (N_40880,N_40423,N_40344);
nor U40881 (N_40881,N_40407,N_40485);
xor U40882 (N_40882,N_40030,N_40253);
or U40883 (N_40883,N_40225,N_40419);
and U40884 (N_40884,N_40360,N_40067);
and U40885 (N_40885,N_40302,N_40372);
and U40886 (N_40886,N_40402,N_40337);
nor U40887 (N_40887,N_40300,N_40266);
and U40888 (N_40888,N_40467,N_40390);
nand U40889 (N_40889,N_40384,N_40299);
and U40890 (N_40890,N_40486,N_40066);
or U40891 (N_40891,N_40051,N_40459);
or U40892 (N_40892,N_40499,N_40493);
xnor U40893 (N_40893,N_40006,N_40490);
or U40894 (N_40894,N_40427,N_40391);
nor U40895 (N_40895,N_40072,N_40020);
and U40896 (N_40896,N_40114,N_40007);
xor U40897 (N_40897,N_40355,N_40326);
or U40898 (N_40898,N_40158,N_40054);
nor U40899 (N_40899,N_40156,N_40007);
xor U40900 (N_40900,N_40190,N_40122);
or U40901 (N_40901,N_40368,N_40350);
nand U40902 (N_40902,N_40158,N_40424);
nor U40903 (N_40903,N_40163,N_40120);
nor U40904 (N_40904,N_40211,N_40155);
nor U40905 (N_40905,N_40471,N_40246);
and U40906 (N_40906,N_40125,N_40464);
or U40907 (N_40907,N_40052,N_40439);
xnor U40908 (N_40908,N_40105,N_40303);
and U40909 (N_40909,N_40276,N_40392);
nor U40910 (N_40910,N_40163,N_40129);
and U40911 (N_40911,N_40225,N_40444);
nand U40912 (N_40912,N_40019,N_40055);
or U40913 (N_40913,N_40038,N_40367);
nand U40914 (N_40914,N_40115,N_40006);
or U40915 (N_40915,N_40361,N_40373);
nand U40916 (N_40916,N_40205,N_40309);
and U40917 (N_40917,N_40143,N_40149);
xor U40918 (N_40918,N_40302,N_40417);
xnor U40919 (N_40919,N_40432,N_40123);
nand U40920 (N_40920,N_40235,N_40372);
and U40921 (N_40921,N_40033,N_40424);
nor U40922 (N_40922,N_40017,N_40334);
and U40923 (N_40923,N_40428,N_40064);
xor U40924 (N_40924,N_40131,N_40104);
or U40925 (N_40925,N_40394,N_40219);
nor U40926 (N_40926,N_40132,N_40032);
or U40927 (N_40927,N_40224,N_40070);
or U40928 (N_40928,N_40388,N_40313);
and U40929 (N_40929,N_40201,N_40232);
nor U40930 (N_40930,N_40056,N_40309);
and U40931 (N_40931,N_40137,N_40095);
nor U40932 (N_40932,N_40423,N_40048);
or U40933 (N_40933,N_40244,N_40357);
or U40934 (N_40934,N_40231,N_40184);
nor U40935 (N_40935,N_40028,N_40342);
and U40936 (N_40936,N_40181,N_40067);
xor U40937 (N_40937,N_40034,N_40367);
and U40938 (N_40938,N_40383,N_40465);
and U40939 (N_40939,N_40026,N_40371);
xnor U40940 (N_40940,N_40126,N_40396);
or U40941 (N_40941,N_40249,N_40110);
nand U40942 (N_40942,N_40435,N_40395);
xnor U40943 (N_40943,N_40222,N_40370);
nor U40944 (N_40944,N_40017,N_40467);
xor U40945 (N_40945,N_40463,N_40480);
nor U40946 (N_40946,N_40283,N_40448);
nor U40947 (N_40947,N_40483,N_40378);
xor U40948 (N_40948,N_40490,N_40309);
or U40949 (N_40949,N_40310,N_40366);
nand U40950 (N_40950,N_40247,N_40016);
xor U40951 (N_40951,N_40074,N_40217);
xnor U40952 (N_40952,N_40461,N_40275);
nand U40953 (N_40953,N_40217,N_40485);
or U40954 (N_40954,N_40162,N_40226);
xnor U40955 (N_40955,N_40073,N_40012);
and U40956 (N_40956,N_40264,N_40465);
nor U40957 (N_40957,N_40104,N_40072);
nand U40958 (N_40958,N_40408,N_40081);
xor U40959 (N_40959,N_40261,N_40047);
nor U40960 (N_40960,N_40091,N_40423);
or U40961 (N_40961,N_40150,N_40108);
xnor U40962 (N_40962,N_40379,N_40381);
and U40963 (N_40963,N_40390,N_40210);
and U40964 (N_40964,N_40222,N_40361);
xnor U40965 (N_40965,N_40473,N_40242);
nand U40966 (N_40966,N_40068,N_40195);
nand U40967 (N_40967,N_40022,N_40109);
xor U40968 (N_40968,N_40100,N_40383);
or U40969 (N_40969,N_40243,N_40318);
or U40970 (N_40970,N_40499,N_40153);
xnor U40971 (N_40971,N_40202,N_40008);
nor U40972 (N_40972,N_40330,N_40419);
xnor U40973 (N_40973,N_40069,N_40003);
nand U40974 (N_40974,N_40276,N_40400);
or U40975 (N_40975,N_40361,N_40032);
nor U40976 (N_40976,N_40458,N_40491);
or U40977 (N_40977,N_40021,N_40027);
and U40978 (N_40978,N_40139,N_40167);
nand U40979 (N_40979,N_40401,N_40266);
nor U40980 (N_40980,N_40327,N_40422);
and U40981 (N_40981,N_40390,N_40140);
or U40982 (N_40982,N_40495,N_40458);
nand U40983 (N_40983,N_40149,N_40374);
and U40984 (N_40984,N_40089,N_40125);
nand U40985 (N_40985,N_40145,N_40489);
xnor U40986 (N_40986,N_40157,N_40327);
or U40987 (N_40987,N_40052,N_40326);
nor U40988 (N_40988,N_40042,N_40070);
nor U40989 (N_40989,N_40308,N_40035);
or U40990 (N_40990,N_40154,N_40011);
nor U40991 (N_40991,N_40047,N_40097);
or U40992 (N_40992,N_40434,N_40395);
nand U40993 (N_40993,N_40336,N_40406);
xnor U40994 (N_40994,N_40156,N_40243);
nor U40995 (N_40995,N_40186,N_40103);
xor U40996 (N_40996,N_40487,N_40192);
and U40997 (N_40997,N_40069,N_40090);
or U40998 (N_40998,N_40162,N_40167);
xor U40999 (N_40999,N_40432,N_40313);
xnor U41000 (N_41000,N_40832,N_40611);
or U41001 (N_41001,N_40675,N_40941);
xor U41002 (N_41002,N_40501,N_40576);
and U41003 (N_41003,N_40886,N_40932);
nor U41004 (N_41004,N_40849,N_40503);
or U41005 (N_41005,N_40566,N_40796);
nor U41006 (N_41006,N_40734,N_40936);
nor U41007 (N_41007,N_40723,N_40631);
and U41008 (N_41008,N_40604,N_40909);
and U41009 (N_41009,N_40993,N_40585);
or U41010 (N_41010,N_40568,N_40910);
xnor U41011 (N_41011,N_40882,N_40749);
nand U41012 (N_41012,N_40916,N_40696);
or U41013 (N_41013,N_40816,N_40607);
or U41014 (N_41014,N_40866,N_40740);
or U41015 (N_41015,N_40697,N_40800);
xor U41016 (N_41016,N_40763,N_40814);
xor U41017 (N_41017,N_40807,N_40798);
nor U41018 (N_41018,N_40515,N_40962);
nand U41019 (N_41019,N_40514,N_40757);
or U41020 (N_41020,N_40965,N_40660);
nor U41021 (N_41021,N_40770,N_40843);
xnor U41022 (N_41022,N_40715,N_40626);
xnor U41023 (N_41023,N_40929,N_40971);
nor U41024 (N_41024,N_40803,N_40574);
nor U41025 (N_41025,N_40949,N_40655);
nor U41026 (N_41026,N_40583,N_40957);
or U41027 (N_41027,N_40511,N_40877);
xor U41028 (N_41028,N_40893,N_40592);
or U41029 (N_41029,N_40784,N_40548);
nor U41030 (N_41030,N_40775,N_40711);
nand U41031 (N_41031,N_40658,N_40808);
and U41032 (N_41032,N_40772,N_40978);
xnor U41033 (N_41033,N_40721,N_40828);
and U41034 (N_41034,N_40633,N_40812);
nand U41035 (N_41035,N_40788,N_40533);
xor U41036 (N_41036,N_40844,N_40799);
nand U41037 (N_41037,N_40751,N_40878);
or U41038 (N_41038,N_40516,N_40705);
nand U41039 (N_41039,N_40954,N_40509);
and U41040 (N_41040,N_40989,N_40654);
or U41041 (N_41041,N_40864,N_40896);
nor U41042 (N_41042,N_40756,N_40593);
nand U41043 (N_41043,N_40513,N_40676);
nand U41044 (N_41044,N_40752,N_40507);
and U41045 (N_41045,N_40958,N_40943);
xnor U41046 (N_41046,N_40914,N_40709);
nor U41047 (N_41047,N_40806,N_40739);
and U41048 (N_41048,N_40824,N_40689);
nor U41049 (N_41049,N_40968,N_40865);
nor U41050 (N_41050,N_40570,N_40905);
nor U41051 (N_41051,N_40947,N_40918);
or U41052 (N_41052,N_40782,N_40616);
nand U41053 (N_41053,N_40945,N_40771);
xnor U41054 (N_41054,N_40794,N_40665);
xnor U41055 (N_41055,N_40783,N_40925);
nor U41056 (N_41056,N_40768,N_40950);
xnor U41057 (N_41057,N_40678,N_40541);
or U41058 (N_41058,N_40876,N_40531);
and U41059 (N_41059,N_40935,N_40535);
nor U41060 (N_41060,N_40744,N_40736);
xor U41061 (N_41061,N_40999,N_40786);
nand U41062 (N_41062,N_40617,N_40577);
xnor U41063 (N_41063,N_40995,N_40746);
nand U41064 (N_41064,N_40933,N_40912);
xnor U41065 (N_41065,N_40712,N_40597);
nor U41066 (N_41066,N_40851,N_40815);
nand U41067 (N_41067,N_40765,N_40764);
nand U41068 (N_41068,N_40520,N_40672);
nor U41069 (N_41069,N_40873,N_40902);
and U41070 (N_41070,N_40661,N_40901);
nor U41071 (N_41071,N_40946,N_40990);
or U41072 (N_41072,N_40967,N_40547);
nand U41073 (N_41073,N_40567,N_40526);
nand U41074 (N_41074,N_40907,N_40748);
nor U41075 (N_41075,N_40716,N_40883);
and U41076 (N_41076,N_40701,N_40899);
nor U41077 (N_41077,N_40545,N_40963);
nand U41078 (N_41078,N_40982,N_40802);
or U41079 (N_41079,N_40699,N_40557);
nor U41080 (N_41080,N_40829,N_40924);
or U41081 (N_41081,N_40892,N_40761);
nand U41082 (N_41082,N_40801,N_40836);
nor U41083 (N_41083,N_40826,N_40820);
or U41084 (N_41084,N_40774,N_40522);
and U41085 (N_41085,N_40894,N_40542);
nand U41086 (N_41086,N_40741,N_40972);
xnor U41087 (N_41087,N_40969,N_40966);
nor U41088 (N_41088,N_40529,N_40662);
xnor U41089 (N_41089,N_40641,N_40931);
or U41090 (N_41090,N_40625,N_40605);
xor U41091 (N_41091,N_40805,N_40858);
nand U41092 (N_41092,N_40781,N_40578);
xnor U41093 (N_41093,N_40992,N_40621);
nor U41094 (N_41094,N_40841,N_40952);
xor U41095 (N_41095,N_40615,N_40939);
nor U41096 (N_41096,N_40599,N_40731);
nand U41097 (N_41097,N_40644,N_40732);
and U41098 (N_41098,N_40818,N_40964);
nor U41099 (N_41099,N_40955,N_40906);
nor U41100 (N_41100,N_40852,N_40730);
and U41101 (N_41101,N_40609,N_40543);
and U41102 (N_41102,N_40504,N_40890);
and U41103 (N_41103,N_40667,N_40789);
and U41104 (N_41104,N_40528,N_40724);
nor U41105 (N_41105,N_40759,N_40793);
nor U41106 (N_41106,N_40512,N_40652);
nand U41107 (N_41107,N_40629,N_40944);
or U41108 (N_41108,N_40600,N_40970);
nand U41109 (N_41109,N_40853,N_40663);
or U41110 (N_41110,N_40839,N_40827);
or U41111 (N_41111,N_40536,N_40551);
nand U41112 (N_41112,N_40986,N_40707);
nor U41113 (N_41113,N_40938,N_40926);
or U41114 (N_41114,N_40645,N_40779);
and U41115 (N_41115,N_40842,N_40603);
or U41116 (N_41116,N_40673,N_40552);
or U41117 (N_41117,N_40527,N_40737);
or U41118 (N_41118,N_40703,N_40684);
and U41119 (N_41119,N_40976,N_40722);
xor U41120 (N_41120,N_40871,N_40563);
and U41121 (N_41121,N_40595,N_40564);
and U41122 (N_41122,N_40884,N_40837);
or U41123 (N_41123,N_40694,N_40817);
or U41124 (N_41124,N_40868,N_40917);
nor U41125 (N_41125,N_40650,N_40908);
nor U41126 (N_41126,N_40558,N_40635);
and U41127 (N_41127,N_40643,N_40636);
nor U41128 (N_41128,N_40750,N_40572);
and U41129 (N_41129,N_40614,N_40885);
xor U41130 (N_41130,N_40863,N_40881);
xnor U41131 (N_41131,N_40769,N_40623);
or U41132 (N_41132,N_40546,N_40666);
or U41133 (N_41133,N_40695,N_40897);
nand U41134 (N_41134,N_40948,N_40632);
nand U41135 (N_41135,N_40590,N_40860);
nor U41136 (N_41136,N_40973,N_40559);
or U41137 (N_41137,N_40647,N_40523);
or U41138 (N_41138,N_40525,N_40555);
nor U41139 (N_41139,N_40717,N_40587);
nor U41140 (N_41140,N_40586,N_40638);
nand U41141 (N_41141,N_40726,N_40620);
or U41142 (N_41142,N_40961,N_40693);
xor U41143 (N_41143,N_40813,N_40875);
nand U41144 (N_41144,N_40668,N_40997);
or U41145 (N_41145,N_40857,N_40704);
xnor U41146 (N_41146,N_40561,N_40735);
nor U41147 (N_41147,N_40619,N_40940);
or U41148 (N_41148,N_40510,N_40974);
or U41149 (N_41149,N_40911,N_40669);
nand U41150 (N_41150,N_40872,N_40766);
nor U41151 (N_41151,N_40698,N_40942);
nor U41152 (N_41152,N_40606,N_40549);
and U41153 (N_41153,N_40760,N_40729);
nor U41154 (N_41154,N_40983,N_40710);
and U41155 (N_41155,N_40919,N_40975);
or U41156 (N_41156,N_40850,N_40582);
nand U41157 (N_41157,N_40904,N_40553);
or U41158 (N_41158,N_40825,N_40618);
and U41159 (N_41159,N_40854,N_40856);
nor U41160 (N_41160,N_40500,N_40659);
or U41161 (N_41161,N_40708,N_40996);
xor U41162 (N_41162,N_40791,N_40888);
and U41163 (N_41163,N_40819,N_40679);
and U41164 (N_41164,N_40589,N_40822);
or U41165 (N_41165,N_40637,N_40519);
and U41166 (N_41166,N_40508,N_40922);
nor U41167 (N_41167,N_40874,N_40861);
xnor U41168 (N_41168,N_40517,N_40670);
nor U41169 (N_41169,N_40728,N_40639);
nand U41170 (N_41170,N_40648,N_40534);
or U41171 (N_41171,N_40687,N_40811);
and U41172 (N_41172,N_40706,N_40887);
xnor U41173 (N_41173,N_40700,N_40640);
or U41174 (N_41174,N_40714,N_40846);
and U41175 (N_41175,N_40677,N_40569);
nand U41176 (N_41176,N_40530,N_40506);
and U41177 (N_41177,N_40573,N_40753);
or U41178 (N_41178,N_40634,N_40988);
and U41179 (N_41179,N_40594,N_40930);
nand U41180 (N_41180,N_40718,N_40934);
xnor U41181 (N_41181,N_40610,N_40745);
or U41182 (N_41182,N_40580,N_40538);
nand U41183 (N_41183,N_40994,N_40550);
nand U41184 (N_41184,N_40981,N_40762);
nand U41185 (N_41185,N_40571,N_40845);
or U41186 (N_41186,N_40521,N_40767);
xor U41187 (N_41187,N_40518,N_40862);
or U41188 (N_41188,N_40537,N_40608);
or U41189 (N_41189,N_40977,N_40804);
nand U41190 (N_41190,N_40821,N_40838);
nand U41191 (N_41191,N_40747,N_40913);
xnor U41192 (N_41192,N_40720,N_40776);
nand U41193 (N_41193,N_40831,N_40560);
nand U41194 (N_41194,N_40692,N_40979);
nor U41195 (N_41195,N_40681,N_40575);
or U41196 (N_41196,N_40780,N_40649);
nor U41197 (N_41197,N_40953,N_40664);
xnor U41198 (N_41198,N_40584,N_40880);
xor U41199 (N_41199,N_40937,N_40630);
and U41200 (N_41200,N_40612,N_40562);
xor U41201 (N_41201,N_40960,N_40727);
or U41202 (N_41202,N_40682,N_40987);
nor U41203 (N_41203,N_40556,N_40833);
nor U41204 (N_41204,N_40702,N_40847);
nor U41205 (N_41205,N_40688,N_40898);
or U41206 (N_41206,N_40830,N_40502);
nand U41207 (N_41207,N_40674,N_40581);
or U41208 (N_41208,N_40920,N_40624);
xnor U41209 (N_41209,N_40835,N_40980);
nand U41210 (N_41210,N_40959,N_40869);
nor U41211 (N_41211,N_40809,N_40540);
nand U41212 (N_41212,N_40598,N_40758);
nor U41213 (N_41213,N_40985,N_40915);
xor U41214 (N_41214,N_40601,N_40596);
nand U41215 (N_41215,N_40628,N_40642);
xor U41216 (N_41216,N_40591,N_40956);
xor U41217 (N_41217,N_40787,N_40834);
nand U41218 (N_41218,N_40792,N_40778);
or U41219 (N_41219,N_40646,N_40903);
xnor U41220 (N_41220,N_40733,N_40773);
or U41221 (N_41221,N_40622,N_40588);
nor U41222 (N_41222,N_40719,N_40505);
and U41223 (N_41223,N_40653,N_40754);
and U41224 (N_41224,N_40565,N_40686);
xor U41225 (N_41225,N_40900,N_40785);
or U41226 (N_41226,N_40613,N_40657);
nand U41227 (N_41227,N_40691,N_40544);
and U41228 (N_41228,N_40870,N_40742);
and U41229 (N_41229,N_40651,N_40738);
and U41230 (N_41230,N_40998,N_40627);
or U41231 (N_41231,N_40777,N_40797);
or U41232 (N_41232,N_40810,N_40680);
and U41233 (N_41233,N_40671,N_40713);
nand U41234 (N_41234,N_40656,N_40690);
and U41235 (N_41235,N_40855,N_40579);
or U41236 (N_41236,N_40524,N_40895);
nand U41237 (N_41237,N_40889,N_40532);
nor U41238 (N_41238,N_40823,N_40554);
xor U41239 (N_41239,N_40848,N_40790);
and U41240 (N_41240,N_40755,N_40991);
xor U41241 (N_41241,N_40795,N_40879);
nor U41242 (N_41242,N_40984,N_40859);
and U41243 (N_41243,N_40685,N_40867);
nand U41244 (N_41244,N_40951,N_40602);
xor U41245 (N_41245,N_40539,N_40840);
or U41246 (N_41246,N_40928,N_40891);
xnor U41247 (N_41247,N_40923,N_40683);
xor U41248 (N_41248,N_40725,N_40927);
nor U41249 (N_41249,N_40921,N_40743);
nor U41250 (N_41250,N_40670,N_40814);
or U41251 (N_41251,N_40679,N_40869);
nand U41252 (N_41252,N_40937,N_40584);
and U41253 (N_41253,N_40929,N_40530);
or U41254 (N_41254,N_40630,N_40767);
and U41255 (N_41255,N_40891,N_40904);
nor U41256 (N_41256,N_40946,N_40786);
nor U41257 (N_41257,N_40907,N_40958);
nor U41258 (N_41258,N_40796,N_40926);
xnor U41259 (N_41259,N_40598,N_40939);
or U41260 (N_41260,N_40849,N_40528);
nor U41261 (N_41261,N_40695,N_40527);
and U41262 (N_41262,N_40881,N_40575);
nand U41263 (N_41263,N_40911,N_40612);
and U41264 (N_41264,N_40773,N_40764);
and U41265 (N_41265,N_40545,N_40787);
nand U41266 (N_41266,N_40560,N_40952);
xor U41267 (N_41267,N_40573,N_40719);
or U41268 (N_41268,N_40588,N_40637);
or U41269 (N_41269,N_40817,N_40758);
nor U41270 (N_41270,N_40679,N_40703);
xnor U41271 (N_41271,N_40763,N_40555);
nor U41272 (N_41272,N_40645,N_40933);
xor U41273 (N_41273,N_40813,N_40543);
nor U41274 (N_41274,N_40974,N_40903);
nor U41275 (N_41275,N_40650,N_40632);
or U41276 (N_41276,N_40976,N_40665);
or U41277 (N_41277,N_40738,N_40796);
nor U41278 (N_41278,N_40811,N_40789);
and U41279 (N_41279,N_40556,N_40990);
nor U41280 (N_41280,N_40780,N_40947);
nor U41281 (N_41281,N_40965,N_40729);
and U41282 (N_41282,N_40566,N_40810);
and U41283 (N_41283,N_40748,N_40621);
nor U41284 (N_41284,N_40642,N_40668);
nand U41285 (N_41285,N_40920,N_40809);
or U41286 (N_41286,N_40966,N_40808);
xor U41287 (N_41287,N_40612,N_40688);
or U41288 (N_41288,N_40559,N_40853);
nor U41289 (N_41289,N_40908,N_40744);
xor U41290 (N_41290,N_40994,N_40596);
and U41291 (N_41291,N_40573,N_40994);
nor U41292 (N_41292,N_40731,N_40704);
xor U41293 (N_41293,N_40862,N_40981);
and U41294 (N_41294,N_40971,N_40774);
and U41295 (N_41295,N_40623,N_40702);
or U41296 (N_41296,N_40747,N_40572);
nor U41297 (N_41297,N_40697,N_40930);
or U41298 (N_41298,N_40712,N_40513);
and U41299 (N_41299,N_40913,N_40964);
or U41300 (N_41300,N_40938,N_40785);
and U41301 (N_41301,N_40620,N_40713);
xor U41302 (N_41302,N_40695,N_40608);
xnor U41303 (N_41303,N_40723,N_40954);
nand U41304 (N_41304,N_40771,N_40902);
nand U41305 (N_41305,N_40605,N_40913);
nand U41306 (N_41306,N_40535,N_40946);
and U41307 (N_41307,N_40546,N_40554);
nor U41308 (N_41308,N_40656,N_40712);
nand U41309 (N_41309,N_40544,N_40646);
xor U41310 (N_41310,N_40879,N_40618);
xnor U41311 (N_41311,N_40582,N_40833);
xnor U41312 (N_41312,N_40627,N_40553);
or U41313 (N_41313,N_40660,N_40567);
or U41314 (N_41314,N_40740,N_40518);
and U41315 (N_41315,N_40626,N_40523);
or U41316 (N_41316,N_40823,N_40530);
nand U41317 (N_41317,N_40537,N_40915);
nand U41318 (N_41318,N_40607,N_40896);
nand U41319 (N_41319,N_40727,N_40780);
xnor U41320 (N_41320,N_40770,N_40535);
xnor U41321 (N_41321,N_40639,N_40970);
or U41322 (N_41322,N_40839,N_40968);
nand U41323 (N_41323,N_40515,N_40676);
and U41324 (N_41324,N_40630,N_40657);
nor U41325 (N_41325,N_40604,N_40871);
nand U41326 (N_41326,N_40599,N_40895);
nand U41327 (N_41327,N_40514,N_40886);
nand U41328 (N_41328,N_40638,N_40534);
xor U41329 (N_41329,N_40884,N_40612);
or U41330 (N_41330,N_40818,N_40536);
xor U41331 (N_41331,N_40709,N_40744);
xnor U41332 (N_41332,N_40649,N_40836);
nand U41333 (N_41333,N_40578,N_40574);
and U41334 (N_41334,N_40622,N_40858);
xor U41335 (N_41335,N_40985,N_40804);
and U41336 (N_41336,N_40783,N_40585);
nand U41337 (N_41337,N_40912,N_40712);
and U41338 (N_41338,N_40913,N_40867);
xor U41339 (N_41339,N_40862,N_40899);
nand U41340 (N_41340,N_40879,N_40814);
nand U41341 (N_41341,N_40859,N_40747);
and U41342 (N_41342,N_40804,N_40983);
and U41343 (N_41343,N_40931,N_40767);
and U41344 (N_41344,N_40931,N_40599);
and U41345 (N_41345,N_40838,N_40730);
or U41346 (N_41346,N_40582,N_40921);
and U41347 (N_41347,N_40689,N_40897);
xnor U41348 (N_41348,N_40641,N_40962);
nand U41349 (N_41349,N_40977,N_40916);
or U41350 (N_41350,N_40924,N_40839);
xor U41351 (N_41351,N_40900,N_40929);
nand U41352 (N_41352,N_40961,N_40702);
or U41353 (N_41353,N_40976,N_40834);
and U41354 (N_41354,N_40934,N_40914);
xor U41355 (N_41355,N_40785,N_40584);
or U41356 (N_41356,N_40879,N_40925);
or U41357 (N_41357,N_40603,N_40811);
xor U41358 (N_41358,N_40613,N_40920);
xor U41359 (N_41359,N_40693,N_40767);
and U41360 (N_41360,N_40962,N_40957);
and U41361 (N_41361,N_40520,N_40675);
or U41362 (N_41362,N_40929,N_40603);
xor U41363 (N_41363,N_40965,N_40871);
and U41364 (N_41364,N_40584,N_40888);
nor U41365 (N_41365,N_40664,N_40702);
nor U41366 (N_41366,N_40564,N_40730);
nand U41367 (N_41367,N_40826,N_40582);
nor U41368 (N_41368,N_40682,N_40973);
nand U41369 (N_41369,N_40626,N_40722);
or U41370 (N_41370,N_40966,N_40933);
and U41371 (N_41371,N_40827,N_40597);
or U41372 (N_41372,N_40965,N_40888);
or U41373 (N_41373,N_40600,N_40872);
nor U41374 (N_41374,N_40940,N_40576);
nand U41375 (N_41375,N_40646,N_40935);
nor U41376 (N_41376,N_40918,N_40772);
and U41377 (N_41377,N_40581,N_40893);
and U41378 (N_41378,N_40944,N_40996);
nand U41379 (N_41379,N_40725,N_40618);
and U41380 (N_41380,N_40793,N_40802);
nor U41381 (N_41381,N_40904,N_40809);
nor U41382 (N_41382,N_40669,N_40699);
nor U41383 (N_41383,N_40901,N_40515);
nor U41384 (N_41384,N_40859,N_40887);
nand U41385 (N_41385,N_40883,N_40881);
or U41386 (N_41386,N_40822,N_40563);
or U41387 (N_41387,N_40594,N_40758);
nor U41388 (N_41388,N_40842,N_40615);
and U41389 (N_41389,N_40757,N_40786);
or U41390 (N_41390,N_40595,N_40763);
and U41391 (N_41391,N_40546,N_40813);
nor U41392 (N_41392,N_40534,N_40517);
nor U41393 (N_41393,N_40508,N_40847);
or U41394 (N_41394,N_40914,N_40797);
xnor U41395 (N_41395,N_40754,N_40940);
xor U41396 (N_41396,N_40545,N_40708);
or U41397 (N_41397,N_40944,N_40840);
or U41398 (N_41398,N_40583,N_40773);
and U41399 (N_41399,N_40978,N_40643);
nor U41400 (N_41400,N_40705,N_40661);
and U41401 (N_41401,N_40955,N_40592);
and U41402 (N_41402,N_40988,N_40582);
and U41403 (N_41403,N_40553,N_40794);
nand U41404 (N_41404,N_40912,N_40899);
nor U41405 (N_41405,N_40567,N_40644);
nor U41406 (N_41406,N_40989,N_40726);
or U41407 (N_41407,N_40723,N_40994);
xnor U41408 (N_41408,N_40547,N_40964);
or U41409 (N_41409,N_40890,N_40541);
xor U41410 (N_41410,N_40793,N_40878);
xor U41411 (N_41411,N_40533,N_40993);
and U41412 (N_41412,N_40896,N_40748);
nand U41413 (N_41413,N_40767,N_40717);
xnor U41414 (N_41414,N_40923,N_40976);
nand U41415 (N_41415,N_40876,N_40833);
or U41416 (N_41416,N_40900,N_40958);
nor U41417 (N_41417,N_40742,N_40625);
nor U41418 (N_41418,N_40838,N_40643);
or U41419 (N_41419,N_40927,N_40784);
xnor U41420 (N_41420,N_40519,N_40853);
nor U41421 (N_41421,N_40934,N_40789);
xor U41422 (N_41422,N_40576,N_40674);
xnor U41423 (N_41423,N_40913,N_40763);
nand U41424 (N_41424,N_40686,N_40695);
and U41425 (N_41425,N_40773,N_40867);
and U41426 (N_41426,N_40785,N_40564);
xnor U41427 (N_41427,N_40966,N_40998);
nand U41428 (N_41428,N_40541,N_40918);
or U41429 (N_41429,N_40543,N_40979);
or U41430 (N_41430,N_40906,N_40966);
nand U41431 (N_41431,N_40705,N_40605);
nand U41432 (N_41432,N_40972,N_40776);
and U41433 (N_41433,N_40673,N_40759);
nand U41434 (N_41434,N_40530,N_40538);
nor U41435 (N_41435,N_40610,N_40850);
or U41436 (N_41436,N_40630,N_40833);
nor U41437 (N_41437,N_40824,N_40581);
nand U41438 (N_41438,N_40709,N_40593);
nor U41439 (N_41439,N_40592,N_40670);
and U41440 (N_41440,N_40575,N_40724);
and U41441 (N_41441,N_40506,N_40995);
nor U41442 (N_41442,N_40877,N_40767);
xor U41443 (N_41443,N_40883,N_40680);
and U41444 (N_41444,N_40776,N_40914);
xnor U41445 (N_41445,N_40524,N_40744);
xor U41446 (N_41446,N_40543,N_40670);
xnor U41447 (N_41447,N_40632,N_40723);
and U41448 (N_41448,N_40769,N_40562);
and U41449 (N_41449,N_40589,N_40818);
nand U41450 (N_41450,N_40958,N_40648);
and U41451 (N_41451,N_40821,N_40615);
and U41452 (N_41452,N_40848,N_40947);
and U41453 (N_41453,N_40713,N_40797);
and U41454 (N_41454,N_40989,N_40579);
xnor U41455 (N_41455,N_40810,N_40803);
nand U41456 (N_41456,N_40629,N_40787);
and U41457 (N_41457,N_40997,N_40513);
or U41458 (N_41458,N_40812,N_40835);
nand U41459 (N_41459,N_40995,N_40821);
or U41460 (N_41460,N_40670,N_40601);
and U41461 (N_41461,N_40913,N_40587);
nor U41462 (N_41462,N_40944,N_40874);
and U41463 (N_41463,N_40570,N_40572);
nor U41464 (N_41464,N_40590,N_40683);
or U41465 (N_41465,N_40988,N_40640);
and U41466 (N_41466,N_40591,N_40554);
nand U41467 (N_41467,N_40915,N_40863);
xnor U41468 (N_41468,N_40700,N_40604);
xnor U41469 (N_41469,N_40565,N_40998);
and U41470 (N_41470,N_40756,N_40983);
nor U41471 (N_41471,N_40574,N_40625);
xor U41472 (N_41472,N_40617,N_40656);
or U41473 (N_41473,N_40936,N_40917);
nand U41474 (N_41474,N_40850,N_40796);
or U41475 (N_41475,N_40566,N_40722);
or U41476 (N_41476,N_40832,N_40620);
nand U41477 (N_41477,N_40782,N_40792);
or U41478 (N_41478,N_40888,N_40556);
nand U41479 (N_41479,N_40595,N_40664);
or U41480 (N_41480,N_40560,N_40606);
nand U41481 (N_41481,N_40523,N_40956);
nor U41482 (N_41482,N_40544,N_40878);
xor U41483 (N_41483,N_40962,N_40948);
or U41484 (N_41484,N_40952,N_40503);
and U41485 (N_41485,N_40524,N_40643);
and U41486 (N_41486,N_40597,N_40968);
xor U41487 (N_41487,N_40907,N_40503);
nand U41488 (N_41488,N_40696,N_40896);
nand U41489 (N_41489,N_40668,N_40916);
xnor U41490 (N_41490,N_40931,N_40503);
nand U41491 (N_41491,N_40561,N_40595);
and U41492 (N_41492,N_40711,N_40736);
nand U41493 (N_41493,N_40801,N_40992);
xor U41494 (N_41494,N_40633,N_40814);
nor U41495 (N_41495,N_40759,N_40705);
nand U41496 (N_41496,N_40674,N_40896);
and U41497 (N_41497,N_40515,N_40969);
xnor U41498 (N_41498,N_40744,N_40620);
and U41499 (N_41499,N_40938,N_40702);
nand U41500 (N_41500,N_41213,N_41379);
nor U41501 (N_41501,N_41385,N_41249);
or U41502 (N_41502,N_41287,N_41161);
xnor U41503 (N_41503,N_41234,N_41128);
or U41504 (N_41504,N_41283,N_41009);
nor U41505 (N_41505,N_41433,N_41138);
and U41506 (N_41506,N_41069,N_41493);
and U41507 (N_41507,N_41359,N_41321);
xor U41508 (N_41508,N_41457,N_41084);
and U41509 (N_41509,N_41278,N_41479);
or U41510 (N_41510,N_41390,N_41290);
and U41511 (N_41511,N_41119,N_41416);
nor U41512 (N_41512,N_41118,N_41004);
nor U41513 (N_41513,N_41471,N_41191);
nand U41514 (N_41514,N_41354,N_41149);
and U41515 (N_41515,N_41075,N_41328);
nand U41516 (N_41516,N_41398,N_41150);
or U41517 (N_41517,N_41061,N_41350);
xnor U41518 (N_41518,N_41269,N_41057);
nand U41519 (N_41519,N_41008,N_41243);
xor U41520 (N_41520,N_41233,N_41481);
nor U41521 (N_41521,N_41248,N_41325);
nor U41522 (N_41522,N_41214,N_41116);
and U41523 (N_41523,N_41261,N_41277);
nor U41524 (N_41524,N_41216,N_41125);
xnor U41525 (N_41525,N_41142,N_41303);
xnor U41526 (N_41526,N_41068,N_41000);
nand U41527 (N_41527,N_41441,N_41336);
nor U41528 (N_41528,N_41021,N_41168);
nor U41529 (N_41529,N_41006,N_41461);
nand U41530 (N_41530,N_41268,N_41201);
nor U41531 (N_41531,N_41208,N_41204);
xor U41532 (N_41532,N_41256,N_41447);
nor U41533 (N_41533,N_41140,N_41017);
nor U41534 (N_41534,N_41245,N_41284);
nor U41535 (N_41535,N_41073,N_41473);
nand U41536 (N_41536,N_41039,N_41477);
and U41537 (N_41537,N_41356,N_41037);
nor U41538 (N_41538,N_41247,N_41423);
nand U41539 (N_41539,N_41123,N_41313);
and U41540 (N_41540,N_41023,N_41469);
and U41541 (N_41541,N_41146,N_41436);
xor U41542 (N_41542,N_41047,N_41418);
xor U41543 (N_41543,N_41242,N_41002);
nor U41544 (N_41544,N_41288,N_41485);
or U41545 (N_41545,N_41217,N_41260);
and U41546 (N_41546,N_41082,N_41252);
nand U41547 (N_41547,N_41154,N_41495);
and U41548 (N_41548,N_41387,N_41439);
xnor U41549 (N_41549,N_41368,N_41376);
or U41550 (N_41550,N_41089,N_41200);
and U41551 (N_41551,N_41169,N_41474);
xnor U41552 (N_41552,N_41352,N_41446);
xor U41553 (N_41553,N_41378,N_41113);
nand U41554 (N_41554,N_41358,N_41251);
or U41555 (N_41555,N_41177,N_41038);
nor U41556 (N_41556,N_41183,N_41312);
nor U41557 (N_41557,N_41330,N_41162);
or U41558 (N_41558,N_41266,N_41206);
nand U41559 (N_41559,N_41115,N_41155);
nand U41560 (N_41560,N_41468,N_41319);
and U41561 (N_41561,N_41148,N_41425);
nor U41562 (N_41562,N_41308,N_41417);
nand U41563 (N_41563,N_41276,N_41338);
nand U41564 (N_41564,N_41428,N_41195);
nand U41565 (N_41565,N_41431,N_41373);
and U41566 (N_41566,N_41111,N_41132);
nor U41567 (N_41567,N_41224,N_41029);
nand U41568 (N_41568,N_41483,N_41235);
nor U41569 (N_41569,N_41130,N_41406);
and U41570 (N_41570,N_41326,N_41275);
xnor U41571 (N_41571,N_41120,N_41105);
nor U41572 (N_41572,N_41059,N_41205);
xnor U41573 (N_41573,N_41136,N_41129);
xnor U41574 (N_41574,N_41335,N_41370);
xnor U41575 (N_41575,N_41094,N_41459);
nor U41576 (N_41576,N_41079,N_41221);
nor U41577 (N_41577,N_41498,N_41202);
xor U41578 (N_41578,N_41145,N_41091);
nand U41579 (N_41579,N_41391,N_41011);
or U41580 (N_41580,N_41300,N_41164);
or U41581 (N_41581,N_41380,N_41016);
and U41582 (N_41582,N_41101,N_41044);
or U41583 (N_41583,N_41371,N_41460);
or U41584 (N_41584,N_41384,N_41050);
xnor U41585 (N_41585,N_41219,N_41246);
xnor U41586 (N_41586,N_41403,N_41271);
xor U41587 (N_41587,N_41298,N_41412);
or U41588 (N_41588,N_41014,N_41365);
nand U41589 (N_41589,N_41035,N_41098);
nand U41590 (N_41590,N_41305,N_41020);
nand U41591 (N_41591,N_41315,N_41339);
or U41592 (N_41592,N_41302,N_41156);
and U41593 (N_41593,N_41426,N_41381);
nand U41594 (N_41594,N_41190,N_41215);
or U41595 (N_41595,N_41175,N_41448);
nand U41596 (N_41596,N_41063,N_41364);
or U41597 (N_41597,N_41241,N_41285);
nand U41598 (N_41598,N_41463,N_41341);
xor U41599 (N_41599,N_41184,N_41291);
or U41600 (N_41600,N_41318,N_41158);
xor U41601 (N_41601,N_41317,N_41424);
or U41602 (N_41602,N_41347,N_41244);
and U41603 (N_41603,N_41346,N_41320);
nand U41604 (N_41604,N_41258,N_41117);
nor U41605 (N_41605,N_41226,N_41332);
xor U41606 (N_41606,N_41062,N_41218);
nand U41607 (N_41607,N_41499,N_41440);
nor U41608 (N_41608,N_41452,N_41492);
nor U41609 (N_41609,N_41444,N_41421);
and U41610 (N_41610,N_41081,N_41171);
and U41611 (N_41611,N_41036,N_41345);
or U41612 (N_41612,N_41173,N_41262);
nor U41613 (N_41613,N_41222,N_41405);
and U41614 (N_41614,N_41040,N_41041);
nor U41615 (N_41615,N_41064,N_41465);
xnor U41616 (N_41616,N_41110,N_41211);
nor U41617 (N_41617,N_41311,N_41255);
or U41618 (N_41618,N_41072,N_41180);
xnor U41619 (N_41619,N_41454,N_41297);
nand U41620 (N_41620,N_41450,N_41139);
or U41621 (N_41621,N_41181,N_41170);
and U41622 (N_41622,N_41270,N_41112);
nor U41623 (N_41623,N_41394,N_41010);
nor U41624 (N_41624,N_41395,N_41099);
or U41625 (N_41625,N_41159,N_41080);
and U41626 (N_41626,N_41001,N_41455);
xnor U41627 (N_41627,N_41056,N_41259);
nor U41628 (N_41628,N_41265,N_41028);
or U41629 (N_41629,N_41489,N_41236);
or U41630 (N_41630,N_41163,N_41078);
or U41631 (N_41631,N_41323,N_41166);
and U41632 (N_41632,N_41310,N_41212);
nor U41633 (N_41633,N_41012,N_41022);
or U41634 (N_41634,N_41272,N_41147);
nand U41635 (N_41635,N_41186,N_41467);
or U41636 (N_41636,N_41487,N_41193);
and U41637 (N_41637,N_41227,N_41042);
or U41638 (N_41638,N_41176,N_41194);
and U41639 (N_41639,N_41442,N_41207);
nand U41640 (N_41640,N_41453,N_41360);
xor U41641 (N_41641,N_41470,N_41229);
or U41642 (N_41642,N_41343,N_41427);
xor U41643 (N_41643,N_41490,N_41185);
and U41644 (N_41644,N_41203,N_41296);
xor U41645 (N_41645,N_41051,N_41443);
xnor U41646 (N_41646,N_41414,N_41353);
xnor U41647 (N_41647,N_41374,N_41293);
nand U41648 (N_41648,N_41497,N_41267);
xnor U41649 (N_41649,N_41015,N_41223);
or U41650 (N_41650,N_41389,N_41102);
or U41651 (N_41651,N_41397,N_41104);
xor U41652 (N_41652,N_41400,N_41030);
or U41653 (N_41653,N_41003,N_41239);
or U41654 (N_41654,N_41209,N_41097);
nor U41655 (N_41655,N_41369,N_41449);
and U41656 (N_41656,N_41351,N_41131);
nand U41657 (N_41657,N_41299,N_41445);
nor U41658 (N_41658,N_41034,N_41337);
or U41659 (N_41659,N_41172,N_41107);
nor U41660 (N_41660,N_41486,N_41273);
nand U41661 (N_41661,N_41478,N_41114);
nor U41662 (N_41662,N_41462,N_41198);
or U41663 (N_41663,N_41349,N_41434);
nand U41664 (N_41664,N_41070,N_41342);
and U41665 (N_41665,N_41362,N_41005);
and U41666 (N_41666,N_41357,N_41077);
nand U41667 (N_41667,N_41178,N_41294);
nand U41668 (N_41668,N_41333,N_41152);
nand U41669 (N_41669,N_41157,N_41386);
xnor U41670 (N_41670,N_41438,N_41451);
and U41671 (N_41671,N_41231,N_41230);
or U41672 (N_41672,N_41088,N_41420);
xor U41673 (N_41673,N_41135,N_41188);
nand U41674 (N_41674,N_41174,N_41401);
nand U41675 (N_41675,N_41407,N_41065);
nand U41676 (N_41676,N_41415,N_41264);
nor U41677 (N_41677,N_41052,N_41491);
and U41678 (N_41678,N_41456,N_41437);
or U41679 (N_41679,N_41013,N_41060);
nor U41680 (N_41680,N_41058,N_41482);
xor U41681 (N_41681,N_41254,N_41025);
xnor U41682 (N_41682,N_41329,N_41363);
xnor U41683 (N_41683,N_41429,N_41086);
xor U41684 (N_41684,N_41432,N_41464);
or U41685 (N_41685,N_41340,N_41018);
and U41686 (N_41686,N_41309,N_41043);
xor U41687 (N_41687,N_41192,N_41327);
nor U41688 (N_41688,N_41377,N_41053);
nor U41689 (N_41689,N_41331,N_41253);
or U41690 (N_41690,N_41076,N_41090);
or U41691 (N_41691,N_41109,N_41210);
or U41692 (N_41692,N_41049,N_41334);
and U41693 (N_41693,N_41250,N_41074);
nand U41694 (N_41694,N_41103,N_41422);
or U41695 (N_41695,N_41027,N_41144);
and U41696 (N_41696,N_41304,N_41496);
and U41697 (N_41697,N_41292,N_41095);
and U41698 (N_41698,N_41085,N_41189);
nand U41699 (N_41699,N_41366,N_41388);
nand U41700 (N_41700,N_41430,N_41137);
xnor U41701 (N_41701,N_41143,N_41182);
xor U41702 (N_41702,N_41410,N_41046);
and U41703 (N_41703,N_41494,N_41289);
nand U41704 (N_41704,N_41355,N_41054);
and U41705 (N_41705,N_41096,N_41124);
xor U41706 (N_41706,N_41032,N_41279);
xor U41707 (N_41707,N_41257,N_41083);
or U41708 (N_41708,N_41367,N_41263);
or U41709 (N_41709,N_41484,N_41092);
nand U41710 (N_41710,N_41127,N_41281);
nand U41711 (N_41711,N_41007,N_41225);
nand U41712 (N_41712,N_41419,N_41237);
or U41713 (N_41713,N_41141,N_41382);
or U41714 (N_41714,N_41344,N_41413);
or U41715 (N_41715,N_41108,N_41348);
and U41716 (N_41716,N_41134,N_41196);
nand U41717 (N_41717,N_41071,N_41402);
nand U41718 (N_41718,N_41048,N_41066);
or U41719 (N_41719,N_41024,N_41282);
and U41720 (N_41720,N_41280,N_41045);
and U41721 (N_41721,N_41026,N_41165);
or U41722 (N_41722,N_41411,N_41399);
xor U41723 (N_41723,N_41361,N_41133);
xor U41724 (N_41724,N_41093,N_41274);
nand U41725 (N_41725,N_41232,N_41476);
nand U41726 (N_41726,N_41466,N_41301);
nor U41727 (N_41727,N_41322,N_41167);
nor U41728 (N_41728,N_41286,N_41179);
or U41729 (N_41729,N_41031,N_41055);
nand U41730 (N_41730,N_41106,N_41033);
or U41731 (N_41731,N_41480,N_41121);
nand U41732 (N_41732,N_41151,N_41126);
nor U41733 (N_41733,N_41306,N_41228);
xor U41734 (N_41734,N_41316,N_41324);
or U41735 (N_41735,N_41240,N_41314);
or U41736 (N_41736,N_41392,N_41160);
nor U41737 (N_41737,N_41372,N_41375);
nand U41738 (N_41738,N_41396,N_41404);
nand U41739 (N_41739,N_41458,N_41087);
or U41740 (N_41740,N_41475,N_41472);
or U41741 (N_41741,N_41393,N_41187);
xor U41742 (N_41742,N_41238,N_41197);
and U41743 (N_41743,N_41409,N_41220);
nor U41744 (N_41744,N_41307,N_41295);
or U41745 (N_41745,N_41019,N_41383);
nor U41746 (N_41746,N_41122,N_41100);
or U41747 (N_41747,N_41435,N_41408);
or U41748 (N_41748,N_41153,N_41488);
or U41749 (N_41749,N_41199,N_41067);
xnor U41750 (N_41750,N_41036,N_41355);
xnor U41751 (N_41751,N_41270,N_41458);
xor U41752 (N_41752,N_41310,N_41268);
or U41753 (N_41753,N_41078,N_41360);
nand U41754 (N_41754,N_41359,N_41440);
nor U41755 (N_41755,N_41472,N_41419);
or U41756 (N_41756,N_41187,N_41301);
and U41757 (N_41757,N_41484,N_41110);
xnor U41758 (N_41758,N_41380,N_41388);
and U41759 (N_41759,N_41193,N_41229);
xnor U41760 (N_41760,N_41117,N_41389);
nand U41761 (N_41761,N_41240,N_41382);
or U41762 (N_41762,N_41301,N_41230);
nand U41763 (N_41763,N_41201,N_41299);
nand U41764 (N_41764,N_41179,N_41388);
nand U41765 (N_41765,N_41402,N_41222);
xnor U41766 (N_41766,N_41451,N_41182);
xnor U41767 (N_41767,N_41336,N_41202);
or U41768 (N_41768,N_41486,N_41407);
and U41769 (N_41769,N_41392,N_41449);
xor U41770 (N_41770,N_41278,N_41260);
nand U41771 (N_41771,N_41463,N_41441);
and U41772 (N_41772,N_41324,N_41028);
nand U41773 (N_41773,N_41053,N_41302);
and U41774 (N_41774,N_41170,N_41139);
xor U41775 (N_41775,N_41402,N_41053);
and U41776 (N_41776,N_41000,N_41196);
or U41777 (N_41777,N_41104,N_41455);
nor U41778 (N_41778,N_41163,N_41150);
xor U41779 (N_41779,N_41355,N_41126);
or U41780 (N_41780,N_41036,N_41100);
and U41781 (N_41781,N_41133,N_41083);
nand U41782 (N_41782,N_41448,N_41393);
nand U41783 (N_41783,N_41213,N_41361);
or U41784 (N_41784,N_41006,N_41065);
or U41785 (N_41785,N_41274,N_41008);
nor U41786 (N_41786,N_41254,N_41196);
or U41787 (N_41787,N_41061,N_41386);
or U41788 (N_41788,N_41059,N_41409);
nand U41789 (N_41789,N_41423,N_41103);
xnor U41790 (N_41790,N_41130,N_41308);
nand U41791 (N_41791,N_41159,N_41461);
nand U41792 (N_41792,N_41102,N_41193);
and U41793 (N_41793,N_41216,N_41128);
and U41794 (N_41794,N_41002,N_41346);
xor U41795 (N_41795,N_41224,N_41182);
nand U41796 (N_41796,N_41415,N_41347);
or U41797 (N_41797,N_41090,N_41135);
nand U41798 (N_41798,N_41341,N_41230);
and U41799 (N_41799,N_41478,N_41123);
nand U41800 (N_41800,N_41134,N_41112);
and U41801 (N_41801,N_41262,N_41063);
and U41802 (N_41802,N_41162,N_41383);
and U41803 (N_41803,N_41193,N_41200);
nor U41804 (N_41804,N_41268,N_41288);
nand U41805 (N_41805,N_41405,N_41030);
xnor U41806 (N_41806,N_41223,N_41314);
and U41807 (N_41807,N_41414,N_41276);
or U41808 (N_41808,N_41071,N_41177);
and U41809 (N_41809,N_41241,N_41424);
nor U41810 (N_41810,N_41398,N_41489);
nand U41811 (N_41811,N_41125,N_41370);
xnor U41812 (N_41812,N_41250,N_41413);
nor U41813 (N_41813,N_41469,N_41134);
or U41814 (N_41814,N_41458,N_41041);
nor U41815 (N_41815,N_41277,N_41000);
nor U41816 (N_41816,N_41061,N_41272);
or U41817 (N_41817,N_41036,N_41005);
nor U41818 (N_41818,N_41034,N_41096);
xnor U41819 (N_41819,N_41275,N_41443);
nand U41820 (N_41820,N_41327,N_41411);
and U41821 (N_41821,N_41024,N_41195);
nand U41822 (N_41822,N_41443,N_41011);
and U41823 (N_41823,N_41056,N_41203);
nor U41824 (N_41824,N_41269,N_41164);
xnor U41825 (N_41825,N_41142,N_41153);
xor U41826 (N_41826,N_41296,N_41424);
nor U41827 (N_41827,N_41491,N_41199);
nand U41828 (N_41828,N_41271,N_41495);
and U41829 (N_41829,N_41349,N_41072);
and U41830 (N_41830,N_41231,N_41254);
and U41831 (N_41831,N_41080,N_41029);
xnor U41832 (N_41832,N_41401,N_41395);
nor U41833 (N_41833,N_41106,N_41146);
nand U41834 (N_41834,N_41159,N_41303);
and U41835 (N_41835,N_41005,N_41334);
xor U41836 (N_41836,N_41198,N_41181);
and U41837 (N_41837,N_41218,N_41019);
xor U41838 (N_41838,N_41299,N_41365);
xnor U41839 (N_41839,N_41177,N_41393);
nor U41840 (N_41840,N_41140,N_41165);
xnor U41841 (N_41841,N_41445,N_41026);
nor U41842 (N_41842,N_41108,N_41325);
xor U41843 (N_41843,N_41378,N_41230);
nand U41844 (N_41844,N_41273,N_41259);
nor U41845 (N_41845,N_41360,N_41112);
nor U41846 (N_41846,N_41259,N_41204);
or U41847 (N_41847,N_41183,N_41454);
and U41848 (N_41848,N_41163,N_41155);
nand U41849 (N_41849,N_41000,N_41212);
or U41850 (N_41850,N_41241,N_41157);
and U41851 (N_41851,N_41183,N_41178);
or U41852 (N_41852,N_41248,N_41340);
and U41853 (N_41853,N_41293,N_41378);
nor U41854 (N_41854,N_41438,N_41168);
and U41855 (N_41855,N_41012,N_41296);
xor U41856 (N_41856,N_41230,N_41042);
xor U41857 (N_41857,N_41333,N_41297);
nor U41858 (N_41858,N_41060,N_41482);
or U41859 (N_41859,N_41352,N_41030);
or U41860 (N_41860,N_41297,N_41154);
xnor U41861 (N_41861,N_41285,N_41021);
nand U41862 (N_41862,N_41292,N_41094);
nor U41863 (N_41863,N_41069,N_41317);
nor U41864 (N_41864,N_41318,N_41040);
nand U41865 (N_41865,N_41167,N_41170);
xor U41866 (N_41866,N_41145,N_41410);
xor U41867 (N_41867,N_41470,N_41009);
nor U41868 (N_41868,N_41314,N_41014);
and U41869 (N_41869,N_41406,N_41052);
nand U41870 (N_41870,N_41252,N_41025);
nor U41871 (N_41871,N_41221,N_41323);
nor U41872 (N_41872,N_41449,N_41036);
or U41873 (N_41873,N_41023,N_41442);
and U41874 (N_41874,N_41039,N_41148);
nand U41875 (N_41875,N_41343,N_41476);
or U41876 (N_41876,N_41493,N_41186);
xnor U41877 (N_41877,N_41196,N_41065);
nand U41878 (N_41878,N_41278,N_41203);
and U41879 (N_41879,N_41202,N_41164);
or U41880 (N_41880,N_41185,N_41156);
xor U41881 (N_41881,N_41182,N_41210);
nor U41882 (N_41882,N_41148,N_41152);
or U41883 (N_41883,N_41019,N_41363);
xnor U41884 (N_41884,N_41381,N_41225);
nand U41885 (N_41885,N_41328,N_41415);
or U41886 (N_41886,N_41491,N_41118);
or U41887 (N_41887,N_41497,N_41122);
nor U41888 (N_41888,N_41298,N_41390);
or U41889 (N_41889,N_41480,N_41383);
nand U41890 (N_41890,N_41348,N_41189);
and U41891 (N_41891,N_41405,N_41484);
and U41892 (N_41892,N_41082,N_41442);
nand U41893 (N_41893,N_41447,N_41000);
nor U41894 (N_41894,N_41405,N_41204);
xor U41895 (N_41895,N_41001,N_41226);
nor U41896 (N_41896,N_41409,N_41088);
nand U41897 (N_41897,N_41281,N_41217);
and U41898 (N_41898,N_41315,N_41478);
and U41899 (N_41899,N_41138,N_41218);
nand U41900 (N_41900,N_41273,N_41296);
and U41901 (N_41901,N_41114,N_41158);
nor U41902 (N_41902,N_41277,N_41075);
or U41903 (N_41903,N_41345,N_41446);
nor U41904 (N_41904,N_41052,N_41021);
or U41905 (N_41905,N_41322,N_41143);
nor U41906 (N_41906,N_41392,N_41130);
and U41907 (N_41907,N_41417,N_41264);
nand U41908 (N_41908,N_41356,N_41371);
or U41909 (N_41909,N_41143,N_41111);
nor U41910 (N_41910,N_41363,N_41347);
xnor U41911 (N_41911,N_41367,N_41141);
or U41912 (N_41912,N_41191,N_41285);
nor U41913 (N_41913,N_41453,N_41408);
xnor U41914 (N_41914,N_41133,N_41136);
nor U41915 (N_41915,N_41253,N_41090);
nand U41916 (N_41916,N_41242,N_41391);
and U41917 (N_41917,N_41405,N_41060);
and U41918 (N_41918,N_41362,N_41351);
and U41919 (N_41919,N_41047,N_41483);
xor U41920 (N_41920,N_41191,N_41009);
xor U41921 (N_41921,N_41304,N_41464);
nor U41922 (N_41922,N_41130,N_41182);
nand U41923 (N_41923,N_41163,N_41459);
and U41924 (N_41924,N_41474,N_41295);
or U41925 (N_41925,N_41037,N_41324);
and U41926 (N_41926,N_41240,N_41160);
and U41927 (N_41927,N_41028,N_41236);
nor U41928 (N_41928,N_41167,N_41183);
nor U41929 (N_41929,N_41319,N_41456);
and U41930 (N_41930,N_41492,N_41090);
nand U41931 (N_41931,N_41251,N_41422);
or U41932 (N_41932,N_41487,N_41118);
or U41933 (N_41933,N_41409,N_41248);
nand U41934 (N_41934,N_41429,N_41295);
and U41935 (N_41935,N_41377,N_41496);
nor U41936 (N_41936,N_41247,N_41482);
or U41937 (N_41937,N_41388,N_41463);
and U41938 (N_41938,N_41202,N_41264);
and U41939 (N_41939,N_41322,N_41009);
or U41940 (N_41940,N_41200,N_41239);
nand U41941 (N_41941,N_41013,N_41447);
nand U41942 (N_41942,N_41482,N_41032);
or U41943 (N_41943,N_41490,N_41031);
and U41944 (N_41944,N_41287,N_41084);
or U41945 (N_41945,N_41284,N_41373);
xor U41946 (N_41946,N_41213,N_41099);
or U41947 (N_41947,N_41259,N_41354);
nor U41948 (N_41948,N_41368,N_41212);
and U41949 (N_41949,N_41357,N_41252);
and U41950 (N_41950,N_41323,N_41469);
xor U41951 (N_41951,N_41037,N_41305);
nor U41952 (N_41952,N_41146,N_41238);
xor U41953 (N_41953,N_41052,N_41221);
xor U41954 (N_41954,N_41293,N_41364);
nor U41955 (N_41955,N_41475,N_41459);
or U41956 (N_41956,N_41054,N_41091);
or U41957 (N_41957,N_41459,N_41047);
or U41958 (N_41958,N_41102,N_41012);
nor U41959 (N_41959,N_41369,N_41209);
and U41960 (N_41960,N_41185,N_41276);
nor U41961 (N_41961,N_41279,N_41429);
or U41962 (N_41962,N_41272,N_41173);
nor U41963 (N_41963,N_41018,N_41222);
xnor U41964 (N_41964,N_41225,N_41494);
nand U41965 (N_41965,N_41280,N_41096);
xnor U41966 (N_41966,N_41039,N_41059);
xnor U41967 (N_41967,N_41116,N_41126);
nor U41968 (N_41968,N_41326,N_41067);
xor U41969 (N_41969,N_41417,N_41414);
nor U41970 (N_41970,N_41099,N_41263);
nor U41971 (N_41971,N_41323,N_41225);
and U41972 (N_41972,N_41105,N_41127);
and U41973 (N_41973,N_41050,N_41468);
nand U41974 (N_41974,N_41272,N_41389);
nor U41975 (N_41975,N_41399,N_41265);
or U41976 (N_41976,N_41410,N_41328);
xnor U41977 (N_41977,N_41323,N_41183);
and U41978 (N_41978,N_41132,N_41434);
or U41979 (N_41979,N_41034,N_41451);
xnor U41980 (N_41980,N_41266,N_41017);
xor U41981 (N_41981,N_41379,N_41124);
nand U41982 (N_41982,N_41253,N_41019);
and U41983 (N_41983,N_41410,N_41383);
or U41984 (N_41984,N_41077,N_41110);
or U41985 (N_41985,N_41306,N_41486);
nor U41986 (N_41986,N_41293,N_41235);
or U41987 (N_41987,N_41135,N_41009);
and U41988 (N_41988,N_41005,N_41382);
and U41989 (N_41989,N_41172,N_41354);
and U41990 (N_41990,N_41329,N_41207);
and U41991 (N_41991,N_41000,N_41128);
or U41992 (N_41992,N_41329,N_41390);
nor U41993 (N_41993,N_41203,N_41008);
xor U41994 (N_41994,N_41010,N_41255);
nor U41995 (N_41995,N_41370,N_41378);
and U41996 (N_41996,N_41335,N_41065);
nand U41997 (N_41997,N_41304,N_41239);
or U41998 (N_41998,N_41322,N_41431);
nor U41999 (N_41999,N_41154,N_41032);
and U42000 (N_42000,N_41871,N_41722);
xnor U42001 (N_42001,N_41934,N_41796);
or U42002 (N_42002,N_41838,N_41716);
nand U42003 (N_42003,N_41884,N_41723);
nand U42004 (N_42004,N_41752,N_41683);
xnor U42005 (N_42005,N_41906,N_41867);
nor U42006 (N_42006,N_41902,N_41614);
xnor U42007 (N_42007,N_41880,N_41558);
xnor U42008 (N_42008,N_41692,N_41686);
nor U42009 (N_42009,N_41715,N_41783);
nand U42010 (N_42010,N_41938,N_41735);
xor U42011 (N_42011,N_41744,N_41963);
nor U42012 (N_42012,N_41932,N_41888);
xor U42013 (N_42013,N_41710,N_41632);
xnor U42014 (N_42014,N_41556,N_41916);
nor U42015 (N_42015,N_41584,N_41857);
or U42016 (N_42016,N_41554,N_41506);
nor U42017 (N_42017,N_41661,N_41645);
xor U42018 (N_42018,N_41758,N_41751);
xor U42019 (N_42019,N_41591,N_41619);
and U42020 (N_42020,N_41964,N_41965);
and U42021 (N_42021,N_41756,N_41733);
or U42022 (N_42022,N_41912,N_41621);
and U42023 (N_42023,N_41557,N_41680);
nor U42024 (N_42024,N_41581,N_41882);
and U42025 (N_42025,N_41775,N_41768);
nor U42026 (N_42026,N_41595,N_41507);
nand U42027 (N_42027,N_41772,N_41656);
nand U42028 (N_42028,N_41620,N_41812);
and U42029 (N_42029,N_41875,N_41674);
or U42030 (N_42030,N_41523,N_41845);
or U42031 (N_42031,N_41908,N_41839);
or U42032 (N_42032,N_41573,N_41699);
xnor U42033 (N_42033,N_41663,N_41910);
or U42034 (N_42034,N_41571,N_41760);
and U42035 (N_42035,N_41983,N_41693);
xnor U42036 (N_42036,N_41860,N_41864);
and U42037 (N_42037,N_41708,N_41815);
nor U42038 (N_42038,N_41555,N_41515);
nor U42039 (N_42039,N_41791,N_41724);
or U42040 (N_42040,N_41813,N_41535);
nor U42041 (N_42041,N_41691,N_41956);
xor U42042 (N_42042,N_41585,N_41625);
nand U42043 (N_42043,N_41905,N_41779);
xor U42044 (N_42044,N_41781,N_41930);
xor U42045 (N_42045,N_41918,N_41830);
and U42046 (N_42046,N_41915,N_41823);
or U42047 (N_42047,N_41842,N_41953);
xor U42048 (N_42048,N_41745,N_41738);
and U42049 (N_42049,N_41968,N_41970);
nand U42050 (N_42050,N_41821,N_41741);
xnor U42051 (N_42051,N_41748,N_41705);
nor U42052 (N_42052,N_41695,N_41978);
and U42053 (N_42053,N_41509,N_41911);
and U42054 (N_42054,N_41998,N_41609);
and U42055 (N_42055,N_41866,N_41924);
xor U42056 (N_42056,N_41909,N_41980);
xor U42057 (N_42057,N_41633,N_41826);
nand U42058 (N_42058,N_41634,N_41975);
and U42059 (N_42059,N_41746,N_41540);
nand U42060 (N_42060,N_41928,N_41567);
and U42061 (N_42061,N_41836,N_41954);
xor U42062 (N_42062,N_41808,N_41870);
or U42063 (N_42063,N_41536,N_41732);
nor U42064 (N_42064,N_41501,N_41827);
nor U42065 (N_42065,N_41769,N_41720);
nor U42066 (N_42066,N_41546,N_41873);
nor U42067 (N_42067,N_41858,N_41721);
nand U42068 (N_42068,N_41869,N_41767);
and U42069 (N_42069,N_41513,N_41832);
xnor U42070 (N_42070,N_41898,N_41766);
nand U42071 (N_42071,N_41936,N_41500);
or U42072 (N_42072,N_41647,N_41629);
nor U42073 (N_42073,N_41681,N_41841);
and U42074 (N_42074,N_41933,N_41712);
nor U42075 (N_42075,N_41706,N_41999);
xnor U42076 (N_42076,N_41755,N_41587);
nand U42077 (N_42077,N_41804,N_41747);
xnor U42078 (N_42078,N_41921,N_41807);
nand U42079 (N_42079,N_41658,N_41868);
nor U42080 (N_42080,N_41923,N_41895);
nor U42081 (N_42081,N_41840,N_41574);
nor U42082 (N_42082,N_41816,N_41725);
xor U42083 (N_42083,N_41763,N_41668);
nor U42084 (N_42084,N_41987,N_41613);
xnor U42085 (N_42085,N_41590,N_41577);
and U42086 (N_42086,N_41525,N_41750);
and U42087 (N_42087,N_41774,N_41865);
and U42088 (N_42088,N_41889,N_41568);
nor U42089 (N_42089,N_41800,N_41913);
or U42090 (N_42090,N_41818,N_41639);
and U42091 (N_42091,N_41597,N_41743);
and U42092 (N_42092,N_41951,N_41520);
nor U42093 (N_42093,N_41662,N_41603);
nor U42094 (N_42094,N_41992,N_41739);
or U42095 (N_42095,N_41679,N_41717);
or U42096 (N_42096,N_41967,N_41979);
and U42097 (N_42097,N_41637,N_41797);
nand U42098 (N_42098,N_41892,N_41801);
xor U42099 (N_42099,N_41569,N_41641);
or U42100 (N_42100,N_41799,N_41922);
nand U42101 (N_42101,N_41731,N_41726);
nand U42102 (N_42102,N_41599,N_41631);
xnor U42103 (N_42103,N_41885,N_41939);
xnor U42104 (N_42104,N_41605,N_41795);
xor U42105 (N_42105,N_41886,N_41958);
and U42106 (N_42106,N_41765,N_41601);
xnor U42107 (N_42107,N_41794,N_41977);
and U42108 (N_42108,N_41896,N_41891);
and U42109 (N_42109,N_41986,N_41862);
and U42110 (N_42110,N_41657,N_41698);
nor U42111 (N_42111,N_41787,N_41802);
nor U42112 (N_42112,N_41988,N_41583);
nor U42113 (N_42113,N_41907,N_41952);
and U42114 (N_42114,N_41843,N_41773);
and U42115 (N_42115,N_41685,N_41701);
nand U42116 (N_42116,N_41789,N_41949);
nor U42117 (N_42117,N_41654,N_41602);
and U42118 (N_42118,N_41829,N_41814);
xnor U42119 (N_42119,N_41596,N_41671);
nand U42120 (N_42120,N_41677,N_41655);
xnor U42121 (N_42121,N_41920,N_41516);
or U42122 (N_42122,N_41576,N_41749);
nand U42123 (N_42123,N_41904,N_41586);
and U42124 (N_42124,N_41510,N_41976);
nand U42125 (N_42125,N_41572,N_41607);
nor U42126 (N_42126,N_41973,N_41610);
nand U42127 (N_42127,N_41955,N_41694);
nand U42128 (N_42128,N_41650,N_41861);
and U42129 (N_42129,N_41901,N_41673);
nor U42130 (N_42130,N_41856,N_41618);
nor U42131 (N_42131,N_41810,N_41505);
or U42132 (N_42132,N_41853,N_41672);
and U42133 (N_42133,N_41727,N_41778);
or U42134 (N_42134,N_41788,N_41897);
nor U42135 (N_42135,N_41899,N_41944);
and U42136 (N_42136,N_41529,N_41847);
xnor U42137 (N_42137,N_41811,N_41636);
nor U42138 (N_42138,N_41990,N_41664);
or U42139 (N_42139,N_41919,N_41713);
and U42140 (N_42140,N_41817,N_41534);
xor U42141 (N_42141,N_41530,N_41640);
xnor U42142 (N_42142,N_41517,N_41642);
nand U42143 (N_42143,N_41638,N_41552);
and U42144 (N_42144,N_41564,N_41854);
xnor U42145 (N_42145,N_41687,N_41579);
and U42146 (N_42146,N_41511,N_41914);
and U42147 (N_42147,N_41690,N_41876);
nand U42148 (N_42148,N_41543,N_41524);
or U42149 (N_42149,N_41784,N_41562);
nand U42150 (N_42150,N_41890,N_41960);
nor U42151 (N_42151,N_41604,N_41643);
nand U42152 (N_42152,N_41544,N_41753);
xor U42153 (N_42153,N_41995,N_41809);
or U42154 (N_42154,N_41600,N_41945);
nand U42155 (N_42155,N_41996,N_41803);
nor U42156 (N_42156,N_41611,N_41550);
xnor U42157 (N_42157,N_41793,N_41728);
nand U42158 (N_42158,N_41833,N_41859);
nor U42159 (N_42159,N_41948,N_41874);
or U42160 (N_42160,N_41644,N_41759);
or U42161 (N_42161,N_41652,N_41545);
nor U42162 (N_42162,N_41563,N_41561);
and U42163 (N_42163,N_41659,N_41969);
or U42164 (N_42164,N_41514,N_41592);
or U42165 (N_42165,N_41792,N_41612);
or U42166 (N_42166,N_41559,N_41961);
nand U42167 (N_42167,N_41531,N_41730);
and U42168 (N_42168,N_41835,N_41831);
or U42169 (N_42169,N_41972,N_41503);
xor U42170 (N_42170,N_41627,N_41508);
and U42171 (N_42171,N_41648,N_41700);
xor U42172 (N_42172,N_41957,N_41761);
nor U42173 (N_42173,N_41593,N_41624);
and U42174 (N_42174,N_41855,N_41719);
nor U42175 (N_42175,N_41966,N_41688);
or U42176 (N_42176,N_41580,N_41740);
xnor U42177 (N_42177,N_41736,N_41900);
or U42178 (N_42178,N_41670,N_41844);
nand U42179 (N_42179,N_41849,N_41806);
nand U42180 (N_42180,N_41651,N_41626);
and U42181 (N_42181,N_41737,N_41714);
nor U42182 (N_42182,N_41927,N_41834);
nand U42183 (N_42183,N_41635,N_41893);
or U42184 (N_42184,N_41962,N_41837);
and U42185 (N_42185,N_41521,N_41606);
or U42186 (N_42186,N_41929,N_41974);
and U42187 (N_42187,N_41548,N_41863);
nor U42188 (N_42188,N_41780,N_41702);
or U42189 (N_42189,N_41819,N_41764);
and U42190 (N_42190,N_41941,N_41785);
nand U42191 (N_42191,N_41711,N_41993);
xor U42192 (N_42192,N_41532,N_41985);
xor U42193 (N_42193,N_41989,N_41649);
nor U42194 (N_42194,N_41825,N_41771);
and U42195 (N_42195,N_41786,N_41937);
and U42196 (N_42196,N_41935,N_41617);
nand U42197 (N_42197,N_41665,N_41926);
xor U42198 (N_42198,N_41528,N_41527);
and U42199 (N_42199,N_41917,N_41950);
nand U42200 (N_42200,N_41757,N_41729);
xnor U42201 (N_42201,N_41805,N_41566);
xnor U42202 (N_42202,N_41676,N_41894);
nand U42203 (N_42203,N_41946,N_41997);
or U42204 (N_42204,N_41991,N_41519);
nand U42205 (N_42205,N_41852,N_41660);
xnor U42206 (N_42206,N_41615,N_41547);
xnor U42207 (N_42207,N_41542,N_41942);
xor U42208 (N_42208,N_41850,N_41589);
and U42209 (N_42209,N_41533,N_41707);
and U42210 (N_42210,N_41943,N_41628);
nor U42211 (N_42211,N_41984,N_41947);
xor U42212 (N_42212,N_41824,N_41959);
xor U42213 (N_42213,N_41689,N_41770);
and U42214 (N_42214,N_41696,N_41678);
and U42215 (N_42215,N_41931,N_41848);
and U42216 (N_42216,N_41553,N_41704);
and U42217 (N_42217,N_41940,N_41551);
nand U42218 (N_42218,N_41878,N_41675);
and U42219 (N_42219,N_41881,N_41518);
nor U42220 (N_42220,N_41570,N_41982);
xor U42221 (N_42221,N_41653,N_41877);
xor U42222 (N_42222,N_41539,N_41820);
nor U42223 (N_42223,N_41666,N_41537);
nand U42224 (N_42224,N_41565,N_41682);
xnor U42225 (N_42225,N_41502,N_41622);
nor U42226 (N_42226,N_41549,N_41822);
xor U42227 (N_42227,N_41504,N_41887);
and U42228 (N_42228,N_41971,N_41782);
or U42229 (N_42229,N_41994,N_41594);
and U42230 (N_42230,N_41538,N_41703);
nor U42231 (N_42231,N_41762,N_41734);
xor U42232 (N_42232,N_41560,N_41646);
or U42233 (N_42233,N_41828,N_41851);
or U42234 (N_42234,N_41776,N_41630);
or U42235 (N_42235,N_41925,N_41616);
nand U42236 (N_42236,N_41754,N_41541);
nor U42237 (N_42237,N_41575,N_41522);
nor U42238 (N_42238,N_41623,N_41777);
nand U42239 (N_42239,N_41790,N_41709);
nand U42240 (N_42240,N_41582,N_41846);
xor U42241 (N_42241,N_41598,N_41697);
nor U42242 (N_42242,N_41684,N_41588);
and U42243 (N_42243,N_41512,N_41872);
nand U42244 (N_42244,N_41718,N_41578);
nand U42245 (N_42245,N_41669,N_41981);
or U42246 (N_42246,N_41742,N_41526);
and U42247 (N_42247,N_41798,N_41667);
or U42248 (N_42248,N_41608,N_41883);
or U42249 (N_42249,N_41879,N_41903);
or U42250 (N_42250,N_41546,N_41789);
or U42251 (N_42251,N_41779,N_41810);
xnor U42252 (N_42252,N_41857,N_41878);
xor U42253 (N_42253,N_41713,N_41833);
xor U42254 (N_42254,N_41949,N_41768);
nor U42255 (N_42255,N_41690,N_41608);
or U42256 (N_42256,N_41905,N_41567);
nor U42257 (N_42257,N_41537,N_41618);
nor U42258 (N_42258,N_41733,N_41557);
or U42259 (N_42259,N_41760,N_41860);
nor U42260 (N_42260,N_41594,N_41735);
nand U42261 (N_42261,N_41760,N_41639);
or U42262 (N_42262,N_41907,N_41875);
and U42263 (N_42263,N_41841,N_41514);
nor U42264 (N_42264,N_41859,N_41581);
xnor U42265 (N_42265,N_41745,N_41627);
nand U42266 (N_42266,N_41770,N_41676);
and U42267 (N_42267,N_41792,N_41836);
xnor U42268 (N_42268,N_41782,N_41750);
xnor U42269 (N_42269,N_41634,N_41810);
xnor U42270 (N_42270,N_41630,N_41999);
nor U42271 (N_42271,N_41978,N_41814);
or U42272 (N_42272,N_41925,N_41845);
nor U42273 (N_42273,N_41786,N_41614);
and U42274 (N_42274,N_41675,N_41722);
or U42275 (N_42275,N_41646,N_41955);
xor U42276 (N_42276,N_41557,N_41533);
xnor U42277 (N_42277,N_41836,N_41549);
nor U42278 (N_42278,N_41751,N_41952);
or U42279 (N_42279,N_41565,N_41533);
xor U42280 (N_42280,N_41686,N_41768);
xor U42281 (N_42281,N_41731,N_41657);
xnor U42282 (N_42282,N_41532,N_41898);
or U42283 (N_42283,N_41748,N_41592);
and U42284 (N_42284,N_41555,N_41746);
nand U42285 (N_42285,N_41547,N_41710);
or U42286 (N_42286,N_41829,N_41633);
xor U42287 (N_42287,N_41592,N_41538);
and U42288 (N_42288,N_41590,N_41982);
and U42289 (N_42289,N_41777,N_41921);
or U42290 (N_42290,N_41874,N_41674);
nor U42291 (N_42291,N_41667,N_41840);
and U42292 (N_42292,N_41558,N_41855);
and U42293 (N_42293,N_41827,N_41554);
and U42294 (N_42294,N_41813,N_41602);
and U42295 (N_42295,N_41584,N_41622);
and U42296 (N_42296,N_41598,N_41548);
nand U42297 (N_42297,N_41694,N_41701);
xor U42298 (N_42298,N_41523,N_41597);
and U42299 (N_42299,N_41966,N_41530);
or U42300 (N_42300,N_41754,N_41824);
xor U42301 (N_42301,N_41924,N_41774);
or U42302 (N_42302,N_41511,N_41976);
and U42303 (N_42303,N_41938,N_41913);
and U42304 (N_42304,N_41871,N_41814);
xor U42305 (N_42305,N_41900,N_41699);
xnor U42306 (N_42306,N_41660,N_41756);
nor U42307 (N_42307,N_41908,N_41966);
or U42308 (N_42308,N_41869,N_41596);
or U42309 (N_42309,N_41737,N_41577);
or U42310 (N_42310,N_41512,N_41765);
or U42311 (N_42311,N_41608,N_41598);
nand U42312 (N_42312,N_41953,N_41965);
or U42313 (N_42313,N_41729,N_41941);
nor U42314 (N_42314,N_41783,N_41877);
nand U42315 (N_42315,N_41804,N_41674);
xnor U42316 (N_42316,N_41979,N_41920);
or U42317 (N_42317,N_41549,N_41841);
nand U42318 (N_42318,N_41550,N_41818);
and U42319 (N_42319,N_41846,N_41965);
and U42320 (N_42320,N_41525,N_41821);
xor U42321 (N_42321,N_41784,N_41827);
nand U42322 (N_42322,N_41985,N_41853);
and U42323 (N_42323,N_41980,N_41725);
nand U42324 (N_42324,N_41675,N_41863);
xnor U42325 (N_42325,N_41800,N_41518);
or U42326 (N_42326,N_41916,N_41890);
nand U42327 (N_42327,N_41795,N_41947);
xnor U42328 (N_42328,N_41923,N_41837);
nor U42329 (N_42329,N_41513,N_41962);
and U42330 (N_42330,N_41618,N_41580);
nand U42331 (N_42331,N_41858,N_41631);
and U42332 (N_42332,N_41507,N_41533);
xnor U42333 (N_42333,N_41987,N_41965);
nor U42334 (N_42334,N_41651,N_41919);
xnor U42335 (N_42335,N_41938,N_41594);
xor U42336 (N_42336,N_41774,N_41722);
and U42337 (N_42337,N_41595,N_41917);
or U42338 (N_42338,N_41810,N_41670);
and U42339 (N_42339,N_41606,N_41501);
nor U42340 (N_42340,N_41521,N_41685);
xor U42341 (N_42341,N_41829,N_41540);
nor U42342 (N_42342,N_41876,N_41830);
nor U42343 (N_42343,N_41866,N_41842);
nand U42344 (N_42344,N_41615,N_41544);
or U42345 (N_42345,N_41514,N_41989);
and U42346 (N_42346,N_41835,N_41860);
nand U42347 (N_42347,N_41916,N_41832);
or U42348 (N_42348,N_41638,N_41816);
and U42349 (N_42349,N_41750,N_41663);
or U42350 (N_42350,N_41944,N_41925);
xnor U42351 (N_42351,N_41845,N_41753);
nor U42352 (N_42352,N_41521,N_41538);
and U42353 (N_42353,N_41609,N_41658);
and U42354 (N_42354,N_41593,N_41976);
nor U42355 (N_42355,N_41707,N_41857);
nand U42356 (N_42356,N_41830,N_41669);
and U42357 (N_42357,N_41791,N_41532);
nor U42358 (N_42358,N_41630,N_41939);
xnor U42359 (N_42359,N_41865,N_41810);
nand U42360 (N_42360,N_41650,N_41942);
and U42361 (N_42361,N_41665,N_41944);
nand U42362 (N_42362,N_41766,N_41515);
nor U42363 (N_42363,N_41665,N_41969);
nor U42364 (N_42364,N_41873,N_41939);
or U42365 (N_42365,N_41615,N_41780);
and U42366 (N_42366,N_41533,N_41505);
nor U42367 (N_42367,N_41915,N_41854);
nor U42368 (N_42368,N_41625,N_41793);
nand U42369 (N_42369,N_41715,N_41898);
nand U42370 (N_42370,N_41887,N_41834);
xnor U42371 (N_42371,N_41618,N_41862);
nor U42372 (N_42372,N_41993,N_41682);
and U42373 (N_42373,N_41899,N_41706);
nand U42374 (N_42374,N_41600,N_41830);
and U42375 (N_42375,N_41513,N_41585);
or U42376 (N_42376,N_41852,N_41539);
or U42377 (N_42377,N_41748,N_41996);
nor U42378 (N_42378,N_41564,N_41751);
nand U42379 (N_42379,N_41555,N_41952);
xnor U42380 (N_42380,N_41766,N_41658);
nand U42381 (N_42381,N_41804,N_41533);
or U42382 (N_42382,N_41903,N_41712);
and U42383 (N_42383,N_41804,N_41719);
xor U42384 (N_42384,N_41899,N_41876);
nand U42385 (N_42385,N_41911,N_41996);
xor U42386 (N_42386,N_41849,N_41762);
xor U42387 (N_42387,N_41620,N_41629);
xnor U42388 (N_42388,N_41524,N_41774);
nor U42389 (N_42389,N_41990,N_41659);
or U42390 (N_42390,N_41552,N_41621);
and U42391 (N_42391,N_41991,N_41536);
and U42392 (N_42392,N_41940,N_41531);
and U42393 (N_42393,N_41805,N_41572);
or U42394 (N_42394,N_41679,N_41561);
nor U42395 (N_42395,N_41698,N_41592);
nand U42396 (N_42396,N_41538,N_41672);
nor U42397 (N_42397,N_41744,N_41659);
or U42398 (N_42398,N_41573,N_41967);
nand U42399 (N_42399,N_41931,N_41936);
or U42400 (N_42400,N_41924,N_41918);
and U42401 (N_42401,N_41621,N_41866);
nor U42402 (N_42402,N_41780,N_41732);
xor U42403 (N_42403,N_41810,N_41878);
and U42404 (N_42404,N_41966,N_41594);
and U42405 (N_42405,N_41593,N_41978);
xor U42406 (N_42406,N_41529,N_41575);
or U42407 (N_42407,N_41931,N_41597);
or U42408 (N_42408,N_41532,N_41802);
nor U42409 (N_42409,N_41818,N_41885);
nand U42410 (N_42410,N_41517,N_41654);
nor U42411 (N_42411,N_41871,N_41777);
or U42412 (N_42412,N_41871,N_41589);
xnor U42413 (N_42413,N_41533,N_41710);
or U42414 (N_42414,N_41744,N_41829);
nor U42415 (N_42415,N_41613,N_41933);
xor U42416 (N_42416,N_41945,N_41852);
xnor U42417 (N_42417,N_41953,N_41531);
nand U42418 (N_42418,N_41993,N_41983);
or U42419 (N_42419,N_41608,N_41526);
or U42420 (N_42420,N_41920,N_41724);
and U42421 (N_42421,N_41672,N_41824);
and U42422 (N_42422,N_41853,N_41772);
and U42423 (N_42423,N_41997,N_41916);
and U42424 (N_42424,N_41576,N_41596);
nor U42425 (N_42425,N_41915,N_41768);
and U42426 (N_42426,N_41595,N_41746);
and U42427 (N_42427,N_41656,N_41578);
and U42428 (N_42428,N_41861,N_41888);
and U42429 (N_42429,N_41649,N_41524);
nand U42430 (N_42430,N_41716,N_41549);
or U42431 (N_42431,N_41574,N_41823);
and U42432 (N_42432,N_41848,N_41899);
xor U42433 (N_42433,N_41954,N_41765);
or U42434 (N_42434,N_41856,N_41502);
and U42435 (N_42435,N_41934,N_41952);
xnor U42436 (N_42436,N_41785,N_41641);
xor U42437 (N_42437,N_41885,N_41898);
nor U42438 (N_42438,N_41641,N_41561);
or U42439 (N_42439,N_41629,N_41719);
nor U42440 (N_42440,N_41517,N_41594);
xnor U42441 (N_42441,N_41930,N_41747);
or U42442 (N_42442,N_41991,N_41768);
or U42443 (N_42443,N_41835,N_41824);
xnor U42444 (N_42444,N_41903,N_41543);
or U42445 (N_42445,N_41982,N_41744);
nor U42446 (N_42446,N_41697,N_41666);
or U42447 (N_42447,N_41706,N_41613);
and U42448 (N_42448,N_41755,N_41711);
nor U42449 (N_42449,N_41753,N_41996);
nor U42450 (N_42450,N_41895,N_41594);
nand U42451 (N_42451,N_41745,N_41560);
and U42452 (N_42452,N_41621,N_41584);
xnor U42453 (N_42453,N_41799,N_41849);
nand U42454 (N_42454,N_41926,N_41616);
or U42455 (N_42455,N_41747,N_41999);
and U42456 (N_42456,N_41638,N_41662);
or U42457 (N_42457,N_41935,N_41928);
xnor U42458 (N_42458,N_41579,N_41632);
or U42459 (N_42459,N_41764,N_41506);
nor U42460 (N_42460,N_41769,N_41980);
and U42461 (N_42461,N_41688,N_41762);
xor U42462 (N_42462,N_41634,N_41788);
xnor U42463 (N_42463,N_41534,N_41891);
nand U42464 (N_42464,N_41748,N_41514);
nor U42465 (N_42465,N_41926,N_41591);
or U42466 (N_42466,N_41881,N_41884);
and U42467 (N_42467,N_41911,N_41829);
nand U42468 (N_42468,N_41595,N_41870);
nor U42469 (N_42469,N_41961,N_41577);
and U42470 (N_42470,N_41991,N_41585);
and U42471 (N_42471,N_41517,N_41593);
nand U42472 (N_42472,N_41697,N_41676);
nand U42473 (N_42473,N_41897,N_41832);
xor U42474 (N_42474,N_41808,N_41630);
nand U42475 (N_42475,N_41691,N_41611);
nand U42476 (N_42476,N_41764,N_41939);
nor U42477 (N_42477,N_41918,N_41966);
xnor U42478 (N_42478,N_41890,N_41808);
nor U42479 (N_42479,N_41750,N_41565);
or U42480 (N_42480,N_41551,N_41911);
or U42481 (N_42481,N_41826,N_41600);
or U42482 (N_42482,N_41970,N_41829);
xor U42483 (N_42483,N_41993,N_41560);
nor U42484 (N_42484,N_41634,N_41876);
nor U42485 (N_42485,N_41918,N_41601);
nand U42486 (N_42486,N_41854,N_41758);
and U42487 (N_42487,N_41566,N_41879);
xor U42488 (N_42488,N_41801,N_41677);
or U42489 (N_42489,N_41969,N_41543);
xnor U42490 (N_42490,N_41820,N_41652);
and U42491 (N_42491,N_41815,N_41840);
and U42492 (N_42492,N_41506,N_41594);
nand U42493 (N_42493,N_41644,N_41980);
nor U42494 (N_42494,N_41816,N_41813);
nor U42495 (N_42495,N_41518,N_41838);
nand U42496 (N_42496,N_41686,N_41644);
and U42497 (N_42497,N_41688,N_41950);
nor U42498 (N_42498,N_41722,N_41684);
or U42499 (N_42499,N_41604,N_41530);
and U42500 (N_42500,N_42011,N_42348);
xnor U42501 (N_42501,N_42355,N_42202);
or U42502 (N_42502,N_42057,N_42450);
nand U42503 (N_42503,N_42016,N_42052);
nand U42504 (N_42504,N_42363,N_42373);
nor U42505 (N_42505,N_42331,N_42115);
or U42506 (N_42506,N_42490,N_42127);
nand U42507 (N_42507,N_42376,N_42163);
nand U42508 (N_42508,N_42413,N_42256);
nand U42509 (N_42509,N_42224,N_42046);
xor U42510 (N_42510,N_42273,N_42103);
xor U42511 (N_42511,N_42381,N_42346);
and U42512 (N_42512,N_42310,N_42368);
nand U42513 (N_42513,N_42404,N_42002);
and U42514 (N_42514,N_42461,N_42492);
and U42515 (N_42515,N_42317,N_42491);
or U42516 (N_42516,N_42200,N_42457);
nand U42517 (N_42517,N_42184,N_42322);
nand U42518 (N_42518,N_42054,N_42214);
nand U42519 (N_42519,N_42481,N_42364);
xnor U42520 (N_42520,N_42397,N_42033);
nor U42521 (N_42521,N_42274,N_42099);
nand U42522 (N_42522,N_42291,N_42332);
and U42523 (N_42523,N_42183,N_42328);
nor U42524 (N_42524,N_42255,N_42309);
and U42525 (N_42525,N_42408,N_42107);
nor U42526 (N_42526,N_42437,N_42014);
xnor U42527 (N_42527,N_42170,N_42323);
nor U42528 (N_42528,N_42295,N_42372);
and U42529 (N_42529,N_42407,N_42341);
nor U42530 (N_42530,N_42118,N_42379);
nand U42531 (N_42531,N_42320,N_42003);
nor U42532 (N_42532,N_42210,N_42117);
nand U42533 (N_42533,N_42306,N_42292);
and U42534 (N_42534,N_42173,N_42488);
xnor U42535 (N_42535,N_42185,N_42130);
and U42536 (N_42536,N_42497,N_42037);
nand U42537 (N_42537,N_42121,N_42019);
or U42538 (N_42538,N_42122,N_42165);
and U42539 (N_42539,N_42300,N_42276);
xnor U42540 (N_42540,N_42411,N_42208);
or U42541 (N_42541,N_42010,N_42431);
or U42542 (N_42542,N_42412,N_42409);
nor U42543 (N_42543,N_42100,N_42043);
nand U42544 (N_42544,N_42063,N_42098);
or U42545 (N_42545,N_42246,N_42394);
nand U42546 (N_42546,N_42294,N_42311);
and U42547 (N_42547,N_42469,N_42489);
or U42548 (N_42548,N_42134,N_42172);
nor U42549 (N_42549,N_42056,N_42349);
xnor U42550 (N_42550,N_42433,N_42371);
nand U42551 (N_42551,N_42204,N_42125);
nand U42552 (N_42552,N_42177,N_42179);
xor U42553 (N_42553,N_42382,N_42478);
or U42554 (N_42554,N_42201,N_42499);
nand U42555 (N_42555,N_42402,N_42158);
or U42556 (N_42556,N_42329,N_42321);
or U42557 (N_42557,N_42226,N_42240);
nor U42558 (N_42558,N_42106,N_42047);
or U42559 (N_42559,N_42384,N_42076);
and U42560 (N_42560,N_42024,N_42211);
and U42561 (N_42561,N_42171,N_42314);
xor U42562 (N_42562,N_42001,N_42393);
or U42563 (N_42563,N_42479,N_42474);
xnor U42564 (N_42564,N_42388,N_42426);
or U42565 (N_42565,N_42216,N_42161);
nor U42566 (N_42566,N_42428,N_42406);
nand U42567 (N_42567,N_42187,N_42195);
nor U42568 (N_42568,N_42458,N_42167);
nor U42569 (N_42569,N_42164,N_42465);
xnor U42570 (N_42570,N_42105,N_42041);
or U42571 (N_42571,N_42302,N_42160);
or U42572 (N_42572,N_42079,N_42220);
or U42573 (N_42573,N_42059,N_42207);
nand U42574 (N_42574,N_42283,N_42451);
and U42575 (N_42575,N_42401,N_42205);
nor U42576 (N_42576,N_42385,N_42141);
or U42577 (N_42577,N_42250,N_42042);
xor U42578 (N_42578,N_42088,N_42225);
xor U42579 (N_42579,N_42000,N_42445);
and U42580 (N_42580,N_42039,N_42138);
nor U42581 (N_42581,N_42425,N_42257);
and U42582 (N_42582,N_42447,N_42070);
or U42583 (N_42583,N_42085,N_42155);
nor U42584 (N_42584,N_42441,N_42420);
and U42585 (N_42585,N_42061,N_42152);
xor U42586 (N_42586,N_42367,N_42303);
nand U42587 (N_42587,N_42045,N_42199);
nor U42588 (N_42588,N_42415,N_42254);
xnor U42589 (N_42589,N_42154,N_42053);
or U42590 (N_42590,N_42082,N_42239);
nand U42591 (N_42591,N_42149,N_42496);
and U42592 (N_42592,N_42464,N_42140);
or U42593 (N_42593,N_42071,N_42083);
nand U42594 (N_42594,N_42108,N_42077);
xnor U42595 (N_42595,N_42350,N_42110);
nand U42596 (N_42596,N_42198,N_42351);
xor U42597 (N_42597,N_42383,N_42482);
and U42598 (N_42598,N_42217,N_42233);
nor U42599 (N_42599,N_42442,N_42470);
and U42600 (N_42600,N_42288,N_42222);
nand U42601 (N_42601,N_42398,N_42290);
and U42602 (N_42602,N_42213,N_42315);
or U42603 (N_42603,N_42020,N_42008);
nand U42604 (N_42604,N_42245,N_42009);
nand U42605 (N_42605,N_42378,N_42467);
or U42606 (N_42606,N_42137,N_42060);
nor U42607 (N_42607,N_42074,N_42209);
nor U42608 (N_42608,N_42175,N_42305);
nand U42609 (N_42609,N_42416,N_42440);
or U42610 (N_42610,N_42247,N_42051);
nor U42611 (N_42611,N_42444,N_42284);
and U42612 (N_42612,N_42230,N_42090);
nand U42613 (N_42613,N_42129,N_42307);
nor U42614 (N_42614,N_42234,N_42013);
xnor U42615 (N_42615,N_42472,N_42270);
nand U42616 (N_42616,N_42073,N_42400);
or U42617 (N_42617,N_42410,N_42448);
nor U42618 (N_42618,N_42387,N_42089);
xor U42619 (N_42619,N_42271,N_42035);
or U42620 (N_42620,N_42261,N_42301);
nor U42621 (N_42621,N_42093,N_42443);
or U42622 (N_42622,N_42361,N_42162);
nor U42623 (N_42623,N_42264,N_42258);
or U42624 (N_42624,N_42174,N_42352);
or U42625 (N_42625,N_42259,N_42480);
and U42626 (N_42626,N_42072,N_42206);
xor U42627 (N_42627,N_42265,N_42025);
xor U42628 (N_42628,N_42078,N_42075);
nor U42629 (N_42629,N_42463,N_42417);
nor U42630 (N_42630,N_42181,N_42080);
nand U42631 (N_42631,N_42169,N_42267);
nand U42632 (N_42632,N_42473,N_42111);
nand U42633 (N_42633,N_42021,N_42395);
or U42634 (N_42634,N_42278,N_42439);
or U42635 (N_42635,N_42068,N_42485);
or U42636 (N_42636,N_42414,N_42342);
xnor U42637 (N_42637,N_42203,N_42150);
or U42638 (N_42638,N_42453,N_42285);
xnor U42639 (N_42639,N_42369,N_42116);
and U42640 (N_42640,N_42251,N_42244);
xor U42641 (N_42641,N_42452,N_42124);
and U42642 (N_42642,N_42197,N_42109);
and U42643 (N_42643,N_42036,N_42142);
or U42644 (N_42644,N_42475,N_42038);
nand U42645 (N_42645,N_42242,N_42194);
xor U42646 (N_42646,N_42260,N_42374);
nand U42647 (N_42647,N_42102,N_42293);
and U42648 (N_42648,N_42015,N_42026);
nor U42649 (N_42649,N_42392,N_42421);
and U42650 (N_42650,N_42396,N_42316);
nand U42651 (N_42651,N_42133,N_42139);
nand U42652 (N_42652,N_42029,N_42159);
nor U42653 (N_42653,N_42252,N_42324);
and U42654 (N_42654,N_42178,N_42229);
nor U42655 (N_42655,N_42028,N_42438);
nand U42656 (N_42656,N_42048,N_42196);
xnor U42657 (N_42657,N_42299,N_42319);
nand U42658 (N_42658,N_42269,N_42403);
xor U42659 (N_42659,N_42120,N_42494);
nand U42660 (N_42660,N_42434,N_42031);
nand U42661 (N_42661,N_42455,N_42272);
nor U42662 (N_42662,N_42389,N_42238);
nand U42663 (N_42663,N_42219,N_42241);
nor U42664 (N_42664,N_42237,N_42215);
or U42665 (N_42665,N_42065,N_42468);
or U42666 (N_42666,N_42281,N_42062);
nor U42667 (N_42667,N_42227,N_42484);
nor U42668 (N_42668,N_42427,N_42104);
xor U42669 (N_42669,N_42432,N_42218);
xor U42670 (N_42670,N_42466,N_42249);
nand U42671 (N_42671,N_42146,N_42081);
xor U42672 (N_42672,N_42044,N_42498);
nand U42673 (N_42673,N_42326,N_42359);
and U42674 (N_42674,N_42232,N_42193);
xor U42675 (N_42675,N_42362,N_42212);
nand U42676 (N_42676,N_42275,N_42476);
or U42677 (N_42677,N_42405,N_42049);
nor U42678 (N_42678,N_42188,N_42144);
nand U42679 (N_42679,N_42423,N_42424);
nand U42680 (N_42680,N_42248,N_42366);
xnor U42681 (N_42681,N_42135,N_42223);
and U42682 (N_42682,N_42279,N_42231);
xor U42683 (N_42683,N_42262,N_42131);
nor U42684 (N_42684,N_42114,N_42006);
or U42685 (N_42685,N_42454,N_42330);
and U42686 (N_42686,N_42487,N_42228);
xor U42687 (N_42687,N_42221,N_42112);
xor U42688 (N_42688,N_42486,N_42012);
xor U42689 (N_42689,N_42034,N_42449);
or U42690 (N_42690,N_42493,N_42477);
and U42691 (N_42691,N_42338,N_42189);
or U42692 (N_42692,N_42148,N_42253);
or U42693 (N_42693,N_42176,N_42166);
or U42694 (N_42694,N_42132,N_42419);
and U42695 (N_42695,N_42343,N_42282);
xnor U42696 (N_42696,N_42312,N_42168);
nand U42697 (N_42697,N_42086,N_42182);
xor U42698 (N_42698,N_42483,N_42429);
and U42699 (N_42699,N_42180,N_42345);
or U42700 (N_42700,N_42356,N_42298);
nor U42701 (N_42701,N_42143,N_42296);
nand U42702 (N_42702,N_42235,N_42391);
nor U42703 (N_42703,N_42087,N_42005);
nand U42704 (N_42704,N_42084,N_42308);
or U42705 (N_42705,N_42456,N_42377);
xor U42706 (N_42706,N_42418,N_42095);
nand U42707 (N_42707,N_42268,N_42340);
and U42708 (N_42708,N_42436,N_42058);
nor U42709 (N_42709,N_42286,N_42091);
or U42710 (N_42710,N_42030,N_42069);
nand U42711 (N_42711,N_42337,N_42101);
xor U42712 (N_42712,N_42018,N_42151);
nand U42713 (N_42713,N_42066,N_42017);
nand U42714 (N_42714,N_42190,N_42399);
nor U42715 (N_42715,N_42459,N_42094);
or U42716 (N_42716,N_42263,N_42067);
nand U42717 (N_42717,N_42236,N_42333);
nand U42718 (N_42718,N_42123,N_42147);
or U42719 (N_42719,N_42096,N_42313);
nand U42720 (N_42720,N_42347,N_42430);
or U42721 (N_42721,N_42092,N_42097);
or U42722 (N_42722,N_42446,N_42023);
nand U42723 (N_42723,N_42336,N_42339);
nor U42724 (N_42724,N_42318,N_42357);
and U42725 (N_42725,N_42344,N_42050);
nand U42726 (N_42726,N_42040,N_42435);
and U42727 (N_42727,N_42128,N_42353);
xor U42728 (N_42728,N_42287,N_42460);
nor U42729 (N_42729,N_42304,N_42280);
or U42730 (N_42730,N_42266,N_42334);
nor U42731 (N_42731,N_42145,N_42422);
and U42732 (N_42732,N_42022,N_42354);
and U42733 (N_42733,N_42365,N_42156);
nor U42734 (N_42734,N_42358,N_42375);
and U42735 (N_42735,N_42386,N_42471);
or U42736 (N_42736,N_42126,N_42157);
nand U42737 (N_42737,N_42495,N_42004);
nor U42738 (N_42738,N_42119,N_42064);
nand U42739 (N_42739,N_42153,N_42192);
or U42740 (N_42740,N_42277,N_42360);
xnor U42741 (N_42741,N_42370,N_42186);
nor U42742 (N_42742,N_42055,N_42289);
or U42743 (N_42743,N_42032,N_42007);
nor U42744 (N_42744,N_42297,N_42325);
nand U42745 (N_42745,N_42390,N_42027);
nor U42746 (N_42746,N_42191,N_42335);
or U42747 (N_42747,N_42327,N_42380);
nor U42748 (N_42748,N_42462,N_42113);
xor U42749 (N_42749,N_42243,N_42136);
or U42750 (N_42750,N_42386,N_42179);
or U42751 (N_42751,N_42178,N_42396);
and U42752 (N_42752,N_42493,N_42079);
and U42753 (N_42753,N_42111,N_42365);
xnor U42754 (N_42754,N_42430,N_42004);
and U42755 (N_42755,N_42158,N_42345);
xor U42756 (N_42756,N_42423,N_42324);
and U42757 (N_42757,N_42007,N_42128);
nor U42758 (N_42758,N_42163,N_42455);
nor U42759 (N_42759,N_42188,N_42089);
nand U42760 (N_42760,N_42146,N_42358);
or U42761 (N_42761,N_42429,N_42039);
and U42762 (N_42762,N_42396,N_42121);
nand U42763 (N_42763,N_42116,N_42389);
and U42764 (N_42764,N_42067,N_42167);
nand U42765 (N_42765,N_42472,N_42025);
nor U42766 (N_42766,N_42393,N_42307);
nand U42767 (N_42767,N_42193,N_42475);
nand U42768 (N_42768,N_42426,N_42488);
or U42769 (N_42769,N_42247,N_42336);
or U42770 (N_42770,N_42090,N_42295);
xor U42771 (N_42771,N_42109,N_42045);
nor U42772 (N_42772,N_42248,N_42386);
or U42773 (N_42773,N_42462,N_42112);
and U42774 (N_42774,N_42323,N_42465);
nand U42775 (N_42775,N_42083,N_42441);
nor U42776 (N_42776,N_42072,N_42427);
xnor U42777 (N_42777,N_42304,N_42177);
or U42778 (N_42778,N_42491,N_42386);
nor U42779 (N_42779,N_42146,N_42258);
and U42780 (N_42780,N_42139,N_42288);
nand U42781 (N_42781,N_42042,N_42475);
xor U42782 (N_42782,N_42329,N_42180);
nand U42783 (N_42783,N_42432,N_42477);
nand U42784 (N_42784,N_42184,N_42374);
or U42785 (N_42785,N_42393,N_42058);
and U42786 (N_42786,N_42373,N_42297);
nand U42787 (N_42787,N_42440,N_42001);
xnor U42788 (N_42788,N_42311,N_42121);
nand U42789 (N_42789,N_42469,N_42187);
nand U42790 (N_42790,N_42272,N_42202);
or U42791 (N_42791,N_42131,N_42060);
xnor U42792 (N_42792,N_42228,N_42371);
xnor U42793 (N_42793,N_42469,N_42041);
nor U42794 (N_42794,N_42254,N_42002);
or U42795 (N_42795,N_42055,N_42059);
or U42796 (N_42796,N_42463,N_42480);
xnor U42797 (N_42797,N_42380,N_42195);
and U42798 (N_42798,N_42432,N_42245);
and U42799 (N_42799,N_42260,N_42070);
xor U42800 (N_42800,N_42056,N_42418);
nor U42801 (N_42801,N_42211,N_42360);
nand U42802 (N_42802,N_42262,N_42399);
xor U42803 (N_42803,N_42316,N_42259);
or U42804 (N_42804,N_42390,N_42103);
and U42805 (N_42805,N_42183,N_42198);
or U42806 (N_42806,N_42027,N_42034);
and U42807 (N_42807,N_42015,N_42242);
nor U42808 (N_42808,N_42138,N_42286);
nor U42809 (N_42809,N_42184,N_42271);
and U42810 (N_42810,N_42120,N_42254);
xnor U42811 (N_42811,N_42454,N_42051);
or U42812 (N_42812,N_42372,N_42247);
nand U42813 (N_42813,N_42175,N_42323);
nor U42814 (N_42814,N_42446,N_42006);
and U42815 (N_42815,N_42234,N_42480);
xor U42816 (N_42816,N_42131,N_42480);
nand U42817 (N_42817,N_42143,N_42439);
nand U42818 (N_42818,N_42107,N_42332);
and U42819 (N_42819,N_42346,N_42283);
xnor U42820 (N_42820,N_42067,N_42463);
or U42821 (N_42821,N_42387,N_42099);
nand U42822 (N_42822,N_42038,N_42160);
or U42823 (N_42823,N_42163,N_42329);
and U42824 (N_42824,N_42378,N_42368);
nand U42825 (N_42825,N_42080,N_42188);
or U42826 (N_42826,N_42377,N_42110);
xnor U42827 (N_42827,N_42073,N_42337);
xnor U42828 (N_42828,N_42037,N_42485);
nor U42829 (N_42829,N_42249,N_42364);
nor U42830 (N_42830,N_42320,N_42479);
and U42831 (N_42831,N_42050,N_42180);
nor U42832 (N_42832,N_42164,N_42441);
xnor U42833 (N_42833,N_42118,N_42025);
xor U42834 (N_42834,N_42042,N_42344);
and U42835 (N_42835,N_42044,N_42397);
xor U42836 (N_42836,N_42200,N_42021);
xor U42837 (N_42837,N_42268,N_42070);
nor U42838 (N_42838,N_42107,N_42090);
xor U42839 (N_42839,N_42167,N_42134);
or U42840 (N_42840,N_42382,N_42197);
xnor U42841 (N_42841,N_42030,N_42335);
and U42842 (N_42842,N_42025,N_42280);
nor U42843 (N_42843,N_42181,N_42414);
nor U42844 (N_42844,N_42243,N_42261);
and U42845 (N_42845,N_42170,N_42166);
nor U42846 (N_42846,N_42197,N_42136);
nand U42847 (N_42847,N_42406,N_42058);
nand U42848 (N_42848,N_42161,N_42230);
nand U42849 (N_42849,N_42072,N_42212);
or U42850 (N_42850,N_42160,N_42061);
and U42851 (N_42851,N_42322,N_42176);
and U42852 (N_42852,N_42279,N_42188);
xnor U42853 (N_42853,N_42015,N_42381);
nor U42854 (N_42854,N_42015,N_42002);
nand U42855 (N_42855,N_42414,N_42431);
or U42856 (N_42856,N_42370,N_42306);
xnor U42857 (N_42857,N_42164,N_42351);
or U42858 (N_42858,N_42461,N_42103);
nand U42859 (N_42859,N_42140,N_42344);
and U42860 (N_42860,N_42417,N_42194);
and U42861 (N_42861,N_42445,N_42312);
nand U42862 (N_42862,N_42387,N_42493);
or U42863 (N_42863,N_42420,N_42055);
nand U42864 (N_42864,N_42194,N_42372);
nand U42865 (N_42865,N_42416,N_42081);
nor U42866 (N_42866,N_42333,N_42346);
nor U42867 (N_42867,N_42274,N_42211);
and U42868 (N_42868,N_42024,N_42049);
nor U42869 (N_42869,N_42402,N_42183);
nand U42870 (N_42870,N_42464,N_42188);
nor U42871 (N_42871,N_42482,N_42431);
nor U42872 (N_42872,N_42280,N_42202);
nand U42873 (N_42873,N_42091,N_42485);
xnor U42874 (N_42874,N_42267,N_42133);
nand U42875 (N_42875,N_42493,N_42354);
nand U42876 (N_42876,N_42365,N_42213);
xnor U42877 (N_42877,N_42160,N_42106);
or U42878 (N_42878,N_42138,N_42449);
or U42879 (N_42879,N_42208,N_42444);
nand U42880 (N_42880,N_42035,N_42413);
and U42881 (N_42881,N_42138,N_42323);
nand U42882 (N_42882,N_42228,N_42322);
nand U42883 (N_42883,N_42249,N_42167);
xnor U42884 (N_42884,N_42207,N_42184);
and U42885 (N_42885,N_42112,N_42132);
nand U42886 (N_42886,N_42001,N_42196);
or U42887 (N_42887,N_42479,N_42089);
nor U42888 (N_42888,N_42053,N_42094);
and U42889 (N_42889,N_42317,N_42333);
nor U42890 (N_42890,N_42100,N_42482);
nand U42891 (N_42891,N_42075,N_42446);
xor U42892 (N_42892,N_42344,N_42456);
xor U42893 (N_42893,N_42268,N_42381);
xnor U42894 (N_42894,N_42209,N_42330);
nor U42895 (N_42895,N_42444,N_42423);
xor U42896 (N_42896,N_42050,N_42098);
nor U42897 (N_42897,N_42489,N_42121);
and U42898 (N_42898,N_42472,N_42265);
nor U42899 (N_42899,N_42141,N_42058);
xnor U42900 (N_42900,N_42280,N_42355);
xnor U42901 (N_42901,N_42435,N_42423);
or U42902 (N_42902,N_42180,N_42402);
or U42903 (N_42903,N_42319,N_42324);
xor U42904 (N_42904,N_42214,N_42456);
nand U42905 (N_42905,N_42122,N_42384);
nor U42906 (N_42906,N_42380,N_42187);
or U42907 (N_42907,N_42040,N_42004);
xor U42908 (N_42908,N_42065,N_42103);
and U42909 (N_42909,N_42134,N_42069);
nor U42910 (N_42910,N_42112,N_42142);
nor U42911 (N_42911,N_42031,N_42250);
and U42912 (N_42912,N_42089,N_42019);
xor U42913 (N_42913,N_42334,N_42268);
or U42914 (N_42914,N_42377,N_42249);
nand U42915 (N_42915,N_42244,N_42416);
nand U42916 (N_42916,N_42315,N_42177);
or U42917 (N_42917,N_42449,N_42391);
xor U42918 (N_42918,N_42122,N_42367);
xor U42919 (N_42919,N_42244,N_42271);
or U42920 (N_42920,N_42480,N_42300);
or U42921 (N_42921,N_42285,N_42006);
xnor U42922 (N_42922,N_42127,N_42265);
and U42923 (N_42923,N_42139,N_42430);
and U42924 (N_42924,N_42052,N_42324);
nand U42925 (N_42925,N_42090,N_42478);
or U42926 (N_42926,N_42055,N_42355);
nand U42927 (N_42927,N_42091,N_42079);
xnor U42928 (N_42928,N_42084,N_42461);
and U42929 (N_42929,N_42116,N_42027);
or U42930 (N_42930,N_42389,N_42077);
xnor U42931 (N_42931,N_42257,N_42200);
or U42932 (N_42932,N_42145,N_42434);
and U42933 (N_42933,N_42021,N_42031);
or U42934 (N_42934,N_42138,N_42203);
or U42935 (N_42935,N_42118,N_42076);
nand U42936 (N_42936,N_42434,N_42243);
or U42937 (N_42937,N_42414,N_42307);
nor U42938 (N_42938,N_42228,N_42288);
or U42939 (N_42939,N_42303,N_42259);
xnor U42940 (N_42940,N_42123,N_42317);
nor U42941 (N_42941,N_42136,N_42443);
nand U42942 (N_42942,N_42064,N_42152);
nand U42943 (N_42943,N_42000,N_42297);
or U42944 (N_42944,N_42178,N_42068);
nor U42945 (N_42945,N_42087,N_42212);
nand U42946 (N_42946,N_42374,N_42288);
nand U42947 (N_42947,N_42133,N_42425);
nand U42948 (N_42948,N_42077,N_42458);
and U42949 (N_42949,N_42065,N_42173);
xnor U42950 (N_42950,N_42037,N_42435);
and U42951 (N_42951,N_42231,N_42263);
nor U42952 (N_42952,N_42453,N_42309);
and U42953 (N_42953,N_42035,N_42112);
nand U42954 (N_42954,N_42410,N_42204);
nand U42955 (N_42955,N_42247,N_42187);
nor U42956 (N_42956,N_42350,N_42384);
or U42957 (N_42957,N_42303,N_42403);
and U42958 (N_42958,N_42154,N_42237);
and U42959 (N_42959,N_42231,N_42227);
nor U42960 (N_42960,N_42210,N_42192);
nor U42961 (N_42961,N_42362,N_42030);
or U42962 (N_42962,N_42295,N_42193);
and U42963 (N_42963,N_42147,N_42090);
or U42964 (N_42964,N_42181,N_42030);
nor U42965 (N_42965,N_42181,N_42067);
nand U42966 (N_42966,N_42440,N_42167);
or U42967 (N_42967,N_42116,N_42200);
and U42968 (N_42968,N_42220,N_42206);
nor U42969 (N_42969,N_42331,N_42391);
nand U42970 (N_42970,N_42349,N_42401);
xnor U42971 (N_42971,N_42188,N_42181);
nor U42972 (N_42972,N_42493,N_42166);
xnor U42973 (N_42973,N_42387,N_42432);
or U42974 (N_42974,N_42104,N_42053);
and U42975 (N_42975,N_42121,N_42197);
or U42976 (N_42976,N_42020,N_42133);
or U42977 (N_42977,N_42453,N_42361);
and U42978 (N_42978,N_42247,N_42285);
xor U42979 (N_42979,N_42173,N_42019);
and U42980 (N_42980,N_42002,N_42188);
xnor U42981 (N_42981,N_42474,N_42125);
and U42982 (N_42982,N_42187,N_42412);
nor U42983 (N_42983,N_42272,N_42142);
xor U42984 (N_42984,N_42441,N_42198);
nor U42985 (N_42985,N_42457,N_42356);
or U42986 (N_42986,N_42184,N_42439);
and U42987 (N_42987,N_42172,N_42484);
nand U42988 (N_42988,N_42034,N_42120);
nor U42989 (N_42989,N_42041,N_42121);
and U42990 (N_42990,N_42339,N_42265);
nand U42991 (N_42991,N_42475,N_42117);
nand U42992 (N_42992,N_42148,N_42112);
nor U42993 (N_42993,N_42025,N_42222);
or U42994 (N_42994,N_42075,N_42415);
and U42995 (N_42995,N_42092,N_42318);
nor U42996 (N_42996,N_42257,N_42272);
nand U42997 (N_42997,N_42263,N_42265);
nand U42998 (N_42998,N_42095,N_42227);
nand U42999 (N_42999,N_42209,N_42438);
xnor U43000 (N_43000,N_42649,N_42787);
nor U43001 (N_43001,N_42611,N_42652);
or U43002 (N_43002,N_42731,N_42749);
and U43003 (N_43003,N_42552,N_42730);
nor U43004 (N_43004,N_42514,N_42501);
xor U43005 (N_43005,N_42642,N_42719);
nand U43006 (N_43006,N_42534,N_42567);
nand U43007 (N_43007,N_42860,N_42743);
and U43008 (N_43008,N_42639,N_42871);
nor U43009 (N_43009,N_42788,N_42765);
xnor U43010 (N_43010,N_42894,N_42671);
or U43011 (N_43011,N_42928,N_42689);
or U43012 (N_43012,N_42880,N_42595);
nor U43013 (N_43013,N_42720,N_42794);
nand U43014 (N_43014,N_42829,N_42902);
xor U43015 (N_43015,N_42695,N_42525);
nand U43016 (N_43016,N_42839,N_42596);
or U43017 (N_43017,N_42949,N_42738);
and U43018 (N_43018,N_42570,N_42760);
nor U43019 (N_43019,N_42887,N_42737);
nand U43020 (N_43020,N_42536,N_42670);
or U43021 (N_43021,N_42950,N_42589);
nor U43022 (N_43022,N_42755,N_42547);
xor U43023 (N_43023,N_42965,N_42597);
nor U43024 (N_43024,N_42840,N_42980);
and U43025 (N_43025,N_42548,N_42684);
or U43026 (N_43026,N_42989,N_42783);
nor U43027 (N_43027,N_42687,N_42975);
xor U43028 (N_43028,N_42680,N_42962);
and U43029 (N_43029,N_42541,N_42591);
xor U43030 (N_43030,N_42568,N_42544);
nand U43031 (N_43031,N_42672,N_42726);
nor U43032 (N_43032,N_42919,N_42833);
xnor U43033 (N_43033,N_42700,N_42575);
and U43034 (N_43034,N_42763,N_42886);
nand U43035 (N_43035,N_42982,N_42948);
nand U43036 (N_43036,N_42777,N_42706);
nor U43037 (N_43037,N_42942,N_42822);
and U43038 (N_43038,N_42924,N_42615);
or U43039 (N_43039,N_42890,N_42842);
nor U43040 (N_43040,N_42657,N_42914);
and U43041 (N_43041,N_42558,N_42804);
nor U43042 (N_43042,N_42869,N_42861);
nand U43043 (N_43043,N_42746,N_42981);
and U43044 (N_43044,N_42898,N_42513);
nand U43045 (N_43045,N_42766,N_42576);
nor U43046 (N_43046,N_42864,N_42773);
xnor U43047 (N_43047,N_42813,N_42709);
nand U43048 (N_43048,N_42958,N_42872);
and U43049 (N_43049,N_42688,N_42978);
nor U43050 (N_43050,N_42632,N_42844);
and U43051 (N_43051,N_42908,N_42776);
and U43052 (N_43052,N_42791,N_42650);
nor U43053 (N_43053,N_42578,N_42505);
nor U43054 (N_43054,N_42526,N_42723);
and U43055 (N_43055,N_42991,N_42518);
and U43056 (N_43056,N_42845,N_42754);
and U43057 (N_43057,N_42748,N_42555);
nand U43058 (N_43058,N_42973,N_42549);
nand U43059 (N_43059,N_42584,N_42952);
xor U43060 (N_43060,N_42905,N_42533);
or U43061 (N_43061,N_42951,N_42992);
nand U43062 (N_43062,N_42874,N_42917);
nor U43063 (N_43063,N_42884,N_42599);
xor U43064 (N_43064,N_42590,N_42588);
nor U43065 (N_43065,N_42583,N_42511);
and U43066 (N_43066,N_42853,N_42532);
nand U43067 (N_43067,N_42598,N_42769);
and U43068 (N_43068,N_42888,N_42560);
nand U43069 (N_43069,N_42970,N_42551);
or U43070 (N_43070,N_42664,N_42637);
xor U43071 (N_43071,N_42734,N_42616);
or U43072 (N_43072,N_42816,N_42814);
and U43073 (N_43073,N_42745,N_42733);
or U43074 (N_43074,N_42711,N_42721);
xnor U43075 (N_43075,N_42638,N_42566);
xor U43076 (N_43076,N_42770,N_42802);
xor U43077 (N_43077,N_42866,N_42622);
xnor U43078 (N_43078,N_42955,N_42781);
or U43079 (N_43079,N_42739,N_42660);
and U43080 (N_43080,N_42640,N_42883);
nand U43081 (N_43081,N_42586,N_42907);
nand U43082 (N_43082,N_42796,N_42805);
nand U43083 (N_43083,N_42520,N_42574);
nor U43084 (N_43084,N_42841,N_42858);
and U43085 (N_43085,N_42939,N_42658);
xnor U43086 (N_43086,N_42545,N_42524);
nor U43087 (N_43087,N_42512,N_42944);
nand U43088 (N_43088,N_42850,N_42529);
xnor U43089 (N_43089,N_42608,N_42537);
xor U43090 (N_43090,N_42885,N_42550);
nor U43091 (N_43091,N_42676,N_42740);
or U43092 (N_43092,N_42943,N_42699);
nand U43093 (N_43093,N_42984,N_42810);
or U43094 (N_43094,N_42929,N_42798);
and U43095 (N_43095,N_42865,N_42517);
or U43096 (N_43096,N_42820,N_42722);
nor U43097 (N_43097,N_42610,N_42582);
nand U43098 (N_43098,N_42623,N_42508);
xor U43099 (N_43099,N_42702,N_42990);
nor U43100 (N_43100,N_42707,N_42602);
nand U43101 (N_43101,N_42785,N_42831);
nand U43102 (N_43102,N_42579,N_42969);
or U43103 (N_43103,N_42636,N_42521);
or U43104 (N_43104,N_42717,N_42971);
nand U43105 (N_43105,N_42895,N_42784);
nand U43106 (N_43106,N_42921,N_42922);
nand U43107 (N_43107,N_42607,N_42979);
xor U43108 (N_43108,N_42806,N_42750);
nor U43109 (N_43109,N_42605,N_42609);
and U43110 (N_43110,N_42851,N_42528);
and U43111 (N_43111,N_42799,N_42875);
and U43112 (N_43112,N_42643,N_42698);
and U43113 (N_43113,N_42729,N_42500);
xnor U43114 (N_43114,N_42911,N_42564);
nor U43115 (N_43115,N_42916,N_42556);
xor U43116 (N_43116,N_42627,N_42857);
and U43117 (N_43117,N_42974,N_42826);
and U43118 (N_43118,N_42604,N_42697);
and U43119 (N_43119,N_42661,N_42538);
and U43120 (N_43120,N_42535,N_42696);
or U43121 (N_43121,N_42987,N_42577);
xnor U43122 (N_43122,N_42912,N_42811);
or U43123 (N_43123,N_42998,N_42782);
xor U43124 (N_43124,N_42600,N_42543);
or U43125 (N_43125,N_42893,N_42531);
nand U43126 (N_43126,N_42587,N_42855);
nand U43127 (N_43127,N_42747,N_42995);
or U43128 (N_43128,N_42808,N_42554);
and U43129 (N_43129,N_42830,N_42562);
xnor U43130 (N_43130,N_42847,N_42879);
or U43131 (N_43131,N_42758,N_42704);
and U43132 (N_43132,N_42827,N_42527);
nand U43133 (N_43133,N_42712,N_42986);
nor U43134 (N_43134,N_42504,N_42581);
nand U43135 (N_43135,N_42735,N_42935);
xnor U43136 (N_43136,N_42646,N_42593);
and U43137 (N_43137,N_42626,N_42753);
or U43138 (N_43138,N_42631,N_42867);
xnor U43139 (N_43139,N_42956,N_42635);
nand U43140 (N_43140,N_42561,N_42876);
or U43141 (N_43141,N_42759,N_42679);
nand U43142 (N_43142,N_42546,N_42507);
and U43143 (N_43143,N_42832,N_42852);
nand U43144 (N_43144,N_42823,N_42837);
nand U43145 (N_43145,N_42778,N_42931);
and U43146 (N_43146,N_42667,N_42834);
nor U43147 (N_43147,N_42644,N_42983);
or U43148 (N_43148,N_42812,N_42946);
and U43149 (N_43149,N_42892,N_42889);
and U43150 (N_43150,N_42937,N_42896);
and U43151 (N_43151,N_42906,N_42648);
and U43152 (N_43152,N_42515,N_42630);
nand U43153 (N_43153,N_42647,N_42620);
or U43154 (N_43154,N_42523,N_42977);
xor U43155 (N_43155,N_42761,N_42961);
nor U43156 (N_43156,N_42553,N_42678);
nand U43157 (N_43157,N_42900,N_42792);
xor U43158 (N_43158,N_42903,N_42817);
and U43159 (N_43159,N_42828,N_42849);
nand U43160 (N_43160,N_42800,N_42881);
nand U43161 (N_43161,N_42868,N_42913);
and U43162 (N_43162,N_42621,N_42742);
nor U43163 (N_43163,N_42634,N_42613);
or U43164 (N_43164,N_42877,N_42617);
xnor U43165 (N_43165,N_42542,N_42744);
nand U43166 (N_43166,N_42601,N_42669);
or U43167 (N_43167,N_42838,N_42918);
nand U43168 (N_43168,N_42927,N_42503);
or U43169 (N_43169,N_42933,N_42563);
xnor U43170 (N_43170,N_42502,N_42967);
and U43171 (N_43171,N_42854,N_42795);
nand U43172 (N_43172,N_42999,N_42651);
xnor U43173 (N_43173,N_42665,N_42752);
xnor U43174 (N_43174,N_42771,N_42509);
and U43175 (N_43175,N_42594,N_42681);
and U43176 (N_43176,N_42920,N_42663);
nor U43177 (N_43177,N_42904,N_42682);
nor U43178 (N_43178,N_42775,N_42724);
nor U43179 (N_43179,N_42690,N_42653);
nand U43180 (N_43180,N_42940,N_42848);
or U43181 (N_43181,N_42945,N_42993);
nor U43182 (N_43182,N_42994,N_42633);
xor U43183 (N_43183,N_42963,N_42655);
and U43184 (N_43184,N_42862,N_42668);
and U43185 (N_43185,N_42941,N_42519);
nand U43186 (N_43186,N_42694,N_42686);
xor U43187 (N_43187,N_42809,N_42934);
or U43188 (N_43188,N_42736,N_42856);
or U43189 (N_43189,N_42530,N_42727);
or U43190 (N_43190,N_42891,N_42824);
nor U43191 (N_43191,N_42930,N_42996);
xor U43192 (N_43192,N_42619,N_42815);
nand U43193 (N_43193,N_42539,N_42618);
xor U43194 (N_43194,N_42715,N_42751);
or U43195 (N_43195,N_42585,N_42522);
nor U43196 (N_43196,N_42843,N_42899);
or U43197 (N_43197,N_42966,N_42797);
or U43198 (N_43198,N_42859,N_42572);
xnor U43199 (N_43199,N_42835,N_42959);
nor U43200 (N_43200,N_42625,N_42685);
xnor U43201 (N_43201,N_42882,N_42540);
nor U43202 (N_43202,N_42953,N_42628);
nor U43203 (N_43203,N_42947,N_42968);
or U43204 (N_43204,N_42654,N_42878);
or U43205 (N_43205,N_42801,N_42819);
xnor U43206 (N_43206,N_42870,N_42677);
xnor U43207 (N_43207,N_42786,N_42645);
or U43208 (N_43208,N_42675,N_42789);
and U43209 (N_43209,N_42938,N_42580);
xor U43210 (N_43210,N_42708,N_42662);
nor U43211 (N_43211,N_42846,N_42674);
nand U43212 (N_43212,N_42923,N_42756);
nand U43213 (N_43213,N_42932,N_42692);
nand U43214 (N_43214,N_42836,N_42954);
and U43215 (N_43215,N_42897,N_42997);
or U43216 (N_43216,N_42780,N_42612);
or U43217 (N_43217,N_42767,N_42516);
nor U43218 (N_43218,N_42741,N_42772);
or U43219 (N_43219,N_42779,N_42926);
or U43220 (N_43220,N_42510,N_42614);
or U43221 (N_43221,N_42818,N_42703);
xor U43222 (N_43222,N_42603,N_42762);
xnor U43223 (N_43223,N_42757,N_42807);
xor U43224 (N_43224,N_42764,N_42659);
and U43225 (N_43225,N_42960,N_42557);
nor U43226 (N_43226,N_42988,N_42569);
nor U43227 (N_43227,N_42683,N_42673);
nor U43228 (N_43228,N_42691,N_42606);
or U43229 (N_43229,N_42873,N_42985);
or U43230 (N_43230,N_42915,N_42863);
and U43231 (N_43231,N_42728,N_42825);
and U43232 (N_43232,N_42774,N_42790);
nor U43233 (N_43233,N_42565,N_42693);
or U43234 (N_43234,N_42821,N_42701);
xnor U43235 (N_43235,N_42768,N_42714);
and U43236 (N_43236,N_42716,N_42624);
and U43237 (N_43237,N_42936,N_42718);
or U43238 (N_43238,N_42793,N_42725);
and U43239 (N_43239,N_42571,N_42976);
xor U43240 (N_43240,N_42972,N_42910);
nor U43241 (N_43241,N_42964,N_42656);
nand U43242 (N_43242,N_42957,N_42803);
nand U43243 (N_43243,N_42925,N_42592);
nand U43244 (N_43244,N_42573,N_42713);
nand U43245 (N_43245,N_42901,N_42629);
nor U43246 (N_43246,N_42705,N_42559);
nand U43247 (N_43247,N_42506,N_42641);
nand U43248 (N_43248,N_42666,N_42732);
xor U43249 (N_43249,N_42710,N_42909);
nor U43250 (N_43250,N_42863,N_42623);
nand U43251 (N_43251,N_42886,N_42771);
xnor U43252 (N_43252,N_42942,N_42699);
nor U43253 (N_43253,N_42646,N_42612);
and U43254 (N_43254,N_42797,N_42970);
nand U43255 (N_43255,N_42970,N_42685);
xor U43256 (N_43256,N_42775,N_42761);
xnor U43257 (N_43257,N_42757,N_42533);
or U43258 (N_43258,N_42625,N_42571);
or U43259 (N_43259,N_42517,N_42782);
or U43260 (N_43260,N_42859,N_42611);
nand U43261 (N_43261,N_42586,N_42576);
or U43262 (N_43262,N_42604,N_42549);
or U43263 (N_43263,N_42857,N_42610);
and U43264 (N_43264,N_42794,N_42742);
and U43265 (N_43265,N_42641,N_42509);
nand U43266 (N_43266,N_42845,N_42965);
or U43267 (N_43267,N_42623,N_42947);
or U43268 (N_43268,N_42738,N_42679);
and U43269 (N_43269,N_42968,N_42932);
nor U43270 (N_43270,N_42768,N_42504);
xor U43271 (N_43271,N_42688,N_42555);
nor U43272 (N_43272,N_42901,N_42509);
xnor U43273 (N_43273,N_42758,N_42926);
nor U43274 (N_43274,N_42784,N_42853);
nor U43275 (N_43275,N_42584,N_42878);
nor U43276 (N_43276,N_42777,N_42786);
or U43277 (N_43277,N_42592,N_42686);
xor U43278 (N_43278,N_42877,N_42747);
or U43279 (N_43279,N_42703,N_42654);
nand U43280 (N_43280,N_42985,N_42929);
xor U43281 (N_43281,N_42537,N_42565);
or U43282 (N_43282,N_42729,N_42691);
xnor U43283 (N_43283,N_42599,N_42522);
and U43284 (N_43284,N_42861,N_42622);
or U43285 (N_43285,N_42895,N_42579);
or U43286 (N_43286,N_42754,N_42815);
and U43287 (N_43287,N_42904,N_42523);
xnor U43288 (N_43288,N_42850,N_42966);
xnor U43289 (N_43289,N_42899,N_42764);
xor U43290 (N_43290,N_42714,N_42927);
nand U43291 (N_43291,N_42966,N_42815);
nor U43292 (N_43292,N_42536,N_42919);
or U43293 (N_43293,N_42813,N_42652);
xnor U43294 (N_43294,N_42713,N_42744);
or U43295 (N_43295,N_42966,N_42897);
nand U43296 (N_43296,N_42556,N_42979);
nand U43297 (N_43297,N_42791,N_42560);
or U43298 (N_43298,N_42774,N_42641);
nand U43299 (N_43299,N_42682,N_42954);
nand U43300 (N_43300,N_42747,N_42608);
nor U43301 (N_43301,N_42693,N_42902);
nor U43302 (N_43302,N_42595,N_42733);
nand U43303 (N_43303,N_42891,N_42727);
or U43304 (N_43304,N_42659,N_42710);
and U43305 (N_43305,N_42717,N_42680);
nor U43306 (N_43306,N_42506,N_42587);
nor U43307 (N_43307,N_42781,N_42546);
xnor U43308 (N_43308,N_42913,N_42781);
xor U43309 (N_43309,N_42862,N_42937);
nor U43310 (N_43310,N_42815,N_42549);
and U43311 (N_43311,N_42542,N_42501);
nand U43312 (N_43312,N_42902,N_42751);
and U43313 (N_43313,N_42611,N_42870);
xor U43314 (N_43314,N_42842,N_42752);
nand U43315 (N_43315,N_42827,N_42584);
xor U43316 (N_43316,N_42846,N_42889);
nand U43317 (N_43317,N_42779,N_42516);
xor U43318 (N_43318,N_42680,N_42841);
xnor U43319 (N_43319,N_42910,N_42933);
nor U43320 (N_43320,N_42639,N_42882);
or U43321 (N_43321,N_42578,N_42958);
and U43322 (N_43322,N_42503,N_42774);
or U43323 (N_43323,N_42931,N_42557);
nand U43324 (N_43324,N_42637,N_42854);
or U43325 (N_43325,N_42614,N_42575);
and U43326 (N_43326,N_42614,N_42603);
xor U43327 (N_43327,N_42926,N_42940);
nand U43328 (N_43328,N_42622,N_42732);
xor U43329 (N_43329,N_42687,N_42795);
or U43330 (N_43330,N_42517,N_42925);
and U43331 (N_43331,N_42884,N_42613);
and U43332 (N_43332,N_42758,N_42879);
and U43333 (N_43333,N_42504,N_42923);
or U43334 (N_43334,N_42800,N_42628);
nand U43335 (N_43335,N_42817,N_42685);
or U43336 (N_43336,N_42648,N_42914);
nor U43337 (N_43337,N_42735,N_42822);
and U43338 (N_43338,N_42799,N_42968);
and U43339 (N_43339,N_42508,N_42820);
xor U43340 (N_43340,N_42708,N_42872);
or U43341 (N_43341,N_42571,N_42716);
and U43342 (N_43342,N_42889,N_42839);
nand U43343 (N_43343,N_42886,N_42842);
nor U43344 (N_43344,N_42818,N_42831);
nor U43345 (N_43345,N_42877,N_42920);
and U43346 (N_43346,N_42647,N_42897);
xnor U43347 (N_43347,N_42594,N_42954);
nor U43348 (N_43348,N_42681,N_42576);
nor U43349 (N_43349,N_42988,N_42552);
nor U43350 (N_43350,N_42829,N_42755);
and U43351 (N_43351,N_42889,N_42693);
nor U43352 (N_43352,N_42635,N_42556);
and U43353 (N_43353,N_42800,N_42762);
xnor U43354 (N_43354,N_42753,N_42580);
or U43355 (N_43355,N_42901,N_42764);
nand U43356 (N_43356,N_42934,N_42806);
and U43357 (N_43357,N_42963,N_42587);
xnor U43358 (N_43358,N_42754,N_42681);
xnor U43359 (N_43359,N_42740,N_42620);
and U43360 (N_43360,N_42629,N_42573);
nand U43361 (N_43361,N_42802,N_42912);
or U43362 (N_43362,N_42731,N_42963);
and U43363 (N_43363,N_42942,N_42613);
nand U43364 (N_43364,N_42549,N_42847);
xor U43365 (N_43365,N_42559,N_42977);
xnor U43366 (N_43366,N_42616,N_42507);
and U43367 (N_43367,N_42998,N_42665);
nor U43368 (N_43368,N_42660,N_42921);
nand U43369 (N_43369,N_42654,N_42951);
nand U43370 (N_43370,N_42537,N_42557);
xnor U43371 (N_43371,N_42736,N_42803);
nand U43372 (N_43372,N_42609,N_42751);
xor U43373 (N_43373,N_42501,N_42965);
xor U43374 (N_43374,N_42543,N_42697);
and U43375 (N_43375,N_42588,N_42585);
xnor U43376 (N_43376,N_42570,N_42700);
or U43377 (N_43377,N_42717,N_42939);
nand U43378 (N_43378,N_42557,N_42749);
or U43379 (N_43379,N_42866,N_42859);
nand U43380 (N_43380,N_42614,N_42980);
and U43381 (N_43381,N_42869,N_42503);
and U43382 (N_43382,N_42673,N_42995);
nor U43383 (N_43383,N_42976,N_42742);
nor U43384 (N_43384,N_42665,N_42648);
nand U43385 (N_43385,N_42904,N_42995);
nor U43386 (N_43386,N_42939,N_42817);
nand U43387 (N_43387,N_42983,N_42759);
xor U43388 (N_43388,N_42521,N_42591);
nand U43389 (N_43389,N_42695,N_42535);
or U43390 (N_43390,N_42506,N_42951);
nor U43391 (N_43391,N_42651,N_42900);
nand U43392 (N_43392,N_42621,N_42974);
and U43393 (N_43393,N_42943,N_42716);
or U43394 (N_43394,N_42664,N_42772);
or U43395 (N_43395,N_42869,N_42623);
or U43396 (N_43396,N_42736,N_42850);
or U43397 (N_43397,N_42670,N_42759);
nand U43398 (N_43398,N_42695,N_42566);
or U43399 (N_43399,N_42536,N_42893);
nor U43400 (N_43400,N_42754,N_42803);
nor U43401 (N_43401,N_42786,N_42962);
nand U43402 (N_43402,N_42620,N_42865);
nand U43403 (N_43403,N_42829,N_42733);
or U43404 (N_43404,N_42786,N_42631);
nor U43405 (N_43405,N_42886,N_42850);
or U43406 (N_43406,N_42747,N_42951);
nor U43407 (N_43407,N_42640,N_42873);
and U43408 (N_43408,N_42544,N_42858);
nor U43409 (N_43409,N_42894,N_42700);
and U43410 (N_43410,N_42606,N_42824);
nand U43411 (N_43411,N_42764,N_42979);
or U43412 (N_43412,N_42859,N_42621);
nand U43413 (N_43413,N_42883,N_42939);
nor U43414 (N_43414,N_42911,N_42748);
or U43415 (N_43415,N_42924,N_42878);
or U43416 (N_43416,N_42683,N_42693);
or U43417 (N_43417,N_42751,N_42935);
nor U43418 (N_43418,N_42630,N_42876);
or U43419 (N_43419,N_42648,N_42659);
nor U43420 (N_43420,N_42532,N_42857);
xor U43421 (N_43421,N_42527,N_42852);
nor U43422 (N_43422,N_42880,N_42605);
nor U43423 (N_43423,N_42780,N_42593);
or U43424 (N_43424,N_42811,N_42532);
nor U43425 (N_43425,N_42739,N_42790);
nand U43426 (N_43426,N_42905,N_42893);
xor U43427 (N_43427,N_42875,N_42753);
nor U43428 (N_43428,N_42807,N_42865);
or U43429 (N_43429,N_42941,N_42583);
and U43430 (N_43430,N_42943,N_42688);
nor U43431 (N_43431,N_42740,N_42558);
and U43432 (N_43432,N_42913,N_42873);
and U43433 (N_43433,N_42722,N_42581);
nor U43434 (N_43434,N_42965,N_42559);
xor U43435 (N_43435,N_42635,N_42527);
xnor U43436 (N_43436,N_42663,N_42898);
and U43437 (N_43437,N_42982,N_42816);
xor U43438 (N_43438,N_42531,N_42539);
xnor U43439 (N_43439,N_42941,N_42600);
nor U43440 (N_43440,N_42609,N_42822);
xnor U43441 (N_43441,N_42556,N_42872);
nand U43442 (N_43442,N_42889,N_42502);
xnor U43443 (N_43443,N_42616,N_42788);
nor U43444 (N_43444,N_42857,N_42585);
or U43445 (N_43445,N_42731,N_42712);
nand U43446 (N_43446,N_42829,N_42594);
or U43447 (N_43447,N_42992,N_42635);
and U43448 (N_43448,N_42615,N_42894);
and U43449 (N_43449,N_42613,N_42991);
xor U43450 (N_43450,N_42507,N_42989);
nand U43451 (N_43451,N_42584,N_42710);
and U43452 (N_43452,N_42731,N_42876);
nand U43453 (N_43453,N_42729,N_42749);
nor U43454 (N_43454,N_42920,N_42702);
nor U43455 (N_43455,N_42683,N_42533);
xor U43456 (N_43456,N_42751,N_42554);
nand U43457 (N_43457,N_42710,N_42575);
xor U43458 (N_43458,N_42785,N_42848);
or U43459 (N_43459,N_42864,N_42812);
nand U43460 (N_43460,N_42517,N_42722);
or U43461 (N_43461,N_42697,N_42569);
xor U43462 (N_43462,N_42933,N_42897);
xnor U43463 (N_43463,N_42544,N_42872);
nor U43464 (N_43464,N_42646,N_42982);
nor U43465 (N_43465,N_42587,N_42546);
xor U43466 (N_43466,N_42576,N_42696);
xor U43467 (N_43467,N_42610,N_42531);
or U43468 (N_43468,N_42887,N_42674);
nand U43469 (N_43469,N_42766,N_42792);
xor U43470 (N_43470,N_42532,N_42564);
and U43471 (N_43471,N_42627,N_42672);
or U43472 (N_43472,N_42835,N_42574);
and U43473 (N_43473,N_42749,N_42997);
or U43474 (N_43474,N_42919,N_42557);
or U43475 (N_43475,N_42918,N_42860);
nand U43476 (N_43476,N_42622,N_42593);
and U43477 (N_43477,N_42605,N_42734);
nand U43478 (N_43478,N_42846,N_42653);
nand U43479 (N_43479,N_42940,N_42641);
nand U43480 (N_43480,N_42926,N_42996);
or U43481 (N_43481,N_42732,N_42582);
or U43482 (N_43482,N_42993,N_42763);
nor U43483 (N_43483,N_42554,N_42571);
xnor U43484 (N_43484,N_42855,N_42943);
and U43485 (N_43485,N_42593,N_42581);
nor U43486 (N_43486,N_42503,N_42738);
and U43487 (N_43487,N_42760,N_42912);
nand U43488 (N_43488,N_42993,N_42671);
nand U43489 (N_43489,N_42838,N_42884);
nand U43490 (N_43490,N_42944,N_42868);
xor U43491 (N_43491,N_42903,N_42877);
and U43492 (N_43492,N_42832,N_42726);
nor U43493 (N_43493,N_42606,N_42878);
nand U43494 (N_43494,N_42952,N_42843);
nand U43495 (N_43495,N_42500,N_42905);
xnor U43496 (N_43496,N_42795,N_42971);
xnor U43497 (N_43497,N_42508,N_42551);
and U43498 (N_43498,N_42788,N_42778);
nor U43499 (N_43499,N_42669,N_42870);
and U43500 (N_43500,N_43386,N_43079);
nor U43501 (N_43501,N_43342,N_43279);
nand U43502 (N_43502,N_43480,N_43004);
xor U43503 (N_43503,N_43315,N_43312);
nor U43504 (N_43504,N_43120,N_43154);
and U43505 (N_43505,N_43038,N_43437);
nor U43506 (N_43506,N_43493,N_43284);
or U43507 (N_43507,N_43141,N_43113);
nor U43508 (N_43508,N_43155,N_43186);
nand U43509 (N_43509,N_43267,N_43462);
xor U43510 (N_43510,N_43081,N_43161);
and U43511 (N_43511,N_43395,N_43045);
and U43512 (N_43512,N_43160,N_43418);
nand U43513 (N_43513,N_43227,N_43291);
and U43514 (N_43514,N_43010,N_43104);
nand U43515 (N_43515,N_43457,N_43020);
and U43516 (N_43516,N_43373,N_43427);
xor U43517 (N_43517,N_43217,N_43230);
or U43518 (N_43518,N_43429,N_43093);
and U43519 (N_43519,N_43261,N_43371);
nor U43520 (N_43520,N_43002,N_43456);
and U43521 (N_43521,N_43269,N_43233);
nor U43522 (N_43522,N_43087,N_43080);
and U43523 (N_43523,N_43276,N_43363);
nor U43524 (N_43524,N_43182,N_43253);
xor U43525 (N_43525,N_43460,N_43213);
nand U43526 (N_43526,N_43466,N_43320);
and U43527 (N_43527,N_43194,N_43376);
nand U43528 (N_43528,N_43127,N_43056);
or U43529 (N_43529,N_43058,N_43409);
xnor U43530 (N_43530,N_43417,N_43378);
nor U43531 (N_43531,N_43325,N_43072);
or U43532 (N_43532,N_43359,N_43412);
nor U43533 (N_43533,N_43467,N_43064);
nor U43534 (N_43534,N_43228,N_43132);
nor U43535 (N_43535,N_43135,N_43201);
and U43536 (N_43536,N_43381,N_43245);
and U43537 (N_43537,N_43257,N_43030);
nor U43538 (N_43538,N_43443,N_43482);
nor U43539 (N_43539,N_43259,N_43232);
and U43540 (N_43540,N_43111,N_43470);
and U43541 (N_43541,N_43098,N_43049);
xor U43542 (N_43542,N_43024,N_43164);
nand U43543 (N_43543,N_43102,N_43313);
xor U43544 (N_43544,N_43190,N_43203);
or U43545 (N_43545,N_43234,N_43296);
nor U43546 (N_43546,N_43198,N_43212);
and U43547 (N_43547,N_43413,N_43444);
nand U43548 (N_43548,N_43076,N_43174);
nor U43549 (N_43549,N_43214,N_43177);
nand U43550 (N_43550,N_43235,N_43299);
and U43551 (N_43551,N_43314,N_43026);
xnor U43552 (N_43552,N_43294,N_43389);
xor U43553 (N_43553,N_43490,N_43035);
and U43554 (N_43554,N_43330,N_43481);
nand U43555 (N_43555,N_43398,N_43451);
xor U43556 (N_43556,N_43239,N_43472);
xor U43557 (N_43557,N_43434,N_43083);
nor U43558 (N_43558,N_43463,N_43420);
xnor U43559 (N_43559,N_43143,N_43303);
nor U43560 (N_43560,N_43000,N_43370);
or U43561 (N_43561,N_43461,N_43029);
and U43562 (N_43562,N_43331,N_43032);
xor U43563 (N_43563,N_43069,N_43277);
or U43564 (N_43564,N_43345,N_43290);
nor U43565 (N_43565,N_43175,N_43243);
and U43566 (N_43566,N_43487,N_43469);
xnor U43567 (N_43567,N_43326,N_43268);
xor U43568 (N_43568,N_43005,N_43116);
xor U43569 (N_43569,N_43343,N_43388);
nor U43570 (N_43570,N_43438,N_43131);
nor U43571 (N_43571,N_43448,N_43248);
and U43572 (N_43572,N_43360,N_43210);
and U43573 (N_43573,N_43014,N_43484);
xor U43574 (N_43574,N_43346,N_43393);
xnor U43575 (N_43575,N_43258,N_43496);
xnor U43576 (N_43576,N_43163,N_43109);
nand U43577 (N_43577,N_43282,N_43449);
xor U43578 (N_43578,N_43464,N_43138);
nand U43579 (N_43579,N_43415,N_43452);
or U43580 (N_43580,N_43231,N_43297);
nand U43581 (N_43581,N_43183,N_43051);
or U43582 (N_43582,N_43317,N_43099);
nand U43583 (N_43583,N_43421,N_43157);
nor U43584 (N_43584,N_43324,N_43499);
nand U43585 (N_43585,N_43065,N_43125);
nand U43586 (N_43586,N_43059,N_43355);
nand U43587 (N_43587,N_43329,N_43424);
xor U43588 (N_43588,N_43139,N_43216);
nand U43589 (N_43589,N_43105,N_43226);
and U43590 (N_43590,N_43328,N_43078);
nor U43591 (N_43591,N_43274,N_43488);
nand U43592 (N_43592,N_43357,N_43218);
nor U43593 (N_43593,N_43436,N_43430);
and U43594 (N_43594,N_43492,N_43319);
nand U43595 (N_43595,N_43077,N_43341);
or U43596 (N_43596,N_43396,N_43361);
nor U43597 (N_43597,N_43440,N_43273);
nand U43598 (N_43598,N_43364,N_43044);
nor U43599 (N_43599,N_43455,N_43205);
nor U43600 (N_43600,N_43095,N_43407);
or U43601 (N_43601,N_43408,N_43298);
or U43602 (N_43602,N_43247,N_43433);
nand U43603 (N_43603,N_43073,N_43166);
or U43604 (N_43604,N_43411,N_43318);
nor U43605 (N_43605,N_43327,N_43285);
nor U43606 (N_43606,N_43442,N_43144);
and U43607 (N_43607,N_43167,N_43446);
xnor U43608 (N_43608,N_43074,N_43366);
and U43609 (N_43609,N_43375,N_43292);
nand U43610 (N_43610,N_43251,N_43071);
nor U43611 (N_43611,N_43018,N_43097);
xor U43612 (N_43612,N_43075,N_43220);
or U43613 (N_43613,N_43060,N_43252);
nand U43614 (N_43614,N_43088,N_43196);
and U43615 (N_43615,N_43170,N_43333);
and U43616 (N_43616,N_43459,N_43255);
or U43617 (N_43617,N_43124,N_43180);
and U43618 (N_43618,N_43383,N_43053);
xor U43619 (N_43619,N_43265,N_43392);
or U43620 (N_43620,N_43256,N_43221);
xnor U43621 (N_43621,N_43168,N_43114);
and U43622 (N_43622,N_43202,N_43382);
nor U43623 (N_43623,N_43070,N_43305);
xor U43624 (N_43624,N_43391,N_43184);
nand U43625 (N_43625,N_43181,N_43435);
nor U43626 (N_43626,N_43385,N_43066);
nor U43627 (N_43627,N_43414,N_43300);
nand U43628 (N_43628,N_43036,N_43169);
nor U43629 (N_43629,N_43108,N_43179);
or U43630 (N_43630,N_43445,N_43034);
and U43631 (N_43631,N_43263,N_43050);
or U43632 (N_43632,N_43368,N_43009);
nand U43633 (N_43633,N_43309,N_43339);
xor U43634 (N_43634,N_43483,N_43468);
nand U43635 (N_43635,N_43426,N_43023);
nor U43636 (N_43636,N_43416,N_43047);
xnor U43637 (N_43637,N_43473,N_43195);
nor U43638 (N_43638,N_43362,N_43063);
xnor U43639 (N_43639,N_43046,N_43447);
nor U43640 (N_43640,N_43206,N_43374);
or U43641 (N_43641,N_43377,N_43260);
xnor U43642 (N_43642,N_43062,N_43117);
nand U43643 (N_43643,N_43092,N_43402);
and U43644 (N_43644,N_43208,N_43275);
nor U43645 (N_43645,N_43061,N_43241);
xnor U43646 (N_43646,N_43441,N_43096);
and U43647 (N_43647,N_43478,N_43187);
and U43648 (N_43648,N_43338,N_43089);
nor U43649 (N_43649,N_43425,N_43021);
and U43650 (N_43650,N_43013,N_43367);
nor U43651 (N_43651,N_43107,N_43025);
or U43652 (N_43652,N_43335,N_43322);
or U43653 (N_43653,N_43146,N_43489);
or U43654 (N_43654,N_43240,N_43118);
and U43655 (N_43655,N_43136,N_43110);
nand U43656 (N_43656,N_43176,N_43085);
xnor U43657 (N_43657,N_43165,N_43281);
and U43658 (N_43658,N_43308,N_43067);
xnor U43659 (N_43659,N_43011,N_43207);
and U43660 (N_43660,N_43422,N_43498);
or U43661 (N_43661,N_43151,N_43140);
xor U43662 (N_43662,N_43115,N_43171);
or U43663 (N_43663,N_43348,N_43310);
and U43664 (N_43664,N_43204,N_43497);
xor U43665 (N_43665,N_43152,N_43185);
nand U43666 (N_43666,N_43121,N_43428);
nor U43667 (N_43667,N_43399,N_43017);
xnor U43668 (N_43668,N_43350,N_43307);
xnor U43669 (N_43669,N_43304,N_43356);
or U43670 (N_43670,N_43254,N_43486);
xor U43671 (N_43671,N_43271,N_43145);
and U43672 (N_43672,N_43380,N_43028);
nor U43673 (N_43673,N_43354,N_43055);
nand U43674 (N_43674,N_43323,N_43397);
nand U43675 (N_43675,N_43090,N_43224);
nor U43676 (N_43676,N_43403,N_43142);
nand U43677 (N_43677,N_43321,N_43037);
nand U43678 (N_43678,N_43008,N_43122);
xnor U43679 (N_43679,N_43134,N_43347);
and U43680 (N_43680,N_43494,N_43130);
nand U43681 (N_43681,N_43178,N_43236);
or U43682 (N_43682,N_43302,N_43401);
or U43683 (N_43683,N_43003,N_43400);
xnor U43684 (N_43684,N_43027,N_43293);
or U43685 (N_43685,N_43040,N_43148);
or U43686 (N_43686,N_43351,N_43015);
nand U43687 (N_43687,N_43340,N_43172);
xor U43688 (N_43688,N_43225,N_43439);
xnor U43689 (N_43689,N_43129,N_43237);
xor U43690 (N_43690,N_43147,N_43474);
nor U43691 (N_43691,N_43068,N_43091);
or U43692 (N_43692,N_43458,N_43280);
nand U43693 (N_43693,N_43272,N_43344);
or U43694 (N_43694,N_43001,N_43287);
or U43695 (N_43695,N_43211,N_43485);
or U43696 (N_43696,N_43336,N_43229);
xnor U43697 (N_43697,N_43126,N_43301);
and U43698 (N_43698,N_43406,N_43054);
nor U43699 (N_43699,N_43453,N_43387);
nand U43700 (N_43700,N_43188,N_43016);
xor U43701 (N_43701,N_43223,N_43153);
or U43702 (N_43702,N_43365,N_43192);
or U43703 (N_43703,N_43022,N_43082);
nor U43704 (N_43704,N_43286,N_43238);
xnor U43705 (N_43705,N_43222,N_43033);
nand U43706 (N_43706,N_43283,N_43158);
and U43707 (N_43707,N_43423,N_43191);
or U43708 (N_43708,N_43100,N_43173);
and U43709 (N_43709,N_43159,N_43103);
xnor U43710 (N_43710,N_43244,N_43052);
nand U43711 (N_43711,N_43193,N_43012);
nor U43712 (N_43712,N_43200,N_43479);
nand U43713 (N_43713,N_43048,N_43316);
xnor U43714 (N_43714,N_43431,N_43379);
nor U43715 (N_43715,N_43197,N_43476);
nand U43716 (N_43716,N_43358,N_43289);
and U43717 (N_43717,N_43369,N_43199);
xnor U43718 (N_43718,N_43349,N_43128);
or U43719 (N_43719,N_43306,N_43043);
nand U43720 (N_43720,N_43086,N_43019);
nand U43721 (N_43721,N_43311,N_43249);
and U43722 (N_43722,N_43278,N_43133);
or U43723 (N_43723,N_43465,N_43123);
nor U43724 (N_43724,N_43006,N_43041);
nand U43725 (N_43725,N_43264,N_43150);
nand U43726 (N_43726,N_43334,N_43390);
and U43727 (N_43727,N_43353,N_43262);
and U43728 (N_43728,N_43372,N_43394);
or U43729 (N_43729,N_43112,N_43471);
nand U43730 (N_43730,N_43162,N_43491);
nor U43731 (N_43731,N_43242,N_43219);
nand U43732 (N_43732,N_43149,N_43432);
nand U43733 (N_43733,N_43410,N_43495);
xor U43734 (N_43734,N_43137,N_43209);
nand U43735 (N_43735,N_43106,N_43384);
or U43736 (N_43736,N_43405,N_43454);
nand U43737 (N_43737,N_43042,N_43189);
or U43738 (N_43738,N_43404,N_43475);
or U43739 (N_43739,N_43215,N_43352);
nor U43740 (N_43740,N_43094,N_43450);
nor U43741 (N_43741,N_43288,N_43101);
and U43742 (N_43742,N_43031,N_43332);
or U43743 (N_43743,N_43084,N_43270);
nor U43744 (N_43744,N_43250,N_43057);
nor U43745 (N_43745,N_43246,N_43119);
nor U43746 (N_43746,N_43337,N_43266);
or U43747 (N_43747,N_43007,N_43295);
and U43748 (N_43748,N_43156,N_43477);
xor U43749 (N_43749,N_43419,N_43039);
or U43750 (N_43750,N_43047,N_43110);
nand U43751 (N_43751,N_43159,N_43358);
nor U43752 (N_43752,N_43138,N_43238);
nand U43753 (N_43753,N_43337,N_43067);
xor U43754 (N_43754,N_43451,N_43304);
or U43755 (N_43755,N_43257,N_43089);
or U43756 (N_43756,N_43468,N_43382);
nand U43757 (N_43757,N_43415,N_43266);
and U43758 (N_43758,N_43029,N_43463);
nor U43759 (N_43759,N_43091,N_43285);
and U43760 (N_43760,N_43256,N_43481);
and U43761 (N_43761,N_43005,N_43203);
and U43762 (N_43762,N_43449,N_43461);
nand U43763 (N_43763,N_43057,N_43232);
or U43764 (N_43764,N_43101,N_43316);
nand U43765 (N_43765,N_43446,N_43116);
and U43766 (N_43766,N_43427,N_43399);
xnor U43767 (N_43767,N_43367,N_43193);
nand U43768 (N_43768,N_43131,N_43284);
or U43769 (N_43769,N_43286,N_43219);
nor U43770 (N_43770,N_43476,N_43442);
and U43771 (N_43771,N_43174,N_43071);
nor U43772 (N_43772,N_43344,N_43049);
xnor U43773 (N_43773,N_43371,N_43320);
nor U43774 (N_43774,N_43221,N_43047);
and U43775 (N_43775,N_43404,N_43004);
or U43776 (N_43776,N_43312,N_43281);
and U43777 (N_43777,N_43036,N_43498);
nor U43778 (N_43778,N_43404,N_43441);
or U43779 (N_43779,N_43336,N_43481);
or U43780 (N_43780,N_43177,N_43357);
or U43781 (N_43781,N_43446,N_43179);
nor U43782 (N_43782,N_43010,N_43036);
and U43783 (N_43783,N_43395,N_43439);
or U43784 (N_43784,N_43326,N_43216);
and U43785 (N_43785,N_43289,N_43051);
and U43786 (N_43786,N_43454,N_43047);
xor U43787 (N_43787,N_43195,N_43239);
nor U43788 (N_43788,N_43293,N_43010);
or U43789 (N_43789,N_43191,N_43186);
or U43790 (N_43790,N_43396,N_43132);
or U43791 (N_43791,N_43187,N_43400);
xor U43792 (N_43792,N_43248,N_43019);
nand U43793 (N_43793,N_43380,N_43434);
nand U43794 (N_43794,N_43461,N_43006);
nor U43795 (N_43795,N_43313,N_43177);
nand U43796 (N_43796,N_43413,N_43027);
nand U43797 (N_43797,N_43348,N_43154);
nor U43798 (N_43798,N_43448,N_43099);
and U43799 (N_43799,N_43201,N_43147);
nand U43800 (N_43800,N_43342,N_43180);
and U43801 (N_43801,N_43101,N_43260);
and U43802 (N_43802,N_43016,N_43174);
nor U43803 (N_43803,N_43277,N_43097);
nand U43804 (N_43804,N_43457,N_43367);
and U43805 (N_43805,N_43191,N_43072);
and U43806 (N_43806,N_43033,N_43398);
and U43807 (N_43807,N_43390,N_43485);
and U43808 (N_43808,N_43247,N_43298);
nand U43809 (N_43809,N_43108,N_43307);
nand U43810 (N_43810,N_43030,N_43208);
or U43811 (N_43811,N_43328,N_43106);
xnor U43812 (N_43812,N_43434,N_43420);
xnor U43813 (N_43813,N_43388,N_43263);
or U43814 (N_43814,N_43140,N_43312);
xor U43815 (N_43815,N_43034,N_43264);
and U43816 (N_43816,N_43218,N_43035);
xor U43817 (N_43817,N_43403,N_43419);
and U43818 (N_43818,N_43192,N_43166);
and U43819 (N_43819,N_43394,N_43366);
and U43820 (N_43820,N_43340,N_43461);
or U43821 (N_43821,N_43471,N_43419);
nor U43822 (N_43822,N_43475,N_43336);
or U43823 (N_43823,N_43409,N_43157);
or U43824 (N_43824,N_43120,N_43106);
xor U43825 (N_43825,N_43387,N_43466);
and U43826 (N_43826,N_43325,N_43160);
and U43827 (N_43827,N_43302,N_43186);
and U43828 (N_43828,N_43361,N_43160);
nor U43829 (N_43829,N_43272,N_43097);
xor U43830 (N_43830,N_43443,N_43093);
and U43831 (N_43831,N_43034,N_43073);
or U43832 (N_43832,N_43313,N_43112);
nand U43833 (N_43833,N_43487,N_43030);
or U43834 (N_43834,N_43363,N_43487);
and U43835 (N_43835,N_43262,N_43467);
and U43836 (N_43836,N_43468,N_43458);
nand U43837 (N_43837,N_43147,N_43456);
nand U43838 (N_43838,N_43442,N_43092);
nor U43839 (N_43839,N_43282,N_43230);
and U43840 (N_43840,N_43005,N_43426);
and U43841 (N_43841,N_43360,N_43288);
and U43842 (N_43842,N_43226,N_43240);
xor U43843 (N_43843,N_43478,N_43278);
and U43844 (N_43844,N_43259,N_43474);
and U43845 (N_43845,N_43351,N_43137);
nor U43846 (N_43846,N_43412,N_43160);
xor U43847 (N_43847,N_43164,N_43034);
and U43848 (N_43848,N_43141,N_43050);
nand U43849 (N_43849,N_43108,N_43185);
or U43850 (N_43850,N_43193,N_43291);
nor U43851 (N_43851,N_43356,N_43065);
nor U43852 (N_43852,N_43414,N_43446);
or U43853 (N_43853,N_43398,N_43449);
and U43854 (N_43854,N_43015,N_43174);
or U43855 (N_43855,N_43372,N_43177);
nand U43856 (N_43856,N_43121,N_43186);
nor U43857 (N_43857,N_43439,N_43327);
xor U43858 (N_43858,N_43290,N_43279);
or U43859 (N_43859,N_43429,N_43087);
and U43860 (N_43860,N_43419,N_43070);
nor U43861 (N_43861,N_43475,N_43101);
nand U43862 (N_43862,N_43363,N_43040);
and U43863 (N_43863,N_43030,N_43052);
or U43864 (N_43864,N_43212,N_43335);
xor U43865 (N_43865,N_43421,N_43023);
or U43866 (N_43866,N_43147,N_43367);
xnor U43867 (N_43867,N_43495,N_43317);
and U43868 (N_43868,N_43352,N_43194);
nor U43869 (N_43869,N_43282,N_43026);
nor U43870 (N_43870,N_43486,N_43255);
nand U43871 (N_43871,N_43097,N_43218);
xor U43872 (N_43872,N_43135,N_43091);
and U43873 (N_43873,N_43128,N_43463);
nand U43874 (N_43874,N_43291,N_43211);
nand U43875 (N_43875,N_43423,N_43253);
xor U43876 (N_43876,N_43256,N_43052);
and U43877 (N_43877,N_43314,N_43193);
nor U43878 (N_43878,N_43172,N_43237);
nor U43879 (N_43879,N_43081,N_43121);
nand U43880 (N_43880,N_43309,N_43009);
and U43881 (N_43881,N_43264,N_43300);
xnor U43882 (N_43882,N_43378,N_43233);
and U43883 (N_43883,N_43070,N_43351);
and U43884 (N_43884,N_43032,N_43034);
xnor U43885 (N_43885,N_43299,N_43158);
or U43886 (N_43886,N_43246,N_43121);
nand U43887 (N_43887,N_43166,N_43222);
nor U43888 (N_43888,N_43332,N_43416);
nor U43889 (N_43889,N_43227,N_43161);
nand U43890 (N_43890,N_43005,N_43141);
nand U43891 (N_43891,N_43196,N_43010);
nor U43892 (N_43892,N_43090,N_43189);
and U43893 (N_43893,N_43405,N_43469);
nor U43894 (N_43894,N_43258,N_43144);
and U43895 (N_43895,N_43101,N_43395);
or U43896 (N_43896,N_43057,N_43446);
nand U43897 (N_43897,N_43204,N_43102);
nor U43898 (N_43898,N_43265,N_43466);
or U43899 (N_43899,N_43426,N_43192);
or U43900 (N_43900,N_43113,N_43365);
nor U43901 (N_43901,N_43469,N_43483);
xor U43902 (N_43902,N_43014,N_43375);
or U43903 (N_43903,N_43052,N_43387);
or U43904 (N_43904,N_43199,N_43465);
or U43905 (N_43905,N_43471,N_43188);
xor U43906 (N_43906,N_43442,N_43138);
or U43907 (N_43907,N_43486,N_43220);
xor U43908 (N_43908,N_43053,N_43001);
and U43909 (N_43909,N_43185,N_43010);
xnor U43910 (N_43910,N_43329,N_43068);
xnor U43911 (N_43911,N_43182,N_43446);
nor U43912 (N_43912,N_43027,N_43461);
or U43913 (N_43913,N_43136,N_43315);
nand U43914 (N_43914,N_43458,N_43489);
xnor U43915 (N_43915,N_43080,N_43453);
nand U43916 (N_43916,N_43054,N_43486);
nand U43917 (N_43917,N_43100,N_43075);
or U43918 (N_43918,N_43499,N_43221);
nor U43919 (N_43919,N_43056,N_43159);
nand U43920 (N_43920,N_43111,N_43340);
nand U43921 (N_43921,N_43010,N_43482);
nor U43922 (N_43922,N_43244,N_43437);
nand U43923 (N_43923,N_43166,N_43396);
nor U43924 (N_43924,N_43191,N_43471);
and U43925 (N_43925,N_43456,N_43220);
or U43926 (N_43926,N_43126,N_43487);
or U43927 (N_43927,N_43211,N_43142);
nor U43928 (N_43928,N_43372,N_43174);
xor U43929 (N_43929,N_43154,N_43393);
xor U43930 (N_43930,N_43409,N_43299);
and U43931 (N_43931,N_43303,N_43190);
nor U43932 (N_43932,N_43454,N_43255);
nand U43933 (N_43933,N_43336,N_43196);
nand U43934 (N_43934,N_43019,N_43332);
and U43935 (N_43935,N_43461,N_43156);
or U43936 (N_43936,N_43382,N_43466);
or U43937 (N_43937,N_43077,N_43199);
xor U43938 (N_43938,N_43311,N_43490);
nor U43939 (N_43939,N_43489,N_43141);
nand U43940 (N_43940,N_43282,N_43305);
nor U43941 (N_43941,N_43285,N_43476);
or U43942 (N_43942,N_43206,N_43086);
nor U43943 (N_43943,N_43460,N_43040);
or U43944 (N_43944,N_43067,N_43484);
and U43945 (N_43945,N_43011,N_43470);
nand U43946 (N_43946,N_43332,N_43078);
and U43947 (N_43947,N_43372,N_43478);
nand U43948 (N_43948,N_43053,N_43176);
xnor U43949 (N_43949,N_43140,N_43145);
xnor U43950 (N_43950,N_43324,N_43283);
or U43951 (N_43951,N_43365,N_43071);
and U43952 (N_43952,N_43470,N_43160);
nor U43953 (N_43953,N_43437,N_43429);
nor U43954 (N_43954,N_43003,N_43292);
or U43955 (N_43955,N_43240,N_43405);
and U43956 (N_43956,N_43448,N_43138);
nor U43957 (N_43957,N_43042,N_43296);
nor U43958 (N_43958,N_43018,N_43374);
nor U43959 (N_43959,N_43375,N_43377);
nor U43960 (N_43960,N_43151,N_43084);
or U43961 (N_43961,N_43197,N_43115);
xnor U43962 (N_43962,N_43141,N_43028);
xor U43963 (N_43963,N_43115,N_43396);
and U43964 (N_43964,N_43153,N_43481);
and U43965 (N_43965,N_43264,N_43467);
or U43966 (N_43966,N_43367,N_43043);
nor U43967 (N_43967,N_43428,N_43409);
nand U43968 (N_43968,N_43355,N_43171);
or U43969 (N_43969,N_43292,N_43425);
nand U43970 (N_43970,N_43126,N_43470);
nand U43971 (N_43971,N_43436,N_43105);
nand U43972 (N_43972,N_43023,N_43391);
nor U43973 (N_43973,N_43286,N_43309);
xnor U43974 (N_43974,N_43362,N_43485);
or U43975 (N_43975,N_43399,N_43043);
or U43976 (N_43976,N_43273,N_43469);
xor U43977 (N_43977,N_43111,N_43291);
or U43978 (N_43978,N_43448,N_43069);
and U43979 (N_43979,N_43407,N_43268);
and U43980 (N_43980,N_43479,N_43345);
or U43981 (N_43981,N_43066,N_43084);
nor U43982 (N_43982,N_43210,N_43475);
nand U43983 (N_43983,N_43343,N_43004);
or U43984 (N_43984,N_43258,N_43285);
or U43985 (N_43985,N_43374,N_43416);
nand U43986 (N_43986,N_43445,N_43278);
nand U43987 (N_43987,N_43010,N_43055);
or U43988 (N_43988,N_43498,N_43052);
nand U43989 (N_43989,N_43086,N_43171);
xnor U43990 (N_43990,N_43415,N_43441);
nand U43991 (N_43991,N_43321,N_43285);
or U43992 (N_43992,N_43099,N_43282);
xor U43993 (N_43993,N_43010,N_43422);
and U43994 (N_43994,N_43064,N_43179);
xnor U43995 (N_43995,N_43249,N_43298);
nand U43996 (N_43996,N_43075,N_43032);
or U43997 (N_43997,N_43310,N_43261);
nor U43998 (N_43998,N_43131,N_43088);
or U43999 (N_43999,N_43326,N_43361);
nor U44000 (N_44000,N_43900,N_43576);
nor U44001 (N_44001,N_43536,N_43727);
xnor U44002 (N_44002,N_43748,N_43679);
nor U44003 (N_44003,N_43511,N_43983);
and U44004 (N_44004,N_43724,N_43729);
nand U44005 (N_44005,N_43858,N_43598);
xor U44006 (N_44006,N_43938,N_43730);
or U44007 (N_44007,N_43524,N_43537);
nor U44008 (N_44008,N_43774,N_43844);
nor U44009 (N_44009,N_43696,N_43712);
nand U44010 (N_44010,N_43606,N_43892);
nor U44011 (N_44011,N_43761,N_43830);
or U44012 (N_44012,N_43801,N_43673);
nand U44013 (N_44013,N_43957,N_43765);
and U44014 (N_44014,N_43716,N_43921);
and U44015 (N_44015,N_43776,N_43956);
xnor U44016 (N_44016,N_43602,N_43969);
nor U44017 (N_44017,N_43722,N_43790);
nand U44018 (N_44018,N_43793,N_43914);
nand U44019 (N_44019,N_43740,N_43670);
xor U44020 (N_44020,N_43661,N_43936);
and U44021 (N_44021,N_43820,N_43944);
and U44022 (N_44022,N_43866,N_43757);
or U44023 (N_44023,N_43982,N_43720);
xor U44024 (N_44024,N_43996,N_43648);
nor U44025 (N_44025,N_43539,N_43630);
nand U44026 (N_44026,N_43633,N_43706);
nor U44027 (N_44027,N_43736,N_43711);
and U44028 (N_44028,N_43547,N_43560);
nand U44029 (N_44029,N_43591,N_43840);
xnor U44030 (N_44030,N_43680,N_43526);
or U44031 (N_44031,N_43521,N_43718);
or U44032 (N_44032,N_43653,N_43886);
or U44033 (N_44033,N_43584,N_43566);
nand U44034 (N_44034,N_43752,N_43565);
xor U44035 (N_44035,N_43617,N_43906);
and U44036 (N_44036,N_43616,N_43703);
and U44037 (N_44037,N_43932,N_43814);
and U44038 (N_44038,N_43753,N_43762);
xnor U44039 (N_44039,N_43634,N_43658);
or U44040 (N_44040,N_43891,N_43802);
xor U44041 (N_44041,N_43845,N_43501);
nor U44042 (N_44042,N_43502,N_43843);
or U44043 (N_44043,N_43636,N_43555);
nor U44044 (N_44044,N_43698,N_43756);
nand U44045 (N_44045,N_43940,N_43933);
or U44046 (N_44046,N_43950,N_43794);
nor U44047 (N_44047,N_43859,N_43846);
nor U44048 (N_44048,N_43901,N_43682);
nand U44049 (N_44049,N_43963,N_43855);
or U44050 (N_44050,N_43717,N_43702);
xnor U44051 (N_44051,N_43595,N_43553);
nand U44052 (N_44052,N_43918,N_43807);
and U44053 (N_44053,N_43659,N_43579);
nand U44054 (N_44054,N_43784,N_43640);
and U44055 (N_44055,N_43990,N_43671);
nand U44056 (N_44056,N_43764,N_43614);
xor U44057 (N_44057,N_43934,N_43751);
and U44058 (N_44058,N_43734,N_43500);
xnor U44059 (N_44059,N_43687,N_43834);
and U44060 (N_44060,N_43719,N_43985);
nand U44061 (N_44061,N_43898,N_43625);
and U44062 (N_44062,N_43605,N_43828);
or U44063 (N_44063,N_43979,N_43540);
and U44064 (N_44064,N_43758,N_43541);
or U44065 (N_44065,N_43667,N_43574);
and U44066 (N_44066,N_43577,N_43709);
xnor U44067 (N_44067,N_43604,N_43533);
xor U44068 (N_44068,N_43965,N_43905);
and U44069 (N_44069,N_43833,N_43903);
or U44070 (N_44070,N_43563,N_43582);
nor U44071 (N_44071,N_43767,N_43980);
nand U44072 (N_44072,N_43791,N_43863);
and U44073 (N_44073,N_43554,N_43623);
and U44074 (N_44074,N_43657,N_43975);
nor U44075 (N_44075,N_43699,N_43650);
nor U44076 (N_44076,N_43781,N_43885);
nor U44077 (N_44077,N_43988,N_43912);
and U44078 (N_44078,N_43690,N_43745);
and U44079 (N_44079,N_43970,N_43949);
nor U44080 (N_44080,N_43775,N_43947);
or U44081 (N_44081,N_43742,N_43763);
nand U44082 (N_44082,N_43622,N_43773);
xor U44083 (N_44083,N_43964,N_43888);
nand U44084 (N_44084,N_43824,N_43816);
nor U44085 (N_44085,N_43839,N_43894);
and U44086 (N_44086,N_43851,N_43655);
nand U44087 (N_44087,N_43935,N_43631);
xor U44088 (N_44088,N_43989,N_43545);
xor U44089 (N_44089,N_43779,N_43798);
nand U44090 (N_44090,N_43946,N_43731);
and U44091 (N_44091,N_43860,N_43583);
nor U44092 (N_44092,N_43567,N_43676);
nor U44093 (N_44093,N_43660,N_43805);
nor U44094 (N_44094,N_43741,N_43505);
nor U44095 (N_44095,N_43827,N_43662);
xnor U44096 (N_44096,N_43991,N_43564);
nor U44097 (N_44097,N_43873,N_43909);
xnor U44098 (N_44098,N_43506,N_43823);
nor U44099 (N_44099,N_43994,N_43683);
and U44100 (N_44100,N_43872,N_43997);
or U44101 (N_44101,N_43896,N_43869);
nor U44102 (N_44102,N_43966,N_43590);
nand U44103 (N_44103,N_43608,N_43871);
and U44104 (N_44104,N_43684,N_43507);
and U44105 (N_44105,N_43677,N_43962);
and U44106 (N_44106,N_43516,N_43948);
and U44107 (N_44107,N_43715,N_43927);
xnor U44108 (N_44108,N_43857,N_43530);
nor U44109 (N_44109,N_43899,N_43854);
and U44110 (N_44110,N_43951,N_43930);
nand U44111 (N_44111,N_43806,N_43666);
and U44112 (N_44112,N_43726,N_43986);
and U44113 (N_44113,N_43635,N_43675);
and U44114 (N_44114,N_43755,N_43639);
nor U44115 (N_44115,N_43826,N_43800);
or U44116 (N_44116,N_43864,N_43520);
or U44117 (N_44117,N_43572,N_43770);
or U44118 (N_44118,N_43769,N_43743);
or U44119 (N_44119,N_43959,N_43573);
xor U44120 (N_44120,N_43656,N_43508);
xnor U44121 (N_44121,N_43546,N_43613);
xnor U44122 (N_44122,N_43621,N_43937);
nor U44123 (N_44123,N_43600,N_43917);
or U44124 (N_44124,N_43548,N_43895);
or U44125 (N_44125,N_43746,N_43915);
nand U44126 (N_44126,N_43837,N_43714);
and U44127 (N_44127,N_43821,N_43570);
xnor U44128 (N_44128,N_43649,N_43999);
xor U44129 (N_44129,N_43877,N_43812);
nor U44130 (N_44130,N_43597,N_43749);
xor U44131 (N_44131,N_43884,N_43878);
nor U44132 (N_44132,N_43531,N_43562);
nor U44133 (N_44133,N_43929,N_43876);
nor U44134 (N_44134,N_43880,N_43558);
and U44135 (N_44135,N_43931,N_43810);
nor U44136 (N_44136,N_43945,N_43522);
nor U44137 (N_44137,N_43808,N_43841);
nand U44138 (N_44138,N_43967,N_43627);
or U44139 (N_44139,N_43881,N_43708);
or U44140 (N_44140,N_43737,N_43998);
xor U44141 (N_44141,N_43615,N_43738);
xor U44142 (N_44142,N_43607,N_43754);
or U44143 (N_44143,N_43610,N_43620);
and U44144 (N_44144,N_43883,N_43953);
or U44145 (N_44145,N_43534,N_43707);
nand U44146 (N_44146,N_43842,N_43538);
or U44147 (N_44147,N_43971,N_43705);
nor U44148 (N_44148,N_43803,N_43594);
and U44149 (N_44149,N_43695,N_43887);
nand U44150 (N_44150,N_43747,N_43580);
xnor U44151 (N_44151,N_43688,N_43611);
nand U44152 (N_44152,N_43652,N_43550);
and U44153 (N_44153,N_43868,N_43721);
nand U44154 (N_44154,N_43955,N_43907);
nand U44155 (N_44155,N_43691,N_43788);
xnor U44156 (N_44156,N_43529,N_43525);
or U44157 (N_44157,N_43568,N_43993);
and U44158 (N_44158,N_43760,N_43629);
and U44159 (N_44159,N_43628,N_43593);
or U44160 (N_44160,N_43509,N_43694);
nor U44161 (N_44161,N_43587,N_43569);
nor U44162 (N_44162,N_43551,N_43850);
nor U44163 (N_44163,N_43504,N_43586);
nand U44164 (N_44164,N_43759,N_43686);
xnor U44165 (N_44165,N_43543,N_43544);
xor U44166 (N_44166,N_43882,N_43674);
nand U44167 (N_44167,N_43782,N_43575);
or U44168 (N_44168,N_43809,N_43766);
or U44169 (N_44169,N_43972,N_43552);
and U44170 (N_44170,N_43733,N_43644);
and U44171 (N_44171,N_43902,N_43618);
xnor U44172 (N_44172,N_43592,N_43818);
nand U44173 (N_44173,N_43599,N_43958);
nor U44174 (N_44174,N_43861,N_43792);
nand U44175 (N_44175,N_43710,N_43815);
nor U44176 (N_44176,N_43512,N_43778);
nand U44177 (N_44177,N_43897,N_43697);
nand U44178 (N_44178,N_43503,N_43867);
nor U44179 (N_44179,N_43723,N_43641);
and U44180 (N_44180,N_43780,N_43811);
nand U44181 (N_44181,N_43976,N_43713);
nand U44182 (N_44182,N_43725,N_43893);
nand U44183 (N_44183,N_43973,N_43632);
nand U44184 (N_44184,N_43874,N_43603);
nor U44185 (N_44185,N_43926,N_43685);
and U44186 (N_44186,N_43692,N_43922);
or U44187 (N_44187,N_43923,N_43799);
or U44188 (N_44188,N_43928,N_43515);
nor U44189 (N_44189,N_43924,N_43904);
nor U44190 (N_44190,N_43783,N_43638);
nor U44191 (N_44191,N_43925,N_43941);
xor U44192 (N_44192,N_43911,N_43813);
or U44193 (N_44193,N_43664,N_43977);
or U44194 (N_44194,N_43961,N_43527);
nor U44195 (N_44195,N_43836,N_43647);
nand U44196 (N_44196,N_43995,N_43870);
xor U44197 (N_44197,N_43987,N_43889);
and U44198 (N_44198,N_43831,N_43849);
nand U44199 (N_44199,N_43968,N_43681);
nand U44200 (N_44200,N_43848,N_43651);
and U44201 (N_44201,N_43750,N_43549);
or U44202 (N_44202,N_43518,N_43825);
and U44203 (N_44203,N_43609,N_43822);
xnor U44204 (N_44204,N_43612,N_43942);
nor U44205 (N_44205,N_43960,N_43772);
nor U44206 (N_44206,N_43678,N_43559);
or U44207 (N_44207,N_43919,N_43626);
xnor U44208 (N_44208,N_43879,N_43847);
and U44209 (N_44209,N_43643,N_43557);
or U44210 (N_44210,N_43637,N_43785);
or U44211 (N_44211,N_43853,N_43581);
and U44212 (N_44212,N_43804,N_43744);
nand U44213 (N_44213,N_43517,N_43974);
xor U44214 (N_44214,N_43992,N_43596);
and U44215 (N_44215,N_43789,N_43862);
or U44216 (N_44216,N_43510,N_43795);
xor U44217 (N_44217,N_43939,N_43642);
nor U44218 (N_44218,N_43819,N_43669);
xor U44219 (N_44219,N_43732,N_43771);
nor U44220 (N_44220,N_43585,N_43890);
xor U44221 (N_44221,N_43619,N_43817);
and U44222 (N_44222,N_43910,N_43943);
and U44223 (N_44223,N_43578,N_43665);
and U44224 (N_44224,N_43908,N_43571);
nand U44225 (N_44225,N_43624,N_43689);
and U44226 (N_44226,N_43920,N_43532);
nand U44227 (N_44227,N_43913,N_43735);
and U44228 (N_44228,N_43786,N_43797);
nor U44229 (N_44229,N_43672,N_43663);
nor U44230 (N_44230,N_43561,N_43535);
or U44231 (N_44231,N_43875,N_43693);
and U44232 (N_44232,N_43588,N_43700);
xor U44233 (N_44233,N_43856,N_43646);
nand U44234 (N_44234,N_43952,N_43556);
nor U44235 (N_44235,N_43768,N_43519);
and U44236 (N_44236,N_43984,N_43589);
xnor U44237 (N_44237,N_43865,N_43739);
and U44238 (N_44238,N_43838,N_43645);
or U44239 (N_44239,N_43704,N_43916);
xnor U44240 (N_44240,N_43829,N_43954);
nand U44241 (N_44241,N_43796,N_43514);
xor U44242 (N_44242,N_43542,N_43513);
nand U44243 (N_44243,N_43852,N_43528);
xor U44244 (N_44244,N_43701,N_43981);
or U44245 (N_44245,N_43668,N_43654);
or U44246 (N_44246,N_43787,N_43835);
and U44247 (N_44247,N_43601,N_43832);
or U44248 (N_44248,N_43777,N_43978);
nand U44249 (N_44249,N_43523,N_43728);
and U44250 (N_44250,N_43648,N_43861);
nor U44251 (N_44251,N_43735,N_43616);
xor U44252 (N_44252,N_43854,N_43550);
nand U44253 (N_44253,N_43525,N_43996);
nand U44254 (N_44254,N_43586,N_43949);
nor U44255 (N_44255,N_43805,N_43921);
and U44256 (N_44256,N_43657,N_43840);
nor U44257 (N_44257,N_43934,N_43551);
xnor U44258 (N_44258,N_43893,N_43510);
xnor U44259 (N_44259,N_43886,N_43720);
nand U44260 (N_44260,N_43809,N_43612);
or U44261 (N_44261,N_43805,N_43636);
or U44262 (N_44262,N_43719,N_43967);
or U44263 (N_44263,N_43783,N_43704);
and U44264 (N_44264,N_43770,N_43762);
and U44265 (N_44265,N_43813,N_43993);
nor U44266 (N_44266,N_43538,N_43828);
xor U44267 (N_44267,N_43669,N_43586);
nor U44268 (N_44268,N_43591,N_43560);
or U44269 (N_44269,N_43979,N_43919);
and U44270 (N_44270,N_43954,N_43798);
nand U44271 (N_44271,N_43683,N_43809);
xor U44272 (N_44272,N_43948,N_43756);
and U44273 (N_44273,N_43849,N_43629);
and U44274 (N_44274,N_43722,N_43812);
xor U44275 (N_44275,N_43749,N_43564);
and U44276 (N_44276,N_43785,N_43910);
nor U44277 (N_44277,N_43660,N_43723);
nand U44278 (N_44278,N_43649,N_43797);
nand U44279 (N_44279,N_43614,N_43804);
and U44280 (N_44280,N_43573,N_43635);
nand U44281 (N_44281,N_43688,N_43896);
nor U44282 (N_44282,N_43670,N_43989);
and U44283 (N_44283,N_43519,N_43938);
xor U44284 (N_44284,N_43737,N_43667);
nor U44285 (N_44285,N_43935,N_43703);
nand U44286 (N_44286,N_43665,N_43791);
nor U44287 (N_44287,N_43884,N_43918);
xnor U44288 (N_44288,N_43687,N_43678);
xor U44289 (N_44289,N_43571,N_43687);
xnor U44290 (N_44290,N_43854,N_43631);
or U44291 (N_44291,N_43657,N_43613);
or U44292 (N_44292,N_43919,N_43685);
nor U44293 (N_44293,N_43991,N_43509);
xor U44294 (N_44294,N_43616,N_43578);
nand U44295 (N_44295,N_43742,N_43821);
nor U44296 (N_44296,N_43860,N_43976);
xor U44297 (N_44297,N_43758,N_43598);
xor U44298 (N_44298,N_43903,N_43823);
xnor U44299 (N_44299,N_43723,N_43510);
nand U44300 (N_44300,N_43932,N_43889);
nand U44301 (N_44301,N_43528,N_43985);
and U44302 (N_44302,N_43852,N_43764);
and U44303 (N_44303,N_43962,N_43803);
xor U44304 (N_44304,N_43545,N_43756);
and U44305 (N_44305,N_43695,N_43501);
nand U44306 (N_44306,N_43692,N_43981);
or U44307 (N_44307,N_43977,N_43811);
and U44308 (N_44308,N_43508,N_43993);
nand U44309 (N_44309,N_43953,N_43859);
nand U44310 (N_44310,N_43907,N_43868);
or U44311 (N_44311,N_43990,N_43710);
xnor U44312 (N_44312,N_43811,N_43529);
nand U44313 (N_44313,N_43757,N_43557);
or U44314 (N_44314,N_43738,N_43906);
xor U44315 (N_44315,N_43965,N_43892);
nand U44316 (N_44316,N_43545,N_43955);
xnor U44317 (N_44317,N_43796,N_43620);
and U44318 (N_44318,N_43578,N_43776);
nor U44319 (N_44319,N_43714,N_43589);
nor U44320 (N_44320,N_43521,N_43567);
xnor U44321 (N_44321,N_43894,N_43524);
nand U44322 (N_44322,N_43560,N_43948);
and U44323 (N_44323,N_43754,N_43843);
or U44324 (N_44324,N_43884,N_43721);
nand U44325 (N_44325,N_43612,N_43772);
and U44326 (N_44326,N_43672,N_43994);
nor U44327 (N_44327,N_43806,N_43514);
and U44328 (N_44328,N_43665,N_43559);
nor U44329 (N_44329,N_43681,N_43827);
nor U44330 (N_44330,N_43595,N_43727);
nand U44331 (N_44331,N_43726,N_43704);
xnor U44332 (N_44332,N_43562,N_43658);
and U44333 (N_44333,N_43764,N_43688);
and U44334 (N_44334,N_43760,N_43611);
nor U44335 (N_44335,N_43958,N_43779);
and U44336 (N_44336,N_43789,N_43637);
xor U44337 (N_44337,N_43729,N_43906);
xor U44338 (N_44338,N_43500,N_43792);
or U44339 (N_44339,N_43520,N_43892);
nor U44340 (N_44340,N_43555,N_43891);
nor U44341 (N_44341,N_43906,N_43946);
nand U44342 (N_44342,N_43524,N_43715);
and U44343 (N_44343,N_43871,N_43677);
nor U44344 (N_44344,N_43784,N_43702);
and U44345 (N_44345,N_43812,N_43691);
nand U44346 (N_44346,N_43649,N_43885);
and U44347 (N_44347,N_43950,N_43802);
or U44348 (N_44348,N_43511,N_43957);
nor U44349 (N_44349,N_43770,N_43740);
xnor U44350 (N_44350,N_43637,N_43623);
nor U44351 (N_44351,N_43558,N_43513);
xnor U44352 (N_44352,N_43929,N_43918);
nor U44353 (N_44353,N_43555,N_43582);
or U44354 (N_44354,N_43740,N_43662);
nand U44355 (N_44355,N_43732,N_43951);
nor U44356 (N_44356,N_43955,N_43620);
or U44357 (N_44357,N_43610,N_43558);
xor U44358 (N_44358,N_43804,N_43928);
nor U44359 (N_44359,N_43723,N_43711);
and U44360 (N_44360,N_43733,N_43858);
nor U44361 (N_44361,N_43976,N_43876);
and U44362 (N_44362,N_43769,N_43942);
nor U44363 (N_44363,N_43678,N_43686);
or U44364 (N_44364,N_43739,N_43593);
or U44365 (N_44365,N_43563,N_43645);
and U44366 (N_44366,N_43811,N_43691);
nand U44367 (N_44367,N_43957,N_43865);
nand U44368 (N_44368,N_43658,N_43593);
or U44369 (N_44369,N_43953,N_43991);
nand U44370 (N_44370,N_43962,N_43814);
and U44371 (N_44371,N_43649,N_43975);
xnor U44372 (N_44372,N_43503,N_43881);
or U44373 (N_44373,N_43703,N_43811);
or U44374 (N_44374,N_43711,N_43714);
nand U44375 (N_44375,N_43733,N_43586);
and U44376 (N_44376,N_43931,N_43910);
xnor U44377 (N_44377,N_43996,N_43988);
and U44378 (N_44378,N_43548,N_43847);
xnor U44379 (N_44379,N_43931,N_43580);
or U44380 (N_44380,N_43627,N_43757);
xnor U44381 (N_44381,N_43737,N_43647);
nand U44382 (N_44382,N_43824,N_43899);
nor U44383 (N_44383,N_43954,N_43542);
xor U44384 (N_44384,N_43635,N_43909);
and U44385 (N_44385,N_43981,N_43802);
xor U44386 (N_44386,N_43851,N_43623);
and U44387 (N_44387,N_43852,N_43582);
or U44388 (N_44388,N_43838,N_43965);
or U44389 (N_44389,N_43765,N_43897);
nand U44390 (N_44390,N_43952,N_43724);
nand U44391 (N_44391,N_43635,N_43696);
or U44392 (N_44392,N_43991,N_43861);
and U44393 (N_44393,N_43948,N_43795);
and U44394 (N_44394,N_43743,N_43741);
nand U44395 (N_44395,N_43719,N_43807);
nand U44396 (N_44396,N_43620,N_43656);
nor U44397 (N_44397,N_43546,N_43879);
xnor U44398 (N_44398,N_43828,N_43720);
nand U44399 (N_44399,N_43525,N_43903);
and U44400 (N_44400,N_43518,N_43745);
and U44401 (N_44401,N_43500,N_43959);
xor U44402 (N_44402,N_43989,N_43736);
xor U44403 (N_44403,N_43563,N_43555);
or U44404 (N_44404,N_43829,N_43791);
xnor U44405 (N_44405,N_43761,N_43554);
xnor U44406 (N_44406,N_43738,N_43843);
and U44407 (N_44407,N_43808,N_43562);
or U44408 (N_44408,N_43530,N_43550);
or U44409 (N_44409,N_43625,N_43759);
or U44410 (N_44410,N_43869,N_43815);
nand U44411 (N_44411,N_43972,N_43587);
or U44412 (N_44412,N_43840,N_43888);
nand U44413 (N_44413,N_43937,N_43811);
xor U44414 (N_44414,N_43533,N_43579);
and U44415 (N_44415,N_43553,N_43708);
xor U44416 (N_44416,N_43769,N_43618);
nand U44417 (N_44417,N_43956,N_43553);
nor U44418 (N_44418,N_43783,N_43790);
nor U44419 (N_44419,N_43958,N_43895);
and U44420 (N_44420,N_43652,N_43986);
or U44421 (N_44421,N_43991,N_43694);
xnor U44422 (N_44422,N_43688,N_43815);
and U44423 (N_44423,N_43999,N_43781);
nand U44424 (N_44424,N_43874,N_43624);
nand U44425 (N_44425,N_43894,N_43695);
nor U44426 (N_44426,N_43655,N_43889);
or U44427 (N_44427,N_43877,N_43870);
xnor U44428 (N_44428,N_43576,N_43661);
or U44429 (N_44429,N_43982,N_43927);
or U44430 (N_44430,N_43860,N_43717);
and U44431 (N_44431,N_43798,N_43946);
nor U44432 (N_44432,N_43689,N_43701);
or U44433 (N_44433,N_43801,N_43653);
nand U44434 (N_44434,N_43894,N_43866);
nand U44435 (N_44435,N_43744,N_43905);
nand U44436 (N_44436,N_43796,N_43917);
and U44437 (N_44437,N_43814,N_43853);
nand U44438 (N_44438,N_43682,N_43847);
or U44439 (N_44439,N_43652,N_43647);
xnor U44440 (N_44440,N_43723,N_43939);
nor U44441 (N_44441,N_43615,N_43803);
xor U44442 (N_44442,N_43569,N_43671);
nor U44443 (N_44443,N_43754,N_43870);
nand U44444 (N_44444,N_43769,N_43549);
nand U44445 (N_44445,N_43747,N_43943);
and U44446 (N_44446,N_43984,N_43668);
and U44447 (N_44447,N_43912,N_43577);
xnor U44448 (N_44448,N_43906,N_43766);
xnor U44449 (N_44449,N_43681,N_43698);
xor U44450 (N_44450,N_43658,N_43856);
and U44451 (N_44451,N_43588,N_43676);
xnor U44452 (N_44452,N_43892,N_43605);
nor U44453 (N_44453,N_43758,N_43636);
or U44454 (N_44454,N_43768,N_43791);
xnor U44455 (N_44455,N_43840,N_43544);
and U44456 (N_44456,N_43753,N_43609);
or U44457 (N_44457,N_43523,N_43755);
and U44458 (N_44458,N_43947,N_43701);
and U44459 (N_44459,N_43664,N_43781);
xnor U44460 (N_44460,N_43734,N_43965);
and U44461 (N_44461,N_43845,N_43770);
nor U44462 (N_44462,N_43767,N_43979);
or U44463 (N_44463,N_43832,N_43793);
nand U44464 (N_44464,N_43630,N_43660);
xor U44465 (N_44465,N_43815,N_43516);
xor U44466 (N_44466,N_43898,N_43835);
nand U44467 (N_44467,N_43512,N_43949);
xnor U44468 (N_44468,N_43539,N_43550);
nand U44469 (N_44469,N_43772,N_43827);
nand U44470 (N_44470,N_43820,N_43910);
nand U44471 (N_44471,N_43511,N_43960);
and U44472 (N_44472,N_43689,N_43752);
nor U44473 (N_44473,N_43687,N_43815);
nor U44474 (N_44474,N_43598,N_43961);
xnor U44475 (N_44475,N_43796,N_43671);
xnor U44476 (N_44476,N_43990,N_43501);
xor U44477 (N_44477,N_43940,N_43575);
nor U44478 (N_44478,N_43663,N_43860);
nor U44479 (N_44479,N_43898,N_43639);
nand U44480 (N_44480,N_43656,N_43948);
and U44481 (N_44481,N_43553,N_43567);
xnor U44482 (N_44482,N_43905,N_43947);
xor U44483 (N_44483,N_43912,N_43631);
xnor U44484 (N_44484,N_43913,N_43905);
nand U44485 (N_44485,N_43537,N_43990);
and U44486 (N_44486,N_43753,N_43848);
nor U44487 (N_44487,N_43626,N_43928);
nand U44488 (N_44488,N_43895,N_43781);
xor U44489 (N_44489,N_43668,N_43710);
nand U44490 (N_44490,N_43844,N_43799);
or U44491 (N_44491,N_43725,N_43655);
nand U44492 (N_44492,N_43718,N_43542);
xor U44493 (N_44493,N_43614,N_43833);
xnor U44494 (N_44494,N_43673,N_43862);
nor U44495 (N_44495,N_43937,N_43538);
xnor U44496 (N_44496,N_43646,N_43966);
xnor U44497 (N_44497,N_43837,N_43740);
xnor U44498 (N_44498,N_43710,N_43564);
and U44499 (N_44499,N_43933,N_43794);
nand U44500 (N_44500,N_44215,N_44316);
nand U44501 (N_44501,N_44112,N_44005);
nand U44502 (N_44502,N_44206,N_44450);
nor U44503 (N_44503,N_44198,N_44442);
or U44504 (N_44504,N_44460,N_44083);
or U44505 (N_44505,N_44169,N_44261);
or U44506 (N_44506,N_44413,N_44447);
and U44507 (N_44507,N_44201,N_44362);
or U44508 (N_44508,N_44392,N_44411);
and U44509 (N_44509,N_44283,N_44243);
and U44510 (N_44510,N_44485,N_44221);
xnor U44511 (N_44511,N_44276,N_44330);
nand U44512 (N_44512,N_44191,N_44388);
and U44513 (N_44513,N_44098,N_44094);
and U44514 (N_44514,N_44246,N_44019);
nor U44515 (N_44515,N_44279,N_44224);
and U44516 (N_44516,N_44126,N_44158);
xor U44517 (N_44517,N_44018,N_44202);
nor U44518 (N_44518,N_44376,N_44285);
and U44519 (N_44519,N_44227,N_44280);
nand U44520 (N_44520,N_44284,N_44179);
nor U44521 (N_44521,N_44311,N_44327);
or U44522 (N_44522,N_44162,N_44070);
and U44523 (N_44523,N_44475,N_44410);
or U44524 (N_44524,N_44080,N_44183);
nor U44525 (N_44525,N_44434,N_44248);
and U44526 (N_44526,N_44455,N_44312);
and U44527 (N_44527,N_44136,N_44291);
xor U44528 (N_44528,N_44104,N_44043);
or U44529 (N_44529,N_44372,N_44457);
and U44530 (N_44530,N_44218,N_44121);
or U44531 (N_44531,N_44028,N_44433);
and U44532 (N_44532,N_44289,N_44012);
nor U44533 (N_44533,N_44440,N_44030);
xor U44534 (N_44534,N_44190,N_44439);
nor U44535 (N_44535,N_44443,N_44099);
nand U44536 (N_44536,N_44247,N_44383);
nand U44537 (N_44537,N_44303,N_44236);
xnor U44538 (N_44538,N_44421,N_44103);
and U44539 (N_44539,N_44220,N_44431);
nor U44540 (N_44540,N_44301,N_44459);
and U44541 (N_44541,N_44233,N_44346);
nor U44542 (N_44542,N_44398,N_44016);
nand U44543 (N_44543,N_44196,N_44319);
xnor U44544 (N_44544,N_44155,N_44110);
nor U44545 (N_44545,N_44156,N_44370);
xor U44546 (N_44546,N_44125,N_44085);
or U44547 (N_44547,N_44051,N_44356);
or U44548 (N_44548,N_44483,N_44002);
xor U44549 (N_44549,N_44288,N_44037);
nand U44550 (N_44550,N_44174,N_44153);
xor U44551 (N_44551,N_44195,N_44258);
nand U44552 (N_44552,N_44160,N_44453);
nor U44553 (N_44553,N_44046,N_44393);
or U44554 (N_44554,N_44142,N_44444);
nand U44555 (N_44555,N_44122,N_44368);
or U44556 (N_44556,N_44058,N_44355);
nand U44557 (N_44557,N_44401,N_44203);
nand U44558 (N_44558,N_44467,N_44360);
nand U44559 (N_44559,N_44363,N_44095);
nand U44560 (N_44560,N_44304,N_44000);
xor U44561 (N_44561,N_44272,N_44417);
nor U44562 (N_44562,N_44014,N_44065);
xor U44563 (N_44563,N_44409,N_44146);
or U44564 (N_44564,N_44254,N_44415);
and U44565 (N_44565,N_44396,N_44296);
xor U44566 (N_44566,N_44208,N_44449);
nand U44567 (N_44567,N_44349,N_44143);
nand U44568 (N_44568,N_44205,N_44499);
xnor U44569 (N_44569,N_44265,N_44302);
or U44570 (N_44570,N_44177,N_44337);
or U44571 (N_44571,N_44259,N_44317);
and U44572 (N_44572,N_44150,N_44361);
nand U44573 (N_44573,N_44050,N_44386);
xnor U44574 (N_44574,N_44022,N_44130);
nand U44575 (N_44575,N_44322,N_44029);
nand U44576 (N_44576,N_44239,N_44400);
or U44577 (N_44577,N_44192,N_44141);
or U44578 (N_44578,N_44364,N_44397);
or U44579 (N_44579,N_44482,N_44152);
nand U44580 (N_44580,N_44222,N_44277);
nor U44581 (N_44581,N_44039,N_44036);
nand U44582 (N_44582,N_44340,N_44270);
nor U44583 (N_44583,N_44041,N_44448);
and U44584 (N_44584,N_44424,N_44314);
nand U44585 (N_44585,N_44154,N_44127);
or U44586 (N_44586,N_44225,N_44318);
or U44587 (N_44587,N_44348,N_44049);
and U44588 (N_44588,N_44033,N_44034);
or U44589 (N_44589,N_44105,N_44017);
nor U44590 (N_44590,N_44427,N_44230);
and U44591 (N_44591,N_44486,N_44406);
nand U44592 (N_44592,N_44040,N_44306);
nand U44593 (N_44593,N_44266,N_44101);
or U44594 (N_44594,N_44114,N_44297);
nand U44595 (N_44595,N_44463,N_44075);
xnor U44596 (N_44596,N_44476,N_44235);
and U44597 (N_44597,N_44387,N_44445);
nor U44598 (N_44598,N_44088,N_44271);
nor U44599 (N_44599,N_44001,N_44117);
nor U44600 (N_44600,N_44176,N_44458);
nor U44601 (N_44601,N_44059,N_44377);
xnor U44602 (N_44602,N_44256,N_44015);
nand U44603 (N_44603,N_44347,N_44237);
nor U44604 (N_44604,N_44074,N_44404);
nor U44605 (N_44605,N_44321,N_44045);
or U44606 (N_44606,N_44328,N_44009);
nand U44607 (N_44607,N_44374,N_44473);
xnor U44608 (N_44608,N_44140,N_44358);
nor U44609 (N_44609,N_44339,N_44062);
or U44610 (N_44610,N_44468,N_44175);
nor U44611 (N_44611,N_44269,N_44390);
nand U44612 (N_44612,N_44129,N_44123);
and U44613 (N_44613,N_44484,N_44255);
or U44614 (N_44614,N_44441,N_44275);
nor U44615 (N_44615,N_44294,N_44164);
and U44616 (N_44616,N_44054,N_44004);
nand U44617 (N_44617,N_44428,N_44477);
or U44618 (N_44618,N_44278,N_44373);
nand U44619 (N_44619,N_44166,N_44325);
and U44620 (N_44620,N_44038,N_44011);
nor U44621 (N_44621,N_44429,N_44023);
nand U44622 (N_44622,N_44371,N_44207);
and U44623 (N_44623,N_44490,N_44232);
and U44624 (N_44624,N_44170,N_44096);
nand U44625 (N_44625,N_44064,N_44055);
nor U44626 (N_44626,N_44488,N_44214);
nor U44627 (N_44627,N_44188,N_44335);
or U44628 (N_44628,N_44326,N_44056);
and U44629 (N_44629,N_44430,N_44133);
xnor U44630 (N_44630,N_44182,N_44305);
and U44631 (N_44631,N_44134,N_44149);
xor U44632 (N_44632,N_44086,N_44008);
nand U44633 (N_44633,N_44384,N_44031);
xnor U44634 (N_44634,N_44006,N_44353);
and U44635 (N_44635,N_44115,N_44210);
or U44636 (N_44636,N_44437,N_44298);
and U44637 (N_44637,N_44226,N_44189);
nand U44638 (N_44638,N_44240,N_44229);
and U44639 (N_44639,N_44389,N_44111);
nor U44640 (N_44640,N_44481,N_44242);
and U44641 (N_44641,N_44184,N_44422);
xnor U44642 (N_44642,N_44351,N_44307);
nor U44643 (N_44643,N_44426,N_44492);
nand U44644 (N_44644,N_44217,N_44352);
nor U44645 (N_44645,N_44412,N_44167);
and U44646 (N_44646,N_44241,N_44451);
and U44647 (N_44647,N_44109,N_44081);
xor U44648 (N_44648,N_44161,N_44379);
nor U44649 (N_44649,N_44071,N_44472);
nand U44650 (N_44650,N_44234,N_44309);
nand U44651 (N_44651,N_44021,N_44200);
nor U44652 (N_44652,N_44308,N_44178);
and U44653 (N_44653,N_44165,N_44252);
xor U44654 (N_44654,N_44181,N_44432);
or U44655 (N_44655,N_44102,N_44343);
nor U44656 (N_44656,N_44090,N_44257);
xor U44657 (N_44657,N_44456,N_44382);
and U44658 (N_44658,N_44197,N_44106);
and U44659 (N_44659,N_44375,N_44454);
xor U44660 (N_44660,N_44338,N_44128);
and U44661 (N_44661,N_44497,N_44171);
xor U44662 (N_44662,N_44498,N_44478);
nand U44663 (N_44663,N_44173,N_44027);
nor U44664 (N_44664,N_44491,N_44342);
nand U44665 (N_44665,N_44333,N_44107);
nand U44666 (N_44666,N_44186,N_44391);
and U44667 (N_44667,N_44300,N_44151);
nor U44668 (N_44668,N_44407,N_44359);
or U44669 (N_44669,N_44344,N_44135);
and U44670 (N_44670,N_44209,N_44394);
nor U44671 (N_44671,N_44087,N_44323);
nand U44672 (N_44672,N_44244,N_44097);
nand U44673 (N_44673,N_44079,N_44299);
nor U44674 (N_44674,N_44470,N_44395);
or U44675 (N_44675,N_44494,N_44320);
and U44676 (N_44676,N_44466,N_44489);
or U44677 (N_44677,N_44365,N_44063);
or U44678 (N_44678,N_44120,N_44060);
and U44679 (N_44679,N_44007,N_44053);
nor U44680 (N_44680,N_44025,N_44003);
nor U44681 (N_44681,N_44047,N_44245);
xnor U44682 (N_44682,N_44223,N_44436);
and U44683 (N_44683,N_44496,N_44493);
nand U44684 (N_44684,N_44035,N_44157);
nor U44685 (N_44685,N_44471,N_44148);
nand U44686 (N_44686,N_44066,N_44290);
or U44687 (N_44687,N_44249,N_44403);
or U44688 (N_44688,N_44211,N_44461);
and U44689 (N_44689,N_44313,N_44100);
nand U44690 (N_44690,N_44267,N_44274);
or U44691 (N_44691,N_44089,N_44042);
nand U44692 (N_44692,N_44180,N_44119);
nor U44693 (N_44693,N_44465,N_44334);
and U44694 (N_44694,N_44350,N_44078);
xnor U44695 (N_44695,N_44048,N_44052);
and U44696 (N_44696,N_44452,N_44228);
and U44697 (N_44697,N_44420,N_44260);
or U44698 (N_44698,N_44113,N_44138);
or U44699 (N_44699,N_44385,N_44399);
xnor U44700 (N_44700,N_44282,N_44324);
or U44701 (N_44701,N_44076,N_44010);
nor U44702 (N_44702,N_44108,N_44073);
nor U44703 (N_44703,N_44067,N_44462);
and U44704 (N_44704,N_44116,N_44144);
xnor U44705 (N_44705,N_44057,N_44366);
and U44706 (N_44706,N_44032,N_44072);
and U44707 (N_44707,N_44212,N_44163);
nor U44708 (N_44708,N_44213,N_44013);
xnor U44709 (N_44709,N_44118,N_44131);
nand U44710 (N_44710,N_44286,N_44268);
nor U44711 (N_44711,N_44281,N_44124);
xor U44712 (N_44712,N_44238,N_44438);
and U44713 (N_44713,N_44077,N_44367);
or U44714 (N_44714,N_44378,N_44341);
nor U44715 (N_44715,N_44369,N_44480);
nor U44716 (N_44716,N_44159,N_44145);
nand U44717 (N_44717,N_44474,N_44068);
and U44718 (N_44718,N_44147,N_44357);
nor U44719 (N_44719,N_44435,N_44292);
or U44720 (N_44720,N_44139,N_44310);
or U44721 (N_44721,N_44345,N_44380);
or U44722 (N_44722,N_44381,N_44293);
and U44723 (N_44723,N_44329,N_44199);
nor U44724 (N_44724,N_44082,N_44219);
and U44725 (N_44725,N_44332,N_44061);
xor U44726 (N_44726,N_44250,N_44020);
xnor U44727 (N_44727,N_44418,N_44044);
or U44728 (N_44728,N_44425,N_44168);
nand U44729 (N_44729,N_44423,N_44414);
nand U44730 (N_44730,N_44287,N_44092);
xnor U44731 (N_44731,N_44253,N_44419);
nor U44732 (N_44732,N_44331,N_44132);
xor U44733 (N_44733,N_44024,N_44185);
and U44734 (N_44734,N_44172,N_44263);
xor U44735 (N_44735,N_44495,N_44408);
nand U44736 (N_44736,N_44193,N_44137);
and U44737 (N_44737,N_44402,N_44446);
or U44738 (N_44738,N_44416,N_44273);
xor U44739 (N_44739,N_44487,N_44336);
nand U44740 (N_44740,N_44405,N_44479);
or U44741 (N_44741,N_44069,N_44295);
or U44742 (N_44742,N_44026,N_44469);
nand U44743 (N_44743,N_44354,N_44204);
or U44744 (N_44744,N_44216,N_44093);
and U44745 (N_44745,N_44264,N_44464);
nor U44746 (N_44746,N_44231,N_44315);
nor U44747 (N_44747,N_44251,N_44084);
xor U44748 (N_44748,N_44262,N_44194);
xnor U44749 (N_44749,N_44091,N_44187);
xnor U44750 (N_44750,N_44199,N_44438);
nand U44751 (N_44751,N_44007,N_44454);
or U44752 (N_44752,N_44367,N_44133);
xnor U44753 (N_44753,N_44211,N_44186);
xnor U44754 (N_44754,N_44047,N_44253);
or U44755 (N_44755,N_44373,N_44168);
and U44756 (N_44756,N_44044,N_44174);
and U44757 (N_44757,N_44061,N_44168);
xor U44758 (N_44758,N_44490,N_44298);
and U44759 (N_44759,N_44161,N_44166);
nand U44760 (N_44760,N_44080,N_44015);
nor U44761 (N_44761,N_44411,N_44187);
nor U44762 (N_44762,N_44337,N_44422);
nand U44763 (N_44763,N_44317,N_44001);
nor U44764 (N_44764,N_44439,N_44322);
nand U44765 (N_44765,N_44490,N_44218);
nor U44766 (N_44766,N_44289,N_44393);
nand U44767 (N_44767,N_44479,N_44023);
nand U44768 (N_44768,N_44108,N_44241);
xnor U44769 (N_44769,N_44404,N_44152);
xnor U44770 (N_44770,N_44004,N_44277);
and U44771 (N_44771,N_44232,N_44215);
or U44772 (N_44772,N_44075,N_44092);
xor U44773 (N_44773,N_44452,N_44266);
nand U44774 (N_44774,N_44355,N_44048);
nor U44775 (N_44775,N_44102,N_44130);
nand U44776 (N_44776,N_44304,N_44013);
or U44777 (N_44777,N_44160,N_44055);
xnor U44778 (N_44778,N_44461,N_44206);
and U44779 (N_44779,N_44331,N_44109);
or U44780 (N_44780,N_44048,N_44466);
xnor U44781 (N_44781,N_44497,N_44117);
nor U44782 (N_44782,N_44327,N_44132);
nor U44783 (N_44783,N_44366,N_44183);
nor U44784 (N_44784,N_44447,N_44152);
nor U44785 (N_44785,N_44220,N_44041);
or U44786 (N_44786,N_44211,N_44119);
or U44787 (N_44787,N_44387,N_44413);
and U44788 (N_44788,N_44080,N_44410);
nor U44789 (N_44789,N_44116,N_44369);
and U44790 (N_44790,N_44283,N_44304);
nand U44791 (N_44791,N_44158,N_44373);
or U44792 (N_44792,N_44083,N_44140);
and U44793 (N_44793,N_44211,N_44077);
and U44794 (N_44794,N_44174,N_44047);
nand U44795 (N_44795,N_44433,N_44405);
and U44796 (N_44796,N_44317,N_44463);
or U44797 (N_44797,N_44204,N_44333);
nand U44798 (N_44798,N_44263,N_44226);
or U44799 (N_44799,N_44406,N_44373);
and U44800 (N_44800,N_44361,N_44232);
or U44801 (N_44801,N_44048,N_44366);
or U44802 (N_44802,N_44196,N_44342);
xor U44803 (N_44803,N_44415,N_44272);
nand U44804 (N_44804,N_44214,N_44386);
and U44805 (N_44805,N_44337,N_44401);
nand U44806 (N_44806,N_44218,N_44007);
and U44807 (N_44807,N_44074,N_44418);
or U44808 (N_44808,N_44372,N_44226);
xor U44809 (N_44809,N_44364,N_44112);
nand U44810 (N_44810,N_44371,N_44307);
or U44811 (N_44811,N_44480,N_44436);
nor U44812 (N_44812,N_44024,N_44219);
nor U44813 (N_44813,N_44233,N_44493);
nand U44814 (N_44814,N_44239,N_44302);
or U44815 (N_44815,N_44240,N_44300);
xnor U44816 (N_44816,N_44203,N_44272);
nor U44817 (N_44817,N_44385,N_44254);
nand U44818 (N_44818,N_44280,N_44420);
nand U44819 (N_44819,N_44022,N_44326);
xor U44820 (N_44820,N_44111,N_44255);
or U44821 (N_44821,N_44095,N_44091);
nand U44822 (N_44822,N_44295,N_44119);
and U44823 (N_44823,N_44218,N_44189);
and U44824 (N_44824,N_44475,N_44122);
nor U44825 (N_44825,N_44285,N_44246);
nor U44826 (N_44826,N_44202,N_44489);
and U44827 (N_44827,N_44313,N_44234);
and U44828 (N_44828,N_44342,N_44263);
or U44829 (N_44829,N_44261,N_44383);
nor U44830 (N_44830,N_44140,N_44309);
nor U44831 (N_44831,N_44129,N_44221);
or U44832 (N_44832,N_44442,N_44433);
nor U44833 (N_44833,N_44476,N_44117);
nor U44834 (N_44834,N_44047,N_44156);
nand U44835 (N_44835,N_44227,N_44406);
nor U44836 (N_44836,N_44479,N_44135);
xnor U44837 (N_44837,N_44379,N_44417);
nor U44838 (N_44838,N_44224,N_44271);
nor U44839 (N_44839,N_44297,N_44487);
or U44840 (N_44840,N_44031,N_44214);
nor U44841 (N_44841,N_44064,N_44122);
nand U44842 (N_44842,N_44094,N_44384);
nand U44843 (N_44843,N_44119,N_44168);
nand U44844 (N_44844,N_44462,N_44072);
or U44845 (N_44845,N_44230,N_44117);
and U44846 (N_44846,N_44300,N_44174);
xnor U44847 (N_44847,N_44143,N_44024);
nand U44848 (N_44848,N_44351,N_44002);
or U44849 (N_44849,N_44088,N_44318);
nor U44850 (N_44850,N_44411,N_44017);
nor U44851 (N_44851,N_44350,N_44485);
nor U44852 (N_44852,N_44451,N_44042);
nand U44853 (N_44853,N_44412,N_44068);
nor U44854 (N_44854,N_44258,N_44390);
or U44855 (N_44855,N_44325,N_44416);
or U44856 (N_44856,N_44397,N_44134);
and U44857 (N_44857,N_44439,N_44192);
or U44858 (N_44858,N_44234,N_44495);
and U44859 (N_44859,N_44368,N_44055);
or U44860 (N_44860,N_44311,N_44185);
nand U44861 (N_44861,N_44017,N_44036);
nand U44862 (N_44862,N_44193,N_44146);
xnor U44863 (N_44863,N_44269,N_44098);
nor U44864 (N_44864,N_44099,N_44293);
nand U44865 (N_44865,N_44040,N_44366);
and U44866 (N_44866,N_44130,N_44159);
or U44867 (N_44867,N_44069,N_44297);
and U44868 (N_44868,N_44353,N_44379);
xnor U44869 (N_44869,N_44124,N_44312);
xor U44870 (N_44870,N_44488,N_44109);
nand U44871 (N_44871,N_44032,N_44346);
or U44872 (N_44872,N_44311,N_44049);
xor U44873 (N_44873,N_44151,N_44068);
xnor U44874 (N_44874,N_44309,N_44365);
nand U44875 (N_44875,N_44443,N_44354);
nor U44876 (N_44876,N_44348,N_44149);
nand U44877 (N_44877,N_44182,N_44112);
and U44878 (N_44878,N_44095,N_44307);
or U44879 (N_44879,N_44182,N_44321);
xor U44880 (N_44880,N_44020,N_44182);
xnor U44881 (N_44881,N_44103,N_44284);
nand U44882 (N_44882,N_44367,N_44377);
nor U44883 (N_44883,N_44269,N_44478);
nor U44884 (N_44884,N_44325,N_44192);
nand U44885 (N_44885,N_44388,N_44312);
nor U44886 (N_44886,N_44169,N_44430);
xor U44887 (N_44887,N_44443,N_44496);
nand U44888 (N_44888,N_44292,N_44140);
or U44889 (N_44889,N_44488,N_44203);
or U44890 (N_44890,N_44398,N_44372);
and U44891 (N_44891,N_44329,N_44033);
and U44892 (N_44892,N_44078,N_44409);
nand U44893 (N_44893,N_44096,N_44216);
xor U44894 (N_44894,N_44031,N_44346);
xor U44895 (N_44895,N_44173,N_44024);
and U44896 (N_44896,N_44195,N_44291);
and U44897 (N_44897,N_44037,N_44440);
xnor U44898 (N_44898,N_44325,N_44077);
xor U44899 (N_44899,N_44457,N_44456);
and U44900 (N_44900,N_44440,N_44366);
and U44901 (N_44901,N_44046,N_44492);
xnor U44902 (N_44902,N_44192,N_44026);
nor U44903 (N_44903,N_44296,N_44312);
or U44904 (N_44904,N_44079,N_44246);
or U44905 (N_44905,N_44102,N_44367);
nor U44906 (N_44906,N_44462,N_44061);
xor U44907 (N_44907,N_44052,N_44466);
xnor U44908 (N_44908,N_44090,N_44384);
nor U44909 (N_44909,N_44395,N_44371);
nor U44910 (N_44910,N_44278,N_44053);
and U44911 (N_44911,N_44101,N_44124);
or U44912 (N_44912,N_44002,N_44355);
xnor U44913 (N_44913,N_44472,N_44286);
or U44914 (N_44914,N_44351,N_44250);
and U44915 (N_44915,N_44191,N_44477);
nor U44916 (N_44916,N_44270,N_44115);
xor U44917 (N_44917,N_44404,N_44488);
xnor U44918 (N_44918,N_44471,N_44177);
or U44919 (N_44919,N_44153,N_44191);
and U44920 (N_44920,N_44266,N_44172);
and U44921 (N_44921,N_44178,N_44497);
xor U44922 (N_44922,N_44430,N_44392);
and U44923 (N_44923,N_44162,N_44454);
xnor U44924 (N_44924,N_44497,N_44390);
or U44925 (N_44925,N_44163,N_44471);
nor U44926 (N_44926,N_44117,N_44037);
nand U44927 (N_44927,N_44487,N_44255);
or U44928 (N_44928,N_44203,N_44377);
or U44929 (N_44929,N_44241,N_44354);
xor U44930 (N_44930,N_44426,N_44009);
or U44931 (N_44931,N_44267,N_44229);
nand U44932 (N_44932,N_44331,N_44362);
or U44933 (N_44933,N_44454,N_44118);
nand U44934 (N_44934,N_44038,N_44465);
xor U44935 (N_44935,N_44230,N_44476);
or U44936 (N_44936,N_44183,N_44255);
nor U44937 (N_44937,N_44455,N_44160);
nor U44938 (N_44938,N_44287,N_44356);
and U44939 (N_44939,N_44382,N_44054);
xor U44940 (N_44940,N_44451,N_44424);
nand U44941 (N_44941,N_44270,N_44454);
xnor U44942 (N_44942,N_44263,N_44478);
or U44943 (N_44943,N_44341,N_44482);
or U44944 (N_44944,N_44087,N_44125);
xnor U44945 (N_44945,N_44483,N_44464);
nor U44946 (N_44946,N_44465,N_44238);
xor U44947 (N_44947,N_44380,N_44311);
nor U44948 (N_44948,N_44429,N_44176);
xor U44949 (N_44949,N_44204,N_44021);
and U44950 (N_44950,N_44334,N_44486);
or U44951 (N_44951,N_44085,N_44220);
or U44952 (N_44952,N_44170,N_44029);
nand U44953 (N_44953,N_44060,N_44220);
nand U44954 (N_44954,N_44460,N_44466);
and U44955 (N_44955,N_44212,N_44231);
and U44956 (N_44956,N_44095,N_44249);
nor U44957 (N_44957,N_44253,N_44220);
nand U44958 (N_44958,N_44259,N_44059);
nor U44959 (N_44959,N_44217,N_44317);
nand U44960 (N_44960,N_44175,N_44368);
xor U44961 (N_44961,N_44359,N_44466);
nor U44962 (N_44962,N_44014,N_44016);
or U44963 (N_44963,N_44330,N_44057);
and U44964 (N_44964,N_44181,N_44118);
or U44965 (N_44965,N_44130,N_44454);
and U44966 (N_44966,N_44126,N_44300);
nor U44967 (N_44967,N_44374,N_44036);
xnor U44968 (N_44968,N_44120,N_44000);
nor U44969 (N_44969,N_44430,N_44100);
nor U44970 (N_44970,N_44270,N_44014);
xor U44971 (N_44971,N_44306,N_44003);
or U44972 (N_44972,N_44394,N_44358);
nand U44973 (N_44973,N_44122,N_44200);
xnor U44974 (N_44974,N_44317,N_44080);
and U44975 (N_44975,N_44165,N_44048);
or U44976 (N_44976,N_44025,N_44278);
nor U44977 (N_44977,N_44177,N_44106);
nor U44978 (N_44978,N_44075,N_44318);
and U44979 (N_44979,N_44466,N_44243);
nor U44980 (N_44980,N_44149,N_44265);
or U44981 (N_44981,N_44273,N_44345);
and U44982 (N_44982,N_44386,N_44162);
xor U44983 (N_44983,N_44247,N_44285);
xnor U44984 (N_44984,N_44258,N_44467);
nor U44985 (N_44985,N_44389,N_44374);
or U44986 (N_44986,N_44074,N_44496);
or U44987 (N_44987,N_44060,N_44410);
and U44988 (N_44988,N_44432,N_44062);
and U44989 (N_44989,N_44269,N_44155);
nand U44990 (N_44990,N_44399,N_44395);
or U44991 (N_44991,N_44005,N_44386);
nand U44992 (N_44992,N_44439,N_44407);
or U44993 (N_44993,N_44133,N_44057);
nand U44994 (N_44994,N_44193,N_44143);
xor U44995 (N_44995,N_44364,N_44357);
and U44996 (N_44996,N_44410,N_44008);
nand U44997 (N_44997,N_44404,N_44287);
and U44998 (N_44998,N_44441,N_44115);
and U44999 (N_44999,N_44486,N_44246);
or U45000 (N_45000,N_44673,N_44820);
and U45001 (N_45001,N_44906,N_44876);
nor U45002 (N_45002,N_44525,N_44654);
nand U45003 (N_45003,N_44921,N_44635);
nor U45004 (N_45004,N_44824,N_44701);
xor U45005 (N_45005,N_44903,N_44968);
or U45006 (N_45006,N_44777,N_44993);
nor U45007 (N_45007,N_44848,N_44996);
xnor U45008 (N_45008,N_44947,N_44704);
nand U45009 (N_45009,N_44856,N_44956);
nor U45010 (N_45010,N_44928,N_44513);
xor U45011 (N_45011,N_44564,N_44606);
xnor U45012 (N_45012,N_44748,N_44678);
and U45013 (N_45013,N_44573,N_44730);
xor U45014 (N_45014,N_44534,N_44512);
xor U45015 (N_45015,N_44645,N_44822);
nor U45016 (N_45016,N_44954,N_44516);
nor U45017 (N_45017,N_44842,N_44631);
nor U45018 (N_45018,N_44858,N_44891);
nand U45019 (N_45019,N_44924,N_44682);
nor U45020 (N_45020,N_44557,N_44549);
nor U45021 (N_45021,N_44752,N_44505);
or U45022 (N_45022,N_44640,N_44849);
xnor U45023 (N_45023,N_44980,N_44530);
nor U45024 (N_45024,N_44655,N_44625);
or U45025 (N_45025,N_44901,N_44543);
and U45026 (N_45026,N_44818,N_44642);
xnor U45027 (N_45027,N_44694,N_44997);
xnor U45028 (N_45028,N_44602,N_44857);
nor U45029 (N_45029,N_44548,N_44617);
and U45030 (N_45030,N_44584,N_44605);
or U45031 (N_45031,N_44755,N_44560);
nand U45032 (N_45032,N_44799,N_44869);
or U45033 (N_45033,N_44950,N_44874);
nand U45034 (N_45034,N_44902,N_44990);
nand U45035 (N_45035,N_44600,N_44737);
and U45036 (N_45036,N_44506,N_44646);
or U45037 (N_45037,N_44863,N_44609);
nor U45038 (N_45038,N_44805,N_44575);
or U45039 (N_45039,N_44637,N_44942);
nand U45040 (N_45040,N_44782,N_44853);
nand U45041 (N_45041,N_44964,N_44572);
nand U45042 (N_45042,N_44514,N_44638);
or U45043 (N_45043,N_44890,N_44961);
nand U45044 (N_45044,N_44962,N_44973);
xnor U45045 (N_45045,N_44815,N_44697);
xor U45046 (N_45046,N_44798,N_44615);
and U45047 (N_45047,N_44801,N_44554);
nor U45048 (N_45048,N_44909,N_44970);
or U45049 (N_45049,N_44541,N_44597);
nand U45050 (N_45050,N_44766,N_44598);
or U45051 (N_45051,N_44894,N_44596);
nor U45052 (N_45052,N_44868,N_44674);
and U45053 (N_45053,N_44946,N_44657);
nand U45054 (N_45054,N_44603,N_44660);
or U45055 (N_45055,N_44937,N_44831);
nand U45056 (N_45056,N_44938,N_44811);
or U45057 (N_45057,N_44834,N_44887);
nand U45058 (N_45058,N_44716,N_44763);
nand U45059 (N_45059,N_44914,N_44983);
xor U45060 (N_45060,N_44727,N_44710);
xor U45061 (N_45061,N_44951,N_44563);
nand U45062 (N_45062,N_44567,N_44877);
nor U45063 (N_45063,N_44531,N_44911);
nor U45064 (N_45064,N_44593,N_44523);
nor U45065 (N_45065,N_44639,N_44886);
xor U45066 (N_45066,N_44994,N_44544);
nor U45067 (N_45067,N_44623,N_44532);
xnor U45068 (N_45068,N_44743,N_44529);
and U45069 (N_45069,N_44840,N_44975);
nor U45070 (N_45070,N_44713,N_44916);
or U45071 (N_45071,N_44957,N_44574);
xor U45072 (N_45072,N_44501,N_44885);
or U45073 (N_45073,N_44562,N_44963);
nor U45074 (N_45074,N_44618,N_44832);
or U45075 (N_45075,N_44816,N_44851);
xor U45076 (N_45076,N_44566,N_44714);
xor U45077 (N_45077,N_44536,N_44992);
and U45078 (N_45078,N_44898,N_44619);
and U45079 (N_45079,N_44881,N_44935);
nand U45080 (N_45080,N_44847,N_44936);
or U45081 (N_45081,N_44601,N_44852);
nand U45082 (N_45082,N_44932,N_44860);
xor U45083 (N_45083,N_44583,N_44800);
or U45084 (N_45084,N_44991,N_44565);
and U45085 (N_45085,N_44949,N_44729);
or U45086 (N_45086,N_44510,N_44725);
nor U45087 (N_45087,N_44841,N_44806);
or U45088 (N_45088,N_44533,N_44582);
nor U45089 (N_45089,N_44742,N_44979);
or U45090 (N_45090,N_44571,N_44895);
xnor U45091 (N_45091,N_44518,N_44828);
or U45092 (N_45092,N_44783,N_44896);
xor U45093 (N_45093,N_44795,N_44717);
or U45094 (N_45094,N_44698,N_44808);
nand U45095 (N_45095,N_44879,N_44839);
and U45096 (N_45096,N_44681,N_44662);
nor U45097 (N_45097,N_44844,N_44519);
and U45098 (N_45098,N_44693,N_44703);
nand U45099 (N_45099,N_44788,N_44836);
nor U45100 (N_45100,N_44837,N_44592);
nor U45101 (N_45101,N_44621,N_44826);
and U45102 (N_45102,N_44680,N_44794);
and U45103 (N_45103,N_44649,N_44611);
nor U45104 (N_45104,N_44897,N_44521);
nand U45105 (N_45105,N_44508,N_44803);
and U45106 (N_45106,N_44629,N_44527);
nor U45107 (N_45107,N_44723,N_44733);
and U45108 (N_45108,N_44689,N_44578);
and U45109 (N_45109,N_44789,N_44920);
nand U45110 (N_45110,N_44982,N_44977);
nand U45111 (N_45111,N_44741,N_44555);
xor U45112 (N_45112,N_44792,N_44870);
xor U45113 (N_45113,N_44864,N_44995);
nand U45114 (N_45114,N_44705,N_44939);
nand U45115 (N_45115,N_44960,N_44653);
nand U45116 (N_45116,N_44882,N_44759);
or U45117 (N_45117,N_44827,N_44819);
xnor U45118 (N_45118,N_44595,N_44685);
and U45119 (N_45119,N_44775,N_44712);
nand U45120 (N_45120,N_44738,N_44802);
xnor U45121 (N_45121,N_44987,N_44652);
xnor U45122 (N_45122,N_44976,N_44612);
or U45123 (N_45123,N_44669,N_44958);
nand U45124 (N_45124,N_44658,N_44665);
xnor U45125 (N_45125,N_44812,N_44684);
and U45126 (N_45126,N_44644,N_44735);
nor U45127 (N_45127,N_44884,N_44966);
nor U45128 (N_45128,N_44721,N_44918);
nor U45129 (N_45129,N_44569,N_44627);
and U45130 (N_45130,N_44659,N_44913);
nor U45131 (N_45131,N_44579,N_44756);
and U45132 (N_45132,N_44668,N_44650);
nand U45133 (N_45133,N_44700,N_44751);
and U45134 (N_45134,N_44767,N_44647);
nand U45135 (N_45135,N_44610,N_44679);
nand U45136 (N_45136,N_44702,N_44807);
or U45137 (N_45137,N_44880,N_44707);
nand U45138 (N_45138,N_44528,N_44944);
nor U45139 (N_45139,N_44943,N_44522);
and U45140 (N_45140,N_44585,N_44999);
or U45141 (N_45141,N_44604,N_44875);
nor U45142 (N_45142,N_44833,N_44607);
nor U45143 (N_45143,N_44545,N_44628);
and U45144 (N_45144,N_44503,N_44769);
nand U45145 (N_45145,N_44633,N_44687);
or U45146 (N_45146,N_44570,N_44930);
or U45147 (N_45147,N_44757,N_44675);
and U45148 (N_45148,N_44590,N_44919);
xnor U45149 (N_45149,N_44825,N_44586);
xnor U45150 (N_45150,N_44764,N_44690);
or U45151 (N_45151,N_44587,N_44754);
and U45152 (N_45152,N_44835,N_44969);
nand U45153 (N_45153,N_44925,N_44591);
nor U45154 (N_45154,N_44576,N_44888);
nor U45155 (N_45155,N_44829,N_44796);
xnor U45156 (N_45156,N_44866,N_44667);
nor U45157 (N_45157,N_44683,N_44632);
nand U45158 (N_45158,N_44988,N_44677);
xor U45159 (N_45159,N_44912,N_44648);
nor U45160 (N_45160,N_44744,N_44762);
nand U45161 (N_45161,N_44580,N_44780);
nand U45162 (N_45162,N_44846,N_44589);
or U45163 (N_45163,N_44641,N_44927);
xor U45164 (N_45164,N_44781,N_44814);
and U45165 (N_45165,N_44599,N_44787);
or U45166 (N_45166,N_44747,N_44552);
nand U45167 (N_45167,N_44843,N_44854);
nand U45168 (N_45168,N_44797,N_44984);
nand U45169 (N_45169,N_44923,N_44905);
or U45170 (N_45170,N_44671,N_44753);
nor U45171 (N_45171,N_44981,N_44940);
or U45172 (N_45172,N_44778,N_44666);
and U45173 (N_45173,N_44974,N_44551);
nor U45174 (N_45174,N_44651,N_44556);
nand U45175 (N_45175,N_44577,N_44965);
and U45176 (N_45176,N_44878,N_44883);
nor U45177 (N_45177,N_44517,N_44770);
xor U45178 (N_45178,N_44719,N_44986);
nor U45179 (N_45179,N_44538,N_44971);
nand U45180 (N_45180,N_44626,N_44540);
nor U45181 (N_45181,N_44749,N_44830);
nand U45182 (N_45182,N_44515,N_44622);
nand U45183 (N_45183,N_44809,N_44959);
and U45184 (N_45184,N_44934,N_44790);
and U45185 (N_45185,N_44941,N_44594);
or U45186 (N_45186,N_44873,N_44670);
xnor U45187 (N_45187,N_44568,N_44581);
nand U45188 (N_45188,N_44904,N_44804);
nand U45189 (N_45189,N_44758,N_44535);
nor U45190 (N_45190,N_44774,N_44630);
xor U45191 (N_45191,N_44711,N_44823);
xor U45192 (N_45192,N_44872,N_44731);
nand U45193 (N_45193,N_44917,N_44726);
and U45194 (N_45194,N_44720,N_44740);
and U45195 (N_45195,N_44634,N_44750);
nand U45196 (N_45196,N_44871,N_44550);
or U45197 (N_45197,N_44526,N_44972);
xnor U45198 (N_45198,N_44656,N_44537);
and U45199 (N_45199,N_44893,N_44838);
nand U45200 (N_45200,N_44985,N_44945);
and U45201 (N_45201,N_44907,N_44892);
xor U45202 (N_45202,N_44561,N_44760);
and U45203 (N_45203,N_44661,N_44899);
xnor U45204 (N_45204,N_44850,N_44948);
or U45205 (N_45205,N_44588,N_44817);
or U45206 (N_45206,N_44616,N_44672);
or U45207 (N_45207,N_44715,N_44709);
xnor U45208 (N_45208,N_44614,N_44865);
or U45209 (N_45209,N_44859,N_44746);
or U45210 (N_45210,N_44855,N_44664);
and U45211 (N_45211,N_44998,N_44509);
or U45212 (N_45212,N_44931,N_44613);
and U45213 (N_45213,N_44728,N_44953);
and U45214 (N_45214,N_44663,N_44821);
nor U45215 (N_45215,N_44845,N_44511);
nand U45216 (N_45216,N_44500,N_44718);
and U45217 (N_45217,N_44900,N_44691);
or U45218 (N_45218,N_44608,N_44520);
xor U45219 (N_45219,N_44559,N_44688);
nand U45220 (N_45220,N_44722,N_44791);
nor U45221 (N_45221,N_44724,N_44889);
and U45222 (N_45222,N_44558,N_44952);
or U45223 (N_45223,N_44507,N_44524);
xnor U45224 (N_45224,N_44771,N_44978);
nand U45225 (N_45225,N_44624,N_44547);
and U45226 (N_45226,N_44734,N_44676);
and U45227 (N_45227,N_44922,N_44695);
or U45228 (N_45228,N_44786,N_44862);
and U45229 (N_45229,N_44708,N_44686);
nor U45230 (N_45230,N_44955,N_44933);
or U45231 (N_45231,N_44620,N_44810);
nor U45232 (N_45232,N_44915,N_44539);
xnor U45233 (N_45233,N_44910,N_44692);
and U45234 (N_45234,N_44785,N_44706);
nor U45235 (N_45235,N_44542,N_44779);
nor U45236 (N_45236,N_44699,N_44867);
nor U45237 (N_45237,N_44546,N_44732);
and U45238 (N_45238,N_44761,N_44773);
xor U45239 (N_45239,N_44784,N_44989);
xnor U45240 (N_45240,N_44776,N_44813);
nand U45241 (N_45241,N_44929,N_44793);
and U45242 (N_45242,N_44772,N_44736);
or U45243 (N_45243,N_44861,N_44967);
xnor U45244 (N_45244,N_44745,N_44765);
nor U45245 (N_45245,N_44643,N_44908);
and U45246 (N_45246,N_44636,N_44739);
or U45247 (N_45247,N_44553,N_44502);
xor U45248 (N_45248,N_44504,N_44768);
or U45249 (N_45249,N_44696,N_44926);
nor U45250 (N_45250,N_44775,N_44722);
nor U45251 (N_45251,N_44921,N_44993);
nor U45252 (N_45252,N_44709,N_44518);
nor U45253 (N_45253,N_44619,N_44994);
or U45254 (N_45254,N_44523,N_44599);
or U45255 (N_45255,N_44807,N_44972);
nand U45256 (N_45256,N_44606,N_44814);
nor U45257 (N_45257,N_44673,N_44573);
or U45258 (N_45258,N_44556,N_44782);
or U45259 (N_45259,N_44930,N_44836);
xor U45260 (N_45260,N_44807,N_44980);
nor U45261 (N_45261,N_44911,N_44830);
xnor U45262 (N_45262,N_44644,N_44993);
nor U45263 (N_45263,N_44787,N_44550);
and U45264 (N_45264,N_44740,N_44629);
xor U45265 (N_45265,N_44983,N_44927);
nor U45266 (N_45266,N_44713,N_44824);
and U45267 (N_45267,N_44924,N_44767);
and U45268 (N_45268,N_44875,N_44745);
xor U45269 (N_45269,N_44915,N_44700);
nor U45270 (N_45270,N_44933,N_44843);
nand U45271 (N_45271,N_44816,N_44735);
or U45272 (N_45272,N_44555,N_44825);
and U45273 (N_45273,N_44829,N_44674);
nand U45274 (N_45274,N_44752,N_44723);
or U45275 (N_45275,N_44817,N_44603);
or U45276 (N_45276,N_44932,N_44779);
and U45277 (N_45277,N_44975,N_44973);
and U45278 (N_45278,N_44915,N_44753);
and U45279 (N_45279,N_44785,N_44904);
or U45280 (N_45280,N_44880,N_44702);
nand U45281 (N_45281,N_44821,N_44519);
or U45282 (N_45282,N_44713,N_44811);
nor U45283 (N_45283,N_44524,N_44570);
xnor U45284 (N_45284,N_44952,N_44814);
or U45285 (N_45285,N_44889,N_44924);
and U45286 (N_45286,N_44869,N_44640);
nand U45287 (N_45287,N_44636,N_44845);
or U45288 (N_45288,N_44714,N_44919);
nor U45289 (N_45289,N_44815,N_44922);
nand U45290 (N_45290,N_44593,N_44783);
xor U45291 (N_45291,N_44522,N_44616);
nand U45292 (N_45292,N_44976,N_44826);
or U45293 (N_45293,N_44586,N_44687);
xor U45294 (N_45294,N_44512,N_44776);
or U45295 (N_45295,N_44774,N_44652);
xnor U45296 (N_45296,N_44971,N_44750);
and U45297 (N_45297,N_44899,N_44826);
nor U45298 (N_45298,N_44940,N_44893);
nand U45299 (N_45299,N_44964,N_44769);
xnor U45300 (N_45300,N_44546,N_44709);
and U45301 (N_45301,N_44748,N_44646);
xor U45302 (N_45302,N_44730,N_44980);
xnor U45303 (N_45303,N_44538,N_44926);
nor U45304 (N_45304,N_44523,N_44689);
or U45305 (N_45305,N_44894,N_44847);
nor U45306 (N_45306,N_44933,N_44891);
nand U45307 (N_45307,N_44948,N_44627);
xor U45308 (N_45308,N_44976,N_44591);
or U45309 (N_45309,N_44657,N_44863);
and U45310 (N_45310,N_44690,N_44657);
or U45311 (N_45311,N_44680,N_44913);
nor U45312 (N_45312,N_44953,N_44564);
or U45313 (N_45313,N_44661,N_44563);
nand U45314 (N_45314,N_44808,N_44695);
or U45315 (N_45315,N_44690,N_44992);
nor U45316 (N_45316,N_44969,N_44905);
and U45317 (N_45317,N_44527,N_44706);
nand U45318 (N_45318,N_44540,N_44817);
nor U45319 (N_45319,N_44533,N_44519);
nand U45320 (N_45320,N_44861,N_44668);
nor U45321 (N_45321,N_44798,N_44595);
or U45322 (N_45322,N_44655,N_44650);
or U45323 (N_45323,N_44859,N_44947);
or U45324 (N_45324,N_44906,N_44880);
and U45325 (N_45325,N_44805,N_44545);
or U45326 (N_45326,N_44922,N_44555);
nor U45327 (N_45327,N_44928,N_44962);
or U45328 (N_45328,N_44980,N_44623);
nor U45329 (N_45329,N_44786,N_44808);
nor U45330 (N_45330,N_44869,N_44828);
nand U45331 (N_45331,N_44913,N_44881);
nor U45332 (N_45332,N_44690,N_44876);
nand U45333 (N_45333,N_44909,N_44605);
and U45334 (N_45334,N_44806,N_44545);
nor U45335 (N_45335,N_44948,N_44557);
nand U45336 (N_45336,N_44576,N_44951);
or U45337 (N_45337,N_44703,N_44821);
or U45338 (N_45338,N_44814,N_44948);
and U45339 (N_45339,N_44586,N_44615);
and U45340 (N_45340,N_44684,N_44769);
or U45341 (N_45341,N_44957,N_44987);
or U45342 (N_45342,N_44813,N_44626);
and U45343 (N_45343,N_44721,N_44905);
xor U45344 (N_45344,N_44937,N_44771);
xor U45345 (N_45345,N_44918,N_44750);
nand U45346 (N_45346,N_44856,N_44564);
nand U45347 (N_45347,N_44745,N_44580);
and U45348 (N_45348,N_44978,N_44511);
xor U45349 (N_45349,N_44960,N_44760);
or U45350 (N_45350,N_44715,N_44621);
nand U45351 (N_45351,N_44784,N_44889);
nand U45352 (N_45352,N_44768,N_44932);
nor U45353 (N_45353,N_44719,N_44912);
xnor U45354 (N_45354,N_44659,N_44800);
or U45355 (N_45355,N_44545,N_44820);
and U45356 (N_45356,N_44518,N_44689);
or U45357 (N_45357,N_44767,N_44838);
xnor U45358 (N_45358,N_44700,N_44758);
and U45359 (N_45359,N_44677,N_44652);
xor U45360 (N_45360,N_44931,N_44732);
xor U45361 (N_45361,N_44970,N_44577);
or U45362 (N_45362,N_44959,N_44545);
nand U45363 (N_45363,N_44932,N_44775);
or U45364 (N_45364,N_44963,N_44535);
and U45365 (N_45365,N_44997,N_44779);
or U45366 (N_45366,N_44972,N_44594);
nor U45367 (N_45367,N_44933,N_44736);
nor U45368 (N_45368,N_44578,N_44594);
or U45369 (N_45369,N_44893,N_44956);
xnor U45370 (N_45370,N_44860,N_44961);
or U45371 (N_45371,N_44806,N_44877);
xor U45372 (N_45372,N_44696,N_44769);
nand U45373 (N_45373,N_44586,N_44568);
xor U45374 (N_45374,N_44987,N_44800);
and U45375 (N_45375,N_44843,N_44985);
and U45376 (N_45376,N_44640,N_44776);
nor U45377 (N_45377,N_44754,N_44712);
nor U45378 (N_45378,N_44689,N_44989);
nand U45379 (N_45379,N_44887,N_44919);
nand U45380 (N_45380,N_44897,N_44816);
and U45381 (N_45381,N_44666,N_44727);
or U45382 (N_45382,N_44744,N_44507);
nor U45383 (N_45383,N_44932,N_44695);
and U45384 (N_45384,N_44545,N_44622);
or U45385 (N_45385,N_44897,N_44741);
nor U45386 (N_45386,N_44634,N_44562);
or U45387 (N_45387,N_44683,N_44752);
xnor U45388 (N_45388,N_44787,N_44794);
and U45389 (N_45389,N_44780,N_44890);
and U45390 (N_45390,N_44919,N_44660);
xnor U45391 (N_45391,N_44549,N_44676);
nand U45392 (N_45392,N_44706,N_44883);
nand U45393 (N_45393,N_44760,N_44579);
or U45394 (N_45394,N_44587,N_44816);
nor U45395 (N_45395,N_44694,N_44600);
nor U45396 (N_45396,N_44707,N_44712);
nand U45397 (N_45397,N_44642,N_44875);
or U45398 (N_45398,N_44998,N_44670);
nor U45399 (N_45399,N_44877,N_44812);
and U45400 (N_45400,N_44700,N_44699);
and U45401 (N_45401,N_44668,N_44597);
nand U45402 (N_45402,N_44900,N_44927);
nand U45403 (N_45403,N_44734,N_44729);
nand U45404 (N_45404,N_44792,N_44963);
nor U45405 (N_45405,N_44960,N_44687);
nor U45406 (N_45406,N_44728,N_44987);
and U45407 (N_45407,N_44503,N_44760);
xor U45408 (N_45408,N_44909,N_44890);
and U45409 (N_45409,N_44699,N_44859);
nand U45410 (N_45410,N_44951,N_44623);
xnor U45411 (N_45411,N_44993,N_44817);
or U45412 (N_45412,N_44880,N_44763);
nor U45413 (N_45413,N_44678,N_44797);
nand U45414 (N_45414,N_44529,N_44772);
or U45415 (N_45415,N_44730,N_44881);
nand U45416 (N_45416,N_44669,N_44813);
nand U45417 (N_45417,N_44695,N_44969);
and U45418 (N_45418,N_44540,N_44811);
xnor U45419 (N_45419,N_44855,N_44563);
xor U45420 (N_45420,N_44630,N_44629);
and U45421 (N_45421,N_44589,N_44958);
nand U45422 (N_45422,N_44725,N_44796);
nor U45423 (N_45423,N_44895,N_44680);
or U45424 (N_45424,N_44924,N_44973);
nor U45425 (N_45425,N_44628,N_44521);
or U45426 (N_45426,N_44530,N_44655);
xor U45427 (N_45427,N_44540,N_44721);
xor U45428 (N_45428,N_44936,N_44920);
xnor U45429 (N_45429,N_44855,N_44711);
nor U45430 (N_45430,N_44589,N_44938);
or U45431 (N_45431,N_44948,N_44637);
and U45432 (N_45432,N_44736,N_44575);
and U45433 (N_45433,N_44759,N_44802);
xor U45434 (N_45434,N_44830,N_44641);
nand U45435 (N_45435,N_44996,N_44903);
xnor U45436 (N_45436,N_44994,N_44694);
or U45437 (N_45437,N_44668,N_44745);
or U45438 (N_45438,N_44659,N_44742);
nor U45439 (N_45439,N_44819,N_44633);
and U45440 (N_45440,N_44740,N_44852);
xor U45441 (N_45441,N_44818,N_44599);
nand U45442 (N_45442,N_44622,N_44522);
xor U45443 (N_45443,N_44824,N_44809);
nand U45444 (N_45444,N_44660,N_44973);
nor U45445 (N_45445,N_44638,N_44531);
nor U45446 (N_45446,N_44589,N_44584);
and U45447 (N_45447,N_44944,N_44536);
or U45448 (N_45448,N_44595,N_44835);
xor U45449 (N_45449,N_44960,N_44574);
or U45450 (N_45450,N_44697,N_44678);
nand U45451 (N_45451,N_44522,N_44705);
nand U45452 (N_45452,N_44705,N_44759);
nand U45453 (N_45453,N_44810,N_44623);
or U45454 (N_45454,N_44974,N_44882);
nor U45455 (N_45455,N_44561,N_44876);
or U45456 (N_45456,N_44993,N_44759);
or U45457 (N_45457,N_44881,N_44598);
xnor U45458 (N_45458,N_44689,N_44532);
and U45459 (N_45459,N_44638,N_44716);
and U45460 (N_45460,N_44713,N_44934);
nand U45461 (N_45461,N_44868,N_44557);
or U45462 (N_45462,N_44752,N_44843);
nor U45463 (N_45463,N_44546,N_44929);
nor U45464 (N_45464,N_44539,N_44508);
nand U45465 (N_45465,N_44920,N_44654);
nor U45466 (N_45466,N_44541,N_44996);
nand U45467 (N_45467,N_44792,N_44629);
nor U45468 (N_45468,N_44706,N_44812);
and U45469 (N_45469,N_44962,N_44858);
and U45470 (N_45470,N_44708,N_44890);
and U45471 (N_45471,N_44958,N_44807);
nand U45472 (N_45472,N_44693,N_44748);
or U45473 (N_45473,N_44960,N_44883);
or U45474 (N_45474,N_44753,N_44909);
and U45475 (N_45475,N_44671,N_44978);
or U45476 (N_45476,N_44663,N_44825);
and U45477 (N_45477,N_44555,N_44816);
nor U45478 (N_45478,N_44520,N_44894);
nor U45479 (N_45479,N_44655,N_44780);
nand U45480 (N_45480,N_44524,N_44919);
nor U45481 (N_45481,N_44500,N_44892);
nand U45482 (N_45482,N_44963,N_44701);
and U45483 (N_45483,N_44655,N_44626);
xor U45484 (N_45484,N_44928,N_44836);
xor U45485 (N_45485,N_44737,N_44824);
or U45486 (N_45486,N_44880,N_44630);
and U45487 (N_45487,N_44670,N_44813);
and U45488 (N_45488,N_44847,N_44601);
nor U45489 (N_45489,N_44815,N_44692);
nor U45490 (N_45490,N_44786,N_44520);
xnor U45491 (N_45491,N_44530,N_44541);
nand U45492 (N_45492,N_44798,N_44980);
and U45493 (N_45493,N_44640,N_44757);
nand U45494 (N_45494,N_44982,N_44955);
or U45495 (N_45495,N_44591,N_44747);
xor U45496 (N_45496,N_44941,N_44980);
nand U45497 (N_45497,N_44680,N_44917);
nand U45498 (N_45498,N_44578,N_44874);
xnor U45499 (N_45499,N_44879,N_44530);
nor U45500 (N_45500,N_45421,N_45397);
nor U45501 (N_45501,N_45072,N_45135);
and U45502 (N_45502,N_45271,N_45231);
nand U45503 (N_45503,N_45483,N_45185);
and U45504 (N_45504,N_45443,N_45149);
nor U45505 (N_45505,N_45468,N_45109);
xnor U45506 (N_45506,N_45199,N_45493);
xnor U45507 (N_45507,N_45080,N_45101);
nor U45508 (N_45508,N_45300,N_45254);
and U45509 (N_45509,N_45447,N_45337);
or U45510 (N_45510,N_45037,N_45496);
and U45511 (N_45511,N_45154,N_45031);
nor U45512 (N_45512,N_45157,N_45373);
or U45513 (N_45513,N_45480,N_45352);
nor U45514 (N_45514,N_45347,N_45115);
nand U45515 (N_45515,N_45329,N_45438);
nor U45516 (N_45516,N_45224,N_45490);
nand U45517 (N_45517,N_45471,N_45140);
nand U45518 (N_45518,N_45497,N_45425);
and U45519 (N_45519,N_45469,N_45048);
nor U45520 (N_45520,N_45086,N_45121);
xor U45521 (N_45521,N_45244,N_45200);
xnor U45522 (N_45522,N_45420,N_45124);
and U45523 (N_45523,N_45044,N_45348);
and U45524 (N_45524,N_45257,N_45171);
nand U45525 (N_45525,N_45407,N_45188);
nor U45526 (N_45526,N_45223,N_45293);
or U45527 (N_45527,N_45378,N_45346);
nor U45528 (N_45528,N_45298,N_45019);
nor U45529 (N_45529,N_45301,N_45082);
and U45530 (N_45530,N_45391,N_45266);
nand U45531 (N_45531,N_45477,N_45056);
nand U45532 (N_45532,N_45076,N_45345);
or U45533 (N_45533,N_45498,N_45302);
or U45534 (N_45534,N_45470,N_45032);
or U45535 (N_45535,N_45398,N_45338);
nand U45536 (N_45536,N_45023,N_45330);
xor U45537 (N_45537,N_45191,N_45047);
and U45538 (N_45538,N_45299,N_45160);
xnor U45539 (N_45539,N_45116,N_45046);
nand U45540 (N_45540,N_45325,N_45487);
and U45541 (N_45541,N_45451,N_45041);
nand U45542 (N_45542,N_45077,N_45022);
nand U45543 (N_45543,N_45435,N_45152);
and U45544 (N_45544,N_45297,N_45351);
and U45545 (N_45545,N_45144,N_45416);
nor U45546 (N_45546,N_45370,N_45312);
xor U45547 (N_45547,N_45102,N_45481);
xor U45548 (N_45548,N_45081,N_45214);
nand U45549 (N_45549,N_45476,N_45075);
or U45550 (N_45550,N_45431,N_45392);
nand U45551 (N_45551,N_45353,N_45227);
xor U45552 (N_45552,N_45426,N_45473);
nand U45553 (N_45553,N_45276,N_45326);
and U45554 (N_45554,N_45052,N_45073);
xor U45555 (N_45555,N_45317,N_45156);
xnor U45556 (N_45556,N_45252,N_45179);
nor U45557 (N_45557,N_45050,N_45058);
nor U45558 (N_45558,N_45369,N_45226);
nor U45559 (N_45559,N_45322,N_45389);
and U45560 (N_45560,N_45485,N_45452);
and U45561 (N_45561,N_45403,N_45111);
and U45562 (N_45562,N_45122,N_45279);
or U45563 (N_45563,N_45357,N_45282);
and U45564 (N_45564,N_45335,N_45371);
xor U45565 (N_45565,N_45410,N_45368);
nand U45566 (N_45566,N_45098,N_45089);
nand U45567 (N_45567,N_45100,N_45422);
nand U45568 (N_45568,N_45383,N_45139);
and U45569 (N_45569,N_45463,N_45002);
nand U45570 (N_45570,N_45461,N_45495);
and U45571 (N_45571,N_45184,N_45007);
xor U45572 (N_45572,N_45429,N_45021);
xnor U45573 (N_45573,N_45108,N_45138);
and U45574 (N_45574,N_45377,N_45310);
nand U45575 (N_45575,N_45482,N_45183);
nor U45576 (N_45576,N_45024,N_45285);
and U45577 (N_45577,N_45456,N_45268);
or U45578 (N_45578,N_45068,N_45159);
nor U45579 (N_45579,N_45078,N_45394);
or U45580 (N_45580,N_45478,N_45251);
nand U45581 (N_45581,N_45163,N_45363);
xor U45582 (N_45582,N_45386,N_45362);
xnor U45583 (N_45583,N_45492,N_45284);
xor U45584 (N_45584,N_45372,N_45264);
nand U45585 (N_45585,N_45079,N_45265);
nor U45586 (N_45586,N_45256,N_45165);
nand U45587 (N_45587,N_45339,N_45120);
nor U45588 (N_45588,N_45281,N_45094);
xnor U45589 (N_45589,N_45164,N_45187);
and U45590 (N_45590,N_45006,N_45117);
nor U45591 (N_45591,N_45240,N_45074);
and U45592 (N_45592,N_45419,N_45113);
or U45593 (N_45593,N_45427,N_45374);
or U45594 (N_45594,N_45355,N_45143);
and U45595 (N_45595,N_45066,N_45150);
nor U45596 (N_45596,N_45375,N_45393);
and U45597 (N_45597,N_45209,N_45202);
xor U45598 (N_45598,N_45241,N_45270);
nor U45599 (N_45599,N_45408,N_45168);
nor U45600 (N_45600,N_45259,N_45195);
nor U45601 (N_45601,N_45376,N_45177);
xnor U45602 (N_45602,N_45499,N_45258);
nor U45603 (N_45603,N_45027,N_45436);
nor U45604 (N_45604,N_45017,N_45417);
nand U45605 (N_45605,N_45087,N_45071);
nor U45606 (N_45606,N_45475,N_45344);
xnor U45607 (N_45607,N_45448,N_45412);
xnor U45608 (N_45608,N_45083,N_45008);
and U45609 (N_45609,N_45396,N_45439);
xnor U45610 (N_45610,N_45380,N_45367);
and U45611 (N_45611,N_45036,N_45466);
nor U45612 (N_45612,N_45142,N_45220);
and U45613 (N_45613,N_45009,N_45198);
or U45614 (N_45614,N_45053,N_45228);
nand U45615 (N_45615,N_45126,N_45203);
nor U45616 (N_45616,N_45166,N_45016);
or U45617 (N_45617,N_45409,N_45018);
nor U45618 (N_45618,N_45273,N_45324);
or U45619 (N_45619,N_45162,N_45382);
nor U45620 (N_45620,N_45424,N_45028);
xnor U45621 (N_45621,N_45449,N_45494);
nand U45622 (N_45622,N_45360,N_45026);
nand U45623 (N_45623,N_45196,N_45306);
nand U45624 (N_45624,N_45103,N_45385);
and U45625 (N_45625,N_45118,N_45434);
nand U45626 (N_45626,N_45043,N_45450);
xnor U45627 (N_45627,N_45379,N_45356);
nor U45628 (N_45628,N_45381,N_45194);
nand U45629 (N_45629,N_45015,N_45432);
nand U45630 (N_45630,N_45457,N_45446);
nand U45631 (N_45631,N_45000,N_45366);
xnor U45632 (N_45632,N_45328,N_45206);
or U45633 (N_45633,N_45182,N_45211);
nand U45634 (N_45634,N_45225,N_45091);
nor U45635 (N_45635,N_45230,N_45153);
nor U45636 (N_45636,N_45255,N_45405);
xor U45637 (N_45637,N_45316,N_45308);
nor U45638 (N_45638,N_45486,N_45280);
nor U45639 (N_45639,N_45313,N_45004);
xor U45640 (N_45640,N_45218,N_45137);
nand U45641 (N_45641,N_45132,N_45404);
xnor U45642 (N_45642,N_45365,N_45229);
nand U45643 (N_45643,N_45128,N_45092);
nand U45644 (N_45644,N_45341,N_45488);
nand U45645 (N_45645,N_45484,N_45390);
nor U45646 (N_45646,N_45400,N_45105);
and U45647 (N_45647,N_45388,N_45275);
xor U45648 (N_45648,N_45242,N_45296);
and U45649 (N_45649,N_45012,N_45070);
and U45650 (N_45650,N_45084,N_45454);
nand U45651 (N_45651,N_45321,N_45458);
nor U45652 (N_45652,N_45235,N_45472);
nand U45653 (N_45653,N_45358,N_45343);
or U45654 (N_45654,N_45222,N_45148);
nor U45655 (N_45655,N_45042,N_45295);
and U45656 (N_45656,N_45013,N_45130);
xor U45657 (N_45657,N_45181,N_45146);
nor U45658 (N_45658,N_45401,N_45030);
xnor U45659 (N_45659,N_45239,N_45430);
nor U45660 (N_45660,N_45119,N_45413);
or U45661 (N_45661,N_45445,N_45005);
nor U45662 (N_45662,N_45110,N_45263);
or U45663 (N_45663,N_45062,N_45327);
xnor U45664 (N_45664,N_45029,N_45033);
xnor U45665 (N_45665,N_45104,N_45063);
and U45666 (N_45666,N_45272,N_45249);
xnor U45667 (N_45667,N_45387,N_45039);
or U45668 (N_45668,N_45315,N_45290);
and U45669 (N_45669,N_45035,N_45145);
nand U45670 (N_45670,N_45361,N_45215);
xnor U45671 (N_45671,N_45011,N_45020);
nand U45672 (N_45672,N_45283,N_45248);
nor U45673 (N_45673,N_45180,N_45292);
xnor U45674 (N_45674,N_45291,N_45232);
nand U45675 (N_45675,N_45213,N_45418);
nor U45676 (N_45676,N_45437,N_45464);
nor U45677 (N_45677,N_45207,N_45189);
xor U45678 (N_45678,N_45192,N_45141);
nor U45679 (N_45679,N_45267,N_45399);
xor U45680 (N_45680,N_45288,N_45455);
xor U45681 (N_45681,N_45186,N_45136);
nand U45682 (N_45682,N_45287,N_45359);
and U45683 (N_45683,N_45204,N_45061);
nand U45684 (N_45684,N_45057,N_45131);
nor U45685 (N_45685,N_45003,N_45489);
xnor U45686 (N_45686,N_45402,N_45201);
nand U45687 (N_45687,N_45253,N_45233);
nand U45688 (N_45688,N_45054,N_45428);
and U45689 (N_45689,N_45250,N_45114);
nor U45690 (N_45690,N_45085,N_45261);
and U45691 (N_45691,N_45107,N_45190);
nand U45692 (N_45692,N_45155,N_45123);
nand U45693 (N_45693,N_45049,N_45243);
xnor U45694 (N_45694,N_45334,N_45193);
and U45695 (N_45695,N_45034,N_45205);
nor U45696 (N_45696,N_45320,N_45051);
nand U45697 (N_45697,N_45208,N_45350);
or U45698 (N_45698,N_45246,N_45309);
and U45699 (N_45699,N_45414,N_45014);
or U45700 (N_45700,N_45055,N_45133);
nor U45701 (N_45701,N_45197,N_45453);
or U45702 (N_45702,N_45462,N_45169);
nand U45703 (N_45703,N_45170,N_45067);
nor U45704 (N_45704,N_45010,N_45305);
nand U45705 (N_45705,N_45289,N_45444);
xor U45706 (N_45706,N_45090,N_45269);
or U45707 (N_45707,N_45134,N_45040);
or U45708 (N_45708,N_45474,N_45423);
and U45709 (N_45709,N_45060,N_45216);
nand U45710 (N_45710,N_45491,N_45460);
nor U45711 (N_45711,N_45093,N_45440);
or U45712 (N_45712,N_45274,N_45172);
nor U45713 (N_45713,N_45099,N_45314);
nor U45714 (N_45714,N_45178,N_45364);
xnor U45715 (N_45715,N_45059,N_45065);
nor U45716 (N_45716,N_45088,N_45459);
or U45717 (N_45717,N_45095,N_45219);
xnor U45718 (N_45718,N_45303,N_45236);
nor U45719 (N_45719,N_45175,N_45384);
or U45720 (N_45720,N_45415,N_45167);
nand U45721 (N_45721,N_45433,N_45176);
xnor U45722 (N_45722,N_45307,N_45221);
nand U45723 (N_45723,N_45465,N_45411);
xor U45724 (N_45724,N_45262,N_45247);
nor U45725 (N_45725,N_45245,N_45151);
xnor U45726 (N_45726,N_45278,N_45318);
nor U45727 (N_45727,N_45294,N_45277);
and U45728 (N_45728,N_45333,N_45332);
xnor U45729 (N_45729,N_45174,N_45331);
xor U45730 (N_45730,N_45304,N_45349);
and U45731 (N_45731,N_45234,N_45045);
and U45732 (N_45732,N_45237,N_45260);
or U45733 (N_45733,N_45336,N_45323);
nor U45734 (N_45734,N_45106,N_45064);
nand U45735 (N_45735,N_45354,N_45479);
nand U45736 (N_45736,N_45173,N_45311);
or U45737 (N_45737,N_45038,N_45319);
or U45738 (N_45738,N_45467,N_45129);
nand U45739 (N_45739,N_45147,N_45395);
and U45740 (N_45740,N_45340,N_45406);
and U45741 (N_45741,N_45158,N_45441);
nor U45742 (N_45742,N_45001,N_45112);
or U45743 (N_45743,N_45286,N_45442);
or U45744 (N_45744,N_45069,N_45096);
nand U45745 (N_45745,N_45125,N_45217);
and U45746 (N_45746,N_45161,N_45127);
nor U45747 (N_45747,N_45238,N_45025);
nand U45748 (N_45748,N_45097,N_45342);
nand U45749 (N_45749,N_45210,N_45212);
xnor U45750 (N_45750,N_45374,N_45005);
nor U45751 (N_45751,N_45345,N_45304);
xnor U45752 (N_45752,N_45044,N_45459);
and U45753 (N_45753,N_45250,N_45085);
nor U45754 (N_45754,N_45369,N_45160);
xor U45755 (N_45755,N_45149,N_45018);
and U45756 (N_45756,N_45292,N_45147);
xor U45757 (N_45757,N_45451,N_45279);
xnor U45758 (N_45758,N_45156,N_45423);
nand U45759 (N_45759,N_45192,N_45044);
xor U45760 (N_45760,N_45255,N_45187);
nand U45761 (N_45761,N_45351,N_45087);
nor U45762 (N_45762,N_45159,N_45000);
nor U45763 (N_45763,N_45285,N_45052);
xnor U45764 (N_45764,N_45244,N_45331);
xor U45765 (N_45765,N_45377,N_45010);
or U45766 (N_45766,N_45260,N_45261);
or U45767 (N_45767,N_45311,N_45367);
nor U45768 (N_45768,N_45026,N_45186);
or U45769 (N_45769,N_45020,N_45102);
xnor U45770 (N_45770,N_45029,N_45376);
xnor U45771 (N_45771,N_45335,N_45026);
or U45772 (N_45772,N_45364,N_45043);
and U45773 (N_45773,N_45048,N_45407);
xnor U45774 (N_45774,N_45107,N_45049);
nand U45775 (N_45775,N_45198,N_45206);
and U45776 (N_45776,N_45142,N_45499);
nand U45777 (N_45777,N_45151,N_45250);
nor U45778 (N_45778,N_45069,N_45359);
or U45779 (N_45779,N_45355,N_45120);
or U45780 (N_45780,N_45230,N_45312);
or U45781 (N_45781,N_45244,N_45196);
nand U45782 (N_45782,N_45261,N_45464);
xnor U45783 (N_45783,N_45079,N_45117);
or U45784 (N_45784,N_45161,N_45404);
nor U45785 (N_45785,N_45011,N_45059);
and U45786 (N_45786,N_45450,N_45065);
nor U45787 (N_45787,N_45254,N_45087);
nand U45788 (N_45788,N_45364,N_45072);
and U45789 (N_45789,N_45419,N_45269);
xor U45790 (N_45790,N_45339,N_45337);
xnor U45791 (N_45791,N_45088,N_45023);
or U45792 (N_45792,N_45496,N_45043);
or U45793 (N_45793,N_45009,N_45450);
and U45794 (N_45794,N_45120,N_45337);
and U45795 (N_45795,N_45053,N_45381);
xnor U45796 (N_45796,N_45017,N_45428);
and U45797 (N_45797,N_45223,N_45372);
and U45798 (N_45798,N_45095,N_45358);
and U45799 (N_45799,N_45201,N_45188);
xnor U45800 (N_45800,N_45196,N_45157);
nor U45801 (N_45801,N_45472,N_45486);
or U45802 (N_45802,N_45438,N_45082);
or U45803 (N_45803,N_45140,N_45134);
and U45804 (N_45804,N_45025,N_45368);
xnor U45805 (N_45805,N_45397,N_45476);
or U45806 (N_45806,N_45197,N_45155);
nor U45807 (N_45807,N_45084,N_45221);
xnor U45808 (N_45808,N_45140,N_45076);
nor U45809 (N_45809,N_45010,N_45007);
and U45810 (N_45810,N_45490,N_45265);
and U45811 (N_45811,N_45392,N_45169);
nor U45812 (N_45812,N_45207,N_45440);
xor U45813 (N_45813,N_45341,N_45300);
xor U45814 (N_45814,N_45454,N_45133);
or U45815 (N_45815,N_45117,N_45331);
nand U45816 (N_45816,N_45274,N_45385);
or U45817 (N_45817,N_45043,N_45122);
or U45818 (N_45818,N_45085,N_45455);
and U45819 (N_45819,N_45381,N_45356);
nand U45820 (N_45820,N_45108,N_45225);
nor U45821 (N_45821,N_45117,N_45296);
nor U45822 (N_45822,N_45333,N_45321);
and U45823 (N_45823,N_45321,N_45236);
nor U45824 (N_45824,N_45261,N_45416);
or U45825 (N_45825,N_45142,N_45355);
nor U45826 (N_45826,N_45356,N_45158);
and U45827 (N_45827,N_45016,N_45376);
nand U45828 (N_45828,N_45199,N_45293);
xor U45829 (N_45829,N_45313,N_45471);
nor U45830 (N_45830,N_45036,N_45239);
xnor U45831 (N_45831,N_45308,N_45441);
and U45832 (N_45832,N_45432,N_45227);
and U45833 (N_45833,N_45476,N_45230);
xor U45834 (N_45834,N_45303,N_45078);
or U45835 (N_45835,N_45454,N_45370);
and U45836 (N_45836,N_45005,N_45107);
nand U45837 (N_45837,N_45091,N_45430);
xnor U45838 (N_45838,N_45057,N_45053);
or U45839 (N_45839,N_45472,N_45011);
xnor U45840 (N_45840,N_45208,N_45412);
nand U45841 (N_45841,N_45051,N_45283);
nor U45842 (N_45842,N_45107,N_45240);
and U45843 (N_45843,N_45299,N_45296);
xnor U45844 (N_45844,N_45367,N_45420);
and U45845 (N_45845,N_45275,N_45424);
xnor U45846 (N_45846,N_45406,N_45303);
nor U45847 (N_45847,N_45408,N_45308);
nor U45848 (N_45848,N_45379,N_45313);
nor U45849 (N_45849,N_45412,N_45206);
or U45850 (N_45850,N_45130,N_45451);
nand U45851 (N_45851,N_45357,N_45198);
xor U45852 (N_45852,N_45440,N_45417);
xnor U45853 (N_45853,N_45122,N_45169);
or U45854 (N_45854,N_45486,N_45451);
and U45855 (N_45855,N_45447,N_45174);
and U45856 (N_45856,N_45213,N_45307);
nand U45857 (N_45857,N_45066,N_45095);
xnor U45858 (N_45858,N_45290,N_45185);
xor U45859 (N_45859,N_45267,N_45348);
xnor U45860 (N_45860,N_45496,N_45082);
or U45861 (N_45861,N_45201,N_45023);
or U45862 (N_45862,N_45429,N_45197);
and U45863 (N_45863,N_45361,N_45000);
xor U45864 (N_45864,N_45278,N_45454);
and U45865 (N_45865,N_45295,N_45202);
or U45866 (N_45866,N_45261,N_45246);
nand U45867 (N_45867,N_45062,N_45036);
or U45868 (N_45868,N_45393,N_45124);
nand U45869 (N_45869,N_45172,N_45055);
nor U45870 (N_45870,N_45325,N_45089);
xor U45871 (N_45871,N_45419,N_45362);
nor U45872 (N_45872,N_45386,N_45405);
xor U45873 (N_45873,N_45453,N_45336);
and U45874 (N_45874,N_45127,N_45149);
or U45875 (N_45875,N_45460,N_45429);
and U45876 (N_45876,N_45393,N_45100);
nand U45877 (N_45877,N_45083,N_45180);
nand U45878 (N_45878,N_45367,N_45373);
or U45879 (N_45879,N_45093,N_45017);
and U45880 (N_45880,N_45468,N_45149);
xor U45881 (N_45881,N_45039,N_45436);
or U45882 (N_45882,N_45268,N_45476);
nor U45883 (N_45883,N_45230,N_45076);
nor U45884 (N_45884,N_45148,N_45391);
or U45885 (N_45885,N_45025,N_45465);
and U45886 (N_45886,N_45398,N_45418);
nand U45887 (N_45887,N_45229,N_45302);
nand U45888 (N_45888,N_45037,N_45205);
xnor U45889 (N_45889,N_45098,N_45483);
xnor U45890 (N_45890,N_45210,N_45235);
nand U45891 (N_45891,N_45084,N_45169);
and U45892 (N_45892,N_45273,N_45306);
nor U45893 (N_45893,N_45139,N_45394);
xnor U45894 (N_45894,N_45233,N_45227);
nor U45895 (N_45895,N_45185,N_45025);
xor U45896 (N_45896,N_45497,N_45050);
xnor U45897 (N_45897,N_45188,N_45119);
or U45898 (N_45898,N_45481,N_45028);
nand U45899 (N_45899,N_45417,N_45346);
nand U45900 (N_45900,N_45279,N_45278);
and U45901 (N_45901,N_45363,N_45048);
or U45902 (N_45902,N_45178,N_45437);
nor U45903 (N_45903,N_45497,N_45074);
nand U45904 (N_45904,N_45472,N_45189);
nand U45905 (N_45905,N_45236,N_45378);
or U45906 (N_45906,N_45302,N_45269);
and U45907 (N_45907,N_45373,N_45224);
xnor U45908 (N_45908,N_45177,N_45430);
or U45909 (N_45909,N_45368,N_45473);
nand U45910 (N_45910,N_45049,N_45420);
nand U45911 (N_45911,N_45426,N_45219);
and U45912 (N_45912,N_45012,N_45347);
or U45913 (N_45913,N_45492,N_45206);
or U45914 (N_45914,N_45319,N_45238);
nor U45915 (N_45915,N_45399,N_45170);
xnor U45916 (N_45916,N_45455,N_45320);
and U45917 (N_45917,N_45458,N_45388);
nand U45918 (N_45918,N_45121,N_45124);
nand U45919 (N_45919,N_45497,N_45062);
and U45920 (N_45920,N_45120,N_45036);
or U45921 (N_45921,N_45233,N_45400);
xor U45922 (N_45922,N_45386,N_45160);
xor U45923 (N_45923,N_45192,N_45109);
nor U45924 (N_45924,N_45161,N_45423);
nor U45925 (N_45925,N_45231,N_45066);
nand U45926 (N_45926,N_45362,N_45135);
xor U45927 (N_45927,N_45025,N_45278);
xor U45928 (N_45928,N_45288,N_45238);
xnor U45929 (N_45929,N_45051,N_45334);
and U45930 (N_45930,N_45295,N_45257);
nand U45931 (N_45931,N_45374,N_45112);
or U45932 (N_45932,N_45382,N_45173);
nand U45933 (N_45933,N_45102,N_45030);
xnor U45934 (N_45934,N_45302,N_45340);
xor U45935 (N_45935,N_45497,N_45449);
nand U45936 (N_45936,N_45421,N_45280);
nand U45937 (N_45937,N_45253,N_45065);
and U45938 (N_45938,N_45284,N_45440);
nand U45939 (N_45939,N_45079,N_45377);
nor U45940 (N_45940,N_45381,N_45173);
or U45941 (N_45941,N_45415,N_45142);
nor U45942 (N_45942,N_45027,N_45427);
nand U45943 (N_45943,N_45204,N_45443);
nor U45944 (N_45944,N_45331,N_45057);
nand U45945 (N_45945,N_45098,N_45270);
nor U45946 (N_45946,N_45394,N_45025);
xnor U45947 (N_45947,N_45375,N_45363);
xor U45948 (N_45948,N_45338,N_45368);
or U45949 (N_45949,N_45243,N_45468);
and U45950 (N_45950,N_45302,N_45495);
nor U45951 (N_45951,N_45269,N_45190);
or U45952 (N_45952,N_45432,N_45061);
nand U45953 (N_45953,N_45340,N_45323);
and U45954 (N_45954,N_45486,N_45052);
or U45955 (N_45955,N_45100,N_45089);
or U45956 (N_45956,N_45146,N_45114);
or U45957 (N_45957,N_45391,N_45462);
nand U45958 (N_45958,N_45240,N_45191);
or U45959 (N_45959,N_45030,N_45017);
xnor U45960 (N_45960,N_45293,N_45264);
nor U45961 (N_45961,N_45039,N_45393);
or U45962 (N_45962,N_45244,N_45266);
and U45963 (N_45963,N_45467,N_45100);
nor U45964 (N_45964,N_45228,N_45149);
nor U45965 (N_45965,N_45103,N_45280);
nor U45966 (N_45966,N_45350,N_45026);
nor U45967 (N_45967,N_45045,N_45328);
nor U45968 (N_45968,N_45282,N_45064);
nor U45969 (N_45969,N_45158,N_45457);
xnor U45970 (N_45970,N_45090,N_45485);
xor U45971 (N_45971,N_45049,N_45444);
nor U45972 (N_45972,N_45352,N_45455);
or U45973 (N_45973,N_45067,N_45137);
nand U45974 (N_45974,N_45183,N_45043);
and U45975 (N_45975,N_45412,N_45327);
xor U45976 (N_45976,N_45147,N_45210);
xnor U45977 (N_45977,N_45494,N_45031);
nor U45978 (N_45978,N_45172,N_45025);
nand U45979 (N_45979,N_45203,N_45072);
nor U45980 (N_45980,N_45280,N_45390);
or U45981 (N_45981,N_45017,N_45242);
nor U45982 (N_45982,N_45129,N_45154);
nor U45983 (N_45983,N_45483,N_45065);
and U45984 (N_45984,N_45022,N_45383);
or U45985 (N_45985,N_45432,N_45349);
or U45986 (N_45986,N_45300,N_45090);
or U45987 (N_45987,N_45063,N_45424);
nor U45988 (N_45988,N_45073,N_45264);
xor U45989 (N_45989,N_45183,N_45327);
or U45990 (N_45990,N_45160,N_45218);
xnor U45991 (N_45991,N_45164,N_45170);
xor U45992 (N_45992,N_45432,N_45261);
or U45993 (N_45993,N_45140,N_45235);
or U45994 (N_45994,N_45481,N_45420);
xnor U45995 (N_45995,N_45408,N_45145);
nand U45996 (N_45996,N_45159,N_45281);
nand U45997 (N_45997,N_45368,N_45322);
xor U45998 (N_45998,N_45314,N_45386);
or U45999 (N_45999,N_45085,N_45012);
and U46000 (N_46000,N_45840,N_45568);
nor U46001 (N_46001,N_45848,N_45996);
xor U46002 (N_46002,N_45917,N_45944);
xor U46003 (N_46003,N_45652,N_45882);
or U46004 (N_46004,N_45660,N_45961);
xnor U46005 (N_46005,N_45936,N_45622);
nand U46006 (N_46006,N_45763,N_45619);
nor U46007 (N_46007,N_45635,N_45862);
nand U46008 (N_46008,N_45927,N_45623);
nand U46009 (N_46009,N_45574,N_45722);
xnor U46010 (N_46010,N_45863,N_45953);
and U46011 (N_46011,N_45657,N_45867);
and U46012 (N_46012,N_45877,N_45891);
nor U46013 (N_46013,N_45771,N_45933);
xor U46014 (N_46014,N_45922,N_45779);
xor U46015 (N_46015,N_45699,N_45500);
nor U46016 (N_46016,N_45975,N_45904);
xor U46017 (N_46017,N_45666,N_45564);
nand U46018 (N_46018,N_45931,N_45675);
xor U46019 (N_46019,N_45876,N_45719);
nand U46020 (N_46020,N_45560,N_45994);
nand U46021 (N_46021,N_45770,N_45600);
nand U46022 (N_46022,N_45939,N_45769);
xor U46023 (N_46023,N_45506,N_45659);
or U46024 (N_46024,N_45811,N_45875);
and U46025 (N_46025,N_45597,N_45563);
or U46026 (N_46026,N_45911,N_45624);
or U46027 (N_46027,N_45617,N_45578);
and U46028 (N_46028,N_45818,N_45942);
and U46029 (N_46029,N_45856,N_45864);
or U46030 (N_46030,N_45838,N_45705);
nor U46031 (N_46031,N_45787,N_45716);
and U46032 (N_46032,N_45883,N_45805);
and U46033 (N_46033,N_45878,N_45592);
xnor U46034 (N_46034,N_45605,N_45515);
and U46035 (N_46035,N_45648,N_45702);
nor U46036 (N_46036,N_45866,N_45509);
and U46037 (N_46037,N_45566,N_45603);
nor U46038 (N_46038,N_45925,N_45930);
and U46039 (N_46039,N_45545,N_45638);
nand U46040 (N_46040,N_45688,N_45611);
nor U46041 (N_46041,N_45929,N_45681);
nor U46042 (N_46042,N_45541,N_45814);
or U46043 (N_46043,N_45559,N_45663);
nand U46044 (N_46044,N_45923,N_45531);
or U46045 (N_46045,N_45978,N_45621);
and U46046 (N_46046,N_45781,N_45881);
or U46047 (N_46047,N_45569,N_45973);
nand U46048 (N_46048,N_45830,N_45565);
nand U46049 (N_46049,N_45872,N_45668);
and U46050 (N_46050,N_45752,N_45865);
xnor U46051 (N_46051,N_45587,N_45747);
or U46052 (N_46052,N_45520,N_45829);
xor U46053 (N_46053,N_45971,N_45723);
or U46054 (N_46054,N_45616,N_45932);
nand U46055 (N_46055,N_45637,N_45803);
or U46056 (N_46056,N_45573,N_45631);
or U46057 (N_46057,N_45977,N_45860);
nand U46058 (N_46058,N_45711,N_45701);
nor U46059 (N_46059,N_45740,N_45645);
or U46060 (N_46060,N_45679,N_45644);
or U46061 (N_46061,N_45812,N_45780);
xor U46062 (N_46062,N_45585,N_45596);
nand U46063 (N_46063,N_45748,N_45642);
nand U46064 (N_46064,N_45999,N_45976);
and U46065 (N_46065,N_45717,N_45630);
and U46066 (N_46066,N_45698,N_45757);
nor U46067 (N_46067,N_45762,N_45899);
and U46068 (N_46068,N_45547,N_45572);
and U46069 (N_46069,N_45987,N_45553);
xor U46070 (N_46070,N_45767,N_45733);
xor U46071 (N_46071,N_45590,N_45834);
nand U46072 (N_46072,N_45732,N_45676);
xnor U46073 (N_46073,N_45807,N_45993);
nand U46074 (N_46074,N_45998,N_45907);
nor U46075 (N_46075,N_45850,N_45873);
nor U46076 (N_46076,N_45720,N_45709);
and U46077 (N_46077,N_45522,N_45724);
xnor U46078 (N_46078,N_45695,N_45844);
and U46079 (N_46079,N_45949,N_45894);
or U46080 (N_46080,N_45809,N_45859);
nand U46081 (N_46081,N_45888,N_45794);
and U46082 (N_46082,N_45798,N_45683);
xnor U46083 (N_46083,N_45626,N_45627);
and U46084 (N_46084,N_45591,N_45914);
and U46085 (N_46085,N_45649,N_45599);
xnor U46086 (N_46086,N_45754,N_45831);
or U46087 (N_46087,N_45921,N_45575);
and U46088 (N_46088,N_45552,N_45697);
and U46089 (N_46089,N_45963,N_45915);
nor U46090 (N_46090,N_45633,N_45725);
xnor U46091 (N_46091,N_45737,N_45868);
xnor U46092 (N_46092,N_45989,N_45950);
nand U46093 (N_46093,N_45982,N_45728);
nand U46094 (N_46094,N_45775,N_45514);
nand U46095 (N_46095,N_45718,N_45744);
nand U46096 (N_46096,N_45710,N_45551);
and U46097 (N_46097,N_45784,N_45589);
nor U46098 (N_46098,N_45960,N_45510);
or U46099 (N_46099,N_45730,N_45696);
nor U46100 (N_46100,N_45893,N_45693);
xor U46101 (N_46101,N_45952,N_45905);
xnor U46102 (N_46102,N_45542,N_45580);
or U46103 (N_46103,N_45833,N_45595);
and U46104 (N_46104,N_45526,N_45854);
nand U46105 (N_46105,N_45912,N_45614);
xor U46106 (N_46106,N_45707,N_45988);
nand U46107 (N_46107,N_45804,N_45937);
and U46108 (N_46108,N_45581,N_45938);
nand U46109 (N_46109,N_45613,N_45503);
xnor U46110 (N_46110,N_45793,N_45792);
and U46111 (N_46111,N_45691,N_45620);
nor U46112 (N_46112,N_45782,N_45742);
nor U46113 (N_46113,N_45890,N_45667);
or U46114 (N_46114,N_45651,N_45816);
xor U46115 (N_46115,N_45577,N_45874);
or U46116 (N_46116,N_45983,N_45523);
or U46117 (N_46117,N_45682,N_45602);
xor U46118 (N_46118,N_45857,N_45991);
or U46119 (N_46119,N_45897,N_45773);
and U46120 (N_46120,N_45704,N_45632);
nor U46121 (N_46121,N_45579,N_45845);
nand U46122 (N_46122,N_45802,N_45940);
nand U46123 (N_46123,N_45884,N_45653);
nor U46124 (N_46124,N_45511,N_45928);
and U46125 (N_46125,N_45768,N_45760);
nor U46126 (N_46126,N_45822,N_45909);
nand U46127 (N_46127,N_45540,N_45544);
xnor U46128 (N_46128,N_45934,N_45570);
nand U46129 (N_46129,N_45727,N_45828);
or U46130 (N_46130,N_45968,N_45647);
nor U46131 (N_46131,N_45751,N_45690);
nand U46132 (N_46132,N_45734,N_45530);
xor U46133 (N_46133,N_45554,N_45539);
xor U46134 (N_46134,N_45820,N_45819);
xor U46135 (N_46135,N_45549,N_45518);
or U46136 (N_46136,N_45943,N_45853);
and U46137 (N_46137,N_45964,N_45636);
nor U46138 (N_46138,N_45671,N_45835);
or U46139 (N_46139,N_45924,N_45919);
or U46140 (N_46140,N_45852,N_45941);
xor U46141 (N_46141,N_45686,N_45985);
nor U46142 (N_46142,N_45981,N_45684);
nand U46143 (N_46143,N_45995,N_45571);
xnor U46144 (N_46144,N_45516,N_45721);
nand U46145 (N_46145,N_45766,N_45714);
nor U46146 (N_46146,N_45920,N_45739);
xor U46147 (N_46147,N_45821,N_45758);
nand U46148 (N_46148,N_45959,N_45594);
xor U46149 (N_46149,N_45685,N_45629);
or U46150 (N_46150,N_45525,N_45846);
nand U46151 (N_46151,N_45521,N_45532);
nand U46152 (N_46152,N_45741,N_45665);
nand U46153 (N_46153,N_45843,N_45608);
and U46154 (N_46154,N_45745,N_45900);
nand U46155 (N_46155,N_45958,N_45926);
nor U46156 (N_46156,N_45810,N_45842);
or U46157 (N_46157,N_45783,N_45947);
or U46158 (N_46158,N_45885,N_45869);
nor U46159 (N_46159,N_45823,N_45593);
xnor U46160 (N_46160,N_45556,N_45898);
nor U46161 (N_46161,N_45646,N_45508);
and U46162 (N_46162,N_45528,N_45501);
nand U46163 (N_46163,N_45655,N_45913);
xnor U46164 (N_46164,N_45851,N_45796);
xnor U46165 (N_46165,N_45765,N_45533);
xnor U46166 (N_46166,N_45562,N_45678);
or U46167 (N_46167,N_45607,N_45618);
nor U46168 (N_46168,N_45598,N_45965);
xor U46169 (N_46169,N_45650,N_45969);
nor U46170 (N_46170,N_45935,N_45673);
or U46171 (N_46171,N_45896,N_45610);
and U46172 (N_46172,N_45849,N_45847);
or U46173 (N_46173,N_45759,N_45735);
nand U46174 (N_46174,N_45546,N_45827);
nor U46175 (N_46175,N_45879,N_45664);
or U46176 (N_46176,N_45871,N_45756);
or U46177 (N_46177,N_45543,N_45639);
and U46178 (N_46178,N_45708,N_45641);
nand U46179 (N_46179,N_45558,N_45918);
xnor U46180 (N_46180,N_45654,N_45555);
and U46181 (N_46181,N_45791,N_45826);
xnor U46182 (N_46182,N_45670,N_45990);
and U46183 (N_46183,N_45801,N_45946);
nand U46184 (N_46184,N_45538,N_45855);
or U46185 (N_46185,N_45790,N_45750);
nor U46186 (N_46186,N_45910,N_45903);
nand U46187 (N_46187,N_45536,N_45908);
nor U46188 (N_46188,N_45870,N_45601);
and U46189 (N_46189,N_45813,N_45800);
or U46190 (N_46190,N_45797,N_45980);
and U46191 (N_46191,N_45700,N_45956);
and U46192 (N_46192,N_45746,N_45583);
nand U46193 (N_46193,N_45916,N_45502);
nand U46194 (N_46194,N_45694,N_45861);
nand U46195 (N_46195,N_45548,N_45755);
xor U46196 (N_46196,N_45513,N_45764);
or U46197 (N_46197,N_45535,N_45713);
nand U46198 (N_46198,N_45832,N_45776);
nand U46199 (N_46199,N_45886,N_45505);
and U46200 (N_46200,N_45839,N_45966);
xnor U46201 (N_46201,N_45954,N_45517);
xnor U46202 (N_46202,N_45729,N_45625);
nor U46203 (N_46203,N_45692,N_45825);
xor U46204 (N_46204,N_45789,N_45997);
nor U46205 (N_46205,N_45527,N_45836);
or U46206 (N_46206,N_45586,N_45672);
xnor U46207 (N_46207,N_45712,N_45588);
or U46208 (N_46208,N_45512,N_45955);
and U46209 (N_46209,N_45507,N_45680);
nand U46210 (N_46210,N_45529,N_45786);
nand U46211 (N_46211,N_45967,N_45689);
and U46212 (N_46212,N_45669,N_45887);
nand U46213 (N_46213,N_45808,N_45609);
nor U46214 (N_46214,N_45677,N_45992);
xor U46215 (N_46215,N_45726,N_45656);
nand U46216 (N_46216,N_45892,N_45687);
or U46217 (N_46217,N_45615,N_45703);
or U46218 (N_46218,N_45534,N_45902);
xor U46219 (N_46219,N_45761,N_45799);
xnor U46220 (N_46220,N_45785,N_45612);
nand U46221 (N_46221,N_45824,N_45674);
nand U46222 (N_46222,N_45837,N_45906);
nor U46223 (N_46223,N_45582,N_45640);
nand U46224 (N_46224,N_45561,N_45795);
nor U46225 (N_46225,N_45736,N_45972);
nand U46226 (N_46226,N_45979,N_45817);
or U46227 (N_46227,N_45643,N_45524);
xnor U46228 (N_46228,N_45880,N_45895);
nand U46229 (N_46229,N_45628,N_45778);
nor U46230 (N_46230,N_45550,N_45962);
nor U46231 (N_46231,N_45858,N_45634);
and U46232 (N_46232,N_45715,N_45731);
nor U46233 (N_46233,N_45567,N_45604);
and U46234 (N_46234,N_45537,N_45504);
and U46235 (N_46235,N_45519,N_45901);
or U46236 (N_46236,N_45584,N_45970);
and U46237 (N_46237,N_45806,N_45986);
xor U46238 (N_46238,N_45841,N_45576);
and U46239 (N_46239,N_45706,N_45974);
nor U46240 (N_46240,N_45777,N_45945);
nand U46241 (N_46241,N_45889,N_45772);
or U46242 (N_46242,N_45606,N_45984);
or U46243 (N_46243,N_45774,N_45753);
nand U46244 (N_46244,N_45662,N_45948);
and U46245 (N_46245,N_45957,N_45951);
nor U46246 (N_46246,N_45743,N_45788);
or U46247 (N_46247,N_45658,N_45749);
or U46248 (N_46248,N_45815,N_45738);
nand U46249 (N_46249,N_45661,N_45557);
xor U46250 (N_46250,N_45578,N_45557);
nand U46251 (N_46251,N_45644,N_45512);
and U46252 (N_46252,N_45935,N_45956);
xor U46253 (N_46253,N_45707,N_45749);
or U46254 (N_46254,N_45705,N_45505);
nand U46255 (N_46255,N_45612,N_45691);
or U46256 (N_46256,N_45965,N_45843);
and U46257 (N_46257,N_45695,N_45874);
nand U46258 (N_46258,N_45990,N_45969);
or U46259 (N_46259,N_45999,N_45962);
or U46260 (N_46260,N_45628,N_45723);
and U46261 (N_46261,N_45743,N_45796);
xor U46262 (N_46262,N_45877,N_45651);
nor U46263 (N_46263,N_45751,N_45925);
and U46264 (N_46264,N_45897,N_45807);
nand U46265 (N_46265,N_45917,N_45793);
or U46266 (N_46266,N_45636,N_45915);
xnor U46267 (N_46267,N_45931,N_45796);
xnor U46268 (N_46268,N_45779,N_45928);
nand U46269 (N_46269,N_45629,N_45605);
nor U46270 (N_46270,N_45617,N_45830);
xor U46271 (N_46271,N_45868,N_45931);
nor U46272 (N_46272,N_45636,N_45583);
and U46273 (N_46273,N_45800,N_45627);
nand U46274 (N_46274,N_45807,N_45809);
and U46275 (N_46275,N_45526,N_45961);
or U46276 (N_46276,N_45862,N_45905);
nor U46277 (N_46277,N_45750,N_45883);
or U46278 (N_46278,N_45793,N_45895);
nor U46279 (N_46279,N_45679,N_45945);
and U46280 (N_46280,N_45907,N_45934);
xor U46281 (N_46281,N_45972,N_45825);
xnor U46282 (N_46282,N_45802,N_45842);
nand U46283 (N_46283,N_45769,N_45531);
nand U46284 (N_46284,N_45954,N_45869);
nor U46285 (N_46285,N_45953,N_45576);
xor U46286 (N_46286,N_45624,N_45670);
nor U46287 (N_46287,N_45990,N_45755);
and U46288 (N_46288,N_45508,N_45687);
nand U46289 (N_46289,N_45915,N_45938);
or U46290 (N_46290,N_45854,N_45744);
or U46291 (N_46291,N_45937,N_45805);
nor U46292 (N_46292,N_45815,N_45797);
nor U46293 (N_46293,N_45958,N_45835);
nand U46294 (N_46294,N_45878,N_45695);
nor U46295 (N_46295,N_45545,N_45608);
nor U46296 (N_46296,N_45671,N_45668);
and U46297 (N_46297,N_45571,N_45945);
nor U46298 (N_46298,N_45738,N_45729);
xnor U46299 (N_46299,N_45941,N_45743);
xnor U46300 (N_46300,N_45957,N_45789);
xnor U46301 (N_46301,N_45926,N_45749);
or U46302 (N_46302,N_45587,N_45721);
xnor U46303 (N_46303,N_45617,N_45955);
nor U46304 (N_46304,N_45551,N_45650);
nand U46305 (N_46305,N_45547,N_45665);
or U46306 (N_46306,N_45780,N_45986);
or U46307 (N_46307,N_45758,N_45730);
or U46308 (N_46308,N_45795,N_45860);
and U46309 (N_46309,N_45630,N_45632);
and U46310 (N_46310,N_45970,N_45817);
or U46311 (N_46311,N_45867,N_45605);
xnor U46312 (N_46312,N_45749,N_45938);
nor U46313 (N_46313,N_45933,N_45942);
xor U46314 (N_46314,N_45835,N_45629);
xnor U46315 (N_46315,N_45603,N_45598);
nand U46316 (N_46316,N_45775,N_45948);
nand U46317 (N_46317,N_45832,N_45990);
nor U46318 (N_46318,N_45814,N_45628);
nor U46319 (N_46319,N_45711,N_45821);
or U46320 (N_46320,N_45668,N_45587);
and U46321 (N_46321,N_45639,N_45765);
or U46322 (N_46322,N_45522,N_45533);
nand U46323 (N_46323,N_45813,N_45505);
xnor U46324 (N_46324,N_45556,N_45786);
and U46325 (N_46325,N_45758,N_45872);
xor U46326 (N_46326,N_45985,N_45525);
xnor U46327 (N_46327,N_45898,N_45530);
nand U46328 (N_46328,N_45840,N_45791);
xnor U46329 (N_46329,N_45758,N_45628);
xnor U46330 (N_46330,N_45646,N_45582);
xnor U46331 (N_46331,N_45509,N_45850);
xnor U46332 (N_46332,N_45657,N_45856);
or U46333 (N_46333,N_45825,N_45841);
and U46334 (N_46334,N_45620,N_45762);
xnor U46335 (N_46335,N_45810,N_45840);
nand U46336 (N_46336,N_45780,N_45880);
nand U46337 (N_46337,N_45600,N_45868);
and U46338 (N_46338,N_45868,N_45581);
nand U46339 (N_46339,N_45568,N_45703);
or U46340 (N_46340,N_45886,N_45791);
or U46341 (N_46341,N_45616,N_45570);
or U46342 (N_46342,N_45532,N_45851);
or U46343 (N_46343,N_45773,N_45541);
xor U46344 (N_46344,N_45803,N_45751);
xor U46345 (N_46345,N_45883,N_45585);
and U46346 (N_46346,N_45678,N_45858);
nand U46347 (N_46347,N_45818,N_45878);
nor U46348 (N_46348,N_45665,N_45956);
xor U46349 (N_46349,N_45991,N_45628);
nand U46350 (N_46350,N_45649,N_45590);
nand U46351 (N_46351,N_45560,N_45691);
or U46352 (N_46352,N_45926,N_45778);
nor U46353 (N_46353,N_45607,N_45830);
or U46354 (N_46354,N_45868,N_45919);
xnor U46355 (N_46355,N_45515,N_45998);
nor U46356 (N_46356,N_45841,N_45875);
or U46357 (N_46357,N_45825,N_45677);
nand U46358 (N_46358,N_45783,N_45945);
or U46359 (N_46359,N_45910,N_45647);
nand U46360 (N_46360,N_45627,N_45721);
nor U46361 (N_46361,N_45545,N_45826);
and U46362 (N_46362,N_45728,N_45553);
or U46363 (N_46363,N_45593,N_45765);
nand U46364 (N_46364,N_45645,N_45944);
or U46365 (N_46365,N_45790,N_45972);
and U46366 (N_46366,N_45818,N_45904);
and U46367 (N_46367,N_45858,N_45772);
and U46368 (N_46368,N_45660,N_45936);
nand U46369 (N_46369,N_45580,N_45944);
and U46370 (N_46370,N_45677,N_45890);
xor U46371 (N_46371,N_45949,N_45504);
xor U46372 (N_46372,N_45736,N_45716);
nor U46373 (N_46373,N_45742,N_45628);
nand U46374 (N_46374,N_45526,N_45675);
and U46375 (N_46375,N_45947,N_45627);
xor U46376 (N_46376,N_45869,N_45651);
xor U46377 (N_46377,N_45839,N_45697);
xnor U46378 (N_46378,N_45838,N_45902);
xnor U46379 (N_46379,N_45626,N_45546);
nand U46380 (N_46380,N_45761,N_45877);
nand U46381 (N_46381,N_45743,N_45777);
nand U46382 (N_46382,N_45661,N_45931);
or U46383 (N_46383,N_45708,N_45634);
or U46384 (N_46384,N_45699,N_45825);
or U46385 (N_46385,N_45589,N_45978);
or U46386 (N_46386,N_45834,N_45784);
and U46387 (N_46387,N_45915,N_45801);
nand U46388 (N_46388,N_45996,N_45962);
xor U46389 (N_46389,N_45756,N_45758);
and U46390 (N_46390,N_45736,N_45801);
nand U46391 (N_46391,N_45792,N_45648);
and U46392 (N_46392,N_45918,N_45543);
or U46393 (N_46393,N_45782,N_45625);
and U46394 (N_46394,N_45777,N_45955);
xnor U46395 (N_46395,N_45782,N_45951);
and U46396 (N_46396,N_45960,N_45655);
nand U46397 (N_46397,N_45740,N_45612);
nand U46398 (N_46398,N_45957,N_45563);
xor U46399 (N_46399,N_45863,N_45798);
or U46400 (N_46400,N_45564,N_45962);
or U46401 (N_46401,N_45911,N_45584);
and U46402 (N_46402,N_45588,N_45626);
or U46403 (N_46403,N_45516,N_45730);
nand U46404 (N_46404,N_45663,N_45596);
xor U46405 (N_46405,N_45501,N_45730);
or U46406 (N_46406,N_45939,N_45819);
and U46407 (N_46407,N_45542,N_45804);
or U46408 (N_46408,N_45886,N_45766);
and U46409 (N_46409,N_45643,N_45531);
xor U46410 (N_46410,N_45711,N_45781);
or U46411 (N_46411,N_45611,N_45865);
or U46412 (N_46412,N_45808,N_45872);
and U46413 (N_46413,N_45966,N_45537);
and U46414 (N_46414,N_45986,N_45551);
or U46415 (N_46415,N_45806,N_45972);
and U46416 (N_46416,N_45996,N_45528);
and U46417 (N_46417,N_45621,N_45586);
or U46418 (N_46418,N_45517,N_45759);
nor U46419 (N_46419,N_45576,N_45503);
xnor U46420 (N_46420,N_45568,N_45649);
nand U46421 (N_46421,N_45724,N_45747);
xor U46422 (N_46422,N_45907,N_45690);
and U46423 (N_46423,N_45895,N_45692);
xor U46424 (N_46424,N_45523,N_45733);
nand U46425 (N_46425,N_45808,N_45543);
nand U46426 (N_46426,N_45812,N_45866);
nand U46427 (N_46427,N_45796,N_45537);
nor U46428 (N_46428,N_45732,N_45731);
or U46429 (N_46429,N_45809,N_45535);
or U46430 (N_46430,N_45575,N_45799);
or U46431 (N_46431,N_45564,N_45704);
and U46432 (N_46432,N_45518,N_45858);
nor U46433 (N_46433,N_45928,N_45743);
and U46434 (N_46434,N_45822,N_45847);
nand U46435 (N_46435,N_45814,N_45970);
and U46436 (N_46436,N_45746,N_45562);
and U46437 (N_46437,N_45899,N_45837);
and U46438 (N_46438,N_45697,N_45792);
and U46439 (N_46439,N_45688,N_45542);
nor U46440 (N_46440,N_45602,N_45797);
or U46441 (N_46441,N_45599,N_45693);
xor U46442 (N_46442,N_45549,N_45829);
nor U46443 (N_46443,N_45860,N_45632);
nand U46444 (N_46444,N_45836,N_45918);
nand U46445 (N_46445,N_45558,N_45512);
xor U46446 (N_46446,N_45673,N_45577);
nor U46447 (N_46447,N_45847,N_45756);
xnor U46448 (N_46448,N_45637,N_45880);
xnor U46449 (N_46449,N_45697,N_45932);
and U46450 (N_46450,N_45895,N_45885);
xor U46451 (N_46451,N_45747,N_45532);
and U46452 (N_46452,N_45840,N_45930);
nor U46453 (N_46453,N_45697,N_45639);
and U46454 (N_46454,N_45626,N_45631);
nand U46455 (N_46455,N_45643,N_45875);
xnor U46456 (N_46456,N_45916,N_45519);
nand U46457 (N_46457,N_45850,N_45986);
nor U46458 (N_46458,N_45932,N_45755);
nor U46459 (N_46459,N_45940,N_45900);
and U46460 (N_46460,N_45701,N_45900);
or U46461 (N_46461,N_45805,N_45840);
nor U46462 (N_46462,N_45928,N_45864);
or U46463 (N_46463,N_45710,N_45645);
xor U46464 (N_46464,N_45500,N_45612);
nor U46465 (N_46465,N_45707,N_45898);
xor U46466 (N_46466,N_45996,N_45779);
and U46467 (N_46467,N_45576,N_45568);
nor U46468 (N_46468,N_45591,N_45840);
nor U46469 (N_46469,N_45940,N_45567);
xnor U46470 (N_46470,N_45532,N_45984);
and U46471 (N_46471,N_45836,N_45652);
xor U46472 (N_46472,N_45824,N_45529);
and U46473 (N_46473,N_45781,N_45600);
or U46474 (N_46474,N_45843,N_45828);
or U46475 (N_46475,N_45531,N_45663);
nand U46476 (N_46476,N_45626,N_45761);
and U46477 (N_46477,N_45875,N_45898);
nand U46478 (N_46478,N_45963,N_45719);
xor U46479 (N_46479,N_45701,N_45876);
or U46480 (N_46480,N_45564,N_45836);
xnor U46481 (N_46481,N_45926,N_45546);
nor U46482 (N_46482,N_45541,N_45846);
and U46483 (N_46483,N_45657,N_45806);
nand U46484 (N_46484,N_45560,N_45819);
xor U46485 (N_46485,N_45703,N_45778);
xnor U46486 (N_46486,N_45524,N_45642);
xor U46487 (N_46487,N_45883,N_45852);
and U46488 (N_46488,N_45626,N_45872);
nand U46489 (N_46489,N_45736,N_45831);
nor U46490 (N_46490,N_45556,N_45698);
nor U46491 (N_46491,N_45875,N_45974);
or U46492 (N_46492,N_45954,N_45552);
or U46493 (N_46493,N_45631,N_45824);
or U46494 (N_46494,N_45930,N_45650);
xor U46495 (N_46495,N_45872,N_45926);
nand U46496 (N_46496,N_45965,N_45503);
xnor U46497 (N_46497,N_45824,N_45581);
xnor U46498 (N_46498,N_45815,N_45954);
nand U46499 (N_46499,N_45704,N_45976);
nor U46500 (N_46500,N_46393,N_46273);
xor U46501 (N_46501,N_46223,N_46143);
or U46502 (N_46502,N_46050,N_46421);
nand U46503 (N_46503,N_46458,N_46205);
xnor U46504 (N_46504,N_46460,N_46031);
nand U46505 (N_46505,N_46170,N_46336);
nand U46506 (N_46506,N_46209,N_46203);
nor U46507 (N_46507,N_46395,N_46478);
nand U46508 (N_46508,N_46383,N_46037);
and U46509 (N_46509,N_46448,N_46069);
and U46510 (N_46510,N_46285,N_46319);
or U46511 (N_46511,N_46021,N_46218);
and U46512 (N_46512,N_46434,N_46369);
and U46513 (N_46513,N_46374,N_46229);
nand U46514 (N_46514,N_46049,N_46165);
nor U46515 (N_46515,N_46488,N_46217);
nor U46516 (N_46516,N_46116,N_46292);
nor U46517 (N_46517,N_46061,N_46423);
and U46518 (N_46518,N_46122,N_46243);
or U46519 (N_46519,N_46459,N_46269);
or U46520 (N_46520,N_46462,N_46175);
or U46521 (N_46521,N_46258,N_46083);
nand U46522 (N_46522,N_46246,N_46178);
or U46523 (N_46523,N_46358,N_46142);
or U46524 (N_46524,N_46315,N_46445);
nand U46525 (N_46525,N_46343,N_46044);
nor U46526 (N_46526,N_46120,N_46264);
nor U46527 (N_46527,N_46291,N_46431);
or U46528 (N_46528,N_46360,N_46411);
and U46529 (N_46529,N_46361,N_46414);
xor U46530 (N_46530,N_46412,N_46146);
xor U46531 (N_46531,N_46331,N_46215);
nand U46532 (N_46532,N_46059,N_46039);
nand U46533 (N_46533,N_46224,N_46316);
and U46534 (N_46534,N_46125,N_46276);
nand U46535 (N_46535,N_46441,N_46477);
and U46536 (N_46536,N_46326,N_46359);
nor U46537 (N_46537,N_46232,N_46317);
and U46538 (N_46538,N_46440,N_46363);
xor U46539 (N_46539,N_46072,N_46156);
or U46540 (N_46540,N_46446,N_46334);
or U46541 (N_46541,N_46192,N_46227);
xor U46542 (N_46542,N_46228,N_46046);
or U46543 (N_46543,N_46389,N_46490);
and U46544 (N_46544,N_46025,N_46270);
xnor U46545 (N_46545,N_46475,N_46275);
nor U46546 (N_46546,N_46307,N_46036);
xor U46547 (N_46547,N_46309,N_46417);
and U46548 (N_46548,N_46087,N_46499);
or U46549 (N_46549,N_46098,N_46457);
nand U46550 (N_46550,N_46282,N_46381);
or U46551 (N_46551,N_46140,N_46211);
or U46552 (N_46552,N_46076,N_46378);
and U46553 (N_46553,N_46220,N_46126);
nor U46554 (N_46554,N_46057,N_46029);
xor U46555 (N_46555,N_46396,N_46377);
nand U46556 (N_46556,N_46207,N_46109);
nand U46557 (N_46557,N_46151,N_46265);
xor U46558 (N_46558,N_46053,N_46296);
and U46559 (N_46559,N_46012,N_46158);
and U46560 (N_46560,N_46118,N_46193);
nor U46561 (N_46561,N_46268,N_46281);
and U46562 (N_46562,N_46333,N_46108);
nand U46563 (N_46563,N_46052,N_46245);
nor U46564 (N_46564,N_46148,N_46006);
and U46565 (N_46565,N_46495,N_46356);
nor U46566 (N_46566,N_46386,N_46241);
nand U46567 (N_46567,N_46035,N_46274);
xor U46568 (N_46568,N_46324,N_46144);
nor U46569 (N_46569,N_46267,N_46402);
and U46570 (N_46570,N_46321,N_46255);
xor U46571 (N_46571,N_46043,N_46107);
nand U46572 (N_46572,N_46106,N_46119);
or U46573 (N_46573,N_46272,N_46452);
nor U46574 (N_46574,N_46449,N_46304);
nand U46575 (N_46575,N_46095,N_46048);
nand U46576 (N_46576,N_46425,N_46420);
or U46577 (N_46577,N_46435,N_46182);
and U46578 (N_46578,N_46014,N_46342);
or U46579 (N_46579,N_46391,N_46066);
nand U46580 (N_46580,N_46300,N_46055);
nand U46581 (N_46581,N_46100,N_46468);
or U46582 (N_46582,N_46442,N_46212);
nand U46583 (N_46583,N_46338,N_46152);
and U46584 (N_46584,N_46432,N_46104);
nor U46585 (N_46585,N_46181,N_46487);
xnor U46586 (N_46586,N_46250,N_46426);
or U46587 (N_46587,N_46210,N_46470);
xnor U46588 (N_46588,N_46347,N_46465);
xnor U46589 (N_46589,N_46485,N_46473);
or U46590 (N_46590,N_46011,N_46026);
or U46591 (N_46591,N_46266,N_46362);
xor U46592 (N_46592,N_46045,N_46413);
nor U46593 (N_46593,N_46332,N_46160);
xnor U46594 (N_46594,N_46350,N_46262);
or U46595 (N_46595,N_46354,N_46364);
and U46596 (N_46596,N_46486,N_46074);
or U46597 (N_46597,N_46213,N_46190);
and U46598 (N_46598,N_46252,N_46344);
nand U46599 (N_46599,N_46009,N_46271);
nor U46600 (N_46600,N_46088,N_46008);
nor U46601 (N_46601,N_46180,N_46173);
and U46602 (N_46602,N_46123,N_46498);
or U46603 (N_46603,N_46279,N_46060);
or U46604 (N_46604,N_46138,N_46067);
nor U46605 (N_46605,N_46091,N_46474);
nand U46606 (N_46606,N_46287,N_46234);
xnor U46607 (N_46607,N_46018,N_46439);
nor U46608 (N_46608,N_46041,N_46171);
xnor U46609 (N_46609,N_46139,N_46033);
or U46610 (N_46610,N_46201,N_46032);
and U46611 (N_46611,N_46040,N_46424);
nand U46612 (N_46612,N_46284,N_46303);
and U46613 (N_46613,N_46065,N_46134);
and U46614 (N_46614,N_46376,N_46038);
and U46615 (N_46615,N_46349,N_46368);
or U46616 (N_46616,N_46236,N_46231);
or U46617 (N_46617,N_46382,N_46208);
or U46618 (N_46618,N_46403,N_46308);
and U46619 (N_46619,N_46051,N_46010);
nand U46620 (N_46620,N_46169,N_46071);
nor U46621 (N_46621,N_46103,N_46384);
nor U46622 (N_46622,N_46482,N_46249);
and U46623 (N_46623,N_46070,N_46323);
xnor U46624 (N_46624,N_46017,N_46114);
and U46625 (N_46625,N_46493,N_46244);
and U46626 (N_46626,N_46277,N_46313);
or U46627 (N_46627,N_46145,N_46310);
nor U46628 (N_46628,N_46484,N_46199);
and U46629 (N_46629,N_46093,N_46078);
and U46630 (N_46630,N_46312,N_46251);
nand U46631 (N_46631,N_46352,N_46022);
or U46632 (N_46632,N_46188,N_46124);
nand U46633 (N_46633,N_46204,N_46082);
or U46634 (N_46634,N_46075,N_46121);
xnor U46635 (N_46635,N_46427,N_46339);
nand U46636 (N_46636,N_46128,N_46177);
nor U46637 (N_46637,N_46016,N_46187);
and U46638 (N_46638,N_46328,N_46346);
nor U46639 (N_46639,N_46283,N_46235);
or U46640 (N_46640,N_46030,N_46133);
nor U46641 (N_46641,N_46102,N_46240);
nor U46642 (N_46642,N_46410,N_46259);
or U46643 (N_46643,N_46409,N_46365);
xnor U46644 (N_46644,N_46353,N_46254);
nor U46645 (N_46645,N_46163,N_46115);
xor U46646 (N_46646,N_46341,N_46099);
nand U46647 (N_46647,N_46166,N_46454);
nand U46648 (N_46648,N_46174,N_46295);
and U46649 (N_46649,N_46222,N_46216);
xor U46650 (N_46650,N_46392,N_46325);
or U46651 (N_46651,N_46497,N_46297);
or U46652 (N_46652,N_46371,N_46164);
and U46653 (N_46653,N_46127,N_46194);
or U46654 (N_46654,N_46429,N_46068);
nand U46655 (N_46655,N_46430,N_46094);
nand U46656 (N_46656,N_46172,N_46206);
nand U46657 (N_46657,N_46280,N_46388);
xor U46658 (N_46658,N_46257,N_46253);
or U46659 (N_46659,N_46379,N_46340);
xor U46660 (N_46660,N_46327,N_46130);
nand U46661 (N_46661,N_46237,N_46000);
nand U46662 (N_46662,N_46183,N_46461);
xnor U46663 (N_46663,N_46176,N_46318);
xor U46664 (N_46664,N_46408,N_46097);
nor U46665 (N_46665,N_46219,N_46242);
nand U46666 (N_46666,N_46054,N_46117);
nor U46667 (N_46667,N_46444,N_46191);
and U46668 (N_46668,N_46004,N_46112);
nor U46669 (N_46669,N_46136,N_46469);
nor U46670 (N_46670,N_46195,N_46404);
xor U46671 (N_46671,N_46034,N_46479);
nand U46672 (N_46672,N_46418,N_46380);
xor U46673 (N_46673,N_46080,N_46185);
nor U46674 (N_46674,N_46320,N_46355);
or U46675 (N_46675,N_46020,N_46314);
and U46676 (N_46676,N_46263,N_46483);
nor U46677 (N_46677,N_46101,N_46077);
or U46678 (N_46678,N_46301,N_46401);
xor U46679 (N_46679,N_46394,N_46003);
and U46680 (N_46680,N_46290,N_46463);
xor U46681 (N_46681,N_46063,N_46436);
nor U46682 (N_46682,N_46248,N_46278);
and U46683 (N_46683,N_46196,N_46351);
nand U46684 (N_46684,N_46005,N_46400);
xor U46685 (N_46685,N_46288,N_46225);
xor U46686 (N_46686,N_46451,N_46289);
nand U46687 (N_46687,N_46042,N_46491);
xor U46688 (N_46688,N_46357,N_46397);
and U46689 (N_46689,N_46024,N_46084);
xor U46690 (N_46690,N_46154,N_46155);
nand U46691 (N_46691,N_46387,N_46492);
nor U46692 (N_46692,N_46322,N_46073);
and U46693 (N_46693,N_46019,N_46481);
and U46694 (N_46694,N_46226,N_46367);
or U46695 (N_46695,N_46476,N_46161);
nor U46696 (N_46696,N_46023,N_46375);
or U46697 (N_46697,N_46455,N_46111);
and U46698 (N_46698,N_46132,N_46416);
nor U46699 (N_46699,N_46447,N_46214);
nand U46700 (N_46700,N_46147,N_46399);
nor U46701 (N_46701,N_46390,N_46233);
and U46702 (N_46702,N_46489,N_46348);
nor U46703 (N_46703,N_46256,N_46096);
nor U46704 (N_46704,N_46089,N_46141);
nand U46705 (N_46705,N_46415,N_46081);
and U46706 (N_46706,N_46467,N_46085);
nor U46707 (N_46707,N_46238,N_46001);
and U46708 (N_46708,N_46406,N_46179);
nor U46709 (N_46709,N_46433,N_46189);
or U46710 (N_46710,N_46456,N_46305);
or U46711 (N_46711,N_46157,N_46330);
nand U46712 (N_46712,N_46239,N_46137);
and U46713 (N_46713,N_46472,N_46370);
xnor U46714 (N_46714,N_46013,N_46015);
and U46715 (N_46715,N_46329,N_46221);
and U46716 (N_46716,N_46202,N_46064);
and U46717 (N_46717,N_46129,N_46466);
and U46718 (N_46718,N_46230,N_46131);
nand U46719 (N_46719,N_46294,N_46480);
or U46720 (N_46720,N_46198,N_46047);
or U46721 (N_46721,N_46437,N_46366);
xor U46722 (N_46722,N_46247,N_46135);
nand U46723 (N_46723,N_46186,N_46405);
nor U46724 (N_46724,N_46335,N_46496);
xor U46725 (N_46725,N_46153,N_46113);
and U46726 (N_46726,N_46260,N_46105);
xnor U46727 (N_46727,N_46398,N_46345);
and U46728 (N_46728,N_46028,N_46419);
xor U46729 (N_46729,N_46007,N_46197);
nor U46730 (N_46730,N_46162,N_46428);
and U46731 (N_46731,N_46200,N_46407);
nor U46732 (N_46732,N_46337,N_46090);
xor U46733 (N_46733,N_46438,N_46471);
nor U46734 (N_46734,N_46002,N_46306);
or U46735 (N_46735,N_46149,N_46453);
or U46736 (N_46736,N_46027,N_46056);
nand U46737 (N_46737,N_46373,N_46494);
nor U46738 (N_46738,N_46150,N_46062);
xnor U46739 (N_46739,N_46311,N_46184);
and U46740 (N_46740,N_46464,N_46299);
nor U46741 (N_46741,N_46159,N_46422);
nor U46742 (N_46742,N_46372,N_46058);
nand U46743 (N_46743,N_46302,N_46079);
nand U46744 (N_46744,N_46450,N_46286);
and U46745 (N_46745,N_46086,N_46168);
nor U46746 (N_46746,N_46092,N_46261);
xnor U46747 (N_46747,N_46167,N_46385);
or U46748 (N_46748,N_46293,N_46298);
nand U46749 (N_46749,N_46443,N_46110);
and U46750 (N_46750,N_46205,N_46360);
nor U46751 (N_46751,N_46305,N_46201);
nor U46752 (N_46752,N_46236,N_46385);
xnor U46753 (N_46753,N_46101,N_46386);
nand U46754 (N_46754,N_46315,N_46451);
nand U46755 (N_46755,N_46292,N_46433);
or U46756 (N_46756,N_46187,N_46253);
xor U46757 (N_46757,N_46399,N_46455);
nor U46758 (N_46758,N_46075,N_46007);
nor U46759 (N_46759,N_46260,N_46154);
or U46760 (N_46760,N_46462,N_46487);
and U46761 (N_46761,N_46365,N_46056);
and U46762 (N_46762,N_46460,N_46002);
nand U46763 (N_46763,N_46028,N_46242);
nor U46764 (N_46764,N_46008,N_46090);
xor U46765 (N_46765,N_46425,N_46496);
and U46766 (N_46766,N_46068,N_46099);
nor U46767 (N_46767,N_46482,N_46195);
xor U46768 (N_46768,N_46035,N_46284);
nor U46769 (N_46769,N_46358,N_46250);
nand U46770 (N_46770,N_46436,N_46374);
xor U46771 (N_46771,N_46393,N_46289);
or U46772 (N_46772,N_46450,N_46289);
xnor U46773 (N_46773,N_46425,N_46171);
or U46774 (N_46774,N_46420,N_46486);
nor U46775 (N_46775,N_46392,N_46005);
or U46776 (N_46776,N_46380,N_46319);
xor U46777 (N_46777,N_46263,N_46298);
or U46778 (N_46778,N_46032,N_46021);
xor U46779 (N_46779,N_46136,N_46371);
xnor U46780 (N_46780,N_46132,N_46287);
xnor U46781 (N_46781,N_46160,N_46268);
nand U46782 (N_46782,N_46127,N_46368);
and U46783 (N_46783,N_46238,N_46365);
nor U46784 (N_46784,N_46162,N_46493);
and U46785 (N_46785,N_46380,N_46318);
or U46786 (N_46786,N_46238,N_46348);
nor U46787 (N_46787,N_46234,N_46105);
xor U46788 (N_46788,N_46076,N_46018);
xor U46789 (N_46789,N_46294,N_46216);
xnor U46790 (N_46790,N_46301,N_46052);
nand U46791 (N_46791,N_46147,N_46382);
nor U46792 (N_46792,N_46274,N_46232);
nand U46793 (N_46793,N_46300,N_46278);
and U46794 (N_46794,N_46241,N_46073);
xor U46795 (N_46795,N_46137,N_46445);
xnor U46796 (N_46796,N_46241,N_46425);
and U46797 (N_46797,N_46124,N_46217);
xnor U46798 (N_46798,N_46099,N_46345);
or U46799 (N_46799,N_46335,N_46087);
nor U46800 (N_46800,N_46239,N_46153);
or U46801 (N_46801,N_46228,N_46175);
nor U46802 (N_46802,N_46288,N_46469);
or U46803 (N_46803,N_46019,N_46208);
or U46804 (N_46804,N_46129,N_46433);
nand U46805 (N_46805,N_46029,N_46079);
nand U46806 (N_46806,N_46365,N_46126);
and U46807 (N_46807,N_46316,N_46471);
and U46808 (N_46808,N_46346,N_46417);
nand U46809 (N_46809,N_46023,N_46097);
xnor U46810 (N_46810,N_46048,N_46297);
nor U46811 (N_46811,N_46112,N_46013);
or U46812 (N_46812,N_46153,N_46059);
and U46813 (N_46813,N_46381,N_46488);
nand U46814 (N_46814,N_46302,N_46387);
and U46815 (N_46815,N_46314,N_46471);
and U46816 (N_46816,N_46331,N_46381);
or U46817 (N_46817,N_46080,N_46274);
and U46818 (N_46818,N_46105,N_46330);
and U46819 (N_46819,N_46345,N_46402);
nand U46820 (N_46820,N_46405,N_46480);
and U46821 (N_46821,N_46354,N_46112);
or U46822 (N_46822,N_46404,N_46220);
nand U46823 (N_46823,N_46189,N_46159);
nor U46824 (N_46824,N_46010,N_46401);
xor U46825 (N_46825,N_46113,N_46173);
nor U46826 (N_46826,N_46345,N_46095);
xor U46827 (N_46827,N_46116,N_46246);
xnor U46828 (N_46828,N_46311,N_46407);
nand U46829 (N_46829,N_46152,N_46403);
nand U46830 (N_46830,N_46104,N_46158);
nand U46831 (N_46831,N_46471,N_46228);
nand U46832 (N_46832,N_46038,N_46100);
nor U46833 (N_46833,N_46258,N_46404);
nand U46834 (N_46834,N_46184,N_46344);
and U46835 (N_46835,N_46466,N_46211);
xor U46836 (N_46836,N_46239,N_46408);
or U46837 (N_46837,N_46344,N_46229);
xor U46838 (N_46838,N_46182,N_46397);
xnor U46839 (N_46839,N_46368,N_46048);
or U46840 (N_46840,N_46428,N_46054);
nand U46841 (N_46841,N_46309,N_46439);
or U46842 (N_46842,N_46045,N_46242);
xor U46843 (N_46843,N_46268,N_46006);
nand U46844 (N_46844,N_46387,N_46197);
nor U46845 (N_46845,N_46019,N_46199);
nand U46846 (N_46846,N_46029,N_46091);
nor U46847 (N_46847,N_46371,N_46063);
and U46848 (N_46848,N_46048,N_46121);
nor U46849 (N_46849,N_46091,N_46057);
nand U46850 (N_46850,N_46065,N_46489);
xor U46851 (N_46851,N_46430,N_46021);
and U46852 (N_46852,N_46084,N_46192);
nor U46853 (N_46853,N_46109,N_46446);
and U46854 (N_46854,N_46206,N_46164);
nand U46855 (N_46855,N_46493,N_46429);
nand U46856 (N_46856,N_46143,N_46491);
xnor U46857 (N_46857,N_46310,N_46432);
and U46858 (N_46858,N_46128,N_46129);
and U46859 (N_46859,N_46121,N_46028);
xor U46860 (N_46860,N_46491,N_46098);
or U46861 (N_46861,N_46421,N_46404);
xor U46862 (N_46862,N_46231,N_46438);
nand U46863 (N_46863,N_46105,N_46398);
and U46864 (N_46864,N_46076,N_46380);
nand U46865 (N_46865,N_46322,N_46385);
or U46866 (N_46866,N_46152,N_46333);
xor U46867 (N_46867,N_46034,N_46052);
xnor U46868 (N_46868,N_46145,N_46072);
or U46869 (N_46869,N_46093,N_46077);
and U46870 (N_46870,N_46175,N_46182);
xor U46871 (N_46871,N_46082,N_46487);
or U46872 (N_46872,N_46088,N_46076);
or U46873 (N_46873,N_46356,N_46110);
xnor U46874 (N_46874,N_46151,N_46267);
xnor U46875 (N_46875,N_46341,N_46209);
nor U46876 (N_46876,N_46039,N_46007);
nand U46877 (N_46877,N_46164,N_46297);
nand U46878 (N_46878,N_46400,N_46000);
or U46879 (N_46879,N_46336,N_46167);
nand U46880 (N_46880,N_46224,N_46416);
nor U46881 (N_46881,N_46456,N_46317);
nand U46882 (N_46882,N_46477,N_46412);
nand U46883 (N_46883,N_46095,N_46435);
nand U46884 (N_46884,N_46000,N_46012);
and U46885 (N_46885,N_46053,N_46320);
nor U46886 (N_46886,N_46376,N_46102);
or U46887 (N_46887,N_46086,N_46284);
nand U46888 (N_46888,N_46042,N_46062);
nand U46889 (N_46889,N_46161,N_46368);
nor U46890 (N_46890,N_46015,N_46308);
nor U46891 (N_46891,N_46323,N_46374);
and U46892 (N_46892,N_46382,N_46381);
and U46893 (N_46893,N_46083,N_46228);
xnor U46894 (N_46894,N_46020,N_46138);
nand U46895 (N_46895,N_46498,N_46065);
xor U46896 (N_46896,N_46411,N_46221);
and U46897 (N_46897,N_46056,N_46344);
xnor U46898 (N_46898,N_46125,N_46116);
or U46899 (N_46899,N_46219,N_46323);
or U46900 (N_46900,N_46075,N_46107);
xnor U46901 (N_46901,N_46186,N_46084);
xor U46902 (N_46902,N_46165,N_46464);
xor U46903 (N_46903,N_46118,N_46286);
xnor U46904 (N_46904,N_46408,N_46310);
nand U46905 (N_46905,N_46232,N_46055);
or U46906 (N_46906,N_46395,N_46317);
and U46907 (N_46907,N_46293,N_46134);
and U46908 (N_46908,N_46342,N_46008);
nand U46909 (N_46909,N_46192,N_46101);
or U46910 (N_46910,N_46435,N_46446);
or U46911 (N_46911,N_46365,N_46156);
and U46912 (N_46912,N_46296,N_46337);
or U46913 (N_46913,N_46155,N_46125);
nor U46914 (N_46914,N_46104,N_46120);
nor U46915 (N_46915,N_46093,N_46218);
nor U46916 (N_46916,N_46300,N_46423);
and U46917 (N_46917,N_46494,N_46336);
nor U46918 (N_46918,N_46142,N_46486);
or U46919 (N_46919,N_46135,N_46150);
xnor U46920 (N_46920,N_46188,N_46288);
xor U46921 (N_46921,N_46070,N_46197);
nor U46922 (N_46922,N_46441,N_46037);
xor U46923 (N_46923,N_46285,N_46476);
and U46924 (N_46924,N_46003,N_46396);
and U46925 (N_46925,N_46018,N_46427);
or U46926 (N_46926,N_46015,N_46455);
nand U46927 (N_46927,N_46223,N_46406);
xor U46928 (N_46928,N_46463,N_46398);
nor U46929 (N_46929,N_46171,N_46351);
and U46930 (N_46930,N_46423,N_46406);
xor U46931 (N_46931,N_46430,N_46066);
nand U46932 (N_46932,N_46088,N_46033);
nand U46933 (N_46933,N_46068,N_46284);
or U46934 (N_46934,N_46061,N_46414);
or U46935 (N_46935,N_46023,N_46417);
and U46936 (N_46936,N_46466,N_46353);
nand U46937 (N_46937,N_46347,N_46325);
and U46938 (N_46938,N_46337,N_46009);
xnor U46939 (N_46939,N_46404,N_46086);
nor U46940 (N_46940,N_46058,N_46343);
and U46941 (N_46941,N_46495,N_46322);
and U46942 (N_46942,N_46055,N_46246);
nor U46943 (N_46943,N_46179,N_46234);
nand U46944 (N_46944,N_46298,N_46481);
xnor U46945 (N_46945,N_46117,N_46109);
nor U46946 (N_46946,N_46285,N_46420);
or U46947 (N_46947,N_46199,N_46052);
nand U46948 (N_46948,N_46001,N_46050);
xor U46949 (N_46949,N_46480,N_46291);
and U46950 (N_46950,N_46067,N_46050);
or U46951 (N_46951,N_46381,N_46304);
nand U46952 (N_46952,N_46381,N_46245);
or U46953 (N_46953,N_46279,N_46187);
and U46954 (N_46954,N_46101,N_46157);
nand U46955 (N_46955,N_46498,N_46192);
or U46956 (N_46956,N_46214,N_46262);
nand U46957 (N_46957,N_46226,N_46026);
and U46958 (N_46958,N_46335,N_46264);
or U46959 (N_46959,N_46015,N_46386);
xnor U46960 (N_46960,N_46398,N_46371);
or U46961 (N_46961,N_46357,N_46406);
or U46962 (N_46962,N_46134,N_46328);
nand U46963 (N_46963,N_46205,N_46300);
and U46964 (N_46964,N_46488,N_46218);
nor U46965 (N_46965,N_46431,N_46464);
nor U46966 (N_46966,N_46240,N_46022);
or U46967 (N_46967,N_46356,N_46153);
nand U46968 (N_46968,N_46191,N_46280);
xnor U46969 (N_46969,N_46238,N_46029);
and U46970 (N_46970,N_46428,N_46292);
and U46971 (N_46971,N_46294,N_46164);
nand U46972 (N_46972,N_46114,N_46231);
nor U46973 (N_46973,N_46148,N_46342);
nand U46974 (N_46974,N_46348,N_46391);
or U46975 (N_46975,N_46154,N_46199);
or U46976 (N_46976,N_46349,N_46473);
nand U46977 (N_46977,N_46282,N_46167);
or U46978 (N_46978,N_46128,N_46240);
or U46979 (N_46979,N_46314,N_46201);
xnor U46980 (N_46980,N_46300,N_46287);
xor U46981 (N_46981,N_46233,N_46014);
and U46982 (N_46982,N_46094,N_46368);
and U46983 (N_46983,N_46370,N_46170);
nand U46984 (N_46984,N_46439,N_46206);
nand U46985 (N_46985,N_46441,N_46348);
nor U46986 (N_46986,N_46086,N_46438);
and U46987 (N_46987,N_46064,N_46075);
or U46988 (N_46988,N_46369,N_46021);
and U46989 (N_46989,N_46493,N_46378);
nor U46990 (N_46990,N_46326,N_46342);
xor U46991 (N_46991,N_46497,N_46247);
nand U46992 (N_46992,N_46498,N_46199);
xor U46993 (N_46993,N_46119,N_46370);
nor U46994 (N_46994,N_46342,N_46017);
and U46995 (N_46995,N_46216,N_46282);
nand U46996 (N_46996,N_46263,N_46183);
xnor U46997 (N_46997,N_46293,N_46056);
and U46998 (N_46998,N_46298,N_46418);
nor U46999 (N_46999,N_46176,N_46055);
xnor U47000 (N_47000,N_46548,N_46511);
nand U47001 (N_47001,N_46736,N_46561);
xor U47002 (N_47002,N_46546,N_46934);
nand U47003 (N_47003,N_46635,N_46835);
or U47004 (N_47004,N_46792,N_46952);
nor U47005 (N_47005,N_46570,N_46790);
xor U47006 (N_47006,N_46622,N_46559);
nand U47007 (N_47007,N_46823,N_46647);
nand U47008 (N_47008,N_46667,N_46637);
and U47009 (N_47009,N_46735,N_46911);
nor U47010 (N_47010,N_46687,N_46756);
nor U47011 (N_47011,N_46646,N_46603);
nand U47012 (N_47012,N_46560,N_46761);
xor U47013 (N_47013,N_46581,N_46827);
or U47014 (N_47014,N_46583,N_46942);
nor U47015 (N_47015,N_46946,N_46696);
and U47016 (N_47016,N_46973,N_46662);
or U47017 (N_47017,N_46732,N_46728);
xor U47018 (N_47018,N_46650,N_46562);
or U47019 (N_47019,N_46563,N_46680);
xor U47020 (N_47020,N_46980,N_46709);
xnor U47021 (N_47021,N_46584,N_46975);
xnor U47022 (N_47022,N_46956,N_46825);
xor U47023 (N_47023,N_46982,N_46530);
nand U47024 (N_47024,N_46840,N_46710);
and U47025 (N_47025,N_46846,N_46886);
and U47026 (N_47026,N_46912,N_46829);
nand U47027 (N_47027,N_46895,N_46532);
and U47028 (N_47028,N_46970,N_46888);
nor U47029 (N_47029,N_46826,N_46990);
xor U47030 (N_47030,N_46595,N_46923);
nand U47031 (N_47031,N_46742,N_46638);
nor U47032 (N_47032,N_46882,N_46738);
or U47033 (N_47033,N_46705,N_46887);
or U47034 (N_47034,N_46612,N_46586);
and U47035 (N_47035,N_46995,N_46905);
xnor U47036 (N_47036,N_46865,N_46787);
or U47037 (N_47037,N_46971,N_46500);
nand U47038 (N_47038,N_46889,N_46831);
xor U47039 (N_47039,N_46566,N_46943);
xor U47040 (N_47040,N_46516,N_46931);
and U47041 (N_47041,N_46844,N_46610);
nand U47042 (N_47042,N_46978,N_46789);
or U47043 (N_47043,N_46645,N_46554);
nand U47044 (N_47044,N_46691,N_46820);
nand U47045 (N_47045,N_46655,N_46753);
and U47046 (N_47046,N_46556,N_46656);
nand U47047 (N_47047,N_46998,N_46620);
nand U47048 (N_47048,N_46513,N_46766);
and U47049 (N_47049,N_46737,N_46585);
or U47050 (N_47050,N_46918,N_46988);
and U47051 (N_47051,N_46676,N_46537);
and U47052 (N_47052,N_46621,N_46945);
and U47053 (N_47053,N_46576,N_46994);
nand U47054 (N_47054,N_46922,N_46900);
nand U47055 (N_47055,N_46692,N_46953);
nor U47056 (N_47056,N_46799,N_46929);
nand U47057 (N_47057,N_46701,N_46854);
or U47058 (N_47058,N_46526,N_46860);
xnor U47059 (N_47059,N_46949,N_46632);
xor U47060 (N_47060,N_46991,N_46925);
or U47061 (N_47061,N_46885,N_46781);
nand U47062 (N_47062,N_46883,N_46804);
nand U47063 (N_47063,N_46599,N_46947);
or U47064 (N_47064,N_46601,N_46718);
and U47065 (N_47065,N_46702,N_46876);
or U47066 (N_47066,N_46750,N_46745);
xor U47067 (N_47067,N_46573,N_46754);
or U47068 (N_47068,N_46981,N_46503);
and U47069 (N_47069,N_46594,N_46534);
or U47070 (N_47070,N_46941,N_46741);
or U47071 (N_47071,N_46915,N_46626);
nand U47072 (N_47072,N_46731,N_46760);
or U47073 (N_47073,N_46993,N_46510);
or U47074 (N_47074,N_46729,N_46514);
nor U47075 (N_47075,N_46613,N_46674);
nand U47076 (N_47076,N_46958,N_46877);
nor U47077 (N_47077,N_46747,N_46751);
xor U47078 (N_47078,N_46553,N_46608);
nand U47079 (N_47079,N_46961,N_46727);
nand U47080 (N_47080,N_46661,N_46932);
or U47081 (N_47081,N_46939,N_46814);
and U47082 (N_47082,N_46870,N_46572);
and U47083 (N_47083,N_46801,N_46706);
and U47084 (N_47084,N_46755,N_46868);
nand U47085 (N_47085,N_46630,N_46757);
or U47086 (N_47086,N_46588,N_46780);
or U47087 (N_47087,N_46640,N_46967);
or U47088 (N_47088,N_46904,N_46614);
xor U47089 (N_47089,N_46624,N_46596);
nand U47090 (N_47090,N_46808,N_46765);
nand U47091 (N_47091,N_46506,N_46507);
and U47092 (N_47092,N_46806,N_46502);
nand U47093 (N_47093,N_46693,N_46896);
or U47094 (N_47094,N_46903,N_46733);
and U47095 (N_47095,N_46714,N_46893);
xnor U47096 (N_47096,N_46522,N_46587);
or U47097 (N_47097,N_46545,N_46748);
nor U47098 (N_47098,N_46504,N_46558);
or U47099 (N_47099,N_46816,N_46824);
nor U47100 (N_47100,N_46660,N_46633);
nor U47101 (N_47101,N_46541,N_46786);
xnor U47102 (N_47102,N_46832,N_46670);
and U47103 (N_47103,N_46658,N_46724);
xnor U47104 (N_47104,N_46550,N_46858);
or U47105 (N_47105,N_46817,N_46564);
xnor U47106 (N_47106,N_46798,N_46579);
nand U47107 (N_47107,N_46683,N_46963);
nand U47108 (N_47108,N_46726,N_46589);
xor U47109 (N_47109,N_46521,N_46935);
and U47110 (N_47110,N_46773,N_46856);
or U47111 (N_47111,N_46851,N_46807);
or U47112 (N_47112,N_46833,N_46703);
xnor U47113 (N_47113,N_46697,N_46725);
nand U47114 (N_47114,N_46721,N_46763);
nand U47115 (N_47115,N_46892,N_46758);
xnor U47116 (N_47116,N_46857,N_46834);
or U47117 (N_47117,N_46966,N_46880);
and U47118 (N_47118,N_46713,N_46933);
nor U47119 (N_47119,N_46805,N_46776);
and U47120 (N_47120,N_46771,N_46782);
or U47121 (N_47121,N_46864,N_46591);
or U47122 (N_47122,N_46779,N_46715);
nor U47123 (N_47123,N_46636,N_46678);
or U47124 (N_47124,N_46759,N_46902);
nand U47125 (N_47125,N_46509,N_46657);
nor U47126 (N_47126,N_46879,N_46695);
nor U47127 (N_47127,N_46527,N_46672);
nand U47128 (N_47128,N_46623,N_46785);
nand U47129 (N_47129,N_46653,N_46850);
nand U47130 (N_47130,N_46688,N_46690);
or U47131 (N_47131,N_46539,N_46987);
nor U47132 (N_47132,N_46666,N_46772);
xor U47133 (N_47133,N_46954,N_46890);
nor U47134 (N_47134,N_46839,N_46938);
nor U47135 (N_47135,N_46796,N_46997);
and U47136 (N_47136,N_46959,N_46628);
nor U47137 (N_47137,N_46602,N_46853);
or U47138 (N_47138,N_46684,N_46862);
and U47139 (N_47139,N_46884,N_46871);
and U47140 (N_47140,N_46571,N_46616);
xor U47141 (N_47141,N_46767,N_46663);
nor U47142 (N_47142,N_46762,N_46968);
nand U47143 (N_47143,N_46659,N_46818);
nand U47144 (N_47144,N_46848,N_46768);
or U47145 (N_47145,N_46811,N_46924);
xnor U47146 (N_47146,N_46671,N_46783);
and U47147 (N_47147,N_46999,N_46567);
xor U47148 (N_47148,N_46664,N_46578);
nand U47149 (N_47149,N_46813,N_46605);
nand U47150 (N_47150,N_46979,N_46543);
and U47151 (N_47151,N_46752,N_46520);
and U47152 (N_47152,N_46836,N_46649);
nand U47153 (N_47153,N_46803,N_46845);
and U47154 (N_47154,N_46679,N_46770);
or U47155 (N_47155,N_46863,N_46764);
or U47156 (N_47156,N_46535,N_46704);
nand U47157 (N_47157,N_46569,N_46609);
or U47158 (N_47158,N_46866,N_46910);
nor U47159 (N_47159,N_46643,N_46686);
or U47160 (N_47160,N_46810,N_46574);
nor U47161 (N_47161,N_46575,N_46996);
xor U47162 (N_47162,N_46689,N_46617);
nor U47163 (N_47163,N_46847,N_46631);
nand U47164 (N_47164,N_46597,N_46897);
nand U47165 (N_47165,N_46694,N_46909);
xnor U47166 (N_47166,N_46878,N_46518);
nor U47167 (N_47167,N_46775,N_46791);
and U47168 (N_47168,N_46852,N_46699);
nand U47169 (N_47169,N_46627,N_46654);
or U47170 (N_47170,N_46673,N_46580);
nor U47171 (N_47171,N_46986,N_46730);
and U47172 (N_47172,N_46739,N_46809);
nand U47173 (N_47173,N_46914,N_46951);
nand U47174 (N_47174,N_46577,N_46606);
nor U47175 (N_47175,N_46965,N_46957);
nor U47176 (N_47176,N_46802,N_46716);
xnor U47177 (N_47177,N_46907,N_46920);
xor U47178 (N_47178,N_46743,N_46593);
nand U47179 (N_47179,N_46819,N_46874);
nor U47180 (N_47180,N_46960,N_46557);
xnor U47181 (N_47181,N_46749,N_46568);
or U47182 (N_47182,N_46642,N_46682);
and U47183 (N_47183,N_46841,N_46913);
xnor U47184 (N_47184,N_46669,N_46927);
or U47185 (N_47185,N_46707,N_46719);
nand U47186 (N_47186,N_46536,N_46875);
nor U47187 (N_47187,N_46969,N_46644);
nand U47188 (N_47188,N_46604,N_46618);
xor U47189 (N_47189,N_46919,N_46976);
nor U47190 (N_47190,N_46677,N_46740);
nor U47191 (N_47191,N_46734,N_46940);
nor U47192 (N_47192,N_46720,N_46598);
or U47193 (N_47193,N_46722,N_46505);
and U47194 (N_47194,N_46926,N_46843);
nor U47195 (N_47195,N_46812,N_46517);
nor U47196 (N_47196,N_46681,N_46600);
nand U47197 (N_47197,N_46652,N_46992);
and U47198 (N_47198,N_46512,N_46822);
nor U47199 (N_47199,N_46540,N_46744);
and U47200 (N_47200,N_46937,N_46711);
nand U47201 (N_47201,N_46977,N_46861);
nor U47202 (N_47202,N_46972,N_46592);
xnor U47203 (N_47203,N_46565,N_46778);
nor U47204 (N_47204,N_46828,N_46881);
nor U47205 (N_47205,N_46615,N_46698);
or U47206 (N_47206,N_46547,N_46788);
nor U47207 (N_47207,N_46542,N_46634);
nand U47208 (N_47208,N_46629,N_46989);
xor U47209 (N_47209,N_46639,N_46675);
nor U47210 (N_47210,N_46974,N_46908);
nor U47211 (N_47211,N_46590,N_46898);
and U47212 (N_47212,N_46508,N_46774);
and U47213 (N_47213,N_46531,N_46830);
nor U47214 (N_47214,N_46544,N_46894);
nand U47215 (N_47215,N_46665,N_46891);
nor U47216 (N_47216,N_46529,N_46555);
or U47217 (N_47217,N_46985,N_46984);
nand U47218 (N_47218,N_46648,N_46769);
nand U47219 (N_47219,N_46525,N_46651);
xnor U47220 (N_47220,N_46685,N_46936);
nor U47221 (N_47221,N_46921,N_46916);
nand U47222 (N_47222,N_46524,N_46944);
or U47223 (N_47223,N_46501,N_46800);
and U47224 (N_47224,N_46928,N_46948);
nand U47225 (N_47225,N_46837,N_46523);
nand U47226 (N_47226,N_46917,N_46528);
nand U47227 (N_47227,N_46859,N_46855);
or U47228 (N_47228,N_46717,N_46582);
xnor U47229 (N_47229,N_46869,N_46515);
nand U47230 (N_47230,N_46619,N_46700);
nand U47231 (N_47231,N_46962,N_46983);
nor U47232 (N_47232,N_46552,N_46842);
nand U47233 (N_47233,N_46668,N_46815);
nand U47234 (N_47234,N_46821,N_46784);
and U47235 (N_47235,N_46551,N_46849);
xor U47236 (N_47236,N_46625,N_46955);
and U47237 (N_47237,N_46906,N_46794);
or U47238 (N_47238,N_46777,N_46611);
nor U47239 (N_47239,N_46607,N_46746);
nand U47240 (N_47240,N_46930,N_46519);
and U47241 (N_47241,N_46538,N_46712);
or U47242 (N_47242,N_46872,N_46899);
xor U47243 (N_47243,N_46549,N_46793);
nor U47244 (N_47244,N_46867,N_46950);
nand U47245 (N_47245,N_46533,N_46873);
nor U47246 (N_47246,N_46797,N_46964);
or U47247 (N_47247,N_46838,N_46641);
nor U47248 (N_47248,N_46723,N_46708);
nor U47249 (N_47249,N_46901,N_46795);
and U47250 (N_47250,N_46998,N_46649);
nand U47251 (N_47251,N_46819,N_46965);
nor U47252 (N_47252,N_46941,N_46907);
or U47253 (N_47253,N_46780,N_46659);
xor U47254 (N_47254,N_46998,N_46848);
xor U47255 (N_47255,N_46807,N_46572);
or U47256 (N_47256,N_46658,N_46717);
and U47257 (N_47257,N_46631,N_46524);
nor U47258 (N_47258,N_46542,N_46582);
or U47259 (N_47259,N_46649,N_46534);
or U47260 (N_47260,N_46736,N_46966);
or U47261 (N_47261,N_46847,N_46512);
and U47262 (N_47262,N_46851,N_46904);
nor U47263 (N_47263,N_46879,N_46910);
and U47264 (N_47264,N_46995,N_46538);
xor U47265 (N_47265,N_46903,N_46532);
and U47266 (N_47266,N_46585,N_46594);
nand U47267 (N_47267,N_46668,N_46796);
nor U47268 (N_47268,N_46913,N_46962);
or U47269 (N_47269,N_46613,N_46746);
nor U47270 (N_47270,N_46872,N_46648);
nor U47271 (N_47271,N_46574,N_46673);
nor U47272 (N_47272,N_46652,N_46522);
xor U47273 (N_47273,N_46994,N_46894);
and U47274 (N_47274,N_46940,N_46542);
or U47275 (N_47275,N_46606,N_46991);
or U47276 (N_47276,N_46734,N_46597);
nand U47277 (N_47277,N_46994,N_46505);
nand U47278 (N_47278,N_46500,N_46629);
and U47279 (N_47279,N_46537,N_46661);
and U47280 (N_47280,N_46691,N_46745);
nor U47281 (N_47281,N_46581,N_46668);
nand U47282 (N_47282,N_46928,N_46733);
xnor U47283 (N_47283,N_46835,N_46960);
or U47284 (N_47284,N_46718,N_46900);
nand U47285 (N_47285,N_46808,N_46663);
or U47286 (N_47286,N_46894,N_46825);
nor U47287 (N_47287,N_46745,N_46994);
nand U47288 (N_47288,N_46564,N_46770);
or U47289 (N_47289,N_46908,N_46880);
or U47290 (N_47290,N_46773,N_46802);
nor U47291 (N_47291,N_46757,N_46815);
nor U47292 (N_47292,N_46985,N_46936);
nor U47293 (N_47293,N_46731,N_46704);
nand U47294 (N_47294,N_46600,N_46552);
nor U47295 (N_47295,N_46908,N_46796);
and U47296 (N_47296,N_46951,N_46776);
and U47297 (N_47297,N_46722,N_46713);
xor U47298 (N_47298,N_46555,N_46583);
nand U47299 (N_47299,N_46865,N_46588);
nor U47300 (N_47300,N_46740,N_46794);
nor U47301 (N_47301,N_46732,N_46641);
and U47302 (N_47302,N_46590,N_46885);
nand U47303 (N_47303,N_46947,N_46950);
and U47304 (N_47304,N_46682,N_46508);
nand U47305 (N_47305,N_46746,N_46911);
or U47306 (N_47306,N_46697,N_46530);
nand U47307 (N_47307,N_46644,N_46639);
xnor U47308 (N_47308,N_46959,N_46744);
or U47309 (N_47309,N_46933,N_46629);
xor U47310 (N_47310,N_46515,N_46680);
or U47311 (N_47311,N_46664,N_46770);
and U47312 (N_47312,N_46926,N_46741);
nand U47313 (N_47313,N_46669,N_46713);
and U47314 (N_47314,N_46751,N_46712);
xnor U47315 (N_47315,N_46562,N_46713);
nand U47316 (N_47316,N_46768,N_46857);
nor U47317 (N_47317,N_46917,N_46764);
nand U47318 (N_47318,N_46666,N_46687);
nor U47319 (N_47319,N_46749,N_46653);
and U47320 (N_47320,N_46693,N_46702);
and U47321 (N_47321,N_46983,N_46985);
and U47322 (N_47322,N_46889,N_46933);
nor U47323 (N_47323,N_46842,N_46505);
or U47324 (N_47324,N_46943,N_46787);
and U47325 (N_47325,N_46515,N_46806);
nor U47326 (N_47326,N_46947,N_46995);
and U47327 (N_47327,N_46833,N_46980);
nand U47328 (N_47328,N_46582,N_46594);
nand U47329 (N_47329,N_46922,N_46552);
nor U47330 (N_47330,N_46913,N_46676);
and U47331 (N_47331,N_46963,N_46665);
nand U47332 (N_47332,N_46557,N_46616);
and U47333 (N_47333,N_46725,N_46510);
or U47334 (N_47334,N_46749,N_46889);
and U47335 (N_47335,N_46864,N_46501);
nand U47336 (N_47336,N_46989,N_46657);
nor U47337 (N_47337,N_46894,N_46569);
or U47338 (N_47338,N_46542,N_46886);
xnor U47339 (N_47339,N_46730,N_46611);
nor U47340 (N_47340,N_46732,N_46688);
and U47341 (N_47341,N_46669,N_46682);
or U47342 (N_47342,N_46906,N_46560);
or U47343 (N_47343,N_46725,N_46525);
and U47344 (N_47344,N_46818,N_46917);
nor U47345 (N_47345,N_46749,N_46730);
nand U47346 (N_47346,N_46543,N_46795);
and U47347 (N_47347,N_46676,N_46800);
and U47348 (N_47348,N_46556,N_46969);
and U47349 (N_47349,N_46524,N_46832);
nor U47350 (N_47350,N_46645,N_46640);
xor U47351 (N_47351,N_46595,N_46855);
nand U47352 (N_47352,N_46783,N_46662);
nor U47353 (N_47353,N_46525,N_46569);
and U47354 (N_47354,N_46876,N_46681);
and U47355 (N_47355,N_46590,N_46839);
nor U47356 (N_47356,N_46658,N_46854);
nor U47357 (N_47357,N_46623,N_46961);
nor U47358 (N_47358,N_46547,N_46857);
nor U47359 (N_47359,N_46650,N_46770);
or U47360 (N_47360,N_46861,N_46886);
or U47361 (N_47361,N_46591,N_46957);
nand U47362 (N_47362,N_46719,N_46791);
xnor U47363 (N_47363,N_46888,N_46660);
nand U47364 (N_47364,N_46647,N_46986);
nand U47365 (N_47365,N_46872,N_46584);
xnor U47366 (N_47366,N_46603,N_46977);
and U47367 (N_47367,N_46710,N_46839);
xor U47368 (N_47368,N_46517,N_46787);
xnor U47369 (N_47369,N_46945,N_46563);
and U47370 (N_47370,N_46713,N_46847);
or U47371 (N_47371,N_46762,N_46883);
nand U47372 (N_47372,N_46666,N_46796);
xor U47373 (N_47373,N_46718,N_46848);
nor U47374 (N_47374,N_46586,N_46652);
or U47375 (N_47375,N_46550,N_46791);
xor U47376 (N_47376,N_46712,N_46886);
nor U47377 (N_47377,N_46624,N_46540);
nand U47378 (N_47378,N_46772,N_46791);
nand U47379 (N_47379,N_46613,N_46890);
or U47380 (N_47380,N_46990,N_46764);
and U47381 (N_47381,N_46533,N_46572);
nor U47382 (N_47382,N_46539,N_46808);
xor U47383 (N_47383,N_46924,N_46645);
or U47384 (N_47384,N_46519,N_46914);
xnor U47385 (N_47385,N_46842,N_46652);
and U47386 (N_47386,N_46855,N_46513);
nor U47387 (N_47387,N_46670,N_46653);
nor U47388 (N_47388,N_46681,N_46607);
nor U47389 (N_47389,N_46884,N_46989);
and U47390 (N_47390,N_46723,N_46747);
nor U47391 (N_47391,N_46758,N_46744);
xor U47392 (N_47392,N_46990,N_46892);
nand U47393 (N_47393,N_46667,N_46820);
and U47394 (N_47394,N_46884,N_46789);
nor U47395 (N_47395,N_46724,N_46654);
nand U47396 (N_47396,N_46628,N_46730);
xnor U47397 (N_47397,N_46608,N_46971);
nand U47398 (N_47398,N_46935,N_46559);
xor U47399 (N_47399,N_46504,N_46781);
xor U47400 (N_47400,N_46960,N_46737);
xor U47401 (N_47401,N_46710,N_46861);
or U47402 (N_47402,N_46819,N_46803);
nor U47403 (N_47403,N_46520,N_46663);
nand U47404 (N_47404,N_46678,N_46925);
nand U47405 (N_47405,N_46997,N_46534);
nor U47406 (N_47406,N_46925,N_46785);
nand U47407 (N_47407,N_46831,N_46801);
xor U47408 (N_47408,N_46787,N_46678);
nor U47409 (N_47409,N_46847,N_46880);
or U47410 (N_47410,N_46734,N_46555);
xnor U47411 (N_47411,N_46602,N_46811);
xor U47412 (N_47412,N_46976,N_46683);
and U47413 (N_47413,N_46700,N_46739);
nand U47414 (N_47414,N_46583,N_46637);
or U47415 (N_47415,N_46940,N_46883);
xor U47416 (N_47416,N_46735,N_46831);
and U47417 (N_47417,N_46764,N_46895);
and U47418 (N_47418,N_46945,N_46846);
nand U47419 (N_47419,N_46801,N_46692);
nor U47420 (N_47420,N_46893,N_46517);
nor U47421 (N_47421,N_46823,N_46681);
and U47422 (N_47422,N_46546,N_46883);
nor U47423 (N_47423,N_46580,N_46804);
nand U47424 (N_47424,N_46524,N_46688);
xnor U47425 (N_47425,N_46947,N_46801);
and U47426 (N_47426,N_46652,N_46813);
xor U47427 (N_47427,N_46719,N_46692);
nor U47428 (N_47428,N_46932,N_46954);
xor U47429 (N_47429,N_46895,N_46696);
or U47430 (N_47430,N_46794,N_46642);
or U47431 (N_47431,N_46588,N_46876);
nor U47432 (N_47432,N_46962,N_46569);
nand U47433 (N_47433,N_46669,N_46888);
xor U47434 (N_47434,N_46772,N_46501);
nand U47435 (N_47435,N_46960,N_46813);
or U47436 (N_47436,N_46875,N_46780);
nor U47437 (N_47437,N_46676,N_46825);
xnor U47438 (N_47438,N_46574,N_46949);
or U47439 (N_47439,N_46675,N_46764);
nor U47440 (N_47440,N_46733,N_46789);
or U47441 (N_47441,N_46810,N_46814);
and U47442 (N_47442,N_46827,N_46665);
xor U47443 (N_47443,N_46826,N_46995);
or U47444 (N_47444,N_46704,N_46723);
nor U47445 (N_47445,N_46665,N_46982);
xnor U47446 (N_47446,N_46785,N_46833);
nor U47447 (N_47447,N_46694,N_46641);
nor U47448 (N_47448,N_46720,N_46508);
nor U47449 (N_47449,N_46744,N_46707);
xor U47450 (N_47450,N_46523,N_46680);
nor U47451 (N_47451,N_46938,N_46688);
nand U47452 (N_47452,N_46826,N_46501);
xor U47453 (N_47453,N_46565,N_46803);
nand U47454 (N_47454,N_46732,N_46763);
xor U47455 (N_47455,N_46785,N_46511);
and U47456 (N_47456,N_46793,N_46923);
nor U47457 (N_47457,N_46629,N_46795);
nor U47458 (N_47458,N_46916,N_46603);
or U47459 (N_47459,N_46917,N_46826);
xnor U47460 (N_47460,N_46789,N_46581);
xor U47461 (N_47461,N_46727,N_46636);
or U47462 (N_47462,N_46714,N_46967);
nor U47463 (N_47463,N_46786,N_46701);
xnor U47464 (N_47464,N_46844,N_46945);
or U47465 (N_47465,N_46844,N_46912);
and U47466 (N_47466,N_46859,N_46543);
xnor U47467 (N_47467,N_46631,N_46957);
nor U47468 (N_47468,N_46545,N_46537);
nand U47469 (N_47469,N_46599,N_46575);
nand U47470 (N_47470,N_46619,N_46923);
xor U47471 (N_47471,N_46901,N_46632);
nor U47472 (N_47472,N_46573,N_46562);
and U47473 (N_47473,N_46958,N_46915);
or U47474 (N_47474,N_46643,N_46599);
and U47475 (N_47475,N_46660,N_46587);
nand U47476 (N_47476,N_46881,N_46599);
nor U47477 (N_47477,N_46556,N_46927);
and U47478 (N_47478,N_46515,N_46786);
nand U47479 (N_47479,N_46732,N_46757);
or U47480 (N_47480,N_46751,N_46681);
nor U47481 (N_47481,N_46623,N_46957);
nor U47482 (N_47482,N_46543,N_46619);
xor U47483 (N_47483,N_46945,N_46758);
nand U47484 (N_47484,N_46968,N_46961);
nor U47485 (N_47485,N_46608,N_46646);
nor U47486 (N_47486,N_46702,N_46889);
xor U47487 (N_47487,N_46740,N_46839);
or U47488 (N_47488,N_46631,N_46914);
and U47489 (N_47489,N_46509,N_46637);
nor U47490 (N_47490,N_46534,N_46547);
xnor U47491 (N_47491,N_46770,N_46786);
nand U47492 (N_47492,N_46726,N_46855);
or U47493 (N_47493,N_46506,N_46502);
xnor U47494 (N_47494,N_46984,N_46720);
xor U47495 (N_47495,N_46609,N_46805);
xnor U47496 (N_47496,N_46664,N_46960);
nand U47497 (N_47497,N_46597,N_46978);
and U47498 (N_47498,N_46986,N_46748);
nand U47499 (N_47499,N_46921,N_46703);
xnor U47500 (N_47500,N_47084,N_47264);
nand U47501 (N_47501,N_47087,N_47338);
nor U47502 (N_47502,N_47353,N_47400);
and U47503 (N_47503,N_47437,N_47430);
xor U47504 (N_47504,N_47054,N_47395);
xor U47505 (N_47505,N_47002,N_47132);
and U47506 (N_47506,N_47361,N_47076);
nand U47507 (N_47507,N_47456,N_47357);
and U47508 (N_47508,N_47309,N_47131);
and U47509 (N_47509,N_47021,N_47426);
and U47510 (N_47510,N_47033,N_47249);
nor U47511 (N_47511,N_47252,N_47205);
nand U47512 (N_47512,N_47261,N_47200);
nand U47513 (N_47513,N_47049,N_47274);
and U47514 (N_47514,N_47052,N_47152);
xnor U47515 (N_47515,N_47148,N_47053);
and U47516 (N_47516,N_47417,N_47399);
xnor U47517 (N_47517,N_47432,N_47320);
nor U47518 (N_47518,N_47050,N_47292);
nand U47519 (N_47519,N_47459,N_47276);
or U47520 (N_47520,N_47317,N_47204);
nand U47521 (N_47521,N_47032,N_47476);
nand U47522 (N_47522,N_47368,N_47420);
nor U47523 (N_47523,N_47123,N_47161);
nand U47524 (N_47524,N_47043,N_47405);
nor U47525 (N_47525,N_47070,N_47210);
or U47526 (N_47526,N_47051,N_47477);
or U47527 (N_47527,N_47362,N_47063);
nand U47528 (N_47528,N_47281,N_47128);
or U47529 (N_47529,N_47019,N_47270);
or U47530 (N_47530,N_47190,N_47453);
or U47531 (N_47531,N_47248,N_47209);
and U47532 (N_47532,N_47315,N_47055);
and U47533 (N_47533,N_47073,N_47351);
or U47534 (N_47534,N_47046,N_47316);
nor U47535 (N_47535,N_47157,N_47017);
or U47536 (N_47536,N_47085,N_47191);
nor U47537 (N_47537,N_47438,N_47402);
or U47538 (N_47538,N_47179,N_47170);
xnor U47539 (N_47539,N_47192,N_47067);
xnor U47540 (N_47540,N_47360,N_47334);
xnor U47541 (N_47541,N_47140,N_47375);
xor U47542 (N_47542,N_47306,N_47401);
and U47543 (N_47543,N_47197,N_47275);
or U47544 (N_47544,N_47410,N_47378);
and U47545 (N_47545,N_47178,N_47162);
and U47546 (N_47546,N_47236,N_47010);
xor U47547 (N_47547,N_47431,N_47117);
and U47548 (N_47548,N_47451,N_47327);
and U47549 (N_47549,N_47221,N_47044);
xnor U47550 (N_47550,N_47096,N_47314);
xnor U47551 (N_47551,N_47189,N_47089);
xor U47552 (N_47552,N_47484,N_47255);
and U47553 (N_47553,N_47020,N_47481);
and U47554 (N_47554,N_47290,N_47271);
nor U47555 (N_47555,N_47372,N_47244);
nor U47556 (N_47556,N_47294,N_47233);
xnor U47557 (N_47557,N_47134,N_47377);
or U47558 (N_47558,N_47074,N_47155);
xor U47559 (N_47559,N_47078,N_47038);
and U47560 (N_47560,N_47196,N_47268);
nor U47561 (N_47561,N_47245,N_47100);
or U47562 (N_47562,N_47416,N_47068);
or U47563 (N_47563,N_47120,N_47494);
xnor U47564 (N_47564,N_47339,N_47103);
nor U47565 (N_47565,N_47231,N_47411);
xor U47566 (N_47566,N_47203,N_47165);
or U47567 (N_47567,N_47222,N_47267);
and U47568 (N_47568,N_47141,N_47390);
or U47569 (N_47569,N_47007,N_47090);
xor U47570 (N_47570,N_47319,N_47279);
xor U47571 (N_47571,N_47452,N_47408);
or U47572 (N_47572,N_47313,N_47036);
nand U47573 (N_47573,N_47440,N_47124);
xor U47574 (N_47574,N_47455,N_47163);
nor U47575 (N_47575,N_47235,N_47119);
nor U47576 (N_47576,N_47150,N_47482);
nand U47577 (N_47577,N_47355,N_47146);
xnor U47578 (N_47578,N_47018,N_47356);
and U47579 (N_47579,N_47116,N_47006);
nor U47580 (N_47580,N_47158,N_47487);
or U47581 (N_47581,N_47139,N_47135);
xnor U47582 (N_47582,N_47181,N_47121);
and U47583 (N_47583,N_47444,N_47262);
and U47584 (N_47584,N_47365,N_47393);
or U47585 (N_47585,N_47156,N_47412);
or U47586 (N_47586,N_47228,N_47154);
nor U47587 (N_47587,N_47391,N_47492);
nor U47588 (N_47588,N_47238,N_47212);
and U47589 (N_47589,N_47387,N_47213);
and U47590 (N_47590,N_47498,N_47218);
nor U47591 (N_47591,N_47024,N_47422);
and U47592 (N_47592,N_47079,N_47081);
nand U47593 (N_47593,N_47407,N_47436);
and U47594 (N_47594,N_47464,N_47388);
and U47595 (N_47595,N_47095,N_47297);
or U47596 (N_47596,N_47376,N_47035);
nand U47597 (N_47597,N_47369,N_47042);
xnor U47598 (N_47598,N_47225,N_47045);
xor U47599 (N_47599,N_47047,N_47478);
xnor U47600 (N_47600,N_47461,N_47465);
xor U47601 (N_47601,N_47475,N_47112);
nand U47602 (N_47602,N_47256,N_47187);
xor U47603 (N_47603,N_47347,N_47130);
nor U47604 (N_47604,N_47489,N_47058);
xnor U47605 (N_47605,N_47182,N_47237);
xnor U47606 (N_47606,N_47424,N_47349);
or U47607 (N_47607,N_47291,N_47384);
nand U47608 (N_47608,N_47083,N_47341);
and U47609 (N_47609,N_47031,N_47293);
nor U47610 (N_47610,N_47447,N_47115);
and U47611 (N_47611,N_47202,N_47258);
and U47612 (N_47612,N_47460,N_47499);
and U47613 (N_47613,N_47318,N_47380);
xor U47614 (N_47614,N_47092,N_47323);
nand U47615 (N_47615,N_47015,N_47295);
or U47616 (N_47616,N_47488,N_47427);
or U47617 (N_47617,N_47324,N_47423);
or U47618 (N_47618,N_47345,N_47304);
and U47619 (N_47619,N_47396,N_47253);
xnor U47620 (N_47620,N_47136,N_47030);
or U47621 (N_47621,N_47126,N_47449);
xnor U47622 (N_47622,N_47298,N_47001);
nor U47623 (N_47623,N_47137,N_47188);
nor U47624 (N_47624,N_47025,N_47207);
xor U47625 (N_47625,N_47113,N_47075);
or U47626 (N_47626,N_47344,N_47160);
nand U47627 (N_47627,N_47057,N_47493);
nand U47628 (N_47628,N_47004,N_47346);
nand U47629 (N_47629,N_47138,N_47288);
nor U47630 (N_47630,N_47348,N_47448);
nor U47631 (N_47631,N_47485,N_47370);
and U47632 (N_47632,N_47382,N_47082);
or U47633 (N_47633,N_47056,N_47127);
nor U47634 (N_47634,N_47091,N_47326);
nand U47635 (N_47635,N_47180,N_47220);
nand U47636 (N_47636,N_47446,N_47143);
nor U47637 (N_47637,N_47234,N_47230);
xnor U47638 (N_47638,N_47098,N_47342);
xnor U47639 (N_47639,N_47468,N_47419);
nand U47640 (N_47640,N_47337,N_47022);
nand U47641 (N_47641,N_47110,N_47273);
xor U47642 (N_47642,N_47284,N_47201);
or U47643 (N_47643,N_47097,N_47443);
nand U47644 (N_47644,N_47166,N_47389);
or U47645 (N_47645,N_47217,N_47149);
and U47646 (N_47646,N_47172,N_47107);
nor U47647 (N_47647,N_47198,N_47027);
or U47648 (N_47648,N_47287,N_47462);
nand U47649 (N_47649,N_47232,N_47173);
xor U47650 (N_47650,N_47397,N_47094);
and U47651 (N_47651,N_47403,N_47214);
or U47652 (N_47652,N_47229,N_47026);
xor U47653 (N_47653,N_47077,N_47226);
nand U47654 (N_47654,N_47216,N_47206);
or U47655 (N_47655,N_47479,N_47414);
or U47656 (N_47656,N_47394,N_47219);
or U47657 (N_47657,N_47223,N_47330);
nor U47658 (N_47658,N_47069,N_47061);
or U47659 (N_47659,N_47308,N_47491);
and U47660 (N_47660,N_47406,N_47260);
or U47661 (N_47661,N_47254,N_47003);
xnor U47662 (N_47662,N_47208,N_47147);
or U47663 (N_47663,N_47373,N_47159);
xnor U47664 (N_47664,N_47144,N_47343);
and U47665 (N_47665,N_47301,N_47215);
and U47666 (N_47666,N_47005,N_47183);
xnor U47667 (N_47667,N_47102,N_47305);
or U47668 (N_47668,N_47106,N_47280);
or U47669 (N_47669,N_47329,N_47433);
xor U47670 (N_47670,N_47474,N_47088);
nand U47671 (N_47671,N_47366,N_47310);
nand U47672 (N_47672,N_47122,N_47413);
or U47673 (N_47673,N_47383,N_47016);
xor U47674 (N_47674,N_47059,N_47064);
and U47675 (N_47675,N_47333,N_47358);
nand U47676 (N_47676,N_47086,N_47014);
and U47677 (N_47677,N_47250,N_47177);
nand U47678 (N_47678,N_47466,N_47335);
and U47679 (N_47679,N_47142,N_47296);
nand U47680 (N_47680,N_47429,N_47379);
xnor U47681 (N_47681,N_47496,N_47392);
nand U47682 (N_47682,N_47224,N_47193);
nor U47683 (N_47683,N_47381,N_47167);
nor U47684 (N_47684,N_47286,N_47269);
xnor U47685 (N_47685,N_47041,N_47425);
nor U47686 (N_47686,N_47463,N_47171);
or U47687 (N_47687,N_47263,N_47108);
xor U47688 (N_47688,N_47458,N_47325);
nor U47689 (N_47689,N_47299,N_47359);
or U47690 (N_47690,N_47328,N_47145);
nand U47691 (N_47691,N_47243,N_47114);
and U47692 (N_47692,N_47247,N_47374);
xor U47693 (N_47693,N_47282,N_47289);
and U47694 (N_47694,N_47457,N_47454);
or U47695 (N_47695,N_47104,N_47009);
and U47696 (N_47696,N_47239,N_47164);
xor U47697 (N_47697,N_47013,N_47311);
nor U47698 (N_47698,N_47278,N_47418);
xor U47699 (N_47699,N_47008,N_47495);
nor U47700 (N_47700,N_47011,N_47272);
and U47701 (N_47701,N_47241,N_47490);
and U47702 (N_47702,N_47386,N_47012);
or U47703 (N_47703,N_47153,N_47322);
xnor U47704 (N_47704,N_47111,N_47065);
nor U47705 (N_47705,N_47099,N_47450);
nor U47706 (N_47706,N_47340,N_47168);
and U47707 (N_47707,N_47133,N_47175);
or U47708 (N_47708,N_47093,N_47277);
and U47709 (N_47709,N_47415,N_47385);
xor U47710 (N_47710,N_47404,N_47303);
nand U47711 (N_47711,N_47442,N_47435);
nor U47712 (N_47712,N_47251,N_47473);
or U47713 (N_47713,N_47028,N_47101);
and U47714 (N_47714,N_47039,N_47125);
and U47715 (N_47715,N_47363,N_47354);
or U47716 (N_47716,N_47023,N_47000);
nand U47717 (N_47717,N_47497,N_47048);
and U47718 (N_47718,N_47037,N_47060);
and U47719 (N_47719,N_47409,N_47195);
and U47720 (N_47720,N_47472,N_47129);
xor U47721 (N_47721,N_47118,N_47441);
xor U47722 (N_47722,N_47350,N_47176);
or U47723 (N_47723,N_47194,N_47398);
nor U47724 (N_47724,N_47109,N_47227);
nand U47725 (N_47725,N_47421,N_47467);
or U47726 (N_47726,N_47312,N_47300);
and U47727 (N_47727,N_47364,N_47321);
nand U47728 (N_47728,N_47471,N_47439);
nor U47729 (N_47729,N_47470,N_47445);
nand U47730 (N_47730,N_47034,N_47105);
nand U47731 (N_47731,N_47480,N_47040);
or U47732 (N_47732,N_47266,N_47080);
and U47733 (N_47733,N_47332,N_47211);
and U47734 (N_47734,N_47029,N_47071);
xor U47735 (N_47735,N_47483,N_47186);
and U47736 (N_47736,N_47062,N_47199);
and U47737 (N_47737,N_47242,N_47352);
and U47738 (N_47738,N_47486,N_47174);
nand U47739 (N_47739,N_47367,N_47257);
xnor U47740 (N_47740,N_47285,N_47434);
and U47741 (N_47741,N_47259,N_47428);
or U47742 (N_47742,N_47184,N_47469);
xor U47743 (N_47743,N_47151,N_47331);
nand U47744 (N_47744,N_47185,N_47283);
or U47745 (N_47745,N_47265,N_47302);
nor U47746 (N_47746,N_47066,N_47336);
or U47747 (N_47747,N_47169,N_47240);
nand U47748 (N_47748,N_47371,N_47072);
nor U47749 (N_47749,N_47307,N_47246);
nor U47750 (N_47750,N_47438,N_47197);
or U47751 (N_47751,N_47150,N_47134);
nor U47752 (N_47752,N_47342,N_47211);
nor U47753 (N_47753,N_47247,N_47262);
and U47754 (N_47754,N_47093,N_47223);
nor U47755 (N_47755,N_47288,N_47112);
nand U47756 (N_47756,N_47438,N_47414);
xor U47757 (N_47757,N_47349,N_47047);
nor U47758 (N_47758,N_47453,N_47394);
nand U47759 (N_47759,N_47339,N_47155);
and U47760 (N_47760,N_47192,N_47133);
and U47761 (N_47761,N_47381,N_47430);
and U47762 (N_47762,N_47015,N_47284);
and U47763 (N_47763,N_47075,N_47416);
nand U47764 (N_47764,N_47330,N_47025);
nand U47765 (N_47765,N_47284,N_47489);
xor U47766 (N_47766,N_47152,N_47104);
nor U47767 (N_47767,N_47047,N_47393);
or U47768 (N_47768,N_47453,N_47166);
or U47769 (N_47769,N_47349,N_47432);
or U47770 (N_47770,N_47097,N_47227);
nand U47771 (N_47771,N_47385,N_47246);
or U47772 (N_47772,N_47073,N_47269);
nand U47773 (N_47773,N_47401,N_47167);
nor U47774 (N_47774,N_47151,N_47239);
nand U47775 (N_47775,N_47384,N_47104);
and U47776 (N_47776,N_47307,N_47139);
or U47777 (N_47777,N_47313,N_47090);
xnor U47778 (N_47778,N_47263,N_47450);
xor U47779 (N_47779,N_47389,N_47261);
or U47780 (N_47780,N_47410,N_47079);
nand U47781 (N_47781,N_47447,N_47346);
nand U47782 (N_47782,N_47076,N_47153);
or U47783 (N_47783,N_47214,N_47222);
nor U47784 (N_47784,N_47040,N_47032);
nand U47785 (N_47785,N_47257,N_47337);
nand U47786 (N_47786,N_47369,N_47054);
nor U47787 (N_47787,N_47061,N_47403);
or U47788 (N_47788,N_47068,N_47299);
xor U47789 (N_47789,N_47137,N_47254);
nand U47790 (N_47790,N_47236,N_47348);
and U47791 (N_47791,N_47061,N_47395);
nor U47792 (N_47792,N_47338,N_47275);
and U47793 (N_47793,N_47212,N_47464);
and U47794 (N_47794,N_47350,N_47067);
and U47795 (N_47795,N_47489,N_47064);
nand U47796 (N_47796,N_47252,N_47286);
or U47797 (N_47797,N_47104,N_47151);
xor U47798 (N_47798,N_47017,N_47440);
and U47799 (N_47799,N_47367,N_47047);
nand U47800 (N_47800,N_47136,N_47492);
nand U47801 (N_47801,N_47055,N_47343);
or U47802 (N_47802,N_47451,N_47137);
nor U47803 (N_47803,N_47347,N_47466);
xor U47804 (N_47804,N_47264,N_47158);
and U47805 (N_47805,N_47271,N_47419);
nand U47806 (N_47806,N_47307,N_47313);
xor U47807 (N_47807,N_47342,N_47262);
xor U47808 (N_47808,N_47379,N_47109);
and U47809 (N_47809,N_47094,N_47136);
and U47810 (N_47810,N_47326,N_47380);
nor U47811 (N_47811,N_47496,N_47441);
and U47812 (N_47812,N_47077,N_47378);
or U47813 (N_47813,N_47305,N_47110);
or U47814 (N_47814,N_47196,N_47445);
and U47815 (N_47815,N_47405,N_47040);
nor U47816 (N_47816,N_47194,N_47392);
nand U47817 (N_47817,N_47380,N_47196);
or U47818 (N_47818,N_47109,N_47104);
nand U47819 (N_47819,N_47084,N_47383);
xor U47820 (N_47820,N_47302,N_47321);
nand U47821 (N_47821,N_47143,N_47320);
and U47822 (N_47822,N_47251,N_47247);
or U47823 (N_47823,N_47389,N_47422);
nor U47824 (N_47824,N_47326,N_47154);
xnor U47825 (N_47825,N_47075,N_47445);
nand U47826 (N_47826,N_47055,N_47107);
and U47827 (N_47827,N_47382,N_47014);
or U47828 (N_47828,N_47218,N_47065);
nor U47829 (N_47829,N_47015,N_47185);
nand U47830 (N_47830,N_47431,N_47342);
nand U47831 (N_47831,N_47331,N_47341);
nand U47832 (N_47832,N_47218,N_47484);
nand U47833 (N_47833,N_47248,N_47188);
or U47834 (N_47834,N_47366,N_47119);
and U47835 (N_47835,N_47157,N_47446);
and U47836 (N_47836,N_47123,N_47326);
and U47837 (N_47837,N_47074,N_47445);
nor U47838 (N_47838,N_47331,N_47055);
and U47839 (N_47839,N_47106,N_47039);
nand U47840 (N_47840,N_47304,N_47450);
or U47841 (N_47841,N_47280,N_47093);
or U47842 (N_47842,N_47328,N_47132);
or U47843 (N_47843,N_47002,N_47192);
and U47844 (N_47844,N_47049,N_47252);
xnor U47845 (N_47845,N_47072,N_47263);
nand U47846 (N_47846,N_47159,N_47279);
or U47847 (N_47847,N_47011,N_47113);
and U47848 (N_47848,N_47400,N_47371);
nand U47849 (N_47849,N_47443,N_47369);
and U47850 (N_47850,N_47232,N_47426);
xor U47851 (N_47851,N_47317,N_47458);
xor U47852 (N_47852,N_47160,N_47353);
nand U47853 (N_47853,N_47241,N_47354);
or U47854 (N_47854,N_47035,N_47275);
nor U47855 (N_47855,N_47367,N_47448);
and U47856 (N_47856,N_47387,N_47293);
xor U47857 (N_47857,N_47031,N_47485);
nor U47858 (N_47858,N_47461,N_47326);
or U47859 (N_47859,N_47029,N_47477);
nor U47860 (N_47860,N_47418,N_47378);
nor U47861 (N_47861,N_47449,N_47083);
or U47862 (N_47862,N_47208,N_47217);
and U47863 (N_47863,N_47158,N_47068);
nor U47864 (N_47864,N_47438,N_47257);
and U47865 (N_47865,N_47146,N_47482);
or U47866 (N_47866,N_47413,N_47218);
or U47867 (N_47867,N_47307,N_47430);
and U47868 (N_47868,N_47195,N_47075);
nor U47869 (N_47869,N_47428,N_47110);
xnor U47870 (N_47870,N_47322,N_47356);
nand U47871 (N_47871,N_47017,N_47367);
and U47872 (N_47872,N_47459,N_47416);
nor U47873 (N_47873,N_47029,N_47301);
and U47874 (N_47874,N_47183,N_47014);
and U47875 (N_47875,N_47010,N_47056);
xnor U47876 (N_47876,N_47401,N_47346);
or U47877 (N_47877,N_47493,N_47084);
xor U47878 (N_47878,N_47389,N_47031);
nand U47879 (N_47879,N_47184,N_47460);
xnor U47880 (N_47880,N_47107,N_47193);
nand U47881 (N_47881,N_47039,N_47100);
xor U47882 (N_47882,N_47351,N_47009);
nor U47883 (N_47883,N_47401,N_47422);
or U47884 (N_47884,N_47484,N_47284);
xnor U47885 (N_47885,N_47145,N_47401);
and U47886 (N_47886,N_47419,N_47377);
and U47887 (N_47887,N_47295,N_47173);
nor U47888 (N_47888,N_47030,N_47254);
nand U47889 (N_47889,N_47218,N_47497);
or U47890 (N_47890,N_47393,N_47211);
nand U47891 (N_47891,N_47053,N_47495);
or U47892 (N_47892,N_47297,N_47428);
nor U47893 (N_47893,N_47454,N_47118);
or U47894 (N_47894,N_47326,N_47297);
or U47895 (N_47895,N_47090,N_47198);
xnor U47896 (N_47896,N_47339,N_47109);
or U47897 (N_47897,N_47303,N_47209);
or U47898 (N_47898,N_47111,N_47291);
nand U47899 (N_47899,N_47339,N_47436);
nor U47900 (N_47900,N_47044,N_47060);
xor U47901 (N_47901,N_47140,N_47167);
nor U47902 (N_47902,N_47066,N_47496);
xor U47903 (N_47903,N_47008,N_47437);
xor U47904 (N_47904,N_47345,N_47369);
or U47905 (N_47905,N_47464,N_47184);
and U47906 (N_47906,N_47192,N_47387);
nor U47907 (N_47907,N_47289,N_47375);
nand U47908 (N_47908,N_47496,N_47168);
xor U47909 (N_47909,N_47233,N_47394);
nor U47910 (N_47910,N_47239,N_47478);
and U47911 (N_47911,N_47321,N_47332);
nor U47912 (N_47912,N_47183,N_47033);
nor U47913 (N_47913,N_47453,N_47255);
xor U47914 (N_47914,N_47134,N_47289);
nand U47915 (N_47915,N_47397,N_47493);
xnor U47916 (N_47916,N_47331,N_47272);
or U47917 (N_47917,N_47410,N_47284);
and U47918 (N_47918,N_47278,N_47300);
nand U47919 (N_47919,N_47450,N_47171);
or U47920 (N_47920,N_47113,N_47193);
xor U47921 (N_47921,N_47107,N_47472);
or U47922 (N_47922,N_47266,N_47346);
or U47923 (N_47923,N_47284,N_47072);
or U47924 (N_47924,N_47084,N_47249);
xnor U47925 (N_47925,N_47319,N_47202);
nor U47926 (N_47926,N_47495,N_47288);
and U47927 (N_47927,N_47366,N_47062);
or U47928 (N_47928,N_47203,N_47142);
and U47929 (N_47929,N_47305,N_47082);
and U47930 (N_47930,N_47302,N_47244);
nor U47931 (N_47931,N_47379,N_47445);
nand U47932 (N_47932,N_47498,N_47334);
nor U47933 (N_47933,N_47210,N_47336);
and U47934 (N_47934,N_47356,N_47162);
xor U47935 (N_47935,N_47196,N_47138);
xnor U47936 (N_47936,N_47098,N_47174);
nand U47937 (N_47937,N_47249,N_47369);
xnor U47938 (N_47938,N_47040,N_47155);
nand U47939 (N_47939,N_47267,N_47002);
nand U47940 (N_47940,N_47475,N_47169);
xnor U47941 (N_47941,N_47292,N_47470);
and U47942 (N_47942,N_47160,N_47299);
and U47943 (N_47943,N_47074,N_47381);
xnor U47944 (N_47944,N_47001,N_47145);
xnor U47945 (N_47945,N_47444,N_47175);
nor U47946 (N_47946,N_47145,N_47189);
nor U47947 (N_47947,N_47462,N_47050);
and U47948 (N_47948,N_47367,N_47224);
nand U47949 (N_47949,N_47485,N_47310);
or U47950 (N_47950,N_47443,N_47005);
nor U47951 (N_47951,N_47170,N_47107);
nand U47952 (N_47952,N_47475,N_47258);
nand U47953 (N_47953,N_47474,N_47353);
nor U47954 (N_47954,N_47482,N_47177);
nor U47955 (N_47955,N_47109,N_47319);
nor U47956 (N_47956,N_47362,N_47082);
and U47957 (N_47957,N_47197,N_47153);
nor U47958 (N_47958,N_47138,N_47427);
nand U47959 (N_47959,N_47418,N_47300);
nand U47960 (N_47960,N_47107,N_47098);
and U47961 (N_47961,N_47169,N_47345);
and U47962 (N_47962,N_47080,N_47061);
xnor U47963 (N_47963,N_47376,N_47049);
nand U47964 (N_47964,N_47261,N_47230);
and U47965 (N_47965,N_47112,N_47173);
nand U47966 (N_47966,N_47254,N_47193);
nand U47967 (N_47967,N_47467,N_47087);
and U47968 (N_47968,N_47455,N_47291);
and U47969 (N_47969,N_47400,N_47159);
and U47970 (N_47970,N_47048,N_47112);
nor U47971 (N_47971,N_47498,N_47182);
nand U47972 (N_47972,N_47396,N_47256);
nor U47973 (N_47973,N_47325,N_47102);
nand U47974 (N_47974,N_47218,N_47021);
xnor U47975 (N_47975,N_47185,N_47357);
or U47976 (N_47976,N_47163,N_47179);
and U47977 (N_47977,N_47103,N_47435);
nand U47978 (N_47978,N_47388,N_47335);
or U47979 (N_47979,N_47038,N_47356);
or U47980 (N_47980,N_47005,N_47459);
nor U47981 (N_47981,N_47419,N_47447);
or U47982 (N_47982,N_47020,N_47152);
nor U47983 (N_47983,N_47322,N_47167);
xnor U47984 (N_47984,N_47492,N_47152);
or U47985 (N_47985,N_47414,N_47218);
or U47986 (N_47986,N_47045,N_47397);
nand U47987 (N_47987,N_47326,N_47230);
or U47988 (N_47988,N_47094,N_47337);
and U47989 (N_47989,N_47052,N_47370);
and U47990 (N_47990,N_47401,N_47075);
nand U47991 (N_47991,N_47199,N_47090);
xnor U47992 (N_47992,N_47391,N_47168);
xnor U47993 (N_47993,N_47122,N_47141);
nor U47994 (N_47994,N_47082,N_47108);
or U47995 (N_47995,N_47104,N_47463);
and U47996 (N_47996,N_47367,N_47465);
or U47997 (N_47997,N_47372,N_47015);
or U47998 (N_47998,N_47471,N_47045);
and U47999 (N_47999,N_47032,N_47169);
nor U48000 (N_48000,N_47631,N_47837);
xor U48001 (N_48001,N_47684,N_47556);
and U48002 (N_48002,N_47740,N_47530);
nor U48003 (N_48003,N_47725,N_47735);
nand U48004 (N_48004,N_47944,N_47750);
or U48005 (N_48005,N_47905,N_47644);
nor U48006 (N_48006,N_47538,N_47649);
nand U48007 (N_48007,N_47659,N_47570);
and U48008 (N_48008,N_47799,N_47707);
or U48009 (N_48009,N_47935,N_47857);
or U48010 (N_48010,N_47965,N_47507);
xor U48011 (N_48011,N_47950,N_47625);
nor U48012 (N_48012,N_47545,N_47918);
nor U48013 (N_48013,N_47709,N_47984);
and U48014 (N_48014,N_47894,N_47689);
nor U48015 (N_48015,N_47879,N_47923);
nand U48016 (N_48016,N_47563,N_47974);
or U48017 (N_48017,N_47737,N_47827);
and U48018 (N_48018,N_47620,N_47742);
or U48019 (N_48019,N_47616,N_47517);
or U48020 (N_48020,N_47568,N_47623);
nor U48021 (N_48021,N_47895,N_47774);
or U48022 (N_48022,N_47912,N_47940);
nand U48023 (N_48023,N_47520,N_47738);
and U48024 (N_48024,N_47762,N_47825);
nand U48025 (N_48025,N_47772,N_47856);
nor U48026 (N_48026,N_47942,N_47964);
nor U48027 (N_48027,N_47686,N_47701);
or U48028 (N_48028,N_47578,N_47654);
xnor U48029 (N_48029,N_47501,N_47915);
and U48030 (N_48030,N_47830,N_47829);
and U48031 (N_48031,N_47613,N_47593);
xor U48032 (N_48032,N_47632,N_47758);
or U48033 (N_48033,N_47702,N_47589);
nand U48034 (N_48034,N_47533,N_47693);
or U48035 (N_48035,N_47720,N_47933);
nor U48036 (N_48036,N_47853,N_47989);
nand U48037 (N_48037,N_47892,N_47877);
and U48038 (N_48038,N_47549,N_47551);
and U48039 (N_48039,N_47711,N_47636);
nor U48040 (N_48040,N_47721,N_47931);
nor U48041 (N_48041,N_47559,N_47565);
and U48042 (N_48042,N_47662,N_47717);
or U48043 (N_48043,N_47751,N_47675);
nand U48044 (N_48044,N_47951,N_47767);
and U48045 (N_48045,N_47775,N_47987);
xor U48046 (N_48046,N_47528,N_47618);
nand U48047 (N_48047,N_47511,N_47722);
nor U48048 (N_48048,N_47922,N_47876);
nand U48049 (N_48049,N_47692,N_47843);
nand U48050 (N_48050,N_47847,N_47599);
and U48051 (N_48051,N_47865,N_47582);
nor U48052 (N_48052,N_47901,N_47907);
xor U48053 (N_48053,N_47956,N_47805);
and U48054 (N_48054,N_47777,N_47954);
and U48055 (N_48055,N_47808,N_47588);
xnor U48056 (N_48056,N_47803,N_47560);
nand U48057 (N_48057,N_47878,N_47855);
and U48058 (N_48058,N_47836,N_47985);
nand U48059 (N_48059,N_47612,N_47748);
nor U48060 (N_48060,N_47888,N_47873);
or U48061 (N_48061,N_47884,N_47890);
or U48062 (N_48062,N_47869,N_47605);
xnor U48063 (N_48063,N_47575,N_47976);
xor U48064 (N_48064,N_47997,N_47561);
xnor U48065 (N_48065,N_47866,N_47999);
nor U48066 (N_48066,N_47790,N_47713);
nor U48067 (N_48067,N_47630,N_47848);
nand U48068 (N_48068,N_47728,N_47506);
and U48069 (N_48069,N_47945,N_47546);
nor U48070 (N_48070,N_47595,N_47586);
nor U48071 (N_48071,N_47900,N_47990);
or U48072 (N_48072,N_47973,N_47862);
xor U48073 (N_48073,N_47801,N_47638);
xor U48074 (N_48074,N_47883,N_47844);
and U48075 (N_48075,N_47733,N_47606);
nor U48076 (N_48076,N_47591,N_47510);
nor U48077 (N_48077,N_47696,N_47641);
nor U48078 (N_48078,N_47508,N_47840);
nand U48079 (N_48079,N_47513,N_47726);
xnor U48080 (N_48080,N_47664,N_47668);
nand U48081 (N_48081,N_47723,N_47946);
xnor U48082 (N_48082,N_47859,N_47809);
xor U48083 (N_48083,N_47665,N_47779);
nand U48084 (N_48084,N_47712,N_47653);
nand U48085 (N_48085,N_47695,N_47972);
xor U48086 (N_48086,N_47786,N_47534);
nand U48087 (N_48087,N_47705,N_47953);
nor U48088 (N_48088,N_47962,N_47650);
nor U48089 (N_48089,N_47567,N_47754);
or U48090 (N_48090,N_47979,N_47542);
or U48091 (N_48091,N_47646,N_47681);
xor U48092 (N_48092,N_47724,N_47746);
xor U48093 (N_48093,N_47532,N_47634);
xor U48094 (N_48094,N_47562,N_47887);
or U48095 (N_48095,N_47991,N_47832);
and U48096 (N_48096,N_47503,N_47755);
xor U48097 (N_48097,N_47581,N_47903);
xnor U48098 (N_48098,N_47908,N_47967);
nand U48099 (N_48099,N_47604,N_47958);
xnor U48100 (N_48100,N_47594,N_47937);
and U48101 (N_48101,N_47739,N_47708);
or U48102 (N_48102,N_47614,N_47670);
xor U48103 (N_48103,N_47917,N_47525);
xnor U48104 (N_48104,N_47863,N_47926);
or U48105 (N_48105,N_47858,N_47988);
nor U48106 (N_48106,N_47592,N_47679);
nand U48107 (N_48107,N_47909,N_47934);
xor U48108 (N_48108,N_47698,N_47615);
or U48109 (N_48109,N_47536,N_47704);
or U48110 (N_48110,N_47544,N_47672);
xor U48111 (N_48111,N_47732,N_47687);
nor U48112 (N_48112,N_47813,N_47761);
xnor U48113 (N_48113,N_47524,N_47669);
and U48114 (N_48114,N_47998,N_47502);
and U48115 (N_48115,N_47763,N_47769);
xor U48116 (N_48116,N_47941,N_47854);
xor U48117 (N_48117,N_47910,N_47817);
and U48118 (N_48118,N_47948,N_47831);
nand U48119 (N_48119,N_47685,N_47655);
nand U48120 (N_48120,N_47509,N_47656);
nor U48121 (N_48121,N_47554,N_47785);
nand U48122 (N_48122,N_47804,N_47798);
xnor U48123 (N_48123,N_47872,N_47519);
xnor U48124 (N_48124,N_47572,N_47810);
nand U48125 (N_48125,N_47826,N_47752);
nor U48126 (N_48126,N_47573,N_47885);
and U48127 (N_48127,N_47791,N_47504);
xnor U48128 (N_48128,N_47743,N_47602);
nor U48129 (N_48129,N_47842,N_47821);
nand U48130 (N_48130,N_47811,N_47778);
xnor U48131 (N_48131,N_47930,N_47947);
and U48132 (N_48132,N_47577,N_47643);
or U48133 (N_48133,N_47626,N_47784);
or U48134 (N_48134,N_47677,N_47986);
nor U48135 (N_48135,N_47526,N_47658);
and U48136 (N_48136,N_47640,N_47579);
or U48137 (N_48137,N_47652,N_47610);
nand U48138 (N_48138,N_47523,N_47527);
nor U48139 (N_48139,N_47812,N_47794);
xnor U48140 (N_48140,N_47860,N_47793);
nand U48141 (N_48141,N_47943,N_47764);
nor U48142 (N_48142,N_47555,N_47768);
nor U48143 (N_48143,N_47874,N_47939);
xnor U48144 (N_48144,N_47906,N_47928);
and U48145 (N_48145,N_47982,N_47787);
and U48146 (N_48146,N_47564,N_47897);
nand U48147 (N_48147,N_47674,N_47637);
and U48148 (N_48148,N_47795,N_47929);
and U48149 (N_48149,N_47667,N_47603);
xor U48150 (N_48150,N_47896,N_47963);
and U48151 (N_48151,N_47970,N_47642);
nor U48152 (N_48152,N_47816,N_47920);
and U48153 (N_48153,N_47961,N_47714);
or U48154 (N_48154,N_47727,N_47518);
xor U48155 (N_48155,N_47835,N_47584);
nand U48156 (N_48156,N_47516,N_47512);
and U48157 (N_48157,N_47719,N_47938);
and U48158 (N_48158,N_47776,N_47601);
nand U48159 (N_48159,N_47797,N_47870);
or U48160 (N_48160,N_47959,N_47760);
and U48161 (N_48161,N_47557,N_47780);
or U48162 (N_48162,N_47992,N_47569);
or U48163 (N_48163,N_47932,N_47690);
nand U48164 (N_48164,N_47741,N_47770);
or U48165 (N_48165,N_47541,N_47807);
or U48166 (N_48166,N_47757,N_47834);
or U48167 (N_48167,N_47745,N_47846);
nand U48168 (N_48168,N_47773,N_47683);
nor U48169 (N_48169,N_47529,N_47782);
and U48170 (N_48170,N_47676,N_47949);
nor U48171 (N_48171,N_47971,N_47680);
nand U48172 (N_48172,N_47839,N_47585);
or U48173 (N_48173,N_47522,N_47688);
xor U48174 (N_48174,N_47747,N_47871);
xnor U48175 (N_48175,N_47633,N_47600);
or U48176 (N_48176,N_47734,N_47868);
xnor U48177 (N_48177,N_47815,N_47994);
xor U48178 (N_48178,N_47925,N_47823);
nor U48179 (N_48179,N_47596,N_47898);
xnor U48180 (N_48180,N_47715,N_47911);
nand U48181 (N_48181,N_47771,N_47766);
and U48182 (N_48182,N_47703,N_47818);
and U48183 (N_48183,N_47983,N_47966);
xnor U48184 (N_48184,N_47730,N_47648);
or U48185 (N_48185,N_47700,N_47913);
and U48186 (N_48186,N_47587,N_47663);
or U48187 (N_48187,N_47597,N_47753);
nand U48188 (N_48188,N_47736,N_47783);
or U48189 (N_48189,N_47574,N_47550);
and U48190 (N_48190,N_47828,N_47851);
nor U48191 (N_48191,N_47968,N_47617);
xnor U48192 (N_48192,N_47678,N_47980);
or U48193 (N_48193,N_47802,N_47820);
and U48194 (N_48194,N_47889,N_47647);
nand U48195 (N_48195,N_47543,N_47861);
and U48196 (N_48196,N_47622,N_47919);
nor U48197 (N_48197,N_47850,N_47629);
and U48198 (N_48198,N_47552,N_47792);
or U48199 (N_48199,N_47539,N_47800);
nor U48200 (N_48200,N_47661,N_47796);
and U48201 (N_48201,N_47881,N_47838);
nor U48202 (N_48202,N_47759,N_47819);
nand U48203 (N_48203,N_47558,N_47657);
xnor U48204 (N_48204,N_47718,N_47660);
nand U48205 (N_48205,N_47936,N_47628);
xnor U48206 (N_48206,N_47849,N_47531);
and U48207 (N_48207,N_47822,N_47814);
nor U48208 (N_48208,N_47619,N_47639);
nor U48209 (N_48209,N_47880,N_47789);
and U48210 (N_48210,N_47960,N_47598);
or U48211 (N_48211,N_47535,N_47731);
nor U48212 (N_48212,N_47975,N_47891);
xnor U48213 (N_48213,N_47788,N_47924);
xor U48214 (N_48214,N_47571,N_47977);
nor U48215 (N_48215,N_47694,N_47608);
or U48216 (N_48216,N_47540,N_47621);
xnor U48217 (N_48217,N_47993,N_47904);
xnor U48218 (N_48218,N_47624,N_47893);
and U48219 (N_48219,N_47978,N_47580);
xnor U48220 (N_48220,N_47607,N_47500);
or U48221 (N_48221,N_47867,N_47852);
and U48222 (N_48222,N_47716,N_47765);
or U48223 (N_48223,N_47864,N_47921);
nor U48224 (N_48224,N_47537,N_47651);
xnor U48225 (N_48225,N_47627,N_47673);
nand U48226 (N_48226,N_47729,N_47710);
nand U48227 (N_48227,N_47845,N_47882);
xor U48228 (N_48228,N_47841,N_47611);
xor U48229 (N_48229,N_47553,N_47682);
nor U48230 (N_48230,N_47756,N_47609);
or U48231 (N_48231,N_47515,N_47547);
or U48232 (N_48232,N_47666,N_47902);
xnor U48233 (N_48233,N_47996,N_47514);
xnor U48234 (N_48234,N_47706,N_47583);
xnor U48235 (N_48235,N_47548,N_47914);
and U48236 (N_48236,N_47671,N_47916);
nand U48237 (N_48237,N_47886,N_47875);
nor U48238 (N_48238,N_47521,N_47749);
or U48239 (N_48239,N_47697,N_47981);
and U48240 (N_48240,N_47824,N_47645);
nand U48241 (N_48241,N_47927,N_47806);
nor U48242 (N_48242,N_47566,N_47635);
nor U48243 (N_48243,N_47899,N_47955);
and U48244 (N_48244,N_47969,N_47781);
nor U48245 (N_48245,N_47505,N_47699);
nor U48246 (N_48246,N_47957,N_47576);
nor U48247 (N_48247,N_47833,N_47691);
nor U48248 (N_48248,N_47952,N_47744);
or U48249 (N_48249,N_47995,N_47590);
nand U48250 (N_48250,N_47755,N_47935);
xnor U48251 (N_48251,N_47696,N_47961);
nand U48252 (N_48252,N_47652,N_47998);
or U48253 (N_48253,N_47684,N_47729);
xor U48254 (N_48254,N_47856,N_47738);
xor U48255 (N_48255,N_47502,N_47973);
xor U48256 (N_48256,N_47940,N_47968);
nor U48257 (N_48257,N_47948,N_47655);
and U48258 (N_48258,N_47750,N_47665);
and U48259 (N_48259,N_47679,N_47783);
or U48260 (N_48260,N_47972,N_47909);
nor U48261 (N_48261,N_47606,N_47759);
and U48262 (N_48262,N_47987,N_47733);
nand U48263 (N_48263,N_47804,N_47643);
nand U48264 (N_48264,N_47712,N_47869);
xnor U48265 (N_48265,N_47852,N_47883);
and U48266 (N_48266,N_47689,N_47840);
or U48267 (N_48267,N_47797,N_47656);
xor U48268 (N_48268,N_47994,N_47674);
xnor U48269 (N_48269,N_47947,N_47869);
or U48270 (N_48270,N_47645,N_47623);
xnor U48271 (N_48271,N_47782,N_47818);
or U48272 (N_48272,N_47809,N_47678);
nand U48273 (N_48273,N_47655,N_47722);
xor U48274 (N_48274,N_47625,N_47657);
nor U48275 (N_48275,N_47568,N_47528);
or U48276 (N_48276,N_47659,N_47997);
or U48277 (N_48277,N_47608,N_47642);
and U48278 (N_48278,N_47730,N_47638);
or U48279 (N_48279,N_47555,N_47958);
or U48280 (N_48280,N_47584,N_47725);
nor U48281 (N_48281,N_47809,N_47607);
and U48282 (N_48282,N_47724,N_47642);
or U48283 (N_48283,N_47770,N_47666);
xnor U48284 (N_48284,N_47703,N_47914);
nor U48285 (N_48285,N_47751,N_47805);
and U48286 (N_48286,N_47686,N_47664);
xor U48287 (N_48287,N_47519,N_47887);
or U48288 (N_48288,N_47921,N_47946);
nor U48289 (N_48289,N_47614,N_47633);
nand U48290 (N_48290,N_47798,N_47779);
nor U48291 (N_48291,N_47662,N_47546);
nor U48292 (N_48292,N_47919,N_47511);
or U48293 (N_48293,N_47744,N_47849);
nor U48294 (N_48294,N_47585,N_47519);
xor U48295 (N_48295,N_47729,N_47711);
nand U48296 (N_48296,N_47963,N_47712);
or U48297 (N_48297,N_47846,N_47780);
nand U48298 (N_48298,N_47925,N_47666);
xnor U48299 (N_48299,N_47940,N_47867);
nor U48300 (N_48300,N_47952,N_47542);
nor U48301 (N_48301,N_47606,N_47682);
and U48302 (N_48302,N_47726,N_47861);
or U48303 (N_48303,N_47708,N_47868);
nor U48304 (N_48304,N_47721,N_47597);
or U48305 (N_48305,N_47905,N_47746);
and U48306 (N_48306,N_47950,N_47967);
and U48307 (N_48307,N_47787,N_47687);
or U48308 (N_48308,N_47527,N_47757);
xor U48309 (N_48309,N_47591,N_47784);
nand U48310 (N_48310,N_47979,N_47625);
and U48311 (N_48311,N_47654,N_47992);
xor U48312 (N_48312,N_47992,N_47689);
or U48313 (N_48313,N_47559,N_47953);
or U48314 (N_48314,N_47992,N_47877);
or U48315 (N_48315,N_47853,N_47816);
or U48316 (N_48316,N_47717,N_47856);
nor U48317 (N_48317,N_47736,N_47576);
nand U48318 (N_48318,N_47556,N_47867);
and U48319 (N_48319,N_47651,N_47842);
or U48320 (N_48320,N_47588,N_47766);
and U48321 (N_48321,N_47643,N_47906);
or U48322 (N_48322,N_47731,N_47564);
nand U48323 (N_48323,N_47850,N_47557);
nand U48324 (N_48324,N_47734,N_47698);
nor U48325 (N_48325,N_47867,N_47724);
xor U48326 (N_48326,N_47592,N_47675);
and U48327 (N_48327,N_47767,N_47629);
xnor U48328 (N_48328,N_47870,N_47931);
and U48329 (N_48329,N_47575,N_47950);
nand U48330 (N_48330,N_47668,N_47569);
xnor U48331 (N_48331,N_47956,N_47766);
nor U48332 (N_48332,N_47739,N_47825);
nor U48333 (N_48333,N_47760,N_47743);
nand U48334 (N_48334,N_47642,N_47685);
nor U48335 (N_48335,N_47646,N_47626);
or U48336 (N_48336,N_47788,N_47833);
and U48337 (N_48337,N_47513,N_47739);
or U48338 (N_48338,N_47521,N_47766);
xnor U48339 (N_48339,N_47767,N_47947);
xnor U48340 (N_48340,N_47736,N_47599);
nor U48341 (N_48341,N_47510,N_47843);
nand U48342 (N_48342,N_47859,N_47960);
nand U48343 (N_48343,N_47663,N_47614);
nand U48344 (N_48344,N_47664,N_47950);
xnor U48345 (N_48345,N_47753,N_47687);
xnor U48346 (N_48346,N_47580,N_47739);
nor U48347 (N_48347,N_47749,N_47635);
and U48348 (N_48348,N_47755,N_47945);
or U48349 (N_48349,N_47781,N_47752);
and U48350 (N_48350,N_47547,N_47723);
or U48351 (N_48351,N_47815,N_47818);
nand U48352 (N_48352,N_47812,N_47973);
xor U48353 (N_48353,N_47822,N_47767);
and U48354 (N_48354,N_47863,N_47816);
or U48355 (N_48355,N_47812,N_47507);
xor U48356 (N_48356,N_47831,N_47714);
or U48357 (N_48357,N_47901,N_47816);
and U48358 (N_48358,N_47755,N_47786);
nor U48359 (N_48359,N_47747,N_47574);
or U48360 (N_48360,N_47665,N_47953);
and U48361 (N_48361,N_47829,N_47723);
or U48362 (N_48362,N_47861,N_47794);
xor U48363 (N_48363,N_47643,N_47655);
nand U48364 (N_48364,N_47655,N_47911);
xnor U48365 (N_48365,N_47715,N_47694);
and U48366 (N_48366,N_47682,N_47861);
nand U48367 (N_48367,N_47755,N_47789);
and U48368 (N_48368,N_47527,N_47522);
xor U48369 (N_48369,N_47774,N_47843);
nor U48370 (N_48370,N_47778,N_47984);
nor U48371 (N_48371,N_47899,N_47528);
or U48372 (N_48372,N_47541,N_47759);
nand U48373 (N_48373,N_47712,N_47533);
nor U48374 (N_48374,N_47834,N_47833);
and U48375 (N_48375,N_47795,N_47906);
and U48376 (N_48376,N_47679,N_47882);
or U48377 (N_48377,N_47770,N_47882);
and U48378 (N_48378,N_47934,N_47815);
nand U48379 (N_48379,N_47870,N_47903);
xor U48380 (N_48380,N_47718,N_47851);
nor U48381 (N_48381,N_47864,N_47840);
xor U48382 (N_48382,N_47782,N_47866);
nor U48383 (N_48383,N_47586,N_47645);
nor U48384 (N_48384,N_47822,N_47852);
or U48385 (N_48385,N_47766,N_47595);
or U48386 (N_48386,N_47632,N_47906);
nand U48387 (N_48387,N_47750,N_47745);
nor U48388 (N_48388,N_47843,N_47683);
nand U48389 (N_48389,N_47822,N_47634);
xnor U48390 (N_48390,N_47597,N_47552);
nand U48391 (N_48391,N_47796,N_47663);
xor U48392 (N_48392,N_47902,N_47755);
or U48393 (N_48393,N_47978,N_47635);
nand U48394 (N_48394,N_47722,N_47697);
xnor U48395 (N_48395,N_47623,N_47833);
nand U48396 (N_48396,N_47665,N_47741);
nand U48397 (N_48397,N_47833,N_47636);
or U48398 (N_48398,N_47956,N_47753);
nand U48399 (N_48399,N_47601,N_47577);
xor U48400 (N_48400,N_47584,N_47807);
xor U48401 (N_48401,N_47729,N_47828);
and U48402 (N_48402,N_47830,N_47688);
nor U48403 (N_48403,N_47862,N_47846);
nor U48404 (N_48404,N_47608,N_47969);
nand U48405 (N_48405,N_47876,N_47810);
nor U48406 (N_48406,N_47928,N_47536);
or U48407 (N_48407,N_47532,N_47932);
nor U48408 (N_48408,N_47580,N_47953);
xnor U48409 (N_48409,N_47627,N_47776);
and U48410 (N_48410,N_47646,N_47873);
or U48411 (N_48411,N_47916,N_47922);
or U48412 (N_48412,N_47676,N_47831);
xnor U48413 (N_48413,N_47719,N_47507);
nand U48414 (N_48414,N_47878,N_47621);
nor U48415 (N_48415,N_47634,N_47900);
nor U48416 (N_48416,N_47762,N_47618);
and U48417 (N_48417,N_47878,N_47526);
and U48418 (N_48418,N_47951,N_47817);
nand U48419 (N_48419,N_47810,N_47929);
or U48420 (N_48420,N_47749,N_47996);
and U48421 (N_48421,N_47888,N_47789);
xnor U48422 (N_48422,N_47929,N_47570);
or U48423 (N_48423,N_47628,N_47647);
xor U48424 (N_48424,N_47863,N_47538);
or U48425 (N_48425,N_47944,N_47899);
xor U48426 (N_48426,N_47690,N_47794);
and U48427 (N_48427,N_47955,N_47916);
and U48428 (N_48428,N_47950,N_47728);
nor U48429 (N_48429,N_47520,N_47582);
or U48430 (N_48430,N_47594,N_47994);
xnor U48431 (N_48431,N_47781,N_47667);
or U48432 (N_48432,N_47941,N_47588);
xnor U48433 (N_48433,N_47505,N_47984);
xnor U48434 (N_48434,N_47901,N_47971);
xor U48435 (N_48435,N_47635,N_47602);
or U48436 (N_48436,N_47568,N_47592);
xor U48437 (N_48437,N_47680,N_47737);
xnor U48438 (N_48438,N_47991,N_47601);
nor U48439 (N_48439,N_47879,N_47797);
xor U48440 (N_48440,N_47877,N_47836);
nor U48441 (N_48441,N_47763,N_47681);
nand U48442 (N_48442,N_47734,N_47877);
or U48443 (N_48443,N_47546,N_47725);
nor U48444 (N_48444,N_47516,N_47767);
or U48445 (N_48445,N_47655,N_47994);
or U48446 (N_48446,N_47965,N_47527);
or U48447 (N_48447,N_47840,N_47672);
and U48448 (N_48448,N_47703,N_47633);
or U48449 (N_48449,N_47987,N_47714);
and U48450 (N_48450,N_47905,N_47548);
or U48451 (N_48451,N_47757,N_47552);
xnor U48452 (N_48452,N_47704,N_47918);
or U48453 (N_48453,N_47772,N_47752);
xnor U48454 (N_48454,N_47616,N_47995);
and U48455 (N_48455,N_47795,N_47675);
and U48456 (N_48456,N_47504,N_47641);
nand U48457 (N_48457,N_47871,N_47717);
nor U48458 (N_48458,N_47814,N_47984);
nand U48459 (N_48459,N_47955,N_47683);
and U48460 (N_48460,N_47917,N_47675);
nand U48461 (N_48461,N_47712,N_47730);
xnor U48462 (N_48462,N_47543,N_47501);
nor U48463 (N_48463,N_47973,N_47524);
and U48464 (N_48464,N_47550,N_47541);
nor U48465 (N_48465,N_47957,N_47708);
nand U48466 (N_48466,N_47528,N_47642);
and U48467 (N_48467,N_47535,N_47507);
nor U48468 (N_48468,N_47731,N_47927);
nand U48469 (N_48469,N_47613,N_47656);
nand U48470 (N_48470,N_47811,N_47624);
or U48471 (N_48471,N_47660,N_47939);
nand U48472 (N_48472,N_47614,N_47807);
and U48473 (N_48473,N_47656,N_47984);
or U48474 (N_48474,N_47950,N_47919);
nand U48475 (N_48475,N_47749,N_47995);
nor U48476 (N_48476,N_47804,N_47742);
nor U48477 (N_48477,N_47658,N_47693);
nor U48478 (N_48478,N_47900,N_47670);
nor U48479 (N_48479,N_47949,N_47959);
or U48480 (N_48480,N_47933,N_47587);
and U48481 (N_48481,N_47865,N_47625);
nor U48482 (N_48482,N_47781,N_47831);
and U48483 (N_48483,N_47680,N_47793);
or U48484 (N_48484,N_47570,N_47594);
nand U48485 (N_48485,N_47721,N_47910);
or U48486 (N_48486,N_47583,N_47599);
xnor U48487 (N_48487,N_47604,N_47781);
xor U48488 (N_48488,N_47914,N_47670);
or U48489 (N_48489,N_47584,N_47744);
nor U48490 (N_48490,N_47534,N_47821);
and U48491 (N_48491,N_47911,N_47728);
nand U48492 (N_48492,N_47960,N_47764);
nand U48493 (N_48493,N_47514,N_47703);
and U48494 (N_48494,N_47687,N_47997);
and U48495 (N_48495,N_47943,N_47552);
nand U48496 (N_48496,N_47652,N_47922);
and U48497 (N_48497,N_47895,N_47622);
xnor U48498 (N_48498,N_47906,N_47657);
nand U48499 (N_48499,N_47856,N_47616);
nor U48500 (N_48500,N_48438,N_48159);
nor U48501 (N_48501,N_48371,N_48043);
and U48502 (N_48502,N_48423,N_48497);
xor U48503 (N_48503,N_48055,N_48327);
nor U48504 (N_48504,N_48218,N_48446);
nand U48505 (N_48505,N_48053,N_48316);
or U48506 (N_48506,N_48239,N_48168);
nand U48507 (N_48507,N_48472,N_48311);
nand U48508 (N_48508,N_48282,N_48058);
and U48509 (N_48509,N_48137,N_48437);
xor U48510 (N_48510,N_48460,N_48300);
nand U48511 (N_48511,N_48077,N_48443);
nand U48512 (N_48512,N_48075,N_48238);
nand U48513 (N_48513,N_48083,N_48378);
or U48514 (N_48514,N_48246,N_48324);
nor U48515 (N_48515,N_48090,N_48177);
nand U48516 (N_48516,N_48171,N_48136);
and U48517 (N_48517,N_48392,N_48455);
nor U48518 (N_48518,N_48005,N_48457);
nand U48519 (N_48519,N_48045,N_48328);
nor U48520 (N_48520,N_48233,N_48337);
xnor U48521 (N_48521,N_48074,N_48334);
nor U48522 (N_48522,N_48485,N_48073);
xnor U48523 (N_48523,N_48291,N_48336);
xor U48524 (N_48524,N_48139,N_48416);
and U48525 (N_48525,N_48204,N_48130);
xor U48526 (N_48526,N_48338,N_48463);
nor U48527 (N_48527,N_48242,N_48332);
xnor U48528 (N_48528,N_48102,N_48290);
or U48529 (N_48529,N_48088,N_48280);
and U48530 (N_48530,N_48036,N_48142);
nand U48531 (N_48531,N_48361,N_48176);
nor U48532 (N_48532,N_48106,N_48266);
xor U48533 (N_48533,N_48089,N_48192);
nor U48534 (N_48534,N_48217,N_48165);
nor U48535 (N_48535,N_48359,N_48220);
or U48536 (N_48536,N_48293,N_48464);
nand U48537 (N_48537,N_48284,N_48418);
or U48538 (N_48538,N_48317,N_48235);
nor U48539 (N_48539,N_48400,N_48352);
and U48540 (N_48540,N_48279,N_48478);
nor U48541 (N_48541,N_48228,N_48301);
xor U48542 (N_48542,N_48208,N_48350);
xnor U48543 (N_48543,N_48000,N_48281);
nand U48544 (N_48544,N_48329,N_48323);
nand U48545 (N_48545,N_48029,N_48158);
nand U48546 (N_48546,N_48452,N_48013);
xor U48547 (N_48547,N_48333,N_48057);
nand U48548 (N_48548,N_48185,N_48330);
nor U48549 (N_48549,N_48143,N_48188);
or U48550 (N_48550,N_48493,N_48366);
xnor U48551 (N_48551,N_48150,N_48313);
nand U48552 (N_48552,N_48249,N_48288);
xnor U48553 (N_48553,N_48269,N_48014);
nor U48554 (N_48554,N_48436,N_48078);
nand U48555 (N_48555,N_48098,N_48095);
xor U48556 (N_48556,N_48433,N_48321);
nor U48557 (N_48557,N_48212,N_48061);
and U48558 (N_48558,N_48450,N_48383);
xnor U48559 (N_48559,N_48178,N_48174);
xnor U48560 (N_48560,N_48243,N_48357);
nand U48561 (N_48561,N_48345,N_48146);
xor U48562 (N_48562,N_48236,N_48138);
or U48563 (N_48563,N_48064,N_48194);
or U48564 (N_48564,N_48099,N_48270);
and U48565 (N_48565,N_48355,N_48440);
nor U48566 (N_48566,N_48203,N_48035);
xnor U48567 (N_48567,N_48495,N_48002);
nor U48568 (N_48568,N_48369,N_48271);
xor U48569 (N_48569,N_48484,N_48051);
nor U48570 (N_48570,N_48474,N_48109);
and U48571 (N_48571,N_48066,N_48020);
nor U48572 (N_48572,N_48342,N_48386);
nor U48573 (N_48573,N_48145,N_48054);
xor U48574 (N_48574,N_48067,N_48257);
nand U48575 (N_48575,N_48399,N_48219);
xor U48576 (N_48576,N_48287,N_48314);
nor U48577 (N_48577,N_48199,N_48133);
xnor U48578 (N_48578,N_48408,N_48473);
and U48579 (N_48579,N_48286,N_48385);
nor U48580 (N_48580,N_48273,N_48319);
nor U48581 (N_48581,N_48297,N_48475);
and U48582 (N_48582,N_48456,N_48389);
or U48583 (N_48583,N_48004,N_48009);
nor U48584 (N_48584,N_48312,N_48047);
xnor U48585 (N_48585,N_48380,N_48131);
or U48586 (N_48586,N_48122,N_48044);
nor U48587 (N_48587,N_48372,N_48059);
or U48588 (N_48588,N_48458,N_48234);
nand U48589 (N_48589,N_48412,N_48413);
or U48590 (N_48590,N_48011,N_48092);
nand U48591 (N_48591,N_48490,N_48391);
and U48592 (N_48592,N_48190,N_48201);
and U48593 (N_48593,N_48197,N_48492);
nor U48594 (N_48594,N_48015,N_48153);
xor U48595 (N_48595,N_48181,N_48261);
xnor U48596 (N_48596,N_48360,N_48213);
nor U48597 (N_48597,N_48162,N_48172);
nor U48598 (N_48598,N_48275,N_48274);
nand U48599 (N_48599,N_48250,N_48040);
nand U48600 (N_48600,N_48039,N_48193);
xor U48601 (N_48601,N_48259,N_48393);
and U48602 (N_48602,N_48048,N_48227);
nor U48603 (N_48603,N_48435,N_48119);
or U48604 (N_48604,N_48260,N_48224);
or U48605 (N_48605,N_48365,N_48308);
and U48606 (N_48606,N_48071,N_48289);
xnor U48607 (N_48607,N_48094,N_48373);
xor U48608 (N_48608,N_48247,N_48346);
nor U48609 (N_48609,N_48245,N_48395);
and U48610 (N_48610,N_48028,N_48184);
nor U48611 (N_48611,N_48422,N_48255);
and U48612 (N_48612,N_48232,N_48231);
and U48613 (N_48613,N_48498,N_48030);
or U48614 (N_48614,N_48425,N_48396);
or U48615 (N_48615,N_48052,N_48023);
and U48616 (N_48616,N_48295,N_48226);
and U48617 (N_48617,N_48144,N_48430);
and U48618 (N_48618,N_48488,N_48244);
xnor U48619 (N_48619,N_48349,N_48296);
and U48620 (N_48620,N_48241,N_48072);
nor U48621 (N_48621,N_48445,N_48049);
xnor U48622 (N_48622,N_48149,N_48222);
xnor U48623 (N_48623,N_48462,N_48079);
nor U48624 (N_48624,N_48398,N_48363);
and U48625 (N_48625,N_48081,N_48180);
xnor U48626 (N_48626,N_48434,N_48348);
and U48627 (N_48627,N_48367,N_48179);
nand U48628 (N_48628,N_48283,N_48123);
and U48629 (N_48629,N_48344,N_48353);
nand U48630 (N_48630,N_48093,N_48407);
xor U48631 (N_48631,N_48254,N_48421);
nor U48632 (N_48632,N_48128,N_48448);
nor U48633 (N_48633,N_48209,N_48124);
and U48634 (N_48634,N_48496,N_48267);
nor U48635 (N_48635,N_48205,N_48156);
or U48636 (N_48636,N_48277,N_48354);
or U48637 (N_48637,N_48211,N_48410);
xor U48638 (N_48638,N_48129,N_48063);
nand U48639 (N_48639,N_48467,N_48263);
nand U48640 (N_48640,N_48251,N_48307);
and U48641 (N_48641,N_48070,N_48225);
and U48642 (N_48642,N_48229,N_48304);
nor U48643 (N_48643,N_48026,N_48221);
nor U48644 (N_48644,N_48008,N_48198);
or U48645 (N_48645,N_48351,N_48453);
or U48646 (N_48646,N_48340,N_48499);
nor U48647 (N_48647,N_48157,N_48439);
and U48648 (N_48648,N_48034,N_48134);
or U48649 (N_48649,N_48268,N_48202);
nand U48650 (N_48650,N_48409,N_48085);
xor U48651 (N_48651,N_48031,N_48292);
and U48652 (N_48652,N_48170,N_48097);
or U48653 (N_48653,N_48424,N_48294);
xnor U48654 (N_48654,N_48147,N_48431);
or U48655 (N_48655,N_48082,N_48169);
or U48656 (N_48656,N_48022,N_48406);
xor U48657 (N_48657,N_48096,N_48486);
nand U48658 (N_48658,N_48309,N_48050);
xnor U48659 (N_48659,N_48320,N_48021);
or U48660 (N_48660,N_48347,N_48414);
nand U48661 (N_48661,N_48163,N_48032);
xnor U48662 (N_48662,N_48384,N_48103);
nand U48663 (N_48663,N_48482,N_48258);
and U48664 (N_48664,N_48299,N_48387);
nor U48665 (N_48665,N_48056,N_48272);
and U48666 (N_48666,N_48120,N_48480);
xor U48667 (N_48667,N_48069,N_48397);
or U48668 (N_48668,N_48335,N_48252);
nand U48669 (N_48669,N_48117,N_48016);
nor U48670 (N_48670,N_48494,N_48491);
nand U48671 (N_48671,N_48166,N_48191);
or U48672 (N_48672,N_48411,N_48368);
and U48673 (N_48673,N_48444,N_48042);
xnor U48674 (N_48674,N_48018,N_48305);
nor U48675 (N_48675,N_48479,N_48285);
nor U48676 (N_48676,N_48449,N_48362);
nand U48677 (N_48677,N_48046,N_48113);
nand U48678 (N_48678,N_48476,N_48404);
or U48679 (N_48679,N_48196,N_48152);
and U48680 (N_48680,N_48326,N_48167);
or U48681 (N_48681,N_48451,N_48216);
nand U48682 (N_48682,N_48186,N_48466);
xor U48683 (N_48683,N_48148,N_48012);
nand U48684 (N_48684,N_48160,N_48265);
and U48685 (N_48685,N_48339,N_48111);
xnor U48686 (N_48686,N_48155,N_48010);
or U48687 (N_48687,N_48356,N_48429);
nand U48688 (N_48688,N_48477,N_48112);
nand U48689 (N_48689,N_48426,N_48127);
and U48690 (N_48690,N_48230,N_48135);
or U48691 (N_48691,N_48187,N_48038);
and U48692 (N_48692,N_48104,N_48182);
nor U48693 (N_48693,N_48033,N_48173);
or U48694 (N_48694,N_48101,N_48164);
nand U48695 (N_48695,N_48427,N_48381);
nor U48696 (N_48696,N_48417,N_48007);
xnor U48697 (N_48697,N_48207,N_48003);
nor U48698 (N_48698,N_48114,N_48256);
and U48699 (N_48699,N_48428,N_48432);
nor U48700 (N_48700,N_48331,N_48200);
or U48701 (N_48701,N_48310,N_48076);
nor U48702 (N_48702,N_48465,N_48405);
and U48703 (N_48703,N_48370,N_48420);
xor U48704 (N_48704,N_48377,N_48390);
or U48705 (N_48705,N_48240,N_48318);
xnor U48706 (N_48706,N_48223,N_48161);
xor U48707 (N_48707,N_48303,N_48116);
nor U48708 (N_48708,N_48062,N_48489);
and U48709 (N_48709,N_48001,N_48419);
nand U48710 (N_48710,N_48306,N_48065);
and U48711 (N_48711,N_48322,N_48132);
nand U48712 (N_48712,N_48262,N_48091);
and U48713 (N_48713,N_48379,N_48401);
nor U48714 (N_48714,N_48403,N_48019);
nor U48715 (N_48715,N_48154,N_48461);
nand U48716 (N_48716,N_48110,N_48105);
nor U48717 (N_48717,N_48175,N_48343);
and U48718 (N_48718,N_48087,N_48100);
nor U48719 (N_48719,N_48121,N_48470);
or U48720 (N_48720,N_48108,N_48402);
nand U48721 (N_48721,N_48382,N_48237);
xor U48722 (N_48722,N_48006,N_48415);
and U48723 (N_48723,N_48454,N_48183);
and U48724 (N_48724,N_48068,N_48017);
nor U48725 (N_48725,N_48298,N_48325);
or U48726 (N_48726,N_48358,N_48487);
or U48727 (N_48727,N_48388,N_48341);
nand U48728 (N_48728,N_48086,N_48469);
or U48729 (N_48729,N_48253,N_48315);
nand U48730 (N_48730,N_48214,N_48302);
and U48731 (N_48731,N_48140,N_48107);
nand U48732 (N_48732,N_48141,N_48151);
or U48733 (N_48733,N_48481,N_48125);
xor U48734 (N_48734,N_48080,N_48195);
xnor U48735 (N_48735,N_48024,N_48206);
or U48736 (N_48736,N_48210,N_48189);
xnor U48737 (N_48737,N_48041,N_48278);
xnor U48738 (N_48738,N_48126,N_48248);
nand U48739 (N_48739,N_48115,N_48364);
nand U48740 (N_48740,N_48375,N_48394);
xor U48741 (N_48741,N_48483,N_48276);
nor U48742 (N_48742,N_48447,N_48025);
and U48743 (N_48743,N_48118,N_48027);
and U48744 (N_48744,N_48374,N_48215);
nand U48745 (N_48745,N_48441,N_48084);
and U48746 (N_48746,N_48471,N_48442);
and U48747 (N_48747,N_48037,N_48468);
or U48748 (N_48748,N_48459,N_48264);
or U48749 (N_48749,N_48060,N_48376);
and U48750 (N_48750,N_48425,N_48278);
nand U48751 (N_48751,N_48042,N_48265);
nand U48752 (N_48752,N_48150,N_48051);
nor U48753 (N_48753,N_48351,N_48271);
nor U48754 (N_48754,N_48300,N_48195);
and U48755 (N_48755,N_48023,N_48447);
or U48756 (N_48756,N_48227,N_48117);
nand U48757 (N_48757,N_48058,N_48006);
xor U48758 (N_48758,N_48431,N_48375);
xor U48759 (N_48759,N_48226,N_48017);
xor U48760 (N_48760,N_48098,N_48403);
nand U48761 (N_48761,N_48485,N_48493);
nor U48762 (N_48762,N_48147,N_48293);
and U48763 (N_48763,N_48136,N_48472);
nand U48764 (N_48764,N_48023,N_48338);
and U48765 (N_48765,N_48405,N_48299);
nand U48766 (N_48766,N_48436,N_48195);
xor U48767 (N_48767,N_48302,N_48476);
nor U48768 (N_48768,N_48330,N_48427);
and U48769 (N_48769,N_48040,N_48232);
nor U48770 (N_48770,N_48350,N_48432);
xnor U48771 (N_48771,N_48157,N_48126);
nand U48772 (N_48772,N_48320,N_48372);
and U48773 (N_48773,N_48024,N_48497);
xnor U48774 (N_48774,N_48009,N_48225);
nor U48775 (N_48775,N_48348,N_48034);
and U48776 (N_48776,N_48200,N_48035);
or U48777 (N_48777,N_48018,N_48104);
xnor U48778 (N_48778,N_48161,N_48185);
or U48779 (N_48779,N_48490,N_48281);
and U48780 (N_48780,N_48256,N_48060);
nand U48781 (N_48781,N_48017,N_48230);
nand U48782 (N_48782,N_48290,N_48497);
xor U48783 (N_48783,N_48339,N_48132);
nand U48784 (N_48784,N_48251,N_48341);
and U48785 (N_48785,N_48256,N_48103);
nand U48786 (N_48786,N_48291,N_48444);
and U48787 (N_48787,N_48166,N_48203);
or U48788 (N_48788,N_48179,N_48413);
xnor U48789 (N_48789,N_48207,N_48253);
nand U48790 (N_48790,N_48216,N_48260);
nand U48791 (N_48791,N_48426,N_48265);
and U48792 (N_48792,N_48099,N_48139);
nor U48793 (N_48793,N_48174,N_48203);
and U48794 (N_48794,N_48372,N_48054);
or U48795 (N_48795,N_48066,N_48445);
or U48796 (N_48796,N_48225,N_48165);
or U48797 (N_48797,N_48202,N_48436);
nor U48798 (N_48798,N_48393,N_48231);
and U48799 (N_48799,N_48480,N_48472);
nand U48800 (N_48800,N_48360,N_48075);
and U48801 (N_48801,N_48338,N_48063);
xor U48802 (N_48802,N_48422,N_48386);
nor U48803 (N_48803,N_48081,N_48173);
xor U48804 (N_48804,N_48302,N_48430);
nor U48805 (N_48805,N_48420,N_48403);
xor U48806 (N_48806,N_48155,N_48435);
nor U48807 (N_48807,N_48442,N_48433);
nor U48808 (N_48808,N_48149,N_48323);
xor U48809 (N_48809,N_48345,N_48030);
and U48810 (N_48810,N_48086,N_48206);
nand U48811 (N_48811,N_48342,N_48332);
nand U48812 (N_48812,N_48394,N_48212);
nor U48813 (N_48813,N_48047,N_48020);
nand U48814 (N_48814,N_48281,N_48460);
nor U48815 (N_48815,N_48157,N_48086);
or U48816 (N_48816,N_48372,N_48255);
nor U48817 (N_48817,N_48248,N_48472);
nand U48818 (N_48818,N_48376,N_48192);
nor U48819 (N_48819,N_48442,N_48452);
and U48820 (N_48820,N_48288,N_48458);
xor U48821 (N_48821,N_48147,N_48377);
or U48822 (N_48822,N_48445,N_48432);
nand U48823 (N_48823,N_48137,N_48286);
xnor U48824 (N_48824,N_48215,N_48135);
and U48825 (N_48825,N_48315,N_48367);
or U48826 (N_48826,N_48439,N_48115);
and U48827 (N_48827,N_48358,N_48132);
and U48828 (N_48828,N_48239,N_48218);
nand U48829 (N_48829,N_48027,N_48101);
and U48830 (N_48830,N_48167,N_48455);
and U48831 (N_48831,N_48321,N_48303);
and U48832 (N_48832,N_48275,N_48218);
nand U48833 (N_48833,N_48244,N_48324);
or U48834 (N_48834,N_48462,N_48025);
nor U48835 (N_48835,N_48174,N_48181);
nor U48836 (N_48836,N_48432,N_48381);
nand U48837 (N_48837,N_48475,N_48375);
or U48838 (N_48838,N_48140,N_48209);
nor U48839 (N_48839,N_48072,N_48220);
nand U48840 (N_48840,N_48267,N_48241);
and U48841 (N_48841,N_48473,N_48025);
nor U48842 (N_48842,N_48221,N_48493);
xnor U48843 (N_48843,N_48046,N_48470);
nand U48844 (N_48844,N_48237,N_48399);
nor U48845 (N_48845,N_48127,N_48130);
nor U48846 (N_48846,N_48480,N_48482);
nor U48847 (N_48847,N_48305,N_48114);
and U48848 (N_48848,N_48104,N_48069);
nand U48849 (N_48849,N_48117,N_48356);
nor U48850 (N_48850,N_48470,N_48377);
nand U48851 (N_48851,N_48165,N_48144);
nor U48852 (N_48852,N_48022,N_48415);
xor U48853 (N_48853,N_48004,N_48246);
nand U48854 (N_48854,N_48125,N_48091);
or U48855 (N_48855,N_48495,N_48405);
or U48856 (N_48856,N_48447,N_48387);
nor U48857 (N_48857,N_48281,N_48179);
nand U48858 (N_48858,N_48168,N_48344);
nand U48859 (N_48859,N_48017,N_48196);
xor U48860 (N_48860,N_48232,N_48368);
or U48861 (N_48861,N_48074,N_48245);
and U48862 (N_48862,N_48490,N_48404);
xnor U48863 (N_48863,N_48247,N_48102);
nand U48864 (N_48864,N_48302,N_48010);
nand U48865 (N_48865,N_48238,N_48174);
nor U48866 (N_48866,N_48187,N_48204);
xnor U48867 (N_48867,N_48494,N_48098);
nor U48868 (N_48868,N_48217,N_48237);
or U48869 (N_48869,N_48168,N_48002);
xor U48870 (N_48870,N_48204,N_48383);
nand U48871 (N_48871,N_48290,N_48135);
and U48872 (N_48872,N_48364,N_48317);
nand U48873 (N_48873,N_48151,N_48278);
nor U48874 (N_48874,N_48161,N_48085);
xnor U48875 (N_48875,N_48071,N_48197);
xor U48876 (N_48876,N_48397,N_48155);
xnor U48877 (N_48877,N_48175,N_48122);
nor U48878 (N_48878,N_48488,N_48340);
or U48879 (N_48879,N_48442,N_48287);
or U48880 (N_48880,N_48408,N_48314);
nand U48881 (N_48881,N_48490,N_48147);
or U48882 (N_48882,N_48147,N_48344);
or U48883 (N_48883,N_48432,N_48333);
nor U48884 (N_48884,N_48016,N_48362);
nand U48885 (N_48885,N_48428,N_48368);
nor U48886 (N_48886,N_48005,N_48323);
xnor U48887 (N_48887,N_48423,N_48325);
nand U48888 (N_48888,N_48156,N_48184);
nand U48889 (N_48889,N_48062,N_48264);
nor U48890 (N_48890,N_48176,N_48032);
nand U48891 (N_48891,N_48038,N_48291);
nand U48892 (N_48892,N_48484,N_48305);
xor U48893 (N_48893,N_48425,N_48288);
nor U48894 (N_48894,N_48320,N_48376);
xor U48895 (N_48895,N_48171,N_48440);
nor U48896 (N_48896,N_48285,N_48373);
or U48897 (N_48897,N_48235,N_48150);
and U48898 (N_48898,N_48321,N_48195);
nand U48899 (N_48899,N_48079,N_48223);
xnor U48900 (N_48900,N_48469,N_48310);
nand U48901 (N_48901,N_48444,N_48269);
nand U48902 (N_48902,N_48013,N_48167);
or U48903 (N_48903,N_48167,N_48145);
and U48904 (N_48904,N_48456,N_48175);
and U48905 (N_48905,N_48480,N_48497);
or U48906 (N_48906,N_48359,N_48288);
nor U48907 (N_48907,N_48119,N_48282);
xor U48908 (N_48908,N_48061,N_48036);
nor U48909 (N_48909,N_48128,N_48389);
xor U48910 (N_48910,N_48056,N_48126);
and U48911 (N_48911,N_48436,N_48132);
and U48912 (N_48912,N_48303,N_48164);
or U48913 (N_48913,N_48014,N_48081);
xor U48914 (N_48914,N_48032,N_48409);
nand U48915 (N_48915,N_48258,N_48022);
xor U48916 (N_48916,N_48388,N_48024);
nand U48917 (N_48917,N_48436,N_48385);
nand U48918 (N_48918,N_48215,N_48055);
nand U48919 (N_48919,N_48221,N_48242);
xnor U48920 (N_48920,N_48484,N_48338);
xor U48921 (N_48921,N_48334,N_48382);
and U48922 (N_48922,N_48133,N_48182);
nor U48923 (N_48923,N_48208,N_48036);
nand U48924 (N_48924,N_48428,N_48237);
xnor U48925 (N_48925,N_48234,N_48023);
and U48926 (N_48926,N_48266,N_48021);
xnor U48927 (N_48927,N_48324,N_48363);
xor U48928 (N_48928,N_48386,N_48086);
xnor U48929 (N_48929,N_48154,N_48123);
or U48930 (N_48930,N_48017,N_48112);
or U48931 (N_48931,N_48011,N_48327);
xor U48932 (N_48932,N_48131,N_48294);
or U48933 (N_48933,N_48398,N_48315);
and U48934 (N_48934,N_48058,N_48187);
nand U48935 (N_48935,N_48328,N_48450);
xnor U48936 (N_48936,N_48473,N_48067);
xnor U48937 (N_48937,N_48392,N_48376);
xnor U48938 (N_48938,N_48391,N_48005);
nor U48939 (N_48939,N_48271,N_48273);
and U48940 (N_48940,N_48020,N_48447);
nor U48941 (N_48941,N_48189,N_48030);
xor U48942 (N_48942,N_48484,N_48102);
and U48943 (N_48943,N_48059,N_48240);
xnor U48944 (N_48944,N_48225,N_48012);
or U48945 (N_48945,N_48461,N_48419);
nand U48946 (N_48946,N_48155,N_48289);
nor U48947 (N_48947,N_48007,N_48487);
or U48948 (N_48948,N_48313,N_48498);
nand U48949 (N_48949,N_48094,N_48257);
nor U48950 (N_48950,N_48361,N_48367);
nand U48951 (N_48951,N_48395,N_48447);
nor U48952 (N_48952,N_48144,N_48319);
or U48953 (N_48953,N_48081,N_48151);
xnor U48954 (N_48954,N_48228,N_48328);
or U48955 (N_48955,N_48180,N_48444);
xor U48956 (N_48956,N_48275,N_48193);
or U48957 (N_48957,N_48212,N_48475);
and U48958 (N_48958,N_48298,N_48313);
nor U48959 (N_48959,N_48150,N_48271);
nand U48960 (N_48960,N_48397,N_48061);
xor U48961 (N_48961,N_48336,N_48173);
nand U48962 (N_48962,N_48375,N_48224);
nand U48963 (N_48963,N_48436,N_48488);
xor U48964 (N_48964,N_48107,N_48392);
or U48965 (N_48965,N_48429,N_48137);
xor U48966 (N_48966,N_48060,N_48331);
and U48967 (N_48967,N_48080,N_48491);
or U48968 (N_48968,N_48158,N_48294);
and U48969 (N_48969,N_48174,N_48427);
xor U48970 (N_48970,N_48445,N_48232);
xnor U48971 (N_48971,N_48017,N_48474);
and U48972 (N_48972,N_48452,N_48363);
or U48973 (N_48973,N_48448,N_48023);
or U48974 (N_48974,N_48130,N_48421);
nand U48975 (N_48975,N_48051,N_48045);
and U48976 (N_48976,N_48111,N_48423);
or U48977 (N_48977,N_48089,N_48232);
or U48978 (N_48978,N_48272,N_48413);
and U48979 (N_48979,N_48161,N_48397);
nand U48980 (N_48980,N_48323,N_48264);
and U48981 (N_48981,N_48073,N_48456);
and U48982 (N_48982,N_48137,N_48168);
nor U48983 (N_48983,N_48197,N_48156);
nor U48984 (N_48984,N_48471,N_48044);
xnor U48985 (N_48985,N_48175,N_48078);
nand U48986 (N_48986,N_48168,N_48076);
nand U48987 (N_48987,N_48141,N_48066);
nor U48988 (N_48988,N_48297,N_48014);
and U48989 (N_48989,N_48154,N_48300);
xor U48990 (N_48990,N_48472,N_48299);
xor U48991 (N_48991,N_48186,N_48114);
nand U48992 (N_48992,N_48212,N_48231);
and U48993 (N_48993,N_48241,N_48338);
and U48994 (N_48994,N_48454,N_48133);
xor U48995 (N_48995,N_48018,N_48121);
nor U48996 (N_48996,N_48084,N_48039);
or U48997 (N_48997,N_48482,N_48474);
and U48998 (N_48998,N_48166,N_48057);
xor U48999 (N_48999,N_48030,N_48096);
or U49000 (N_49000,N_48849,N_48564);
or U49001 (N_49001,N_48923,N_48741);
or U49002 (N_49002,N_48649,N_48531);
nor U49003 (N_49003,N_48569,N_48855);
xor U49004 (N_49004,N_48537,N_48573);
or U49005 (N_49005,N_48613,N_48610);
and U49006 (N_49006,N_48747,N_48919);
and U49007 (N_49007,N_48520,N_48935);
nand U49008 (N_49008,N_48570,N_48699);
xnor U49009 (N_49009,N_48571,N_48836);
or U49010 (N_49010,N_48921,N_48828);
nand U49011 (N_49011,N_48586,N_48793);
xor U49012 (N_49012,N_48985,N_48763);
and U49013 (N_49013,N_48915,N_48731);
nand U49014 (N_49014,N_48994,N_48627);
xnor U49015 (N_49015,N_48865,N_48956);
nand U49016 (N_49016,N_48727,N_48660);
nand U49017 (N_49017,N_48834,N_48514);
nor U49018 (N_49018,N_48628,N_48854);
or U49019 (N_49019,N_48951,N_48847);
nor U49020 (N_49020,N_48942,N_48823);
xnor U49021 (N_49021,N_48687,N_48709);
nor U49022 (N_49022,N_48639,N_48661);
and U49023 (N_49023,N_48707,N_48995);
and U49024 (N_49024,N_48901,N_48533);
xor U49025 (N_49025,N_48593,N_48601);
nor U49026 (N_49026,N_48954,N_48623);
and U49027 (N_49027,N_48987,N_48524);
and U49028 (N_49028,N_48812,N_48736);
nor U49029 (N_49029,N_48842,N_48883);
xnor U49030 (N_49030,N_48800,N_48578);
xnor U49031 (N_49031,N_48637,N_48924);
nor U49032 (N_49032,N_48691,N_48519);
and U49033 (N_49033,N_48965,N_48549);
or U49034 (N_49034,N_48887,N_48587);
or U49035 (N_49035,N_48698,N_48650);
xnor U49036 (N_49036,N_48960,N_48890);
or U49037 (N_49037,N_48703,N_48543);
and U49038 (N_49038,N_48645,N_48635);
xnor U49039 (N_49039,N_48723,N_48590);
or U49040 (N_49040,N_48600,N_48974);
nand U49041 (N_49041,N_48766,N_48585);
xor U49042 (N_49042,N_48922,N_48563);
or U49043 (N_49043,N_48932,N_48872);
nand U49044 (N_49044,N_48721,N_48595);
and U49045 (N_49045,N_48534,N_48668);
or U49046 (N_49046,N_48512,N_48925);
and U49047 (N_49047,N_48827,N_48545);
or U49048 (N_49048,N_48914,N_48976);
nor U49049 (N_49049,N_48769,N_48981);
xor U49050 (N_49050,N_48523,N_48990);
nand U49051 (N_49051,N_48943,N_48695);
nor U49052 (N_49052,N_48562,N_48806);
xnor U49053 (N_49053,N_48809,N_48666);
and U49054 (N_49054,N_48936,N_48715);
and U49055 (N_49055,N_48756,N_48556);
nand U49056 (N_49056,N_48605,N_48513);
nand U49057 (N_49057,N_48770,N_48778);
and U49058 (N_49058,N_48900,N_48930);
and U49059 (N_49059,N_48546,N_48833);
xnor U49060 (N_49060,N_48962,N_48878);
xor U49061 (N_49061,N_48853,N_48724);
and U49062 (N_49062,N_48944,N_48726);
nand U49063 (N_49063,N_48801,N_48680);
or U49064 (N_49064,N_48898,N_48772);
or U49065 (N_49065,N_48704,N_48642);
nor U49066 (N_49066,N_48711,N_48963);
nand U49067 (N_49067,N_48961,N_48577);
xnor U49068 (N_49068,N_48893,N_48767);
and U49069 (N_49069,N_48619,N_48941);
xor U49070 (N_49070,N_48819,N_48748);
and U49071 (N_49071,N_48972,N_48988);
nand U49072 (N_49072,N_48894,N_48896);
nand U49073 (N_49073,N_48567,N_48810);
xnor U49074 (N_49074,N_48581,N_48592);
or U49075 (N_49075,N_48621,N_48576);
xor U49076 (N_49076,N_48818,N_48575);
xor U49077 (N_49077,N_48572,N_48653);
nand U49078 (N_49078,N_48760,N_48967);
nor U49079 (N_49079,N_48751,N_48879);
nor U49080 (N_49080,N_48630,N_48913);
and U49081 (N_49081,N_48937,N_48688);
nand U49082 (N_49082,N_48841,N_48622);
xor U49083 (N_49083,N_48808,N_48968);
nand U49084 (N_49084,N_48732,N_48996);
nor U49085 (N_49085,N_48651,N_48978);
nand U49086 (N_49086,N_48897,N_48529);
nor U49087 (N_49087,N_48881,N_48904);
xnor U49088 (N_49088,N_48507,N_48796);
or U49089 (N_49089,N_48541,N_48658);
xnor U49090 (N_49090,N_48905,N_48648);
and U49091 (N_49091,N_48501,N_48544);
or U49092 (N_49092,N_48993,N_48617);
nor U49093 (N_49093,N_48557,N_48877);
xnor U49094 (N_49094,N_48862,N_48844);
and U49095 (N_49095,N_48782,N_48934);
xnor U49096 (N_49096,N_48977,N_48591);
nand U49097 (N_49097,N_48735,N_48843);
or U49098 (N_49098,N_48874,N_48582);
xnor U49099 (N_49099,N_48789,N_48588);
or U49100 (N_49100,N_48596,N_48697);
xor U49101 (N_49101,N_48710,N_48989);
xnor U49102 (N_49102,N_48521,N_48560);
xor U49103 (N_49103,N_48532,N_48912);
or U49104 (N_49104,N_48868,N_48788);
nand U49105 (N_49105,N_48850,N_48685);
or U49106 (N_49106,N_48720,N_48526);
nand U49107 (N_49107,N_48714,N_48670);
nand U49108 (N_49108,N_48550,N_48784);
and U49109 (N_49109,N_48927,N_48656);
nor U49110 (N_49110,N_48753,N_48774);
or U49111 (N_49111,N_48603,N_48826);
nor U49112 (N_49112,N_48555,N_48831);
nand U49113 (N_49113,N_48616,N_48597);
or U49114 (N_49114,N_48908,N_48970);
nor U49115 (N_49115,N_48739,N_48502);
nand U49116 (N_49116,N_48690,N_48561);
or U49117 (N_49117,N_48848,N_48629);
xnor U49118 (N_49118,N_48762,N_48719);
nand U49119 (N_49119,N_48676,N_48667);
nor U49120 (N_49120,N_48536,N_48539);
or U49121 (N_49121,N_48955,N_48787);
or U49122 (N_49122,N_48683,N_48505);
nor U49123 (N_49123,N_48939,N_48821);
xnor U49124 (N_49124,N_48798,N_48920);
and U49125 (N_49125,N_48659,N_48750);
nand U49126 (N_49126,N_48779,N_48681);
or U49127 (N_49127,N_48712,N_48693);
xor U49128 (N_49128,N_48559,N_48895);
nor U49129 (N_49129,N_48705,N_48509);
and U49130 (N_49130,N_48515,N_48547);
nand U49131 (N_49131,N_48986,N_48641);
or U49132 (N_49132,N_48644,N_48608);
nand U49133 (N_49133,N_48999,N_48737);
and U49134 (N_49134,N_48888,N_48655);
and U49135 (N_49135,N_48729,N_48861);
nand U49136 (N_49136,N_48632,N_48746);
nor U49137 (N_49137,N_48816,N_48949);
and U49138 (N_49138,N_48840,N_48730);
xor U49139 (N_49139,N_48907,N_48566);
nor U49140 (N_49140,N_48633,N_48640);
nand U49141 (N_49141,N_48899,N_48837);
nor U49142 (N_49142,N_48846,N_48643);
and U49143 (N_49143,N_48759,N_48947);
xnor U49144 (N_49144,N_48884,N_48579);
nor U49145 (N_49145,N_48752,N_48743);
or U49146 (N_49146,N_48785,N_48946);
xnor U49147 (N_49147,N_48964,N_48672);
nor U49148 (N_49148,N_48889,N_48882);
and U49149 (N_49149,N_48860,N_48984);
xor U49150 (N_49150,N_48832,N_48811);
or U49151 (N_49151,N_48953,N_48876);
or U49152 (N_49152,N_48945,N_48771);
nor U49153 (N_49153,N_48794,N_48506);
or U49154 (N_49154,N_48775,N_48792);
nor U49155 (N_49155,N_48802,N_48742);
and U49156 (N_49156,N_48875,N_48702);
nor U49157 (N_49157,N_48673,N_48991);
xnor U49158 (N_49158,N_48903,N_48754);
xor U49159 (N_49159,N_48599,N_48694);
nand U49160 (N_49160,N_48791,N_48892);
xor U49161 (N_49161,N_48510,N_48538);
xnor U49162 (N_49162,N_48765,N_48745);
and U49163 (N_49163,N_48527,N_48696);
nor U49164 (N_49164,N_48554,N_48508);
or U49165 (N_49165,N_48856,N_48679);
nor U49166 (N_49166,N_48814,N_48869);
nand U49167 (N_49167,N_48646,N_48783);
xor U49168 (N_49168,N_48612,N_48857);
or U49169 (N_49169,N_48503,N_48631);
or U49170 (N_49170,N_48568,N_48535);
nand U49171 (N_49171,N_48761,N_48864);
nand U49172 (N_49172,N_48817,N_48807);
or U49173 (N_49173,N_48528,N_48992);
or U49174 (N_49174,N_48553,N_48665);
and U49175 (N_49175,N_48795,N_48758);
and U49176 (N_49176,N_48799,N_48983);
or U49177 (N_49177,N_48867,N_48609);
nand U49178 (N_49178,N_48825,N_48518);
and U49179 (N_49179,N_48542,N_48552);
or U49180 (N_49180,N_48777,N_48851);
xor U49181 (N_49181,N_48614,N_48606);
xnor U49182 (N_49182,N_48625,N_48873);
xnor U49183 (N_49183,N_48540,N_48734);
or U49184 (N_49184,N_48638,N_48933);
xor U49185 (N_49185,N_48813,N_48708);
or U49186 (N_49186,N_48871,N_48598);
nand U49187 (N_49187,N_48803,N_48626);
nand U49188 (N_49188,N_48839,N_48776);
or U49189 (N_49189,N_48584,N_48551);
nand U49190 (N_49190,N_48716,N_48773);
and U49191 (N_49191,N_48583,N_48845);
nand U49192 (N_49192,N_48940,N_48740);
and U49193 (N_49193,N_48971,N_48815);
or U49194 (N_49194,N_48998,N_48931);
nand U49195 (N_49195,N_48786,N_48652);
xnor U49196 (N_49196,N_48733,N_48558);
or U49197 (N_49197,N_48863,N_48997);
and U49198 (N_49198,N_48669,N_48664);
nor U49199 (N_49199,N_48548,N_48959);
nor U49200 (N_49200,N_48790,N_48725);
nand U49201 (N_49201,N_48738,N_48749);
nor U49202 (N_49202,N_48938,N_48858);
and U49203 (N_49203,N_48700,N_48866);
nor U49204 (N_49204,N_48689,N_48870);
and U49205 (N_49205,N_48701,N_48957);
and U49206 (N_49206,N_48980,N_48969);
nor U49207 (N_49207,N_48657,N_48918);
nand U49208 (N_49208,N_48902,N_48618);
and U49209 (N_49209,N_48718,N_48909);
xnor U49210 (N_49210,N_48911,N_48982);
or U49211 (N_49211,N_48926,N_48910);
xor U49212 (N_49212,N_48973,N_48820);
and U49213 (N_49213,N_48757,N_48602);
or U49214 (N_49214,N_48522,N_48517);
or U49215 (N_49215,N_48859,N_48677);
nor U49216 (N_49216,N_48835,N_48804);
xor U49217 (N_49217,N_48950,N_48636);
and U49218 (N_49218,N_48565,N_48574);
and U49219 (N_49219,N_48675,N_48692);
or U49220 (N_49220,N_48917,N_48829);
and U49221 (N_49221,N_48717,N_48764);
and U49222 (N_49222,N_48830,N_48663);
and U49223 (N_49223,N_48744,N_48580);
xor U49224 (N_49224,N_48928,N_48615);
and U49225 (N_49225,N_48852,N_48500);
nand U49226 (N_49226,N_48885,N_48682);
or U49227 (N_49227,N_48797,N_48511);
or U49228 (N_49228,N_48671,N_48634);
nand U49229 (N_49229,N_48979,N_48781);
nand U49230 (N_49230,N_48891,N_48684);
nand U49231 (N_49231,N_48780,N_48654);
xor U49232 (N_49232,N_48886,N_48768);
nor U49233 (N_49233,N_48838,N_48525);
nor U49234 (N_49234,N_48728,N_48589);
and U49235 (N_49235,N_48755,N_48686);
nor U49236 (N_49236,N_48722,N_48674);
and U49237 (N_49237,N_48713,N_48906);
or U49238 (N_49238,N_48824,N_48805);
nor U49239 (N_49239,N_48880,N_48516);
nand U49240 (N_49240,N_48916,N_48948);
nor U49241 (N_49241,N_48624,N_48620);
nand U49242 (N_49242,N_48975,N_48958);
nand U49243 (N_49243,N_48929,N_48607);
nand U49244 (N_49244,N_48604,N_48647);
xor U49245 (N_49245,N_48611,N_48662);
or U49246 (N_49246,N_48952,N_48822);
nor U49247 (N_49247,N_48594,N_48678);
nor U49248 (N_49248,N_48706,N_48530);
nor U49249 (N_49249,N_48966,N_48504);
nor U49250 (N_49250,N_48650,N_48559);
nand U49251 (N_49251,N_48550,N_48662);
nand U49252 (N_49252,N_48964,N_48644);
nor U49253 (N_49253,N_48899,N_48501);
and U49254 (N_49254,N_48998,N_48823);
and U49255 (N_49255,N_48768,N_48654);
nand U49256 (N_49256,N_48620,N_48693);
or U49257 (N_49257,N_48601,N_48918);
and U49258 (N_49258,N_48510,N_48823);
xor U49259 (N_49259,N_48598,N_48785);
nand U49260 (N_49260,N_48844,N_48845);
nand U49261 (N_49261,N_48756,N_48661);
nand U49262 (N_49262,N_48758,N_48927);
nand U49263 (N_49263,N_48621,N_48953);
or U49264 (N_49264,N_48866,N_48721);
nand U49265 (N_49265,N_48607,N_48644);
nor U49266 (N_49266,N_48512,N_48635);
nand U49267 (N_49267,N_48725,N_48818);
or U49268 (N_49268,N_48987,N_48728);
xor U49269 (N_49269,N_48920,N_48848);
or U49270 (N_49270,N_48618,N_48500);
and U49271 (N_49271,N_48648,N_48675);
xor U49272 (N_49272,N_48529,N_48548);
and U49273 (N_49273,N_48549,N_48534);
xnor U49274 (N_49274,N_48696,N_48764);
or U49275 (N_49275,N_48987,N_48857);
or U49276 (N_49276,N_48709,N_48875);
and U49277 (N_49277,N_48567,N_48713);
and U49278 (N_49278,N_48502,N_48698);
xor U49279 (N_49279,N_48572,N_48717);
and U49280 (N_49280,N_48744,N_48896);
nor U49281 (N_49281,N_48644,N_48974);
nor U49282 (N_49282,N_48522,N_48944);
nor U49283 (N_49283,N_48758,N_48940);
nand U49284 (N_49284,N_48579,N_48881);
nor U49285 (N_49285,N_48891,N_48548);
xor U49286 (N_49286,N_48600,N_48755);
and U49287 (N_49287,N_48529,N_48987);
nand U49288 (N_49288,N_48657,N_48955);
nor U49289 (N_49289,N_48639,N_48602);
or U49290 (N_49290,N_48716,N_48597);
and U49291 (N_49291,N_48596,N_48658);
nand U49292 (N_49292,N_48594,N_48936);
nor U49293 (N_49293,N_48916,N_48502);
and U49294 (N_49294,N_48522,N_48669);
nor U49295 (N_49295,N_48884,N_48553);
and U49296 (N_49296,N_48838,N_48884);
nor U49297 (N_49297,N_48900,N_48620);
nand U49298 (N_49298,N_48855,N_48779);
or U49299 (N_49299,N_48660,N_48962);
and U49300 (N_49300,N_48697,N_48667);
nand U49301 (N_49301,N_48555,N_48604);
or U49302 (N_49302,N_48716,N_48581);
or U49303 (N_49303,N_48678,N_48542);
nor U49304 (N_49304,N_48734,N_48940);
xnor U49305 (N_49305,N_48660,N_48820);
and U49306 (N_49306,N_48621,N_48847);
nor U49307 (N_49307,N_48677,N_48998);
xor U49308 (N_49308,N_48921,N_48500);
nand U49309 (N_49309,N_48576,N_48777);
nand U49310 (N_49310,N_48909,N_48949);
and U49311 (N_49311,N_48805,N_48731);
and U49312 (N_49312,N_48521,N_48816);
nor U49313 (N_49313,N_48875,N_48640);
or U49314 (N_49314,N_48911,N_48745);
or U49315 (N_49315,N_48656,N_48758);
and U49316 (N_49316,N_48935,N_48712);
nand U49317 (N_49317,N_48651,N_48690);
nand U49318 (N_49318,N_48666,N_48801);
xnor U49319 (N_49319,N_48567,N_48606);
or U49320 (N_49320,N_48973,N_48520);
nand U49321 (N_49321,N_48755,N_48551);
and U49322 (N_49322,N_48501,N_48662);
xnor U49323 (N_49323,N_48807,N_48837);
xor U49324 (N_49324,N_48595,N_48527);
or U49325 (N_49325,N_48696,N_48963);
nor U49326 (N_49326,N_48655,N_48504);
or U49327 (N_49327,N_48813,N_48515);
nand U49328 (N_49328,N_48571,N_48713);
and U49329 (N_49329,N_48593,N_48919);
nand U49330 (N_49330,N_48824,N_48827);
and U49331 (N_49331,N_48611,N_48606);
xor U49332 (N_49332,N_48817,N_48571);
and U49333 (N_49333,N_48881,N_48807);
xnor U49334 (N_49334,N_48845,N_48593);
and U49335 (N_49335,N_48576,N_48845);
and U49336 (N_49336,N_48885,N_48908);
or U49337 (N_49337,N_48558,N_48608);
xnor U49338 (N_49338,N_48781,N_48909);
or U49339 (N_49339,N_48835,N_48600);
nor U49340 (N_49340,N_48929,N_48849);
or U49341 (N_49341,N_48807,N_48922);
xor U49342 (N_49342,N_48588,N_48979);
nand U49343 (N_49343,N_48945,N_48545);
or U49344 (N_49344,N_48569,N_48506);
xor U49345 (N_49345,N_48518,N_48902);
or U49346 (N_49346,N_48670,N_48610);
nand U49347 (N_49347,N_48683,N_48612);
or U49348 (N_49348,N_48953,N_48820);
or U49349 (N_49349,N_48647,N_48746);
xnor U49350 (N_49350,N_48620,N_48774);
xor U49351 (N_49351,N_48698,N_48886);
nand U49352 (N_49352,N_48741,N_48717);
or U49353 (N_49353,N_48948,N_48791);
xor U49354 (N_49354,N_48623,N_48764);
xnor U49355 (N_49355,N_48822,N_48870);
or U49356 (N_49356,N_48916,N_48903);
nor U49357 (N_49357,N_48672,N_48957);
or U49358 (N_49358,N_48871,N_48964);
or U49359 (N_49359,N_48889,N_48706);
and U49360 (N_49360,N_48535,N_48538);
and U49361 (N_49361,N_48710,N_48731);
nand U49362 (N_49362,N_48932,N_48569);
xnor U49363 (N_49363,N_48707,N_48513);
nor U49364 (N_49364,N_48797,N_48932);
and U49365 (N_49365,N_48661,N_48581);
and U49366 (N_49366,N_48833,N_48547);
nand U49367 (N_49367,N_48915,N_48506);
and U49368 (N_49368,N_48846,N_48869);
nor U49369 (N_49369,N_48646,N_48566);
nor U49370 (N_49370,N_48693,N_48887);
xor U49371 (N_49371,N_48507,N_48619);
nand U49372 (N_49372,N_48632,N_48635);
xor U49373 (N_49373,N_48863,N_48907);
nand U49374 (N_49374,N_48537,N_48843);
and U49375 (N_49375,N_48982,N_48877);
or U49376 (N_49376,N_48809,N_48881);
and U49377 (N_49377,N_48957,N_48797);
xnor U49378 (N_49378,N_48515,N_48581);
and U49379 (N_49379,N_48963,N_48521);
nor U49380 (N_49380,N_48703,N_48608);
or U49381 (N_49381,N_48834,N_48996);
or U49382 (N_49382,N_48516,N_48827);
xor U49383 (N_49383,N_48830,N_48976);
xor U49384 (N_49384,N_48952,N_48721);
nand U49385 (N_49385,N_48694,N_48763);
nand U49386 (N_49386,N_48583,N_48775);
nand U49387 (N_49387,N_48743,N_48997);
or U49388 (N_49388,N_48682,N_48551);
or U49389 (N_49389,N_48500,N_48601);
xor U49390 (N_49390,N_48704,N_48702);
or U49391 (N_49391,N_48544,N_48597);
or U49392 (N_49392,N_48710,N_48968);
and U49393 (N_49393,N_48964,N_48525);
nor U49394 (N_49394,N_48993,N_48665);
nand U49395 (N_49395,N_48819,N_48599);
nor U49396 (N_49396,N_48504,N_48580);
nor U49397 (N_49397,N_48643,N_48957);
nor U49398 (N_49398,N_48924,N_48775);
nand U49399 (N_49399,N_48617,N_48817);
nand U49400 (N_49400,N_48532,N_48957);
nand U49401 (N_49401,N_48739,N_48988);
nor U49402 (N_49402,N_48909,N_48740);
and U49403 (N_49403,N_48746,N_48598);
or U49404 (N_49404,N_48553,N_48504);
or U49405 (N_49405,N_48959,N_48847);
nand U49406 (N_49406,N_48822,N_48883);
xor U49407 (N_49407,N_48882,N_48564);
nand U49408 (N_49408,N_48710,N_48638);
nand U49409 (N_49409,N_48744,N_48825);
nor U49410 (N_49410,N_48552,N_48869);
and U49411 (N_49411,N_48589,N_48878);
xnor U49412 (N_49412,N_48860,N_48707);
nand U49413 (N_49413,N_48868,N_48941);
nor U49414 (N_49414,N_48826,N_48900);
and U49415 (N_49415,N_48548,N_48679);
xor U49416 (N_49416,N_48631,N_48967);
and U49417 (N_49417,N_48737,N_48795);
or U49418 (N_49418,N_48961,N_48570);
and U49419 (N_49419,N_48873,N_48702);
and U49420 (N_49420,N_48766,N_48883);
xor U49421 (N_49421,N_48982,N_48858);
and U49422 (N_49422,N_48786,N_48702);
nor U49423 (N_49423,N_48560,N_48546);
xor U49424 (N_49424,N_48580,N_48598);
and U49425 (N_49425,N_48826,N_48680);
or U49426 (N_49426,N_48646,N_48956);
or U49427 (N_49427,N_48884,N_48626);
and U49428 (N_49428,N_48899,N_48998);
and U49429 (N_49429,N_48559,N_48944);
or U49430 (N_49430,N_48702,N_48552);
nand U49431 (N_49431,N_48757,N_48515);
nand U49432 (N_49432,N_48788,N_48647);
and U49433 (N_49433,N_48560,N_48851);
nor U49434 (N_49434,N_48853,N_48600);
or U49435 (N_49435,N_48682,N_48751);
xor U49436 (N_49436,N_48741,N_48926);
xnor U49437 (N_49437,N_48975,N_48900);
or U49438 (N_49438,N_48736,N_48733);
nor U49439 (N_49439,N_48905,N_48700);
or U49440 (N_49440,N_48527,N_48725);
xnor U49441 (N_49441,N_48832,N_48736);
or U49442 (N_49442,N_48896,N_48671);
nand U49443 (N_49443,N_48956,N_48684);
xor U49444 (N_49444,N_48877,N_48855);
nand U49445 (N_49445,N_48933,N_48686);
nand U49446 (N_49446,N_48840,N_48648);
nor U49447 (N_49447,N_48612,N_48928);
nand U49448 (N_49448,N_48915,N_48738);
and U49449 (N_49449,N_48951,N_48669);
and U49450 (N_49450,N_48715,N_48540);
nand U49451 (N_49451,N_48569,N_48764);
nand U49452 (N_49452,N_48974,N_48935);
or U49453 (N_49453,N_48783,N_48565);
xnor U49454 (N_49454,N_48827,N_48896);
or U49455 (N_49455,N_48942,N_48676);
and U49456 (N_49456,N_48839,N_48864);
nor U49457 (N_49457,N_48927,N_48849);
xnor U49458 (N_49458,N_48570,N_48626);
or U49459 (N_49459,N_48755,N_48679);
nand U49460 (N_49460,N_48890,N_48858);
and U49461 (N_49461,N_48655,N_48539);
nand U49462 (N_49462,N_48681,N_48635);
nor U49463 (N_49463,N_48503,N_48599);
and U49464 (N_49464,N_48551,N_48651);
nand U49465 (N_49465,N_48762,N_48602);
nor U49466 (N_49466,N_48953,N_48919);
nand U49467 (N_49467,N_48604,N_48657);
or U49468 (N_49468,N_48943,N_48945);
and U49469 (N_49469,N_48601,N_48760);
or U49470 (N_49470,N_48518,N_48932);
or U49471 (N_49471,N_48557,N_48616);
or U49472 (N_49472,N_48960,N_48837);
nand U49473 (N_49473,N_48852,N_48922);
or U49474 (N_49474,N_48789,N_48559);
nand U49475 (N_49475,N_48565,N_48583);
nor U49476 (N_49476,N_48554,N_48760);
nand U49477 (N_49477,N_48963,N_48687);
and U49478 (N_49478,N_48949,N_48623);
nor U49479 (N_49479,N_48514,N_48790);
or U49480 (N_49480,N_48731,N_48707);
and U49481 (N_49481,N_48879,N_48741);
nor U49482 (N_49482,N_48873,N_48807);
or U49483 (N_49483,N_48937,N_48924);
and U49484 (N_49484,N_48966,N_48621);
or U49485 (N_49485,N_48538,N_48648);
xor U49486 (N_49486,N_48952,N_48787);
xor U49487 (N_49487,N_48769,N_48757);
xor U49488 (N_49488,N_48980,N_48589);
xnor U49489 (N_49489,N_48781,N_48522);
nand U49490 (N_49490,N_48849,N_48512);
xnor U49491 (N_49491,N_48839,N_48878);
nor U49492 (N_49492,N_48749,N_48866);
nor U49493 (N_49493,N_48535,N_48610);
or U49494 (N_49494,N_48610,N_48625);
nand U49495 (N_49495,N_48680,N_48527);
nand U49496 (N_49496,N_48986,N_48661);
or U49497 (N_49497,N_48842,N_48972);
and U49498 (N_49498,N_48898,N_48508);
and U49499 (N_49499,N_48856,N_48750);
xor U49500 (N_49500,N_49244,N_49181);
and U49501 (N_49501,N_49326,N_49229);
nor U49502 (N_49502,N_49389,N_49331);
and U49503 (N_49503,N_49015,N_49104);
xnor U49504 (N_49504,N_49067,N_49363);
or U49505 (N_49505,N_49129,N_49075);
xnor U49506 (N_49506,N_49279,N_49442);
or U49507 (N_49507,N_49484,N_49174);
or U49508 (N_49508,N_49076,N_49246);
nor U49509 (N_49509,N_49108,N_49355);
xnor U49510 (N_49510,N_49032,N_49204);
and U49511 (N_49511,N_49154,N_49328);
and U49512 (N_49512,N_49380,N_49155);
xnor U49513 (N_49513,N_49082,N_49411);
and U49514 (N_49514,N_49377,N_49258);
or U49515 (N_49515,N_49496,N_49308);
or U49516 (N_49516,N_49419,N_49459);
and U49517 (N_49517,N_49054,N_49121);
nand U49518 (N_49518,N_49226,N_49233);
and U49519 (N_49519,N_49271,N_49418);
nor U49520 (N_49520,N_49044,N_49143);
xor U49521 (N_49521,N_49083,N_49309);
nand U49522 (N_49522,N_49238,N_49159);
or U49523 (N_49523,N_49491,N_49109);
nor U49524 (N_49524,N_49281,N_49190);
or U49525 (N_49525,N_49357,N_49046);
nand U49526 (N_49526,N_49250,N_49147);
or U49527 (N_49527,N_49180,N_49035);
or U49528 (N_49528,N_49049,N_49257);
nor U49529 (N_49529,N_49058,N_49414);
and U49530 (N_49530,N_49351,N_49406);
nand U49531 (N_49531,N_49381,N_49292);
or U49532 (N_49532,N_49086,N_49362);
nor U49533 (N_49533,N_49408,N_49077);
xnor U49534 (N_49534,N_49300,N_49350);
xnor U49535 (N_49535,N_49068,N_49495);
and U49536 (N_49536,N_49353,N_49405);
and U49537 (N_49537,N_49303,N_49119);
and U49538 (N_49538,N_49220,N_49367);
xor U49539 (N_49539,N_49236,N_49449);
and U49540 (N_49540,N_49088,N_49285);
and U49541 (N_49541,N_49436,N_49024);
nand U49542 (N_49542,N_49092,N_49070);
nand U49543 (N_49543,N_49313,N_49269);
and U49544 (N_49544,N_49208,N_49451);
nor U49545 (N_49545,N_49304,N_49274);
nand U49546 (N_49546,N_49492,N_49234);
xnor U49547 (N_49547,N_49456,N_49441);
nand U49548 (N_49548,N_49420,N_49342);
xnor U49549 (N_49549,N_49005,N_49305);
xnor U49550 (N_49550,N_49402,N_49057);
xor U49551 (N_49551,N_49487,N_49467);
nand U49552 (N_49552,N_49360,N_49162);
nor U49553 (N_49553,N_49332,N_49125);
or U49554 (N_49554,N_49018,N_49117);
and U49555 (N_49555,N_49315,N_49283);
nand U49556 (N_49556,N_49020,N_49065);
nand U49557 (N_49557,N_49217,N_49282);
xnor U49558 (N_49558,N_49163,N_49011);
or U49559 (N_49559,N_49232,N_49369);
and U49560 (N_49560,N_49319,N_49066);
and U49561 (N_49561,N_49266,N_49063);
nor U49562 (N_49562,N_49434,N_49242);
nand U49563 (N_49563,N_49422,N_49412);
xor U49564 (N_49564,N_49223,N_49019);
or U49565 (N_49565,N_49100,N_49297);
nand U49566 (N_49566,N_49383,N_49392);
or U49567 (N_49567,N_49179,N_49134);
and U49568 (N_49568,N_49106,N_49173);
xnor U49569 (N_49569,N_49316,N_49059);
nand U49570 (N_49570,N_49069,N_49037);
nand U49571 (N_49571,N_49373,N_49477);
and U49572 (N_49572,N_49293,N_49384);
or U49573 (N_49573,N_49382,N_49146);
nor U49574 (N_49574,N_49391,N_49178);
and U49575 (N_49575,N_49317,N_49062);
nand U49576 (N_49576,N_49177,N_49337);
and U49577 (N_49577,N_49352,N_49201);
nor U49578 (N_49578,N_49499,N_49288);
or U49579 (N_49579,N_49335,N_49031);
xor U49580 (N_49580,N_49343,N_49324);
nor U49581 (N_49581,N_49094,N_49004);
or U49582 (N_49582,N_49465,N_49435);
nor U49583 (N_49583,N_49152,N_49008);
nand U49584 (N_49584,N_49284,N_49206);
and U49585 (N_49585,N_49338,N_49395);
nand U49586 (N_49586,N_49424,N_49452);
or U49587 (N_49587,N_49053,N_49023);
or U49588 (N_49588,N_49267,N_49371);
and U49589 (N_49589,N_49454,N_49221);
nor U49590 (N_49590,N_49368,N_49041);
xor U49591 (N_49591,N_49196,N_49349);
and U49592 (N_49592,N_49334,N_49047);
or U49593 (N_49593,N_49014,N_49128);
nand U49594 (N_49594,N_49137,N_49055);
nor U49595 (N_49595,N_49445,N_49141);
or U49596 (N_49596,N_49481,N_49421);
xor U49597 (N_49597,N_49123,N_49160);
xor U49598 (N_49598,N_49097,N_49056);
and U49599 (N_49599,N_49472,N_49039);
nor U49600 (N_49600,N_49458,N_49443);
or U49601 (N_49601,N_49051,N_49156);
xor U49602 (N_49602,N_49401,N_49264);
and U49603 (N_49603,N_49262,N_49361);
nor U49604 (N_49604,N_49192,N_49333);
or U49605 (N_49605,N_49400,N_49322);
and U49606 (N_49606,N_49183,N_49398);
nor U49607 (N_49607,N_49142,N_49112);
nor U49608 (N_49608,N_49022,N_49040);
xor U49609 (N_49609,N_49488,N_49375);
nand U49610 (N_49610,N_49093,N_49139);
xor U49611 (N_49611,N_49095,N_49016);
nand U49612 (N_49612,N_49164,N_49034);
xnor U49613 (N_49613,N_49429,N_49149);
xor U49614 (N_49614,N_49036,N_49078);
xnor U49615 (N_49615,N_49189,N_49348);
xor U49616 (N_49616,N_49222,N_49038);
or U49617 (N_49617,N_49275,N_49224);
nand U49618 (N_49618,N_49476,N_49209);
nor U49619 (N_49619,N_49431,N_49425);
and U49620 (N_49620,N_49253,N_49199);
or U49621 (N_49621,N_49071,N_49494);
nor U49622 (N_49622,N_49111,N_49176);
nand U49623 (N_49623,N_49365,N_49268);
nor U49624 (N_49624,N_49294,N_49493);
xor U49625 (N_49625,N_49193,N_49376);
xnor U49626 (N_49626,N_49072,N_49290);
and U49627 (N_49627,N_49000,N_49336);
nand U49628 (N_49628,N_49430,N_49460);
nand U49629 (N_49629,N_49248,N_49455);
xor U49630 (N_49630,N_49245,N_49158);
nand U49631 (N_49631,N_49140,N_49415);
nor U49632 (N_49632,N_49347,N_49272);
nor U49633 (N_49633,N_49374,N_49026);
xor U49634 (N_49634,N_49330,N_49354);
or U49635 (N_49635,N_49265,N_49052);
xnor U49636 (N_49636,N_49498,N_49261);
nor U49637 (N_49637,N_49416,N_49218);
xor U49638 (N_49638,N_49203,N_49230);
nor U49639 (N_49639,N_49187,N_49085);
xor U49640 (N_49640,N_49237,N_49437);
xor U49641 (N_49641,N_49466,N_49298);
xor U49642 (N_49642,N_49243,N_49027);
and U49643 (N_49643,N_49457,N_49273);
and U49644 (N_49644,N_49145,N_49251);
or U49645 (N_49645,N_49438,N_49200);
nor U49646 (N_49646,N_49359,N_49385);
xor U49647 (N_49647,N_49122,N_49479);
xor U49648 (N_49648,N_49195,N_49132);
or U49649 (N_49649,N_49194,N_49341);
xor U49650 (N_49650,N_49482,N_49329);
nand U49651 (N_49651,N_49219,N_49228);
nor U49652 (N_49652,N_49169,N_49296);
nor U49653 (N_49653,N_49186,N_49386);
or U49654 (N_49654,N_49118,N_49399);
nand U49655 (N_49655,N_49302,N_49320);
and U49656 (N_49656,N_49126,N_49478);
nand U49657 (N_49657,N_49182,N_49247);
nor U49658 (N_49658,N_49388,N_49346);
xnor U49659 (N_49659,N_49061,N_49098);
nand U49660 (N_49660,N_49311,N_49090);
xor U49661 (N_49661,N_49387,N_49471);
or U49662 (N_49662,N_49409,N_49151);
or U49663 (N_49663,N_49105,N_49453);
and U49664 (N_49664,N_49364,N_49136);
nand U49665 (N_49665,N_49073,N_49107);
and U49666 (N_49666,N_49207,N_49447);
nor U49667 (N_49667,N_49252,N_49497);
and U49668 (N_49668,N_49115,N_49113);
nor U49669 (N_49669,N_49396,N_49116);
xnor U49670 (N_49670,N_49161,N_49130);
nand U49671 (N_49671,N_49259,N_49433);
nand U49672 (N_49672,N_49241,N_49295);
xnor U49673 (N_49673,N_49210,N_49301);
nand U49674 (N_49674,N_49184,N_49050);
or U49675 (N_49675,N_49366,N_49148);
or U49676 (N_49676,N_49213,N_49091);
or U49677 (N_49677,N_49468,N_49214);
or U49678 (N_49678,N_49045,N_49426);
and U49679 (N_49679,N_49102,N_49440);
nand U49680 (N_49680,N_49255,N_49114);
nor U49681 (N_49681,N_49165,N_49314);
or U49682 (N_49682,N_49240,N_49256);
nand U49683 (N_49683,N_49432,N_49216);
nand U49684 (N_49684,N_49299,N_49017);
or U49685 (N_49685,N_49356,N_49306);
or U49686 (N_49686,N_49413,N_49171);
xnor U49687 (N_49687,N_49135,N_49007);
xnor U49688 (N_49688,N_49394,N_49474);
and U49689 (N_49689,N_49231,N_49463);
and U49690 (N_49690,N_49080,N_49215);
xor U49691 (N_49691,N_49167,N_49470);
or U49692 (N_49692,N_49340,N_49370);
nand U49693 (N_49693,N_49327,N_49263);
nor U49694 (N_49694,N_49043,N_49225);
nand U49695 (N_49695,N_49025,N_49287);
nor U49696 (N_49696,N_49427,N_49099);
nor U49697 (N_49697,N_49461,N_49450);
and U49698 (N_49698,N_49172,N_49397);
xnor U49699 (N_49699,N_49168,N_49480);
xnor U49700 (N_49700,N_49048,N_49087);
nor U49701 (N_49701,N_49010,N_49021);
xor U49702 (N_49702,N_49033,N_49096);
nand U49703 (N_49703,N_49138,N_49310);
or U49704 (N_49704,N_49428,N_49278);
and U49705 (N_49705,N_49249,N_49339);
or U49706 (N_49706,N_49188,N_49013);
and U49707 (N_49707,N_49103,N_49410);
or U49708 (N_49708,N_49191,N_49133);
xor U49709 (N_49709,N_49289,N_49175);
xor U49710 (N_49710,N_49312,N_49464);
and U49711 (N_49711,N_49344,N_49202);
xor U49712 (N_49712,N_49157,N_49286);
and U49713 (N_49713,N_49089,N_49101);
nand U49714 (N_49714,N_49475,N_49064);
or U49715 (N_49715,N_49473,N_49489);
and U49716 (N_49716,N_49469,N_49003);
and U49717 (N_49717,N_49483,N_49291);
and U49718 (N_49718,N_49404,N_49110);
or U49719 (N_49719,N_49127,N_49235);
nor U49720 (N_49720,N_49197,N_49144);
and U49721 (N_49721,N_49205,N_49486);
xnor U49722 (N_49722,N_49439,N_49153);
and U49723 (N_49723,N_49006,N_49084);
or U49724 (N_49724,N_49323,N_49060);
nand U49725 (N_49725,N_49042,N_49407);
nor U49726 (N_49726,N_49009,N_49170);
nor U49727 (N_49727,N_49227,N_49030);
and U49728 (N_49728,N_49307,N_49260);
nand U49729 (N_49729,N_49325,N_49345);
nand U49730 (N_49730,N_49239,N_49446);
nand U49731 (N_49731,N_49074,N_49211);
xor U49732 (N_49732,N_49212,N_49393);
nand U49733 (N_49733,N_49390,N_49372);
and U49734 (N_49734,N_49131,N_49254);
nor U49735 (N_49735,N_49378,N_49198);
nor U49736 (N_49736,N_49277,N_49081);
xnor U49737 (N_49737,N_49485,N_49028);
nor U49738 (N_49738,N_49166,N_49150);
nand U49739 (N_49739,N_49379,N_49270);
nand U49740 (N_49740,N_49462,N_49120);
and U49741 (N_49741,N_49417,N_49001);
nor U49742 (N_49742,N_49321,N_49448);
or U49743 (N_49743,N_49002,N_49012);
or U49744 (N_49744,N_49276,N_49185);
and U49745 (N_49745,N_49029,N_49403);
and U49746 (N_49746,N_49280,N_49490);
nand U49747 (N_49747,N_49318,N_49124);
xor U49748 (N_49748,N_49444,N_49358);
nor U49749 (N_49749,N_49423,N_49079);
nand U49750 (N_49750,N_49015,N_49392);
xnor U49751 (N_49751,N_49488,N_49395);
nand U49752 (N_49752,N_49116,N_49380);
xor U49753 (N_49753,N_49346,N_49108);
nand U49754 (N_49754,N_49306,N_49362);
nor U49755 (N_49755,N_49256,N_49103);
nand U49756 (N_49756,N_49052,N_49312);
xor U49757 (N_49757,N_49385,N_49054);
or U49758 (N_49758,N_49394,N_49410);
and U49759 (N_49759,N_49280,N_49408);
and U49760 (N_49760,N_49425,N_49050);
and U49761 (N_49761,N_49378,N_49317);
nor U49762 (N_49762,N_49071,N_49276);
xnor U49763 (N_49763,N_49133,N_49252);
nor U49764 (N_49764,N_49326,N_49380);
nor U49765 (N_49765,N_49357,N_49231);
xnor U49766 (N_49766,N_49038,N_49085);
nor U49767 (N_49767,N_49265,N_49235);
nor U49768 (N_49768,N_49444,N_49487);
or U49769 (N_49769,N_49483,N_49109);
nand U49770 (N_49770,N_49269,N_49320);
and U49771 (N_49771,N_49328,N_49127);
or U49772 (N_49772,N_49149,N_49096);
or U49773 (N_49773,N_49364,N_49146);
nand U49774 (N_49774,N_49075,N_49303);
or U49775 (N_49775,N_49331,N_49397);
nand U49776 (N_49776,N_49006,N_49338);
or U49777 (N_49777,N_49327,N_49257);
nand U49778 (N_49778,N_49035,N_49016);
nor U49779 (N_49779,N_49011,N_49112);
and U49780 (N_49780,N_49017,N_49255);
and U49781 (N_49781,N_49254,N_49279);
nor U49782 (N_49782,N_49328,N_49412);
and U49783 (N_49783,N_49432,N_49279);
and U49784 (N_49784,N_49107,N_49437);
xor U49785 (N_49785,N_49116,N_49299);
nand U49786 (N_49786,N_49136,N_49058);
and U49787 (N_49787,N_49416,N_49113);
nor U49788 (N_49788,N_49269,N_49114);
or U49789 (N_49789,N_49060,N_49416);
nand U49790 (N_49790,N_49206,N_49052);
and U49791 (N_49791,N_49082,N_49126);
xor U49792 (N_49792,N_49404,N_49152);
or U49793 (N_49793,N_49469,N_49158);
nor U49794 (N_49794,N_49488,N_49148);
xnor U49795 (N_49795,N_49332,N_49101);
xnor U49796 (N_49796,N_49234,N_49056);
nand U49797 (N_49797,N_49377,N_49160);
and U49798 (N_49798,N_49371,N_49104);
xnor U49799 (N_49799,N_49199,N_49366);
or U49800 (N_49800,N_49128,N_49195);
nor U49801 (N_49801,N_49203,N_49146);
xor U49802 (N_49802,N_49069,N_49401);
or U49803 (N_49803,N_49319,N_49286);
nand U49804 (N_49804,N_49363,N_49018);
xnor U49805 (N_49805,N_49143,N_49005);
or U49806 (N_49806,N_49191,N_49123);
nor U49807 (N_49807,N_49484,N_49182);
and U49808 (N_49808,N_49356,N_49444);
xnor U49809 (N_49809,N_49101,N_49019);
xnor U49810 (N_49810,N_49370,N_49363);
and U49811 (N_49811,N_49336,N_49256);
xor U49812 (N_49812,N_49080,N_49481);
xor U49813 (N_49813,N_49489,N_49163);
nand U49814 (N_49814,N_49241,N_49089);
nand U49815 (N_49815,N_49469,N_49392);
or U49816 (N_49816,N_49103,N_49451);
nand U49817 (N_49817,N_49442,N_49463);
and U49818 (N_49818,N_49301,N_49442);
or U49819 (N_49819,N_49017,N_49455);
xor U49820 (N_49820,N_49257,N_49364);
xnor U49821 (N_49821,N_49037,N_49211);
xor U49822 (N_49822,N_49206,N_49129);
and U49823 (N_49823,N_49214,N_49352);
or U49824 (N_49824,N_49137,N_49207);
or U49825 (N_49825,N_49286,N_49013);
and U49826 (N_49826,N_49118,N_49321);
nand U49827 (N_49827,N_49307,N_49217);
xor U49828 (N_49828,N_49005,N_49264);
nand U49829 (N_49829,N_49116,N_49233);
xnor U49830 (N_49830,N_49177,N_49002);
or U49831 (N_49831,N_49013,N_49369);
or U49832 (N_49832,N_49496,N_49290);
or U49833 (N_49833,N_49324,N_49106);
nand U49834 (N_49834,N_49087,N_49353);
or U49835 (N_49835,N_49077,N_49029);
xor U49836 (N_49836,N_49091,N_49287);
or U49837 (N_49837,N_49131,N_49360);
xor U49838 (N_49838,N_49171,N_49352);
xnor U49839 (N_49839,N_49276,N_49465);
nor U49840 (N_49840,N_49213,N_49175);
nor U49841 (N_49841,N_49469,N_49108);
or U49842 (N_49842,N_49272,N_49047);
xor U49843 (N_49843,N_49405,N_49264);
xor U49844 (N_49844,N_49471,N_49001);
nor U49845 (N_49845,N_49253,N_49186);
and U49846 (N_49846,N_49396,N_49383);
nor U49847 (N_49847,N_49380,N_49374);
or U49848 (N_49848,N_49213,N_49037);
nor U49849 (N_49849,N_49370,N_49499);
nor U49850 (N_49850,N_49120,N_49471);
nand U49851 (N_49851,N_49245,N_49354);
or U49852 (N_49852,N_49092,N_49438);
and U49853 (N_49853,N_49481,N_49173);
and U49854 (N_49854,N_49282,N_49249);
and U49855 (N_49855,N_49286,N_49257);
nand U49856 (N_49856,N_49183,N_49315);
nor U49857 (N_49857,N_49138,N_49233);
nand U49858 (N_49858,N_49321,N_49398);
nand U49859 (N_49859,N_49331,N_49352);
xnor U49860 (N_49860,N_49364,N_49259);
and U49861 (N_49861,N_49244,N_49198);
and U49862 (N_49862,N_49101,N_49129);
and U49863 (N_49863,N_49166,N_49255);
xor U49864 (N_49864,N_49211,N_49179);
nor U49865 (N_49865,N_49056,N_49012);
and U49866 (N_49866,N_49474,N_49297);
xnor U49867 (N_49867,N_49334,N_49199);
and U49868 (N_49868,N_49041,N_49359);
nand U49869 (N_49869,N_49472,N_49431);
or U49870 (N_49870,N_49277,N_49297);
xor U49871 (N_49871,N_49237,N_49019);
xor U49872 (N_49872,N_49137,N_49240);
nand U49873 (N_49873,N_49348,N_49224);
xor U49874 (N_49874,N_49224,N_49234);
nand U49875 (N_49875,N_49401,N_49326);
nand U49876 (N_49876,N_49019,N_49333);
nor U49877 (N_49877,N_49445,N_49316);
and U49878 (N_49878,N_49332,N_49275);
or U49879 (N_49879,N_49331,N_49127);
and U49880 (N_49880,N_49223,N_49329);
or U49881 (N_49881,N_49268,N_49066);
xor U49882 (N_49882,N_49469,N_49006);
nor U49883 (N_49883,N_49049,N_49115);
nand U49884 (N_49884,N_49426,N_49185);
and U49885 (N_49885,N_49263,N_49253);
xor U49886 (N_49886,N_49393,N_49201);
nor U49887 (N_49887,N_49056,N_49104);
nor U49888 (N_49888,N_49383,N_49422);
xor U49889 (N_49889,N_49203,N_49216);
nor U49890 (N_49890,N_49073,N_49379);
xor U49891 (N_49891,N_49247,N_49406);
or U49892 (N_49892,N_49110,N_49137);
xnor U49893 (N_49893,N_49394,N_49347);
xnor U49894 (N_49894,N_49203,N_49244);
nand U49895 (N_49895,N_49189,N_49051);
nor U49896 (N_49896,N_49076,N_49413);
nand U49897 (N_49897,N_49204,N_49368);
or U49898 (N_49898,N_49149,N_49089);
nand U49899 (N_49899,N_49125,N_49221);
and U49900 (N_49900,N_49016,N_49475);
and U49901 (N_49901,N_49458,N_49411);
and U49902 (N_49902,N_49184,N_49007);
and U49903 (N_49903,N_49480,N_49130);
and U49904 (N_49904,N_49471,N_49113);
and U49905 (N_49905,N_49451,N_49452);
and U49906 (N_49906,N_49399,N_49107);
nand U49907 (N_49907,N_49264,N_49364);
or U49908 (N_49908,N_49446,N_49162);
nand U49909 (N_49909,N_49000,N_49094);
or U49910 (N_49910,N_49196,N_49384);
nor U49911 (N_49911,N_49260,N_49358);
nand U49912 (N_49912,N_49218,N_49151);
and U49913 (N_49913,N_49032,N_49037);
or U49914 (N_49914,N_49296,N_49497);
or U49915 (N_49915,N_49387,N_49030);
xnor U49916 (N_49916,N_49472,N_49349);
nand U49917 (N_49917,N_49116,N_49150);
xor U49918 (N_49918,N_49421,N_49006);
or U49919 (N_49919,N_49134,N_49394);
xor U49920 (N_49920,N_49053,N_49093);
and U49921 (N_49921,N_49279,N_49343);
xnor U49922 (N_49922,N_49491,N_49242);
xor U49923 (N_49923,N_49466,N_49173);
nand U49924 (N_49924,N_49021,N_49161);
nand U49925 (N_49925,N_49298,N_49393);
or U49926 (N_49926,N_49246,N_49350);
and U49927 (N_49927,N_49045,N_49105);
xor U49928 (N_49928,N_49267,N_49178);
xnor U49929 (N_49929,N_49047,N_49091);
nor U49930 (N_49930,N_49244,N_49222);
nand U49931 (N_49931,N_49323,N_49486);
nor U49932 (N_49932,N_49474,N_49482);
xnor U49933 (N_49933,N_49105,N_49134);
xnor U49934 (N_49934,N_49147,N_49294);
xor U49935 (N_49935,N_49030,N_49078);
and U49936 (N_49936,N_49268,N_49258);
xnor U49937 (N_49937,N_49012,N_49319);
or U49938 (N_49938,N_49306,N_49151);
or U49939 (N_49939,N_49170,N_49188);
nand U49940 (N_49940,N_49304,N_49176);
nor U49941 (N_49941,N_49053,N_49055);
xnor U49942 (N_49942,N_49466,N_49318);
or U49943 (N_49943,N_49158,N_49155);
xnor U49944 (N_49944,N_49487,N_49222);
nor U49945 (N_49945,N_49442,N_49208);
xor U49946 (N_49946,N_49234,N_49107);
or U49947 (N_49947,N_49210,N_49356);
nand U49948 (N_49948,N_49181,N_49298);
and U49949 (N_49949,N_49135,N_49008);
nand U49950 (N_49950,N_49059,N_49041);
nor U49951 (N_49951,N_49269,N_49193);
xor U49952 (N_49952,N_49186,N_49393);
or U49953 (N_49953,N_49442,N_49381);
nand U49954 (N_49954,N_49338,N_49380);
and U49955 (N_49955,N_49049,N_49019);
nand U49956 (N_49956,N_49251,N_49298);
nand U49957 (N_49957,N_49271,N_49029);
nor U49958 (N_49958,N_49281,N_49146);
or U49959 (N_49959,N_49376,N_49409);
or U49960 (N_49960,N_49429,N_49409);
xnor U49961 (N_49961,N_49458,N_49227);
nand U49962 (N_49962,N_49120,N_49092);
xnor U49963 (N_49963,N_49091,N_49476);
nand U49964 (N_49964,N_49193,N_49325);
xnor U49965 (N_49965,N_49188,N_49447);
xor U49966 (N_49966,N_49082,N_49119);
xnor U49967 (N_49967,N_49036,N_49421);
or U49968 (N_49968,N_49166,N_49276);
and U49969 (N_49969,N_49134,N_49419);
nand U49970 (N_49970,N_49403,N_49070);
and U49971 (N_49971,N_49181,N_49091);
or U49972 (N_49972,N_49249,N_49414);
xnor U49973 (N_49973,N_49432,N_49182);
and U49974 (N_49974,N_49481,N_49468);
and U49975 (N_49975,N_49163,N_49223);
and U49976 (N_49976,N_49244,N_49140);
nand U49977 (N_49977,N_49430,N_49359);
nand U49978 (N_49978,N_49063,N_49150);
or U49979 (N_49979,N_49269,N_49022);
nor U49980 (N_49980,N_49242,N_49475);
nor U49981 (N_49981,N_49437,N_49499);
and U49982 (N_49982,N_49244,N_49074);
and U49983 (N_49983,N_49448,N_49096);
nand U49984 (N_49984,N_49079,N_49209);
or U49985 (N_49985,N_49095,N_49063);
nand U49986 (N_49986,N_49458,N_49116);
xnor U49987 (N_49987,N_49389,N_49398);
nand U49988 (N_49988,N_49120,N_49228);
nand U49989 (N_49989,N_49442,N_49140);
and U49990 (N_49990,N_49277,N_49207);
nor U49991 (N_49991,N_49019,N_49460);
and U49992 (N_49992,N_49090,N_49378);
or U49993 (N_49993,N_49208,N_49399);
nand U49994 (N_49994,N_49444,N_49201);
and U49995 (N_49995,N_49205,N_49127);
xnor U49996 (N_49996,N_49032,N_49091);
or U49997 (N_49997,N_49106,N_49286);
and U49998 (N_49998,N_49440,N_49216);
nand U49999 (N_49999,N_49443,N_49380);
xor UO_0 (O_0,N_49821,N_49755);
nand UO_1 (O_1,N_49757,N_49671);
xnor UO_2 (O_2,N_49882,N_49588);
or UO_3 (O_3,N_49772,N_49928);
nor UO_4 (O_4,N_49577,N_49846);
nand UO_5 (O_5,N_49946,N_49625);
nand UO_6 (O_6,N_49764,N_49869);
nor UO_7 (O_7,N_49579,N_49594);
or UO_8 (O_8,N_49566,N_49921);
xnor UO_9 (O_9,N_49822,N_49975);
xnor UO_10 (O_10,N_49521,N_49780);
and UO_11 (O_11,N_49918,N_49617);
xnor UO_12 (O_12,N_49578,N_49626);
nand UO_13 (O_13,N_49845,N_49902);
or UO_14 (O_14,N_49952,N_49690);
xnor UO_15 (O_15,N_49874,N_49799);
or UO_16 (O_16,N_49761,N_49887);
and UO_17 (O_17,N_49677,N_49587);
and UO_18 (O_18,N_49865,N_49858);
or UO_19 (O_19,N_49993,N_49929);
or UO_20 (O_20,N_49836,N_49752);
and UO_21 (O_21,N_49738,N_49814);
nor UO_22 (O_22,N_49991,N_49525);
and UO_23 (O_23,N_49835,N_49842);
xnor UO_24 (O_24,N_49610,N_49703);
nor UO_25 (O_25,N_49619,N_49965);
xor UO_26 (O_26,N_49976,N_49633);
nand UO_27 (O_27,N_49853,N_49652);
xor UO_28 (O_28,N_49723,N_49642);
nand UO_29 (O_29,N_49564,N_49771);
nand UO_30 (O_30,N_49568,N_49581);
nor UO_31 (O_31,N_49540,N_49701);
nor UO_32 (O_32,N_49923,N_49693);
xnor UO_33 (O_33,N_49951,N_49529);
or UO_34 (O_34,N_49927,N_49616);
nand UO_35 (O_35,N_49732,N_49582);
xnor UO_36 (O_36,N_49979,N_49724);
nand UO_37 (O_37,N_49503,N_49974);
nor UO_38 (O_38,N_49550,N_49562);
or UO_39 (O_39,N_49856,N_49609);
and UO_40 (O_40,N_49675,N_49641);
and UO_41 (O_41,N_49645,N_49828);
nand UO_42 (O_42,N_49913,N_49754);
nor UO_43 (O_43,N_49673,N_49802);
xnor UO_44 (O_44,N_49580,N_49999);
and UO_45 (O_45,N_49637,N_49765);
or UO_46 (O_46,N_49973,N_49680);
and UO_47 (O_47,N_49713,N_49942);
or UO_48 (O_48,N_49934,N_49632);
xnor UO_49 (O_49,N_49994,N_49702);
nor UO_50 (O_50,N_49877,N_49744);
nand UO_51 (O_51,N_49978,N_49995);
or UO_52 (O_52,N_49689,N_49825);
and UO_53 (O_53,N_49571,N_49599);
nor UO_54 (O_54,N_49792,N_49962);
or UO_55 (O_55,N_49733,N_49852);
and UO_56 (O_56,N_49507,N_49788);
xnor UO_57 (O_57,N_49914,N_49696);
or UO_58 (O_58,N_49627,N_49750);
and UO_59 (O_59,N_49572,N_49516);
nor UO_60 (O_60,N_49800,N_49669);
nor UO_61 (O_61,N_49982,N_49924);
or UO_62 (O_62,N_49504,N_49532);
nor UO_63 (O_63,N_49807,N_49762);
nand UO_64 (O_64,N_49546,N_49520);
nand UO_65 (O_65,N_49700,N_49998);
nand UO_66 (O_66,N_49506,N_49980);
xor UO_67 (O_67,N_49688,N_49658);
nor UO_68 (O_68,N_49657,N_49816);
xnor UO_69 (O_69,N_49868,N_49873);
nor UO_70 (O_70,N_49538,N_49718);
nor UO_71 (O_71,N_49785,N_49990);
xnor UO_72 (O_72,N_49889,N_49901);
nand UO_73 (O_73,N_49984,N_49751);
xor UO_74 (O_74,N_49900,N_49871);
xor UO_75 (O_75,N_49639,N_49730);
or UO_76 (O_76,N_49570,N_49518);
nand UO_77 (O_77,N_49593,N_49681);
nor UO_78 (O_78,N_49857,N_49911);
and UO_79 (O_79,N_49715,N_49548);
xnor UO_80 (O_80,N_49968,N_49945);
or UO_81 (O_81,N_49940,N_49985);
or UO_82 (O_82,N_49555,N_49551);
nand UO_83 (O_83,N_49937,N_49653);
nand UO_84 (O_84,N_49692,N_49784);
or UO_85 (O_85,N_49584,N_49654);
and UO_86 (O_86,N_49830,N_49563);
xor UO_87 (O_87,N_49848,N_49763);
and UO_88 (O_88,N_49864,N_49508);
nor UO_89 (O_89,N_49971,N_49554);
or UO_90 (O_90,N_49547,N_49988);
and UO_91 (O_91,N_49794,N_49560);
and UO_92 (O_92,N_49808,N_49840);
xnor UO_93 (O_93,N_49589,N_49963);
nor UO_94 (O_94,N_49997,N_49576);
xor UO_95 (O_95,N_49812,N_49523);
and UO_96 (O_96,N_49892,N_49725);
or UO_97 (O_97,N_49904,N_49638);
or UO_98 (O_98,N_49957,N_49829);
and UO_99 (O_99,N_49810,N_49969);
and UO_100 (O_100,N_49967,N_49741);
nor UO_101 (O_101,N_49586,N_49631);
and UO_102 (O_102,N_49820,N_49896);
or UO_103 (O_103,N_49801,N_49668);
nand UO_104 (O_104,N_49909,N_49815);
or UO_105 (O_105,N_49595,N_49666);
nor UO_106 (O_106,N_49517,N_49682);
xor UO_107 (O_107,N_49781,N_49933);
and UO_108 (O_108,N_49742,N_49833);
nor UO_109 (O_109,N_49708,N_49533);
nand UO_110 (O_110,N_49501,N_49987);
and UO_111 (O_111,N_49583,N_49760);
and UO_112 (O_112,N_49542,N_49620);
and UO_113 (O_113,N_49970,N_49512);
nand UO_114 (O_114,N_49736,N_49664);
and UO_115 (O_115,N_49676,N_49950);
and UO_116 (O_116,N_49734,N_49651);
nand UO_117 (O_117,N_49510,N_49849);
or UO_118 (O_118,N_49818,N_49932);
nor UO_119 (O_119,N_49678,N_49726);
xor UO_120 (O_120,N_49522,N_49606);
or UO_121 (O_121,N_49743,N_49679);
or UO_122 (O_122,N_49832,N_49886);
nand UO_123 (O_123,N_49607,N_49798);
nand UO_124 (O_124,N_49981,N_49956);
and UO_125 (O_125,N_49809,N_49731);
and UO_126 (O_126,N_49854,N_49611);
xnor UO_127 (O_127,N_49655,N_49888);
nand UO_128 (O_128,N_49608,N_49526);
or UO_129 (O_129,N_49819,N_49735);
xnor UO_130 (O_130,N_49793,N_49813);
and UO_131 (O_131,N_49767,N_49649);
or UO_132 (O_132,N_49838,N_49686);
or UO_133 (O_133,N_49894,N_49590);
xor UO_134 (O_134,N_49515,N_49876);
or UO_135 (O_135,N_49753,N_49740);
nand UO_136 (O_136,N_49665,N_49710);
xor UO_137 (O_137,N_49843,N_49683);
or UO_138 (O_138,N_49806,N_49804);
nand UO_139 (O_139,N_49776,N_49936);
nor UO_140 (O_140,N_49646,N_49539);
xnor UO_141 (O_141,N_49907,N_49960);
xor UO_142 (O_142,N_49749,N_49720);
nor UO_143 (O_143,N_49596,N_49916);
xnor UO_144 (O_144,N_49541,N_49603);
nand UO_145 (O_145,N_49556,N_49791);
nand UO_146 (O_146,N_49648,N_49716);
nor UO_147 (O_147,N_49943,N_49880);
or UO_148 (O_148,N_49795,N_49779);
xnor UO_149 (O_149,N_49519,N_49543);
or UO_150 (O_150,N_49899,N_49903);
nand UO_151 (O_151,N_49769,N_49640);
nor UO_152 (O_152,N_49817,N_49629);
and UO_153 (O_153,N_49803,N_49513);
nor UO_154 (O_154,N_49919,N_49890);
nor UO_155 (O_155,N_49850,N_49613);
and UO_156 (O_156,N_49672,N_49643);
xor UO_157 (O_157,N_49747,N_49574);
or UO_158 (O_158,N_49511,N_49774);
nor UO_159 (O_159,N_49746,N_49561);
xor UO_160 (O_160,N_49931,N_49558);
nor UO_161 (O_161,N_49958,N_49691);
nor UO_162 (O_162,N_49824,N_49660);
nand UO_163 (O_163,N_49697,N_49775);
and UO_164 (O_164,N_49647,N_49778);
or UO_165 (O_165,N_49863,N_49662);
and UO_166 (O_166,N_49839,N_49851);
nand UO_167 (O_167,N_49552,N_49897);
xnor UO_168 (O_168,N_49948,N_49860);
and UO_169 (O_169,N_49912,N_49674);
xor UO_170 (O_170,N_49949,N_49955);
nand UO_171 (O_171,N_49601,N_49727);
nor UO_172 (O_172,N_49972,N_49527);
or UO_173 (O_173,N_49910,N_49954);
and UO_174 (O_174,N_49714,N_49841);
nor UO_175 (O_175,N_49536,N_49847);
nand UO_176 (O_176,N_49528,N_49695);
or UO_177 (O_177,N_49908,N_49862);
nor UO_178 (O_178,N_49557,N_49935);
and UO_179 (O_179,N_49861,N_49630);
or UO_180 (O_180,N_49567,N_49789);
nand UO_181 (O_181,N_49719,N_49553);
nand UO_182 (O_182,N_49953,N_49786);
xnor UO_183 (O_183,N_49867,N_49694);
nor UO_184 (O_184,N_49895,N_49624);
xor UO_185 (O_185,N_49986,N_49614);
and UO_186 (O_186,N_49621,N_49706);
nand UO_187 (O_187,N_49922,N_49811);
xnor UO_188 (O_188,N_49721,N_49500);
xnor UO_189 (O_189,N_49906,N_49699);
or UO_190 (O_190,N_49623,N_49707);
xor UO_191 (O_191,N_49944,N_49687);
nand UO_192 (O_192,N_49870,N_49745);
nor UO_193 (O_193,N_49917,N_49711);
nor UO_194 (O_194,N_49941,N_49549);
nand UO_195 (O_195,N_49502,N_49717);
xor UO_196 (O_196,N_49855,N_49644);
and UO_197 (O_197,N_49704,N_49905);
nand UO_198 (O_198,N_49939,N_49989);
nor UO_199 (O_199,N_49650,N_49636);
and UO_200 (O_200,N_49530,N_49826);
or UO_201 (O_201,N_49592,N_49670);
xor UO_202 (O_202,N_49866,N_49667);
xor UO_203 (O_203,N_49783,N_49983);
nand UO_204 (O_204,N_49712,N_49926);
or UO_205 (O_205,N_49545,N_49805);
nor UO_206 (O_206,N_49881,N_49615);
and UO_207 (O_207,N_49597,N_49915);
or UO_208 (O_208,N_49612,N_49823);
nand UO_209 (O_209,N_49634,N_49759);
or UO_210 (O_210,N_49604,N_49898);
xor UO_211 (O_211,N_49748,N_49782);
or UO_212 (O_212,N_49509,N_49827);
and UO_213 (O_213,N_49739,N_49883);
xnor UO_214 (O_214,N_49961,N_49959);
nand UO_215 (O_215,N_49966,N_49756);
and UO_216 (O_216,N_49758,N_49796);
and UO_217 (O_217,N_49729,N_49569);
nand UO_218 (O_218,N_49605,N_49505);
nand UO_219 (O_219,N_49534,N_49770);
and UO_220 (O_220,N_49925,N_49709);
nor UO_221 (O_221,N_49879,N_49628);
xnor UO_222 (O_222,N_49872,N_49728);
nand UO_223 (O_223,N_49661,N_49930);
nand UO_224 (O_224,N_49996,N_49722);
and UO_225 (O_225,N_49875,N_49797);
xor UO_226 (O_226,N_49834,N_49684);
nand UO_227 (O_227,N_49602,N_49585);
nand UO_228 (O_228,N_49544,N_49831);
nand UO_229 (O_229,N_49766,N_49537);
or UO_230 (O_230,N_49656,N_49777);
nor UO_231 (O_231,N_49698,N_49885);
nor UO_232 (O_232,N_49768,N_49565);
nand UO_233 (O_233,N_49837,N_49575);
nor UO_234 (O_234,N_49573,N_49514);
nand UO_235 (O_235,N_49598,N_49737);
and UO_236 (O_236,N_49947,N_49559);
nand UO_237 (O_237,N_49591,N_49635);
xor UO_238 (O_238,N_49938,N_49600);
or UO_239 (O_239,N_49535,N_49878);
or UO_240 (O_240,N_49844,N_49977);
and UO_241 (O_241,N_49773,N_49663);
nand UO_242 (O_242,N_49884,N_49859);
xor UO_243 (O_243,N_49787,N_49992);
nand UO_244 (O_244,N_49524,N_49920);
and UO_245 (O_245,N_49705,N_49618);
xnor UO_246 (O_246,N_49685,N_49531);
nand UO_247 (O_247,N_49893,N_49964);
or UO_248 (O_248,N_49891,N_49790);
nor UO_249 (O_249,N_49659,N_49622);
nand UO_250 (O_250,N_49631,N_49806);
and UO_251 (O_251,N_49754,N_49926);
xnor UO_252 (O_252,N_49890,N_49696);
xnor UO_253 (O_253,N_49844,N_49534);
nand UO_254 (O_254,N_49710,N_49666);
nor UO_255 (O_255,N_49511,N_49797);
xor UO_256 (O_256,N_49519,N_49685);
nor UO_257 (O_257,N_49959,N_49892);
and UO_258 (O_258,N_49666,N_49912);
xor UO_259 (O_259,N_49891,N_49877);
or UO_260 (O_260,N_49679,N_49530);
nand UO_261 (O_261,N_49713,N_49963);
nor UO_262 (O_262,N_49855,N_49663);
or UO_263 (O_263,N_49771,N_49807);
xor UO_264 (O_264,N_49672,N_49533);
nand UO_265 (O_265,N_49865,N_49657);
nand UO_266 (O_266,N_49750,N_49573);
and UO_267 (O_267,N_49819,N_49749);
xnor UO_268 (O_268,N_49869,N_49717);
or UO_269 (O_269,N_49885,N_49646);
or UO_270 (O_270,N_49560,N_49750);
nand UO_271 (O_271,N_49700,N_49847);
xor UO_272 (O_272,N_49960,N_49704);
and UO_273 (O_273,N_49674,N_49611);
nand UO_274 (O_274,N_49652,N_49581);
or UO_275 (O_275,N_49760,N_49779);
nand UO_276 (O_276,N_49662,N_49755);
or UO_277 (O_277,N_49972,N_49505);
and UO_278 (O_278,N_49854,N_49552);
xnor UO_279 (O_279,N_49727,N_49672);
nor UO_280 (O_280,N_49827,N_49616);
nor UO_281 (O_281,N_49622,N_49724);
and UO_282 (O_282,N_49650,N_49546);
xnor UO_283 (O_283,N_49896,N_49795);
nor UO_284 (O_284,N_49824,N_49892);
nor UO_285 (O_285,N_49893,N_49994);
nand UO_286 (O_286,N_49876,N_49685);
or UO_287 (O_287,N_49551,N_49984);
or UO_288 (O_288,N_49948,N_49756);
nor UO_289 (O_289,N_49687,N_49837);
or UO_290 (O_290,N_49596,N_49799);
nor UO_291 (O_291,N_49681,N_49690);
nor UO_292 (O_292,N_49878,N_49815);
nand UO_293 (O_293,N_49640,N_49541);
nand UO_294 (O_294,N_49592,N_49545);
nor UO_295 (O_295,N_49714,N_49679);
or UO_296 (O_296,N_49982,N_49946);
or UO_297 (O_297,N_49899,N_49622);
nor UO_298 (O_298,N_49622,N_49840);
xor UO_299 (O_299,N_49655,N_49618);
xnor UO_300 (O_300,N_49936,N_49504);
or UO_301 (O_301,N_49686,N_49540);
xnor UO_302 (O_302,N_49507,N_49758);
and UO_303 (O_303,N_49932,N_49951);
and UO_304 (O_304,N_49703,N_49542);
and UO_305 (O_305,N_49875,N_49837);
and UO_306 (O_306,N_49836,N_49653);
and UO_307 (O_307,N_49623,N_49592);
and UO_308 (O_308,N_49652,N_49774);
and UO_309 (O_309,N_49747,N_49763);
nand UO_310 (O_310,N_49898,N_49909);
nand UO_311 (O_311,N_49975,N_49978);
nand UO_312 (O_312,N_49599,N_49894);
nand UO_313 (O_313,N_49629,N_49627);
nand UO_314 (O_314,N_49742,N_49616);
xor UO_315 (O_315,N_49882,N_49560);
xnor UO_316 (O_316,N_49544,N_49651);
nand UO_317 (O_317,N_49539,N_49535);
nand UO_318 (O_318,N_49505,N_49854);
or UO_319 (O_319,N_49874,N_49977);
xor UO_320 (O_320,N_49645,N_49846);
or UO_321 (O_321,N_49930,N_49558);
or UO_322 (O_322,N_49632,N_49946);
and UO_323 (O_323,N_49750,N_49587);
and UO_324 (O_324,N_49877,N_49896);
or UO_325 (O_325,N_49714,N_49816);
and UO_326 (O_326,N_49837,N_49711);
nor UO_327 (O_327,N_49963,N_49875);
or UO_328 (O_328,N_49813,N_49703);
or UO_329 (O_329,N_49811,N_49500);
nor UO_330 (O_330,N_49964,N_49710);
and UO_331 (O_331,N_49565,N_49639);
nor UO_332 (O_332,N_49562,N_49648);
or UO_333 (O_333,N_49870,N_49596);
xor UO_334 (O_334,N_49505,N_49838);
nor UO_335 (O_335,N_49500,N_49577);
xor UO_336 (O_336,N_49946,N_49581);
and UO_337 (O_337,N_49697,N_49803);
nand UO_338 (O_338,N_49530,N_49900);
or UO_339 (O_339,N_49796,N_49956);
xor UO_340 (O_340,N_49874,N_49880);
xor UO_341 (O_341,N_49858,N_49860);
xnor UO_342 (O_342,N_49687,N_49865);
nand UO_343 (O_343,N_49631,N_49904);
nand UO_344 (O_344,N_49766,N_49783);
or UO_345 (O_345,N_49680,N_49679);
nor UO_346 (O_346,N_49841,N_49939);
nor UO_347 (O_347,N_49971,N_49734);
and UO_348 (O_348,N_49768,N_49722);
and UO_349 (O_349,N_49549,N_49505);
xnor UO_350 (O_350,N_49520,N_49566);
nand UO_351 (O_351,N_49771,N_49843);
nor UO_352 (O_352,N_49875,N_49784);
and UO_353 (O_353,N_49924,N_49786);
and UO_354 (O_354,N_49856,N_49984);
or UO_355 (O_355,N_49751,N_49900);
nand UO_356 (O_356,N_49762,N_49737);
and UO_357 (O_357,N_49926,N_49910);
nor UO_358 (O_358,N_49545,N_49863);
nor UO_359 (O_359,N_49651,N_49523);
nand UO_360 (O_360,N_49890,N_49594);
or UO_361 (O_361,N_49952,N_49524);
and UO_362 (O_362,N_49760,N_49709);
and UO_363 (O_363,N_49610,N_49689);
xnor UO_364 (O_364,N_49880,N_49715);
nor UO_365 (O_365,N_49619,N_49904);
nor UO_366 (O_366,N_49918,N_49621);
nand UO_367 (O_367,N_49989,N_49675);
and UO_368 (O_368,N_49677,N_49647);
nor UO_369 (O_369,N_49725,N_49995);
nand UO_370 (O_370,N_49926,N_49631);
nor UO_371 (O_371,N_49557,N_49674);
or UO_372 (O_372,N_49695,N_49906);
nor UO_373 (O_373,N_49521,N_49501);
or UO_374 (O_374,N_49761,N_49759);
or UO_375 (O_375,N_49560,N_49600);
or UO_376 (O_376,N_49869,N_49802);
xnor UO_377 (O_377,N_49979,N_49694);
or UO_378 (O_378,N_49557,N_49835);
xor UO_379 (O_379,N_49529,N_49942);
or UO_380 (O_380,N_49763,N_49919);
and UO_381 (O_381,N_49813,N_49634);
or UO_382 (O_382,N_49934,N_49680);
nand UO_383 (O_383,N_49822,N_49930);
or UO_384 (O_384,N_49777,N_49671);
and UO_385 (O_385,N_49759,N_49851);
and UO_386 (O_386,N_49712,N_49958);
or UO_387 (O_387,N_49949,N_49531);
nor UO_388 (O_388,N_49616,N_49990);
nand UO_389 (O_389,N_49575,N_49932);
xnor UO_390 (O_390,N_49592,N_49716);
nor UO_391 (O_391,N_49658,N_49544);
nand UO_392 (O_392,N_49870,N_49716);
nor UO_393 (O_393,N_49595,N_49671);
nor UO_394 (O_394,N_49979,N_49659);
nand UO_395 (O_395,N_49802,N_49751);
nor UO_396 (O_396,N_49798,N_49919);
xor UO_397 (O_397,N_49781,N_49937);
and UO_398 (O_398,N_49877,N_49619);
or UO_399 (O_399,N_49584,N_49516);
or UO_400 (O_400,N_49796,N_49822);
nand UO_401 (O_401,N_49620,N_49619);
nand UO_402 (O_402,N_49790,N_49896);
and UO_403 (O_403,N_49677,N_49722);
nor UO_404 (O_404,N_49877,N_49975);
xor UO_405 (O_405,N_49972,N_49718);
and UO_406 (O_406,N_49815,N_49882);
nand UO_407 (O_407,N_49857,N_49513);
and UO_408 (O_408,N_49757,N_49933);
nor UO_409 (O_409,N_49710,N_49982);
nor UO_410 (O_410,N_49894,N_49737);
or UO_411 (O_411,N_49517,N_49884);
and UO_412 (O_412,N_49820,N_49981);
or UO_413 (O_413,N_49606,N_49656);
nor UO_414 (O_414,N_49700,N_49772);
xnor UO_415 (O_415,N_49519,N_49812);
or UO_416 (O_416,N_49673,N_49895);
and UO_417 (O_417,N_49836,N_49862);
or UO_418 (O_418,N_49572,N_49804);
nor UO_419 (O_419,N_49503,N_49778);
xnor UO_420 (O_420,N_49800,N_49732);
and UO_421 (O_421,N_49931,N_49868);
or UO_422 (O_422,N_49993,N_49779);
nor UO_423 (O_423,N_49576,N_49728);
nand UO_424 (O_424,N_49740,N_49736);
or UO_425 (O_425,N_49736,N_49632);
or UO_426 (O_426,N_49557,N_49654);
xor UO_427 (O_427,N_49740,N_49904);
or UO_428 (O_428,N_49674,N_49576);
or UO_429 (O_429,N_49899,N_49784);
xnor UO_430 (O_430,N_49551,N_49801);
nand UO_431 (O_431,N_49576,N_49699);
nor UO_432 (O_432,N_49638,N_49700);
and UO_433 (O_433,N_49905,N_49883);
or UO_434 (O_434,N_49793,N_49897);
nand UO_435 (O_435,N_49716,N_49541);
or UO_436 (O_436,N_49688,N_49624);
and UO_437 (O_437,N_49532,N_49547);
nand UO_438 (O_438,N_49819,N_49658);
nand UO_439 (O_439,N_49998,N_49596);
nand UO_440 (O_440,N_49896,N_49829);
nor UO_441 (O_441,N_49934,N_49648);
or UO_442 (O_442,N_49956,N_49732);
nand UO_443 (O_443,N_49678,N_49745);
nor UO_444 (O_444,N_49809,N_49810);
and UO_445 (O_445,N_49761,N_49733);
nor UO_446 (O_446,N_49672,N_49531);
or UO_447 (O_447,N_49800,N_49584);
xor UO_448 (O_448,N_49787,N_49939);
or UO_449 (O_449,N_49521,N_49676);
nor UO_450 (O_450,N_49717,N_49849);
xor UO_451 (O_451,N_49737,N_49694);
and UO_452 (O_452,N_49976,N_49517);
xor UO_453 (O_453,N_49928,N_49925);
nor UO_454 (O_454,N_49688,N_49570);
or UO_455 (O_455,N_49845,N_49875);
xor UO_456 (O_456,N_49654,N_49529);
nor UO_457 (O_457,N_49753,N_49803);
nand UO_458 (O_458,N_49923,N_49799);
xnor UO_459 (O_459,N_49971,N_49621);
or UO_460 (O_460,N_49794,N_49814);
xnor UO_461 (O_461,N_49703,N_49906);
or UO_462 (O_462,N_49911,N_49635);
nand UO_463 (O_463,N_49714,N_49818);
nand UO_464 (O_464,N_49686,N_49699);
xnor UO_465 (O_465,N_49724,N_49858);
xnor UO_466 (O_466,N_49836,N_49886);
nand UO_467 (O_467,N_49926,N_49909);
xnor UO_468 (O_468,N_49950,N_49939);
and UO_469 (O_469,N_49627,N_49550);
nor UO_470 (O_470,N_49788,N_49778);
and UO_471 (O_471,N_49692,N_49930);
nand UO_472 (O_472,N_49701,N_49520);
nand UO_473 (O_473,N_49732,N_49729);
nand UO_474 (O_474,N_49747,N_49555);
or UO_475 (O_475,N_49768,N_49670);
xor UO_476 (O_476,N_49755,N_49759);
xor UO_477 (O_477,N_49930,N_49638);
xor UO_478 (O_478,N_49755,N_49505);
nor UO_479 (O_479,N_49786,N_49898);
xnor UO_480 (O_480,N_49845,N_49529);
nor UO_481 (O_481,N_49588,N_49558);
and UO_482 (O_482,N_49542,N_49910);
nor UO_483 (O_483,N_49794,N_49619);
or UO_484 (O_484,N_49670,N_49711);
nand UO_485 (O_485,N_49539,N_49988);
nand UO_486 (O_486,N_49883,N_49644);
nor UO_487 (O_487,N_49644,N_49711);
nand UO_488 (O_488,N_49512,N_49501);
nor UO_489 (O_489,N_49769,N_49720);
nor UO_490 (O_490,N_49705,N_49941);
xnor UO_491 (O_491,N_49873,N_49782);
nor UO_492 (O_492,N_49764,N_49683);
and UO_493 (O_493,N_49812,N_49720);
xnor UO_494 (O_494,N_49694,N_49843);
xor UO_495 (O_495,N_49613,N_49770);
nand UO_496 (O_496,N_49791,N_49840);
and UO_497 (O_497,N_49619,N_49837);
xnor UO_498 (O_498,N_49618,N_49852);
xor UO_499 (O_499,N_49716,N_49777);
and UO_500 (O_500,N_49879,N_49959);
and UO_501 (O_501,N_49736,N_49720);
nor UO_502 (O_502,N_49719,N_49804);
and UO_503 (O_503,N_49627,N_49937);
or UO_504 (O_504,N_49693,N_49655);
nor UO_505 (O_505,N_49622,N_49845);
and UO_506 (O_506,N_49812,N_49808);
xor UO_507 (O_507,N_49892,N_49902);
or UO_508 (O_508,N_49656,N_49513);
or UO_509 (O_509,N_49946,N_49596);
xor UO_510 (O_510,N_49504,N_49728);
xor UO_511 (O_511,N_49734,N_49747);
nor UO_512 (O_512,N_49696,N_49737);
xnor UO_513 (O_513,N_49675,N_49610);
and UO_514 (O_514,N_49681,N_49619);
and UO_515 (O_515,N_49825,N_49939);
and UO_516 (O_516,N_49617,N_49688);
nand UO_517 (O_517,N_49640,N_49602);
nand UO_518 (O_518,N_49992,N_49867);
nand UO_519 (O_519,N_49934,N_49562);
or UO_520 (O_520,N_49893,N_49772);
nor UO_521 (O_521,N_49637,N_49858);
or UO_522 (O_522,N_49988,N_49689);
and UO_523 (O_523,N_49930,N_49958);
nor UO_524 (O_524,N_49747,N_49791);
nor UO_525 (O_525,N_49854,N_49923);
and UO_526 (O_526,N_49834,N_49993);
xor UO_527 (O_527,N_49526,N_49827);
nand UO_528 (O_528,N_49947,N_49765);
and UO_529 (O_529,N_49868,N_49549);
or UO_530 (O_530,N_49716,N_49815);
xor UO_531 (O_531,N_49826,N_49568);
nand UO_532 (O_532,N_49790,N_49976);
xnor UO_533 (O_533,N_49706,N_49522);
xnor UO_534 (O_534,N_49724,N_49618);
and UO_535 (O_535,N_49683,N_49514);
xnor UO_536 (O_536,N_49651,N_49574);
nor UO_537 (O_537,N_49540,N_49590);
nand UO_538 (O_538,N_49557,N_49802);
nand UO_539 (O_539,N_49684,N_49577);
xnor UO_540 (O_540,N_49701,N_49595);
and UO_541 (O_541,N_49971,N_49944);
xor UO_542 (O_542,N_49595,N_49609);
nor UO_543 (O_543,N_49527,N_49927);
xor UO_544 (O_544,N_49943,N_49865);
xor UO_545 (O_545,N_49948,N_49899);
or UO_546 (O_546,N_49559,N_49858);
xnor UO_547 (O_547,N_49890,N_49728);
nor UO_548 (O_548,N_49559,N_49788);
and UO_549 (O_549,N_49802,N_49735);
xor UO_550 (O_550,N_49940,N_49720);
nand UO_551 (O_551,N_49975,N_49634);
and UO_552 (O_552,N_49643,N_49957);
and UO_553 (O_553,N_49661,N_49842);
and UO_554 (O_554,N_49789,N_49647);
xor UO_555 (O_555,N_49901,N_49611);
nand UO_556 (O_556,N_49749,N_49566);
nor UO_557 (O_557,N_49703,N_49547);
nand UO_558 (O_558,N_49667,N_49607);
nand UO_559 (O_559,N_49521,N_49627);
nor UO_560 (O_560,N_49527,N_49876);
or UO_561 (O_561,N_49991,N_49905);
xnor UO_562 (O_562,N_49970,N_49709);
nand UO_563 (O_563,N_49928,N_49950);
nand UO_564 (O_564,N_49571,N_49882);
and UO_565 (O_565,N_49905,N_49559);
xor UO_566 (O_566,N_49638,N_49712);
and UO_567 (O_567,N_49799,N_49681);
or UO_568 (O_568,N_49551,N_49511);
xor UO_569 (O_569,N_49975,N_49539);
xnor UO_570 (O_570,N_49611,N_49761);
or UO_571 (O_571,N_49583,N_49754);
nor UO_572 (O_572,N_49906,N_49874);
nand UO_573 (O_573,N_49673,N_49785);
nand UO_574 (O_574,N_49729,N_49854);
nand UO_575 (O_575,N_49502,N_49591);
xor UO_576 (O_576,N_49554,N_49855);
or UO_577 (O_577,N_49736,N_49731);
or UO_578 (O_578,N_49998,N_49620);
nand UO_579 (O_579,N_49545,N_49922);
nand UO_580 (O_580,N_49939,N_49567);
xor UO_581 (O_581,N_49604,N_49721);
xnor UO_582 (O_582,N_49839,N_49804);
nand UO_583 (O_583,N_49754,N_49875);
and UO_584 (O_584,N_49892,N_49686);
and UO_585 (O_585,N_49911,N_49998);
nor UO_586 (O_586,N_49962,N_49912);
xor UO_587 (O_587,N_49745,N_49505);
xor UO_588 (O_588,N_49700,N_49508);
xor UO_589 (O_589,N_49997,N_49604);
nand UO_590 (O_590,N_49884,N_49946);
or UO_591 (O_591,N_49540,N_49527);
nand UO_592 (O_592,N_49795,N_49902);
nor UO_593 (O_593,N_49836,N_49670);
nor UO_594 (O_594,N_49905,N_49628);
nor UO_595 (O_595,N_49892,N_49562);
or UO_596 (O_596,N_49778,N_49599);
nand UO_597 (O_597,N_49537,N_49945);
nor UO_598 (O_598,N_49810,N_49838);
or UO_599 (O_599,N_49875,N_49840);
or UO_600 (O_600,N_49682,N_49993);
nor UO_601 (O_601,N_49713,N_49980);
xor UO_602 (O_602,N_49852,N_49761);
nor UO_603 (O_603,N_49576,N_49828);
or UO_604 (O_604,N_49907,N_49982);
nand UO_605 (O_605,N_49791,N_49818);
xnor UO_606 (O_606,N_49933,N_49734);
nor UO_607 (O_607,N_49876,N_49863);
nor UO_608 (O_608,N_49549,N_49957);
nand UO_609 (O_609,N_49645,N_49558);
and UO_610 (O_610,N_49637,N_49883);
and UO_611 (O_611,N_49666,N_49648);
nand UO_612 (O_612,N_49612,N_49845);
nand UO_613 (O_613,N_49574,N_49696);
or UO_614 (O_614,N_49737,N_49750);
xnor UO_615 (O_615,N_49715,N_49934);
nor UO_616 (O_616,N_49619,N_49724);
or UO_617 (O_617,N_49827,N_49511);
xnor UO_618 (O_618,N_49985,N_49954);
or UO_619 (O_619,N_49931,N_49799);
xor UO_620 (O_620,N_49635,N_49573);
or UO_621 (O_621,N_49808,N_49674);
or UO_622 (O_622,N_49566,N_49556);
xor UO_623 (O_623,N_49763,N_49672);
nor UO_624 (O_624,N_49727,N_49963);
nor UO_625 (O_625,N_49963,N_49609);
nor UO_626 (O_626,N_49673,N_49638);
or UO_627 (O_627,N_49953,N_49992);
or UO_628 (O_628,N_49899,N_49994);
nand UO_629 (O_629,N_49564,N_49758);
xnor UO_630 (O_630,N_49522,N_49771);
or UO_631 (O_631,N_49787,N_49549);
nor UO_632 (O_632,N_49697,N_49784);
nor UO_633 (O_633,N_49997,N_49904);
xor UO_634 (O_634,N_49729,N_49741);
and UO_635 (O_635,N_49889,N_49878);
nor UO_636 (O_636,N_49579,N_49946);
nor UO_637 (O_637,N_49754,N_49544);
nor UO_638 (O_638,N_49687,N_49987);
nor UO_639 (O_639,N_49541,N_49626);
xor UO_640 (O_640,N_49679,N_49831);
or UO_641 (O_641,N_49768,N_49931);
xnor UO_642 (O_642,N_49666,N_49713);
xnor UO_643 (O_643,N_49530,N_49922);
xor UO_644 (O_644,N_49847,N_49546);
and UO_645 (O_645,N_49966,N_49906);
nor UO_646 (O_646,N_49552,N_49526);
or UO_647 (O_647,N_49814,N_49918);
nand UO_648 (O_648,N_49990,N_49552);
xor UO_649 (O_649,N_49545,N_49762);
nor UO_650 (O_650,N_49697,N_49724);
nor UO_651 (O_651,N_49571,N_49880);
nor UO_652 (O_652,N_49566,N_49644);
xnor UO_653 (O_653,N_49716,N_49649);
and UO_654 (O_654,N_49667,N_49986);
xor UO_655 (O_655,N_49760,N_49946);
or UO_656 (O_656,N_49547,N_49652);
or UO_657 (O_657,N_49941,N_49902);
and UO_658 (O_658,N_49785,N_49502);
nand UO_659 (O_659,N_49561,N_49601);
and UO_660 (O_660,N_49621,N_49546);
or UO_661 (O_661,N_49763,N_49583);
or UO_662 (O_662,N_49500,N_49851);
or UO_663 (O_663,N_49501,N_49725);
nor UO_664 (O_664,N_49548,N_49902);
or UO_665 (O_665,N_49629,N_49757);
nor UO_666 (O_666,N_49922,N_49981);
nand UO_667 (O_667,N_49574,N_49860);
and UO_668 (O_668,N_49958,N_49807);
xnor UO_669 (O_669,N_49817,N_49713);
nor UO_670 (O_670,N_49637,N_49846);
nor UO_671 (O_671,N_49820,N_49503);
and UO_672 (O_672,N_49880,N_49763);
and UO_673 (O_673,N_49908,N_49834);
nor UO_674 (O_674,N_49932,N_49565);
nand UO_675 (O_675,N_49667,N_49942);
nor UO_676 (O_676,N_49811,N_49799);
and UO_677 (O_677,N_49847,N_49826);
and UO_678 (O_678,N_49972,N_49906);
or UO_679 (O_679,N_49779,N_49741);
and UO_680 (O_680,N_49612,N_49514);
nand UO_681 (O_681,N_49741,N_49928);
nor UO_682 (O_682,N_49885,N_49958);
and UO_683 (O_683,N_49581,N_49606);
or UO_684 (O_684,N_49672,N_49897);
nand UO_685 (O_685,N_49819,N_49900);
or UO_686 (O_686,N_49560,N_49736);
xnor UO_687 (O_687,N_49591,N_49694);
nor UO_688 (O_688,N_49866,N_49895);
nor UO_689 (O_689,N_49877,N_49592);
or UO_690 (O_690,N_49988,N_49606);
and UO_691 (O_691,N_49789,N_49806);
nand UO_692 (O_692,N_49763,N_49869);
and UO_693 (O_693,N_49610,N_49803);
nand UO_694 (O_694,N_49698,N_49536);
or UO_695 (O_695,N_49932,N_49745);
nor UO_696 (O_696,N_49912,N_49878);
nor UO_697 (O_697,N_49977,N_49519);
or UO_698 (O_698,N_49623,N_49546);
nand UO_699 (O_699,N_49961,N_49807);
nor UO_700 (O_700,N_49545,N_49965);
and UO_701 (O_701,N_49900,N_49768);
xor UO_702 (O_702,N_49847,N_49686);
and UO_703 (O_703,N_49561,N_49618);
and UO_704 (O_704,N_49896,N_49593);
nor UO_705 (O_705,N_49856,N_49546);
xor UO_706 (O_706,N_49737,N_49968);
nor UO_707 (O_707,N_49624,N_49799);
xor UO_708 (O_708,N_49761,N_49836);
xnor UO_709 (O_709,N_49962,N_49533);
xor UO_710 (O_710,N_49524,N_49747);
nor UO_711 (O_711,N_49794,N_49591);
nand UO_712 (O_712,N_49985,N_49694);
or UO_713 (O_713,N_49507,N_49845);
and UO_714 (O_714,N_49988,N_49950);
nand UO_715 (O_715,N_49743,N_49896);
nand UO_716 (O_716,N_49679,N_49730);
or UO_717 (O_717,N_49746,N_49820);
and UO_718 (O_718,N_49954,N_49536);
nor UO_719 (O_719,N_49685,N_49788);
or UO_720 (O_720,N_49863,N_49619);
nor UO_721 (O_721,N_49945,N_49993);
and UO_722 (O_722,N_49638,N_49539);
and UO_723 (O_723,N_49620,N_49713);
nor UO_724 (O_724,N_49625,N_49955);
nor UO_725 (O_725,N_49656,N_49608);
and UO_726 (O_726,N_49697,N_49512);
nor UO_727 (O_727,N_49661,N_49786);
nand UO_728 (O_728,N_49584,N_49720);
and UO_729 (O_729,N_49988,N_49813);
and UO_730 (O_730,N_49690,N_49557);
and UO_731 (O_731,N_49562,N_49680);
nand UO_732 (O_732,N_49588,N_49932);
nand UO_733 (O_733,N_49663,N_49521);
nand UO_734 (O_734,N_49846,N_49842);
xnor UO_735 (O_735,N_49785,N_49692);
nor UO_736 (O_736,N_49999,N_49889);
nand UO_737 (O_737,N_49696,N_49749);
and UO_738 (O_738,N_49596,N_49923);
xnor UO_739 (O_739,N_49755,N_49687);
nor UO_740 (O_740,N_49653,N_49750);
or UO_741 (O_741,N_49645,N_49691);
and UO_742 (O_742,N_49774,N_49681);
nand UO_743 (O_743,N_49820,N_49851);
or UO_744 (O_744,N_49880,N_49964);
xnor UO_745 (O_745,N_49902,N_49971);
xnor UO_746 (O_746,N_49603,N_49660);
nand UO_747 (O_747,N_49615,N_49895);
nor UO_748 (O_748,N_49747,N_49591);
nand UO_749 (O_749,N_49711,N_49912);
or UO_750 (O_750,N_49586,N_49776);
nor UO_751 (O_751,N_49725,N_49843);
or UO_752 (O_752,N_49672,N_49543);
nor UO_753 (O_753,N_49635,N_49845);
xor UO_754 (O_754,N_49539,N_49734);
and UO_755 (O_755,N_49815,N_49668);
or UO_756 (O_756,N_49973,N_49954);
and UO_757 (O_757,N_49580,N_49956);
xnor UO_758 (O_758,N_49745,N_49950);
xor UO_759 (O_759,N_49544,N_49784);
nor UO_760 (O_760,N_49732,N_49791);
or UO_761 (O_761,N_49683,N_49614);
and UO_762 (O_762,N_49553,N_49604);
xnor UO_763 (O_763,N_49748,N_49753);
nand UO_764 (O_764,N_49688,N_49611);
nand UO_765 (O_765,N_49879,N_49521);
and UO_766 (O_766,N_49509,N_49830);
xnor UO_767 (O_767,N_49837,N_49887);
xor UO_768 (O_768,N_49990,N_49559);
nand UO_769 (O_769,N_49858,N_49527);
and UO_770 (O_770,N_49617,N_49888);
xnor UO_771 (O_771,N_49637,N_49842);
xor UO_772 (O_772,N_49551,N_49754);
xor UO_773 (O_773,N_49916,N_49859);
nand UO_774 (O_774,N_49679,N_49685);
xor UO_775 (O_775,N_49549,N_49978);
nor UO_776 (O_776,N_49672,N_49751);
or UO_777 (O_777,N_49962,N_49507);
and UO_778 (O_778,N_49638,N_49994);
xor UO_779 (O_779,N_49642,N_49949);
nand UO_780 (O_780,N_49817,N_49998);
xor UO_781 (O_781,N_49677,N_49563);
and UO_782 (O_782,N_49500,N_49871);
nor UO_783 (O_783,N_49770,N_49773);
xnor UO_784 (O_784,N_49826,N_49727);
xnor UO_785 (O_785,N_49761,N_49874);
and UO_786 (O_786,N_49767,N_49679);
or UO_787 (O_787,N_49800,N_49796);
nor UO_788 (O_788,N_49694,N_49666);
xor UO_789 (O_789,N_49858,N_49561);
xnor UO_790 (O_790,N_49983,N_49733);
and UO_791 (O_791,N_49924,N_49855);
or UO_792 (O_792,N_49934,N_49902);
nor UO_793 (O_793,N_49889,N_49515);
xor UO_794 (O_794,N_49751,N_49843);
and UO_795 (O_795,N_49947,N_49666);
xor UO_796 (O_796,N_49695,N_49926);
or UO_797 (O_797,N_49590,N_49989);
nand UO_798 (O_798,N_49564,N_49903);
or UO_799 (O_799,N_49866,N_49892);
or UO_800 (O_800,N_49644,N_49715);
nor UO_801 (O_801,N_49661,N_49998);
nor UO_802 (O_802,N_49584,N_49628);
or UO_803 (O_803,N_49552,N_49644);
nand UO_804 (O_804,N_49971,N_49977);
and UO_805 (O_805,N_49810,N_49756);
nand UO_806 (O_806,N_49689,N_49591);
xor UO_807 (O_807,N_49906,N_49738);
and UO_808 (O_808,N_49713,N_49629);
xnor UO_809 (O_809,N_49717,N_49552);
nand UO_810 (O_810,N_49617,N_49894);
and UO_811 (O_811,N_49952,N_49976);
xnor UO_812 (O_812,N_49965,N_49714);
and UO_813 (O_813,N_49696,N_49967);
nor UO_814 (O_814,N_49579,N_49790);
nand UO_815 (O_815,N_49849,N_49603);
nor UO_816 (O_816,N_49808,N_49677);
xnor UO_817 (O_817,N_49973,N_49523);
nor UO_818 (O_818,N_49565,N_49695);
nor UO_819 (O_819,N_49701,N_49582);
or UO_820 (O_820,N_49581,N_49633);
or UO_821 (O_821,N_49637,N_49841);
or UO_822 (O_822,N_49948,N_49629);
xor UO_823 (O_823,N_49534,N_49812);
nand UO_824 (O_824,N_49690,N_49671);
nor UO_825 (O_825,N_49855,N_49994);
nand UO_826 (O_826,N_49943,N_49580);
or UO_827 (O_827,N_49949,N_49950);
nor UO_828 (O_828,N_49522,N_49869);
or UO_829 (O_829,N_49641,N_49797);
or UO_830 (O_830,N_49522,N_49854);
and UO_831 (O_831,N_49626,N_49746);
or UO_832 (O_832,N_49608,N_49793);
xnor UO_833 (O_833,N_49685,N_49677);
nor UO_834 (O_834,N_49997,N_49955);
and UO_835 (O_835,N_49539,N_49502);
nor UO_836 (O_836,N_49987,N_49846);
nand UO_837 (O_837,N_49696,N_49986);
nand UO_838 (O_838,N_49615,N_49830);
nand UO_839 (O_839,N_49962,N_49567);
or UO_840 (O_840,N_49771,N_49762);
or UO_841 (O_841,N_49548,N_49884);
xnor UO_842 (O_842,N_49711,N_49880);
nor UO_843 (O_843,N_49594,N_49742);
nor UO_844 (O_844,N_49781,N_49889);
xnor UO_845 (O_845,N_49670,N_49534);
nand UO_846 (O_846,N_49738,N_49928);
and UO_847 (O_847,N_49710,N_49685);
xnor UO_848 (O_848,N_49630,N_49532);
xnor UO_849 (O_849,N_49756,N_49692);
and UO_850 (O_850,N_49697,N_49943);
xor UO_851 (O_851,N_49922,N_49741);
nor UO_852 (O_852,N_49786,N_49976);
xor UO_853 (O_853,N_49773,N_49629);
nand UO_854 (O_854,N_49791,N_49522);
or UO_855 (O_855,N_49902,N_49998);
or UO_856 (O_856,N_49580,N_49553);
nand UO_857 (O_857,N_49635,N_49558);
nor UO_858 (O_858,N_49655,N_49743);
and UO_859 (O_859,N_49816,N_49771);
or UO_860 (O_860,N_49574,N_49985);
and UO_861 (O_861,N_49607,N_49976);
xnor UO_862 (O_862,N_49559,N_49714);
or UO_863 (O_863,N_49742,N_49505);
nor UO_864 (O_864,N_49887,N_49577);
nor UO_865 (O_865,N_49744,N_49559);
nand UO_866 (O_866,N_49820,N_49675);
nand UO_867 (O_867,N_49822,N_49602);
and UO_868 (O_868,N_49727,N_49628);
and UO_869 (O_869,N_49741,N_49988);
nor UO_870 (O_870,N_49500,N_49541);
nor UO_871 (O_871,N_49579,N_49533);
nand UO_872 (O_872,N_49865,N_49985);
and UO_873 (O_873,N_49967,N_49657);
nor UO_874 (O_874,N_49833,N_49713);
and UO_875 (O_875,N_49867,N_49708);
nor UO_876 (O_876,N_49779,N_49945);
xor UO_877 (O_877,N_49683,N_49845);
or UO_878 (O_878,N_49663,N_49726);
and UO_879 (O_879,N_49694,N_49972);
nand UO_880 (O_880,N_49888,N_49507);
and UO_881 (O_881,N_49545,N_49875);
nand UO_882 (O_882,N_49859,N_49541);
xnor UO_883 (O_883,N_49828,N_49591);
nor UO_884 (O_884,N_49673,N_49565);
nor UO_885 (O_885,N_49941,N_49630);
xor UO_886 (O_886,N_49748,N_49565);
and UO_887 (O_887,N_49936,N_49915);
nand UO_888 (O_888,N_49773,N_49761);
and UO_889 (O_889,N_49910,N_49747);
xor UO_890 (O_890,N_49511,N_49739);
nor UO_891 (O_891,N_49647,N_49566);
xor UO_892 (O_892,N_49666,N_49696);
or UO_893 (O_893,N_49611,N_49509);
nor UO_894 (O_894,N_49606,N_49952);
nand UO_895 (O_895,N_49801,N_49830);
nor UO_896 (O_896,N_49564,N_49673);
or UO_897 (O_897,N_49645,N_49885);
nor UO_898 (O_898,N_49925,N_49962);
nand UO_899 (O_899,N_49724,N_49664);
and UO_900 (O_900,N_49750,N_49837);
nor UO_901 (O_901,N_49653,N_49823);
or UO_902 (O_902,N_49706,N_49500);
nor UO_903 (O_903,N_49872,N_49787);
and UO_904 (O_904,N_49625,N_49593);
or UO_905 (O_905,N_49867,N_49741);
or UO_906 (O_906,N_49914,N_49900);
nor UO_907 (O_907,N_49748,N_49879);
xor UO_908 (O_908,N_49958,N_49995);
nor UO_909 (O_909,N_49854,N_49827);
and UO_910 (O_910,N_49994,N_49622);
xnor UO_911 (O_911,N_49606,N_49883);
or UO_912 (O_912,N_49716,N_49657);
nand UO_913 (O_913,N_49751,N_49711);
xor UO_914 (O_914,N_49937,N_49994);
or UO_915 (O_915,N_49763,N_49841);
nor UO_916 (O_916,N_49694,N_49659);
xnor UO_917 (O_917,N_49656,N_49813);
nor UO_918 (O_918,N_49844,N_49838);
or UO_919 (O_919,N_49889,N_49737);
and UO_920 (O_920,N_49524,N_49976);
or UO_921 (O_921,N_49927,N_49754);
nor UO_922 (O_922,N_49611,N_49769);
nor UO_923 (O_923,N_49969,N_49842);
and UO_924 (O_924,N_49769,N_49505);
nor UO_925 (O_925,N_49719,N_49958);
or UO_926 (O_926,N_49892,N_49777);
nand UO_927 (O_927,N_49829,N_49836);
nand UO_928 (O_928,N_49892,N_49581);
nor UO_929 (O_929,N_49504,N_49911);
xnor UO_930 (O_930,N_49673,N_49629);
nor UO_931 (O_931,N_49627,N_49900);
xor UO_932 (O_932,N_49624,N_49574);
nor UO_933 (O_933,N_49507,N_49571);
or UO_934 (O_934,N_49876,N_49833);
nor UO_935 (O_935,N_49867,N_49995);
or UO_936 (O_936,N_49876,N_49956);
nand UO_937 (O_937,N_49812,N_49958);
xor UO_938 (O_938,N_49756,N_49657);
nand UO_939 (O_939,N_49719,N_49592);
or UO_940 (O_940,N_49844,N_49782);
and UO_941 (O_941,N_49633,N_49876);
nor UO_942 (O_942,N_49632,N_49811);
xor UO_943 (O_943,N_49811,N_49906);
and UO_944 (O_944,N_49930,N_49698);
nor UO_945 (O_945,N_49678,N_49683);
nor UO_946 (O_946,N_49892,N_49780);
nor UO_947 (O_947,N_49944,N_49710);
xor UO_948 (O_948,N_49822,N_49949);
nor UO_949 (O_949,N_49933,N_49565);
nor UO_950 (O_950,N_49988,N_49514);
xor UO_951 (O_951,N_49905,N_49963);
or UO_952 (O_952,N_49566,N_49684);
nor UO_953 (O_953,N_49785,N_49594);
and UO_954 (O_954,N_49846,N_49761);
and UO_955 (O_955,N_49943,N_49924);
or UO_956 (O_956,N_49969,N_49586);
nand UO_957 (O_957,N_49872,N_49717);
or UO_958 (O_958,N_49753,N_49780);
nor UO_959 (O_959,N_49670,N_49785);
or UO_960 (O_960,N_49525,N_49806);
or UO_961 (O_961,N_49761,N_49620);
nor UO_962 (O_962,N_49705,N_49697);
or UO_963 (O_963,N_49784,N_49904);
and UO_964 (O_964,N_49933,N_49917);
xnor UO_965 (O_965,N_49716,N_49503);
nand UO_966 (O_966,N_49504,N_49765);
nand UO_967 (O_967,N_49728,N_49572);
and UO_968 (O_968,N_49591,N_49549);
nand UO_969 (O_969,N_49646,N_49867);
and UO_970 (O_970,N_49937,N_49943);
xor UO_971 (O_971,N_49989,N_49920);
nand UO_972 (O_972,N_49790,N_49748);
xnor UO_973 (O_973,N_49974,N_49577);
or UO_974 (O_974,N_49613,N_49942);
or UO_975 (O_975,N_49524,N_49713);
and UO_976 (O_976,N_49667,N_49872);
and UO_977 (O_977,N_49991,N_49943);
or UO_978 (O_978,N_49877,N_49787);
and UO_979 (O_979,N_49593,N_49501);
nor UO_980 (O_980,N_49607,N_49726);
xnor UO_981 (O_981,N_49789,N_49926);
or UO_982 (O_982,N_49919,N_49996);
nand UO_983 (O_983,N_49669,N_49580);
or UO_984 (O_984,N_49852,N_49776);
nor UO_985 (O_985,N_49892,N_49971);
xor UO_986 (O_986,N_49731,N_49840);
xor UO_987 (O_987,N_49506,N_49655);
nand UO_988 (O_988,N_49853,N_49844);
nor UO_989 (O_989,N_49786,N_49821);
or UO_990 (O_990,N_49664,N_49892);
xor UO_991 (O_991,N_49531,N_49588);
xnor UO_992 (O_992,N_49927,N_49693);
or UO_993 (O_993,N_49869,N_49513);
xor UO_994 (O_994,N_49743,N_49566);
or UO_995 (O_995,N_49864,N_49801);
or UO_996 (O_996,N_49752,N_49772);
or UO_997 (O_997,N_49582,N_49913);
and UO_998 (O_998,N_49624,N_49611);
nand UO_999 (O_999,N_49708,N_49615);
xor UO_1000 (O_1000,N_49911,N_49546);
xor UO_1001 (O_1001,N_49991,N_49716);
and UO_1002 (O_1002,N_49597,N_49998);
or UO_1003 (O_1003,N_49507,N_49863);
nor UO_1004 (O_1004,N_49536,N_49923);
xor UO_1005 (O_1005,N_49612,N_49588);
nand UO_1006 (O_1006,N_49743,N_49945);
nand UO_1007 (O_1007,N_49672,N_49656);
nand UO_1008 (O_1008,N_49707,N_49579);
or UO_1009 (O_1009,N_49635,N_49535);
or UO_1010 (O_1010,N_49863,N_49804);
or UO_1011 (O_1011,N_49598,N_49950);
or UO_1012 (O_1012,N_49609,N_49551);
nand UO_1013 (O_1013,N_49505,N_49945);
and UO_1014 (O_1014,N_49956,N_49615);
or UO_1015 (O_1015,N_49633,N_49833);
xor UO_1016 (O_1016,N_49806,N_49915);
or UO_1017 (O_1017,N_49620,N_49588);
nand UO_1018 (O_1018,N_49593,N_49688);
and UO_1019 (O_1019,N_49920,N_49893);
nor UO_1020 (O_1020,N_49819,N_49976);
nor UO_1021 (O_1021,N_49766,N_49565);
nor UO_1022 (O_1022,N_49979,N_49922);
or UO_1023 (O_1023,N_49954,N_49779);
nor UO_1024 (O_1024,N_49615,N_49620);
xnor UO_1025 (O_1025,N_49612,N_49582);
or UO_1026 (O_1026,N_49830,N_49657);
and UO_1027 (O_1027,N_49950,N_49884);
nand UO_1028 (O_1028,N_49909,N_49605);
and UO_1029 (O_1029,N_49813,N_49849);
or UO_1030 (O_1030,N_49962,N_49591);
xnor UO_1031 (O_1031,N_49806,N_49646);
nor UO_1032 (O_1032,N_49878,N_49938);
xnor UO_1033 (O_1033,N_49966,N_49972);
nand UO_1034 (O_1034,N_49500,N_49654);
or UO_1035 (O_1035,N_49851,N_49895);
nor UO_1036 (O_1036,N_49891,N_49539);
xnor UO_1037 (O_1037,N_49623,N_49910);
or UO_1038 (O_1038,N_49502,N_49880);
nand UO_1039 (O_1039,N_49700,N_49774);
nand UO_1040 (O_1040,N_49761,N_49989);
and UO_1041 (O_1041,N_49653,N_49859);
and UO_1042 (O_1042,N_49730,N_49594);
or UO_1043 (O_1043,N_49897,N_49977);
nand UO_1044 (O_1044,N_49568,N_49979);
nand UO_1045 (O_1045,N_49791,N_49994);
or UO_1046 (O_1046,N_49533,N_49577);
or UO_1047 (O_1047,N_49873,N_49721);
xnor UO_1048 (O_1048,N_49915,N_49687);
and UO_1049 (O_1049,N_49719,N_49555);
or UO_1050 (O_1050,N_49853,N_49669);
and UO_1051 (O_1051,N_49914,N_49831);
or UO_1052 (O_1052,N_49793,N_49931);
or UO_1053 (O_1053,N_49864,N_49564);
nor UO_1054 (O_1054,N_49732,N_49560);
nor UO_1055 (O_1055,N_49500,N_49810);
and UO_1056 (O_1056,N_49947,N_49841);
and UO_1057 (O_1057,N_49578,N_49852);
xnor UO_1058 (O_1058,N_49736,N_49951);
nor UO_1059 (O_1059,N_49654,N_49790);
xor UO_1060 (O_1060,N_49722,N_49766);
or UO_1061 (O_1061,N_49982,N_49739);
xor UO_1062 (O_1062,N_49912,N_49722);
nor UO_1063 (O_1063,N_49957,N_49991);
or UO_1064 (O_1064,N_49557,N_49957);
and UO_1065 (O_1065,N_49710,N_49864);
nor UO_1066 (O_1066,N_49989,N_49968);
nand UO_1067 (O_1067,N_49669,N_49672);
nor UO_1068 (O_1068,N_49951,N_49731);
nand UO_1069 (O_1069,N_49550,N_49848);
or UO_1070 (O_1070,N_49762,N_49996);
and UO_1071 (O_1071,N_49705,N_49987);
nand UO_1072 (O_1072,N_49598,N_49995);
and UO_1073 (O_1073,N_49759,N_49820);
nor UO_1074 (O_1074,N_49618,N_49574);
nand UO_1075 (O_1075,N_49550,N_49612);
or UO_1076 (O_1076,N_49523,N_49924);
nor UO_1077 (O_1077,N_49613,N_49779);
or UO_1078 (O_1078,N_49876,N_49744);
nand UO_1079 (O_1079,N_49505,N_49861);
nor UO_1080 (O_1080,N_49661,N_49708);
xor UO_1081 (O_1081,N_49543,N_49958);
nand UO_1082 (O_1082,N_49639,N_49517);
or UO_1083 (O_1083,N_49771,N_49732);
and UO_1084 (O_1084,N_49671,N_49666);
and UO_1085 (O_1085,N_49508,N_49942);
nand UO_1086 (O_1086,N_49829,N_49861);
nor UO_1087 (O_1087,N_49595,N_49685);
and UO_1088 (O_1088,N_49734,N_49958);
or UO_1089 (O_1089,N_49564,N_49515);
nor UO_1090 (O_1090,N_49961,N_49575);
and UO_1091 (O_1091,N_49827,N_49661);
nor UO_1092 (O_1092,N_49582,N_49903);
nand UO_1093 (O_1093,N_49903,N_49911);
and UO_1094 (O_1094,N_49793,N_49540);
nand UO_1095 (O_1095,N_49564,N_49995);
xor UO_1096 (O_1096,N_49907,N_49636);
nor UO_1097 (O_1097,N_49545,N_49851);
nor UO_1098 (O_1098,N_49797,N_49820);
or UO_1099 (O_1099,N_49677,N_49813);
or UO_1100 (O_1100,N_49683,N_49892);
nor UO_1101 (O_1101,N_49872,N_49641);
xnor UO_1102 (O_1102,N_49856,N_49804);
nand UO_1103 (O_1103,N_49881,N_49679);
xnor UO_1104 (O_1104,N_49596,N_49949);
and UO_1105 (O_1105,N_49602,N_49590);
nor UO_1106 (O_1106,N_49535,N_49972);
xnor UO_1107 (O_1107,N_49763,N_49549);
nand UO_1108 (O_1108,N_49598,N_49687);
xnor UO_1109 (O_1109,N_49624,N_49966);
xnor UO_1110 (O_1110,N_49829,N_49999);
nor UO_1111 (O_1111,N_49833,N_49722);
and UO_1112 (O_1112,N_49674,N_49692);
nand UO_1113 (O_1113,N_49560,N_49694);
nor UO_1114 (O_1114,N_49585,N_49532);
and UO_1115 (O_1115,N_49631,N_49895);
xor UO_1116 (O_1116,N_49574,N_49541);
or UO_1117 (O_1117,N_49809,N_49608);
nor UO_1118 (O_1118,N_49638,N_49583);
and UO_1119 (O_1119,N_49709,N_49790);
or UO_1120 (O_1120,N_49950,N_49532);
xnor UO_1121 (O_1121,N_49719,N_49544);
nand UO_1122 (O_1122,N_49683,N_49739);
nor UO_1123 (O_1123,N_49632,N_49702);
and UO_1124 (O_1124,N_49911,N_49551);
xnor UO_1125 (O_1125,N_49792,N_49838);
nand UO_1126 (O_1126,N_49974,N_49705);
nand UO_1127 (O_1127,N_49744,N_49662);
or UO_1128 (O_1128,N_49802,N_49501);
nand UO_1129 (O_1129,N_49550,N_49515);
xor UO_1130 (O_1130,N_49696,N_49709);
and UO_1131 (O_1131,N_49840,N_49513);
or UO_1132 (O_1132,N_49742,N_49961);
or UO_1133 (O_1133,N_49571,N_49988);
nand UO_1134 (O_1134,N_49973,N_49883);
nor UO_1135 (O_1135,N_49637,N_49517);
and UO_1136 (O_1136,N_49825,N_49700);
xnor UO_1137 (O_1137,N_49724,N_49778);
nor UO_1138 (O_1138,N_49652,N_49583);
or UO_1139 (O_1139,N_49724,N_49937);
and UO_1140 (O_1140,N_49760,N_49949);
and UO_1141 (O_1141,N_49597,N_49755);
or UO_1142 (O_1142,N_49687,N_49940);
and UO_1143 (O_1143,N_49756,N_49666);
nor UO_1144 (O_1144,N_49825,N_49978);
nand UO_1145 (O_1145,N_49959,N_49552);
xnor UO_1146 (O_1146,N_49702,N_49552);
and UO_1147 (O_1147,N_49731,N_49685);
and UO_1148 (O_1148,N_49522,N_49839);
and UO_1149 (O_1149,N_49981,N_49686);
nor UO_1150 (O_1150,N_49772,N_49519);
xnor UO_1151 (O_1151,N_49605,N_49827);
nor UO_1152 (O_1152,N_49868,N_49552);
or UO_1153 (O_1153,N_49503,N_49840);
xnor UO_1154 (O_1154,N_49559,N_49635);
or UO_1155 (O_1155,N_49770,N_49664);
and UO_1156 (O_1156,N_49544,N_49897);
nor UO_1157 (O_1157,N_49514,N_49629);
nand UO_1158 (O_1158,N_49799,N_49643);
nand UO_1159 (O_1159,N_49690,N_49960);
and UO_1160 (O_1160,N_49783,N_49811);
xnor UO_1161 (O_1161,N_49853,N_49978);
or UO_1162 (O_1162,N_49766,N_49734);
or UO_1163 (O_1163,N_49711,N_49834);
or UO_1164 (O_1164,N_49964,N_49624);
xor UO_1165 (O_1165,N_49907,N_49775);
nor UO_1166 (O_1166,N_49791,N_49937);
nor UO_1167 (O_1167,N_49708,N_49740);
nor UO_1168 (O_1168,N_49500,N_49597);
nor UO_1169 (O_1169,N_49612,N_49580);
or UO_1170 (O_1170,N_49848,N_49858);
xnor UO_1171 (O_1171,N_49659,N_49883);
nor UO_1172 (O_1172,N_49710,N_49844);
and UO_1173 (O_1173,N_49645,N_49721);
xor UO_1174 (O_1174,N_49689,N_49556);
or UO_1175 (O_1175,N_49992,N_49628);
xor UO_1176 (O_1176,N_49644,N_49546);
and UO_1177 (O_1177,N_49781,N_49645);
xor UO_1178 (O_1178,N_49928,N_49978);
or UO_1179 (O_1179,N_49979,N_49650);
nor UO_1180 (O_1180,N_49585,N_49561);
nor UO_1181 (O_1181,N_49539,N_49746);
nor UO_1182 (O_1182,N_49636,N_49753);
nand UO_1183 (O_1183,N_49795,N_49614);
nor UO_1184 (O_1184,N_49946,N_49931);
xor UO_1185 (O_1185,N_49710,N_49646);
and UO_1186 (O_1186,N_49893,N_49624);
xnor UO_1187 (O_1187,N_49802,N_49707);
nor UO_1188 (O_1188,N_49934,N_49591);
nor UO_1189 (O_1189,N_49810,N_49798);
nand UO_1190 (O_1190,N_49961,N_49605);
and UO_1191 (O_1191,N_49852,N_49754);
or UO_1192 (O_1192,N_49695,N_49515);
and UO_1193 (O_1193,N_49976,N_49619);
xnor UO_1194 (O_1194,N_49554,N_49591);
or UO_1195 (O_1195,N_49818,N_49757);
xnor UO_1196 (O_1196,N_49800,N_49739);
nand UO_1197 (O_1197,N_49685,N_49525);
nor UO_1198 (O_1198,N_49641,N_49552);
nor UO_1199 (O_1199,N_49696,N_49730);
or UO_1200 (O_1200,N_49782,N_49764);
nand UO_1201 (O_1201,N_49870,N_49529);
nor UO_1202 (O_1202,N_49756,N_49639);
nor UO_1203 (O_1203,N_49947,N_49871);
xnor UO_1204 (O_1204,N_49890,N_49694);
and UO_1205 (O_1205,N_49682,N_49535);
and UO_1206 (O_1206,N_49978,N_49933);
or UO_1207 (O_1207,N_49512,N_49725);
nor UO_1208 (O_1208,N_49812,N_49554);
or UO_1209 (O_1209,N_49788,N_49718);
and UO_1210 (O_1210,N_49930,N_49739);
nor UO_1211 (O_1211,N_49733,N_49548);
nand UO_1212 (O_1212,N_49599,N_49943);
xor UO_1213 (O_1213,N_49910,N_49953);
and UO_1214 (O_1214,N_49606,N_49686);
nand UO_1215 (O_1215,N_49980,N_49565);
or UO_1216 (O_1216,N_49705,N_49845);
nand UO_1217 (O_1217,N_49564,N_49710);
xor UO_1218 (O_1218,N_49755,N_49560);
and UO_1219 (O_1219,N_49945,N_49835);
nand UO_1220 (O_1220,N_49975,N_49675);
nand UO_1221 (O_1221,N_49561,N_49656);
nand UO_1222 (O_1222,N_49885,N_49844);
nand UO_1223 (O_1223,N_49678,N_49659);
or UO_1224 (O_1224,N_49790,N_49728);
nand UO_1225 (O_1225,N_49567,N_49751);
or UO_1226 (O_1226,N_49885,N_49705);
xnor UO_1227 (O_1227,N_49992,N_49766);
or UO_1228 (O_1228,N_49850,N_49829);
nand UO_1229 (O_1229,N_49991,N_49723);
nand UO_1230 (O_1230,N_49959,N_49797);
or UO_1231 (O_1231,N_49729,N_49788);
or UO_1232 (O_1232,N_49622,N_49876);
nand UO_1233 (O_1233,N_49876,N_49931);
xnor UO_1234 (O_1234,N_49533,N_49916);
xnor UO_1235 (O_1235,N_49850,N_49956);
or UO_1236 (O_1236,N_49967,N_49641);
xnor UO_1237 (O_1237,N_49879,N_49834);
nand UO_1238 (O_1238,N_49748,N_49966);
or UO_1239 (O_1239,N_49710,N_49975);
and UO_1240 (O_1240,N_49627,N_49648);
nor UO_1241 (O_1241,N_49962,N_49870);
xnor UO_1242 (O_1242,N_49819,N_49990);
and UO_1243 (O_1243,N_49808,N_49657);
or UO_1244 (O_1244,N_49554,N_49623);
nor UO_1245 (O_1245,N_49527,N_49505);
nand UO_1246 (O_1246,N_49969,N_49640);
and UO_1247 (O_1247,N_49508,N_49528);
and UO_1248 (O_1248,N_49963,N_49565);
or UO_1249 (O_1249,N_49895,N_49874);
and UO_1250 (O_1250,N_49773,N_49946);
and UO_1251 (O_1251,N_49987,N_49616);
xor UO_1252 (O_1252,N_49528,N_49713);
nor UO_1253 (O_1253,N_49671,N_49500);
nor UO_1254 (O_1254,N_49636,N_49641);
xnor UO_1255 (O_1255,N_49911,N_49818);
or UO_1256 (O_1256,N_49618,N_49713);
or UO_1257 (O_1257,N_49821,N_49623);
nand UO_1258 (O_1258,N_49526,N_49775);
and UO_1259 (O_1259,N_49716,N_49517);
nand UO_1260 (O_1260,N_49644,N_49588);
nand UO_1261 (O_1261,N_49549,N_49656);
or UO_1262 (O_1262,N_49561,N_49902);
or UO_1263 (O_1263,N_49586,N_49710);
nor UO_1264 (O_1264,N_49695,N_49809);
nor UO_1265 (O_1265,N_49998,N_49899);
and UO_1266 (O_1266,N_49949,N_49819);
or UO_1267 (O_1267,N_49753,N_49551);
nor UO_1268 (O_1268,N_49737,N_49848);
nand UO_1269 (O_1269,N_49503,N_49668);
and UO_1270 (O_1270,N_49707,N_49677);
nand UO_1271 (O_1271,N_49537,N_49540);
and UO_1272 (O_1272,N_49676,N_49616);
and UO_1273 (O_1273,N_49882,N_49904);
and UO_1274 (O_1274,N_49693,N_49867);
or UO_1275 (O_1275,N_49848,N_49507);
nand UO_1276 (O_1276,N_49825,N_49752);
and UO_1277 (O_1277,N_49895,N_49754);
and UO_1278 (O_1278,N_49752,N_49957);
xor UO_1279 (O_1279,N_49906,N_49870);
nand UO_1280 (O_1280,N_49848,N_49600);
and UO_1281 (O_1281,N_49726,N_49888);
xor UO_1282 (O_1282,N_49661,N_49992);
nor UO_1283 (O_1283,N_49570,N_49900);
xnor UO_1284 (O_1284,N_49659,N_49662);
or UO_1285 (O_1285,N_49574,N_49526);
or UO_1286 (O_1286,N_49990,N_49613);
or UO_1287 (O_1287,N_49629,N_49722);
and UO_1288 (O_1288,N_49924,N_49543);
or UO_1289 (O_1289,N_49553,N_49642);
nor UO_1290 (O_1290,N_49805,N_49705);
nand UO_1291 (O_1291,N_49505,N_49954);
xor UO_1292 (O_1292,N_49517,N_49654);
and UO_1293 (O_1293,N_49524,N_49784);
nor UO_1294 (O_1294,N_49565,N_49515);
xor UO_1295 (O_1295,N_49706,N_49506);
or UO_1296 (O_1296,N_49547,N_49969);
and UO_1297 (O_1297,N_49692,N_49665);
or UO_1298 (O_1298,N_49820,N_49899);
nor UO_1299 (O_1299,N_49995,N_49699);
and UO_1300 (O_1300,N_49516,N_49701);
and UO_1301 (O_1301,N_49748,N_49812);
or UO_1302 (O_1302,N_49780,N_49773);
or UO_1303 (O_1303,N_49686,N_49804);
and UO_1304 (O_1304,N_49978,N_49740);
nor UO_1305 (O_1305,N_49817,N_49502);
and UO_1306 (O_1306,N_49577,N_49558);
xor UO_1307 (O_1307,N_49922,N_49923);
nor UO_1308 (O_1308,N_49647,N_49936);
and UO_1309 (O_1309,N_49890,N_49563);
nor UO_1310 (O_1310,N_49819,N_49805);
nor UO_1311 (O_1311,N_49602,N_49972);
nor UO_1312 (O_1312,N_49627,N_49617);
and UO_1313 (O_1313,N_49797,N_49910);
xnor UO_1314 (O_1314,N_49802,N_49593);
or UO_1315 (O_1315,N_49956,N_49924);
xnor UO_1316 (O_1316,N_49746,N_49966);
nand UO_1317 (O_1317,N_49844,N_49928);
nand UO_1318 (O_1318,N_49832,N_49959);
or UO_1319 (O_1319,N_49792,N_49545);
xor UO_1320 (O_1320,N_49585,N_49600);
nor UO_1321 (O_1321,N_49914,N_49987);
nor UO_1322 (O_1322,N_49828,N_49776);
or UO_1323 (O_1323,N_49791,N_49578);
and UO_1324 (O_1324,N_49655,N_49855);
or UO_1325 (O_1325,N_49849,N_49904);
and UO_1326 (O_1326,N_49576,N_49793);
nand UO_1327 (O_1327,N_49713,N_49806);
nor UO_1328 (O_1328,N_49715,N_49598);
and UO_1329 (O_1329,N_49770,N_49517);
or UO_1330 (O_1330,N_49853,N_49647);
and UO_1331 (O_1331,N_49983,N_49895);
xor UO_1332 (O_1332,N_49803,N_49641);
nand UO_1333 (O_1333,N_49933,N_49658);
nand UO_1334 (O_1334,N_49715,N_49996);
xnor UO_1335 (O_1335,N_49708,N_49670);
or UO_1336 (O_1336,N_49568,N_49605);
nand UO_1337 (O_1337,N_49585,N_49530);
nand UO_1338 (O_1338,N_49893,N_49815);
or UO_1339 (O_1339,N_49858,N_49849);
and UO_1340 (O_1340,N_49800,N_49642);
and UO_1341 (O_1341,N_49544,N_49744);
and UO_1342 (O_1342,N_49952,N_49745);
nand UO_1343 (O_1343,N_49657,N_49530);
nand UO_1344 (O_1344,N_49671,N_49552);
nor UO_1345 (O_1345,N_49625,N_49579);
nand UO_1346 (O_1346,N_49743,N_49642);
nand UO_1347 (O_1347,N_49830,N_49754);
nor UO_1348 (O_1348,N_49682,N_49760);
and UO_1349 (O_1349,N_49634,N_49674);
nor UO_1350 (O_1350,N_49708,N_49963);
nor UO_1351 (O_1351,N_49860,N_49740);
nand UO_1352 (O_1352,N_49981,N_49918);
xor UO_1353 (O_1353,N_49828,N_49928);
nor UO_1354 (O_1354,N_49832,N_49687);
or UO_1355 (O_1355,N_49741,N_49515);
xor UO_1356 (O_1356,N_49926,N_49729);
or UO_1357 (O_1357,N_49973,N_49873);
nor UO_1358 (O_1358,N_49627,N_49685);
or UO_1359 (O_1359,N_49809,N_49803);
nand UO_1360 (O_1360,N_49849,N_49600);
nand UO_1361 (O_1361,N_49863,N_49884);
nor UO_1362 (O_1362,N_49744,N_49702);
xnor UO_1363 (O_1363,N_49514,N_49616);
or UO_1364 (O_1364,N_49511,N_49909);
nand UO_1365 (O_1365,N_49539,N_49930);
nor UO_1366 (O_1366,N_49548,N_49591);
xor UO_1367 (O_1367,N_49511,N_49703);
xnor UO_1368 (O_1368,N_49557,N_49982);
nor UO_1369 (O_1369,N_49789,N_49782);
nand UO_1370 (O_1370,N_49683,N_49536);
or UO_1371 (O_1371,N_49841,N_49986);
nand UO_1372 (O_1372,N_49757,N_49589);
or UO_1373 (O_1373,N_49916,N_49524);
or UO_1374 (O_1374,N_49909,N_49623);
nor UO_1375 (O_1375,N_49932,N_49879);
nor UO_1376 (O_1376,N_49859,N_49695);
nand UO_1377 (O_1377,N_49552,N_49758);
xnor UO_1378 (O_1378,N_49605,N_49649);
or UO_1379 (O_1379,N_49930,N_49812);
and UO_1380 (O_1380,N_49930,N_49641);
nor UO_1381 (O_1381,N_49894,N_49723);
nor UO_1382 (O_1382,N_49582,N_49937);
and UO_1383 (O_1383,N_49844,N_49544);
nand UO_1384 (O_1384,N_49856,N_49872);
xnor UO_1385 (O_1385,N_49759,N_49708);
and UO_1386 (O_1386,N_49785,N_49861);
nor UO_1387 (O_1387,N_49655,N_49603);
xor UO_1388 (O_1388,N_49622,N_49500);
and UO_1389 (O_1389,N_49963,N_49741);
or UO_1390 (O_1390,N_49593,N_49746);
nand UO_1391 (O_1391,N_49584,N_49917);
nor UO_1392 (O_1392,N_49527,N_49574);
or UO_1393 (O_1393,N_49980,N_49771);
nor UO_1394 (O_1394,N_49987,N_49539);
xor UO_1395 (O_1395,N_49731,N_49968);
nand UO_1396 (O_1396,N_49781,N_49568);
xnor UO_1397 (O_1397,N_49808,N_49811);
nor UO_1398 (O_1398,N_49518,N_49632);
and UO_1399 (O_1399,N_49750,N_49902);
nor UO_1400 (O_1400,N_49685,N_49997);
nand UO_1401 (O_1401,N_49748,N_49777);
or UO_1402 (O_1402,N_49657,N_49665);
nor UO_1403 (O_1403,N_49528,N_49687);
and UO_1404 (O_1404,N_49787,N_49527);
or UO_1405 (O_1405,N_49873,N_49874);
and UO_1406 (O_1406,N_49804,N_49934);
and UO_1407 (O_1407,N_49516,N_49828);
nor UO_1408 (O_1408,N_49677,N_49829);
and UO_1409 (O_1409,N_49882,N_49578);
xor UO_1410 (O_1410,N_49845,N_49581);
and UO_1411 (O_1411,N_49836,N_49739);
and UO_1412 (O_1412,N_49683,N_49839);
or UO_1413 (O_1413,N_49771,N_49982);
xnor UO_1414 (O_1414,N_49947,N_49905);
or UO_1415 (O_1415,N_49932,N_49545);
or UO_1416 (O_1416,N_49604,N_49560);
nor UO_1417 (O_1417,N_49582,N_49748);
xnor UO_1418 (O_1418,N_49600,N_49804);
xor UO_1419 (O_1419,N_49731,N_49845);
and UO_1420 (O_1420,N_49626,N_49908);
and UO_1421 (O_1421,N_49526,N_49990);
nor UO_1422 (O_1422,N_49827,N_49855);
or UO_1423 (O_1423,N_49887,N_49742);
and UO_1424 (O_1424,N_49897,N_49858);
xnor UO_1425 (O_1425,N_49798,N_49554);
nand UO_1426 (O_1426,N_49688,N_49572);
or UO_1427 (O_1427,N_49503,N_49664);
or UO_1428 (O_1428,N_49927,N_49730);
xor UO_1429 (O_1429,N_49865,N_49661);
nor UO_1430 (O_1430,N_49894,N_49696);
nand UO_1431 (O_1431,N_49790,N_49606);
xor UO_1432 (O_1432,N_49998,N_49629);
nand UO_1433 (O_1433,N_49900,N_49770);
or UO_1434 (O_1434,N_49901,N_49556);
xnor UO_1435 (O_1435,N_49990,N_49502);
nand UO_1436 (O_1436,N_49779,N_49669);
nor UO_1437 (O_1437,N_49852,N_49940);
xor UO_1438 (O_1438,N_49855,N_49848);
xor UO_1439 (O_1439,N_49508,N_49698);
and UO_1440 (O_1440,N_49554,N_49594);
nand UO_1441 (O_1441,N_49718,N_49554);
and UO_1442 (O_1442,N_49726,N_49983);
nand UO_1443 (O_1443,N_49981,N_49946);
nand UO_1444 (O_1444,N_49753,N_49714);
nand UO_1445 (O_1445,N_49665,N_49566);
and UO_1446 (O_1446,N_49504,N_49977);
nor UO_1447 (O_1447,N_49800,N_49985);
and UO_1448 (O_1448,N_49600,N_49665);
or UO_1449 (O_1449,N_49502,N_49555);
and UO_1450 (O_1450,N_49622,N_49690);
or UO_1451 (O_1451,N_49657,N_49587);
xnor UO_1452 (O_1452,N_49537,N_49956);
nor UO_1453 (O_1453,N_49517,N_49565);
and UO_1454 (O_1454,N_49804,N_49985);
and UO_1455 (O_1455,N_49892,N_49874);
or UO_1456 (O_1456,N_49617,N_49638);
nand UO_1457 (O_1457,N_49844,N_49925);
or UO_1458 (O_1458,N_49654,N_49788);
nor UO_1459 (O_1459,N_49575,N_49519);
xor UO_1460 (O_1460,N_49727,N_49840);
nor UO_1461 (O_1461,N_49636,N_49710);
xor UO_1462 (O_1462,N_49995,N_49813);
nor UO_1463 (O_1463,N_49738,N_49601);
or UO_1464 (O_1464,N_49902,N_49775);
nand UO_1465 (O_1465,N_49514,N_49563);
xor UO_1466 (O_1466,N_49785,N_49991);
xnor UO_1467 (O_1467,N_49609,N_49776);
nand UO_1468 (O_1468,N_49722,N_49680);
and UO_1469 (O_1469,N_49579,N_49962);
nor UO_1470 (O_1470,N_49511,N_49824);
nand UO_1471 (O_1471,N_49787,N_49677);
xor UO_1472 (O_1472,N_49950,N_49701);
xor UO_1473 (O_1473,N_49557,N_49516);
or UO_1474 (O_1474,N_49730,N_49850);
nor UO_1475 (O_1475,N_49885,N_49783);
xor UO_1476 (O_1476,N_49569,N_49943);
or UO_1477 (O_1477,N_49607,N_49952);
and UO_1478 (O_1478,N_49946,N_49660);
xnor UO_1479 (O_1479,N_49926,N_49801);
or UO_1480 (O_1480,N_49505,N_49589);
nor UO_1481 (O_1481,N_49695,N_49618);
nand UO_1482 (O_1482,N_49899,N_49847);
nand UO_1483 (O_1483,N_49923,N_49809);
xnor UO_1484 (O_1484,N_49522,N_49996);
and UO_1485 (O_1485,N_49837,N_49503);
nor UO_1486 (O_1486,N_49582,N_49805);
xor UO_1487 (O_1487,N_49505,N_49739);
nand UO_1488 (O_1488,N_49687,N_49947);
and UO_1489 (O_1489,N_49641,N_49834);
and UO_1490 (O_1490,N_49594,N_49873);
nor UO_1491 (O_1491,N_49641,N_49723);
xnor UO_1492 (O_1492,N_49542,N_49933);
or UO_1493 (O_1493,N_49902,N_49670);
xnor UO_1494 (O_1494,N_49634,N_49803);
or UO_1495 (O_1495,N_49584,N_49546);
nand UO_1496 (O_1496,N_49904,N_49986);
xor UO_1497 (O_1497,N_49984,N_49939);
nor UO_1498 (O_1498,N_49579,N_49819);
xor UO_1499 (O_1499,N_49915,N_49769);
and UO_1500 (O_1500,N_49886,N_49572);
nor UO_1501 (O_1501,N_49951,N_49966);
nand UO_1502 (O_1502,N_49646,N_49616);
nor UO_1503 (O_1503,N_49891,N_49536);
xor UO_1504 (O_1504,N_49687,N_49874);
and UO_1505 (O_1505,N_49582,N_49753);
nor UO_1506 (O_1506,N_49959,N_49689);
and UO_1507 (O_1507,N_49940,N_49530);
nor UO_1508 (O_1508,N_49688,N_49705);
or UO_1509 (O_1509,N_49561,N_49510);
and UO_1510 (O_1510,N_49749,N_49879);
or UO_1511 (O_1511,N_49597,N_49817);
xor UO_1512 (O_1512,N_49684,N_49996);
or UO_1513 (O_1513,N_49938,N_49667);
xor UO_1514 (O_1514,N_49953,N_49866);
or UO_1515 (O_1515,N_49616,N_49982);
and UO_1516 (O_1516,N_49772,N_49787);
nor UO_1517 (O_1517,N_49649,N_49843);
xnor UO_1518 (O_1518,N_49627,N_49942);
xnor UO_1519 (O_1519,N_49910,N_49959);
and UO_1520 (O_1520,N_49575,N_49869);
and UO_1521 (O_1521,N_49549,N_49580);
xor UO_1522 (O_1522,N_49879,N_49785);
xnor UO_1523 (O_1523,N_49616,N_49835);
or UO_1524 (O_1524,N_49517,N_49807);
or UO_1525 (O_1525,N_49914,N_49506);
xor UO_1526 (O_1526,N_49797,N_49650);
nor UO_1527 (O_1527,N_49673,N_49711);
xor UO_1528 (O_1528,N_49772,N_49596);
xnor UO_1529 (O_1529,N_49666,N_49682);
nor UO_1530 (O_1530,N_49519,N_49522);
xnor UO_1531 (O_1531,N_49828,N_49599);
xor UO_1532 (O_1532,N_49533,N_49591);
nor UO_1533 (O_1533,N_49633,N_49884);
or UO_1534 (O_1534,N_49775,N_49604);
nor UO_1535 (O_1535,N_49694,N_49962);
or UO_1536 (O_1536,N_49842,N_49600);
and UO_1537 (O_1537,N_49746,N_49871);
or UO_1538 (O_1538,N_49940,N_49703);
or UO_1539 (O_1539,N_49782,N_49680);
xor UO_1540 (O_1540,N_49700,N_49990);
nand UO_1541 (O_1541,N_49650,N_49988);
and UO_1542 (O_1542,N_49964,N_49796);
nand UO_1543 (O_1543,N_49552,N_49697);
and UO_1544 (O_1544,N_49919,N_49876);
nand UO_1545 (O_1545,N_49656,N_49501);
or UO_1546 (O_1546,N_49556,N_49861);
or UO_1547 (O_1547,N_49624,N_49673);
nand UO_1548 (O_1548,N_49607,N_49987);
or UO_1549 (O_1549,N_49529,N_49944);
nand UO_1550 (O_1550,N_49746,N_49738);
xor UO_1551 (O_1551,N_49716,N_49692);
and UO_1552 (O_1552,N_49651,N_49749);
xnor UO_1553 (O_1553,N_49657,N_49671);
nor UO_1554 (O_1554,N_49926,N_49846);
xor UO_1555 (O_1555,N_49820,N_49681);
xor UO_1556 (O_1556,N_49995,N_49904);
nand UO_1557 (O_1557,N_49812,N_49631);
xor UO_1558 (O_1558,N_49805,N_49709);
nor UO_1559 (O_1559,N_49960,N_49598);
xor UO_1560 (O_1560,N_49912,N_49764);
nor UO_1561 (O_1561,N_49892,N_49541);
or UO_1562 (O_1562,N_49577,N_49845);
nor UO_1563 (O_1563,N_49527,N_49659);
nand UO_1564 (O_1564,N_49840,N_49647);
xnor UO_1565 (O_1565,N_49544,N_49894);
and UO_1566 (O_1566,N_49961,N_49520);
and UO_1567 (O_1567,N_49732,N_49993);
or UO_1568 (O_1568,N_49651,N_49565);
nand UO_1569 (O_1569,N_49856,N_49707);
or UO_1570 (O_1570,N_49889,N_49857);
and UO_1571 (O_1571,N_49765,N_49703);
xor UO_1572 (O_1572,N_49886,N_49955);
nand UO_1573 (O_1573,N_49507,N_49953);
or UO_1574 (O_1574,N_49578,N_49656);
and UO_1575 (O_1575,N_49804,N_49898);
and UO_1576 (O_1576,N_49894,N_49791);
or UO_1577 (O_1577,N_49875,N_49609);
nand UO_1578 (O_1578,N_49704,N_49843);
xor UO_1579 (O_1579,N_49935,N_49518);
xnor UO_1580 (O_1580,N_49638,N_49857);
nor UO_1581 (O_1581,N_49758,N_49802);
nand UO_1582 (O_1582,N_49515,N_49532);
or UO_1583 (O_1583,N_49978,N_49582);
xor UO_1584 (O_1584,N_49589,N_49737);
xnor UO_1585 (O_1585,N_49698,N_49719);
or UO_1586 (O_1586,N_49811,N_49954);
xor UO_1587 (O_1587,N_49561,N_49541);
xor UO_1588 (O_1588,N_49583,N_49501);
or UO_1589 (O_1589,N_49627,N_49689);
and UO_1590 (O_1590,N_49882,N_49525);
nand UO_1591 (O_1591,N_49999,N_49506);
and UO_1592 (O_1592,N_49707,N_49836);
nor UO_1593 (O_1593,N_49939,N_49573);
nor UO_1594 (O_1594,N_49886,N_49907);
xor UO_1595 (O_1595,N_49761,N_49659);
or UO_1596 (O_1596,N_49765,N_49680);
xnor UO_1597 (O_1597,N_49575,N_49713);
and UO_1598 (O_1598,N_49821,N_49650);
xnor UO_1599 (O_1599,N_49836,N_49819);
and UO_1600 (O_1600,N_49746,N_49537);
nor UO_1601 (O_1601,N_49925,N_49794);
nand UO_1602 (O_1602,N_49901,N_49956);
nand UO_1603 (O_1603,N_49643,N_49730);
nor UO_1604 (O_1604,N_49522,N_49921);
or UO_1605 (O_1605,N_49644,N_49683);
nand UO_1606 (O_1606,N_49905,N_49636);
or UO_1607 (O_1607,N_49793,N_49967);
nand UO_1608 (O_1608,N_49807,N_49860);
or UO_1609 (O_1609,N_49935,N_49884);
xor UO_1610 (O_1610,N_49937,N_49575);
nor UO_1611 (O_1611,N_49785,N_49897);
and UO_1612 (O_1612,N_49990,N_49887);
or UO_1613 (O_1613,N_49551,N_49659);
nand UO_1614 (O_1614,N_49694,N_49874);
nor UO_1615 (O_1615,N_49748,N_49770);
nor UO_1616 (O_1616,N_49799,N_49833);
xnor UO_1617 (O_1617,N_49611,N_49738);
nor UO_1618 (O_1618,N_49986,N_49519);
nand UO_1619 (O_1619,N_49649,N_49593);
xor UO_1620 (O_1620,N_49815,N_49610);
xor UO_1621 (O_1621,N_49677,N_49864);
nor UO_1622 (O_1622,N_49819,N_49867);
and UO_1623 (O_1623,N_49870,N_49558);
or UO_1624 (O_1624,N_49624,N_49830);
xnor UO_1625 (O_1625,N_49514,N_49505);
and UO_1626 (O_1626,N_49679,N_49876);
and UO_1627 (O_1627,N_49599,N_49637);
nor UO_1628 (O_1628,N_49997,N_49644);
and UO_1629 (O_1629,N_49929,N_49816);
xor UO_1630 (O_1630,N_49975,N_49761);
and UO_1631 (O_1631,N_49572,N_49522);
or UO_1632 (O_1632,N_49608,N_49965);
nor UO_1633 (O_1633,N_49570,N_49655);
nand UO_1634 (O_1634,N_49709,N_49533);
and UO_1635 (O_1635,N_49699,N_49885);
nand UO_1636 (O_1636,N_49609,N_49798);
xnor UO_1637 (O_1637,N_49555,N_49965);
and UO_1638 (O_1638,N_49659,N_49942);
nor UO_1639 (O_1639,N_49932,N_49528);
and UO_1640 (O_1640,N_49709,N_49573);
or UO_1641 (O_1641,N_49956,N_49666);
nand UO_1642 (O_1642,N_49857,N_49581);
and UO_1643 (O_1643,N_49913,N_49695);
and UO_1644 (O_1644,N_49847,N_49653);
nand UO_1645 (O_1645,N_49993,N_49610);
xor UO_1646 (O_1646,N_49787,N_49539);
and UO_1647 (O_1647,N_49974,N_49575);
nor UO_1648 (O_1648,N_49881,N_49939);
and UO_1649 (O_1649,N_49636,N_49853);
and UO_1650 (O_1650,N_49629,N_49932);
nor UO_1651 (O_1651,N_49510,N_49918);
nor UO_1652 (O_1652,N_49920,N_49654);
xnor UO_1653 (O_1653,N_49539,N_49620);
and UO_1654 (O_1654,N_49821,N_49537);
or UO_1655 (O_1655,N_49610,N_49605);
or UO_1656 (O_1656,N_49657,N_49977);
or UO_1657 (O_1657,N_49652,N_49920);
and UO_1658 (O_1658,N_49728,N_49565);
and UO_1659 (O_1659,N_49983,N_49625);
xnor UO_1660 (O_1660,N_49616,N_49570);
nand UO_1661 (O_1661,N_49876,N_49810);
and UO_1662 (O_1662,N_49757,N_49579);
nor UO_1663 (O_1663,N_49654,N_49553);
nand UO_1664 (O_1664,N_49918,N_49611);
or UO_1665 (O_1665,N_49924,N_49733);
nand UO_1666 (O_1666,N_49932,N_49519);
nand UO_1667 (O_1667,N_49907,N_49734);
and UO_1668 (O_1668,N_49676,N_49877);
xnor UO_1669 (O_1669,N_49958,N_49863);
and UO_1670 (O_1670,N_49668,N_49670);
or UO_1671 (O_1671,N_49765,N_49541);
nor UO_1672 (O_1672,N_49630,N_49810);
nand UO_1673 (O_1673,N_49777,N_49670);
or UO_1674 (O_1674,N_49558,N_49675);
and UO_1675 (O_1675,N_49583,N_49804);
or UO_1676 (O_1676,N_49780,N_49866);
xor UO_1677 (O_1677,N_49879,N_49846);
xnor UO_1678 (O_1678,N_49648,N_49768);
nor UO_1679 (O_1679,N_49508,N_49951);
nand UO_1680 (O_1680,N_49549,N_49525);
xor UO_1681 (O_1681,N_49613,N_49734);
xnor UO_1682 (O_1682,N_49872,N_49827);
and UO_1683 (O_1683,N_49792,N_49617);
xnor UO_1684 (O_1684,N_49555,N_49630);
or UO_1685 (O_1685,N_49799,N_49828);
and UO_1686 (O_1686,N_49719,N_49655);
xnor UO_1687 (O_1687,N_49959,N_49671);
xnor UO_1688 (O_1688,N_49809,N_49871);
nand UO_1689 (O_1689,N_49501,N_49807);
or UO_1690 (O_1690,N_49539,N_49769);
and UO_1691 (O_1691,N_49728,N_49542);
and UO_1692 (O_1692,N_49703,N_49595);
and UO_1693 (O_1693,N_49842,N_49630);
nor UO_1694 (O_1694,N_49764,N_49785);
or UO_1695 (O_1695,N_49808,N_49521);
nor UO_1696 (O_1696,N_49533,N_49994);
xor UO_1697 (O_1697,N_49550,N_49648);
xor UO_1698 (O_1698,N_49760,N_49680);
and UO_1699 (O_1699,N_49502,N_49529);
xor UO_1700 (O_1700,N_49718,N_49739);
or UO_1701 (O_1701,N_49866,N_49726);
xor UO_1702 (O_1702,N_49819,N_49806);
nor UO_1703 (O_1703,N_49693,N_49889);
nor UO_1704 (O_1704,N_49619,N_49922);
nand UO_1705 (O_1705,N_49747,N_49908);
nor UO_1706 (O_1706,N_49579,N_49523);
xor UO_1707 (O_1707,N_49587,N_49918);
nand UO_1708 (O_1708,N_49933,N_49911);
nor UO_1709 (O_1709,N_49757,N_49707);
and UO_1710 (O_1710,N_49811,N_49991);
and UO_1711 (O_1711,N_49705,N_49556);
nand UO_1712 (O_1712,N_49834,N_49523);
and UO_1713 (O_1713,N_49662,N_49899);
nand UO_1714 (O_1714,N_49741,N_49509);
or UO_1715 (O_1715,N_49831,N_49772);
nand UO_1716 (O_1716,N_49809,N_49678);
or UO_1717 (O_1717,N_49697,N_49578);
xnor UO_1718 (O_1718,N_49649,N_49853);
nand UO_1719 (O_1719,N_49726,N_49990);
or UO_1720 (O_1720,N_49900,N_49858);
nand UO_1721 (O_1721,N_49744,N_49897);
nor UO_1722 (O_1722,N_49715,N_49985);
and UO_1723 (O_1723,N_49813,N_49937);
nand UO_1724 (O_1724,N_49690,N_49887);
and UO_1725 (O_1725,N_49528,N_49930);
nand UO_1726 (O_1726,N_49612,N_49966);
and UO_1727 (O_1727,N_49814,N_49791);
nor UO_1728 (O_1728,N_49691,N_49675);
xor UO_1729 (O_1729,N_49932,N_49919);
nand UO_1730 (O_1730,N_49984,N_49838);
nand UO_1731 (O_1731,N_49750,N_49702);
or UO_1732 (O_1732,N_49868,N_49840);
nor UO_1733 (O_1733,N_49925,N_49719);
nand UO_1734 (O_1734,N_49609,N_49763);
nand UO_1735 (O_1735,N_49605,N_49588);
xor UO_1736 (O_1736,N_49844,N_49791);
nand UO_1737 (O_1737,N_49668,N_49693);
xor UO_1738 (O_1738,N_49721,N_49644);
and UO_1739 (O_1739,N_49917,N_49603);
xnor UO_1740 (O_1740,N_49970,N_49892);
nand UO_1741 (O_1741,N_49722,N_49974);
and UO_1742 (O_1742,N_49908,N_49559);
and UO_1743 (O_1743,N_49668,N_49682);
nand UO_1744 (O_1744,N_49873,N_49935);
xnor UO_1745 (O_1745,N_49969,N_49782);
nor UO_1746 (O_1746,N_49758,N_49553);
or UO_1747 (O_1747,N_49680,N_49546);
nor UO_1748 (O_1748,N_49722,N_49921);
or UO_1749 (O_1749,N_49892,N_49569);
nor UO_1750 (O_1750,N_49961,N_49898);
or UO_1751 (O_1751,N_49877,N_49829);
nand UO_1752 (O_1752,N_49677,N_49957);
nand UO_1753 (O_1753,N_49565,N_49732);
nor UO_1754 (O_1754,N_49730,N_49857);
and UO_1755 (O_1755,N_49551,N_49792);
and UO_1756 (O_1756,N_49615,N_49807);
and UO_1757 (O_1757,N_49669,N_49581);
and UO_1758 (O_1758,N_49672,N_49670);
nand UO_1759 (O_1759,N_49500,N_49567);
nand UO_1760 (O_1760,N_49866,N_49566);
and UO_1761 (O_1761,N_49576,N_49722);
nor UO_1762 (O_1762,N_49513,N_49874);
and UO_1763 (O_1763,N_49981,N_49734);
xor UO_1764 (O_1764,N_49949,N_49919);
or UO_1765 (O_1765,N_49673,N_49635);
xnor UO_1766 (O_1766,N_49556,N_49714);
nor UO_1767 (O_1767,N_49509,N_49627);
nor UO_1768 (O_1768,N_49621,N_49822);
and UO_1769 (O_1769,N_49598,N_49527);
or UO_1770 (O_1770,N_49693,N_49509);
or UO_1771 (O_1771,N_49875,N_49982);
or UO_1772 (O_1772,N_49611,N_49580);
and UO_1773 (O_1773,N_49559,N_49915);
and UO_1774 (O_1774,N_49764,N_49776);
nand UO_1775 (O_1775,N_49713,N_49577);
and UO_1776 (O_1776,N_49628,N_49688);
or UO_1777 (O_1777,N_49518,N_49984);
nor UO_1778 (O_1778,N_49596,N_49582);
nand UO_1779 (O_1779,N_49812,N_49501);
xor UO_1780 (O_1780,N_49768,N_49926);
xnor UO_1781 (O_1781,N_49971,N_49668);
nor UO_1782 (O_1782,N_49918,N_49627);
or UO_1783 (O_1783,N_49732,N_49530);
xnor UO_1784 (O_1784,N_49621,N_49595);
nand UO_1785 (O_1785,N_49959,N_49817);
or UO_1786 (O_1786,N_49900,N_49580);
nor UO_1787 (O_1787,N_49571,N_49861);
xnor UO_1788 (O_1788,N_49892,N_49861);
nand UO_1789 (O_1789,N_49901,N_49687);
and UO_1790 (O_1790,N_49898,N_49556);
nor UO_1791 (O_1791,N_49514,N_49710);
nand UO_1792 (O_1792,N_49742,N_49621);
nor UO_1793 (O_1793,N_49551,N_49763);
nand UO_1794 (O_1794,N_49682,N_49785);
xnor UO_1795 (O_1795,N_49664,N_49870);
nor UO_1796 (O_1796,N_49607,N_49981);
nand UO_1797 (O_1797,N_49802,N_49586);
nor UO_1798 (O_1798,N_49717,N_49860);
nor UO_1799 (O_1799,N_49893,N_49968);
xor UO_1800 (O_1800,N_49992,N_49909);
nand UO_1801 (O_1801,N_49693,N_49525);
nor UO_1802 (O_1802,N_49507,N_49739);
nor UO_1803 (O_1803,N_49584,N_49998);
nand UO_1804 (O_1804,N_49927,N_49640);
nand UO_1805 (O_1805,N_49614,N_49695);
nor UO_1806 (O_1806,N_49719,N_49892);
nand UO_1807 (O_1807,N_49638,N_49766);
or UO_1808 (O_1808,N_49927,N_49800);
xnor UO_1809 (O_1809,N_49983,N_49838);
nor UO_1810 (O_1810,N_49611,N_49919);
nand UO_1811 (O_1811,N_49647,N_49977);
xnor UO_1812 (O_1812,N_49960,N_49964);
nand UO_1813 (O_1813,N_49554,N_49843);
nand UO_1814 (O_1814,N_49881,N_49860);
nor UO_1815 (O_1815,N_49536,N_49563);
nor UO_1816 (O_1816,N_49879,N_49903);
and UO_1817 (O_1817,N_49970,N_49779);
or UO_1818 (O_1818,N_49932,N_49688);
xnor UO_1819 (O_1819,N_49805,N_49984);
nand UO_1820 (O_1820,N_49941,N_49841);
or UO_1821 (O_1821,N_49509,N_49676);
or UO_1822 (O_1822,N_49880,N_49976);
nor UO_1823 (O_1823,N_49721,N_49540);
nand UO_1824 (O_1824,N_49667,N_49730);
nor UO_1825 (O_1825,N_49533,N_49802);
nor UO_1826 (O_1826,N_49984,N_49813);
nand UO_1827 (O_1827,N_49782,N_49907);
nor UO_1828 (O_1828,N_49530,N_49508);
and UO_1829 (O_1829,N_49819,N_49597);
or UO_1830 (O_1830,N_49660,N_49501);
and UO_1831 (O_1831,N_49739,N_49845);
nand UO_1832 (O_1832,N_49855,N_49864);
nand UO_1833 (O_1833,N_49807,N_49560);
nor UO_1834 (O_1834,N_49501,N_49818);
xnor UO_1835 (O_1835,N_49546,N_49523);
xor UO_1836 (O_1836,N_49502,N_49618);
xnor UO_1837 (O_1837,N_49558,N_49897);
nor UO_1838 (O_1838,N_49895,N_49602);
nor UO_1839 (O_1839,N_49681,N_49677);
and UO_1840 (O_1840,N_49648,N_49635);
nor UO_1841 (O_1841,N_49827,N_49843);
nor UO_1842 (O_1842,N_49748,N_49730);
or UO_1843 (O_1843,N_49949,N_49514);
and UO_1844 (O_1844,N_49550,N_49780);
or UO_1845 (O_1845,N_49828,N_49835);
or UO_1846 (O_1846,N_49674,N_49592);
or UO_1847 (O_1847,N_49641,N_49774);
nand UO_1848 (O_1848,N_49794,N_49525);
or UO_1849 (O_1849,N_49576,N_49680);
nor UO_1850 (O_1850,N_49686,N_49709);
or UO_1851 (O_1851,N_49691,N_49784);
and UO_1852 (O_1852,N_49856,N_49922);
nand UO_1853 (O_1853,N_49558,N_49729);
nor UO_1854 (O_1854,N_49718,N_49905);
nand UO_1855 (O_1855,N_49525,N_49591);
xnor UO_1856 (O_1856,N_49849,N_49845);
nor UO_1857 (O_1857,N_49544,N_49847);
and UO_1858 (O_1858,N_49560,N_49924);
and UO_1859 (O_1859,N_49773,N_49596);
or UO_1860 (O_1860,N_49693,N_49640);
nand UO_1861 (O_1861,N_49906,N_49521);
nor UO_1862 (O_1862,N_49760,N_49767);
or UO_1863 (O_1863,N_49658,N_49654);
xor UO_1864 (O_1864,N_49762,N_49928);
xor UO_1865 (O_1865,N_49801,N_49500);
or UO_1866 (O_1866,N_49608,N_49988);
or UO_1867 (O_1867,N_49734,N_49964);
nor UO_1868 (O_1868,N_49935,N_49699);
and UO_1869 (O_1869,N_49913,N_49596);
and UO_1870 (O_1870,N_49808,N_49977);
nor UO_1871 (O_1871,N_49810,N_49700);
or UO_1872 (O_1872,N_49793,N_49885);
or UO_1873 (O_1873,N_49677,N_49597);
nand UO_1874 (O_1874,N_49503,N_49922);
nor UO_1875 (O_1875,N_49983,N_49664);
nor UO_1876 (O_1876,N_49635,N_49902);
or UO_1877 (O_1877,N_49983,N_49921);
xor UO_1878 (O_1878,N_49660,N_49724);
or UO_1879 (O_1879,N_49579,N_49799);
and UO_1880 (O_1880,N_49858,N_49974);
nand UO_1881 (O_1881,N_49870,N_49572);
nand UO_1882 (O_1882,N_49778,N_49588);
nor UO_1883 (O_1883,N_49890,N_49790);
xor UO_1884 (O_1884,N_49883,N_49714);
xor UO_1885 (O_1885,N_49587,N_49646);
xnor UO_1886 (O_1886,N_49710,N_49726);
nand UO_1887 (O_1887,N_49872,N_49719);
or UO_1888 (O_1888,N_49765,N_49756);
xnor UO_1889 (O_1889,N_49848,N_49662);
or UO_1890 (O_1890,N_49556,N_49635);
xnor UO_1891 (O_1891,N_49877,N_49509);
nand UO_1892 (O_1892,N_49773,N_49878);
or UO_1893 (O_1893,N_49815,N_49582);
xnor UO_1894 (O_1894,N_49738,N_49827);
xnor UO_1895 (O_1895,N_49887,N_49956);
and UO_1896 (O_1896,N_49500,N_49696);
nor UO_1897 (O_1897,N_49890,N_49791);
xor UO_1898 (O_1898,N_49651,N_49942);
or UO_1899 (O_1899,N_49829,N_49646);
and UO_1900 (O_1900,N_49969,N_49663);
nand UO_1901 (O_1901,N_49735,N_49680);
nor UO_1902 (O_1902,N_49826,N_49866);
xnor UO_1903 (O_1903,N_49731,N_49504);
nand UO_1904 (O_1904,N_49912,N_49500);
and UO_1905 (O_1905,N_49513,N_49618);
nor UO_1906 (O_1906,N_49905,N_49845);
xor UO_1907 (O_1907,N_49875,N_49603);
nand UO_1908 (O_1908,N_49872,N_49724);
xor UO_1909 (O_1909,N_49529,N_49883);
or UO_1910 (O_1910,N_49907,N_49698);
nand UO_1911 (O_1911,N_49698,N_49972);
nor UO_1912 (O_1912,N_49634,N_49958);
nor UO_1913 (O_1913,N_49731,N_49808);
nor UO_1914 (O_1914,N_49851,N_49556);
and UO_1915 (O_1915,N_49544,N_49506);
nand UO_1916 (O_1916,N_49728,N_49811);
or UO_1917 (O_1917,N_49557,N_49841);
and UO_1918 (O_1918,N_49530,N_49924);
xor UO_1919 (O_1919,N_49501,N_49783);
or UO_1920 (O_1920,N_49588,N_49532);
nand UO_1921 (O_1921,N_49784,N_49948);
or UO_1922 (O_1922,N_49761,N_49805);
nor UO_1923 (O_1923,N_49933,N_49873);
or UO_1924 (O_1924,N_49523,N_49797);
nor UO_1925 (O_1925,N_49953,N_49863);
and UO_1926 (O_1926,N_49834,N_49767);
nor UO_1927 (O_1927,N_49775,N_49646);
nor UO_1928 (O_1928,N_49885,N_49548);
and UO_1929 (O_1929,N_49930,N_49541);
nand UO_1930 (O_1930,N_49970,N_49760);
xnor UO_1931 (O_1931,N_49781,N_49820);
or UO_1932 (O_1932,N_49637,N_49946);
or UO_1933 (O_1933,N_49890,N_49605);
or UO_1934 (O_1934,N_49581,N_49796);
and UO_1935 (O_1935,N_49566,N_49723);
and UO_1936 (O_1936,N_49726,N_49603);
nand UO_1937 (O_1937,N_49634,N_49563);
or UO_1938 (O_1938,N_49946,N_49966);
nor UO_1939 (O_1939,N_49878,N_49734);
xor UO_1940 (O_1940,N_49687,N_49974);
xnor UO_1941 (O_1941,N_49587,N_49592);
or UO_1942 (O_1942,N_49636,N_49610);
and UO_1943 (O_1943,N_49550,N_49949);
nor UO_1944 (O_1944,N_49582,N_49878);
and UO_1945 (O_1945,N_49652,N_49688);
or UO_1946 (O_1946,N_49762,N_49583);
and UO_1947 (O_1947,N_49548,N_49963);
xnor UO_1948 (O_1948,N_49718,N_49891);
or UO_1949 (O_1949,N_49753,N_49655);
or UO_1950 (O_1950,N_49845,N_49779);
and UO_1951 (O_1951,N_49547,N_49955);
or UO_1952 (O_1952,N_49932,N_49965);
nor UO_1953 (O_1953,N_49596,N_49766);
or UO_1954 (O_1954,N_49792,N_49721);
xnor UO_1955 (O_1955,N_49861,N_49642);
or UO_1956 (O_1956,N_49893,N_49825);
nor UO_1957 (O_1957,N_49883,N_49674);
or UO_1958 (O_1958,N_49757,N_49965);
nand UO_1959 (O_1959,N_49921,N_49791);
nand UO_1960 (O_1960,N_49860,N_49953);
and UO_1961 (O_1961,N_49778,N_49804);
xnor UO_1962 (O_1962,N_49981,N_49615);
nor UO_1963 (O_1963,N_49580,N_49951);
or UO_1964 (O_1964,N_49686,N_49532);
or UO_1965 (O_1965,N_49700,N_49940);
or UO_1966 (O_1966,N_49527,N_49580);
nor UO_1967 (O_1967,N_49857,N_49809);
nor UO_1968 (O_1968,N_49891,N_49689);
nor UO_1969 (O_1969,N_49567,N_49684);
and UO_1970 (O_1970,N_49741,N_49523);
nand UO_1971 (O_1971,N_49736,N_49600);
and UO_1972 (O_1972,N_49696,N_49658);
xnor UO_1973 (O_1973,N_49903,N_49958);
xnor UO_1974 (O_1974,N_49761,N_49645);
xnor UO_1975 (O_1975,N_49871,N_49816);
nor UO_1976 (O_1976,N_49982,N_49774);
nand UO_1977 (O_1977,N_49681,N_49875);
nand UO_1978 (O_1978,N_49546,N_49618);
nor UO_1979 (O_1979,N_49977,N_49524);
xnor UO_1980 (O_1980,N_49795,N_49702);
and UO_1981 (O_1981,N_49731,N_49658);
nand UO_1982 (O_1982,N_49584,N_49508);
and UO_1983 (O_1983,N_49665,N_49871);
xnor UO_1984 (O_1984,N_49590,N_49679);
and UO_1985 (O_1985,N_49791,N_49815);
xnor UO_1986 (O_1986,N_49994,N_49978);
and UO_1987 (O_1987,N_49849,N_49624);
nor UO_1988 (O_1988,N_49576,N_49838);
nand UO_1989 (O_1989,N_49677,N_49959);
and UO_1990 (O_1990,N_49574,N_49801);
and UO_1991 (O_1991,N_49879,N_49881);
and UO_1992 (O_1992,N_49967,N_49654);
and UO_1993 (O_1993,N_49884,N_49827);
xnor UO_1994 (O_1994,N_49805,N_49593);
and UO_1995 (O_1995,N_49567,N_49721);
or UO_1996 (O_1996,N_49936,N_49577);
and UO_1997 (O_1997,N_49574,N_49865);
nor UO_1998 (O_1998,N_49633,N_49680);
nand UO_1999 (O_1999,N_49933,N_49550);
and UO_2000 (O_2000,N_49662,N_49964);
or UO_2001 (O_2001,N_49647,N_49854);
nand UO_2002 (O_2002,N_49594,N_49749);
or UO_2003 (O_2003,N_49812,N_49765);
xor UO_2004 (O_2004,N_49535,N_49639);
nor UO_2005 (O_2005,N_49782,N_49688);
and UO_2006 (O_2006,N_49980,N_49577);
and UO_2007 (O_2007,N_49773,N_49575);
xnor UO_2008 (O_2008,N_49530,N_49528);
and UO_2009 (O_2009,N_49577,N_49819);
xor UO_2010 (O_2010,N_49659,N_49685);
or UO_2011 (O_2011,N_49910,N_49726);
nor UO_2012 (O_2012,N_49652,N_49655);
nor UO_2013 (O_2013,N_49683,N_49656);
and UO_2014 (O_2014,N_49932,N_49765);
nor UO_2015 (O_2015,N_49911,N_49833);
or UO_2016 (O_2016,N_49726,N_49938);
nand UO_2017 (O_2017,N_49602,N_49879);
and UO_2018 (O_2018,N_49702,N_49599);
nor UO_2019 (O_2019,N_49805,N_49759);
and UO_2020 (O_2020,N_49760,N_49883);
or UO_2021 (O_2021,N_49968,N_49653);
nand UO_2022 (O_2022,N_49707,N_49958);
and UO_2023 (O_2023,N_49672,N_49988);
and UO_2024 (O_2024,N_49853,N_49717);
and UO_2025 (O_2025,N_49833,N_49668);
xnor UO_2026 (O_2026,N_49594,N_49548);
and UO_2027 (O_2027,N_49717,N_49694);
and UO_2028 (O_2028,N_49712,N_49951);
nor UO_2029 (O_2029,N_49813,N_49753);
or UO_2030 (O_2030,N_49813,N_49991);
nor UO_2031 (O_2031,N_49917,N_49788);
or UO_2032 (O_2032,N_49542,N_49697);
or UO_2033 (O_2033,N_49666,N_49633);
nand UO_2034 (O_2034,N_49796,N_49534);
nand UO_2035 (O_2035,N_49708,N_49920);
and UO_2036 (O_2036,N_49707,N_49627);
and UO_2037 (O_2037,N_49770,N_49704);
or UO_2038 (O_2038,N_49977,N_49894);
nor UO_2039 (O_2039,N_49635,N_49707);
xor UO_2040 (O_2040,N_49576,N_49510);
or UO_2041 (O_2041,N_49645,N_49860);
xor UO_2042 (O_2042,N_49915,N_49643);
nor UO_2043 (O_2043,N_49635,N_49692);
nor UO_2044 (O_2044,N_49551,N_49560);
xor UO_2045 (O_2045,N_49549,N_49513);
nor UO_2046 (O_2046,N_49832,N_49941);
nor UO_2047 (O_2047,N_49944,N_49858);
nand UO_2048 (O_2048,N_49558,N_49539);
nor UO_2049 (O_2049,N_49674,N_49793);
and UO_2050 (O_2050,N_49943,N_49558);
nor UO_2051 (O_2051,N_49750,N_49809);
or UO_2052 (O_2052,N_49746,N_49630);
nor UO_2053 (O_2053,N_49870,N_49874);
nor UO_2054 (O_2054,N_49694,N_49731);
xnor UO_2055 (O_2055,N_49977,N_49928);
or UO_2056 (O_2056,N_49928,N_49571);
xnor UO_2057 (O_2057,N_49874,N_49997);
xnor UO_2058 (O_2058,N_49556,N_49669);
and UO_2059 (O_2059,N_49741,N_49957);
or UO_2060 (O_2060,N_49800,N_49632);
nand UO_2061 (O_2061,N_49848,N_49977);
nor UO_2062 (O_2062,N_49873,N_49849);
nand UO_2063 (O_2063,N_49958,N_49723);
nand UO_2064 (O_2064,N_49611,N_49904);
and UO_2065 (O_2065,N_49512,N_49810);
or UO_2066 (O_2066,N_49992,N_49754);
and UO_2067 (O_2067,N_49680,N_49833);
nand UO_2068 (O_2068,N_49815,N_49641);
or UO_2069 (O_2069,N_49511,N_49918);
or UO_2070 (O_2070,N_49803,N_49740);
xnor UO_2071 (O_2071,N_49696,N_49539);
nor UO_2072 (O_2072,N_49954,N_49764);
nand UO_2073 (O_2073,N_49578,N_49945);
or UO_2074 (O_2074,N_49774,N_49666);
nand UO_2075 (O_2075,N_49980,N_49722);
and UO_2076 (O_2076,N_49637,N_49840);
xor UO_2077 (O_2077,N_49895,N_49975);
nand UO_2078 (O_2078,N_49966,N_49713);
nand UO_2079 (O_2079,N_49510,N_49728);
or UO_2080 (O_2080,N_49619,N_49865);
nor UO_2081 (O_2081,N_49696,N_49776);
and UO_2082 (O_2082,N_49901,N_49814);
xor UO_2083 (O_2083,N_49893,N_49765);
nor UO_2084 (O_2084,N_49957,N_49876);
and UO_2085 (O_2085,N_49775,N_49834);
or UO_2086 (O_2086,N_49868,N_49951);
xnor UO_2087 (O_2087,N_49802,N_49849);
nor UO_2088 (O_2088,N_49941,N_49833);
xnor UO_2089 (O_2089,N_49695,N_49548);
and UO_2090 (O_2090,N_49730,N_49865);
nor UO_2091 (O_2091,N_49943,N_49519);
nor UO_2092 (O_2092,N_49501,N_49856);
nor UO_2093 (O_2093,N_49805,N_49637);
nor UO_2094 (O_2094,N_49514,N_49555);
or UO_2095 (O_2095,N_49981,N_49680);
and UO_2096 (O_2096,N_49832,N_49916);
and UO_2097 (O_2097,N_49646,N_49626);
nor UO_2098 (O_2098,N_49887,N_49708);
nand UO_2099 (O_2099,N_49586,N_49772);
nor UO_2100 (O_2100,N_49842,N_49644);
nor UO_2101 (O_2101,N_49982,N_49734);
nor UO_2102 (O_2102,N_49622,N_49592);
nor UO_2103 (O_2103,N_49945,N_49933);
xor UO_2104 (O_2104,N_49993,N_49759);
xor UO_2105 (O_2105,N_49835,N_49539);
or UO_2106 (O_2106,N_49531,N_49919);
nor UO_2107 (O_2107,N_49703,N_49694);
and UO_2108 (O_2108,N_49783,N_49897);
xor UO_2109 (O_2109,N_49584,N_49786);
and UO_2110 (O_2110,N_49884,N_49963);
and UO_2111 (O_2111,N_49926,N_49685);
xor UO_2112 (O_2112,N_49707,N_49972);
nand UO_2113 (O_2113,N_49771,N_49674);
nor UO_2114 (O_2114,N_49813,N_49931);
or UO_2115 (O_2115,N_49839,N_49985);
nor UO_2116 (O_2116,N_49744,N_49576);
or UO_2117 (O_2117,N_49581,N_49972);
nor UO_2118 (O_2118,N_49803,N_49768);
xor UO_2119 (O_2119,N_49544,N_49866);
nand UO_2120 (O_2120,N_49984,N_49705);
and UO_2121 (O_2121,N_49804,N_49773);
nor UO_2122 (O_2122,N_49912,N_49849);
and UO_2123 (O_2123,N_49880,N_49788);
or UO_2124 (O_2124,N_49939,N_49908);
xnor UO_2125 (O_2125,N_49700,N_49956);
and UO_2126 (O_2126,N_49855,N_49999);
or UO_2127 (O_2127,N_49859,N_49852);
nand UO_2128 (O_2128,N_49566,N_49959);
xnor UO_2129 (O_2129,N_49665,N_49897);
xnor UO_2130 (O_2130,N_49744,N_49901);
nor UO_2131 (O_2131,N_49826,N_49675);
xor UO_2132 (O_2132,N_49744,N_49931);
xnor UO_2133 (O_2133,N_49527,N_49925);
and UO_2134 (O_2134,N_49789,N_49757);
and UO_2135 (O_2135,N_49718,N_49967);
and UO_2136 (O_2136,N_49839,N_49543);
nor UO_2137 (O_2137,N_49852,N_49613);
and UO_2138 (O_2138,N_49861,N_49746);
and UO_2139 (O_2139,N_49837,N_49999);
nand UO_2140 (O_2140,N_49570,N_49545);
nand UO_2141 (O_2141,N_49938,N_49840);
or UO_2142 (O_2142,N_49656,N_49647);
and UO_2143 (O_2143,N_49933,N_49838);
and UO_2144 (O_2144,N_49975,N_49881);
and UO_2145 (O_2145,N_49924,N_49701);
or UO_2146 (O_2146,N_49778,N_49969);
or UO_2147 (O_2147,N_49658,N_49838);
and UO_2148 (O_2148,N_49813,N_49705);
nor UO_2149 (O_2149,N_49909,N_49563);
and UO_2150 (O_2150,N_49864,N_49599);
or UO_2151 (O_2151,N_49546,N_49861);
or UO_2152 (O_2152,N_49630,N_49881);
or UO_2153 (O_2153,N_49565,N_49897);
nand UO_2154 (O_2154,N_49573,N_49967);
or UO_2155 (O_2155,N_49679,N_49718);
nor UO_2156 (O_2156,N_49937,N_49972);
nor UO_2157 (O_2157,N_49588,N_49751);
xnor UO_2158 (O_2158,N_49626,N_49570);
nor UO_2159 (O_2159,N_49725,N_49762);
nand UO_2160 (O_2160,N_49640,N_49842);
xnor UO_2161 (O_2161,N_49947,N_49737);
xnor UO_2162 (O_2162,N_49998,N_49917);
nand UO_2163 (O_2163,N_49905,N_49887);
nor UO_2164 (O_2164,N_49791,N_49558);
xnor UO_2165 (O_2165,N_49599,N_49723);
or UO_2166 (O_2166,N_49929,N_49869);
nand UO_2167 (O_2167,N_49766,N_49743);
and UO_2168 (O_2168,N_49839,N_49617);
and UO_2169 (O_2169,N_49769,N_49863);
or UO_2170 (O_2170,N_49978,N_49618);
nand UO_2171 (O_2171,N_49682,N_49749);
xnor UO_2172 (O_2172,N_49594,N_49973);
nor UO_2173 (O_2173,N_49929,N_49623);
or UO_2174 (O_2174,N_49855,N_49598);
or UO_2175 (O_2175,N_49605,N_49613);
xnor UO_2176 (O_2176,N_49904,N_49729);
nand UO_2177 (O_2177,N_49593,N_49738);
or UO_2178 (O_2178,N_49845,N_49647);
or UO_2179 (O_2179,N_49687,N_49529);
nor UO_2180 (O_2180,N_49701,N_49792);
nand UO_2181 (O_2181,N_49900,N_49771);
or UO_2182 (O_2182,N_49881,N_49608);
nand UO_2183 (O_2183,N_49860,N_49862);
nand UO_2184 (O_2184,N_49702,N_49906);
and UO_2185 (O_2185,N_49638,N_49924);
or UO_2186 (O_2186,N_49852,N_49963);
xor UO_2187 (O_2187,N_49825,N_49521);
xnor UO_2188 (O_2188,N_49784,N_49638);
xor UO_2189 (O_2189,N_49982,N_49920);
or UO_2190 (O_2190,N_49691,N_49612);
and UO_2191 (O_2191,N_49810,N_49586);
nand UO_2192 (O_2192,N_49693,N_49502);
nor UO_2193 (O_2193,N_49669,N_49877);
nor UO_2194 (O_2194,N_49760,N_49502);
or UO_2195 (O_2195,N_49730,N_49517);
xor UO_2196 (O_2196,N_49710,N_49980);
nor UO_2197 (O_2197,N_49718,N_49892);
xnor UO_2198 (O_2198,N_49747,N_49793);
nand UO_2199 (O_2199,N_49666,N_49579);
xnor UO_2200 (O_2200,N_49564,N_49766);
and UO_2201 (O_2201,N_49684,N_49854);
nor UO_2202 (O_2202,N_49745,N_49762);
xor UO_2203 (O_2203,N_49742,N_49902);
or UO_2204 (O_2204,N_49692,N_49923);
and UO_2205 (O_2205,N_49699,N_49504);
xor UO_2206 (O_2206,N_49807,N_49832);
and UO_2207 (O_2207,N_49597,N_49793);
or UO_2208 (O_2208,N_49633,N_49801);
or UO_2209 (O_2209,N_49630,N_49548);
nand UO_2210 (O_2210,N_49726,N_49851);
and UO_2211 (O_2211,N_49767,N_49741);
xor UO_2212 (O_2212,N_49729,N_49864);
xnor UO_2213 (O_2213,N_49764,N_49557);
nor UO_2214 (O_2214,N_49839,N_49890);
nand UO_2215 (O_2215,N_49892,N_49875);
nor UO_2216 (O_2216,N_49890,N_49771);
nor UO_2217 (O_2217,N_49893,N_49790);
nand UO_2218 (O_2218,N_49839,N_49798);
xor UO_2219 (O_2219,N_49753,N_49770);
nor UO_2220 (O_2220,N_49823,N_49555);
nand UO_2221 (O_2221,N_49511,N_49746);
xor UO_2222 (O_2222,N_49641,N_49996);
and UO_2223 (O_2223,N_49883,N_49866);
nor UO_2224 (O_2224,N_49877,N_49973);
or UO_2225 (O_2225,N_49600,N_49810);
and UO_2226 (O_2226,N_49986,N_49910);
xor UO_2227 (O_2227,N_49845,N_49996);
and UO_2228 (O_2228,N_49819,N_49998);
and UO_2229 (O_2229,N_49504,N_49888);
and UO_2230 (O_2230,N_49742,N_49920);
nor UO_2231 (O_2231,N_49967,N_49598);
or UO_2232 (O_2232,N_49548,N_49696);
nand UO_2233 (O_2233,N_49622,N_49671);
nand UO_2234 (O_2234,N_49605,N_49690);
nor UO_2235 (O_2235,N_49991,N_49994);
nor UO_2236 (O_2236,N_49784,N_49839);
nor UO_2237 (O_2237,N_49906,N_49587);
nor UO_2238 (O_2238,N_49684,N_49895);
nor UO_2239 (O_2239,N_49917,N_49540);
or UO_2240 (O_2240,N_49674,N_49764);
nor UO_2241 (O_2241,N_49894,N_49640);
nor UO_2242 (O_2242,N_49533,N_49933);
nor UO_2243 (O_2243,N_49575,N_49552);
xnor UO_2244 (O_2244,N_49858,N_49531);
nand UO_2245 (O_2245,N_49980,N_49925);
or UO_2246 (O_2246,N_49612,N_49565);
nand UO_2247 (O_2247,N_49731,N_49558);
nor UO_2248 (O_2248,N_49771,N_49986);
and UO_2249 (O_2249,N_49924,N_49827);
nand UO_2250 (O_2250,N_49673,N_49750);
xor UO_2251 (O_2251,N_49746,N_49898);
or UO_2252 (O_2252,N_49691,N_49549);
nor UO_2253 (O_2253,N_49662,N_49971);
and UO_2254 (O_2254,N_49852,N_49923);
xnor UO_2255 (O_2255,N_49766,N_49730);
nand UO_2256 (O_2256,N_49774,N_49848);
xnor UO_2257 (O_2257,N_49766,N_49628);
nor UO_2258 (O_2258,N_49981,N_49949);
nand UO_2259 (O_2259,N_49597,N_49620);
nor UO_2260 (O_2260,N_49654,N_49727);
nand UO_2261 (O_2261,N_49890,N_49531);
xor UO_2262 (O_2262,N_49658,N_49549);
xnor UO_2263 (O_2263,N_49653,N_49951);
and UO_2264 (O_2264,N_49814,N_49699);
and UO_2265 (O_2265,N_49733,N_49728);
nor UO_2266 (O_2266,N_49957,N_49917);
or UO_2267 (O_2267,N_49703,N_49987);
xnor UO_2268 (O_2268,N_49827,N_49938);
or UO_2269 (O_2269,N_49584,N_49883);
nor UO_2270 (O_2270,N_49816,N_49681);
or UO_2271 (O_2271,N_49820,N_49522);
or UO_2272 (O_2272,N_49985,N_49872);
or UO_2273 (O_2273,N_49923,N_49826);
xnor UO_2274 (O_2274,N_49615,N_49832);
nand UO_2275 (O_2275,N_49574,N_49993);
nor UO_2276 (O_2276,N_49967,N_49644);
nand UO_2277 (O_2277,N_49521,N_49849);
or UO_2278 (O_2278,N_49914,N_49722);
nor UO_2279 (O_2279,N_49981,N_49877);
and UO_2280 (O_2280,N_49686,N_49970);
nor UO_2281 (O_2281,N_49590,N_49920);
and UO_2282 (O_2282,N_49504,N_49605);
nand UO_2283 (O_2283,N_49899,N_49815);
nand UO_2284 (O_2284,N_49994,N_49597);
or UO_2285 (O_2285,N_49812,N_49539);
nor UO_2286 (O_2286,N_49648,N_49790);
and UO_2287 (O_2287,N_49641,N_49780);
nand UO_2288 (O_2288,N_49754,N_49764);
nand UO_2289 (O_2289,N_49897,N_49836);
and UO_2290 (O_2290,N_49695,N_49686);
or UO_2291 (O_2291,N_49649,N_49861);
xnor UO_2292 (O_2292,N_49704,N_49948);
nand UO_2293 (O_2293,N_49680,N_49733);
nand UO_2294 (O_2294,N_49648,N_49835);
and UO_2295 (O_2295,N_49590,N_49759);
or UO_2296 (O_2296,N_49543,N_49730);
nor UO_2297 (O_2297,N_49891,N_49618);
and UO_2298 (O_2298,N_49602,N_49965);
and UO_2299 (O_2299,N_49623,N_49661);
nand UO_2300 (O_2300,N_49654,N_49536);
and UO_2301 (O_2301,N_49578,N_49821);
nor UO_2302 (O_2302,N_49973,N_49608);
and UO_2303 (O_2303,N_49599,N_49956);
or UO_2304 (O_2304,N_49694,N_49939);
xnor UO_2305 (O_2305,N_49772,N_49574);
nor UO_2306 (O_2306,N_49600,N_49778);
and UO_2307 (O_2307,N_49642,N_49682);
xor UO_2308 (O_2308,N_49666,N_49797);
nor UO_2309 (O_2309,N_49585,N_49875);
nor UO_2310 (O_2310,N_49666,N_49968);
nor UO_2311 (O_2311,N_49704,N_49816);
nand UO_2312 (O_2312,N_49640,N_49887);
nand UO_2313 (O_2313,N_49502,N_49999);
and UO_2314 (O_2314,N_49748,N_49962);
or UO_2315 (O_2315,N_49646,N_49963);
nand UO_2316 (O_2316,N_49654,N_49906);
nand UO_2317 (O_2317,N_49705,N_49958);
xnor UO_2318 (O_2318,N_49845,N_49693);
nand UO_2319 (O_2319,N_49663,N_49944);
nor UO_2320 (O_2320,N_49952,N_49699);
nand UO_2321 (O_2321,N_49708,N_49795);
or UO_2322 (O_2322,N_49613,N_49915);
and UO_2323 (O_2323,N_49748,N_49909);
nor UO_2324 (O_2324,N_49727,N_49571);
xor UO_2325 (O_2325,N_49745,N_49784);
nor UO_2326 (O_2326,N_49754,N_49954);
or UO_2327 (O_2327,N_49578,N_49646);
and UO_2328 (O_2328,N_49673,N_49870);
and UO_2329 (O_2329,N_49748,N_49775);
and UO_2330 (O_2330,N_49625,N_49860);
xnor UO_2331 (O_2331,N_49663,N_49665);
or UO_2332 (O_2332,N_49594,N_49946);
nand UO_2333 (O_2333,N_49860,N_49525);
and UO_2334 (O_2334,N_49757,N_49576);
nand UO_2335 (O_2335,N_49750,N_49921);
nand UO_2336 (O_2336,N_49803,N_49880);
nand UO_2337 (O_2337,N_49865,N_49841);
xnor UO_2338 (O_2338,N_49593,N_49508);
nand UO_2339 (O_2339,N_49709,N_49645);
or UO_2340 (O_2340,N_49548,N_49737);
xnor UO_2341 (O_2341,N_49910,N_49885);
xnor UO_2342 (O_2342,N_49609,N_49632);
nand UO_2343 (O_2343,N_49882,N_49774);
nor UO_2344 (O_2344,N_49984,N_49677);
nor UO_2345 (O_2345,N_49916,N_49708);
nor UO_2346 (O_2346,N_49722,N_49534);
xor UO_2347 (O_2347,N_49825,N_49838);
xor UO_2348 (O_2348,N_49974,N_49597);
nand UO_2349 (O_2349,N_49959,N_49917);
and UO_2350 (O_2350,N_49658,N_49726);
nor UO_2351 (O_2351,N_49790,N_49805);
and UO_2352 (O_2352,N_49519,N_49588);
or UO_2353 (O_2353,N_49655,N_49884);
nand UO_2354 (O_2354,N_49606,N_49792);
or UO_2355 (O_2355,N_49694,N_49584);
nor UO_2356 (O_2356,N_49970,N_49949);
xor UO_2357 (O_2357,N_49958,N_49777);
or UO_2358 (O_2358,N_49515,N_49562);
xor UO_2359 (O_2359,N_49869,N_49818);
nor UO_2360 (O_2360,N_49572,N_49893);
or UO_2361 (O_2361,N_49814,N_49847);
or UO_2362 (O_2362,N_49925,N_49596);
and UO_2363 (O_2363,N_49813,N_49875);
nor UO_2364 (O_2364,N_49724,N_49720);
xnor UO_2365 (O_2365,N_49972,N_49589);
and UO_2366 (O_2366,N_49646,N_49583);
nand UO_2367 (O_2367,N_49830,N_49757);
xor UO_2368 (O_2368,N_49587,N_49649);
nor UO_2369 (O_2369,N_49600,N_49522);
nor UO_2370 (O_2370,N_49568,N_49923);
xor UO_2371 (O_2371,N_49601,N_49721);
xor UO_2372 (O_2372,N_49946,N_49796);
or UO_2373 (O_2373,N_49664,N_49995);
and UO_2374 (O_2374,N_49754,N_49731);
or UO_2375 (O_2375,N_49539,N_49775);
and UO_2376 (O_2376,N_49949,N_49675);
or UO_2377 (O_2377,N_49610,N_49814);
or UO_2378 (O_2378,N_49770,N_49562);
and UO_2379 (O_2379,N_49726,N_49718);
or UO_2380 (O_2380,N_49598,N_49590);
xor UO_2381 (O_2381,N_49712,N_49643);
nand UO_2382 (O_2382,N_49771,N_49742);
and UO_2383 (O_2383,N_49639,N_49614);
nand UO_2384 (O_2384,N_49754,N_49882);
xor UO_2385 (O_2385,N_49747,N_49720);
xnor UO_2386 (O_2386,N_49910,N_49504);
or UO_2387 (O_2387,N_49776,N_49502);
xnor UO_2388 (O_2388,N_49802,N_49747);
or UO_2389 (O_2389,N_49825,N_49870);
nor UO_2390 (O_2390,N_49567,N_49623);
nand UO_2391 (O_2391,N_49695,N_49564);
or UO_2392 (O_2392,N_49733,N_49675);
nand UO_2393 (O_2393,N_49584,N_49609);
xor UO_2394 (O_2394,N_49996,N_49667);
nor UO_2395 (O_2395,N_49585,N_49503);
or UO_2396 (O_2396,N_49524,N_49533);
nand UO_2397 (O_2397,N_49788,N_49538);
or UO_2398 (O_2398,N_49844,N_49772);
nand UO_2399 (O_2399,N_49859,N_49874);
nand UO_2400 (O_2400,N_49595,N_49503);
nand UO_2401 (O_2401,N_49911,N_49627);
xnor UO_2402 (O_2402,N_49955,N_49629);
or UO_2403 (O_2403,N_49661,N_49596);
nand UO_2404 (O_2404,N_49747,N_49790);
nand UO_2405 (O_2405,N_49532,N_49969);
or UO_2406 (O_2406,N_49547,N_49998);
xnor UO_2407 (O_2407,N_49544,N_49711);
or UO_2408 (O_2408,N_49636,N_49969);
nor UO_2409 (O_2409,N_49907,N_49863);
xor UO_2410 (O_2410,N_49765,N_49557);
xnor UO_2411 (O_2411,N_49732,N_49942);
or UO_2412 (O_2412,N_49583,N_49607);
nor UO_2413 (O_2413,N_49542,N_49616);
nor UO_2414 (O_2414,N_49772,N_49857);
and UO_2415 (O_2415,N_49903,N_49741);
or UO_2416 (O_2416,N_49643,N_49916);
nand UO_2417 (O_2417,N_49634,N_49688);
xnor UO_2418 (O_2418,N_49746,N_49872);
nand UO_2419 (O_2419,N_49797,N_49532);
xnor UO_2420 (O_2420,N_49554,N_49684);
xnor UO_2421 (O_2421,N_49733,N_49937);
nand UO_2422 (O_2422,N_49587,N_49837);
and UO_2423 (O_2423,N_49953,N_49901);
xnor UO_2424 (O_2424,N_49721,N_49599);
nand UO_2425 (O_2425,N_49663,N_49609);
nand UO_2426 (O_2426,N_49588,N_49802);
nor UO_2427 (O_2427,N_49840,N_49561);
nor UO_2428 (O_2428,N_49981,N_49603);
nor UO_2429 (O_2429,N_49930,N_49808);
nor UO_2430 (O_2430,N_49950,N_49639);
xor UO_2431 (O_2431,N_49520,N_49776);
or UO_2432 (O_2432,N_49595,N_49951);
xor UO_2433 (O_2433,N_49906,N_49552);
nand UO_2434 (O_2434,N_49951,N_49599);
nand UO_2435 (O_2435,N_49602,N_49726);
nor UO_2436 (O_2436,N_49636,N_49767);
nor UO_2437 (O_2437,N_49761,N_49992);
nand UO_2438 (O_2438,N_49899,N_49956);
xor UO_2439 (O_2439,N_49861,N_49949);
and UO_2440 (O_2440,N_49744,N_49960);
or UO_2441 (O_2441,N_49719,N_49661);
or UO_2442 (O_2442,N_49528,N_49785);
and UO_2443 (O_2443,N_49740,N_49931);
or UO_2444 (O_2444,N_49587,N_49560);
or UO_2445 (O_2445,N_49800,N_49870);
nor UO_2446 (O_2446,N_49541,N_49510);
and UO_2447 (O_2447,N_49871,N_49842);
xnor UO_2448 (O_2448,N_49830,N_49818);
nor UO_2449 (O_2449,N_49818,N_49769);
xnor UO_2450 (O_2450,N_49646,N_49812);
xor UO_2451 (O_2451,N_49709,N_49942);
or UO_2452 (O_2452,N_49704,N_49969);
xor UO_2453 (O_2453,N_49607,N_49908);
xor UO_2454 (O_2454,N_49895,N_49724);
and UO_2455 (O_2455,N_49559,N_49912);
nor UO_2456 (O_2456,N_49785,N_49641);
and UO_2457 (O_2457,N_49752,N_49599);
and UO_2458 (O_2458,N_49924,N_49727);
xor UO_2459 (O_2459,N_49793,N_49562);
or UO_2460 (O_2460,N_49879,N_49761);
or UO_2461 (O_2461,N_49763,N_49906);
nor UO_2462 (O_2462,N_49707,N_49910);
nor UO_2463 (O_2463,N_49921,N_49694);
and UO_2464 (O_2464,N_49623,N_49955);
nor UO_2465 (O_2465,N_49587,N_49796);
and UO_2466 (O_2466,N_49933,N_49773);
and UO_2467 (O_2467,N_49753,N_49768);
or UO_2468 (O_2468,N_49800,N_49704);
nor UO_2469 (O_2469,N_49528,N_49948);
nand UO_2470 (O_2470,N_49940,N_49640);
nand UO_2471 (O_2471,N_49943,N_49687);
or UO_2472 (O_2472,N_49525,N_49833);
or UO_2473 (O_2473,N_49540,N_49725);
nand UO_2474 (O_2474,N_49662,N_49718);
or UO_2475 (O_2475,N_49657,N_49924);
and UO_2476 (O_2476,N_49574,N_49862);
or UO_2477 (O_2477,N_49778,N_49951);
or UO_2478 (O_2478,N_49697,N_49629);
nor UO_2479 (O_2479,N_49609,N_49878);
xor UO_2480 (O_2480,N_49976,N_49911);
xnor UO_2481 (O_2481,N_49576,N_49608);
and UO_2482 (O_2482,N_49894,N_49671);
nor UO_2483 (O_2483,N_49835,N_49734);
and UO_2484 (O_2484,N_49839,N_49603);
and UO_2485 (O_2485,N_49793,N_49614);
or UO_2486 (O_2486,N_49708,N_49737);
or UO_2487 (O_2487,N_49809,N_49838);
xor UO_2488 (O_2488,N_49980,N_49838);
and UO_2489 (O_2489,N_49949,N_49931);
nor UO_2490 (O_2490,N_49968,N_49696);
xnor UO_2491 (O_2491,N_49766,N_49613);
nor UO_2492 (O_2492,N_49925,N_49869);
and UO_2493 (O_2493,N_49919,N_49812);
nand UO_2494 (O_2494,N_49872,N_49583);
nand UO_2495 (O_2495,N_49983,N_49735);
xor UO_2496 (O_2496,N_49972,N_49703);
xnor UO_2497 (O_2497,N_49630,N_49654);
or UO_2498 (O_2498,N_49590,N_49588);
xnor UO_2499 (O_2499,N_49961,N_49970);
xor UO_2500 (O_2500,N_49781,N_49915);
or UO_2501 (O_2501,N_49837,N_49572);
and UO_2502 (O_2502,N_49652,N_49693);
nand UO_2503 (O_2503,N_49699,N_49872);
or UO_2504 (O_2504,N_49940,N_49857);
xor UO_2505 (O_2505,N_49800,N_49533);
and UO_2506 (O_2506,N_49597,N_49664);
nand UO_2507 (O_2507,N_49971,N_49992);
or UO_2508 (O_2508,N_49708,N_49799);
nand UO_2509 (O_2509,N_49949,N_49894);
xnor UO_2510 (O_2510,N_49509,N_49656);
nand UO_2511 (O_2511,N_49984,N_49933);
or UO_2512 (O_2512,N_49709,N_49559);
or UO_2513 (O_2513,N_49937,N_49981);
xnor UO_2514 (O_2514,N_49663,N_49946);
nand UO_2515 (O_2515,N_49519,N_49658);
nor UO_2516 (O_2516,N_49833,N_49656);
nand UO_2517 (O_2517,N_49766,N_49782);
nand UO_2518 (O_2518,N_49973,N_49779);
or UO_2519 (O_2519,N_49556,N_49548);
and UO_2520 (O_2520,N_49658,N_49816);
or UO_2521 (O_2521,N_49613,N_49589);
nand UO_2522 (O_2522,N_49767,N_49604);
nand UO_2523 (O_2523,N_49763,N_49630);
nor UO_2524 (O_2524,N_49566,N_49549);
or UO_2525 (O_2525,N_49685,N_49958);
xor UO_2526 (O_2526,N_49570,N_49573);
or UO_2527 (O_2527,N_49629,N_49647);
nand UO_2528 (O_2528,N_49851,N_49529);
and UO_2529 (O_2529,N_49513,N_49679);
or UO_2530 (O_2530,N_49741,N_49521);
nand UO_2531 (O_2531,N_49607,N_49851);
nand UO_2532 (O_2532,N_49863,N_49517);
and UO_2533 (O_2533,N_49856,N_49949);
and UO_2534 (O_2534,N_49821,N_49859);
and UO_2535 (O_2535,N_49723,N_49841);
or UO_2536 (O_2536,N_49992,N_49544);
nor UO_2537 (O_2537,N_49838,N_49867);
nor UO_2538 (O_2538,N_49932,N_49857);
xnor UO_2539 (O_2539,N_49890,N_49539);
nor UO_2540 (O_2540,N_49821,N_49677);
xnor UO_2541 (O_2541,N_49942,N_49670);
and UO_2542 (O_2542,N_49746,N_49968);
nand UO_2543 (O_2543,N_49991,N_49569);
nand UO_2544 (O_2544,N_49736,N_49653);
xor UO_2545 (O_2545,N_49764,N_49730);
nand UO_2546 (O_2546,N_49714,N_49744);
and UO_2547 (O_2547,N_49799,N_49890);
xor UO_2548 (O_2548,N_49742,N_49908);
nor UO_2549 (O_2549,N_49919,N_49935);
nor UO_2550 (O_2550,N_49882,N_49969);
nand UO_2551 (O_2551,N_49736,N_49566);
nor UO_2552 (O_2552,N_49853,N_49875);
xor UO_2553 (O_2553,N_49653,N_49938);
nand UO_2554 (O_2554,N_49779,N_49735);
nor UO_2555 (O_2555,N_49695,N_49826);
nor UO_2556 (O_2556,N_49811,N_49675);
nand UO_2557 (O_2557,N_49538,N_49533);
nor UO_2558 (O_2558,N_49695,N_49982);
and UO_2559 (O_2559,N_49713,N_49645);
and UO_2560 (O_2560,N_49884,N_49885);
and UO_2561 (O_2561,N_49936,N_49749);
nor UO_2562 (O_2562,N_49987,N_49586);
nand UO_2563 (O_2563,N_49500,N_49518);
and UO_2564 (O_2564,N_49850,N_49734);
nor UO_2565 (O_2565,N_49891,N_49992);
and UO_2566 (O_2566,N_49999,N_49777);
and UO_2567 (O_2567,N_49703,N_49733);
and UO_2568 (O_2568,N_49653,N_49969);
nor UO_2569 (O_2569,N_49653,N_49966);
xor UO_2570 (O_2570,N_49853,N_49870);
nor UO_2571 (O_2571,N_49907,N_49677);
nor UO_2572 (O_2572,N_49812,N_49784);
nand UO_2573 (O_2573,N_49633,N_49852);
or UO_2574 (O_2574,N_49772,N_49544);
or UO_2575 (O_2575,N_49591,N_49741);
xor UO_2576 (O_2576,N_49553,N_49861);
nor UO_2577 (O_2577,N_49771,N_49504);
nor UO_2578 (O_2578,N_49580,N_49688);
xor UO_2579 (O_2579,N_49984,N_49837);
nor UO_2580 (O_2580,N_49577,N_49804);
or UO_2581 (O_2581,N_49880,N_49972);
or UO_2582 (O_2582,N_49687,N_49760);
or UO_2583 (O_2583,N_49987,N_49649);
xor UO_2584 (O_2584,N_49824,N_49763);
xor UO_2585 (O_2585,N_49584,N_49551);
xor UO_2586 (O_2586,N_49564,N_49804);
xor UO_2587 (O_2587,N_49788,N_49522);
or UO_2588 (O_2588,N_49925,N_49623);
nor UO_2589 (O_2589,N_49879,N_49617);
and UO_2590 (O_2590,N_49916,N_49757);
or UO_2591 (O_2591,N_49552,N_49869);
or UO_2592 (O_2592,N_49697,N_49992);
xnor UO_2593 (O_2593,N_49857,N_49781);
nor UO_2594 (O_2594,N_49908,N_49597);
and UO_2595 (O_2595,N_49516,N_49983);
and UO_2596 (O_2596,N_49990,N_49858);
xor UO_2597 (O_2597,N_49506,N_49636);
nand UO_2598 (O_2598,N_49567,N_49616);
and UO_2599 (O_2599,N_49658,N_49758);
or UO_2600 (O_2600,N_49960,N_49882);
or UO_2601 (O_2601,N_49869,N_49934);
nand UO_2602 (O_2602,N_49994,N_49784);
and UO_2603 (O_2603,N_49730,N_49585);
and UO_2604 (O_2604,N_49745,N_49749);
xnor UO_2605 (O_2605,N_49981,N_49913);
nor UO_2606 (O_2606,N_49587,N_49935);
and UO_2607 (O_2607,N_49633,N_49694);
or UO_2608 (O_2608,N_49780,N_49533);
nand UO_2609 (O_2609,N_49857,N_49656);
nand UO_2610 (O_2610,N_49915,N_49910);
and UO_2611 (O_2611,N_49604,N_49625);
or UO_2612 (O_2612,N_49792,N_49749);
and UO_2613 (O_2613,N_49889,N_49559);
xnor UO_2614 (O_2614,N_49599,N_49591);
and UO_2615 (O_2615,N_49800,N_49692);
xor UO_2616 (O_2616,N_49848,N_49984);
or UO_2617 (O_2617,N_49562,N_49965);
or UO_2618 (O_2618,N_49679,N_49608);
or UO_2619 (O_2619,N_49511,N_49758);
and UO_2620 (O_2620,N_49938,N_49556);
and UO_2621 (O_2621,N_49911,N_49705);
nand UO_2622 (O_2622,N_49552,N_49563);
or UO_2623 (O_2623,N_49611,N_49683);
or UO_2624 (O_2624,N_49919,N_49623);
xor UO_2625 (O_2625,N_49687,N_49792);
xor UO_2626 (O_2626,N_49681,N_49708);
xnor UO_2627 (O_2627,N_49602,N_49676);
nand UO_2628 (O_2628,N_49620,N_49774);
xor UO_2629 (O_2629,N_49915,N_49793);
nor UO_2630 (O_2630,N_49648,N_49909);
nand UO_2631 (O_2631,N_49952,N_49803);
and UO_2632 (O_2632,N_49618,N_49570);
nand UO_2633 (O_2633,N_49786,N_49714);
and UO_2634 (O_2634,N_49694,N_49565);
or UO_2635 (O_2635,N_49837,N_49510);
xor UO_2636 (O_2636,N_49783,N_49698);
or UO_2637 (O_2637,N_49599,N_49620);
and UO_2638 (O_2638,N_49991,N_49956);
and UO_2639 (O_2639,N_49875,N_49789);
and UO_2640 (O_2640,N_49822,N_49993);
nor UO_2641 (O_2641,N_49702,N_49505);
nand UO_2642 (O_2642,N_49830,N_49904);
nand UO_2643 (O_2643,N_49790,N_49869);
xor UO_2644 (O_2644,N_49609,N_49880);
and UO_2645 (O_2645,N_49628,N_49856);
nor UO_2646 (O_2646,N_49560,N_49622);
or UO_2647 (O_2647,N_49737,N_49678);
xor UO_2648 (O_2648,N_49877,N_49621);
and UO_2649 (O_2649,N_49530,N_49543);
xnor UO_2650 (O_2650,N_49901,N_49944);
nand UO_2651 (O_2651,N_49956,N_49727);
and UO_2652 (O_2652,N_49535,N_49933);
and UO_2653 (O_2653,N_49946,N_49590);
nand UO_2654 (O_2654,N_49519,N_49814);
xor UO_2655 (O_2655,N_49609,N_49738);
or UO_2656 (O_2656,N_49979,N_49955);
xnor UO_2657 (O_2657,N_49590,N_49688);
nand UO_2658 (O_2658,N_49851,N_49863);
nor UO_2659 (O_2659,N_49502,N_49589);
and UO_2660 (O_2660,N_49806,N_49755);
xor UO_2661 (O_2661,N_49587,N_49728);
nor UO_2662 (O_2662,N_49688,N_49577);
and UO_2663 (O_2663,N_49715,N_49730);
nand UO_2664 (O_2664,N_49804,N_49929);
nor UO_2665 (O_2665,N_49610,N_49969);
or UO_2666 (O_2666,N_49861,N_49833);
nor UO_2667 (O_2667,N_49565,N_49718);
and UO_2668 (O_2668,N_49688,N_49821);
and UO_2669 (O_2669,N_49713,N_49536);
xor UO_2670 (O_2670,N_49848,N_49740);
and UO_2671 (O_2671,N_49849,N_49727);
or UO_2672 (O_2672,N_49865,N_49882);
xor UO_2673 (O_2673,N_49638,N_49500);
xor UO_2674 (O_2674,N_49841,N_49650);
nor UO_2675 (O_2675,N_49955,N_49930);
and UO_2676 (O_2676,N_49571,N_49970);
nor UO_2677 (O_2677,N_49552,N_49798);
nor UO_2678 (O_2678,N_49998,N_49826);
nand UO_2679 (O_2679,N_49802,N_49597);
or UO_2680 (O_2680,N_49948,N_49909);
nand UO_2681 (O_2681,N_49807,N_49610);
nor UO_2682 (O_2682,N_49672,N_49626);
nand UO_2683 (O_2683,N_49888,N_49643);
xnor UO_2684 (O_2684,N_49940,N_49569);
or UO_2685 (O_2685,N_49612,N_49995);
and UO_2686 (O_2686,N_49815,N_49649);
or UO_2687 (O_2687,N_49675,N_49822);
nand UO_2688 (O_2688,N_49769,N_49524);
and UO_2689 (O_2689,N_49736,N_49988);
and UO_2690 (O_2690,N_49687,N_49921);
xor UO_2691 (O_2691,N_49803,N_49814);
or UO_2692 (O_2692,N_49964,N_49745);
and UO_2693 (O_2693,N_49741,N_49608);
xnor UO_2694 (O_2694,N_49998,N_49855);
xnor UO_2695 (O_2695,N_49982,N_49535);
nor UO_2696 (O_2696,N_49776,N_49561);
nor UO_2697 (O_2697,N_49637,N_49784);
and UO_2698 (O_2698,N_49549,N_49675);
xnor UO_2699 (O_2699,N_49534,N_49803);
nand UO_2700 (O_2700,N_49677,N_49740);
nor UO_2701 (O_2701,N_49509,N_49587);
or UO_2702 (O_2702,N_49907,N_49571);
xor UO_2703 (O_2703,N_49917,N_49983);
xor UO_2704 (O_2704,N_49940,N_49536);
and UO_2705 (O_2705,N_49664,N_49785);
and UO_2706 (O_2706,N_49761,N_49673);
or UO_2707 (O_2707,N_49651,N_49624);
xor UO_2708 (O_2708,N_49618,N_49921);
or UO_2709 (O_2709,N_49737,N_49673);
xnor UO_2710 (O_2710,N_49648,N_49519);
and UO_2711 (O_2711,N_49589,N_49648);
xor UO_2712 (O_2712,N_49826,N_49988);
and UO_2713 (O_2713,N_49548,N_49571);
or UO_2714 (O_2714,N_49624,N_49619);
xor UO_2715 (O_2715,N_49888,N_49618);
and UO_2716 (O_2716,N_49799,N_49558);
or UO_2717 (O_2717,N_49754,N_49919);
xnor UO_2718 (O_2718,N_49605,N_49700);
or UO_2719 (O_2719,N_49607,N_49839);
nor UO_2720 (O_2720,N_49606,N_49946);
nand UO_2721 (O_2721,N_49574,N_49566);
or UO_2722 (O_2722,N_49521,N_49919);
and UO_2723 (O_2723,N_49901,N_49807);
xor UO_2724 (O_2724,N_49624,N_49757);
xor UO_2725 (O_2725,N_49954,N_49748);
and UO_2726 (O_2726,N_49554,N_49783);
nor UO_2727 (O_2727,N_49679,N_49524);
xnor UO_2728 (O_2728,N_49791,N_49986);
xor UO_2729 (O_2729,N_49508,N_49903);
nor UO_2730 (O_2730,N_49548,N_49500);
nand UO_2731 (O_2731,N_49909,N_49696);
or UO_2732 (O_2732,N_49592,N_49714);
and UO_2733 (O_2733,N_49796,N_49844);
or UO_2734 (O_2734,N_49962,N_49701);
xor UO_2735 (O_2735,N_49860,N_49671);
nand UO_2736 (O_2736,N_49618,N_49521);
and UO_2737 (O_2737,N_49523,N_49836);
nor UO_2738 (O_2738,N_49872,N_49838);
or UO_2739 (O_2739,N_49601,N_49531);
and UO_2740 (O_2740,N_49900,N_49509);
or UO_2741 (O_2741,N_49995,N_49903);
nor UO_2742 (O_2742,N_49800,N_49910);
and UO_2743 (O_2743,N_49686,N_49922);
nor UO_2744 (O_2744,N_49673,N_49778);
nand UO_2745 (O_2745,N_49760,N_49928);
nand UO_2746 (O_2746,N_49754,N_49810);
nor UO_2747 (O_2747,N_49738,N_49926);
xor UO_2748 (O_2748,N_49779,N_49563);
and UO_2749 (O_2749,N_49717,N_49548);
and UO_2750 (O_2750,N_49627,N_49533);
and UO_2751 (O_2751,N_49694,N_49822);
nor UO_2752 (O_2752,N_49691,N_49740);
nor UO_2753 (O_2753,N_49932,N_49652);
and UO_2754 (O_2754,N_49529,N_49573);
nand UO_2755 (O_2755,N_49686,N_49946);
xor UO_2756 (O_2756,N_49826,N_49559);
nand UO_2757 (O_2757,N_49542,N_49762);
nand UO_2758 (O_2758,N_49618,N_49525);
nand UO_2759 (O_2759,N_49566,N_49601);
or UO_2760 (O_2760,N_49578,N_49587);
or UO_2761 (O_2761,N_49772,N_49781);
nand UO_2762 (O_2762,N_49576,N_49925);
xor UO_2763 (O_2763,N_49729,N_49822);
nand UO_2764 (O_2764,N_49614,N_49629);
or UO_2765 (O_2765,N_49887,N_49784);
nor UO_2766 (O_2766,N_49803,N_49961);
or UO_2767 (O_2767,N_49674,N_49920);
nand UO_2768 (O_2768,N_49600,N_49845);
and UO_2769 (O_2769,N_49907,N_49831);
and UO_2770 (O_2770,N_49615,N_49936);
and UO_2771 (O_2771,N_49512,N_49576);
nand UO_2772 (O_2772,N_49972,N_49856);
xor UO_2773 (O_2773,N_49557,N_49980);
and UO_2774 (O_2774,N_49938,N_49926);
xor UO_2775 (O_2775,N_49575,N_49787);
and UO_2776 (O_2776,N_49951,N_49747);
xor UO_2777 (O_2777,N_49653,N_49555);
or UO_2778 (O_2778,N_49836,N_49622);
nand UO_2779 (O_2779,N_49592,N_49777);
nand UO_2780 (O_2780,N_49728,N_49603);
and UO_2781 (O_2781,N_49873,N_49901);
nand UO_2782 (O_2782,N_49619,N_49826);
and UO_2783 (O_2783,N_49738,N_49677);
xor UO_2784 (O_2784,N_49890,N_49856);
xnor UO_2785 (O_2785,N_49822,N_49895);
xnor UO_2786 (O_2786,N_49773,N_49940);
nor UO_2787 (O_2787,N_49625,N_49510);
and UO_2788 (O_2788,N_49700,N_49530);
xor UO_2789 (O_2789,N_49899,N_49652);
xnor UO_2790 (O_2790,N_49597,N_49625);
or UO_2791 (O_2791,N_49823,N_49571);
and UO_2792 (O_2792,N_49866,N_49513);
and UO_2793 (O_2793,N_49956,N_49931);
xnor UO_2794 (O_2794,N_49990,N_49967);
nand UO_2795 (O_2795,N_49514,N_49775);
and UO_2796 (O_2796,N_49605,N_49692);
nand UO_2797 (O_2797,N_49987,N_49922);
and UO_2798 (O_2798,N_49686,N_49801);
nand UO_2799 (O_2799,N_49872,N_49590);
and UO_2800 (O_2800,N_49924,N_49799);
nor UO_2801 (O_2801,N_49807,N_49628);
nand UO_2802 (O_2802,N_49526,N_49648);
nand UO_2803 (O_2803,N_49661,N_49534);
or UO_2804 (O_2804,N_49635,N_49521);
and UO_2805 (O_2805,N_49870,N_49663);
xnor UO_2806 (O_2806,N_49635,N_49657);
or UO_2807 (O_2807,N_49938,N_49789);
nand UO_2808 (O_2808,N_49684,N_49778);
xor UO_2809 (O_2809,N_49965,N_49775);
nor UO_2810 (O_2810,N_49970,N_49661);
or UO_2811 (O_2811,N_49829,N_49602);
nand UO_2812 (O_2812,N_49704,N_49626);
nand UO_2813 (O_2813,N_49674,N_49922);
and UO_2814 (O_2814,N_49767,N_49943);
nor UO_2815 (O_2815,N_49564,N_49581);
nor UO_2816 (O_2816,N_49799,N_49560);
and UO_2817 (O_2817,N_49886,N_49688);
or UO_2818 (O_2818,N_49757,N_49506);
and UO_2819 (O_2819,N_49714,N_49921);
or UO_2820 (O_2820,N_49604,N_49517);
nand UO_2821 (O_2821,N_49502,N_49899);
nand UO_2822 (O_2822,N_49938,N_49715);
nand UO_2823 (O_2823,N_49841,N_49520);
or UO_2824 (O_2824,N_49721,N_49995);
and UO_2825 (O_2825,N_49898,N_49656);
or UO_2826 (O_2826,N_49846,N_49991);
nand UO_2827 (O_2827,N_49891,N_49546);
xor UO_2828 (O_2828,N_49871,N_49639);
and UO_2829 (O_2829,N_49980,N_49581);
or UO_2830 (O_2830,N_49625,N_49748);
nor UO_2831 (O_2831,N_49759,N_49734);
or UO_2832 (O_2832,N_49698,N_49837);
or UO_2833 (O_2833,N_49613,N_49978);
or UO_2834 (O_2834,N_49521,N_49957);
xnor UO_2835 (O_2835,N_49599,N_49803);
nor UO_2836 (O_2836,N_49522,N_49592);
and UO_2837 (O_2837,N_49558,N_49992);
or UO_2838 (O_2838,N_49635,N_49700);
nand UO_2839 (O_2839,N_49543,N_49891);
xor UO_2840 (O_2840,N_49548,N_49595);
xor UO_2841 (O_2841,N_49875,N_49924);
nor UO_2842 (O_2842,N_49891,N_49548);
nand UO_2843 (O_2843,N_49558,N_49528);
nand UO_2844 (O_2844,N_49997,N_49502);
nand UO_2845 (O_2845,N_49948,N_49993);
and UO_2846 (O_2846,N_49528,N_49517);
nor UO_2847 (O_2847,N_49773,N_49624);
and UO_2848 (O_2848,N_49711,N_49963);
or UO_2849 (O_2849,N_49607,N_49721);
nor UO_2850 (O_2850,N_49830,N_49540);
nand UO_2851 (O_2851,N_49577,N_49643);
xor UO_2852 (O_2852,N_49563,N_49554);
xnor UO_2853 (O_2853,N_49654,N_49549);
nor UO_2854 (O_2854,N_49826,N_49595);
nor UO_2855 (O_2855,N_49808,N_49658);
xor UO_2856 (O_2856,N_49674,N_49716);
nor UO_2857 (O_2857,N_49835,N_49930);
and UO_2858 (O_2858,N_49566,N_49898);
nor UO_2859 (O_2859,N_49884,N_49644);
nor UO_2860 (O_2860,N_49930,N_49648);
or UO_2861 (O_2861,N_49762,N_49682);
nor UO_2862 (O_2862,N_49738,N_49777);
nand UO_2863 (O_2863,N_49506,N_49558);
and UO_2864 (O_2864,N_49624,N_49680);
xnor UO_2865 (O_2865,N_49996,N_49787);
and UO_2866 (O_2866,N_49856,N_49573);
and UO_2867 (O_2867,N_49914,N_49794);
or UO_2868 (O_2868,N_49577,N_49878);
nor UO_2869 (O_2869,N_49951,N_49813);
or UO_2870 (O_2870,N_49845,N_49744);
xor UO_2871 (O_2871,N_49540,N_49680);
and UO_2872 (O_2872,N_49981,N_49991);
and UO_2873 (O_2873,N_49670,N_49821);
nor UO_2874 (O_2874,N_49583,N_49624);
xor UO_2875 (O_2875,N_49580,N_49568);
nand UO_2876 (O_2876,N_49592,N_49880);
xnor UO_2877 (O_2877,N_49867,N_49994);
and UO_2878 (O_2878,N_49565,N_49993);
nand UO_2879 (O_2879,N_49899,N_49854);
nand UO_2880 (O_2880,N_49965,N_49588);
nand UO_2881 (O_2881,N_49570,N_49515);
xnor UO_2882 (O_2882,N_49860,N_49980);
nand UO_2883 (O_2883,N_49726,N_49948);
nor UO_2884 (O_2884,N_49867,N_49587);
xor UO_2885 (O_2885,N_49594,N_49924);
and UO_2886 (O_2886,N_49566,N_49809);
and UO_2887 (O_2887,N_49725,N_49575);
nor UO_2888 (O_2888,N_49658,N_49566);
or UO_2889 (O_2889,N_49836,N_49641);
and UO_2890 (O_2890,N_49863,N_49770);
and UO_2891 (O_2891,N_49885,N_49599);
nor UO_2892 (O_2892,N_49757,N_49893);
nand UO_2893 (O_2893,N_49936,N_49943);
and UO_2894 (O_2894,N_49978,N_49991);
nor UO_2895 (O_2895,N_49896,N_49649);
and UO_2896 (O_2896,N_49959,N_49570);
and UO_2897 (O_2897,N_49625,N_49814);
and UO_2898 (O_2898,N_49747,N_49604);
or UO_2899 (O_2899,N_49828,N_49667);
nor UO_2900 (O_2900,N_49623,N_49958);
or UO_2901 (O_2901,N_49790,N_49902);
and UO_2902 (O_2902,N_49626,N_49781);
xor UO_2903 (O_2903,N_49807,N_49743);
and UO_2904 (O_2904,N_49845,N_49801);
xnor UO_2905 (O_2905,N_49927,N_49619);
and UO_2906 (O_2906,N_49774,N_49754);
and UO_2907 (O_2907,N_49941,N_49985);
nor UO_2908 (O_2908,N_49749,N_49869);
and UO_2909 (O_2909,N_49670,N_49809);
xor UO_2910 (O_2910,N_49856,N_49532);
nand UO_2911 (O_2911,N_49602,N_49635);
nor UO_2912 (O_2912,N_49509,N_49928);
nor UO_2913 (O_2913,N_49967,N_49774);
nor UO_2914 (O_2914,N_49936,N_49901);
or UO_2915 (O_2915,N_49896,N_49628);
nor UO_2916 (O_2916,N_49801,N_49629);
and UO_2917 (O_2917,N_49704,N_49775);
nor UO_2918 (O_2918,N_49528,N_49723);
and UO_2919 (O_2919,N_49756,N_49668);
nor UO_2920 (O_2920,N_49756,N_49982);
nor UO_2921 (O_2921,N_49532,N_49652);
and UO_2922 (O_2922,N_49600,N_49739);
and UO_2923 (O_2923,N_49959,N_49584);
nand UO_2924 (O_2924,N_49623,N_49721);
xor UO_2925 (O_2925,N_49785,N_49585);
or UO_2926 (O_2926,N_49912,N_49554);
or UO_2927 (O_2927,N_49956,N_49635);
nor UO_2928 (O_2928,N_49629,N_49876);
nand UO_2929 (O_2929,N_49829,N_49742);
and UO_2930 (O_2930,N_49610,N_49839);
xnor UO_2931 (O_2931,N_49763,N_49858);
nand UO_2932 (O_2932,N_49657,N_49674);
nor UO_2933 (O_2933,N_49655,N_49576);
and UO_2934 (O_2934,N_49902,N_49554);
or UO_2935 (O_2935,N_49796,N_49944);
nand UO_2936 (O_2936,N_49532,N_49658);
nand UO_2937 (O_2937,N_49715,N_49915);
nor UO_2938 (O_2938,N_49697,N_49812);
xnor UO_2939 (O_2939,N_49503,N_49963);
or UO_2940 (O_2940,N_49714,N_49819);
or UO_2941 (O_2941,N_49733,N_49649);
and UO_2942 (O_2942,N_49891,N_49708);
xor UO_2943 (O_2943,N_49902,N_49709);
nor UO_2944 (O_2944,N_49591,N_49534);
xor UO_2945 (O_2945,N_49861,N_49648);
nor UO_2946 (O_2946,N_49680,N_49584);
and UO_2947 (O_2947,N_49790,N_49993);
or UO_2948 (O_2948,N_49610,N_49590);
and UO_2949 (O_2949,N_49926,N_49868);
xnor UO_2950 (O_2950,N_49754,N_49519);
or UO_2951 (O_2951,N_49542,N_49966);
and UO_2952 (O_2952,N_49648,N_49645);
nand UO_2953 (O_2953,N_49898,N_49657);
xnor UO_2954 (O_2954,N_49966,N_49510);
nand UO_2955 (O_2955,N_49905,N_49759);
xor UO_2956 (O_2956,N_49541,N_49527);
and UO_2957 (O_2957,N_49695,N_49999);
nor UO_2958 (O_2958,N_49535,N_49818);
xnor UO_2959 (O_2959,N_49627,N_49992);
xnor UO_2960 (O_2960,N_49556,N_49910);
xor UO_2961 (O_2961,N_49656,N_49691);
nand UO_2962 (O_2962,N_49988,N_49519);
nor UO_2963 (O_2963,N_49733,N_49674);
nand UO_2964 (O_2964,N_49568,N_49937);
and UO_2965 (O_2965,N_49841,N_49738);
nand UO_2966 (O_2966,N_49524,N_49685);
and UO_2967 (O_2967,N_49554,N_49575);
xnor UO_2968 (O_2968,N_49641,N_49913);
or UO_2969 (O_2969,N_49794,N_49577);
nor UO_2970 (O_2970,N_49920,N_49786);
or UO_2971 (O_2971,N_49881,N_49535);
nor UO_2972 (O_2972,N_49802,N_49536);
nand UO_2973 (O_2973,N_49694,N_49856);
nor UO_2974 (O_2974,N_49940,N_49587);
and UO_2975 (O_2975,N_49872,N_49552);
nor UO_2976 (O_2976,N_49861,N_49608);
and UO_2977 (O_2977,N_49847,N_49744);
and UO_2978 (O_2978,N_49632,N_49951);
nor UO_2979 (O_2979,N_49821,N_49953);
nor UO_2980 (O_2980,N_49788,N_49750);
nor UO_2981 (O_2981,N_49832,N_49686);
nor UO_2982 (O_2982,N_49522,N_49705);
or UO_2983 (O_2983,N_49795,N_49784);
or UO_2984 (O_2984,N_49722,N_49928);
and UO_2985 (O_2985,N_49882,N_49965);
or UO_2986 (O_2986,N_49906,N_49779);
and UO_2987 (O_2987,N_49751,N_49835);
nand UO_2988 (O_2988,N_49648,N_49818);
or UO_2989 (O_2989,N_49831,N_49739);
xnor UO_2990 (O_2990,N_49532,N_49908);
nand UO_2991 (O_2991,N_49922,N_49701);
and UO_2992 (O_2992,N_49805,N_49960);
nor UO_2993 (O_2993,N_49710,N_49735);
and UO_2994 (O_2994,N_49692,N_49932);
nor UO_2995 (O_2995,N_49941,N_49917);
xnor UO_2996 (O_2996,N_49881,N_49681);
nor UO_2997 (O_2997,N_49845,N_49783);
nor UO_2998 (O_2998,N_49543,N_49566);
or UO_2999 (O_2999,N_49854,N_49518);
nand UO_3000 (O_3000,N_49795,N_49564);
nand UO_3001 (O_3001,N_49961,N_49858);
and UO_3002 (O_3002,N_49802,N_49631);
nand UO_3003 (O_3003,N_49633,N_49509);
or UO_3004 (O_3004,N_49952,N_49638);
nand UO_3005 (O_3005,N_49798,N_49611);
and UO_3006 (O_3006,N_49759,N_49689);
nand UO_3007 (O_3007,N_49858,N_49516);
nor UO_3008 (O_3008,N_49861,N_49540);
xnor UO_3009 (O_3009,N_49677,N_49560);
nand UO_3010 (O_3010,N_49598,N_49932);
or UO_3011 (O_3011,N_49554,N_49850);
or UO_3012 (O_3012,N_49536,N_49638);
nand UO_3013 (O_3013,N_49658,N_49693);
and UO_3014 (O_3014,N_49718,N_49936);
xnor UO_3015 (O_3015,N_49744,N_49763);
nand UO_3016 (O_3016,N_49836,N_49575);
or UO_3017 (O_3017,N_49772,N_49592);
nand UO_3018 (O_3018,N_49819,N_49848);
or UO_3019 (O_3019,N_49543,N_49865);
nor UO_3020 (O_3020,N_49697,N_49939);
nand UO_3021 (O_3021,N_49856,N_49967);
xor UO_3022 (O_3022,N_49692,N_49964);
xor UO_3023 (O_3023,N_49517,N_49511);
and UO_3024 (O_3024,N_49621,N_49512);
and UO_3025 (O_3025,N_49641,N_49868);
xnor UO_3026 (O_3026,N_49584,N_49839);
xnor UO_3027 (O_3027,N_49724,N_49638);
and UO_3028 (O_3028,N_49515,N_49551);
xor UO_3029 (O_3029,N_49711,N_49599);
nor UO_3030 (O_3030,N_49880,N_49829);
nand UO_3031 (O_3031,N_49849,N_49688);
nor UO_3032 (O_3032,N_49763,N_49973);
and UO_3033 (O_3033,N_49716,N_49904);
nand UO_3034 (O_3034,N_49710,N_49847);
and UO_3035 (O_3035,N_49898,N_49587);
nor UO_3036 (O_3036,N_49866,N_49622);
nand UO_3037 (O_3037,N_49727,N_49554);
nor UO_3038 (O_3038,N_49547,N_49617);
xor UO_3039 (O_3039,N_49887,N_49665);
and UO_3040 (O_3040,N_49969,N_49895);
and UO_3041 (O_3041,N_49747,N_49876);
nor UO_3042 (O_3042,N_49736,N_49891);
nand UO_3043 (O_3043,N_49627,N_49612);
or UO_3044 (O_3044,N_49760,N_49540);
nand UO_3045 (O_3045,N_49973,N_49749);
or UO_3046 (O_3046,N_49531,N_49974);
nand UO_3047 (O_3047,N_49990,N_49824);
and UO_3048 (O_3048,N_49941,N_49763);
xnor UO_3049 (O_3049,N_49940,N_49884);
nor UO_3050 (O_3050,N_49739,N_49652);
or UO_3051 (O_3051,N_49927,N_49936);
xor UO_3052 (O_3052,N_49546,N_49774);
xnor UO_3053 (O_3053,N_49649,N_49922);
nand UO_3054 (O_3054,N_49970,N_49916);
and UO_3055 (O_3055,N_49771,N_49631);
nor UO_3056 (O_3056,N_49566,N_49716);
and UO_3057 (O_3057,N_49619,N_49875);
and UO_3058 (O_3058,N_49852,N_49519);
nor UO_3059 (O_3059,N_49618,N_49810);
nor UO_3060 (O_3060,N_49897,N_49592);
nand UO_3061 (O_3061,N_49908,N_49502);
or UO_3062 (O_3062,N_49818,N_49968);
nor UO_3063 (O_3063,N_49711,N_49999);
or UO_3064 (O_3064,N_49657,N_49809);
or UO_3065 (O_3065,N_49707,N_49745);
nor UO_3066 (O_3066,N_49731,N_49890);
nor UO_3067 (O_3067,N_49623,N_49746);
or UO_3068 (O_3068,N_49904,N_49775);
or UO_3069 (O_3069,N_49989,N_49954);
and UO_3070 (O_3070,N_49970,N_49573);
xor UO_3071 (O_3071,N_49845,N_49870);
nor UO_3072 (O_3072,N_49578,N_49874);
nand UO_3073 (O_3073,N_49894,N_49763);
nand UO_3074 (O_3074,N_49736,N_49706);
and UO_3075 (O_3075,N_49645,N_49844);
xnor UO_3076 (O_3076,N_49992,N_49872);
nor UO_3077 (O_3077,N_49587,N_49736);
or UO_3078 (O_3078,N_49652,N_49603);
nor UO_3079 (O_3079,N_49573,N_49664);
xor UO_3080 (O_3080,N_49838,N_49583);
xnor UO_3081 (O_3081,N_49627,N_49981);
nor UO_3082 (O_3082,N_49705,N_49625);
or UO_3083 (O_3083,N_49934,N_49927);
nor UO_3084 (O_3084,N_49909,N_49937);
xor UO_3085 (O_3085,N_49720,N_49626);
and UO_3086 (O_3086,N_49954,N_49732);
nand UO_3087 (O_3087,N_49972,N_49685);
nand UO_3088 (O_3088,N_49853,N_49855);
and UO_3089 (O_3089,N_49699,N_49597);
nand UO_3090 (O_3090,N_49786,N_49596);
xnor UO_3091 (O_3091,N_49875,N_49656);
nand UO_3092 (O_3092,N_49802,N_49608);
nand UO_3093 (O_3093,N_49854,N_49865);
nand UO_3094 (O_3094,N_49644,N_49654);
or UO_3095 (O_3095,N_49633,N_49999);
nand UO_3096 (O_3096,N_49504,N_49654);
nor UO_3097 (O_3097,N_49518,N_49920);
nor UO_3098 (O_3098,N_49787,N_49874);
xnor UO_3099 (O_3099,N_49614,N_49527);
and UO_3100 (O_3100,N_49810,N_49803);
xnor UO_3101 (O_3101,N_49502,N_49569);
xor UO_3102 (O_3102,N_49623,N_49786);
nand UO_3103 (O_3103,N_49820,N_49984);
nor UO_3104 (O_3104,N_49868,N_49952);
nor UO_3105 (O_3105,N_49581,N_49836);
or UO_3106 (O_3106,N_49590,N_49800);
and UO_3107 (O_3107,N_49510,N_49773);
nand UO_3108 (O_3108,N_49597,N_49934);
nand UO_3109 (O_3109,N_49510,N_49768);
and UO_3110 (O_3110,N_49796,N_49514);
nor UO_3111 (O_3111,N_49930,N_49510);
or UO_3112 (O_3112,N_49798,N_49927);
and UO_3113 (O_3113,N_49779,N_49642);
xor UO_3114 (O_3114,N_49655,N_49672);
nor UO_3115 (O_3115,N_49519,N_49601);
and UO_3116 (O_3116,N_49550,N_49574);
and UO_3117 (O_3117,N_49662,N_49746);
and UO_3118 (O_3118,N_49642,N_49954);
or UO_3119 (O_3119,N_49675,N_49882);
xor UO_3120 (O_3120,N_49608,N_49622);
and UO_3121 (O_3121,N_49566,N_49662);
xor UO_3122 (O_3122,N_49884,N_49513);
or UO_3123 (O_3123,N_49900,N_49531);
or UO_3124 (O_3124,N_49956,N_49632);
or UO_3125 (O_3125,N_49794,N_49852);
nand UO_3126 (O_3126,N_49545,N_49898);
nor UO_3127 (O_3127,N_49892,N_49533);
and UO_3128 (O_3128,N_49749,N_49916);
and UO_3129 (O_3129,N_49612,N_49557);
nor UO_3130 (O_3130,N_49531,N_49924);
nand UO_3131 (O_3131,N_49608,N_49905);
nand UO_3132 (O_3132,N_49737,N_49865);
xnor UO_3133 (O_3133,N_49646,N_49821);
nand UO_3134 (O_3134,N_49818,N_49611);
nand UO_3135 (O_3135,N_49534,N_49608);
and UO_3136 (O_3136,N_49625,N_49619);
xnor UO_3137 (O_3137,N_49698,N_49946);
and UO_3138 (O_3138,N_49662,N_49736);
nand UO_3139 (O_3139,N_49654,N_49911);
or UO_3140 (O_3140,N_49560,N_49960);
xor UO_3141 (O_3141,N_49927,N_49612);
xor UO_3142 (O_3142,N_49718,N_49976);
nand UO_3143 (O_3143,N_49692,N_49518);
xor UO_3144 (O_3144,N_49932,N_49997);
nand UO_3145 (O_3145,N_49782,N_49805);
and UO_3146 (O_3146,N_49703,N_49534);
or UO_3147 (O_3147,N_49829,N_49599);
and UO_3148 (O_3148,N_49568,N_49645);
nor UO_3149 (O_3149,N_49501,N_49857);
or UO_3150 (O_3150,N_49990,N_49648);
or UO_3151 (O_3151,N_49744,N_49535);
nor UO_3152 (O_3152,N_49932,N_49974);
xor UO_3153 (O_3153,N_49704,N_49787);
and UO_3154 (O_3154,N_49574,N_49549);
and UO_3155 (O_3155,N_49922,N_49542);
xnor UO_3156 (O_3156,N_49817,N_49668);
nand UO_3157 (O_3157,N_49745,N_49631);
nand UO_3158 (O_3158,N_49884,N_49711);
or UO_3159 (O_3159,N_49760,N_49756);
or UO_3160 (O_3160,N_49879,N_49566);
xnor UO_3161 (O_3161,N_49720,N_49740);
nor UO_3162 (O_3162,N_49704,N_49680);
and UO_3163 (O_3163,N_49799,N_49507);
nand UO_3164 (O_3164,N_49824,N_49840);
nand UO_3165 (O_3165,N_49970,N_49968);
nor UO_3166 (O_3166,N_49964,N_49750);
xnor UO_3167 (O_3167,N_49742,N_49740);
nand UO_3168 (O_3168,N_49664,N_49670);
or UO_3169 (O_3169,N_49601,N_49674);
or UO_3170 (O_3170,N_49905,N_49740);
xor UO_3171 (O_3171,N_49708,N_49656);
nand UO_3172 (O_3172,N_49865,N_49990);
nor UO_3173 (O_3173,N_49509,N_49813);
and UO_3174 (O_3174,N_49688,N_49963);
nand UO_3175 (O_3175,N_49723,N_49980);
and UO_3176 (O_3176,N_49819,N_49609);
or UO_3177 (O_3177,N_49995,N_49909);
nand UO_3178 (O_3178,N_49844,N_49663);
nor UO_3179 (O_3179,N_49821,N_49718);
xor UO_3180 (O_3180,N_49743,N_49899);
nand UO_3181 (O_3181,N_49840,N_49506);
nand UO_3182 (O_3182,N_49707,N_49921);
nand UO_3183 (O_3183,N_49726,N_49982);
or UO_3184 (O_3184,N_49707,N_49549);
xnor UO_3185 (O_3185,N_49840,N_49797);
nor UO_3186 (O_3186,N_49778,N_49970);
nand UO_3187 (O_3187,N_49957,N_49681);
nand UO_3188 (O_3188,N_49854,N_49975);
nand UO_3189 (O_3189,N_49813,N_49698);
nor UO_3190 (O_3190,N_49998,N_49801);
nor UO_3191 (O_3191,N_49605,N_49704);
nor UO_3192 (O_3192,N_49790,N_49949);
xnor UO_3193 (O_3193,N_49624,N_49917);
xnor UO_3194 (O_3194,N_49917,N_49724);
and UO_3195 (O_3195,N_49786,N_49621);
nor UO_3196 (O_3196,N_49975,N_49750);
nor UO_3197 (O_3197,N_49974,N_49694);
and UO_3198 (O_3198,N_49844,N_49878);
nand UO_3199 (O_3199,N_49893,N_49599);
or UO_3200 (O_3200,N_49626,N_49695);
nor UO_3201 (O_3201,N_49759,N_49773);
or UO_3202 (O_3202,N_49695,N_49837);
xor UO_3203 (O_3203,N_49977,N_49542);
nand UO_3204 (O_3204,N_49529,N_49618);
xor UO_3205 (O_3205,N_49661,N_49731);
or UO_3206 (O_3206,N_49908,N_49621);
nand UO_3207 (O_3207,N_49824,N_49695);
and UO_3208 (O_3208,N_49921,N_49692);
nand UO_3209 (O_3209,N_49663,N_49930);
or UO_3210 (O_3210,N_49693,N_49924);
and UO_3211 (O_3211,N_49615,N_49760);
xor UO_3212 (O_3212,N_49562,N_49918);
nand UO_3213 (O_3213,N_49826,N_49782);
and UO_3214 (O_3214,N_49562,N_49889);
or UO_3215 (O_3215,N_49760,N_49701);
and UO_3216 (O_3216,N_49757,N_49825);
nand UO_3217 (O_3217,N_49702,N_49830);
and UO_3218 (O_3218,N_49531,N_49576);
and UO_3219 (O_3219,N_49805,N_49799);
nor UO_3220 (O_3220,N_49918,N_49865);
xnor UO_3221 (O_3221,N_49890,N_49734);
nand UO_3222 (O_3222,N_49899,N_49794);
xnor UO_3223 (O_3223,N_49936,N_49737);
or UO_3224 (O_3224,N_49863,N_49620);
and UO_3225 (O_3225,N_49771,N_49886);
and UO_3226 (O_3226,N_49689,N_49948);
nand UO_3227 (O_3227,N_49917,N_49903);
xnor UO_3228 (O_3228,N_49848,N_49806);
nand UO_3229 (O_3229,N_49891,N_49799);
xor UO_3230 (O_3230,N_49795,N_49925);
and UO_3231 (O_3231,N_49537,N_49613);
and UO_3232 (O_3232,N_49849,N_49612);
and UO_3233 (O_3233,N_49561,N_49577);
or UO_3234 (O_3234,N_49620,N_49891);
and UO_3235 (O_3235,N_49927,N_49759);
nor UO_3236 (O_3236,N_49702,N_49801);
and UO_3237 (O_3237,N_49958,N_49950);
or UO_3238 (O_3238,N_49992,N_49553);
and UO_3239 (O_3239,N_49500,N_49625);
or UO_3240 (O_3240,N_49956,N_49556);
or UO_3241 (O_3241,N_49783,N_49604);
and UO_3242 (O_3242,N_49525,N_49938);
xor UO_3243 (O_3243,N_49717,N_49514);
nor UO_3244 (O_3244,N_49770,N_49768);
xnor UO_3245 (O_3245,N_49726,N_49545);
nand UO_3246 (O_3246,N_49737,N_49503);
or UO_3247 (O_3247,N_49699,N_49641);
or UO_3248 (O_3248,N_49840,N_49581);
or UO_3249 (O_3249,N_49721,N_49670);
xnor UO_3250 (O_3250,N_49984,N_49537);
and UO_3251 (O_3251,N_49695,N_49576);
or UO_3252 (O_3252,N_49536,N_49754);
nor UO_3253 (O_3253,N_49855,N_49736);
and UO_3254 (O_3254,N_49981,N_49516);
nand UO_3255 (O_3255,N_49871,N_49517);
xnor UO_3256 (O_3256,N_49878,N_49519);
xnor UO_3257 (O_3257,N_49536,N_49636);
nor UO_3258 (O_3258,N_49828,N_49784);
or UO_3259 (O_3259,N_49925,N_49691);
nand UO_3260 (O_3260,N_49907,N_49883);
nor UO_3261 (O_3261,N_49860,N_49837);
nor UO_3262 (O_3262,N_49896,N_49912);
and UO_3263 (O_3263,N_49645,N_49960);
nor UO_3264 (O_3264,N_49795,N_49857);
nand UO_3265 (O_3265,N_49621,N_49704);
nor UO_3266 (O_3266,N_49837,N_49835);
xor UO_3267 (O_3267,N_49527,N_49702);
or UO_3268 (O_3268,N_49601,N_49781);
xnor UO_3269 (O_3269,N_49547,N_49567);
or UO_3270 (O_3270,N_49967,N_49586);
nor UO_3271 (O_3271,N_49960,N_49901);
and UO_3272 (O_3272,N_49771,N_49669);
nor UO_3273 (O_3273,N_49945,N_49709);
and UO_3274 (O_3274,N_49554,N_49544);
and UO_3275 (O_3275,N_49702,N_49875);
nand UO_3276 (O_3276,N_49628,N_49873);
and UO_3277 (O_3277,N_49875,N_49855);
nor UO_3278 (O_3278,N_49645,N_49823);
or UO_3279 (O_3279,N_49923,N_49675);
nand UO_3280 (O_3280,N_49898,N_49783);
or UO_3281 (O_3281,N_49906,N_49802);
nand UO_3282 (O_3282,N_49897,N_49940);
xnor UO_3283 (O_3283,N_49849,N_49990);
xor UO_3284 (O_3284,N_49807,N_49782);
xor UO_3285 (O_3285,N_49798,N_49925);
and UO_3286 (O_3286,N_49797,N_49846);
nand UO_3287 (O_3287,N_49696,N_49999);
nand UO_3288 (O_3288,N_49665,N_49813);
nor UO_3289 (O_3289,N_49905,N_49668);
or UO_3290 (O_3290,N_49880,N_49646);
nor UO_3291 (O_3291,N_49561,N_49759);
or UO_3292 (O_3292,N_49694,N_49602);
nor UO_3293 (O_3293,N_49792,N_49604);
nand UO_3294 (O_3294,N_49845,N_49554);
xor UO_3295 (O_3295,N_49734,N_49900);
xnor UO_3296 (O_3296,N_49714,N_49727);
xor UO_3297 (O_3297,N_49849,N_49890);
and UO_3298 (O_3298,N_49837,N_49895);
xor UO_3299 (O_3299,N_49994,N_49562);
nand UO_3300 (O_3300,N_49650,N_49889);
and UO_3301 (O_3301,N_49609,N_49734);
and UO_3302 (O_3302,N_49731,N_49569);
and UO_3303 (O_3303,N_49524,N_49612);
nor UO_3304 (O_3304,N_49592,N_49953);
xor UO_3305 (O_3305,N_49780,N_49513);
or UO_3306 (O_3306,N_49648,N_49570);
nor UO_3307 (O_3307,N_49854,N_49516);
xnor UO_3308 (O_3308,N_49885,N_49662);
nor UO_3309 (O_3309,N_49669,N_49901);
xnor UO_3310 (O_3310,N_49578,N_49987);
xor UO_3311 (O_3311,N_49714,N_49512);
xor UO_3312 (O_3312,N_49559,N_49949);
nor UO_3313 (O_3313,N_49682,N_49561);
nor UO_3314 (O_3314,N_49812,N_49950);
and UO_3315 (O_3315,N_49937,N_49841);
nand UO_3316 (O_3316,N_49821,N_49651);
nor UO_3317 (O_3317,N_49775,N_49784);
and UO_3318 (O_3318,N_49545,N_49848);
xor UO_3319 (O_3319,N_49664,N_49646);
or UO_3320 (O_3320,N_49827,N_49647);
nand UO_3321 (O_3321,N_49825,N_49997);
or UO_3322 (O_3322,N_49540,N_49767);
xor UO_3323 (O_3323,N_49855,N_49936);
nor UO_3324 (O_3324,N_49523,N_49630);
xnor UO_3325 (O_3325,N_49879,N_49514);
and UO_3326 (O_3326,N_49518,N_49902);
and UO_3327 (O_3327,N_49761,N_49546);
xnor UO_3328 (O_3328,N_49961,N_49763);
nor UO_3329 (O_3329,N_49666,N_49561);
nor UO_3330 (O_3330,N_49714,N_49738);
or UO_3331 (O_3331,N_49786,N_49974);
xor UO_3332 (O_3332,N_49791,N_49708);
nand UO_3333 (O_3333,N_49938,N_49503);
xor UO_3334 (O_3334,N_49803,N_49547);
or UO_3335 (O_3335,N_49526,N_49846);
nor UO_3336 (O_3336,N_49838,N_49647);
nor UO_3337 (O_3337,N_49855,N_49845);
and UO_3338 (O_3338,N_49577,N_49528);
nand UO_3339 (O_3339,N_49630,N_49647);
or UO_3340 (O_3340,N_49573,N_49600);
nand UO_3341 (O_3341,N_49745,N_49895);
nor UO_3342 (O_3342,N_49830,N_49952);
or UO_3343 (O_3343,N_49895,N_49749);
xor UO_3344 (O_3344,N_49533,N_49608);
and UO_3345 (O_3345,N_49863,N_49581);
or UO_3346 (O_3346,N_49738,N_49577);
xnor UO_3347 (O_3347,N_49586,N_49868);
xnor UO_3348 (O_3348,N_49532,N_49628);
nor UO_3349 (O_3349,N_49597,N_49796);
nor UO_3350 (O_3350,N_49507,N_49867);
nand UO_3351 (O_3351,N_49848,N_49689);
xnor UO_3352 (O_3352,N_49543,N_49719);
nor UO_3353 (O_3353,N_49785,N_49504);
xnor UO_3354 (O_3354,N_49771,N_49727);
or UO_3355 (O_3355,N_49616,N_49849);
and UO_3356 (O_3356,N_49734,N_49893);
xor UO_3357 (O_3357,N_49845,N_49820);
or UO_3358 (O_3358,N_49997,N_49579);
nand UO_3359 (O_3359,N_49862,N_49892);
xnor UO_3360 (O_3360,N_49974,N_49591);
xor UO_3361 (O_3361,N_49746,N_49719);
or UO_3362 (O_3362,N_49784,N_49588);
nand UO_3363 (O_3363,N_49898,N_49887);
and UO_3364 (O_3364,N_49671,N_49853);
nor UO_3365 (O_3365,N_49741,N_49678);
nor UO_3366 (O_3366,N_49982,N_49861);
xor UO_3367 (O_3367,N_49786,N_49501);
nand UO_3368 (O_3368,N_49659,N_49904);
xnor UO_3369 (O_3369,N_49735,N_49610);
or UO_3370 (O_3370,N_49857,N_49557);
xnor UO_3371 (O_3371,N_49686,N_49589);
xnor UO_3372 (O_3372,N_49710,N_49773);
nand UO_3373 (O_3373,N_49955,N_49502);
or UO_3374 (O_3374,N_49657,N_49925);
or UO_3375 (O_3375,N_49819,N_49855);
nor UO_3376 (O_3376,N_49759,N_49666);
xor UO_3377 (O_3377,N_49671,N_49829);
nor UO_3378 (O_3378,N_49908,N_49600);
xnor UO_3379 (O_3379,N_49864,N_49513);
xnor UO_3380 (O_3380,N_49950,N_49596);
or UO_3381 (O_3381,N_49513,N_49598);
xor UO_3382 (O_3382,N_49586,N_49519);
xnor UO_3383 (O_3383,N_49713,N_49979);
nand UO_3384 (O_3384,N_49717,N_49554);
nand UO_3385 (O_3385,N_49892,N_49751);
and UO_3386 (O_3386,N_49565,N_49679);
xor UO_3387 (O_3387,N_49897,N_49709);
xnor UO_3388 (O_3388,N_49860,N_49520);
nor UO_3389 (O_3389,N_49523,N_49969);
or UO_3390 (O_3390,N_49925,N_49684);
xnor UO_3391 (O_3391,N_49667,N_49762);
xor UO_3392 (O_3392,N_49655,N_49590);
nor UO_3393 (O_3393,N_49654,N_49625);
xnor UO_3394 (O_3394,N_49609,N_49809);
and UO_3395 (O_3395,N_49801,N_49942);
and UO_3396 (O_3396,N_49672,N_49524);
or UO_3397 (O_3397,N_49649,N_49525);
nor UO_3398 (O_3398,N_49589,N_49748);
or UO_3399 (O_3399,N_49965,N_49692);
or UO_3400 (O_3400,N_49957,N_49740);
or UO_3401 (O_3401,N_49814,N_49983);
and UO_3402 (O_3402,N_49741,N_49835);
xnor UO_3403 (O_3403,N_49514,N_49525);
and UO_3404 (O_3404,N_49627,N_49602);
nand UO_3405 (O_3405,N_49578,N_49941);
and UO_3406 (O_3406,N_49950,N_49601);
and UO_3407 (O_3407,N_49896,N_49812);
xnor UO_3408 (O_3408,N_49656,N_49943);
xor UO_3409 (O_3409,N_49704,N_49700);
nand UO_3410 (O_3410,N_49673,N_49866);
nor UO_3411 (O_3411,N_49890,N_49549);
xor UO_3412 (O_3412,N_49767,N_49898);
xnor UO_3413 (O_3413,N_49953,N_49548);
or UO_3414 (O_3414,N_49760,N_49923);
nand UO_3415 (O_3415,N_49562,N_49715);
nor UO_3416 (O_3416,N_49586,N_49994);
nor UO_3417 (O_3417,N_49743,N_49742);
and UO_3418 (O_3418,N_49962,N_49575);
and UO_3419 (O_3419,N_49827,N_49792);
and UO_3420 (O_3420,N_49573,N_49788);
nor UO_3421 (O_3421,N_49892,N_49746);
or UO_3422 (O_3422,N_49893,N_49918);
or UO_3423 (O_3423,N_49769,N_49678);
xnor UO_3424 (O_3424,N_49652,N_49777);
nor UO_3425 (O_3425,N_49835,N_49645);
or UO_3426 (O_3426,N_49564,N_49833);
nand UO_3427 (O_3427,N_49880,N_49522);
nor UO_3428 (O_3428,N_49715,N_49759);
or UO_3429 (O_3429,N_49959,N_49508);
xnor UO_3430 (O_3430,N_49515,N_49989);
or UO_3431 (O_3431,N_49523,N_49748);
xor UO_3432 (O_3432,N_49969,N_49563);
or UO_3433 (O_3433,N_49969,N_49825);
xor UO_3434 (O_3434,N_49655,N_49724);
and UO_3435 (O_3435,N_49563,N_49505);
and UO_3436 (O_3436,N_49727,N_49594);
nand UO_3437 (O_3437,N_49718,N_49719);
nand UO_3438 (O_3438,N_49763,N_49789);
nand UO_3439 (O_3439,N_49955,N_49743);
xor UO_3440 (O_3440,N_49664,N_49590);
nand UO_3441 (O_3441,N_49858,N_49811);
nor UO_3442 (O_3442,N_49870,N_49875);
xnor UO_3443 (O_3443,N_49503,N_49752);
nand UO_3444 (O_3444,N_49768,N_49804);
nand UO_3445 (O_3445,N_49558,N_49795);
or UO_3446 (O_3446,N_49931,N_49644);
nand UO_3447 (O_3447,N_49983,N_49523);
or UO_3448 (O_3448,N_49911,N_49611);
nor UO_3449 (O_3449,N_49562,N_49671);
xnor UO_3450 (O_3450,N_49955,N_49834);
nor UO_3451 (O_3451,N_49987,N_49886);
nand UO_3452 (O_3452,N_49567,N_49597);
xnor UO_3453 (O_3453,N_49670,N_49983);
or UO_3454 (O_3454,N_49627,N_49703);
nand UO_3455 (O_3455,N_49522,N_49800);
or UO_3456 (O_3456,N_49939,N_49935);
and UO_3457 (O_3457,N_49545,N_49716);
xnor UO_3458 (O_3458,N_49874,N_49962);
xor UO_3459 (O_3459,N_49886,N_49768);
xnor UO_3460 (O_3460,N_49978,N_49895);
and UO_3461 (O_3461,N_49882,N_49894);
nor UO_3462 (O_3462,N_49689,N_49746);
nor UO_3463 (O_3463,N_49814,N_49899);
nor UO_3464 (O_3464,N_49696,N_49615);
nand UO_3465 (O_3465,N_49736,N_49804);
nor UO_3466 (O_3466,N_49608,N_49862);
xnor UO_3467 (O_3467,N_49544,N_49829);
and UO_3468 (O_3468,N_49997,N_49792);
xor UO_3469 (O_3469,N_49928,N_49890);
and UO_3470 (O_3470,N_49903,N_49962);
xor UO_3471 (O_3471,N_49719,N_49585);
xor UO_3472 (O_3472,N_49690,N_49616);
and UO_3473 (O_3473,N_49506,N_49559);
nand UO_3474 (O_3474,N_49790,N_49999);
and UO_3475 (O_3475,N_49966,N_49875);
xor UO_3476 (O_3476,N_49810,N_49743);
or UO_3477 (O_3477,N_49671,N_49726);
xor UO_3478 (O_3478,N_49769,N_49723);
and UO_3479 (O_3479,N_49631,N_49717);
xor UO_3480 (O_3480,N_49790,N_49948);
nand UO_3481 (O_3481,N_49505,N_49924);
xnor UO_3482 (O_3482,N_49500,N_49775);
nand UO_3483 (O_3483,N_49829,N_49970);
xnor UO_3484 (O_3484,N_49758,N_49548);
nand UO_3485 (O_3485,N_49718,N_49684);
and UO_3486 (O_3486,N_49791,N_49637);
and UO_3487 (O_3487,N_49669,N_49810);
xor UO_3488 (O_3488,N_49579,N_49749);
and UO_3489 (O_3489,N_49911,N_49623);
nand UO_3490 (O_3490,N_49765,N_49679);
nor UO_3491 (O_3491,N_49929,N_49759);
xnor UO_3492 (O_3492,N_49623,N_49798);
nor UO_3493 (O_3493,N_49580,N_49682);
and UO_3494 (O_3494,N_49920,N_49896);
nand UO_3495 (O_3495,N_49504,N_49519);
xor UO_3496 (O_3496,N_49793,N_49938);
nor UO_3497 (O_3497,N_49891,N_49674);
nor UO_3498 (O_3498,N_49917,N_49825);
xnor UO_3499 (O_3499,N_49511,N_49541);
nor UO_3500 (O_3500,N_49926,N_49706);
nor UO_3501 (O_3501,N_49506,N_49844);
xnor UO_3502 (O_3502,N_49971,N_49858);
xor UO_3503 (O_3503,N_49656,N_49598);
nand UO_3504 (O_3504,N_49881,N_49570);
and UO_3505 (O_3505,N_49946,N_49965);
nor UO_3506 (O_3506,N_49594,N_49672);
and UO_3507 (O_3507,N_49741,N_49593);
xor UO_3508 (O_3508,N_49575,N_49859);
nand UO_3509 (O_3509,N_49928,N_49512);
and UO_3510 (O_3510,N_49680,N_49942);
xnor UO_3511 (O_3511,N_49966,N_49803);
xnor UO_3512 (O_3512,N_49561,N_49985);
xnor UO_3513 (O_3513,N_49736,N_49906);
nor UO_3514 (O_3514,N_49536,N_49794);
nor UO_3515 (O_3515,N_49595,N_49645);
nor UO_3516 (O_3516,N_49906,N_49850);
or UO_3517 (O_3517,N_49725,N_49724);
nor UO_3518 (O_3518,N_49787,N_49630);
nor UO_3519 (O_3519,N_49591,N_49737);
and UO_3520 (O_3520,N_49615,N_49774);
or UO_3521 (O_3521,N_49919,N_49559);
or UO_3522 (O_3522,N_49717,N_49680);
nand UO_3523 (O_3523,N_49628,N_49935);
nand UO_3524 (O_3524,N_49903,N_49506);
xnor UO_3525 (O_3525,N_49888,N_49960);
xor UO_3526 (O_3526,N_49974,N_49748);
xor UO_3527 (O_3527,N_49705,N_49741);
nor UO_3528 (O_3528,N_49796,N_49741);
and UO_3529 (O_3529,N_49580,N_49755);
nor UO_3530 (O_3530,N_49558,N_49698);
nor UO_3531 (O_3531,N_49507,N_49979);
xor UO_3532 (O_3532,N_49745,N_49886);
or UO_3533 (O_3533,N_49994,N_49569);
nand UO_3534 (O_3534,N_49871,N_49798);
nand UO_3535 (O_3535,N_49676,N_49883);
and UO_3536 (O_3536,N_49935,N_49850);
nand UO_3537 (O_3537,N_49837,N_49596);
and UO_3538 (O_3538,N_49933,N_49940);
nor UO_3539 (O_3539,N_49808,N_49954);
nand UO_3540 (O_3540,N_49988,N_49811);
or UO_3541 (O_3541,N_49940,N_49553);
or UO_3542 (O_3542,N_49624,N_49637);
and UO_3543 (O_3543,N_49939,N_49776);
nor UO_3544 (O_3544,N_49508,N_49981);
nor UO_3545 (O_3545,N_49687,N_49728);
nand UO_3546 (O_3546,N_49933,N_49815);
nor UO_3547 (O_3547,N_49536,N_49543);
or UO_3548 (O_3548,N_49631,N_49991);
nor UO_3549 (O_3549,N_49871,N_49747);
and UO_3550 (O_3550,N_49769,N_49742);
and UO_3551 (O_3551,N_49886,N_49889);
xor UO_3552 (O_3552,N_49620,N_49649);
and UO_3553 (O_3553,N_49811,N_49893);
nand UO_3554 (O_3554,N_49770,N_49624);
or UO_3555 (O_3555,N_49878,N_49688);
xnor UO_3556 (O_3556,N_49643,N_49715);
nand UO_3557 (O_3557,N_49606,N_49709);
and UO_3558 (O_3558,N_49783,N_49857);
nor UO_3559 (O_3559,N_49782,N_49740);
xnor UO_3560 (O_3560,N_49617,N_49757);
nor UO_3561 (O_3561,N_49836,N_49822);
or UO_3562 (O_3562,N_49775,N_49577);
xor UO_3563 (O_3563,N_49553,N_49617);
and UO_3564 (O_3564,N_49741,N_49938);
or UO_3565 (O_3565,N_49912,N_49609);
nand UO_3566 (O_3566,N_49698,N_49659);
and UO_3567 (O_3567,N_49627,N_49925);
nand UO_3568 (O_3568,N_49623,N_49949);
nand UO_3569 (O_3569,N_49648,N_49900);
xor UO_3570 (O_3570,N_49958,N_49804);
xnor UO_3571 (O_3571,N_49910,N_49693);
or UO_3572 (O_3572,N_49633,N_49646);
xnor UO_3573 (O_3573,N_49761,N_49632);
nor UO_3574 (O_3574,N_49791,N_49786);
xor UO_3575 (O_3575,N_49661,N_49568);
nor UO_3576 (O_3576,N_49534,N_49678);
xnor UO_3577 (O_3577,N_49940,N_49716);
xor UO_3578 (O_3578,N_49996,N_49700);
xor UO_3579 (O_3579,N_49910,N_49590);
xor UO_3580 (O_3580,N_49678,N_49822);
and UO_3581 (O_3581,N_49772,N_49557);
and UO_3582 (O_3582,N_49859,N_49633);
nand UO_3583 (O_3583,N_49847,N_49720);
nand UO_3584 (O_3584,N_49713,N_49504);
nand UO_3585 (O_3585,N_49591,N_49808);
or UO_3586 (O_3586,N_49905,N_49816);
and UO_3587 (O_3587,N_49765,N_49950);
and UO_3588 (O_3588,N_49563,N_49652);
nand UO_3589 (O_3589,N_49975,N_49785);
or UO_3590 (O_3590,N_49869,N_49797);
or UO_3591 (O_3591,N_49944,N_49694);
nand UO_3592 (O_3592,N_49742,N_49595);
xnor UO_3593 (O_3593,N_49776,N_49888);
xor UO_3594 (O_3594,N_49631,N_49889);
nor UO_3595 (O_3595,N_49730,N_49571);
nand UO_3596 (O_3596,N_49571,N_49659);
and UO_3597 (O_3597,N_49845,N_49764);
nand UO_3598 (O_3598,N_49711,N_49926);
xnor UO_3599 (O_3599,N_49625,N_49754);
and UO_3600 (O_3600,N_49583,N_49738);
nor UO_3601 (O_3601,N_49911,N_49592);
xor UO_3602 (O_3602,N_49511,N_49946);
xnor UO_3603 (O_3603,N_49848,N_49900);
nor UO_3604 (O_3604,N_49841,N_49855);
or UO_3605 (O_3605,N_49719,N_49978);
and UO_3606 (O_3606,N_49901,N_49718);
xnor UO_3607 (O_3607,N_49741,N_49980);
nand UO_3608 (O_3608,N_49812,N_49632);
xnor UO_3609 (O_3609,N_49827,N_49836);
nor UO_3610 (O_3610,N_49560,N_49954);
or UO_3611 (O_3611,N_49913,N_49710);
nor UO_3612 (O_3612,N_49566,N_49838);
nor UO_3613 (O_3613,N_49587,N_49956);
nand UO_3614 (O_3614,N_49676,N_49613);
and UO_3615 (O_3615,N_49900,N_49507);
and UO_3616 (O_3616,N_49882,N_49706);
or UO_3617 (O_3617,N_49574,N_49885);
or UO_3618 (O_3618,N_49997,N_49782);
nand UO_3619 (O_3619,N_49752,N_49509);
or UO_3620 (O_3620,N_49538,N_49657);
xor UO_3621 (O_3621,N_49923,N_49528);
nand UO_3622 (O_3622,N_49589,N_49767);
xnor UO_3623 (O_3623,N_49674,N_49824);
nor UO_3624 (O_3624,N_49789,N_49538);
nand UO_3625 (O_3625,N_49811,N_49673);
or UO_3626 (O_3626,N_49870,N_49642);
nor UO_3627 (O_3627,N_49902,N_49708);
nand UO_3628 (O_3628,N_49597,N_49754);
xor UO_3629 (O_3629,N_49617,N_49515);
and UO_3630 (O_3630,N_49712,N_49555);
and UO_3631 (O_3631,N_49792,N_49797);
xnor UO_3632 (O_3632,N_49610,N_49999);
nor UO_3633 (O_3633,N_49551,N_49548);
or UO_3634 (O_3634,N_49622,N_49870);
and UO_3635 (O_3635,N_49728,N_49865);
xor UO_3636 (O_3636,N_49544,N_49640);
or UO_3637 (O_3637,N_49969,N_49763);
and UO_3638 (O_3638,N_49811,N_49892);
or UO_3639 (O_3639,N_49923,N_49783);
and UO_3640 (O_3640,N_49637,N_49886);
nand UO_3641 (O_3641,N_49995,N_49998);
or UO_3642 (O_3642,N_49694,N_49901);
nand UO_3643 (O_3643,N_49608,N_49536);
xnor UO_3644 (O_3644,N_49615,N_49565);
nand UO_3645 (O_3645,N_49573,N_49807);
and UO_3646 (O_3646,N_49544,N_49999);
and UO_3647 (O_3647,N_49701,N_49915);
nand UO_3648 (O_3648,N_49990,N_49595);
nor UO_3649 (O_3649,N_49501,N_49570);
xnor UO_3650 (O_3650,N_49549,N_49606);
xor UO_3651 (O_3651,N_49879,N_49972);
nor UO_3652 (O_3652,N_49921,N_49937);
and UO_3653 (O_3653,N_49548,N_49860);
or UO_3654 (O_3654,N_49530,N_49635);
and UO_3655 (O_3655,N_49542,N_49990);
nor UO_3656 (O_3656,N_49793,N_49698);
and UO_3657 (O_3657,N_49703,N_49805);
nor UO_3658 (O_3658,N_49682,N_49759);
xor UO_3659 (O_3659,N_49845,N_49589);
nand UO_3660 (O_3660,N_49522,N_49951);
and UO_3661 (O_3661,N_49950,N_49624);
nand UO_3662 (O_3662,N_49828,N_49593);
or UO_3663 (O_3663,N_49843,N_49587);
nor UO_3664 (O_3664,N_49925,N_49705);
nand UO_3665 (O_3665,N_49757,N_49813);
nand UO_3666 (O_3666,N_49741,N_49841);
and UO_3667 (O_3667,N_49986,N_49787);
xnor UO_3668 (O_3668,N_49865,N_49511);
nor UO_3669 (O_3669,N_49727,N_49853);
nor UO_3670 (O_3670,N_49623,N_49823);
nor UO_3671 (O_3671,N_49551,N_49614);
nor UO_3672 (O_3672,N_49610,N_49720);
nor UO_3673 (O_3673,N_49865,N_49980);
nand UO_3674 (O_3674,N_49668,N_49601);
or UO_3675 (O_3675,N_49532,N_49889);
xnor UO_3676 (O_3676,N_49512,N_49582);
nand UO_3677 (O_3677,N_49653,N_49903);
or UO_3678 (O_3678,N_49963,N_49857);
or UO_3679 (O_3679,N_49604,N_49612);
nand UO_3680 (O_3680,N_49623,N_49544);
nor UO_3681 (O_3681,N_49935,N_49691);
nand UO_3682 (O_3682,N_49711,N_49832);
nor UO_3683 (O_3683,N_49525,N_49721);
nand UO_3684 (O_3684,N_49928,N_49508);
and UO_3685 (O_3685,N_49972,N_49827);
xnor UO_3686 (O_3686,N_49846,N_49586);
or UO_3687 (O_3687,N_49893,N_49822);
or UO_3688 (O_3688,N_49817,N_49847);
xnor UO_3689 (O_3689,N_49716,N_49926);
or UO_3690 (O_3690,N_49696,N_49873);
nand UO_3691 (O_3691,N_49560,N_49952);
or UO_3692 (O_3692,N_49940,N_49850);
or UO_3693 (O_3693,N_49841,N_49574);
nor UO_3694 (O_3694,N_49852,N_49536);
nor UO_3695 (O_3695,N_49804,N_49996);
nand UO_3696 (O_3696,N_49861,N_49587);
or UO_3697 (O_3697,N_49706,N_49502);
nor UO_3698 (O_3698,N_49710,N_49791);
and UO_3699 (O_3699,N_49567,N_49619);
and UO_3700 (O_3700,N_49679,N_49668);
or UO_3701 (O_3701,N_49846,N_49612);
and UO_3702 (O_3702,N_49900,N_49638);
nor UO_3703 (O_3703,N_49918,N_49871);
nor UO_3704 (O_3704,N_49956,N_49926);
and UO_3705 (O_3705,N_49876,N_49814);
xor UO_3706 (O_3706,N_49516,N_49935);
nand UO_3707 (O_3707,N_49552,N_49937);
xnor UO_3708 (O_3708,N_49909,N_49808);
or UO_3709 (O_3709,N_49752,N_49793);
and UO_3710 (O_3710,N_49939,N_49692);
xor UO_3711 (O_3711,N_49790,N_49881);
or UO_3712 (O_3712,N_49859,N_49747);
or UO_3713 (O_3713,N_49996,N_49903);
xnor UO_3714 (O_3714,N_49691,N_49633);
nor UO_3715 (O_3715,N_49973,N_49936);
or UO_3716 (O_3716,N_49717,N_49612);
nor UO_3717 (O_3717,N_49689,N_49903);
or UO_3718 (O_3718,N_49512,N_49759);
and UO_3719 (O_3719,N_49811,N_49696);
nor UO_3720 (O_3720,N_49685,N_49857);
xor UO_3721 (O_3721,N_49602,N_49636);
or UO_3722 (O_3722,N_49568,N_49639);
nor UO_3723 (O_3723,N_49731,N_49746);
and UO_3724 (O_3724,N_49514,N_49598);
or UO_3725 (O_3725,N_49833,N_49781);
nand UO_3726 (O_3726,N_49825,N_49852);
xnor UO_3727 (O_3727,N_49537,N_49739);
xnor UO_3728 (O_3728,N_49706,N_49555);
xor UO_3729 (O_3729,N_49548,N_49948);
and UO_3730 (O_3730,N_49719,N_49517);
and UO_3731 (O_3731,N_49600,N_49502);
xnor UO_3732 (O_3732,N_49641,N_49926);
xor UO_3733 (O_3733,N_49995,N_49936);
and UO_3734 (O_3734,N_49681,N_49835);
nor UO_3735 (O_3735,N_49537,N_49548);
nand UO_3736 (O_3736,N_49885,N_49529);
nand UO_3737 (O_3737,N_49778,N_49745);
xor UO_3738 (O_3738,N_49953,N_49968);
nand UO_3739 (O_3739,N_49651,N_49634);
or UO_3740 (O_3740,N_49983,N_49922);
or UO_3741 (O_3741,N_49627,N_49577);
xor UO_3742 (O_3742,N_49758,N_49819);
or UO_3743 (O_3743,N_49727,N_49780);
nand UO_3744 (O_3744,N_49512,N_49563);
or UO_3745 (O_3745,N_49841,N_49902);
xnor UO_3746 (O_3746,N_49716,N_49646);
nand UO_3747 (O_3747,N_49712,N_49997);
nor UO_3748 (O_3748,N_49767,N_49965);
nand UO_3749 (O_3749,N_49881,N_49808);
nor UO_3750 (O_3750,N_49607,N_49873);
or UO_3751 (O_3751,N_49793,N_49973);
and UO_3752 (O_3752,N_49846,N_49899);
nor UO_3753 (O_3753,N_49951,N_49567);
nor UO_3754 (O_3754,N_49860,N_49755);
nand UO_3755 (O_3755,N_49899,N_49811);
nor UO_3756 (O_3756,N_49603,N_49898);
nor UO_3757 (O_3757,N_49743,N_49541);
nand UO_3758 (O_3758,N_49602,N_49625);
nand UO_3759 (O_3759,N_49572,N_49961);
nor UO_3760 (O_3760,N_49785,N_49657);
nand UO_3761 (O_3761,N_49596,N_49514);
xnor UO_3762 (O_3762,N_49881,N_49898);
or UO_3763 (O_3763,N_49782,N_49839);
nor UO_3764 (O_3764,N_49661,N_49611);
or UO_3765 (O_3765,N_49561,N_49946);
xor UO_3766 (O_3766,N_49546,N_49756);
and UO_3767 (O_3767,N_49997,N_49743);
xor UO_3768 (O_3768,N_49631,N_49561);
and UO_3769 (O_3769,N_49892,N_49879);
nor UO_3770 (O_3770,N_49950,N_49994);
nand UO_3771 (O_3771,N_49787,N_49912);
or UO_3772 (O_3772,N_49941,N_49958);
and UO_3773 (O_3773,N_49881,N_49912);
or UO_3774 (O_3774,N_49910,N_49620);
nor UO_3775 (O_3775,N_49666,N_49589);
nor UO_3776 (O_3776,N_49684,N_49983);
and UO_3777 (O_3777,N_49979,N_49592);
nor UO_3778 (O_3778,N_49871,N_49717);
nand UO_3779 (O_3779,N_49935,N_49868);
nand UO_3780 (O_3780,N_49594,N_49563);
or UO_3781 (O_3781,N_49841,N_49786);
nor UO_3782 (O_3782,N_49749,N_49668);
xor UO_3783 (O_3783,N_49867,N_49586);
xnor UO_3784 (O_3784,N_49894,N_49519);
xnor UO_3785 (O_3785,N_49697,N_49777);
xnor UO_3786 (O_3786,N_49863,N_49837);
and UO_3787 (O_3787,N_49952,N_49511);
xnor UO_3788 (O_3788,N_49644,N_49717);
nor UO_3789 (O_3789,N_49793,N_49943);
xnor UO_3790 (O_3790,N_49670,N_49779);
or UO_3791 (O_3791,N_49992,N_49619);
nand UO_3792 (O_3792,N_49525,N_49537);
nand UO_3793 (O_3793,N_49722,N_49975);
xnor UO_3794 (O_3794,N_49630,N_49741);
nand UO_3795 (O_3795,N_49709,N_49744);
and UO_3796 (O_3796,N_49573,N_49612);
nand UO_3797 (O_3797,N_49556,N_49899);
or UO_3798 (O_3798,N_49502,N_49987);
nand UO_3799 (O_3799,N_49963,N_49602);
xnor UO_3800 (O_3800,N_49821,N_49738);
and UO_3801 (O_3801,N_49618,N_49560);
nand UO_3802 (O_3802,N_49631,N_49681);
or UO_3803 (O_3803,N_49975,N_49742);
nor UO_3804 (O_3804,N_49667,N_49518);
xnor UO_3805 (O_3805,N_49654,N_49647);
xor UO_3806 (O_3806,N_49646,N_49736);
nor UO_3807 (O_3807,N_49571,N_49914);
xor UO_3808 (O_3808,N_49712,N_49609);
and UO_3809 (O_3809,N_49884,N_49804);
nand UO_3810 (O_3810,N_49729,N_49547);
nand UO_3811 (O_3811,N_49901,N_49884);
nand UO_3812 (O_3812,N_49899,N_49933);
xnor UO_3813 (O_3813,N_49580,N_49953);
and UO_3814 (O_3814,N_49740,N_49532);
or UO_3815 (O_3815,N_49990,N_49593);
or UO_3816 (O_3816,N_49716,N_49865);
xor UO_3817 (O_3817,N_49953,N_49891);
and UO_3818 (O_3818,N_49623,N_49892);
or UO_3819 (O_3819,N_49508,N_49971);
nand UO_3820 (O_3820,N_49728,N_49602);
nand UO_3821 (O_3821,N_49633,N_49729);
nor UO_3822 (O_3822,N_49613,N_49519);
xor UO_3823 (O_3823,N_49951,N_49514);
or UO_3824 (O_3824,N_49698,N_49543);
or UO_3825 (O_3825,N_49989,N_49978);
xor UO_3826 (O_3826,N_49554,N_49829);
xor UO_3827 (O_3827,N_49910,N_49824);
nand UO_3828 (O_3828,N_49762,N_49942);
nand UO_3829 (O_3829,N_49669,N_49840);
or UO_3830 (O_3830,N_49541,N_49650);
nor UO_3831 (O_3831,N_49816,N_49819);
nand UO_3832 (O_3832,N_49532,N_49644);
nand UO_3833 (O_3833,N_49875,N_49534);
xor UO_3834 (O_3834,N_49510,N_49813);
and UO_3835 (O_3835,N_49565,N_49761);
xor UO_3836 (O_3836,N_49957,N_49867);
nor UO_3837 (O_3837,N_49941,N_49866);
nor UO_3838 (O_3838,N_49513,N_49741);
or UO_3839 (O_3839,N_49737,N_49738);
and UO_3840 (O_3840,N_49837,N_49932);
xnor UO_3841 (O_3841,N_49864,N_49932);
xnor UO_3842 (O_3842,N_49645,N_49634);
or UO_3843 (O_3843,N_49614,N_49649);
nor UO_3844 (O_3844,N_49705,N_49814);
and UO_3845 (O_3845,N_49628,N_49615);
or UO_3846 (O_3846,N_49851,N_49594);
nor UO_3847 (O_3847,N_49712,N_49634);
xor UO_3848 (O_3848,N_49606,N_49511);
and UO_3849 (O_3849,N_49502,N_49960);
or UO_3850 (O_3850,N_49752,N_49759);
and UO_3851 (O_3851,N_49512,N_49629);
and UO_3852 (O_3852,N_49667,N_49991);
xnor UO_3853 (O_3853,N_49718,N_49996);
nand UO_3854 (O_3854,N_49582,N_49868);
and UO_3855 (O_3855,N_49907,N_49536);
or UO_3856 (O_3856,N_49754,N_49876);
nand UO_3857 (O_3857,N_49654,N_49914);
or UO_3858 (O_3858,N_49782,N_49892);
nand UO_3859 (O_3859,N_49978,N_49757);
and UO_3860 (O_3860,N_49761,N_49928);
and UO_3861 (O_3861,N_49687,N_49512);
or UO_3862 (O_3862,N_49574,N_49586);
or UO_3863 (O_3863,N_49908,N_49660);
or UO_3864 (O_3864,N_49832,N_49757);
or UO_3865 (O_3865,N_49810,N_49848);
or UO_3866 (O_3866,N_49510,N_49829);
nand UO_3867 (O_3867,N_49993,N_49575);
nor UO_3868 (O_3868,N_49984,N_49883);
or UO_3869 (O_3869,N_49537,N_49778);
or UO_3870 (O_3870,N_49527,N_49980);
and UO_3871 (O_3871,N_49753,N_49738);
xor UO_3872 (O_3872,N_49661,N_49847);
and UO_3873 (O_3873,N_49997,N_49829);
nor UO_3874 (O_3874,N_49888,N_49531);
or UO_3875 (O_3875,N_49974,N_49942);
or UO_3876 (O_3876,N_49901,N_49985);
xnor UO_3877 (O_3877,N_49620,N_49696);
or UO_3878 (O_3878,N_49836,N_49506);
nand UO_3879 (O_3879,N_49698,N_49963);
and UO_3880 (O_3880,N_49787,N_49878);
or UO_3881 (O_3881,N_49731,N_49820);
or UO_3882 (O_3882,N_49943,N_49674);
or UO_3883 (O_3883,N_49585,N_49606);
and UO_3884 (O_3884,N_49682,N_49639);
xnor UO_3885 (O_3885,N_49963,N_49772);
xnor UO_3886 (O_3886,N_49992,N_49880);
xor UO_3887 (O_3887,N_49801,N_49953);
or UO_3888 (O_3888,N_49898,N_49637);
or UO_3889 (O_3889,N_49972,N_49775);
xor UO_3890 (O_3890,N_49956,N_49937);
or UO_3891 (O_3891,N_49630,N_49569);
nor UO_3892 (O_3892,N_49607,N_49520);
xnor UO_3893 (O_3893,N_49647,N_49589);
nor UO_3894 (O_3894,N_49581,N_49776);
nand UO_3895 (O_3895,N_49710,N_49630);
xor UO_3896 (O_3896,N_49789,N_49551);
nand UO_3897 (O_3897,N_49551,N_49823);
nand UO_3898 (O_3898,N_49674,N_49507);
nand UO_3899 (O_3899,N_49717,N_49846);
xnor UO_3900 (O_3900,N_49735,N_49867);
nand UO_3901 (O_3901,N_49518,N_49651);
xor UO_3902 (O_3902,N_49957,N_49694);
and UO_3903 (O_3903,N_49642,N_49614);
nor UO_3904 (O_3904,N_49715,N_49688);
or UO_3905 (O_3905,N_49823,N_49784);
nand UO_3906 (O_3906,N_49795,N_49534);
or UO_3907 (O_3907,N_49535,N_49644);
xor UO_3908 (O_3908,N_49970,N_49898);
or UO_3909 (O_3909,N_49608,N_49587);
and UO_3910 (O_3910,N_49697,N_49567);
or UO_3911 (O_3911,N_49757,N_49684);
and UO_3912 (O_3912,N_49824,N_49942);
xor UO_3913 (O_3913,N_49542,N_49938);
and UO_3914 (O_3914,N_49820,N_49957);
nor UO_3915 (O_3915,N_49996,N_49831);
nand UO_3916 (O_3916,N_49783,N_49622);
or UO_3917 (O_3917,N_49587,N_49622);
nor UO_3918 (O_3918,N_49869,N_49574);
nand UO_3919 (O_3919,N_49876,N_49902);
or UO_3920 (O_3920,N_49701,N_49777);
or UO_3921 (O_3921,N_49866,N_49817);
nand UO_3922 (O_3922,N_49673,N_49718);
xnor UO_3923 (O_3923,N_49752,N_49846);
or UO_3924 (O_3924,N_49765,N_49582);
and UO_3925 (O_3925,N_49797,N_49589);
xor UO_3926 (O_3926,N_49805,N_49519);
and UO_3927 (O_3927,N_49919,N_49950);
or UO_3928 (O_3928,N_49991,N_49967);
nor UO_3929 (O_3929,N_49527,N_49813);
xor UO_3930 (O_3930,N_49909,N_49658);
nor UO_3931 (O_3931,N_49692,N_49610);
nor UO_3932 (O_3932,N_49765,N_49754);
or UO_3933 (O_3933,N_49671,N_49890);
xnor UO_3934 (O_3934,N_49696,N_49865);
or UO_3935 (O_3935,N_49804,N_49844);
or UO_3936 (O_3936,N_49872,N_49891);
nor UO_3937 (O_3937,N_49592,N_49758);
xor UO_3938 (O_3938,N_49850,N_49727);
xnor UO_3939 (O_3939,N_49807,N_49651);
nor UO_3940 (O_3940,N_49661,N_49810);
nand UO_3941 (O_3941,N_49512,N_49544);
nor UO_3942 (O_3942,N_49847,N_49640);
and UO_3943 (O_3943,N_49670,N_49520);
and UO_3944 (O_3944,N_49561,N_49994);
xnor UO_3945 (O_3945,N_49789,N_49795);
xor UO_3946 (O_3946,N_49721,N_49859);
and UO_3947 (O_3947,N_49902,N_49727);
and UO_3948 (O_3948,N_49535,N_49622);
and UO_3949 (O_3949,N_49974,N_49884);
and UO_3950 (O_3950,N_49648,N_49717);
nand UO_3951 (O_3951,N_49690,N_49812);
or UO_3952 (O_3952,N_49863,N_49922);
and UO_3953 (O_3953,N_49854,N_49677);
or UO_3954 (O_3954,N_49919,N_49847);
xnor UO_3955 (O_3955,N_49631,N_49502);
xnor UO_3956 (O_3956,N_49970,N_49616);
nor UO_3957 (O_3957,N_49736,N_49865);
xnor UO_3958 (O_3958,N_49709,N_49638);
or UO_3959 (O_3959,N_49981,N_49712);
xnor UO_3960 (O_3960,N_49717,N_49746);
nor UO_3961 (O_3961,N_49907,N_49519);
nand UO_3962 (O_3962,N_49986,N_49810);
nor UO_3963 (O_3963,N_49549,N_49585);
nand UO_3964 (O_3964,N_49670,N_49639);
nor UO_3965 (O_3965,N_49751,N_49750);
or UO_3966 (O_3966,N_49825,N_49918);
xnor UO_3967 (O_3967,N_49788,N_49577);
nor UO_3968 (O_3968,N_49591,N_49593);
or UO_3969 (O_3969,N_49773,N_49547);
xor UO_3970 (O_3970,N_49929,N_49546);
nor UO_3971 (O_3971,N_49705,N_49639);
and UO_3972 (O_3972,N_49602,N_49922);
xnor UO_3973 (O_3973,N_49573,N_49562);
and UO_3974 (O_3974,N_49911,N_49691);
and UO_3975 (O_3975,N_49874,N_49928);
nor UO_3976 (O_3976,N_49586,N_49733);
or UO_3977 (O_3977,N_49506,N_49586);
nand UO_3978 (O_3978,N_49986,N_49592);
or UO_3979 (O_3979,N_49889,N_49745);
nor UO_3980 (O_3980,N_49589,N_49947);
xnor UO_3981 (O_3981,N_49894,N_49855);
nor UO_3982 (O_3982,N_49801,N_49721);
nor UO_3983 (O_3983,N_49849,N_49770);
nor UO_3984 (O_3984,N_49556,N_49941);
nor UO_3985 (O_3985,N_49988,N_49510);
nor UO_3986 (O_3986,N_49508,N_49668);
nor UO_3987 (O_3987,N_49891,N_49551);
and UO_3988 (O_3988,N_49639,N_49992);
xor UO_3989 (O_3989,N_49881,N_49540);
and UO_3990 (O_3990,N_49533,N_49806);
or UO_3991 (O_3991,N_49841,N_49561);
xor UO_3992 (O_3992,N_49527,N_49657);
and UO_3993 (O_3993,N_49926,N_49504);
xor UO_3994 (O_3994,N_49728,N_49505);
xor UO_3995 (O_3995,N_49812,N_49713);
and UO_3996 (O_3996,N_49686,N_49846);
nor UO_3997 (O_3997,N_49710,N_49998);
nor UO_3998 (O_3998,N_49767,N_49784);
nor UO_3999 (O_3999,N_49895,N_49616);
or UO_4000 (O_4000,N_49733,N_49868);
or UO_4001 (O_4001,N_49597,N_49688);
xor UO_4002 (O_4002,N_49897,N_49981);
xnor UO_4003 (O_4003,N_49571,N_49502);
nand UO_4004 (O_4004,N_49695,N_49890);
nand UO_4005 (O_4005,N_49943,N_49755);
nor UO_4006 (O_4006,N_49672,N_49701);
xor UO_4007 (O_4007,N_49582,N_49702);
and UO_4008 (O_4008,N_49642,N_49503);
nand UO_4009 (O_4009,N_49520,N_49842);
and UO_4010 (O_4010,N_49982,N_49571);
or UO_4011 (O_4011,N_49806,N_49599);
xnor UO_4012 (O_4012,N_49552,N_49846);
and UO_4013 (O_4013,N_49656,N_49915);
nor UO_4014 (O_4014,N_49564,N_49869);
or UO_4015 (O_4015,N_49549,N_49878);
or UO_4016 (O_4016,N_49748,N_49605);
xor UO_4017 (O_4017,N_49655,N_49902);
nand UO_4018 (O_4018,N_49908,N_49562);
nor UO_4019 (O_4019,N_49918,N_49931);
nor UO_4020 (O_4020,N_49973,N_49962);
nor UO_4021 (O_4021,N_49580,N_49849);
xnor UO_4022 (O_4022,N_49936,N_49903);
nand UO_4023 (O_4023,N_49774,N_49825);
nor UO_4024 (O_4024,N_49926,N_49964);
nor UO_4025 (O_4025,N_49606,N_49516);
nand UO_4026 (O_4026,N_49758,N_49984);
nand UO_4027 (O_4027,N_49871,N_49527);
xor UO_4028 (O_4028,N_49606,N_49963);
nor UO_4029 (O_4029,N_49898,N_49694);
xor UO_4030 (O_4030,N_49842,N_49822);
and UO_4031 (O_4031,N_49803,N_49595);
nor UO_4032 (O_4032,N_49664,N_49561);
and UO_4033 (O_4033,N_49605,N_49898);
nor UO_4034 (O_4034,N_49765,N_49935);
xnor UO_4035 (O_4035,N_49543,N_49600);
and UO_4036 (O_4036,N_49526,N_49867);
nor UO_4037 (O_4037,N_49576,N_49794);
nor UO_4038 (O_4038,N_49800,N_49808);
nor UO_4039 (O_4039,N_49670,N_49929);
or UO_4040 (O_4040,N_49847,N_49739);
nor UO_4041 (O_4041,N_49937,N_49749);
nand UO_4042 (O_4042,N_49753,N_49733);
xor UO_4043 (O_4043,N_49986,N_49764);
nor UO_4044 (O_4044,N_49998,N_49611);
nor UO_4045 (O_4045,N_49609,N_49804);
or UO_4046 (O_4046,N_49583,N_49584);
nor UO_4047 (O_4047,N_49569,N_49776);
nor UO_4048 (O_4048,N_49627,N_49892);
xor UO_4049 (O_4049,N_49926,N_49890);
xnor UO_4050 (O_4050,N_49675,N_49503);
or UO_4051 (O_4051,N_49502,N_49741);
xor UO_4052 (O_4052,N_49523,N_49771);
xnor UO_4053 (O_4053,N_49877,N_49548);
nand UO_4054 (O_4054,N_49614,N_49831);
xor UO_4055 (O_4055,N_49903,N_49519);
and UO_4056 (O_4056,N_49865,N_49944);
nor UO_4057 (O_4057,N_49948,N_49531);
and UO_4058 (O_4058,N_49759,N_49705);
nand UO_4059 (O_4059,N_49906,N_49892);
nand UO_4060 (O_4060,N_49546,N_49878);
xnor UO_4061 (O_4061,N_49798,N_49851);
or UO_4062 (O_4062,N_49592,N_49927);
and UO_4063 (O_4063,N_49659,N_49916);
nor UO_4064 (O_4064,N_49606,N_49610);
and UO_4065 (O_4065,N_49759,N_49514);
and UO_4066 (O_4066,N_49779,N_49925);
nor UO_4067 (O_4067,N_49826,N_49561);
and UO_4068 (O_4068,N_49769,N_49638);
and UO_4069 (O_4069,N_49503,N_49825);
nand UO_4070 (O_4070,N_49749,N_49672);
nor UO_4071 (O_4071,N_49988,N_49541);
nor UO_4072 (O_4072,N_49659,N_49996);
or UO_4073 (O_4073,N_49592,N_49596);
and UO_4074 (O_4074,N_49519,N_49992);
and UO_4075 (O_4075,N_49825,N_49771);
xor UO_4076 (O_4076,N_49765,N_49677);
nor UO_4077 (O_4077,N_49966,N_49968);
nor UO_4078 (O_4078,N_49902,N_49819);
and UO_4079 (O_4079,N_49979,N_49919);
or UO_4080 (O_4080,N_49539,N_49832);
nor UO_4081 (O_4081,N_49831,N_49657);
and UO_4082 (O_4082,N_49964,N_49546);
nand UO_4083 (O_4083,N_49758,N_49930);
nand UO_4084 (O_4084,N_49585,N_49610);
nand UO_4085 (O_4085,N_49659,N_49749);
nor UO_4086 (O_4086,N_49914,N_49503);
nand UO_4087 (O_4087,N_49615,N_49761);
nor UO_4088 (O_4088,N_49872,N_49624);
xor UO_4089 (O_4089,N_49793,N_49784);
and UO_4090 (O_4090,N_49836,N_49547);
and UO_4091 (O_4091,N_49600,N_49672);
and UO_4092 (O_4092,N_49653,N_49721);
or UO_4093 (O_4093,N_49559,N_49994);
xor UO_4094 (O_4094,N_49528,N_49850);
or UO_4095 (O_4095,N_49780,N_49787);
and UO_4096 (O_4096,N_49905,N_49723);
nor UO_4097 (O_4097,N_49555,N_49667);
xnor UO_4098 (O_4098,N_49806,N_49813);
nor UO_4099 (O_4099,N_49548,N_49755);
or UO_4100 (O_4100,N_49873,N_49645);
nand UO_4101 (O_4101,N_49714,N_49970);
nand UO_4102 (O_4102,N_49699,N_49584);
nand UO_4103 (O_4103,N_49766,N_49928);
nand UO_4104 (O_4104,N_49970,N_49754);
xnor UO_4105 (O_4105,N_49673,N_49766);
or UO_4106 (O_4106,N_49686,N_49549);
and UO_4107 (O_4107,N_49654,N_49636);
nor UO_4108 (O_4108,N_49782,N_49601);
and UO_4109 (O_4109,N_49831,N_49904);
nand UO_4110 (O_4110,N_49932,N_49883);
xor UO_4111 (O_4111,N_49669,N_49867);
xor UO_4112 (O_4112,N_49601,N_49762);
nand UO_4113 (O_4113,N_49988,N_49822);
nor UO_4114 (O_4114,N_49777,N_49644);
nor UO_4115 (O_4115,N_49959,N_49523);
or UO_4116 (O_4116,N_49972,N_49708);
nor UO_4117 (O_4117,N_49886,N_49680);
nor UO_4118 (O_4118,N_49694,N_49526);
or UO_4119 (O_4119,N_49622,N_49751);
nand UO_4120 (O_4120,N_49891,N_49513);
nor UO_4121 (O_4121,N_49957,N_49904);
nand UO_4122 (O_4122,N_49561,N_49835);
or UO_4123 (O_4123,N_49862,N_49927);
and UO_4124 (O_4124,N_49948,N_49703);
or UO_4125 (O_4125,N_49681,N_49912);
xor UO_4126 (O_4126,N_49584,N_49518);
or UO_4127 (O_4127,N_49801,N_49735);
nor UO_4128 (O_4128,N_49945,N_49714);
nand UO_4129 (O_4129,N_49565,N_49997);
and UO_4130 (O_4130,N_49808,N_49990);
nand UO_4131 (O_4131,N_49928,N_49922);
nand UO_4132 (O_4132,N_49872,N_49750);
xor UO_4133 (O_4133,N_49919,N_49677);
and UO_4134 (O_4134,N_49763,N_49697);
xnor UO_4135 (O_4135,N_49785,N_49586);
and UO_4136 (O_4136,N_49666,N_49665);
or UO_4137 (O_4137,N_49790,N_49565);
or UO_4138 (O_4138,N_49536,N_49820);
nor UO_4139 (O_4139,N_49737,N_49938);
nand UO_4140 (O_4140,N_49737,N_49804);
xnor UO_4141 (O_4141,N_49568,N_49959);
xnor UO_4142 (O_4142,N_49812,N_49783);
or UO_4143 (O_4143,N_49679,N_49925);
or UO_4144 (O_4144,N_49560,N_49582);
xnor UO_4145 (O_4145,N_49508,N_49837);
and UO_4146 (O_4146,N_49842,N_49688);
nand UO_4147 (O_4147,N_49600,N_49831);
or UO_4148 (O_4148,N_49536,N_49956);
or UO_4149 (O_4149,N_49767,N_49830);
and UO_4150 (O_4150,N_49985,N_49923);
or UO_4151 (O_4151,N_49930,N_49863);
nand UO_4152 (O_4152,N_49907,N_49611);
xnor UO_4153 (O_4153,N_49582,N_49719);
and UO_4154 (O_4154,N_49644,N_49814);
nor UO_4155 (O_4155,N_49741,N_49574);
nor UO_4156 (O_4156,N_49957,N_49964);
nand UO_4157 (O_4157,N_49651,N_49502);
nor UO_4158 (O_4158,N_49996,N_49675);
or UO_4159 (O_4159,N_49743,N_49788);
xnor UO_4160 (O_4160,N_49633,N_49599);
nor UO_4161 (O_4161,N_49890,N_49841);
and UO_4162 (O_4162,N_49615,N_49618);
nor UO_4163 (O_4163,N_49629,N_49652);
nand UO_4164 (O_4164,N_49680,N_49608);
nand UO_4165 (O_4165,N_49804,N_49674);
nand UO_4166 (O_4166,N_49946,N_49950);
and UO_4167 (O_4167,N_49731,N_49778);
xnor UO_4168 (O_4168,N_49651,N_49830);
nor UO_4169 (O_4169,N_49931,N_49943);
and UO_4170 (O_4170,N_49770,N_49568);
and UO_4171 (O_4171,N_49672,N_49560);
nor UO_4172 (O_4172,N_49748,N_49666);
and UO_4173 (O_4173,N_49645,N_49807);
nor UO_4174 (O_4174,N_49871,N_49601);
xor UO_4175 (O_4175,N_49520,N_49500);
xor UO_4176 (O_4176,N_49594,N_49568);
and UO_4177 (O_4177,N_49770,N_49998);
nand UO_4178 (O_4178,N_49577,N_49961);
nand UO_4179 (O_4179,N_49866,N_49912);
and UO_4180 (O_4180,N_49539,N_49632);
nor UO_4181 (O_4181,N_49641,N_49974);
xnor UO_4182 (O_4182,N_49574,N_49943);
nor UO_4183 (O_4183,N_49737,N_49785);
or UO_4184 (O_4184,N_49709,N_49610);
xnor UO_4185 (O_4185,N_49823,N_49821);
nor UO_4186 (O_4186,N_49864,N_49580);
or UO_4187 (O_4187,N_49872,N_49864);
or UO_4188 (O_4188,N_49980,N_49854);
xnor UO_4189 (O_4189,N_49552,N_49713);
or UO_4190 (O_4190,N_49692,N_49737);
and UO_4191 (O_4191,N_49823,N_49751);
or UO_4192 (O_4192,N_49733,N_49899);
or UO_4193 (O_4193,N_49723,N_49730);
and UO_4194 (O_4194,N_49869,N_49955);
nand UO_4195 (O_4195,N_49530,N_49931);
nand UO_4196 (O_4196,N_49554,N_49552);
and UO_4197 (O_4197,N_49987,N_49814);
xnor UO_4198 (O_4198,N_49520,N_49647);
nor UO_4199 (O_4199,N_49787,N_49510);
nor UO_4200 (O_4200,N_49688,N_49876);
xnor UO_4201 (O_4201,N_49916,N_49871);
or UO_4202 (O_4202,N_49633,N_49738);
or UO_4203 (O_4203,N_49869,N_49576);
xnor UO_4204 (O_4204,N_49612,N_49606);
and UO_4205 (O_4205,N_49660,N_49833);
or UO_4206 (O_4206,N_49905,N_49598);
xor UO_4207 (O_4207,N_49974,N_49967);
or UO_4208 (O_4208,N_49882,N_49616);
nor UO_4209 (O_4209,N_49930,N_49933);
or UO_4210 (O_4210,N_49906,N_49773);
xnor UO_4211 (O_4211,N_49986,N_49854);
or UO_4212 (O_4212,N_49855,N_49873);
nor UO_4213 (O_4213,N_49601,N_49748);
or UO_4214 (O_4214,N_49925,N_49895);
or UO_4215 (O_4215,N_49949,N_49742);
and UO_4216 (O_4216,N_49551,N_49556);
or UO_4217 (O_4217,N_49707,N_49939);
nor UO_4218 (O_4218,N_49837,N_49728);
nor UO_4219 (O_4219,N_49509,N_49669);
nor UO_4220 (O_4220,N_49615,N_49835);
xnor UO_4221 (O_4221,N_49984,N_49617);
xor UO_4222 (O_4222,N_49915,N_49630);
xor UO_4223 (O_4223,N_49997,N_49879);
nand UO_4224 (O_4224,N_49938,N_49755);
nor UO_4225 (O_4225,N_49895,N_49872);
or UO_4226 (O_4226,N_49735,N_49580);
xnor UO_4227 (O_4227,N_49507,N_49666);
and UO_4228 (O_4228,N_49606,N_49897);
nor UO_4229 (O_4229,N_49988,N_49894);
nor UO_4230 (O_4230,N_49826,N_49825);
nand UO_4231 (O_4231,N_49709,N_49762);
and UO_4232 (O_4232,N_49577,N_49732);
xnor UO_4233 (O_4233,N_49509,N_49949);
and UO_4234 (O_4234,N_49991,N_49936);
nand UO_4235 (O_4235,N_49621,N_49564);
xor UO_4236 (O_4236,N_49613,N_49961);
nor UO_4237 (O_4237,N_49942,N_49716);
nand UO_4238 (O_4238,N_49887,N_49702);
nand UO_4239 (O_4239,N_49862,N_49870);
xnor UO_4240 (O_4240,N_49659,N_49585);
and UO_4241 (O_4241,N_49515,N_49690);
nand UO_4242 (O_4242,N_49782,N_49557);
nand UO_4243 (O_4243,N_49870,N_49704);
nor UO_4244 (O_4244,N_49533,N_49516);
xnor UO_4245 (O_4245,N_49871,N_49636);
xnor UO_4246 (O_4246,N_49619,N_49506);
or UO_4247 (O_4247,N_49678,N_49508);
nor UO_4248 (O_4248,N_49719,N_49607);
or UO_4249 (O_4249,N_49712,N_49886);
and UO_4250 (O_4250,N_49731,N_49977);
xor UO_4251 (O_4251,N_49755,N_49882);
nand UO_4252 (O_4252,N_49768,N_49749);
nand UO_4253 (O_4253,N_49711,N_49704);
xnor UO_4254 (O_4254,N_49744,N_49806);
nor UO_4255 (O_4255,N_49806,N_49869);
or UO_4256 (O_4256,N_49833,N_49847);
or UO_4257 (O_4257,N_49743,N_49584);
or UO_4258 (O_4258,N_49651,N_49810);
and UO_4259 (O_4259,N_49707,N_49684);
xnor UO_4260 (O_4260,N_49665,N_49714);
nor UO_4261 (O_4261,N_49895,N_49557);
and UO_4262 (O_4262,N_49888,N_49577);
nand UO_4263 (O_4263,N_49833,N_49937);
nand UO_4264 (O_4264,N_49972,N_49886);
and UO_4265 (O_4265,N_49501,N_49556);
or UO_4266 (O_4266,N_49557,N_49873);
nor UO_4267 (O_4267,N_49707,N_49699);
nand UO_4268 (O_4268,N_49709,N_49991);
and UO_4269 (O_4269,N_49867,N_49706);
and UO_4270 (O_4270,N_49769,N_49558);
or UO_4271 (O_4271,N_49937,N_49674);
nor UO_4272 (O_4272,N_49987,N_49734);
and UO_4273 (O_4273,N_49614,N_49784);
nand UO_4274 (O_4274,N_49796,N_49698);
or UO_4275 (O_4275,N_49927,N_49848);
nor UO_4276 (O_4276,N_49780,N_49721);
xor UO_4277 (O_4277,N_49860,N_49673);
or UO_4278 (O_4278,N_49609,N_49748);
nor UO_4279 (O_4279,N_49941,N_49655);
or UO_4280 (O_4280,N_49749,N_49610);
and UO_4281 (O_4281,N_49991,N_49599);
xor UO_4282 (O_4282,N_49720,N_49815);
nand UO_4283 (O_4283,N_49635,N_49772);
or UO_4284 (O_4284,N_49709,N_49815);
nand UO_4285 (O_4285,N_49930,N_49936);
nand UO_4286 (O_4286,N_49687,N_49804);
or UO_4287 (O_4287,N_49730,N_49555);
nand UO_4288 (O_4288,N_49653,N_49882);
nand UO_4289 (O_4289,N_49905,N_49944);
xor UO_4290 (O_4290,N_49845,N_49761);
nor UO_4291 (O_4291,N_49580,N_49817);
nand UO_4292 (O_4292,N_49607,N_49903);
and UO_4293 (O_4293,N_49805,N_49750);
or UO_4294 (O_4294,N_49693,N_49772);
nor UO_4295 (O_4295,N_49816,N_49702);
nand UO_4296 (O_4296,N_49517,N_49779);
and UO_4297 (O_4297,N_49875,N_49812);
and UO_4298 (O_4298,N_49761,N_49800);
nand UO_4299 (O_4299,N_49973,N_49915);
and UO_4300 (O_4300,N_49633,N_49825);
or UO_4301 (O_4301,N_49831,N_49829);
nor UO_4302 (O_4302,N_49525,N_49557);
and UO_4303 (O_4303,N_49844,N_49689);
and UO_4304 (O_4304,N_49961,N_49621);
nor UO_4305 (O_4305,N_49823,N_49946);
nor UO_4306 (O_4306,N_49592,N_49506);
or UO_4307 (O_4307,N_49615,N_49722);
or UO_4308 (O_4308,N_49700,N_49502);
nand UO_4309 (O_4309,N_49984,N_49961);
and UO_4310 (O_4310,N_49994,N_49888);
or UO_4311 (O_4311,N_49759,N_49774);
xor UO_4312 (O_4312,N_49836,N_49559);
or UO_4313 (O_4313,N_49666,N_49902);
or UO_4314 (O_4314,N_49907,N_49811);
nor UO_4315 (O_4315,N_49897,N_49668);
or UO_4316 (O_4316,N_49749,N_49976);
and UO_4317 (O_4317,N_49948,N_49667);
or UO_4318 (O_4318,N_49902,N_49784);
nor UO_4319 (O_4319,N_49747,N_49757);
nand UO_4320 (O_4320,N_49956,N_49668);
or UO_4321 (O_4321,N_49910,N_49665);
nor UO_4322 (O_4322,N_49636,N_49568);
xnor UO_4323 (O_4323,N_49977,N_49734);
or UO_4324 (O_4324,N_49886,N_49546);
nand UO_4325 (O_4325,N_49800,N_49586);
nor UO_4326 (O_4326,N_49615,N_49553);
nor UO_4327 (O_4327,N_49518,N_49592);
or UO_4328 (O_4328,N_49673,N_49523);
nand UO_4329 (O_4329,N_49697,N_49850);
xor UO_4330 (O_4330,N_49944,N_49551);
and UO_4331 (O_4331,N_49991,N_49701);
xor UO_4332 (O_4332,N_49565,N_49870);
xnor UO_4333 (O_4333,N_49944,N_49800);
xor UO_4334 (O_4334,N_49949,N_49828);
or UO_4335 (O_4335,N_49818,N_49883);
or UO_4336 (O_4336,N_49698,N_49643);
nand UO_4337 (O_4337,N_49829,N_49527);
and UO_4338 (O_4338,N_49727,N_49858);
or UO_4339 (O_4339,N_49849,N_49939);
nor UO_4340 (O_4340,N_49853,N_49866);
xnor UO_4341 (O_4341,N_49544,N_49567);
nor UO_4342 (O_4342,N_49873,N_49751);
and UO_4343 (O_4343,N_49806,N_49517);
or UO_4344 (O_4344,N_49532,N_49521);
xor UO_4345 (O_4345,N_49917,N_49581);
or UO_4346 (O_4346,N_49813,N_49869);
xnor UO_4347 (O_4347,N_49947,N_49509);
xor UO_4348 (O_4348,N_49958,N_49911);
and UO_4349 (O_4349,N_49532,N_49718);
nor UO_4350 (O_4350,N_49528,N_49697);
xnor UO_4351 (O_4351,N_49901,N_49524);
or UO_4352 (O_4352,N_49770,N_49515);
nand UO_4353 (O_4353,N_49525,N_49535);
or UO_4354 (O_4354,N_49505,N_49889);
nand UO_4355 (O_4355,N_49888,N_49640);
nand UO_4356 (O_4356,N_49656,N_49678);
nand UO_4357 (O_4357,N_49527,N_49812);
and UO_4358 (O_4358,N_49889,N_49939);
or UO_4359 (O_4359,N_49672,N_49807);
and UO_4360 (O_4360,N_49886,N_49629);
or UO_4361 (O_4361,N_49532,N_49601);
or UO_4362 (O_4362,N_49888,N_49500);
nor UO_4363 (O_4363,N_49913,N_49711);
nand UO_4364 (O_4364,N_49648,N_49958);
and UO_4365 (O_4365,N_49698,N_49849);
xnor UO_4366 (O_4366,N_49646,N_49779);
or UO_4367 (O_4367,N_49880,N_49767);
and UO_4368 (O_4368,N_49860,N_49663);
or UO_4369 (O_4369,N_49511,N_49789);
nor UO_4370 (O_4370,N_49546,N_49654);
or UO_4371 (O_4371,N_49880,N_49709);
nor UO_4372 (O_4372,N_49812,N_49845);
nand UO_4373 (O_4373,N_49887,N_49666);
xor UO_4374 (O_4374,N_49646,N_49769);
or UO_4375 (O_4375,N_49786,N_49945);
nor UO_4376 (O_4376,N_49608,N_49583);
or UO_4377 (O_4377,N_49634,N_49550);
xnor UO_4378 (O_4378,N_49605,N_49751);
xor UO_4379 (O_4379,N_49886,N_49650);
and UO_4380 (O_4380,N_49934,N_49806);
xnor UO_4381 (O_4381,N_49801,N_49604);
nand UO_4382 (O_4382,N_49858,N_49838);
nor UO_4383 (O_4383,N_49620,N_49720);
nor UO_4384 (O_4384,N_49681,N_49639);
nand UO_4385 (O_4385,N_49862,N_49558);
or UO_4386 (O_4386,N_49774,N_49721);
nand UO_4387 (O_4387,N_49503,N_49539);
or UO_4388 (O_4388,N_49581,N_49647);
and UO_4389 (O_4389,N_49970,N_49950);
xor UO_4390 (O_4390,N_49996,N_49567);
nor UO_4391 (O_4391,N_49974,N_49980);
nor UO_4392 (O_4392,N_49649,N_49778);
nand UO_4393 (O_4393,N_49900,N_49912);
or UO_4394 (O_4394,N_49619,N_49880);
nand UO_4395 (O_4395,N_49903,N_49680);
nand UO_4396 (O_4396,N_49687,N_49977);
nor UO_4397 (O_4397,N_49974,N_49975);
and UO_4398 (O_4398,N_49869,N_49786);
nand UO_4399 (O_4399,N_49992,N_49658);
nor UO_4400 (O_4400,N_49729,N_49957);
nand UO_4401 (O_4401,N_49520,N_49590);
and UO_4402 (O_4402,N_49646,N_49869);
nor UO_4403 (O_4403,N_49667,N_49717);
nand UO_4404 (O_4404,N_49759,N_49610);
nand UO_4405 (O_4405,N_49716,N_49975);
nand UO_4406 (O_4406,N_49863,N_49861);
or UO_4407 (O_4407,N_49805,N_49897);
nand UO_4408 (O_4408,N_49775,N_49609);
and UO_4409 (O_4409,N_49677,N_49550);
nand UO_4410 (O_4410,N_49727,N_49876);
nor UO_4411 (O_4411,N_49806,N_49691);
nor UO_4412 (O_4412,N_49703,N_49567);
nor UO_4413 (O_4413,N_49666,N_49519);
xnor UO_4414 (O_4414,N_49526,N_49754);
xnor UO_4415 (O_4415,N_49994,N_49550);
nor UO_4416 (O_4416,N_49754,N_49647);
nor UO_4417 (O_4417,N_49640,N_49908);
xor UO_4418 (O_4418,N_49953,N_49622);
or UO_4419 (O_4419,N_49525,N_49927);
nand UO_4420 (O_4420,N_49702,N_49835);
nor UO_4421 (O_4421,N_49747,N_49922);
or UO_4422 (O_4422,N_49633,N_49735);
and UO_4423 (O_4423,N_49709,N_49535);
nor UO_4424 (O_4424,N_49553,N_49508);
nor UO_4425 (O_4425,N_49629,N_49550);
xor UO_4426 (O_4426,N_49621,N_49841);
or UO_4427 (O_4427,N_49608,N_49825);
nand UO_4428 (O_4428,N_49739,N_49667);
xor UO_4429 (O_4429,N_49588,N_49635);
nor UO_4430 (O_4430,N_49506,N_49542);
nand UO_4431 (O_4431,N_49777,N_49819);
nand UO_4432 (O_4432,N_49826,N_49600);
nor UO_4433 (O_4433,N_49734,N_49573);
or UO_4434 (O_4434,N_49672,N_49842);
xor UO_4435 (O_4435,N_49837,N_49622);
or UO_4436 (O_4436,N_49995,N_49611);
nor UO_4437 (O_4437,N_49699,N_49674);
nor UO_4438 (O_4438,N_49931,N_49916);
nor UO_4439 (O_4439,N_49780,N_49887);
or UO_4440 (O_4440,N_49587,N_49977);
or UO_4441 (O_4441,N_49706,N_49632);
xnor UO_4442 (O_4442,N_49714,N_49610);
nor UO_4443 (O_4443,N_49739,N_49621);
or UO_4444 (O_4444,N_49635,N_49595);
xor UO_4445 (O_4445,N_49647,N_49816);
nor UO_4446 (O_4446,N_49623,N_49864);
xnor UO_4447 (O_4447,N_49900,N_49641);
or UO_4448 (O_4448,N_49839,N_49786);
nand UO_4449 (O_4449,N_49846,N_49973);
xnor UO_4450 (O_4450,N_49848,N_49560);
or UO_4451 (O_4451,N_49611,N_49737);
xor UO_4452 (O_4452,N_49794,N_49943);
nor UO_4453 (O_4453,N_49919,N_49666);
nand UO_4454 (O_4454,N_49788,N_49516);
nand UO_4455 (O_4455,N_49850,N_49945);
or UO_4456 (O_4456,N_49927,N_49529);
and UO_4457 (O_4457,N_49568,N_49612);
nand UO_4458 (O_4458,N_49688,N_49659);
and UO_4459 (O_4459,N_49654,N_49674);
nor UO_4460 (O_4460,N_49861,N_49627);
xor UO_4461 (O_4461,N_49543,N_49638);
and UO_4462 (O_4462,N_49650,N_49521);
nand UO_4463 (O_4463,N_49815,N_49565);
nor UO_4464 (O_4464,N_49770,N_49882);
and UO_4465 (O_4465,N_49598,N_49983);
nand UO_4466 (O_4466,N_49972,N_49810);
xor UO_4467 (O_4467,N_49928,N_49744);
nor UO_4468 (O_4468,N_49888,N_49574);
nand UO_4469 (O_4469,N_49700,N_49520);
or UO_4470 (O_4470,N_49618,N_49942);
nand UO_4471 (O_4471,N_49625,N_49537);
xnor UO_4472 (O_4472,N_49889,N_49602);
nor UO_4473 (O_4473,N_49535,N_49652);
and UO_4474 (O_4474,N_49519,N_49616);
xnor UO_4475 (O_4475,N_49933,N_49932);
nand UO_4476 (O_4476,N_49638,N_49551);
nor UO_4477 (O_4477,N_49715,N_49521);
nor UO_4478 (O_4478,N_49924,N_49931);
xor UO_4479 (O_4479,N_49795,N_49563);
xnor UO_4480 (O_4480,N_49764,N_49802);
or UO_4481 (O_4481,N_49502,N_49619);
or UO_4482 (O_4482,N_49679,N_49511);
or UO_4483 (O_4483,N_49912,N_49588);
xnor UO_4484 (O_4484,N_49641,N_49556);
nand UO_4485 (O_4485,N_49560,N_49696);
or UO_4486 (O_4486,N_49549,N_49583);
nor UO_4487 (O_4487,N_49573,N_49705);
nand UO_4488 (O_4488,N_49661,N_49653);
and UO_4489 (O_4489,N_49614,N_49650);
or UO_4490 (O_4490,N_49759,N_49830);
nor UO_4491 (O_4491,N_49656,N_49807);
nand UO_4492 (O_4492,N_49711,N_49931);
nor UO_4493 (O_4493,N_49513,N_49893);
xor UO_4494 (O_4494,N_49592,N_49618);
or UO_4495 (O_4495,N_49727,N_49546);
nor UO_4496 (O_4496,N_49820,N_49578);
or UO_4497 (O_4497,N_49798,N_49680);
xor UO_4498 (O_4498,N_49997,N_49628);
xor UO_4499 (O_4499,N_49907,N_49954);
nand UO_4500 (O_4500,N_49870,N_49847);
xor UO_4501 (O_4501,N_49827,N_49959);
xor UO_4502 (O_4502,N_49663,N_49611);
xnor UO_4503 (O_4503,N_49507,N_49854);
nor UO_4504 (O_4504,N_49613,N_49950);
or UO_4505 (O_4505,N_49815,N_49729);
nor UO_4506 (O_4506,N_49666,N_49524);
and UO_4507 (O_4507,N_49937,N_49590);
or UO_4508 (O_4508,N_49722,N_49701);
nor UO_4509 (O_4509,N_49737,N_49635);
xor UO_4510 (O_4510,N_49832,N_49871);
nor UO_4511 (O_4511,N_49910,N_49992);
nor UO_4512 (O_4512,N_49939,N_49783);
or UO_4513 (O_4513,N_49737,N_49599);
nand UO_4514 (O_4514,N_49994,N_49741);
or UO_4515 (O_4515,N_49563,N_49847);
and UO_4516 (O_4516,N_49512,N_49934);
nor UO_4517 (O_4517,N_49530,N_49798);
and UO_4518 (O_4518,N_49882,N_49648);
xnor UO_4519 (O_4519,N_49626,N_49648);
nand UO_4520 (O_4520,N_49815,N_49947);
and UO_4521 (O_4521,N_49801,N_49816);
xor UO_4522 (O_4522,N_49982,N_49997);
and UO_4523 (O_4523,N_49614,N_49777);
nand UO_4524 (O_4524,N_49999,N_49975);
nand UO_4525 (O_4525,N_49974,N_49812);
or UO_4526 (O_4526,N_49626,N_49658);
nand UO_4527 (O_4527,N_49661,N_49904);
or UO_4528 (O_4528,N_49566,N_49590);
nor UO_4529 (O_4529,N_49857,N_49587);
xnor UO_4530 (O_4530,N_49697,N_49936);
nand UO_4531 (O_4531,N_49933,N_49897);
or UO_4532 (O_4532,N_49782,N_49556);
and UO_4533 (O_4533,N_49527,N_49627);
nor UO_4534 (O_4534,N_49511,N_49712);
or UO_4535 (O_4535,N_49576,N_49749);
and UO_4536 (O_4536,N_49871,N_49912);
and UO_4537 (O_4537,N_49683,N_49868);
xor UO_4538 (O_4538,N_49528,N_49522);
or UO_4539 (O_4539,N_49515,N_49641);
and UO_4540 (O_4540,N_49852,N_49523);
and UO_4541 (O_4541,N_49657,N_49848);
nor UO_4542 (O_4542,N_49633,N_49737);
nand UO_4543 (O_4543,N_49992,N_49799);
nor UO_4544 (O_4544,N_49992,N_49514);
or UO_4545 (O_4545,N_49762,N_49641);
nand UO_4546 (O_4546,N_49912,N_49616);
nor UO_4547 (O_4547,N_49573,N_49660);
nor UO_4548 (O_4548,N_49931,N_49576);
and UO_4549 (O_4549,N_49617,N_49749);
xnor UO_4550 (O_4550,N_49658,N_49768);
nor UO_4551 (O_4551,N_49721,N_49837);
nand UO_4552 (O_4552,N_49969,N_49884);
and UO_4553 (O_4553,N_49915,N_49797);
xnor UO_4554 (O_4554,N_49809,N_49959);
nor UO_4555 (O_4555,N_49639,N_49776);
xnor UO_4556 (O_4556,N_49997,N_49828);
or UO_4557 (O_4557,N_49683,N_49647);
nor UO_4558 (O_4558,N_49723,N_49886);
xnor UO_4559 (O_4559,N_49962,N_49593);
or UO_4560 (O_4560,N_49781,N_49851);
xnor UO_4561 (O_4561,N_49807,N_49541);
nand UO_4562 (O_4562,N_49864,N_49699);
or UO_4563 (O_4563,N_49876,N_49936);
nand UO_4564 (O_4564,N_49665,N_49987);
nor UO_4565 (O_4565,N_49860,N_49715);
nand UO_4566 (O_4566,N_49648,N_49549);
and UO_4567 (O_4567,N_49758,N_49685);
nand UO_4568 (O_4568,N_49684,N_49631);
or UO_4569 (O_4569,N_49713,N_49500);
and UO_4570 (O_4570,N_49572,N_49501);
and UO_4571 (O_4571,N_49504,N_49973);
xnor UO_4572 (O_4572,N_49954,N_49666);
nor UO_4573 (O_4573,N_49928,N_49641);
nor UO_4574 (O_4574,N_49749,N_49625);
or UO_4575 (O_4575,N_49539,N_49728);
or UO_4576 (O_4576,N_49620,N_49646);
and UO_4577 (O_4577,N_49909,N_49649);
xor UO_4578 (O_4578,N_49637,N_49769);
xnor UO_4579 (O_4579,N_49569,N_49578);
or UO_4580 (O_4580,N_49588,N_49785);
nor UO_4581 (O_4581,N_49585,N_49539);
and UO_4582 (O_4582,N_49692,N_49638);
or UO_4583 (O_4583,N_49558,N_49592);
and UO_4584 (O_4584,N_49655,N_49988);
xor UO_4585 (O_4585,N_49847,N_49873);
nand UO_4586 (O_4586,N_49919,N_49926);
nor UO_4587 (O_4587,N_49504,N_49990);
or UO_4588 (O_4588,N_49801,N_49963);
nand UO_4589 (O_4589,N_49715,N_49589);
and UO_4590 (O_4590,N_49670,N_49513);
and UO_4591 (O_4591,N_49591,N_49758);
nor UO_4592 (O_4592,N_49665,N_49743);
xnor UO_4593 (O_4593,N_49909,N_49542);
and UO_4594 (O_4594,N_49752,N_49924);
or UO_4595 (O_4595,N_49679,N_49890);
or UO_4596 (O_4596,N_49582,N_49926);
nand UO_4597 (O_4597,N_49670,N_49598);
nor UO_4598 (O_4598,N_49502,N_49541);
nand UO_4599 (O_4599,N_49746,N_49838);
and UO_4600 (O_4600,N_49856,N_49530);
xor UO_4601 (O_4601,N_49636,N_49828);
and UO_4602 (O_4602,N_49717,N_49979);
nand UO_4603 (O_4603,N_49743,N_49500);
nand UO_4604 (O_4604,N_49591,N_49836);
or UO_4605 (O_4605,N_49690,N_49677);
or UO_4606 (O_4606,N_49732,N_49627);
xnor UO_4607 (O_4607,N_49524,N_49614);
nor UO_4608 (O_4608,N_49528,N_49631);
nand UO_4609 (O_4609,N_49652,N_49596);
xnor UO_4610 (O_4610,N_49755,N_49509);
or UO_4611 (O_4611,N_49983,N_49581);
nor UO_4612 (O_4612,N_49717,N_49807);
xor UO_4613 (O_4613,N_49828,N_49781);
or UO_4614 (O_4614,N_49680,N_49920);
nand UO_4615 (O_4615,N_49845,N_49895);
nor UO_4616 (O_4616,N_49638,N_49925);
nor UO_4617 (O_4617,N_49868,N_49908);
or UO_4618 (O_4618,N_49529,N_49996);
xor UO_4619 (O_4619,N_49786,N_49991);
or UO_4620 (O_4620,N_49911,N_49952);
xor UO_4621 (O_4621,N_49714,N_49973);
nand UO_4622 (O_4622,N_49540,N_49826);
or UO_4623 (O_4623,N_49828,N_49814);
xor UO_4624 (O_4624,N_49837,N_49871);
and UO_4625 (O_4625,N_49581,N_49680);
or UO_4626 (O_4626,N_49901,N_49610);
nor UO_4627 (O_4627,N_49779,N_49941);
and UO_4628 (O_4628,N_49655,N_49565);
and UO_4629 (O_4629,N_49607,N_49727);
and UO_4630 (O_4630,N_49544,N_49778);
nand UO_4631 (O_4631,N_49858,N_49934);
and UO_4632 (O_4632,N_49839,N_49800);
or UO_4633 (O_4633,N_49945,N_49641);
nand UO_4634 (O_4634,N_49847,N_49732);
or UO_4635 (O_4635,N_49600,N_49725);
or UO_4636 (O_4636,N_49981,N_49850);
xnor UO_4637 (O_4637,N_49728,N_49765);
or UO_4638 (O_4638,N_49614,N_49619);
nand UO_4639 (O_4639,N_49676,N_49515);
xnor UO_4640 (O_4640,N_49760,N_49546);
nor UO_4641 (O_4641,N_49617,N_49637);
and UO_4642 (O_4642,N_49532,N_49507);
xnor UO_4643 (O_4643,N_49679,N_49607);
or UO_4644 (O_4644,N_49779,N_49546);
nand UO_4645 (O_4645,N_49816,N_49910);
and UO_4646 (O_4646,N_49771,N_49806);
nand UO_4647 (O_4647,N_49873,N_49504);
xnor UO_4648 (O_4648,N_49935,N_49653);
xor UO_4649 (O_4649,N_49627,N_49643);
nor UO_4650 (O_4650,N_49882,N_49854);
xnor UO_4651 (O_4651,N_49626,N_49886);
or UO_4652 (O_4652,N_49625,N_49637);
or UO_4653 (O_4653,N_49830,N_49876);
and UO_4654 (O_4654,N_49762,N_49537);
nor UO_4655 (O_4655,N_49792,N_49853);
and UO_4656 (O_4656,N_49748,N_49902);
nor UO_4657 (O_4657,N_49504,N_49753);
nor UO_4658 (O_4658,N_49783,N_49820);
and UO_4659 (O_4659,N_49579,N_49521);
or UO_4660 (O_4660,N_49713,N_49799);
nor UO_4661 (O_4661,N_49590,N_49693);
nor UO_4662 (O_4662,N_49706,N_49979);
nand UO_4663 (O_4663,N_49890,N_49830);
and UO_4664 (O_4664,N_49981,N_49766);
nand UO_4665 (O_4665,N_49808,N_49915);
xnor UO_4666 (O_4666,N_49889,N_49891);
nor UO_4667 (O_4667,N_49826,N_49925);
nor UO_4668 (O_4668,N_49959,N_49803);
xor UO_4669 (O_4669,N_49632,N_49580);
and UO_4670 (O_4670,N_49786,N_49693);
xnor UO_4671 (O_4671,N_49670,N_49740);
or UO_4672 (O_4672,N_49592,N_49970);
nor UO_4673 (O_4673,N_49632,N_49512);
or UO_4674 (O_4674,N_49745,N_49744);
and UO_4675 (O_4675,N_49971,N_49562);
or UO_4676 (O_4676,N_49519,N_49698);
nor UO_4677 (O_4677,N_49691,N_49919);
nor UO_4678 (O_4678,N_49756,N_49650);
xnor UO_4679 (O_4679,N_49918,N_49719);
and UO_4680 (O_4680,N_49559,N_49801);
and UO_4681 (O_4681,N_49876,N_49709);
and UO_4682 (O_4682,N_49800,N_49701);
nand UO_4683 (O_4683,N_49918,N_49580);
xnor UO_4684 (O_4684,N_49641,N_49625);
or UO_4685 (O_4685,N_49502,N_49932);
xnor UO_4686 (O_4686,N_49626,N_49791);
or UO_4687 (O_4687,N_49962,N_49824);
xnor UO_4688 (O_4688,N_49955,N_49780);
nand UO_4689 (O_4689,N_49941,N_49791);
nand UO_4690 (O_4690,N_49999,N_49659);
and UO_4691 (O_4691,N_49556,N_49844);
xnor UO_4692 (O_4692,N_49837,N_49866);
nand UO_4693 (O_4693,N_49574,N_49714);
xor UO_4694 (O_4694,N_49913,N_49895);
xor UO_4695 (O_4695,N_49677,N_49783);
nor UO_4696 (O_4696,N_49717,N_49822);
or UO_4697 (O_4697,N_49903,N_49656);
nor UO_4698 (O_4698,N_49936,N_49586);
nand UO_4699 (O_4699,N_49708,N_49730);
and UO_4700 (O_4700,N_49599,N_49909);
and UO_4701 (O_4701,N_49827,N_49775);
or UO_4702 (O_4702,N_49820,N_49733);
xor UO_4703 (O_4703,N_49587,N_49818);
nor UO_4704 (O_4704,N_49545,N_49519);
xnor UO_4705 (O_4705,N_49666,N_49529);
nand UO_4706 (O_4706,N_49948,N_49505);
nor UO_4707 (O_4707,N_49821,N_49606);
nand UO_4708 (O_4708,N_49574,N_49579);
xnor UO_4709 (O_4709,N_49948,N_49877);
xor UO_4710 (O_4710,N_49997,N_49678);
nand UO_4711 (O_4711,N_49867,N_49740);
nor UO_4712 (O_4712,N_49746,N_49988);
nor UO_4713 (O_4713,N_49848,N_49849);
xnor UO_4714 (O_4714,N_49741,N_49859);
nand UO_4715 (O_4715,N_49996,N_49978);
nor UO_4716 (O_4716,N_49529,N_49959);
nor UO_4717 (O_4717,N_49822,N_49748);
xor UO_4718 (O_4718,N_49842,N_49820);
or UO_4719 (O_4719,N_49758,N_49500);
or UO_4720 (O_4720,N_49855,N_49505);
nor UO_4721 (O_4721,N_49768,N_49816);
nand UO_4722 (O_4722,N_49567,N_49522);
nand UO_4723 (O_4723,N_49760,N_49836);
nand UO_4724 (O_4724,N_49941,N_49533);
or UO_4725 (O_4725,N_49896,N_49705);
xnor UO_4726 (O_4726,N_49512,N_49722);
and UO_4727 (O_4727,N_49930,N_49842);
or UO_4728 (O_4728,N_49975,N_49691);
xor UO_4729 (O_4729,N_49880,N_49813);
xor UO_4730 (O_4730,N_49750,N_49727);
and UO_4731 (O_4731,N_49687,N_49842);
or UO_4732 (O_4732,N_49903,N_49713);
nor UO_4733 (O_4733,N_49694,N_49504);
nand UO_4734 (O_4734,N_49805,N_49876);
and UO_4735 (O_4735,N_49515,N_49978);
nand UO_4736 (O_4736,N_49704,N_49597);
or UO_4737 (O_4737,N_49922,N_49815);
xnor UO_4738 (O_4738,N_49923,N_49652);
xnor UO_4739 (O_4739,N_49686,N_49743);
nor UO_4740 (O_4740,N_49976,N_49719);
xnor UO_4741 (O_4741,N_49556,N_49949);
nor UO_4742 (O_4742,N_49888,N_49848);
nor UO_4743 (O_4743,N_49988,N_49574);
nand UO_4744 (O_4744,N_49590,N_49742);
nor UO_4745 (O_4745,N_49951,N_49885);
nand UO_4746 (O_4746,N_49781,N_49522);
nand UO_4747 (O_4747,N_49834,N_49631);
xor UO_4748 (O_4748,N_49899,N_49806);
or UO_4749 (O_4749,N_49870,N_49921);
nor UO_4750 (O_4750,N_49946,N_49598);
nor UO_4751 (O_4751,N_49861,N_49784);
and UO_4752 (O_4752,N_49668,N_49580);
nand UO_4753 (O_4753,N_49716,N_49814);
nor UO_4754 (O_4754,N_49665,N_49578);
nand UO_4755 (O_4755,N_49584,N_49655);
nor UO_4756 (O_4756,N_49773,N_49849);
xnor UO_4757 (O_4757,N_49540,N_49883);
or UO_4758 (O_4758,N_49679,N_49677);
and UO_4759 (O_4759,N_49999,N_49527);
nor UO_4760 (O_4760,N_49858,N_49779);
xor UO_4761 (O_4761,N_49506,N_49993);
and UO_4762 (O_4762,N_49545,N_49639);
nand UO_4763 (O_4763,N_49768,N_49974);
nand UO_4764 (O_4764,N_49559,N_49629);
or UO_4765 (O_4765,N_49735,N_49844);
nand UO_4766 (O_4766,N_49903,N_49940);
xnor UO_4767 (O_4767,N_49722,N_49866);
xnor UO_4768 (O_4768,N_49872,N_49995);
nor UO_4769 (O_4769,N_49722,N_49931);
nor UO_4770 (O_4770,N_49524,N_49807);
and UO_4771 (O_4771,N_49675,N_49823);
nand UO_4772 (O_4772,N_49832,N_49668);
nand UO_4773 (O_4773,N_49800,N_49853);
or UO_4774 (O_4774,N_49813,N_49522);
nor UO_4775 (O_4775,N_49929,N_49797);
and UO_4776 (O_4776,N_49740,N_49798);
or UO_4777 (O_4777,N_49986,N_49554);
nand UO_4778 (O_4778,N_49762,N_49773);
and UO_4779 (O_4779,N_49723,N_49944);
or UO_4780 (O_4780,N_49504,N_49793);
nand UO_4781 (O_4781,N_49873,N_49940);
nand UO_4782 (O_4782,N_49990,N_49510);
and UO_4783 (O_4783,N_49551,N_49653);
nor UO_4784 (O_4784,N_49978,N_49787);
xor UO_4785 (O_4785,N_49506,N_49790);
and UO_4786 (O_4786,N_49952,N_49859);
or UO_4787 (O_4787,N_49701,N_49761);
nor UO_4788 (O_4788,N_49693,N_49759);
xor UO_4789 (O_4789,N_49785,N_49973);
or UO_4790 (O_4790,N_49614,N_49622);
or UO_4791 (O_4791,N_49785,N_49592);
xnor UO_4792 (O_4792,N_49904,N_49899);
nand UO_4793 (O_4793,N_49960,N_49597);
nor UO_4794 (O_4794,N_49868,N_49671);
nor UO_4795 (O_4795,N_49962,N_49886);
and UO_4796 (O_4796,N_49844,N_49999);
xor UO_4797 (O_4797,N_49514,N_49952);
xnor UO_4798 (O_4798,N_49877,N_49887);
nand UO_4799 (O_4799,N_49891,N_49566);
nor UO_4800 (O_4800,N_49561,N_49591);
nand UO_4801 (O_4801,N_49552,N_49562);
xor UO_4802 (O_4802,N_49596,N_49567);
or UO_4803 (O_4803,N_49660,N_49777);
and UO_4804 (O_4804,N_49562,N_49678);
nor UO_4805 (O_4805,N_49641,N_49993);
nor UO_4806 (O_4806,N_49521,N_49588);
and UO_4807 (O_4807,N_49919,N_49816);
and UO_4808 (O_4808,N_49897,N_49832);
and UO_4809 (O_4809,N_49614,N_49638);
nor UO_4810 (O_4810,N_49977,N_49823);
nor UO_4811 (O_4811,N_49890,N_49518);
nand UO_4812 (O_4812,N_49920,N_49944);
or UO_4813 (O_4813,N_49561,N_49921);
xnor UO_4814 (O_4814,N_49882,N_49741);
nand UO_4815 (O_4815,N_49854,N_49984);
or UO_4816 (O_4816,N_49648,N_49892);
and UO_4817 (O_4817,N_49537,N_49928);
or UO_4818 (O_4818,N_49545,N_49524);
xor UO_4819 (O_4819,N_49518,N_49817);
nor UO_4820 (O_4820,N_49699,N_49782);
and UO_4821 (O_4821,N_49888,N_49511);
nand UO_4822 (O_4822,N_49881,N_49971);
or UO_4823 (O_4823,N_49614,N_49901);
nand UO_4824 (O_4824,N_49804,N_49859);
xor UO_4825 (O_4825,N_49697,N_49865);
and UO_4826 (O_4826,N_49588,N_49950);
or UO_4827 (O_4827,N_49995,N_49669);
nor UO_4828 (O_4828,N_49991,N_49990);
and UO_4829 (O_4829,N_49938,N_49506);
xor UO_4830 (O_4830,N_49901,N_49742);
xnor UO_4831 (O_4831,N_49717,N_49990);
xnor UO_4832 (O_4832,N_49859,N_49968);
nand UO_4833 (O_4833,N_49890,N_49710);
nor UO_4834 (O_4834,N_49797,N_49503);
or UO_4835 (O_4835,N_49561,N_49979);
nor UO_4836 (O_4836,N_49527,N_49955);
or UO_4837 (O_4837,N_49967,N_49884);
nor UO_4838 (O_4838,N_49669,N_49550);
nor UO_4839 (O_4839,N_49695,N_49788);
nand UO_4840 (O_4840,N_49546,N_49947);
and UO_4841 (O_4841,N_49541,N_49757);
and UO_4842 (O_4842,N_49695,N_49547);
xor UO_4843 (O_4843,N_49952,N_49978);
nor UO_4844 (O_4844,N_49792,N_49533);
or UO_4845 (O_4845,N_49797,N_49856);
nand UO_4846 (O_4846,N_49743,N_49797);
or UO_4847 (O_4847,N_49701,N_49827);
or UO_4848 (O_4848,N_49528,N_49535);
or UO_4849 (O_4849,N_49689,N_49690);
nand UO_4850 (O_4850,N_49764,N_49650);
nor UO_4851 (O_4851,N_49993,N_49865);
or UO_4852 (O_4852,N_49936,N_49788);
and UO_4853 (O_4853,N_49852,N_49501);
and UO_4854 (O_4854,N_49592,N_49825);
xnor UO_4855 (O_4855,N_49840,N_49746);
nor UO_4856 (O_4856,N_49624,N_49694);
xnor UO_4857 (O_4857,N_49818,N_49599);
nor UO_4858 (O_4858,N_49877,N_49651);
and UO_4859 (O_4859,N_49997,N_49556);
nor UO_4860 (O_4860,N_49546,N_49963);
or UO_4861 (O_4861,N_49851,N_49622);
nor UO_4862 (O_4862,N_49696,N_49677);
nor UO_4863 (O_4863,N_49840,N_49736);
and UO_4864 (O_4864,N_49710,N_49938);
and UO_4865 (O_4865,N_49744,N_49611);
or UO_4866 (O_4866,N_49832,N_49921);
xor UO_4867 (O_4867,N_49738,N_49787);
or UO_4868 (O_4868,N_49533,N_49930);
nor UO_4869 (O_4869,N_49760,N_49799);
nand UO_4870 (O_4870,N_49994,N_49739);
and UO_4871 (O_4871,N_49889,N_49746);
or UO_4872 (O_4872,N_49852,N_49753);
and UO_4873 (O_4873,N_49678,N_49770);
or UO_4874 (O_4874,N_49887,N_49639);
nor UO_4875 (O_4875,N_49536,N_49803);
nor UO_4876 (O_4876,N_49845,N_49755);
xor UO_4877 (O_4877,N_49793,N_49892);
and UO_4878 (O_4878,N_49519,N_49846);
and UO_4879 (O_4879,N_49922,N_49623);
nand UO_4880 (O_4880,N_49952,N_49620);
xnor UO_4881 (O_4881,N_49876,N_49862);
and UO_4882 (O_4882,N_49526,N_49875);
nor UO_4883 (O_4883,N_49605,N_49545);
xor UO_4884 (O_4884,N_49524,N_49731);
or UO_4885 (O_4885,N_49901,N_49784);
or UO_4886 (O_4886,N_49743,N_49613);
or UO_4887 (O_4887,N_49552,N_49569);
xnor UO_4888 (O_4888,N_49624,N_49506);
nor UO_4889 (O_4889,N_49727,N_49547);
or UO_4890 (O_4890,N_49760,N_49566);
xor UO_4891 (O_4891,N_49550,N_49530);
nor UO_4892 (O_4892,N_49683,N_49897);
and UO_4893 (O_4893,N_49835,N_49746);
and UO_4894 (O_4894,N_49589,N_49864);
nand UO_4895 (O_4895,N_49571,N_49816);
or UO_4896 (O_4896,N_49613,N_49735);
or UO_4897 (O_4897,N_49652,N_49675);
nand UO_4898 (O_4898,N_49973,N_49650);
xnor UO_4899 (O_4899,N_49817,N_49990);
nor UO_4900 (O_4900,N_49613,N_49551);
or UO_4901 (O_4901,N_49913,N_49980);
xnor UO_4902 (O_4902,N_49759,N_49719);
and UO_4903 (O_4903,N_49563,N_49787);
and UO_4904 (O_4904,N_49526,N_49965);
and UO_4905 (O_4905,N_49741,N_49732);
and UO_4906 (O_4906,N_49986,N_49925);
and UO_4907 (O_4907,N_49748,N_49710);
and UO_4908 (O_4908,N_49726,N_49605);
nor UO_4909 (O_4909,N_49703,N_49623);
xor UO_4910 (O_4910,N_49805,N_49855);
or UO_4911 (O_4911,N_49709,N_49673);
and UO_4912 (O_4912,N_49807,N_49691);
or UO_4913 (O_4913,N_49960,N_49988);
or UO_4914 (O_4914,N_49771,N_49785);
nand UO_4915 (O_4915,N_49773,N_49841);
xor UO_4916 (O_4916,N_49832,N_49966);
nand UO_4917 (O_4917,N_49984,N_49635);
or UO_4918 (O_4918,N_49844,N_49762);
nor UO_4919 (O_4919,N_49860,N_49583);
nand UO_4920 (O_4920,N_49636,N_49703);
or UO_4921 (O_4921,N_49963,N_49811);
nand UO_4922 (O_4922,N_49759,N_49720);
nor UO_4923 (O_4923,N_49626,N_49748);
and UO_4924 (O_4924,N_49684,N_49522);
and UO_4925 (O_4925,N_49885,N_49588);
xnor UO_4926 (O_4926,N_49646,N_49605);
xor UO_4927 (O_4927,N_49635,N_49989);
xnor UO_4928 (O_4928,N_49526,N_49870);
nor UO_4929 (O_4929,N_49655,N_49899);
or UO_4930 (O_4930,N_49704,N_49963);
nand UO_4931 (O_4931,N_49620,N_49614);
or UO_4932 (O_4932,N_49829,N_49521);
or UO_4933 (O_4933,N_49605,N_49639);
nor UO_4934 (O_4934,N_49890,N_49991);
and UO_4935 (O_4935,N_49741,N_49821);
xor UO_4936 (O_4936,N_49969,N_49961);
xnor UO_4937 (O_4937,N_49869,N_49660);
xor UO_4938 (O_4938,N_49626,N_49722);
and UO_4939 (O_4939,N_49872,N_49537);
nand UO_4940 (O_4940,N_49542,N_49835);
nor UO_4941 (O_4941,N_49647,N_49942);
and UO_4942 (O_4942,N_49881,N_49865);
nor UO_4943 (O_4943,N_49911,N_49621);
or UO_4944 (O_4944,N_49588,N_49977);
nand UO_4945 (O_4945,N_49783,N_49979);
nand UO_4946 (O_4946,N_49964,N_49563);
and UO_4947 (O_4947,N_49744,N_49903);
nor UO_4948 (O_4948,N_49843,N_49721);
nor UO_4949 (O_4949,N_49981,N_49715);
and UO_4950 (O_4950,N_49854,N_49583);
or UO_4951 (O_4951,N_49926,N_49661);
or UO_4952 (O_4952,N_49698,N_49661);
or UO_4953 (O_4953,N_49789,N_49837);
xor UO_4954 (O_4954,N_49970,N_49550);
and UO_4955 (O_4955,N_49661,N_49597);
or UO_4956 (O_4956,N_49732,N_49730);
nand UO_4957 (O_4957,N_49787,N_49764);
and UO_4958 (O_4958,N_49675,N_49724);
nor UO_4959 (O_4959,N_49529,N_49974);
or UO_4960 (O_4960,N_49548,N_49849);
and UO_4961 (O_4961,N_49569,N_49746);
xnor UO_4962 (O_4962,N_49868,N_49918);
nand UO_4963 (O_4963,N_49807,N_49735);
xor UO_4964 (O_4964,N_49779,N_49631);
and UO_4965 (O_4965,N_49842,N_49873);
xnor UO_4966 (O_4966,N_49642,N_49685);
nor UO_4967 (O_4967,N_49568,N_49714);
and UO_4968 (O_4968,N_49728,N_49534);
or UO_4969 (O_4969,N_49816,N_49671);
nor UO_4970 (O_4970,N_49790,N_49640);
nand UO_4971 (O_4971,N_49809,N_49633);
or UO_4972 (O_4972,N_49993,N_49689);
xor UO_4973 (O_4973,N_49873,N_49525);
nor UO_4974 (O_4974,N_49716,N_49578);
nand UO_4975 (O_4975,N_49765,N_49784);
or UO_4976 (O_4976,N_49825,N_49935);
or UO_4977 (O_4977,N_49607,N_49728);
and UO_4978 (O_4978,N_49591,N_49769);
nor UO_4979 (O_4979,N_49728,N_49707);
nor UO_4980 (O_4980,N_49842,N_49938);
nand UO_4981 (O_4981,N_49561,N_49887);
nand UO_4982 (O_4982,N_49881,N_49693);
and UO_4983 (O_4983,N_49806,N_49879);
or UO_4984 (O_4984,N_49904,N_49718);
nor UO_4985 (O_4985,N_49682,N_49501);
and UO_4986 (O_4986,N_49762,N_49943);
and UO_4987 (O_4987,N_49742,N_49760);
xnor UO_4988 (O_4988,N_49978,N_49504);
xor UO_4989 (O_4989,N_49967,N_49504);
and UO_4990 (O_4990,N_49821,N_49617);
nand UO_4991 (O_4991,N_49676,N_49769);
nor UO_4992 (O_4992,N_49614,N_49806);
and UO_4993 (O_4993,N_49716,N_49743);
nor UO_4994 (O_4994,N_49650,N_49857);
and UO_4995 (O_4995,N_49884,N_49922);
and UO_4996 (O_4996,N_49972,N_49942);
nand UO_4997 (O_4997,N_49867,N_49920);
xnor UO_4998 (O_4998,N_49683,N_49554);
and UO_4999 (O_4999,N_49610,N_49900);
endmodule