module basic_500_3000_500_30_levels_10xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
xor U0 (N_0,In_209,In_455);
nor U1 (N_1,In_320,In_164);
and U2 (N_2,In_473,In_29);
nand U3 (N_3,In_138,In_293);
xor U4 (N_4,In_441,In_56);
and U5 (N_5,In_171,In_264);
xnor U6 (N_6,In_90,In_329);
and U7 (N_7,In_223,In_351);
xnor U8 (N_8,In_80,In_290);
and U9 (N_9,In_435,In_417);
xor U10 (N_10,In_96,In_428);
xor U11 (N_11,In_477,In_85);
nor U12 (N_12,In_134,In_247);
nand U13 (N_13,In_115,In_284);
xnor U14 (N_14,In_445,In_287);
xnor U15 (N_15,In_265,In_88);
xnor U16 (N_16,In_466,In_470);
or U17 (N_17,In_394,In_268);
nand U18 (N_18,In_222,In_49);
and U19 (N_19,In_73,In_195);
xor U20 (N_20,In_352,In_46);
xnor U21 (N_21,In_464,In_336);
nor U22 (N_22,In_230,In_108);
nor U23 (N_23,In_296,In_388);
xor U24 (N_24,In_135,In_12);
nor U25 (N_25,In_14,In_163);
or U26 (N_26,In_493,In_93);
and U27 (N_27,In_68,In_407);
and U28 (N_28,In_60,In_32);
xnor U29 (N_29,In_0,In_459);
or U30 (N_30,In_308,In_67);
or U31 (N_31,In_468,In_159);
or U32 (N_32,In_316,In_208);
and U33 (N_33,In_201,In_393);
or U34 (N_34,In_259,In_182);
and U35 (N_35,In_349,In_360);
and U36 (N_36,In_101,In_365);
or U37 (N_37,In_430,In_397);
and U38 (N_38,In_144,In_2);
and U39 (N_39,In_147,In_215);
xnor U40 (N_40,In_168,In_494);
nor U41 (N_41,In_160,In_239);
nand U42 (N_42,In_326,In_252);
nor U43 (N_43,In_420,In_406);
nand U44 (N_44,In_399,In_367);
nand U45 (N_45,In_314,In_57);
or U46 (N_46,In_364,In_153);
and U47 (N_47,In_346,In_237);
xor U48 (N_48,In_124,In_234);
xor U49 (N_49,In_26,In_465);
nor U50 (N_50,In_109,In_489);
xor U51 (N_51,In_301,In_43);
xnor U52 (N_52,In_382,In_104);
or U53 (N_53,In_156,In_275);
nand U54 (N_54,In_51,In_184);
nand U55 (N_55,In_288,In_335);
nor U56 (N_56,In_321,In_419);
nand U57 (N_57,In_269,In_169);
or U58 (N_58,In_118,In_61);
nand U59 (N_59,In_220,In_149);
nand U60 (N_60,In_206,In_368);
and U61 (N_61,In_426,In_113);
xnor U62 (N_62,In_392,In_189);
nand U63 (N_63,In_389,In_75);
xnor U64 (N_64,In_436,In_112);
xor U65 (N_65,In_28,In_236);
xor U66 (N_66,In_338,In_83);
or U67 (N_67,In_110,In_272);
xnor U68 (N_68,In_150,In_432);
and U69 (N_69,In_19,In_69);
and U70 (N_70,In_409,In_356);
and U71 (N_71,In_255,In_276);
and U72 (N_72,In_188,In_20);
nor U73 (N_73,In_373,In_345);
xor U74 (N_74,In_421,In_361);
nand U75 (N_75,In_196,In_309);
and U76 (N_76,In_377,In_100);
and U77 (N_77,In_454,In_121);
and U78 (N_78,In_89,In_111);
xnor U79 (N_79,In_327,In_344);
or U80 (N_80,In_337,In_246);
nor U81 (N_81,In_312,In_353);
nand U82 (N_82,In_376,In_241);
nor U83 (N_83,In_490,In_400);
xor U84 (N_84,In_273,In_487);
and U85 (N_85,In_181,In_91);
or U86 (N_86,In_343,In_44);
or U87 (N_87,In_190,In_439);
and U88 (N_88,In_461,In_38);
xor U89 (N_89,In_324,In_257);
or U90 (N_90,In_47,In_292);
nor U91 (N_91,In_205,In_42);
or U92 (N_92,In_45,In_34);
nand U93 (N_93,In_307,In_282);
nor U94 (N_94,In_64,In_281);
nand U95 (N_95,In_262,In_130);
nor U96 (N_96,In_243,In_383);
nand U97 (N_97,In_238,In_175);
xor U98 (N_98,In_18,In_120);
nand U99 (N_99,In_183,In_313);
nor U100 (N_100,N_20,In_418);
and U101 (N_101,N_52,In_192);
or U102 (N_102,N_49,In_10);
nor U103 (N_103,N_23,In_374);
nand U104 (N_104,In_126,In_416);
nor U105 (N_105,In_359,In_232);
or U106 (N_106,In_251,In_289);
nand U107 (N_107,N_19,In_87);
nand U108 (N_108,N_98,In_488);
and U109 (N_109,In_350,In_161);
nand U110 (N_110,In_433,In_178);
or U111 (N_111,N_16,In_261);
xor U112 (N_112,N_31,In_71);
nor U113 (N_113,In_166,In_131);
and U114 (N_114,In_481,In_410);
nand U115 (N_115,In_146,In_244);
nor U116 (N_116,In_363,In_267);
xnor U117 (N_117,In_381,N_99);
and U118 (N_118,In_391,N_62);
xnor U119 (N_119,In_429,N_32);
nor U120 (N_120,N_89,In_200);
xor U121 (N_121,N_68,In_228);
and U122 (N_122,N_9,In_129);
nand U123 (N_123,In_52,N_15);
xor U124 (N_124,In_41,In_362);
nand U125 (N_125,In_6,N_39);
nor U126 (N_126,N_58,In_127);
and U127 (N_127,In_125,In_483);
or U128 (N_128,In_194,N_0);
and U129 (N_129,N_54,In_438);
xnor U130 (N_130,In_491,In_35);
nor U131 (N_131,N_36,In_81);
xor U132 (N_132,In_177,N_75);
nand U133 (N_133,N_91,In_306);
or U134 (N_134,In_425,In_339);
or U135 (N_135,In_385,In_444);
nor U136 (N_136,In_7,In_225);
nor U137 (N_137,N_3,In_453);
xnor U138 (N_138,In_242,N_25);
nand U139 (N_139,In_27,In_97);
xnor U140 (N_140,N_30,In_13);
xnor U141 (N_141,In_423,In_245);
nand U142 (N_142,In_142,In_202);
nor U143 (N_143,In_231,In_58);
or U144 (N_144,In_270,In_498);
and U145 (N_145,In_1,In_133);
and U146 (N_146,N_93,In_250);
and U147 (N_147,In_145,In_63);
nor U148 (N_148,In_132,In_317);
or U149 (N_149,In_198,In_25);
nand U150 (N_150,In_476,In_66);
and U151 (N_151,In_319,In_462);
or U152 (N_152,In_387,N_72);
nand U153 (N_153,In_176,In_357);
xor U154 (N_154,N_78,N_18);
and U155 (N_155,In_229,N_13);
nand U156 (N_156,In_492,In_98);
nor U157 (N_157,In_325,In_180);
xnor U158 (N_158,N_69,In_347);
xor U159 (N_159,N_37,In_154);
nor U160 (N_160,In_213,In_408);
xnor U161 (N_161,In_24,In_17);
nand U162 (N_162,N_22,N_57);
nand U163 (N_163,In_412,In_405);
and U164 (N_164,In_48,In_136);
xor U165 (N_165,In_210,In_370);
nor U166 (N_166,In_65,In_119);
or U167 (N_167,In_499,In_369);
and U168 (N_168,In_170,In_411);
and U169 (N_169,In_260,In_318);
nor U170 (N_170,In_139,In_82);
nor U171 (N_171,N_79,In_114);
or U172 (N_172,In_323,In_186);
nor U173 (N_173,In_141,In_463);
or U174 (N_174,In_271,In_431);
nor U175 (N_175,In_390,In_174);
nand U176 (N_176,In_157,In_50);
nand U177 (N_177,In_76,N_12);
xnor U178 (N_178,In_216,N_60);
nand U179 (N_179,N_51,In_414);
and U180 (N_180,In_62,In_437);
and U181 (N_181,In_446,In_117);
nand U182 (N_182,N_67,N_34);
nor U183 (N_183,In_480,In_92);
xor U184 (N_184,In_106,In_342);
nand U185 (N_185,In_277,In_297);
xor U186 (N_186,In_404,In_137);
xnor U187 (N_187,N_61,In_331);
or U188 (N_188,In_207,In_274);
nor U189 (N_189,In_22,In_280);
nand U190 (N_190,In_116,N_76);
xnor U191 (N_191,In_315,N_43);
nand U192 (N_192,In_122,In_475);
nand U193 (N_193,In_84,In_187);
xnor U194 (N_194,In_224,In_219);
xor U195 (N_195,In_53,In_380);
nand U196 (N_196,In_99,N_44);
nand U197 (N_197,In_330,In_458);
or U198 (N_198,In_31,In_371);
or U199 (N_199,In_451,In_413);
xor U200 (N_200,N_190,In_162);
and U201 (N_201,In_295,In_94);
and U202 (N_202,N_192,N_50);
and U203 (N_203,In_77,In_193);
xnor U204 (N_204,In_4,N_77);
xor U205 (N_205,In_333,In_3);
xor U206 (N_206,N_105,In_403);
xor U207 (N_207,N_96,In_332);
nor U208 (N_208,In_310,N_94);
nand U209 (N_209,N_123,In_298);
or U210 (N_210,N_155,In_442);
nor U211 (N_211,In_203,In_304);
or U212 (N_212,N_156,N_38);
or U213 (N_213,N_198,In_484);
xor U214 (N_214,In_375,N_83);
nor U215 (N_215,In_165,In_128);
nand U216 (N_216,In_221,N_132);
or U217 (N_217,N_128,N_181);
nand U218 (N_218,In_218,In_217);
nand U219 (N_219,N_73,N_119);
or U220 (N_220,N_115,N_174);
or U221 (N_221,N_173,N_176);
xnor U222 (N_222,In_396,In_226);
nand U223 (N_223,N_126,N_189);
xnor U224 (N_224,N_188,In_235);
nand U225 (N_225,N_74,N_171);
or U226 (N_226,N_127,N_162);
nand U227 (N_227,N_35,N_121);
nor U228 (N_228,N_185,In_299);
xnor U229 (N_229,In_434,N_130);
xnor U230 (N_230,In_305,N_138);
nor U231 (N_231,N_116,N_141);
nor U232 (N_232,In_258,In_469);
and U233 (N_233,In_54,N_55);
or U234 (N_234,In_143,N_112);
xnor U235 (N_235,In_212,N_40);
xnor U236 (N_236,In_279,In_158);
nand U237 (N_237,N_195,N_160);
and U238 (N_238,In_378,N_33);
or U239 (N_239,In_263,In_204);
or U240 (N_240,N_8,In_253);
xor U241 (N_241,In_37,N_197);
and U242 (N_242,N_1,In_30);
nand U243 (N_243,N_168,N_97);
and U244 (N_244,In_105,N_199);
or U245 (N_245,N_56,N_87);
or U246 (N_246,In_415,In_16);
or U247 (N_247,N_196,In_355);
or U248 (N_248,N_191,In_155);
nand U249 (N_249,In_256,N_21);
nand U250 (N_250,In_341,N_53);
and U251 (N_251,In_78,In_422);
or U252 (N_252,In_482,In_467);
nor U253 (N_253,In_328,N_28);
and U254 (N_254,In_79,In_398);
xnor U255 (N_255,In_185,In_358);
or U256 (N_256,In_59,In_140);
nor U257 (N_257,In_86,In_74);
or U258 (N_258,In_286,N_179);
xnor U259 (N_259,N_111,N_117);
nor U260 (N_260,In_107,N_106);
nor U261 (N_261,In_322,N_124);
xnor U262 (N_262,In_366,In_21);
xor U263 (N_263,N_10,In_448);
nor U264 (N_264,N_81,N_140);
and U265 (N_265,In_395,N_80);
nor U266 (N_266,In_471,N_82);
and U267 (N_267,In_254,In_179);
or U268 (N_268,In_440,N_88);
nand U269 (N_269,In_291,In_197);
nor U270 (N_270,N_133,N_142);
or U271 (N_271,In_233,N_165);
nor U272 (N_272,In_36,N_177);
nor U273 (N_273,In_449,In_456);
or U274 (N_274,In_283,N_92);
and U275 (N_275,N_100,N_122);
nor U276 (N_276,N_129,N_178);
nor U277 (N_277,N_152,N_108);
and U278 (N_278,In_497,N_134);
and U279 (N_279,In_123,N_180);
or U280 (N_280,In_70,N_135);
nor U281 (N_281,N_11,N_64);
nor U282 (N_282,In_152,In_496);
and U283 (N_283,In_95,N_85);
and U284 (N_284,N_48,In_39);
or U285 (N_285,In_450,N_164);
or U286 (N_286,In_386,N_167);
xor U287 (N_287,N_95,In_348);
xor U288 (N_288,N_17,In_384);
xor U289 (N_289,N_104,N_110);
or U290 (N_290,N_193,In_486);
nand U291 (N_291,N_125,N_2);
and U292 (N_292,N_187,In_478);
nand U293 (N_293,N_120,N_144);
xnor U294 (N_294,In_474,N_163);
and U295 (N_295,N_59,In_72);
and U296 (N_296,In_240,In_15);
nor U297 (N_297,In_167,N_27);
or U298 (N_298,In_266,N_154);
and U299 (N_299,N_24,In_211);
or U300 (N_300,N_29,N_292);
xnor U301 (N_301,N_265,N_143);
and U302 (N_302,N_294,N_66);
or U303 (N_303,N_90,In_248);
nand U304 (N_304,N_159,In_278);
and U305 (N_305,N_236,N_7);
and U306 (N_306,N_224,In_457);
or U307 (N_307,In_249,N_280);
nand U308 (N_308,N_298,N_219);
and U309 (N_309,N_238,N_250);
nor U310 (N_310,N_186,N_71);
nor U311 (N_311,N_260,N_245);
and U312 (N_312,N_281,In_354);
and U313 (N_313,N_175,N_184);
nor U314 (N_314,N_153,N_268);
nand U315 (N_315,N_296,N_4);
xor U316 (N_316,In_452,N_210);
and U317 (N_317,N_259,N_291);
nor U318 (N_318,N_287,N_266);
and U319 (N_319,N_286,In_402);
nand U320 (N_320,N_148,N_299);
and U321 (N_321,N_158,N_256);
or U322 (N_322,N_84,N_146);
nand U323 (N_323,N_215,In_340);
and U324 (N_324,In_148,In_5);
and U325 (N_325,N_253,In_9);
and U326 (N_326,N_262,In_294);
xnor U327 (N_327,N_113,N_271);
or U328 (N_328,In_472,N_150);
nand U329 (N_329,N_254,N_172);
xnor U330 (N_330,N_114,N_213);
and U331 (N_331,N_205,N_6);
and U332 (N_332,In_8,In_300);
nor U333 (N_333,N_293,N_63);
nand U334 (N_334,N_261,In_103);
nor U335 (N_335,N_258,N_284);
nand U336 (N_336,N_101,N_264);
xor U337 (N_337,N_70,N_45);
nand U338 (N_338,N_275,N_220);
or U339 (N_339,In_485,N_206);
or U340 (N_340,N_282,N_109);
and U341 (N_341,N_228,N_243);
or U342 (N_342,In_303,N_248);
nand U343 (N_343,N_277,N_5);
nand U344 (N_344,In_199,In_495);
nor U345 (N_345,In_173,N_239);
nand U346 (N_346,N_170,N_226);
and U347 (N_347,N_14,In_372);
or U348 (N_348,N_288,N_118);
nand U349 (N_349,In_227,N_137);
and U350 (N_350,In_151,N_169);
and U351 (N_351,N_194,In_102);
or U352 (N_352,In_285,N_214);
nor U353 (N_353,N_244,In_447);
or U354 (N_354,In_172,N_65);
or U355 (N_355,In_55,N_263);
or U356 (N_356,N_249,N_207);
nand U357 (N_357,In_334,N_225);
and U358 (N_358,N_204,N_231);
nand U359 (N_359,N_211,N_47);
xnor U360 (N_360,N_232,N_229);
and U361 (N_361,In_424,In_214);
nand U362 (N_362,N_46,N_161);
xor U363 (N_363,N_131,N_139);
nor U364 (N_364,N_41,N_276);
and U365 (N_365,In_11,N_147);
xnor U366 (N_366,N_255,N_42);
xnor U367 (N_367,In_191,N_289);
and U368 (N_368,In_401,N_252);
and U369 (N_369,N_222,N_270);
nor U370 (N_370,N_209,N_297);
nor U371 (N_371,N_269,N_273);
nand U372 (N_372,N_26,N_247);
nand U373 (N_373,In_40,N_242);
or U374 (N_374,N_272,N_251);
nand U375 (N_375,N_203,N_200);
xnor U376 (N_376,N_208,N_102);
and U377 (N_377,N_157,N_290);
or U378 (N_378,N_235,In_302);
nand U379 (N_379,N_201,N_182);
nand U380 (N_380,N_283,N_103);
nand U381 (N_381,In_311,In_427);
or U382 (N_382,N_237,In_23);
and U383 (N_383,N_218,In_33);
xor U384 (N_384,N_149,N_223);
nor U385 (N_385,In_379,N_241);
nand U386 (N_386,N_257,N_145);
or U387 (N_387,N_221,N_166);
or U388 (N_388,N_230,N_86);
nor U389 (N_389,N_278,N_240);
xor U390 (N_390,N_279,N_202);
xor U391 (N_391,N_246,In_460);
nor U392 (N_392,In_479,N_136);
nand U393 (N_393,N_267,N_233);
nor U394 (N_394,N_295,N_234);
nand U395 (N_395,N_107,N_285);
nor U396 (N_396,N_151,N_183);
nand U397 (N_397,N_274,N_216);
nor U398 (N_398,N_217,N_227);
nor U399 (N_399,In_443,N_212);
xor U400 (N_400,N_305,N_344);
or U401 (N_401,N_323,N_333);
xnor U402 (N_402,N_376,N_341);
nor U403 (N_403,N_363,N_391);
and U404 (N_404,N_368,N_335);
and U405 (N_405,N_383,N_309);
xnor U406 (N_406,N_314,N_398);
nand U407 (N_407,N_350,N_359);
nor U408 (N_408,N_393,N_311);
and U409 (N_409,N_360,N_388);
and U410 (N_410,N_394,N_380);
xnor U411 (N_411,N_358,N_349);
or U412 (N_412,N_318,N_346);
nand U413 (N_413,N_312,N_367);
and U414 (N_414,N_386,N_371);
nor U415 (N_415,N_327,N_334);
and U416 (N_416,N_307,N_362);
nand U417 (N_417,N_395,N_343);
or U418 (N_418,N_340,N_306);
nor U419 (N_419,N_373,N_399);
xor U420 (N_420,N_379,N_321);
nor U421 (N_421,N_310,N_304);
xnor U422 (N_422,N_392,N_352);
nor U423 (N_423,N_302,N_331);
xnor U424 (N_424,N_365,N_361);
nor U425 (N_425,N_315,N_336);
or U426 (N_426,N_316,N_374);
nor U427 (N_427,N_317,N_356);
or U428 (N_428,N_375,N_338);
nor U429 (N_429,N_347,N_382);
and U430 (N_430,N_329,N_326);
nand U431 (N_431,N_357,N_320);
or U432 (N_432,N_325,N_387);
nor U433 (N_433,N_337,N_313);
and U434 (N_434,N_330,N_389);
and U435 (N_435,N_369,N_364);
or U436 (N_436,N_353,N_319);
nand U437 (N_437,N_300,N_378);
and U438 (N_438,N_396,N_308);
and U439 (N_439,N_342,N_385);
or U440 (N_440,N_345,N_366);
nor U441 (N_441,N_303,N_332);
and U442 (N_442,N_354,N_372);
and U443 (N_443,N_355,N_301);
and U444 (N_444,N_339,N_377);
nor U445 (N_445,N_322,N_348);
or U446 (N_446,N_390,N_351);
and U447 (N_447,N_324,N_370);
and U448 (N_448,N_384,N_397);
or U449 (N_449,N_381,N_328);
xnor U450 (N_450,N_365,N_366);
nor U451 (N_451,N_310,N_359);
or U452 (N_452,N_303,N_335);
xor U453 (N_453,N_302,N_336);
nor U454 (N_454,N_318,N_393);
xor U455 (N_455,N_305,N_383);
xor U456 (N_456,N_346,N_308);
nor U457 (N_457,N_322,N_332);
xnor U458 (N_458,N_382,N_349);
or U459 (N_459,N_364,N_311);
xor U460 (N_460,N_375,N_343);
nor U461 (N_461,N_306,N_342);
nor U462 (N_462,N_388,N_325);
nand U463 (N_463,N_392,N_351);
or U464 (N_464,N_390,N_391);
or U465 (N_465,N_388,N_322);
xor U466 (N_466,N_354,N_381);
or U467 (N_467,N_309,N_352);
nor U468 (N_468,N_335,N_357);
or U469 (N_469,N_351,N_317);
nand U470 (N_470,N_305,N_387);
or U471 (N_471,N_370,N_342);
nor U472 (N_472,N_381,N_330);
xnor U473 (N_473,N_326,N_303);
nor U474 (N_474,N_322,N_364);
nor U475 (N_475,N_311,N_300);
or U476 (N_476,N_304,N_307);
xor U477 (N_477,N_354,N_312);
and U478 (N_478,N_395,N_333);
xor U479 (N_479,N_310,N_333);
or U480 (N_480,N_329,N_367);
nand U481 (N_481,N_338,N_326);
and U482 (N_482,N_353,N_339);
or U483 (N_483,N_343,N_342);
xor U484 (N_484,N_329,N_319);
nand U485 (N_485,N_348,N_395);
nor U486 (N_486,N_323,N_310);
xnor U487 (N_487,N_383,N_307);
or U488 (N_488,N_349,N_369);
xor U489 (N_489,N_329,N_399);
and U490 (N_490,N_374,N_371);
nand U491 (N_491,N_337,N_332);
or U492 (N_492,N_373,N_386);
nor U493 (N_493,N_365,N_334);
nor U494 (N_494,N_311,N_357);
and U495 (N_495,N_351,N_316);
or U496 (N_496,N_308,N_331);
xor U497 (N_497,N_317,N_349);
and U498 (N_498,N_331,N_373);
xnor U499 (N_499,N_347,N_376);
and U500 (N_500,N_474,N_410);
nand U501 (N_501,N_407,N_444);
xor U502 (N_502,N_429,N_478);
and U503 (N_503,N_436,N_491);
and U504 (N_504,N_488,N_499);
or U505 (N_505,N_440,N_437);
xor U506 (N_506,N_421,N_464);
nand U507 (N_507,N_489,N_459);
or U508 (N_508,N_448,N_465);
nor U509 (N_509,N_401,N_422);
or U510 (N_510,N_466,N_434);
nor U511 (N_511,N_409,N_413);
nand U512 (N_512,N_454,N_405);
and U513 (N_513,N_423,N_486);
nor U514 (N_514,N_443,N_431);
nor U515 (N_515,N_439,N_481);
or U516 (N_516,N_441,N_427);
nand U517 (N_517,N_451,N_473);
nor U518 (N_518,N_463,N_420);
nand U519 (N_519,N_417,N_406);
or U520 (N_520,N_403,N_452);
xor U521 (N_521,N_479,N_435);
or U522 (N_522,N_475,N_447);
and U523 (N_523,N_494,N_495);
or U524 (N_524,N_476,N_445);
and U525 (N_525,N_433,N_432);
and U526 (N_526,N_483,N_480);
or U527 (N_527,N_438,N_496);
xor U528 (N_528,N_484,N_446);
nor U529 (N_529,N_400,N_469);
and U530 (N_530,N_411,N_455);
or U531 (N_531,N_428,N_471);
nor U532 (N_532,N_408,N_461);
or U533 (N_533,N_467,N_424);
and U534 (N_534,N_418,N_498);
nor U535 (N_535,N_470,N_472);
or U536 (N_536,N_449,N_460);
nor U537 (N_537,N_468,N_415);
nor U538 (N_538,N_450,N_426);
or U539 (N_539,N_462,N_453);
xnor U540 (N_540,N_404,N_458);
nand U541 (N_541,N_425,N_492);
and U542 (N_542,N_493,N_430);
and U543 (N_543,N_497,N_490);
and U544 (N_544,N_482,N_412);
nand U545 (N_545,N_457,N_402);
or U546 (N_546,N_442,N_485);
or U547 (N_547,N_487,N_419);
xor U548 (N_548,N_477,N_416);
nor U549 (N_549,N_414,N_456);
nor U550 (N_550,N_428,N_476);
nor U551 (N_551,N_448,N_431);
xnor U552 (N_552,N_443,N_425);
nand U553 (N_553,N_445,N_413);
nand U554 (N_554,N_406,N_489);
xor U555 (N_555,N_497,N_458);
nand U556 (N_556,N_471,N_464);
or U557 (N_557,N_484,N_467);
nor U558 (N_558,N_432,N_440);
xnor U559 (N_559,N_456,N_432);
nor U560 (N_560,N_478,N_468);
nand U561 (N_561,N_492,N_432);
and U562 (N_562,N_486,N_412);
and U563 (N_563,N_436,N_481);
and U564 (N_564,N_470,N_480);
nand U565 (N_565,N_424,N_462);
nand U566 (N_566,N_411,N_466);
and U567 (N_567,N_455,N_429);
nand U568 (N_568,N_449,N_469);
xnor U569 (N_569,N_477,N_422);
and U570 (N_570,N_414,N_469);
nand U571 (N_571,N_481,N_434);
and U572 (N_572,N_472,N_433);
and U573 (N_573,N_439,N_454);
or U574 (N_574,N_498,N_411);
or U575 (N_575,N_498,N_496);
or U576 (N_576,N_416,N_449);
or U577 (N_577,N_401,N_488);
nor U578 (N_578,N_423,N_470);
nand U579 (N_579,N_426,N_472);
nor U580 (N_580,N_489,N_421);
nand U581 (N_581,N_430,N_464);
and U582 (N_582,N_446,N_419);
nor U583 (N_583,N_455,N_440);
xor U584 (N_584,N_473,N_462);
xnor U585 (N_585,N_495,N_401);
or U586 (N_586,N_430,N_478);
nor U587 (N_587,N_435,N_451);
nand U588 (N_588,N_405,N_408);
nand U589 (N_589,N_466,N_412);
nand U590 (N_590,N_457,N_426);
and U591 (N_591,N_476,N_493);
nor U592 (N_592,N_497,N_473);
and U593 (N_593,N_450,N_486);
nor U594 (N_594,N_422,N_408);
nor U595 (N_595,N_435,N_477);
and U596 (N_596,N_475,N_430);
and U597 (N_597,N_431,N_404);
nand U598 (N_598,N_412,N_436);
or U599 (N_599,N_422,N_426);
or U600 (N_600,N_553,N_509);
and U601 (N_601,N_508,N_575);
or U602 (N_602,N_501,N_511);
nand U603 (N_603,N_535,N_523);
nand U604 (N_604,N_549,N_518);
or U605 (N_605,N_510,N_522);
and U606 (N_606,N_583,N_591);
nand U607 (N_607,N_587,N_557);
xor U608 (N_608,N_520,N_547);
nand U609 (N_609,N_590,N_565);
or U610 (N_610,N_505,N_574);
xnor U611 (N_611,N_585,N_526);
xor U612 (N_612,N_592,N_516);
nor U613 (N_613,N_532,N_570);
nand U614 (N_614,N_546,N_515);
nand U615 (N_615,N_559,N_502);
and U616 (N_616,N_576,N_530);
nand U617 (N_617,N_588,N_512);
or U618 (N_618,N_527,N_598);
xnor U619 (N_619,N_524,N_536);
and U620 (N_620,N_533,N_582);
or U621 (N_621,N_504,N_573);
or U622 (N_622,N_566,N_596);
xor U623 (N_623,N_593,N_599);
or U624 (N_624,N_552,N_572);
or U625 (N_625,N_589,N_556);
or U626 (N_626,N_514,N_537);
or U627 (N_627,N_525,N_554);
xor U628 (N_628,N_544,N_519);
nor U629 (N_629,N_595,N_540);
nand U630 (N_630,N_564,N_577);
nor U631 (N_631,N_586,N_594);
xnor U632 (N_632,N_571,N_563);
or U633 (N_633,N_528,N_597);
nor U634 (N_634,N_506,N_580);
nand U635 (N_635,N_567,N_569);
or U636 (N_636,N_560,N_578);
nand U637 (N_637,N_555,N_534);
nand U638 (N_638,N_545,N_579);
nand U639 (N_639,N_551,N_507);
or U640 (N_640,N_531,N_503);
or U641 (N_641,N_541,N_568);
or U642 (N_642,N_558,N_543);
and U643 (N_643,N_517,N_561);
nor U644 (N_644,N_521,N_538);
xor U645 (N_645,N_550,N_529);
xor U646 (N_646,N_581,N_539);
nor U647 (N_647,N_513,N_584);
xor U648 (N_648,N_542,N_500);
and U649 (N_649,N_562,N_548);
and U650 (N_650,N_577,N_553);
or U651 (N_651,N_508,N_568);
xor U652 (N_652,N_589,N_515);
nand U653 (N_653,N_589,N_513);
or U654 (N_654,N_510,N_582);
nand U655 (N_655,N_538,N_535);
nand U656 (N_656,N_568,N_534);
and U657 (N_657,N_501,N_550);
and U658 (N_658,N_507,N_517);
and U659 (N_659,N_537,N_595);
and U660 (N_660,N_553,N_534);
and U661 (N_661,N_576,N_510);
xor U662 (N_662,N_586,N_516);
xor U663 (N_663,N_545,N_540);
nand U664 (N_664,N_523,N_529);
or U665 (N_665,N_533,N_598);
xor U666 (N_666,N_522,N_502);
nor U667 (N_667,N_526,N_521);
nor U668 (N_668,N_513,N_542);
and U669 (N_669,N_544,N_526);
or U670 (N_670,N_528,N_554);
nand U671 (N_671,N_568,N_575);
nand U672 (N_672,N_552,N_567);
xnor U673 (N_673,N_581,N_546);
nor U674 (N_674,N_507,N_510);
and U675 (N_675,N_579,N_503);
nor U676 (N_676,N_574,N_548);
xnor U677 (N_677,N_517,N_599);
xnor U678 (N_678,N_525,N_504);
and U679 (N_679,N_504,N_571);
and U680 (N_680,N_528,N_563);
nor U681 (N_681,N_596,N_565);
nand U682 (N_682,N_598,N_536);
nand U683 (N_683,N_518,N_542);
nand U684 (N_684,N_591,N_506);
nand U685 (N_685,N_507,N_575);
and U686 (N_686,N_566,N_546);
or U687 (N_687,N_512,N_598);
nand U688 (N_688,N_558,N_508);
xnor U689 (N_689,N_586,N_571);
nand U690 (N_690,N_515,N_557);
xor U691 (N_691,N_512,N_516);
nor U692 (N_692,N_500,N_584);
and U693 (N_693,N_513,N_575);
nor U694 (N_694,N_524,N_566);
and U695 (N_695,N_591,N_565);
or U696 (N_696,N_576,N_599);
xnor U697 (N_697,N_529,N_543);
xnor U698 (N_698,N_505,N_508);
nor U699 (N_699,N_592,N_581);
xor U700 (N_700,N_686,N_655);
xnor U701 (N_701,N_691,N_690);
and U702 (N_702,N_696,N_638);
nand U703 (N_703,N_615,N_600);
and U704 (N_704,N_632,N_664);
xnor U705 (N_705,N_611,N_656);
and U706 (N_706,N_614,N_604);
nand U707 (N_707,N_616,N_606);
nor U708 (N_708,N_646,N_640);
nor U709 (N_709,N_676,N_670);
nor U710 (N_710,N_637,N_692);
nor U711 (N_711,N_624,N_659);
nand U712 (N_712,N_663,N_660);
or U713 (N_713,N_650,N_672);
and U714 (N_714,N_643,N_662);
nand U715 (N_715,N_657,N_688);
nand U716 (N_716,N_620,N_648);
and U717 (N_717,N_694,N_678);
and U718 (N_718,N_673,N_684);
nand U719 (N_719,N_639,N_601);
nor U720 (N_720,N_693,N_661);
and U721 (N_721,N_608,N_658);
nand U722 (N_722,N_609,N_679);
nand U723 (N_723,N_677,N_607);
nor U724 (N_724,N_625,N_644);
nor U725 (N_725,N_698,N_634);
nor U726 (N_726,N_633,N_618);
xor U727 (N_727,N_699,N_605);
and U728 (N_728,N_675,N_668);
nor U729 (N_729,N_645,N_610);
and U730 (N_730,N_681,N_683);
xnor U731 (N_731,N_623,N_619);
and U732 (N_732,N_630,N_667);
nor U733 (N_733,N_666,N_636);
or U734 (N_734,N_629,N_682);
nor U735 (N_735,N_680,N_695);
nor U736 (N_736,N_647,N_649);
nand U737 (N_737,N_617,N_674);
or U738 (N_738,N_603,N_652);
or U739 (N_739,N_627,N_669);
nand U740 (N_740,N_665,N_635);
or U741 (N_741,N_612,N_628);
nand U742 (N_742,N_653,N_641);
and U743 (N_743,N_689,N_651);
nor U744 (N_744,N_626,N_621);
nor U745 (N_745,N_654,N_697);
nor U746 (N_746,N_687,N_631);
nand U747 (N_747,N_622,N_685);
nor U748 (N_748,N_671,N_642);
and U749 (N_749,N_613,N_602);
and U750 (N_750,N_694,N_693);
or U751 (N_751,N_618,N_661);
nor U752 (N_752,N_690,N_645);
or U753 (N_753,N_663,N_647);
nor U754 (N_754,N_654,N_698);
xor U755 (N_755,N_617,N_633);
nor U756 (N_756,N_644,N_688);
or U757 (N_757,N_610,N_609);
nor U758 (N_758,N_644,N_652);
nor U759 (N_759,N_613,N_669);
and U760 (N_760,N_657,N_653);
nor U761 (N_761,N_629,N_693);
or U762 (N_762,N_645,N_678);
or U763 (N_763,N_617,N_634);
xor U764 (N_764,N_647,N_650);
nor U765 (N_765,N_639,N_691);
or U766 (N_766,N_632,N_683);
or U767 (N_767,N_612,N_699);
nand U768 (N_768,N_681,N_648);
nand U769 (N_769,N_639,N_636);
xor U770 (N_770,N_663,N_661);
and U771 (N_771,N_630,N_663);
nor U772 (N_772,N_630,N_614);
and U773 (N_773,N_626,N_638);
xnor U774 (N_774,N_672,N_628);
and U775 (N_775,N_681,N_604);
nor U776 (N_776,N_676,N_666);
nand U777 (N_777,N_611,N_621);
xnor U778 (N_778,N_604,N_679);
nor U779 (N_779,N_691,N_616);
xnor U780 (N_780,N_677,N_691);
or U781 (N_781,N_698,N_689);
or U782 (N_782,N_637,N_609);
or U783 (N_783,N_677,N_665);
nand U784 (N_784,N_628,N_693);
or U785 (N_785,N_670,N_645);
nand U786 (N_786,N_670,N_650);
nor U787 (N_787,N_672,N_611);
or U788 (N_788,N_605,N_631);
nor U789 (N_789,N_622,N_688);
and U790 (N_790,N_651,N_628);
nor U791 (N_791,N_645,N_646);
nand U792 (N_792,N_645,N_613);
and U793 (N_793,N_640,N_658);
and U794 (N_794,N_632,N_630);
or U795 (N_795,N_616,N_659);
nor U796 (N_796,N_624,N_633);
nand U797 (N_797,N_608,N_677);
nand U798 (N_798,N_660,N_620);
nand U799 (N_799,N_651,N_605);
nand U800 (N_800,N_786,N_705);
xor U801 (N_801,N_783,N_763);
xor U802 (N_802,N_730,N_714);
nand U803 (N_803,N_794,N_773);
nand U804 (N_804,N_781,N_785);
nand U805 (N_805,N_702,N_784);
or U806 (N_806,N_733,N_772);
and U807 (N_807,N_721,N_738);
xnor U808 (N_808,N_707,N_777);
nand U809 (N_809,N_710,N_704);
or U810 (N_810,N_731,N_766);
nand U811 (N_811,N_797,N_750);
and U812 (N_812,N_729,N_752);
and U813 (N_813,N_728,N_759);
or U814 (N_814,N_734,N_753);
and U815 (N_815,N_740,N_780);
nor U816 (N_816,N_723,N_761);
xnor U817 (N_817,N_736,N_767);
or U818 (N_818,N_722,N_748);
xnor U819 (N_819,N_700,N_737);
xor U820 (N_820,N_727,N_788);
and U821 (N_821,N_717,N_711);
nand U822 (N_822,N_713,N_755);
xnor U823 (N_823,N_732,N_745);
nor U824 (N_824,N_739,N_743);
and U825 (N_825,N_703,N_776);
nand U826 (N_826,N_792,N_770);
nor U827 (N_827,N_760,N_757);
nor U828 (N_828,N_706,N_768);
xnor U829 (N_829,N_712,N_774);
nand U830 (N_830,N_762,N_756);
nand U831 (N_831,N_720,N_741);
or U832 (N_832,N_726,N_769);
or U833 (N_833,N_790,N_791);
xor U834 (N_834,N_758,N_795);
nand U835 (N_835,N_798,N_735);
and U836 (N_836,N_708,N_782);
or U837 (N_837,N_749,N_751);
nor U838 (N_838,N_725,N_718);
or U839 (N_839,N_715,N_719);
or U840 (N_840,N_793,N_724);
and U841 (N_841,N_765,N_742);
xor U842 (N_842,N_775,N_754);
nand U843 (N_843,N_764,N_701);
or U844 (N_844,N_716,N_796);
or U845 (N_845,N_709,N_787);
or U846 (N_846,N_778,N_799);
xor U847 (N_847,N_746,N_744);
and U848 (N_848,N_779,N_789);
xor U849 (N_849,N_771,N_747);
or U850 (N_850,N_738,N_720);
nand U851 (N_851,N_782,N_765);
and U852 (N_852,N_713,N_754);
and U853 (N_853,N_741,N_778);
and U854 (N_854,N_742,N_783);
nand U855 (N_855,N_723,N_799);
and U856 (N_856,N_739,N_799);
xnor U857 (N_857,N_750,N_791);
and U858 (N_858,N_721,N_754);
or U859 (N_859,N_772,N_786);
nor U860 (N_860,N_746,N_707);
nor U861 (N_861,N_786,N_778);
nor U862 (N_862,N_708,N_719);
or U863 (N_863,N_701,N_731);
xnor U864 (N_864,N_795,N_715);
nor U865 (N_865,N_775,N_758);
or U866 (N_866,N_733,N_796);
xor U867 (N_867,N_797,N_740);
nand U868 (N_868,N_729,N_748);
or U869 (N_869,N_798,N_732);
and U870 (N_870,N_737,N_781);
and U871 (N_871,N_706,N_746);
nor U872 (N_872,N_791,N_756);
or U873 (N_873,N_718,N_756);
nor U874 (N_874,N_774,N_786);
and U875 (N_875,N_715,N_704);
nor U876 (N_876,N_706,N_718);
and U877 (N_877,N_719,N_755);
nand U878 (N_878,N_735,N_785);
xnor U879 (N_879,N_761,N_717);
xnor U880 (N_880,N_772,N_771);
and U881 (N_881,N_761,N_770);
nand U882 (N_882,N_754,N_734);
and U883 (N_883,N_711,N_706);
and U884 (N_884,N_752,N_794);
nand U885 (N_885,N_766,N_770);
nand U886 (N_886,N_764,N_759);
nor U887 (N_887,N_759,N_710);
nand U888 (N_888,N_775,N_719);
or U889 (N_889,N_789,N_757);
nand U890 (N_890,N_724,N_767);
nand U891 (N_891,N_707,N_790);
xor U892 (N_892,N_718,N_734);
or U893 (N_893,N_775,N_774);
xnor U894 (N_894,N_724,N_745);
nor U895 (N_895,N_711,N_769);
nand U896 (N_896,N_795,N_775);
and U897 (N_897,N_769,N_760);
xor U898 (N_898,N_722,N_730);
and U899 (N_899,N_757,N_744);
nor U900 (N_900,N_819,N_822);
and U901 (N_901,N_866,N_843);
and U902 (N_902,N_886,N_853);
or U903 (N_903,N_844,N_807);
xor U904 (N_904,N_802,N_829);
nor U905 (N_905,N_860,N_839);
nand U906 (N_906,N_867,N_889);
or U907 (N_907,N_821,N_808);
nand U908 (N_908,N_888,N_837);
nand U909 (N_909,N_803,N_817);
nand U910 (N_910,N_830,N_818);
xnor U911 (N_911,N_873,N_845);
xor U912 (N_912,N_898,N_892);
nand U913 (N_913,N_893,N_855);
and U914 (N_914,N_884,N_850);
nand U915 (N_915,N_864,N_813);
and U916 (N_916,N_896,N_824);
nor U917 (N_917,N_861,N_871);
or U918 (N_918,N_833,N_805);
or U919 (N_919,N_878,N_854);
and U920 (N_920,N_828,N_852);
and U921 (N_921,N_868,N_801);
and U922 (N_922,N_816,N_827);
nor U923 (N_923,N_863,N_823);
and U924 (N_924,N_879,N_831);
and U925 (N_925,N_851,N_848);
nor U926 (N_926,N_842,N_810);
nor U927 (N_927,N_869,N_815);
nor U928 (N_928,N_804,N_847);
nor U929 (N_929,N_800,N_826);
or U930 (N_930,N_874,N_858);
xnor U931 (N_931,N_887,N_806);
nand U932 (N_932,N_877,N_881);
and U933 (N_933,N_885,N_840);
nand U934 (N_934,N_891,N_836);
and U935 (N_935,N_890,N_820);
or U936 (N_936,N_834,N_838);
and U937 (N_937,N_865,N_832);
nor U938 (N_938,N_882,N_835);
and U939 (N_939,N_811,N_862);
nand U940 (N_940,N_857,N_846);
nor U941 (N_941,N_809,N_895);
xnor U942 (N_942,N_841,N_814);
nor U943 (N_943,N_872,N_859);
or U944 (N_944,N_880,N_856);
nand U945 (N_945,N_812,N_876);
nor U946 (N_946,N_899,N_849);
nor U947 (N_947,N_825,N_870);
and U948 (N_948,N_875,N_897);
xnor U949 (N_949,N_883,N_894);
nor U950 (N_950,N_847,N_814);
nand U951 (N_951,N_868,N_840);
and U952 (N_952,N_828,N_870);
and U953 (N_953,N_806,N_862);
or U954 (N_954,N_871,N_895);
and U955 (N_955,N_856,N_861);
or U956 (N_956,N_887,N_875);
and U957 (N_957,N_801,N_857);
or U958 (N_958,N_884,N_877);
xor U959 (N_959,N_868,N_843);
nor U960 (N_960,N_858,N_833);
xnor U961 (N_961,N_881,N_846);
xnor U962 (N_962,N_872,N_884);
nor U963 (N_963,N_801,N_893);
or U964 (N_964,N_862,N_827);
nor U965 (N_965,N_856,N_891);
or U966 (N_966,N_865,N_889);
or U967 (N_967,N_893,N_888);
or U968 (N_968,N_854,N_834);
and U969 (N_969,N_845,N_885);
and U970 (N_970,N_840,N_847);
nor U971 (N_971,N_819,N_809);
nand U972 (N_972,N_871,N_809);
and U973 (N_973,N_885,N_863);
nand U974 (N_974,N_806,N_832);
or U975 (N_975,N_860,N_819);
and U976 (N_976,N_862,N_886);
xnor U977 (N_977,N_868,N_880);
xnor U978 (N_978,N_839,N_885);
xnor U979 (N_979,N_814,N_813);
nand U980 (N_980,N_861,N_870);
nor U981 (N_981,N_808,N_875);
and U982 (N_982,N_818,N_860);
nand U983 (N_983,N_844,N_860);
xnor U984 (N_984,N_833,N_824);
nor U985 (N_985,N_840,N_811);
or U986 (N_986,N_896,N_872);
or U987 (N_987,N_855,N_805);
and U988 (N_988,N_810,N_836);
or U989 (N_989,N_834,N_820);
or U990 (N_990,N_889,N_868);
xor U991 (N_991,N_870,N_854);
nand U992 (N_992,N_869,N_824);
nor U993 (N_993,N_827,N_844);
nor U994 (N_994,N_867,N_841);
nor U995 (N_995,N_876,N_886);
and U996 (N_996,N_895,N_887);
and U997 (N_997,N_891,N_819);
xor U998 (N_998,N_897,N_891);
and U999 (N_999,N_861,N_830);
nand U1000 (N_1000,N_972,N_987);
xnor U1001 (N_1001,N_904,N_927);
and U1002 (N_1002,N_981,N_914);
and U1003 (N_1003,N_996,N_984);
nand U1004 (N_1004,N_922,N_994);
nand U1005 (N_1005,N_946,N_962);
and U1006 (N_1006,N_918,N_932);
or U1007 (N_1007,N_977,N_907);
xnor U1008 (N_1008,N_934,N_967);
and U1009 (N_1009,N_989,N_986);
nand U1010 (N_1010,N_917,N_957);
or U1011 (N_1011,N_910,N_963);
nor U1012 (N_1012,N_905,N_935);
xor U1013 (N_1013,N_919,N_945);
xor U1014 (N_1014,N_969,N_951);
nand U1015 (N_1015,N_901,N_906);
nor U1016 (N_1016,N_953,N_915);
nor U1017 (N_1017,N_909,N_990);
and U1018 (N_1018,N_959,N_955);
nand U1019 (N_1019,N_924,N_936);
or U1020 (N_1020,N_949,N_960);
and U1021 (N_1021,N_903,N_913);
and U1022 (N_1022,N_985,N_937);
nor U1023 (N_1023,N_908,N_999);
xnor U1024 (N_1024,N_980,N_968);
nor U1025 (N_1025,N_966,N_964);
and U1026 (N_1026,N_973,N_954);
nor U1027 (N_1027,N_979,N_912);
nor U1028 (N_1028,N_952,N_998);
and U1029 (N_1029,N_961,N_900);
and U1030 (N_1030,N_995,N_975);
nor U1031 (N_1031,N_911,N_939);
nor U1032 (N_1032,N_926,N_974);
and U1033 (N_1033,N_993,N_971);
nor U1034 (N_1034,N_965,N_978);
xor U1035 (N_1035,N_930,N_938);
nand U1036 (N_1036,N_931,N_916);
nor U1037 (N_1037,N_923,N_943);
or U1038 (N_1038,N_983,N_941);
and U1039 (N_1039,N_970,N_942);
nor U1040 (N_1040,N_948,N_940);
and U1041 (N_1041,N_997,N_982);
xor U1042 (N_1042,N_950,N_991);
nand U1043 (N_1043,N_944,N_929);
or U1044 (N_1044,N_925,N_920);
nand U1045 (N_1045,N_958,N_928);
xnor U1046 (N_1046,N_947,N_976);
xnor U1047 (N_1047,N_902,N_988);
xor U1048 (N_1048,N_933,N_992);
xnor U1049 (N_1049,N_956,N_921);
xor U1050 (N_1050,N_945,N_985);
xnor U1051 (N_1051,N_949,N_990);
or U1052 (N_1052,N_948,N_908);
xor U1053 (N_1053,N_977,N_924);
xnor U1054 (N_1054,N_902,N_930);
xnor U1055 (N_1055,N_973,N_924);
and U1056 (N_1056,N_925,N_909);
nand U1057 (N_1057,N_927,N_913);
nor U1058 (N_1058,N_940,N_946);
or U1059 (N_1059,N_942,N_933);
and U1060 (N_1060,N_993,N_976);
xnor U1061 (N_1061,N_923,N_901);
xnor U1062 (N_1062,N_938,N_964);
and U1063 (N_1063,N_913,N_962);
nor U1064 (N_1064,N_955,N_928);
and U1065 (N_1065,N_904,N_985);
and U1066 (N_1066,N_964,N_973);
xor U1067 (N_1067,N_949,N_905);
nor U1068 (N_1068,N_969,N_907);
or U1069 (N_1069,N_946,N_927);
nor U1070 (N_1070,N_937,N_923);
and U1071 (N_1071,N_939,N_975);
nand U1072 (N_1072,N_939,N_993);
xor U1073 (N_1073,N_980,N_971);
nand U1074 (N_1074,N_946,N_936);
or U1075 (N_1075,N_949,N_917);
nor U1076 (N_1076,N_993,N_921);
and U1077 (N_1077,N_931,N_963);
xor U1078 (N_1078,N_953,N_992);
and U1079 (N_1079,N_909,N_958);
or U1080 (N_1080,N_958,N_926);
and U1081 (N_1081,N_984,N_974);
nand U1082 (N_1082,N_903,N_988);
or U1083 (N_1083,N_911,N_914);
or U1084 (N_1084,N_907,N_972);
or U1085 (N_1085,N_948,N_937);
or U1086 (N_1086,N_995,N_960);
nor U1087 (N_1087,N_911,N_976);
or U1088 (N_1088,N_979,N_951);
nor U1089 (N_1089,N_997,N_957);
or U1090 (N_1090,N_989,N_972);
nor U1091 (N_1091,N_969,N_903);
and U1092 (N_1092,N_993,N_986);
nor U1093 (N_1093,N_982,N_909);
nor U1094 (N_1094,N_937,N_911);
nand U1095 (N_1095,N_909,N_926);
nor U1096 (N_1096,N_939,N_908);
xor U1097 (N_1097,N_954,N_984);
and U1098 (N_1098,N_932,N_999);
nand U1099 (N_1099,N_925,N_911);
xnor U1100 (N_1100,N_1013,N_1033);
nor U1101 (N_1101,N_1054,N_1041);
or U1102 (N_1102,N_1071,N_1068);
or U1103 (N_1103,N_1015,N_1060);
or U1104 (N_1104,N_1052,N_1046);
or U1105 (N_1105,N_1094,N_1045);
or U1106 (N_1106,N_1049,N_1004);
and U1107 (N_1107,N_1081,N_1069);
nor U1108 (N_1108,N_1036,N_1072);
nand U1109 (N_1109,N_1055,N_1024);
nand U1110 (N_1110,N_1028,N_1035);
or U1111 (N_1111,N_1043,N_1014);
nand U1112 (N_1112,N_1002,N_1018);
or U1113 (N_1113,N_1077,N_1078);
xor U1114 (N_1114,N_1001,N_1074);
xnor U1115 (N_1115,N_1087,N_1047);
nand U1116 (N_1116,N_1017,N_1065);
or U1117 (N_1117,N_1029,N_1097);
nor U1118 (N_1118,N_1032,N_1010);
xor U1119 (N_1119,N_1062,N_1022);
xor U1120 (N_1120,N_1009,N_1040);
and U1121 (N_1121,N_1005,N_1067);
nand U1122 (N_1122,N_1053,N_1020);
and U1123 (N_1123,N_1099,N_1063);
nand U1124 (N_1124,N_1012,N_1042);
nand U1125 (N_1125,N_1057,N_1089);
nand U1126 (N_1126,N_1076,N_1023);
xnor U1127 (N_1127,N_1037,N_1085);
xor U1128 (N_1128,N_1079,N_1050);
and U1129 (N_1129,N_1048,N_1030);
nor U1130 (N_1130,N_1066,N_1006);
nand U1131 (N_1131,N_1026,N_1008);
nor U1132 (N_1132,N_1083,N_1091);
and U1133 (N_1133,N_1088,N_1059);
xnor U1134 (N_1134,N_1092,N_1003);
xor U1135 (N_1135,N_1031,N_1007);
or U1136 (N_1136,N_1090,N_1093);
xnor U1137 (N_1137,N_1051,N_1080);
xor U1138 (N_1138,N_1082,N_1000);
xnor U1139 (N_1139,N_1056,N_1039);
nand U1140 (N_1140,N_1058,N_1061);
nor U1141 (N_1141,N_1019,N_1011);
xnor U1142 (N_1142,N_1095,N_1038);
nor U1143 (N_1143,N_1070,N_1025);
nand U1144 (N_1144,N_1064,N_1075);
nand U1145 (N_1145,N_1098,N_1096);
nor U1146 (N_1146,N_1034,N_1073);
xnor U1147 (N_1147,N_1086,N_1027);
or U1148 (N_1148,N_1084,N_1021);
or U1149 (N_1149,N_1016,N_1044);
and U1150 (N_1150,N_1058,N_1057);
xor U1151 (N_1151,N_1013,N_1036);
nor U1152 (N_1152,N_1076,N_1086);
nand U1153 (N_1153,N_1026,N_1046);
or U1154 (N_1154,N_1000,N_1022);
nor U1155 (N_1155,N_1063,N_1013);
or U1156 (N_1156,N_1065,N_1067);
nor U1157 (N_1157,N_1093,N_1025);
xor U1158 (N_1158,N_1020,N_1009);
and U1159 (N_1159,N_1038,N_1079);
nor U1160 (N_1160,N_1013,N_1024);
and U1161 (N_1161,N_1088,N_1009);
nor U1162 (N_1162,N_1034,N_1068);
xnor U1163 (N_1163,N_1073,N_1075);
xnor U1164 (N_1164,N_1090,N_1015);
or U1165 (N_1165,N_1090,N_1065);
nor U1166 (N_1166,N_1080,N_1077);
or U1167 (N_1167,N_1086,N_1042);
xor U1168 (N_1168,N_1071,N_1004);
nand U1169 (N_1169,N_1001,N_1066);
and U1170 (N_1170,N_1072,N_1049);
nand U1171 (N_1171,N_1070,N_1055);
and U1172 (N_1172,N_1004,N_1031);
nor U1173 (N_1173,N_1074,N_1025);
xnor U1174 (N_1174,N_1040,N_1047);
nand U1175 (N_1175,N_1072,N_1032);
or U1176 (N_1176,N_1006,N_1061);
or U1177 (N_1177,N_1084,N_1094);
nor U1178 (N_1178,N_1058,N_1045);
nand U1179 (N_1179,N_1074,N_1063);
or U1180 (N_1180,N_1011,N_1048);
nor U1181 (N_1181,N_1040,N_1086);
or U1182 (N_1182,N_1050,N_1062);
nand U1183 (N_1183,N_1088,N_1083);
xnor U1184 (N_1184,N_1003,N_1052);
nor U1185 (N_1185,N_1006,N_1075);
and U1186 (N_1186,N_1024,N_1046);
nor U1187 (N_1187,N_1027,N_1070);
or U1188 (N_1188,N_1041,N_1076);
or U1189 (N_1189,N_1080,N_1019);
xnor U1190 (N_1190,N_1018,N_1027);
or U1191 (N_1191,N_1020,N_1090);
nor U1192 (N_1192,N_1044,N_1047);
nand U1193 (N_1193,N_1011,N_1089);
or U1194 (N_1194,N_1088,N_1024);
nand U1195 (N_1195,N_1013,N_1022);
nand U1196 (N_1196,N_1006,N_1099);
and U1197 (N_1197,N_1012,N_1021);
nor U1198 (N_1198,N_1072,N_1057);
xor U1199 (N_1199,N_1082,N_1047);
nor U1200 (N_1200,N_1127,N_1162);
xor U1201 (N_1201,N_1164,N_1152);
nor U1202 (N_1202,N_1194,N_1193);
or U1203 (N_1203,N_1176,N_1178);
xor U1204 (N_1204,N_1159,N_1143);
and U1205 (N_1205,N_1180,N_1168);
or U1206 (N_1206,N_1120,N_1187);
xor U1207 (N_1207,N_1139,N_1109);
nor U1208 (N_1208,N_1161,N_1190);
or U1209 (N_1209,N_1101,N_1107);
or U1210 (N_1210,N_1185,N_1163);
nand U1211 (N_1211,N_1170,N_1150);
and U1212 (N_1212,N_1175,N_1141);
nand U1213 (N_1213,N_1145,N_1166);
nand U1214 (N_1214,N_1156,N_1124);
and U1215 (N_1215,N_1137,N_1113);
or U1216 (N_1216,N_1181,N_1119);
or U1217 (N_1217,N_1174,N_1177);
xor U1218 (N_1218,N_1192,N_1135);
or U1219 (N_1219,N_1146,N_1165);
and U1220 (N_1220,N_1167,N_1188);
nand U1221 (N_1221,N_1140,N_1102);
xnor U1222 (N_1222,N_1136,N_1142);
xor U1223 (N_1223,N_1184,N_1171);
nand U1224 (N_1224,N_1198,N_1173);
nor U1225 (N_1225,N_1155,N_1125);
or U1226 (N_1226,N_1104,N_1129);
and U1227 (N_1227,N_1121,N_1189);
and U1228 (N_1228,N_1115,N_1112);
or U1229 (N_1229,N_1144,N_1103);
and U1230 (N_1230,N_1108,N_1130);
xor U1231 (N_1231,N_1138,N_1122);
xor U1232 (N_1232,N_1154,N_1105);
nor U1233 (N_1233,N_1183,N_1117);
and U1234 (N_1234,N_1172,N_1100);
or U1235 (N_1235,N_1182,N_1158);
and U1236 (N_1236,N_1186,N_1126);
nor U1237 (N_1237,N_1153,N_1132);
or U1238 (N_1238,N_1191,N_1160);
or U1239 (N_1239,N_1196,N_1111);
nand U1240 (N_1240,N_1128,N_1195);
and U1241 (N_1241,N_1199,N_1157);
xor U1242 (N_1242,N_1110,N_1197);
nand U1243 (N_1243,N_1114,N_1169);
and U1244 (N_1244,N_1148,N_1133);
nor U1245 (N_1245,N_1118,N_1116);
or U1246 (N_1246,N_1147,N_1151);
xnor U1247 (N_1247,N_1123,N_1149);
and U1248 (N_1248,N_1179,N_1131);
nand U1249 (N_1249,N_1134,N_1106);
nor U1250 (N_1250,N_1188,N_1117);
or U1251 (N_1251,N_1111,N_1112);
nand U1252 (N_1252,N_1148,N_1150);
or U1253 (N_1253,N_1154,N_1151);
nand U1254 (N_1254,N_1142,N_1116);
or U1255 (N_1255,N_1146,N_1128);
nor U1256 (N_1256,N_1140,N_1115);
and U1257 (N_1257,N_1159,N_1160);
and U1258 (N_1258,N_1102,N_1192);
and U1259 (N_1259,N_1129,N_1145);
and U1260 (N_1260,N_1192,N_1147);
or U1261 (N_1261,N_1177,N_1142);
nor U1262 (N_1262,N_1177,N_1141);
or U1263 (N_1263,N_1130,N_1145);
and U1264 (N_1264,N_1139,N_1169);
nor U1265 (N_1265,N_1187,N_1103);
or U1266 (N_1266,N_1163,N_1169);
and U1267 (N_1267,N_1102,N_1104);
or U1268 (N_1268,N_1132,N_1140);
xnor U1269 (N_1269,N_1178,N_1121);
xor U1270 (N_1270,N_1112,N_1184);
or U1271 (N_1271,N_1153,N_1183);
nor U1272 (N_1272,N_1137,N_1166);
nand U1273 (N_1273,N_1101,N_1142);
or U1274 (N_1274,N_1104,N_1143);
nand U1275 (N_1275,N_1162,N_1184);
nand U1276 (N_1276,N_1153,N_1113);
and U1277 (N_1277,N_1135,N_1103);
xnor U1278 (N_1278,N_1166,N_1143);
nand U1279 (N_1279,N_1169,N_1135);
nor U1280 (N_1280,N_1191,N_1130);
nand U1281 (N_1281,N_1160,N_1171);
and U1282 (N_1282,N_1109,N_1170);
and U1283 (N_1283,N_1152,N_1163);
nor U1284 (N_1284,N_1148,N_1144);
nand U1285 (N_1285,N_1188,N_1106);
nand U1286 (N_1286,N_1150,N_1144);
and U1287 (N_1287,N_1118,N_1188);
and U1288 (N_1288,N_1129,N_1176);
nor U1289 (N_1289,N_1134,N_1175);
nor U1290 (N_1290,N_1141,N_1134);
xor U1291 (N_1291,N_1162,N_1181);
nor U1292 (N_1292,N_1162,N_1179);
and U1293 (N_1293,N_1133,N_1153);
nor U1294 (N_1294,N_1112,N_1174);
xor U1295 (N_1295,N_1162,N_1189);
xor U1296 (N_1296,N_1147,N_1118);
nand U1297 (N_1297,N_1149,N_1134);
nor U1298 (N_1298,N_1178,N_1173);
and U1299 (N_1299,N_1192,N_1158);
nor U1300 (N_1300,N_1227,N_1268);
or U1301 (N_1301,N_1200,N_1242);
xor U1302 (N_1302,N_1224,N_1245);
or U1303 (N_1303,N_1221,N_1218);
or U1304 (N_1304,N_1267,N_1289);
nor U1305 (N_1305,N_1209,N_1231);
nor U1306 (N_1306,N_1222,N_1276);
and U1307 (N_1307,N_1219,N_1240);
nor U1308 (N_1308,N_1207,N_1212);
and U1309 (N_1309,N_1249,N_1297);
nor U1310 (N_1310,N_1243,N_1256);
or U1311 (N_1311,N_1283,N_1262);
nor U1312 (N_1312,N_1287,N_1248);
and U1313 (N_1313,N_1239,N_1295);
or U1314 (N_1314,N_1238,N_1216);
and U1315 (N_1315,N_1281,N_1255);
or U1316 (N_1316,N_1241,N_1223);
xnor U1317 (N_1317,N_1251,N_1217);
nand U1318 (N_1318,N_1298,N_1271);
and U1319 (N_1319,N_1253,N_1205);
nand U1320 (N_1320,N_1277,N_1229);
nor U1321 (N_1321,N_1265,N_1254);
xor U1322 (N_1322,N_1233,N_1269);
nor U1323 (N_1323,N_1213,N_1291);
xnor U1324 (N_1324,N_1234,N_1236);
nand U1325 (N_1325,N_1208,N_1203);
or U1326 (N_1326,N_1237,N_1292);
or U1327 (N_1327,N_1278,N_1204);
nor U1328 (N_1328,N_1299,N_1293);
nor U1329 (N_1329,N_1275,N_1294);
xor U1330 (N_1330,N_1272,N_1211);
nand U1331 (N_1331,N_1257,N_1220);
or U1332 (N_1332,N_1246,N_1206);
and U1333 (N_1333,N_1201,N_1279);
nor U1334 (N_1334,N_1230,N_1270);
xor U1335 (N_1335,N_1226,N_1252);
nand U1336 (N_1336,N_1296,N_1286);
and U1337 (N_1337,N_1228,N_1282);
and U1338 (N_1338,N_1261,N_1288);
nand U1339 (N_1339,N_1274,N_1264);
nand U1340 (N_1340,N_1235,N_1290);
xnor U1341 (N_1341,N_1266,N_1225);
nand U1342 (N_1342,N_1258,N_1259);
or U1343 (N_1343,N_1202,N_1214);
or U1344 (N_1344,N_1232,N_1285);
or U1345 (N_1345,N_1244,N_1284);
nand U1346 (N_1346,N_1273,N_1250);
or U1347 (N_1347,N_1210,N_1280);
or U1348 (N_1348,N_1247,N_1260);
nand U1349 (N_1349,N_1215,N_1263);
and U1350 (N_1350,N_1246,N_1234);
and U1351 (N_1351,N_1220,N_1244);
xnor U1352 (N_1352,N_1282,N_1239);
nand U1353 (N_1353,N_1255,N_1295);
or U1354 (N_1354,N_1298,N_1228);
xor U1355 (N_1355,N_1253,N_1257);
and U1356 (N_1356,N_1293,N_1295);
nor U1357 (N_1357,N_1232,N_1281);
nor U1358 (N_1358,N_1204,N_1241);
xnor U1359 (N_1359,N_1203,N_1225);
nor U1360 (N_1360,N_1213,N_1256);
nand U1361 (N_1361,N_1231,N_1256);
xor U1362 (N_1362,N_1290,N_1271);
nor U1363 (N_1363,N_1229,N_1291);
or U1364 (N_1364,N_1269,N_1201);
nor U1365 (N_1365,N_1212,N_1272);
xnor U1366 (N_1366,N_1202,N_1284);
nand U1367 (N_1367,N_1228,N_1223);
and U1368 (N_1368,N_1237,N_1235);
nand U1369 (N_1369,N_1245,N_1227);
or U1370 (N_1370,N_1267,N_1231);
and U1371 (N_1371,N_1272,N_1283);
or U1372 (N_1372,N_1234,N_1296);
and U1373 (N_1373,N_1259,N_1249);
or U1374 (N_1374,N_1287,N_1229);
xnor U1375 (N_1375,N_1263,N_1287);
nand U1376 (N_1376,N_1218,N_1258);
xnor U1377 (N_1377,N_1228,N_1252);
nand U1378 (N_1378,N_1241,N_1254);
nor U1379 (N_1379,N_1224,N_1299);
and U1380 (N_1380,N_1295,N_1207);
xor U1381 (N_1381,N_1285,N_1205);
nor U1382 (N_1382,N_1235,N_1213);
nor U1383 (N_1383,N_1219,N_1277);
or U1384 (N_1384,N_1277,N_1256);
and U1385 (N_1385,N_1262,N_1288);
or U1386 (N_1386,N_1221,N_1262);
nand U1387 (N_1387,N_1206,N_1240);
nand U1388 (N_1388,N_1285,N_1216);
nor U1389 (N_1389,N_1247,N_1285);
and U1390 (N_1390,N_1282,N_1226);
xor U1391 (N_1391,N_1277,N_1289);
nand U1392 (N_1392,N_1258,N_1293);
and U1393 (N_1393,N_1291,N_1272);
nor U1394 (N_1394,N_1247,N_1229);
xor U1395 (N_1395,N_1265,N_1253);
nand U1396 (N_1396,N_1207,N_1247);
xnor U1397 (N_1397,N_1276,N_1281);
and U1398 (N_1398,N_1293,N_1215);
or U1399 (N_1399,N_1220,N_1236);
or U1400 (N_1400,N_1345,N_1384);
or U1401 (N_1401,N_1322,N_1376);
and U1402 (N_1402,N_1319,N_1382);
nand U1403 (N_1403,N_1386,N_1331);
nand U1404 (N_1404,N_1317,N_1335);
nand U1405 (N_1405,N_1350,N_1393);
or U1406 (N_1406,N_1338,N_1328);
and U1407 (N_1407,N_1306,N_1346);
xnor U1408 (N_1408,N_1398,N_1320);
xnor U1409 (N_1409,N_1360,N_1356);
nand U1410 (N_1410,N_1392,N_1369);
and U1411 (N_1411,N_1308,N_1372);
nor U1412 (N_1412,N_1363,N_1355);
xnor U1413 (N_1413,N_1397,N_1336);
nor U1414 (N_1414,N_1301,N_1342);
nand U1415 (N_1415,N_1334,N_1321);
or U1416 (N_1416,N_1347,N_1325);
xnor U1417 (N_1417,N_1316,N_1305);
or U1418 (N_1418,N_1362,N_1307);
or U1419 (N_1419,N_1381,N_1340);
and U1420 (N_1420,N_1388,N_1390);
and U1421 (N_1421,N_1380,N_1383);
nand U1422 (N_1422,N_1314,N_1361);
nor U1423 (N_1423,N_1330,N_1337);
xnor U1424 (N_1424,N_1312,N_1375);
nor U1425 (N_1425,N_1374,N_1348);
xor U1426 (N_1426,N_1379,N_1327);
xnor U1427 (N_1427,N_1315,N_1318);
nor U1428 (N_1428,N_1349,N_1352);
or U1429 (N_1429,N_1368,N_1357);
or U1430 (N_1430,N_1303,N_1365);
nor U1431 (N_1431,N_1324,N_1378);
and U1432 (N_1432,N_1329,N_1302);
or U1433 (N_1433,N_1309,N_1326);
nor U1434 (N_1434,N_1313,N_1332);
or U1435 (N_1435,N_1371,N_1364);
nand U1436 (N_1436,N_1343,N_1341);
and U1437 (N_1437,N_1366,N_1391);
nand U1438 (N_1438,N_1344,N_1339);
nor U1439 (N_1439,N_1353,N_1387);
nor U1440 (N_1440,N_1359,N_1395);
or U1441 (N_1441,N_1396,N_1399);
nor U1442 (N_1442,N_1377,N_1385);
nor U1443 (N_1443,N_1300,N_1310);
or U1444 (N_1444,N_1367,N_1351);
xnor U1445 (N_1445,N_1373,N_1311);
or U1446 (N_1446,N_1304,N_1394);
or U1447 (N_1447,N_1358,N_1333);
nand U1448 (N_1448,N_1323,N_1354);
nor U1449 (N_1449,N_1389,N_1370);
nand U1450 (N_1450,N_1331,N_1345);
xor U1451 (N_1451,N_1352,N_1346);
nand U1452 (N_1452,N_1364,N_1343);
or U1453 (N_1453,N_1333,N_1325);
or U1454 (N_1454,N_1325,N_1358);
xor U1455 (N_1455,N_1367,N_1390);
or U1456 (N_1456,N_1341,N_1375);
xor U1457 (N_1457,N_1377,N_1378);
and U1458 (N_1458,N_1324,N_1383);
xor U1459 (N_1459,N_1369,N_1333);
xor U1460 (N_1460,N_1398,N_1318);
or U1461 (N_1461,N_1385,N_1353);
nor U1462 (N_1462,N_1369,N_1326);
and U1463 (N_1463,N_1372,N_1320);
nand U1464 (N_1464,N_1322,N_1303);
or U1465 (N_1465,N_1321,N_1379);
xnor U1466 (N_1466,N_1382,N_1337);
nand U1467 (N_1467,N_1365,N_1359);
or U1468 (N_1468,N_1344,N_1303);
xnor U1469 (N_1469,N_1310,N_1312);
nor U1470 (N_1470,N_1321,N_1398);
and U1471 (N_1471,N_1333,N_1313);
nor U1472 (N_1472,N_1305,N_1348);
and U1473 (N_1473,N_1316,N_1344);
nor U1474 (N_1474,N_1356,N_1358);
and U1475 (N_1475,N_1354,N_1316);
nand U1476 (N_1476,N_1338,N_1316);
or U1477 (N_1477,N_1363,N_1332);
and U1478 (N_1478,N_1321,N_1368);
nor U1479 (N_1479,N_1367,N_1337);
nand U1480 (N_1480,N_1341,N_1321);
xor U1481 (N_1481,N_1361,N_1312);
or U1482 (N_1482,N_1370,N_1307);
and U1483 (N_1483,N_1305,N_1382);
xor U1484 (N_1484,N_1347,N_1380);
xnor U1485 (N_1485,N_1318,N_1320);
or U1486 (N_1486,N_1369,N_1390);
nand U1487 (N_1487,N_1355,N_1326);
nand U1488 (N_1488,N_1360,N_1399);
or U1489 (N_1489,N_1392,N_1359);
nand U1490 (N_1490,N_1300,N_1393);
nor U1491 (N_1491,N_1339,N_1307);
and U1492 (N_1492,N_1302,N_1363);
or U1493 (N_1493,N_1333,N_1373);
nand U1494 (N_1494,N_1393,N_1370);
or U1495 (N_1495,N_1346,N_1304);
and U1496 (N_1496,N_1312,N_1381);
xor U1497 (N_1497,N_1398,N_1373);
or U1498 (N_1498,N_1387,N_1380);
and U1499 (N_1499,N_1324,N_1374);
or U1500 (N_1500,N_1425,N_1427);
xnor U1501 (N_1501,N_1482,N_1429);
nand U1502 (N_1502,N_1453,N_1471);
and U1503 (N_1503,N_1488,N_1408);
xnor U1504 (N_1504,N_1443,N_1475);
nor U1505 (N_1505,N_1480,N_1478);
nor U1506 (N_1506,N_1459,N_1483);
nor U1507 (N_1507,N_1432,N_1458);
nand U1508 (N_1508,N_1477,N_1494);
or U1509 (N_1509,N_1487,N_1498);
or U1510 (N_1510,N_1416,N_1414);
xnor U1511 (N_1511,N_1493,N_1481);
or U1512 (N_1512,N_1465,N_1433);
nor U1513 (N_1513,N_1407,N_1495);
nand U1514 (N_1514,N_1457,N_1400);
nand U1515 (N_1515,N_1473,N_1499);
xnor U1516 (N_1516,N_1447,N_1474);
nor U1517 (N_1517,N_1437,N_1497);
or U1518 (N_1518,N_1455,N_1406);
nor U1519 (N_1519,N_1441,N_1404);
xor U1520 (N_1520,N_1417,N_1446);
or U1521 (N_1521,N_1435,N_1467);
xnor U1522 (N_1522,N_1491,N_1460);
and U1523 (N_1523,N_1464,N_1470);
nand U1524 (N_1524,N_1426,N_1422);
nor U1525 (N_1525,N_1492,N_1436);
nor U1526 (N_1526,N_1461,N_1410);
xnor U1527 (N_1527,N_1485,N_1442);
xor U1528 (N_1528,N_1456,N_1409);
and U1529 (N_1529,N_1403,N_1472);
nand U1530 (N_1530,N_1430,N_1434);
and U1531 (N_1531,N_1421,N_1439);
nand U1532 (N_1532,N_1423,N_1418);
and U1533 (N_1533,N_1451,N_1463);
and U1534 (N_1534,N_1466,N_1445);
or U1535 (N_1535,N_1450,N_1462);
nand U1536 (N_1536,N_1479,N_1431);
nand U1537 (N_1537,N_1438,N_1486);
nor U1538 (N_1538,N_1419,N_1415);
nor U1539 (N_1539,N_1413,N_1405);
nand U1540 (N_1540,N_1412,N_1411);
and U1541 (N_1541,N_1454,N_1420);
nand U1542 (N_1542,N_1401,N_1490);
nand U1543 (N_1543,N_1484,N_1440);
or U1544 (N_1544,N_1489,N_1452);
and U1545 (N_1545,N_1428,N_1402);
and U1546 (N_1546,N_1468,N_1469);
and U1547 (N_1547,N_1496,N_1476);
or U1548 (N_1548,N_1424,N_1449);
or U1549 (N_1549,N_1444,N_1448);
xor U1550 (N_1550,N_1436,N_1450);
xor U1551 (N_1551,N_1412,N_1475);
xor U1552 (N_1552,N_1481,N_1483);
nand U1553 (N_1553,N_1441,N_1469);
or U1554 (N_1554,N_1498,N_1444);
and U1555 (N_1555,N_1477,N_1400);
xor U1556 (N_1556,N_1432,N_1480);
nor U1557 (N_1557,N_1457,N_1416);
or U1558 (N_1558,N_1456,N_1492);
and U1559 (N_1559,N_1459,N_1492);
xor U1560 (N_1560,N_1418,N_1474);
nor U1561 (N_1561,N_1446,N_1481);
nand U1562 (N_1562,N_1424,N_1459);
or U1563 (N_1563,N_1420,N_1460);
nand U1564 (N_1564,N_1488,N_1493);
xnor U1565 (N_1565,N_1408,N_1496);
and U1566 (N_1566,N_1470,N_1496);
and U1567 (N_1567,N_1418,N_1471);
nand U1568 (N_1568,N_1450,N_1417);
nor U1569 (N_1569,N_1429,N_1484);
or U1570 (N_1570,N_1497,N_1423);
or U1571 (N_1571,N_1433,N_1425);
and U1572 (N_1572,N_1427,N_1494);
or U1573 (N_1573,N_1402,N_1431);
xor U1574 (N_1574,N_1410,N_1438);
xnor U1575 (N_1575,N_1476,N_1481);
or U1576 (N_1576,N_1414,N_1409);
nand U1577 (N_1577,N_1437,N_1463);
xor U1578 (N_1578,N_1424,N_1464);
and U1579 (N_1579,N_1467,N_1474);
nor U1580 (N_1580,N_1457,N_1483);
nor U1581 (N_1581,N_1414,N_1490);
or U1582 (N_1582,N_1461,N_1464);
and U1583 (N_1583,N_1461,N_1417);
nand U1584 (N_1584,N_1471,N_1422);
and U1585 (N_1585,N_1453,N_1482);
nand U1586 (N_1586,N_1488,N_1415);
nand U1587 (N_1587,N_1432,N_1481);
and U1588 (N_1588,N_1462,N_1429);
nor U1589 (N_1589,N_1494,N_1469);
nor U1590 (N_1590,N_1484,N_1424);
and U1591 (N_1591,N_1401,N_1483);
nor U1592 (N_1592,N_1412,N_1410);
or U1593 (N_1593,N_1410,N_1489);
nand U1594 (N_1594,N_1403,N_1498);
xnor U1595 (N_1595,N_1451,N_1406);
and U1596 (N_1596,N_1478,N_1444);
xor U1597 (N_1597,N_1415,N_1439);
xor U1598 (N_1598,N_1485,N_1465);
nand U1599 (N_1599,N_1495,N_1488);
nand U1600 (N_1600,N_1555,N_1503);
or U1601 (N_1601,N_1578,N_1582);
nor U1602 (N_1602,N_1569,N_1529);
nand U1603 (N_1603,N_1544,N_1526);
or U1604 (N_1604,N_1551,N_1570);
nand U1605 (N_1605,N_1574,N_1558);
nor U1606 (N_1606,N_1598,N_1514);
xor U1607 (N_1607,N_1519,N_1556);
and U1608 (N_1608,N_1587,N_1524);
nor U1609 (N_1609,N_1559,N_1515);
and U1610 (N_1610,N_1552,N_1531);
and U1611 (N_1611,N_1594,N_1501);
nor U1612 (N_1612,N_1573,N_1506);
nand U1613 (N_1613,N_1527,N_1576);
or U1614 (N_1614,N_1532,N_1589);
nand U1615 (N_1615,N_1540,N_1572);
nand U1616 (N_1616,N_1561,N_1549);
nor U1617 (N_1617,N_1508,N_1517);
or U1618 (N_1618,N_1591,N_1560);
nor U1619 (N_1619,N_1554,N_1518);
nand U1620 (N_1620,N_1543,N_1523);
nor U1621 (N_1621,N_1563,N_1586);
and U1622 (N_1622,N_1505,N_1580);
xnor U1623 (N_1623,N_1596,N_1546);
nor U1624 (N_1624,N_1541,N_1550);
nor U1625 (N_1625,N_1568,N_1512);
or U1626 (N_1626,N_1539,N_1584);
and U1627 (N_1627,N_1599,N_1588);
nor U1628 (N_1628,N_1581,N_1575);
and U1629 (N_1629,N_1597,N_1536);
nor U1630 (N_1630,N_1530,N_1537);
nor U1631 (N_1631,N_1564,N_1566);
or U1632 (N_1632,N_1547,N_1562);
nor U1633 (N_1633,N_1583,N_1592);
or U1634 (N_1634,N_1535,N_1590);
nor U1635 (N_1635,N_1513,N_1593);
or U1636 (N_1636,N_1548,N_1502);
nor U1637 (N_1637,N_1542,N_1500);
and U1638 (N_1638,N_1553,N_1534);
nand U1639 (N_1639,N_1528,N_1533);
and U1640 (N_1640,N_1507,N_1509);
or U1641 (N_1641,N_1510,N_1511);
xnor U1642 (N_1642,N_1522,N_1595);
nand U1643 (N_1643,N_1520,N_1565);
xnor U1644 (N_1644,N_1579,N_1525);
nand U1645 (N_1645,N_1577,N_1571);
xor U1646 (N_1646,N_1504,N_1557);
or U1647 (N_1647,N_1545,N_1567);
nand U1648 (N_1648,N_1516,N_1585);
nor U1649 (N_1649,N_1521,N_1538);
nand U1650 (N_1650,N_1568,N_1552);
nand U1651 (N_1651,N_1518,N_1574);
nand U1652 (N_1652,N_1595,N_1516);
or U1653 (N_1653,N_1579,N_1581);
or U1654 (N_1654,N_1521,N_1513);
or U1655 (N_1655,N_1561,N_1524);
or U1656 (N_1656,N_1561,N_1514);
nor U1657 (N_1657,N_1538,N_1510);
nand U1658 (N_1658,N_1527,N_1532);
nand U1659 (N_1659,N_1573,N_1576);
xnor U1660 (N_1660,N_1586,N_1591);
and U1661 (N_1661,N_1532,N_1502);
nand U1662 (N_1662,N_1556,N_1560);
nand U1663 (N_1663,N_1529,N_1568);
nor U1664 (N_1664,N_1516,N_1555);
or U1665 (N_1665,N_1549,N_1564);
nor U1666 (N_1666,N_1559,N_1502);
nor U1667 (N_1667,N_1577,N_1509);
nand U1668 (N_1668,N_1513,N_1525);
or U1669 (N_1669,N_1564,N_1575);
xor U1670 (N_1670,N_1567,N_1518);
or U1671 (N_1671,N_1510,N_1536);
and U1672 (N_1672,N_1519,N_1518);
or U1673 (N_1673,N_1591,N_1561);
nor U1674 (N_1674,N_1557,N_1598);
nor U1675 (N_1675,N_1507,N_1557);
xnor U1676 (N_1676,N_1509,N_1555);
xnor U1677 (N_1677,N_1596,N_1543);
or U1678 (N_1678,N_1501,N_1561);
nand U1679 (N_1679,N_1526,N_1571);
and U1680 (N_1680,N_1568,N_1562);
xnor U1681 (N_1681,N_1556,N_1565);
xor U1682 (N_1682,N_1596,N_1554);
nand U1683 (N_1683,N_1557,N_1558);
or U1684 (N_1684,N_1527,N_1504);
nor U1685 (N_1685,N_1559,N_1564);
nor U1686 (N_1686,N_1542,N_1546);
and U1687 (N_1687,N_1525,N_1539);
or U1688 (N_1688,N_1502,N_1500);
nor U1689 (N_1689,N_1548,N_1512);
and U1690 (N_1690,N_1519,N_1587);
or U1691 (N_1691,N_1594,N_1520);
and U1692 (N_1692,N_1559,N_1576);
and U1693 (N_1693,N_1537,N_1542);
nor U1694 (N_1694,N_1593,N_1578);
and U1695 (N_1695,N_1576,N_1519);
or U1696 (N_1696,N_1563,N_1511);
nand U1697 (N_1697,N_1587,N_1505);
nor U1698 (N_1698,N_1564,N_1590);
and U1699 (N_1699,N_1596,N_1598);
and U1700 (N_1700,N_1692,N_1619);
nand U1701 (N_1701,N_1682,N_1673);
and U1702 (N_1702,N_1659,N_1685);
and U1703 (N_1703,N_1615,N_1649);
nor U1704 (N_1704,N_1688,N_1606);
nor U1705 (N_1705,N_1668,N_1686);
nor U1706 (N_1706,N_1616,N_1667);
xnor U1707 (N_1707,N_1680,N_1605);
xor U1708 (N_1708,N_1691,N_1611);
xor U1709 (N_1709,N_1645,N_1623);
and U1710 (N_1710,N_1600,N_1638);
nor U1711 (N_1711,N_1610,N_1695);
nor U1712 (N_1712,N_1614,N_1641);
nor U1713 (N_1713,N_1648,N_1675);
xnor U1714 (N_1714,N_1678,N_1622);
or U1715 (N_1715,N_1602,N_1609);
nand U1716 (N_1716,N_1644,N_1687);
xnor U1717 (N_1717,N_1630,N_1608);
and U1718 (N_1718,N_1690,N_1650);
nor U1719 (N_1719,N_1612,N_1634);
nand U1720 (N_1720,N_1689,N_1642);
or U1721 (N_1721,N_1618,N_1635);
nor U1722 (N_1722,N_1626,N_1683);
or U1723 (N_1723,N_1627,N_1697);
xnor U1724 (N_1724,N_1632,N_1646);
and U1725 (N_1725,N_1693,N_1643);
or U1726 (N_1726,N_1681,N_1633);
nand U1727 (N_1727,N_1664,N_1674);
nor U1728 (N_1728,N_1660,N_1631);
xor U1729 (N_1729,N_1640,N_1671);
xnor U1730 (N_1730,N_1658,N_1677);
or U1731 (N_1731,N_1625,N_1670);
nand U1732 (N_1732,N_1603,N_1654);
nor U1733 (N_1733,N_1657,N_1653);
nand U1734 (N_1734,N_1651,N_1624);
nand U1735 (N_1735,N_1656,N_1694);
or U1736 (N_1736,N_1669,N_1621);
nor U1737 (N_1737,N_1684,N_1637);
nor U1738 (N_1738,N_1604,N_1663);
xor U1739 (N_1739,N_1652,N_1666);
xnor U1740 (N_1740,N_1607,N_1613);
nand U1741 (N_1741,N_1639,N_1676);
or U1742 (N_1742,N_1628,N_1617);
and U1743 (N_1743,N_1601,N_1620);
and U1744 (N_1744,N_1698,N_1662);
nand U1745 (N_1745,N_1636,N_1661);
or U1746 (N_1746,N_1699,N_1629);
and U1747 (N_1747,N_1679,N_1665);
xor U1748 (N_1748,N_1647,N_1696);
xnor U1749 (N_1749,N_1672,N_1655);
nand U1750 (N_1750,N_1666,N_1694);
xnor U1751 (N_1751,N_1681,N_1625);
and U1752 (N_1752,N_1627,N_1670);
nand U1753 (N_1753,N_1613,N_1657);
nand U1754 (N_1754,N_1615,N_1619);
nor U1755 (N_1755,N_1650,N_1675);
nand U1756 (N_1756,N_1685,N_1667);
nor U1757 (N_1757,N_1697,N_1665);
nor U1758 (N_1758,N_1641,N_1640);
or U1759 (N_1759,N_1674,N_1692);
or U1760 (N_1760,N_1692,N_1696);
nand U1761 (N_1761,N_1645,N_1669);
nand U1762 (N_1762,N_1657,N_1698);
or U1763 (N_1763,N_1699,N_1677);
nand U1764 (N_1764,N_1681,N_1667);
or U1765 (N_1765,N_1699,N_1664);
xnor U1766 (N_1766,N_1635,N_1616);
or U1767 (N_1767,N_1673,N_1629);
and U1768 (N_1768,N_1644,N_1603);
xor U1769 (N_1769,N_1673,N_1695);
or U1770 (N_1770,N_1618,N_1673);
or U1771 (N_1771,N_1607,N_1646);
nand U1772 (N_1772,N_1607,N_1655);
and U1773 (N_1773,N_1661,N_1678);
xor U1774 (N_1774,N_1642,N_1660);
xor U1775 (N_1775,N_1691,N_1600);
nor U1776 (N_1776,N_1662,N_1644);
nor U1777 (N_1777,N_1687,N_1658);
nor U1778 (N_1778,N_1629,N_1634);
nand U1779 (N_1779,N_1673,N_1654);
nor U1780 (N_1780,N_1646,N_1642);
nor U1781 (N_1781,N_1695,N_1630);
nand U1782 (N_1782,N_1631,N_1602);
xnor U1783 (N_1783,N_1637,N_1664);
nand U1784 (N_1784,N_1696,N_1632);
and U1785 (N_1785,N_1682,N_1689);
nor U1786 (N_1786,N_1639,N_1634);
xor U1787 (N_1787,N_1655,N_1622);
and U1788 (N_1788,N_1639,N_1651);
nand U1789 (N_1789,N_1642,N_1686);
xnor U1790 (N_1790,N_1605,N_1669);
xnor U1791 (N_1791,N_1687,N_1610);
xor U1792 (N_1792,N_1652,N_1628);
or U1793 (N_1793,N_1650,N_1660);
and U1794 (N_1794,N_1603,N_1651);
or U1795 (N_1795,N_1690,N_1635);
nor U1796 (N_1796,N_1699,N_1651);
xor U1797 (N_1797,N_1626,N_1678);
and U1798 (N_1798,N_1609,N_1642);
xor U1799 (N_1799,N_1648,N_1651);
and U1800 (N_1800,N_1761,N_1760);
nor U1801 (N_1801,N_1784,N_1793);
or U1802 (N_1802,N_1787,N_1799);
nor U1803 (N_1803,N_1750,N_1744);
nor U1804 (N_1804,N_1742,N_1775);
or U1805 (N_1805,N_1713,N_1729);
xor U1806 (N_1806,N_1733,N_1734);
nand U1807 (N_1807,N_1736,N_1743);
nand U1808 (N_1808,N_1720,N_1774);
or U1809 (N_1809,N_1746,N_1702);
nor U1810 (N_1810,N_1779,N_1780);
or U1811 (N_1811,N_1708,N_1786);
or U1812 (N_1812,N_1772,N_1740);
or U1813 (N_1813,N_1752,N_1739);
and U1814 (N_1814,N_1724,N_1759);
and U1815 (N_1815,N_1723,N_1704);
xor U1816 (N_1816,N_1747,N_1718);
and U1817 (N_1817,N_1791,N_1757);
and U1818 (N_1818,N_1738,N_1731);
nand U1819 (N_1819,N_1777,N_1756);
or U1820 (N_1820,N_1730,N_1706);
nor U1821 (N_1821,N_1776,N_1781);
and U1822 (N_1822,N_1783,N_1715);
or U1823 (N_1823,N_1790,N_1722);
xnor U1824 (N_1824,N_1785,N_1732);
nor U1825 (N_1825,N_1794,N_1795);
nor U1826 (N_1826,N_1741,N_1728);
nand U1827 (N_1827,N_1754,N_1727);
nor U1828 (N_1828,N_1768,N_1766);
and U1829 (N_1829,N_1711,N_1745);
or U1830 (N_1830,N_1705,N_1758);
nor U1831 (N_1831,N_1788,N_1796);
and U1832 (N_1832,N_1749,N_1778);
xor U1833 (N_1833,N_1700,N_1717);
or U1834 (N_1834,N_1735,N_1769);
xor U1835 (N_1835,N_1751,N_1782);
or U1836 (N_1836,N_1710,N_1792);
xnor U1837 (N_1837,N_1773,N_1726);
xor U1838 (N_1838,N_1765,N_1763);
and U1839 (N_1839,N_1721,N_1798);
nand U1840 (N_1840,N_1770,N_1712);
xnor U1841 (N_1841,N_1725,N_1762);
xor U1842 (N_1842,N_1709,N_1737);
xor U1843 (N_1843,N_1755,N_1748);
nand U1844 (N_1844,N_1716,N_1701);
and U1845 (N_1845,N_1703,N_1753);
nand U1846 (N_1846,N_1771,N_1767);
nor U1847 (N_1847,N_1789,N_1719);
nor U1848 (N_1848,N_1797,N_1764);
nand U1849 (N_1849,N_1707,N_1714);
xor U1850 (N_1850,N_1736,N_1781);
nand U1851 (N_1851,N_1776,N_1775);
and U1852 (N_1852,N_1741,N_1768);
xnor U1853 (N_1853,N_1795,N_1721);
or U1854 (N_1854,N_1753,N_1784);
xnor U1855 (N_1855,N_1743,N_1742);
or U1856 (N_1856,N_1704,N_1783);
xnor U1857 (N_1857,N_1714,N_1700);
nor U1858 (N_1858,N_1790,N_1773);
xnor U1859 (N_1859,N_1707,N_1713);
xnor U1860 (N_1860,N_1785,N_1724);
and U1861 (N_1861,N_1726,N_1740);
nand U1862 (N_1862,N_1711,N_1704);
or U1863 (N_1863,N_1784,N_1701);
and U1864 (N_1864,N_1715,N_1768);
nor U1865 (N_1865,N_1729,N_1797);
nor U1866 (N_1866,N_1705,N_1706);
nor U1867 (N_1867,N_1742,N_1758);
and U1868 (N_1868,N_1714,N_1728);
and U1869 (N_1869,N_1769,N_1706);
and U1870 (N_1870,N_1717,N_1751);
nor U1871 (N_1871,N_1743,N_1710);
nor U1872 (N_1872,N_1780,N_1783);
nand U1873 (N_1873,N_1700,N_1751);
nand U1874 (N_1874,N_1795,N_1701);
or U1875 (N_1875,N_1748,N_1764);
nand U1876 (N_1876,N_1728,N_1709);
or U1877 (N_1877,N_1771,N_1725);
nand U1878 (N_1878,N_1736,N_1790);
or U1879 (N_1879,N_1731,N_1732);
nor U1880 (N_1880,N_1780,N_1737);
nand U1881 (N_1881,N_1736,N_1716);
xnor U1882 (N_1882,N_1785,N_1746);
nand U1883 (N_1883,N_1772,N_1782);
nand U1884 (N_1884,N_1746,N_1721);
nor U1885 (N_1885,N_1779,N_1701);
nand U1886 (N_1886,N_1795,N_1735);
or U1887 (N_1887,N_1752,N_1771);
nand U1888 (N_1888,N_1742,N_1731);
nor U1889 (N_1889,N_1765,N_1718);
nor U1890 (N_1890,N_1745,N_1779);
and U1891 (N_1891,N_1778,N_1719);
or U1892 (N_1892,N_1748,N_1704);
and U1893 (N_1893,N_1765,N_1793);
and U1894 (N_1894,N_1733,N_1746);
nand U1895 (N_1895,N_1788,N_1789);
nand U1896 (N_1896,N_1721,N_1755);
or U1897 (N_1897,N_1766,N_1762);
or U1898 (N_1898,N_1788,N_1747);
and U1899 (N_1899,N_1718,N_1768);
nor U1900 (N_1900,N_1819,N_1866);
and U1901 (N_1901,N_1882,N_1800);
and U1902 (N_1902,N_1868,N_1893);
or U1903 (N_1903,N_1857,N_1870);
and U1904 (N_1904,N_1890,N_1879);
nand U1905 (N_1905,N_1892,N_1865);
and U1906 (N_1906,N_1899,N_1823);
xor U1907 (N_1907,N_1872,N_1896);
xor U1908 (N_1908,N_1832,N_1881);
or U1909 (N_1909,N_1889,N_1883);
nor U1910 (N_1910,N_1856,N_1806);
nand U1911 (N_1911,N_1840,N_1858);
and U1912 (N_1912,N_1818,N_1817);
nor U1913 (N_1913,N_1803,N_1847);
or U1914 (N_1914,N_1849,N_1864);
and U1915 (N_1915,N_1820,N_1898);
nor U1916 (N_1916,N_1885,N_1836);
and U1917 (N_1917,N_1846,N_1887);
and U1918 (N_1918,N_1854,N_1839);
nor U1919 (N_1919,N_1867,N_1877);
and U1920 (N_1920,N_1852,N_1880);
and U1921 (N_1921,N_1873,N_1848);
and U1922 (N_1922,N_1878,N_1804);
nor U1923 (N_1923,N_1874,N_1855);
or U1924 (N_1924,N_1884,N_1816);
and U1925 (N_1925,N_1888,N_1809);
nand U1926 (N_1926,N_1876,N_1826);
xnor U1927 (N_1927,N_1897,N_1871);
xor U1928 (N_1928,N_1802,N_1812);
xor U1929 (N_1929,N_1821,N_1845);
and U1930 (N_1930,N_1844,N_1810);
nor U1931 (N_1931,N_1842,N_1886);
and U1932 (N_1932,N_1814,N_1813);
nor U1933 (N_1933,N_1837,N_1862);
nand U1934 (N_1934,N_1807,N_1805);
or U1935 (N_1935,N_1808,N_1853);
and U1936 (N_1936,N_1875,N_1838);
or U1937 (N_1937,N_1834,N_1829);
nor U1938 (N_1938,N_1841,N_1824);
or U1939 (N_1939,N_1843,N_1828);
nand U1940 (N_1940,N_1815,N_1860);
xor U1941 (N_1941,N_1895,N_1801);
or U1942 (N_1942,N_1827,N_1850);
nor U1943 (N_1943,N_1835,N_1859);
nand U1944 (N_1944,N_1894,N_1822);
xor U1945 (N_1945,N_1833,N_1851);
nor U1946 (N_1946,N_1861,N_1831);
or U1947 (N_1947,N_1825,N_1811);
nor U1948 (N_1948,N_1869,N_1891);
xnor U1949 (N_1949,N_1863,N_1830);
xor U1950 (N_1950,N_1887,N_1814);
or U1951 (N_1951,N_1838,N_1895);
nand U1952 (N_1952,N_1857,N_1884);
nor U1953 (N_1953,N_1847,N_1882);
and U1954 (N_1954,N_1833,N_1871);
nand U1955 (N_1955,N_1867,N_1879);
xnor U1956 (N_1956,N_1814,N_1893);
xnor U1957 (N_1957,N_1833,N_1893);
or U1958 (N_1958,N_1871,N_1842);
and U1959 (N_1959,N_1826,N_1854);
nand U1960 (N_1960,N_1810,N_1864);
or U1961 (N_1961,N_1894,N_1800);
nand U1962 (N_1962,N_1878,N_1889);
nand U1963 (N_1963,N_1865,N_1809);
nand U1964 (N_1964,N_1834,N_1807);
xnor U1965 (N_1965,N_1896,N_1813);
and U1966 (N_1966,N_1822,N_1824);
nor U1967 (N_1967,N_1889,N_1899);
or U1968 (N_1968,N_1867,N_1807);
nor U1969 (N_1969,N_1801,N_1896);
nand U1970 (N_1970,N_1819,N_1898);
xnor U1971 (N_1971,N_1852,N_1894);
xor U1972 (N_1972,N_1893,N_1850);
and U1973 (N_1973,N_1819,N_1867);
xor U1974 (N_1974,N_1831,N_1892);
nor U1975 (N_1975,N_1825,N_1864);
nand U1976 (N_1976,N_1899,N_1832);
xor U1977 (N_1977,N_1861,N_1830);
nor U1978 (N_1978,N_1893,N_1863);
or U1979 (N_1979,N_1871,N_1827);
or U1980 (N_1980,N_1855,N_1857);
nor U1981 (N_1981,N_1863,N_1845);
or U1982 (N_1982,N_1877,N_1863);
xor U1983 (N_1983,N_1886,N_1811);
xnor U1984 (N_1984,N_1820,N_1828);
xnor U1985 (N_1985,N_1807,N_1847);
nor U1986 (N_1986,N_1845,N_1844);
xor U1987 (N_1987,N_1886,N_1832);
nor U1988 (N_1988,N_1888,N_1894);
nand U1989 (N_1989,N_1897,N_1852);
xnor U1990 (N_1990,N_1884,N_1889);
nand U1991 (N_1991,N_1838,N_1807);
nand U1992 (N_1992,N_1879,N_1838);
and U1993 (N_1993,N_1863,N_1812);
xnor U1994 (N_1994,N_1834,N_1865);
nand U1995 (N_1995,N_1804,N_1877);
nand U1996 (N_1996,N_1853,N_1892);
xor U1997 (N_1997,N_1898,N_1897);
xnor U1998 (N_1998,N_1803,N_1886);
and U1999 (N_1999,N_1801,N_1824);
nor U2000 (N_2000,N_1932,N_1960);
nor U2001 (N_2001,N_1946,N_1911);
or U2002 (N_2002,N_1925,N_1923);
or U2003 (N_2003,N_1921,N_1945);
or U2004 (N_2004,N_1943,N_1978);
nor U2005 (N_2005,N_1912,N_1954);
nand U2006 (N_2006,N_1917,N_1926);
nand U2007 (N_2007,N_1968,N_1929);
nand U2008 (N_2008,N_1983,N_1967);
and U2009 (N_2009,N_1985,N_1992);
or U2010 (N_2010,N_1999,N_1961);
nor U2011 (N_2011,N_1931,N_1918);
or U2012 (N_2012,N_1982,N_1998);
nand U2013 (N_2013,N_1906,N_1959);
or U2014 (N_2014,N_1971,N_1902);
or U2015 (N_2015,N_1904,N_1936);
nor U2016 (N_2016,N_1962,N_1924);
and U2017 (N_2017,N_1974,N_1984);
nand U2018 (N_2018,N_1908,N_1981);
nor U2019 (N_2019,N_1919,N_1995);
nor U2020 (N_2020,N_1939,N_1955);
or U2021 (N_2021,N_1986,N_1965);
and U2022 (N_2022,N_1969,N_1934);
xor U2023 (N_2023,N_1907,N_1935);
nor U2024 (N_2024,N_1979,N_1958);
and U2025 (N_2025,N_1966,N_1937);
or U2026 (N_2026,N_1942,N_1930);
nor U2027 (N_2027,N_1997,N_1922);
and U2028 (N_2028,N_1956,N_1996);
xor U2029 (N_2029,N_1977,N_1972);
nor U2030 (N_2030,N_1951,N_1993);
and U2031 (N_2031,N_1973,N_1914);
xnor U2032 (N_2032,N_1905,N_1901);
xnor U2033 (N_2033,N_1952,N_1980);
nand U2034 (N_2034,N_1994,N_1970);
nand U2035 (N_2035,N_1910,N_1944);
nor U2036 (N_2036,N_1990,N_1988);
xor U2037 (N_2037,N_1953,N_1989);
xnor U2038 (N_2038,N_1949,N_1975);
and U2039 (N_2039,N_1947,N_1938);
xor U2040 (N_2040,N_1909,N_1987);
nand U2041 (N_2041,N_1948,N_1940);
xor U2042 (N_2042,N_1915,N_1913);
xor U2043 (N_2043,N_1927,N_1950);
nand U2044 (N_2044,N_1957,N_1900);
and U2045 (N_2045,N_1964,N_1963);
and U2046 (N_2046,N_1903,N_1920);
nand U2047 (N_2047,N_1933,N_1928);
and U2048 (N_2048,N_1976,N_1941);
and U2049 (N_2049,N_1991,N_1916);
and U2050 (N_2050,N_1901,N_1964);
or U2051 (N_2051,N_1936,N_1982);
or U2052 (N_2052,N_1964,N_1990);
xor U2053 (N_2053,N_1990,N_1969);
or U2054 (N_2054,N_1921,N_1997);
xor U2055 (N_2055,N_1919,N_1965);
and U2056 (N_2056,N_1936,N_1990);
xnor U2057 (N_2057,N_1931,N_1969);
or U2058 (N_2058,N_1986,N_1936);
nor U2059 (N_2059,N_1910,N_1955);
xnor U2060 (N_2060,N_1927,N_1904);
or U2061 (N_2061,N_1957,N_1976);
and U2062 (N_2062,N_1994,N_1942);
nor U2063 (N_2063,N_1900,N_1908);
xnor U2064 (N_2064,N_1911,N_1990);
nor U2065 (N_2065,N_1957,N_1969);
xnor U2066 (N_2066,N_1925,N_1949);
and U2067 (N_2067,N_1969,N_1936);
or U2068 (N_2068,N_1966,N_1982);
or U2069 (N_2069,N_1965,N_1998);
xor U2070 (N_2070,N_1951,N_1959);
nor U2071 (N_2071,N_1984,N_1979);
nand U2072 (N_2072,N_1979,N_1946);
nand U2073 (N_2073,N_1999,N_1977);
nand U2074 (N_2074,N_1934,N_1991);
nor U2075 (N_2075,N_1920,N_1970);
nor U2076 (N_2076,N_1953,N_1950);
and U2077 (N_2077,N_1925,N_1915);
and U2078 (N_2078,N_1970,N_1957);
xnor U2079 (N_2079,N_1939,N_1930);
xnor U2080 (N_2080,N_1946,N_1927);
nand U2081 (N_2081,N_1956,N_1919);
nand U2082 (N_2082,N_1911,N_1978);
nor U2083 (N_2083,N_1985,N_1932);
nor U2084 (N_2084,N_1981,N_1916);
or U2085 (N_2085,N_1949,N_1950);
or U2086 (N_2086,N_1927,N_1948);
nor U2087 (N_2087,N_1991,N_1956);
nand U2088 (N_2088,N_1951,N_1963);
nor U2089 (N_2089,N_1962,N_1935);
nor U2090 (N_2090,N_1990,N_1914);
nor U2091 (N_2091,N_1923,N_1959);
and U2092 (N_2092,N_1923,N_1937);
xor U2093 (N_2093,N_1937,N_1924);
or U2094 (N_2094,N_1930,N_1925);
nor U2095 (N_2095,N_1926,N_1975);
and U2096 (N_2096,N_1952,N_1938);
xnor U2097 (N_2097,N_1910,N_1936);
xnor U2098 (N_2098,N_1970,N_1913);
nand U2099 (N_2099,N_1959,N_1919);
or U2100 (N_2100,N_2015,N_2031);
xnor U2101 (N_2101,N_2010,N_2004);
or U2102 (N_2102,N_2093,N_2036);
nor U2103 (N_2103,N_2017,N_2081);
and U2104 (N_2104,N_2073,N_2069);
nor U2105 (N_2105,N_2089,N_2088);
or U2106 (N_2106,N_2065,N_2028);
xnor U2107 (N_2107,N_2005,N_2096);
nand U2108 (N_2108,N_2006,N_2020);
nor U2109 (N_2109,N_2030,N_2016);
xor U2110 (N_2110,N_2067,N_2033);
or U2111 (N_2111,N_2064,N_2066);
nor U2112 (N_2112,N_2052,N_2034);
nor U2113 (N_2113,N_2029,N_2021);
or U2114 (N_2114,N_2003,N_2086);
xor U2115 (N_2115,N_2072,N_2079);
or U2116 (N_2116,N_2074,N_2057);
nor U2117 (N_2117,N_2077,N_2080);
and U2118 (N_2118,N_2037,N_2019);
nor U2119 (N_2119,N_2055,N_2047);
nand U2120 (N_2120,N_2018,N_2087);
xnor U2121 (N_2121,N_2060,N_2009);
nor U2122 (N_2122,N_2027,N_2061);
and U2123 (N_2123,N_2048,N_2042);
xnor U2124 (N_2124,N_2053,N_2041);
xor U2125 (N_2125,N_2013,N_2097);
nor U2126 (N_2126,N_2076,N_2049);
xnor U2127 (N_2127,N_2000,N_2046);
nor U2128 (N_2128,N_2091,N_2014);
xnor U2129 (N_2129,N_2051,N_2008);
or U2130 (N_2130,N_2044,N_2026);
nand U2131 (N_2131,N_2090,N_2071);
and U2132 (N_2132,N_2043,N_2035);
nand U2133 (N_2133,N_2082,N_2085);
nor U2134 (N_2134,N_2092,N_2032);
or U2135 (N_2135,N_2075,N_2063);
and U2136 (N_2136,N_2038,N_2040);
and U2137 (N_2137,N_2056,N_2012);
nand U2138 (N_2138,N_2002,N_2050);
nor U2139 (N_2139,N_2022,N_2059);
and U2140 (N_2140,N_2007,N_2039);
xnor U2141 (N_2141,N_2054,N_2099);
and U2142 (N_2142,N_2083,N_2095);
or U2143 (N_2143,N_2045,N_2023);
and U2144 (N_2144,N_2094,N_2024);
or U2145 (N_2145,N_2001,N_2078);
nor U2146 (N_2146,N_2062,N_2025);
xor U2147 (N_2147,N_2070,N_2011);
nor U2148 (N_2148,N_2068,N_2084);
nand U2149 (N_2149,N_2098,N_2058);
nand U2150 (N_2150,N_2049,N_2088);
xor U2151 (N_2151,N_2079,N_2046);
or U2152 (N_2152,N_2062,N_2056);
or U2153 (N_2153,N_2028,N_2063);
or U2154 (N_2154,N_2057,N_2000);
xor U2155 (N_2155,N_2013,N_2036);
and U2156 (N_2156,N_2000,N_2016);
xnor U2157 (N_2157,N_2082,N_2044);
and U2158 (N_2158,N_2041,N_2035);
xor U2159 (N_2159,N_2090,N_2011);
nand U2160 (N_2160,N_2083,N_2070);
or U2161 (N_2161,N_2075,N_2012);
nand U2162 (N_2162,N_2038,N_2045);
and U2163 (N_2163,N_2003,N_2038);
or U2164 (N_2164,N_2047,N_2031);
nor U2165 (N_2165,N_2003,N_2090);
nor U2166 (N_2166,N_2023,N_2017);
or U2167 (N_2167,N_2020,N_2045);
nand U2168 (N_2168,N_2082,N_2051);
xor U2169 (N_2169,N_2097,N_2051);
xor U2170 (N_2170,N_2027,N_2028);
nor U2171 (N_2171,N_2054,N_2040);
nand U2172 (N_2172,N_2015,N_2070);
xor U2173 (N_2173,N_2063,N_2055);
nor U2174 (N_2174,N_2095,N_2062);
or U2175 (N_2175,N_2093,N_2037);
or U2176 (N_2176,N_2034,N_2094);
or U2177 (N_2177,N_2033,N_2011);
or U2178 (N_2178,N_2008,N_2094);
nor U2179 (N_2179,N_2028,N_2089);
xnor U2180 (N_2180,N_2034,N_2086);
nand U2181 (N_2181,N_2081,N_2027);
or U2182 (N_2182,N_2060,N_2048);
nor U2183 (N_2183,N_2052,N_2002);
or U2184 (N_2184,N_2096,N_2019);
and U2185 (N_2185,N_2031,N_2070);
and U2186 (N_2186,N_2011,N_2084);
nor U2187 (N_2187,N_2002,N_2013);
nor U2188 (N_2188,N_2092,N_2076);
nand U2189 (N_2189,N_2060,N_2019);
nor U2190 (N_2190,N_2038,N_2005);
or U2191 (N_2191,N_2028,N_2075);
or U2192 (N_2192,N_2030,N_2008);
nand U2193 (N_2193,N_2089,N_2058);
or U2194 (N_2194,N_2028,N_2026);
nand U2195 (N_2195,N_2041,N_2076);
nand U2196 (N_2196,N_2005,N_2089);
nand U2197 (N_2197,N_2069,N_2052);
or U2198 (N_2198,N_2053,N_2088);
or U2199 (N_2199,N_2061,N_2028);
and U2200 (N_2200,N_2155,N_2129);
xnor U2201 (N_2201,N_2111,N_2189);
xnor U2202 (N_2202,N_2153,N_2120);
nand U2203 (N_2203,N_2147,N_2142);
nand U2204 (N_2204,N_2193,N_2190);
nor U2205 (N_2205,N_2128,N_2134);
xor U2206 (N_2206,N_2183,N_2146);
nand U2207 (N_2207,N_2162,N_2101);
or U2208 (N_2208,N_2112,N_2172);
or U2209 (N_2209,N_2158,N_2126);
nand U2210 (N_2210,N_2132,N_2125);
or U2211 (N_2211,N_2184,N_2176);
xor U2212 (N_2212,N_2140,N_2151);
nand U2213 (N_2213,N_2169,N_2173);
nand U2214 (N_2214,N_2137,N_2143);
xor U2215 (N_2215,N_2124,N_2187);
nand U2216 (N_2216,N_2102,N_2199);
nor U2217 (N_2217,N_2106,N_2110);
xor U2218 (N_2218,N_2105,N_2141);
and U2219 (N_2219,N_2174,N_2192);
and U2220 (N_2220,N_2163,N_2182);
and U2221 (N_2221,N_2166,N_2136);
nand U2222 (N_2222,N_2157,N_2103);
nor U2223 (N_2223,N_2160,N_2119);
or U2224 (N_2224,N_2139,N_2115);
nor U2225 (N_2225,N_2175,N_2109);
xor U2226 (N_2226,N_2123,N_2168);
nand U2227 (N_2227,N_2145,N_2104);
and U2228 (N_2228,N_2196,N_2144);
or U2229 (N_2229,N_2114,N_2181);
xor U2230 (N_2230,N_2159,N_2100);
nor U2231 (N_2231,N_2191,N_2156);
nor U2232 (N_2232,N_2127,N_2131);
and U2233 (N_2233,N_2108,N_2150);
xor U2234 (N_2234,N_2116,N_2118);
and U2235 (N_2235,N_2149,N_2164);
and U2236 (N_2236,N_2107,N_2133);
or U2237 (N_2237,N_2154,N_2178);
nor U2238 (N_2238,N_2152,N_2122);
or U2239 (N_2239,N_2197,N_2165);
xor U2240 (N_2240,N_2194,N_2121);
and U2241 (N_2241,N_2185,N_2195);
xor U2242 (N_2242,N_2167,N_2113);
and U2243 (N_2243,N_2177,N_2148);
or U2244 (N_2244,N_2188,N_2198);
and U2245 (N_2245,N_2161,N_2130);
xnor U2246 (N_2246,N_2179,N_2171);
nand U2247 (N_2247,N_2186,N_2138);
or U2248 (N_2248,N_2117,N_2135);
xnor U2249 (N_2249,N_2180,N_2170);
and U2250 (N_2250,N_2101,N_2159);
or U2251 (N_2251,N_2126,N_2184);
nand U2252 (N_2252,N_2136,N_2199);
nand U2253 (N_2253,N_2158,N_2159);
nor U2254 (N_2254,N_2189,N_2115);
xor U2255 (N_2255,N_2192,N_2131);
nor U2256 (N_2256,N_2164,N_2168);
or U2257 (N_2257,N_2171,N_2148);
nor U2258 (N_2258,N_2184,N_2130);
nand U2259 (N_2259,N_2143,N_2152);
nand U2260 (N_2260,N_2100,N_2193);
nor U2261 (N_2261,N_2169,N_2195);
nor U2262 (N_2262,N_2188,N_2104);
xnor U2263 (N_2263,N_2164,N_2136);
xnor U2264 (N_2264,N_2157,N_2161);
or U2265 (N_2265,N_2133,N_2125);
and U2266 (N_2266,N_2162,N_2127);
or U2267 (N_2267,N_2198,N_2166);
nand U2268 (N_2268,N_2119,N_2141);
nand U2269 (N_2269,N_2118,N_2180);
and U2270 (N_2270,N_2161,N_2182);
nor U2271 (N_2271,N_2101,N_2118);
nand U2272 (N_2272,N_2141,N_2161);
nor U2273 (N_2273,N_2182,N_2154);
xor U2274 (N_2274,N_2123,N_2133);
or U2275 (N_2275,N_2176,N_2100);
and U2276 (N_2276,N_2142,N_2163);
xor U2277 (N_2277,N_2107,N_2187);
and U2278 (N_2278,N_2124,N_2146);
nand U2279 (N_2279,N_2199,N_2161);
and U2280 (N_2280,N_2197,N_2181);
xnor U2281 (N_2281,N_2128,N_2183);
or U2282 (N_2282,N_2100,N_2132);
xnor U2283 (N_2283,N_2117,N_2100);
nand U2284 (N_2284,N_2133,N_2121);
and U2285 (N_2285,N_2129,N_2116);
and U2286 (N_2286,N_2153,N_2198);
xor U2287 (N_2287,N_2194,N_2141);
nor U2288 (N_2288,N_2135,N_2112);
nor U2289 (N_2289,N_2140,N_2117);
and U2290 (N_2290,N_2137,N_2125);
or U2291 (N_2291,N_2122,N_2174);
nand U2292 (N_2292,N_2173,N_2188);
nor U2293 (N_2293,N_2188,N_2110);
and U2294 (N_2294,N_2110,N_2193);
nor U2295 (N_2295,N_2140,N_2122);
nand U2296 (N_2296,N_2113,N_2177);
and U2297 (N_2297,N_2167,N_2189);
xor U2298 (N_2298,N_2188,N_2115);
nor U2299 (N_2299,N_2173,N_2116);
nand U2300 (N_2300,N_2283,N_2282);
or U2301 (N_2301,N_2203,N_2233);
nand U2302 (N_2302,N_2244,N_2241);
nor U2303 (N_2303,N_2278,N_2235);
nor U2304 (N_2304,N_2225,N_2201);
and U2305 (N_2305,N_2287,N_2274);
nor U2306 (N_2306,N_2248,N_2262);
and U2307 (N_2307,N_2220,N_2265);
xnor U2308 (N_2308,N_2258,N_2253);
xor U2309 (N_2309,N_2275,N_2240);
nand U2310 (N_2310,N_2288,N_2256);
or U2311 (N_2311,N_2226,N_2297);
or U2312 (N_2312,N_2228,N_2273);
nand U2313 (N_2313,N_2295,N_2218);
nor U2314 (N_2314,N_2231,N_2296);
and U2315 (N_2315,N_2211,N_2289);
and U2316 (N_2316,N_2268,N_2208);
and U2317 (N_2317,N_2279,N_2222);
or U2318 (N_2318,N_2264,N_2285);
or U2319 (N_2319,N_2213,N_2249);
nand U2320 (N_2320,N_2267,N_2209);
xor U2321 (N_2321,N_2259,N_2214);
nor U2322 (N_2322,N_2221,N_2204);
nor U2323 (N_2323,N_2293,N_2294);
nand U2324 (N_2324,N_2281,N_2202);
or U2325 (N_2325,N_2276,N_2257);
and U2326 (N_2326,N_2291,N_2238);
xor U2327 (N_2327,N_2252,N_2298);
and U2328 (N_2328,N_2272,N_2217);
xor U2329 (N_2329,N_2280,N_2234);
and U2330 (N_2330,N_2224,N_2207);
nor U2331 (N_2331,N_2200,N_2277);
and U2332 (N_2332,N_2216,N_2243);
nor U2333 (N_2333,N_2290,N_2246);
and U2334 (N_2334,N_2239,N_2270);
and U2335 (N_2335,N_2212,N_2227);
nor U2336 (N_2336,N_2271,N_2250);
or U2337 (N_2337,N_2299,N_2269);
nor U2338 (N_2338,N_2236,N_2219);
or U2339 (N_2339,N_2205,N_2292);
or U2340 (N_2340,N_2223,N_2254);
nor U2341 (N_2341,N_2260,N_2210);
nor U2342 (N_2342,N_2284,N_2286);
or U2343 (N_2343,N_2255,N_2215);
nand U2344 (N_2344,N_2261,N_2251);
and U2345 (N_2345,N_2230,N_2263);
nand U2346 (N_2346,N_2266,N_2245);
xor U2347 (N_2347,N_2237,N_2229);
nand U2348 (N_2348,N_2247,N_2206);
xor U2349 (N_2349,N_2232,N_2242);
nand U2350 (N_2350,N_2203,N_2285);
xor U2351 (N_2351,N_2203,N_2279);
xor U2352 (N_2352,N_2260,N_2239);
and U2353 (N_2353,N_2289,N_2233);
xnor U2354 (N_2354,N_2239,N_2261);
and U2355 (N_2355,N_2227,N_2264);
xor U2356 (N_2356,N_2286,N_2282);
or U2357 (N_2357,N_2240,N_2213);
nand U2358 (N_2358,N_2261,N_2218);
xnor U2359 (N_2359,N_2271,N_2215);
or U2360 (N_2360,N_2243,N_2206);
nand U2361 (N_2361,N_2219,N_2224);
or U2362 (N_2362,N_2233,N_2241);
xor U2363 (N_2363,N_2224,N_2261);
xnor U2364 (N_2364,N_2215,N_2213);
nand U2365 (N_2365,N_2249,N_2297);
and U2366 (N_2366,N_2202,N_2200);
nor U2367 (N_2367,N_2286,N_2209);
nand U2368 (N_2368,N_2271,N_2200);
and U2369 (N_2369,N_2272,N_2206);
and U2370 (N_2370,N_2245,N_2225);
xor U2371 (N_2371,N_2293,N_2201);
or U2372 (N_2372,N_2291,N_2273);
nand U2373 (N_2373,N_2218,N_2209);
xor U2374 (N_2374,N_2258,N_2234);
nand U2375 (N_2375,N_2265,N_2227);
nor U2376 (N_2376,N_2292,N_2283);
or U2377 (N_2377,N_2288,N_2247);
nand U2378 (N_2378,N_2235,N_2260);
nor U2379 (N_2379,N_2288,N_2245);
nand U2380 (N_2380,N_2266,N_2290);
or U2381 (N_2381,N_2288,N_2248);
nor U2382 (N_2382,N_2277,N_2227);
xor U2383 (N_2383,N_2262,N_2276);
and U2384 (N_2384,N_2218,N_2202);
nor U2385 (N_2385,N_2259,N_2296);
nand U2386 (N_2386,N_2205,N_2217);
xnor U2387 (N_2387,N_2218,N_2281);
and U2388 (N_2388,N_2291,N_2202);
xnor U2389 (N_2389,N_2259,N_2273);
and U2390 (N_2390,N_2228,N_2253);
or U2391 (N_2391,N_2255,N_2284);
nand U2392 (N_2392,N_2251,N_2232);
nor U2393 (N_2393,N_2242,N_2220);
xnor U2394 (N_2394,N_2269,N_2260);
xnor U2395 (N_2395,N_2292,N_2221);
and U2396 (N_2396,N_2227,N_2258);
or U2397 (N_2397,N_2283,N_2200);
or U2398 (N_2398,N_2203,N_2229);
xnor U2399 (N_2399,N_2260,N_2250);
or U2400 (N_2400,N_2381,N_2371);
xor U2401 (N_2401,N_2307,N_2342);
and U2402 (N_2402,N_2354,N_2324);
nand U2403 (N_2403,N_2365,N_2346);
and U2404 (N_2404,N_2305,N_2398);
or U2405 (N_2405,N_2348,N_2396);
nor U2406 (N_2406,N_2377,N_2302);
nand U2407 (N_2407,N_2313,N_2331);
and U2408 (N_2408,N_2343,N_2301);
nand U2409 (N_2409,N_2368,N_2364);
nand U2410 (N_2410,N_2380,N_2300);
xor U2411 (N_2411,N_2385,N_2327);
nand U2412 (N_2412,N_2391,N_2328);
or U2413 (N_2413,N_2347,N_2319);
nor U2414 (N_2414,N_2326,N_2321);
nor U2415 (N_2415,N_2318,N_2373);
xor U2416 (N_2416,N_2370,N_2399);
xnor U2417 (N_2417,N_2323,N_2303);
nand U2418 (N_2418,N_2395,N_2306);
nand U2419 (N_2419,N_2314,N_2378);
nor U2420 (N_2420,N_2352,N_2315);
nor U2421 (N_2421,N_2330,N_2358);
and U2422 (N_2422,N_2350,N_2369);
nor U2423 (N_2423,N_2322,N_2345);
xor U2424 (N_2424,N_2337,N_2388);
and U2425 (N_2425,N_2336,N_2316);
or U2426 (N_2426,N_2332,N_2390);
nand U2427 (N_2427,N_2374,N_2397);
nor U2428 (N_2428,N_2320,N_2310);
or U2429 (N_2429,N_2339,N_2384);
nand U2430 (N_2430,N_2308,N_2351);
nand U2431 (N_2431,N_2383,N_2392);
xnor U2432 (N_2432,N_2387,N_2357);
and U2433 (N_2433,N_2389,N_2372);
nor U2434 (N_2434,N_2360,N_2325);
nor U2435 (N_2435,N_2353,N_2317);
and U2436 (N_2436,N_2344,N_2361);
nor U2437 (N_2437,N_2386,N_2349);
xnor U2438 (N_2438,N_2356,N_2341);
nand U2439 (N_2439,N_2309,N_2375);
nand U2440 (N_2440,N_2355,N_2362);
or U2441 (N_2441,N_2334,N_2394);
or U2442 (N_2442,N_2359,N_2366);
and U2443 (N_2443,N_2329,N_2333);
or U2444 (N_2444,N_2382,N_2312);
nor U2445 (N_2445,N_2363,N_2367);
nand U2446 (N_2446,N_2311,N_2338);
nor U2447 (N_2447,N_2335,N_2393);
or U2448 (N_2448,N_2379,N_2376);
or U2449 (N_2449,N_2340,N_2304);
xnor U2450 (N_2450,N_2324,N_2319);
nor U2451 (N_2451,N_2310,N_2342);
and U2452 (N_2452,N_2399,N_2319);
nor U2453 (N_2453,N_2359,N_2344);
nand U2454 (N_2454,N_2340,N_2337);
and U2455 (N_2455,N_2327,N_2334);
xnor U2456 (N_2456,N_2327,N_2368);
nand U2457 (N_2457,N_2381,N_2395);
xor U2458 (N_2458,N_2363,N_2374);
and U2459 (N_2459,N_2335,N_2336);
xnor U2460 (N_2460,N_2304,N_2358);
xnor U2461 (N_2461,N_2390,N_2313);
and U2462 (N_2462,N_2360,N_2330);
or U2463 (N_2463,N_2339,N_2379);
or U2464 (N_2464,N_2362,N_2310);
and U2465 (N_2465,N_2393,N_2344);
nor U2466 (N_2466,N_2369,N_2372);
or U2467 (N_2467,N_2329,N_2345);
or U2468 (N_2468,N_2334,N_2335);
or U2469 (N_2469,N_2378,N_2374);
xor U2470 (N_2470,N_2354,N_2392);
nor U2471 (N_2471,N_2359,N_2364);
xnor U2472 (N_2472,N_2325,N_2321);
xor U2473 (N_2473,N_2341,N_2363);
nor U2474 (N_2474,N_2339,N_2328);
or U2475 (N_2475,N_2361,N_2337);
or U2476 (N_2476,N_2374,N_2340);
nor U2477 (N_2477,N_2374,N_2344);
and U2478 (N_2478,N_2329,N_2344);
nand U2479 (N_2479,N_2324,N_2345);
and U2480 (N_2480,N_2339,N_2362);
xor U2481 (N_2481,N_2373,N_2330);
xor U2482 (N_2482,N_2355,N_2348);
and U2483 (N_2483,N_2367,N_2312);
xor U2484 (N_2484,N_2383,N_2322);
and U2485 (N_2485,N_2342,N_2377);
and U2486 (N_2486,N_2327,N_2301);
nor U2487 (N_2487,N_2336,N_2308);
and U2488 (N_2488,N_2379,N_2349);
or U2489 (N_2489,N_2347,N_2308);
xnor U2490 (N_2490,N_2347,N_2330);
or U2491 (N_2491,N_2338,N_2308);
nand U2492 (N_2492,N_2351,N_2327);
or U2493 (N_2493,N_2337,N_2339);
nor U2494 (N_2494,N_2396,N_2363);
nand U2495 (N_2495,N_2332,N_2365);
nand U2496 (N_2496,N_2359,N_2361);
xor U2497 (N_2497,N_2325,N_2331);
nor U2498 (N_2498,N_2310,N_2391);
nand U2499 (N_2499,N_2307,N_2309);
xor U2500 (N_2500,N_2442,N_2489);
and U2501 (N_2501,N_2428,N_2470);
nand U2502 (N_2502,N_2443,N_2482);
nand U2503 (N_2503,N_2475,N_2488);
nor U2504 (N_2504,N_2483,N_2431);
xor U2505 (N_2505,N_2459,N_2403);
xor U2506 (N_2506,N_2407,N_2444);
xor U2507 (N_2507,N_2427,N_2435);
xnor U2508 (N_2508,N_2400,N_2404);
or U2509 (N_2509,N_2445,N_2424);
or U2510 (N_2510,N_2474,N_2490);
xnor U2511 (N_2511,N_2454,N_2423);
xor U2512 (N_2512,N_2413,N_2466);
nand U2513 (N_2513,N_2471,N_2452);
or U2514 (N_2514,N_2426,N_2447);
nand U2515 (N_2515,N_2440,N_2477);
xnor U2516 (N_2516,N_2467,N_2455);
nand U2517 (N_2517,N_2494,N_2496);
nand U2518 (N_2518,N_2479,N_2432);
or U2519 (N_2519,N_2433,N_2420);
nor U2520 (N_2520,N_2464,N_2414);
nand U2521 (N_2521,N_2430,N_2458);
or U2522 (N_2522,N_2448,N_2478);
nand U2523 (N_2523,N_2485,N_2491);
and U2524 (N_2524,N_2484,N_2480);
nor U2525 (N_2525,N_2493,N_2499);
nand U2526 (N_2526,N_2422,N_2418);
or U2527 (N_2527,N_2439,N_2481);
nor U2528 (N_2528,N_2497,N_2456);
nand U2529 (N_2529,N_2468,N_2451);
nor U2530 (N_2530,N_2472,N_2408);
nand U2531 (N_2531,N_2463,N_2417);
xor U2532 (N_2532,N_2473,N_2410);
nand U2533 (N_2533,N_2425,N_2453);
or U2534 (N_2534,N_2446,N_2436);
and U2535 (N_2535,N_2415,N_2434);
nand U2536 (N_2536,N_2449,N_2421);
nand U2537 (N_2537,N_2411,N_2429);
nor U2538 (N_2538,N_2498,N_2461);
nand U2539 (N_2539,N_2437,N_2457);
and U2540 (N_2540,N_2416,N_2450);
xnor U2541 (N_2541,N_2460,N_2419);
nor U2542 (N_2542,N_2487,N_2409);
nand U2543 (N_2543,N_2495,N_2441);
and U2544 (N_2544,N_2401,N_2462);
or U2545 (N_2545,N_2438,N_2412);
xor U2546 (N_2546,N_2465,N_2406);
and U2547 (N_2547,N_2486,N_2405);
and U2548 (N_2548,N_2492,N_2469);
or U2549 (N_2549,N_2402,N_2476);
and U2550 (N_2550,N_2443,N_2450);
and U2551 (N_2551,N_2415,N_2421);
nand U2552 (N_2552,N_2485,N_2490);
nand U2553 (N_2553,N_2465,N_2429);
and U2554 (N_2554,N_2446,N_2474);
xor U2555 (N_2555,N_2401,N_2438);
and U2556 (N_2556,N_2426,N_2404);
nor U2557 (N_2557,N_2459,N_2478);
xnor U2558 (N_2558,N_2430,N_2439);
nor U2559 (N_2559,N_2462,N_2470);
and U2560 (N_2560,N_2464,N_2482);
and U2561 (N_2561,N_2494,N_2452);
nor U2562 (N_2562,N_2427,N_2411);
or U2563 (N_2563,N_2468,N_2428);
xnor U2564 (N_2564,N_2420,N_2452);
nand U2565 (N_2565,N_2442,N_2483);
or U2566 (N_2566,N_2476,N_2487);
xor U2567 (N_2567,N_2402,N_2440);
or U2568 (N_2568,N_2454,N_2453);
and U2569 (N_2569,N_2448,N_2488);
nand U2570 (N_2570,N_2466,N_2457);
or U2571 (N_2571,N_2479,N_2402);
nand U2572 (N_2572,N_2482,N_2422);
nand U2573 (N_2573,N_2407,N_2411);
or U2574 (N_2574,N_2403,N_2443);
nand U2575 (N_2575,N_2402,N_2451);
nor U2576 (N_2576,N_2493,N_2436);
nor U2577 (N_2577,N_2400,N_2457);
and U2578 (N_2578,N_2425,N_2496);
nor U2579 (N_2579,N_2494,N_2450);
xor U2580 (N_2580,N_2425,N_2440);
or U2581 (N_2581,N_2460,N_2477);
xor U2582 (N_2582,N_2497,N_2424);
and U2583 (N_2583,N_2414,N_2485);
nand U2584 (N_2584,N_2454,N_2417);
xor U2585 (N_2585,N_2412,N_2423);
and U2586 (N_2586,N_2416,N_2484);
nand U2587 (N_2587,N_2426,N_2465);
xor U2588 (N_2588,N_2483,N_2457);
xnor U2589 (N_2589,N_2488,N_2426);
and U2590 (N_2590,N_2408,N_2489);
xnor U2591 (N_2591,N_2463,N_2474);
nand U2592 (N_2592,N_2426,N_2466);
or U2593 (N_2593,N_2441,N_2413);
and U2594 (N_2594,N_2488,N_2446);
nor U2595 (N_2595,N_2498,N_2426);
nor U2596 (N_2596,N_2412,N_2415);
xnor U2597 (N_2597,N_2420,N_2402);
nor U2598 (N_2598,N_2468,N_2489);
xor U2599 (N_2599,N_2462,N_2435);
nor U2600 (N_2600,N_2572,N_2545);
or U2601 (N_2601,N_2599,N_2540);
nor U2602 (N_2602,N_2524,N_2546);
nor U2603 (N_2603,N_2535,N_2584);
nand U2604 (N_2604,N_2552,N_2590);
or U2605 (N_2605,N_2542,N_2528);
nand U2606 (N_2606,N_2588,N_2580);
and U2607 (N_2607,N_2567,N_2531);
nand U2608 (N_2608,N_2585,N_2562);
nor U2609 (N_2609,N_2500,N_2569);
xor U2610 (N_2610,N_2514,N_2548);
nor U2611 (N_2611,N_2586,N_2593);
or U2612 (N_2612,N_2520,N_2533);
xnor U2613 (N_2613,N_2517,N_2511);
nand U2614 (N_2614,N_2592,N_2519);
or U2615 (N_2615,N_2543,N_2561);
xnor U2616 (N_2616,N_2509,N_2594);
or U2617 (N_2617,N_2502,N_2530);
and U2618 (N_2618,N_2566,N_2510);
and U2619 (N_2619,N_2557,N_2526);
nand U2620 (N_2620,N_2529,N_2508);
nor U2621 (N_2621,N_2554,N_2558);
or U2622 (N_2622,N_2522,N_2571);
or U2623 (N_2623,N_2583,N_2582);
and U2624 (N_2624,N_2523,N_2503);
and U2625 (N_2625,N_2506,N_2544);
nor U2626 (N_2626,N_2518,N_2597);
nand U2627 (N_2627,N_2504,N_2501);
or U2628 (N_2628,N_2553,N_2549);
nor U2629 (N_2629,N_2568,N_2591);
nor U2630 (N_2630,N_2574,N_2559);
nand U2631 (N_2631,N_2551,N_2538);
nand U2632 (N_2632,N_2581,N_2576);
xor U2633 (N_2633,N_2598,N_2515);
nor U2634 (N_2634,N_2527,N_2577);
and U2635 (N_2635,N_2565,N_2536);
nor U2636 (N_2636,N_2596,N_2563);
and U2637 (N_2637,N_2570,N_2556);
xor U2638 (N_2638,N_2516,N_2507);
nand U2639 (N_2639,N_2573,N_2532);
and U2640 (N_2640,N_2595,N_2525);
or U2641 (N_2641,N_2564,N_2547);
nand U2642 (N_2642,N_2560,N_2589);
nor U2643 (N_2643,N_2541,N_2579);
xor U2644 (N_2644,N_2587,N_2550);
or U2645 (N_2645,N_2521,N_2578);
xnor U2646 (N_2646,N_2537,N_2534);
nand U2647 (N_2647,N_2539,N_2555);
or U2648 (N_2648,N_2513,N_2512);
and U2649 (N_2649,N_2575,N_2505);
xor U2650 (N_2650,N_2504,N_2568);
and U2651 (N_2651,N_2595,N_2535);
nor U2652 (N_2652,N_2533,N_2547);
or U2653 (N_2653,N_2507,N_2548);
or U2654 (N_2654,N_2520,N_2521);
or U2655 (N_2655,N_2559,N_2506);
and U2656 (N_2656,N_2500,N_2573);
xor U2657 (N_2657,N_2519,N_2564);
and U2658 (N_2658,N_2570,N_2527);
nand U2659 (N_2659,N_2516,N_2534);
or U2660 (N_2660,N_2571,N_2558);
or U2661 (N_2661,N_2550,N_2537);
nand U2662 (N_2662,N_2581,N_2588);
and U2663 (N_2663,N_2542,N_2500);
xnor U2664 (N_2664,N_2595,N_2560);
or U2665 (N_2665,N_2589,N_2551);
xor U2666 (N_2666,N_2542,N_2501);
and U2667 (N_2667,N_2563,N_2552);
or U2668 (N_2668,N_2590,N_2527);
and U2669 (N_2669,N_2537,N_2581);
xor U2670 (N_2670,N_2526,N_2554);
xor U2671 (N_2671,N_2558,N_2504);
or U2672 (N_2672,N_2539,N_2552);
or U2673 (N_2673,N_2552,N_2582);
nand U2674 (N_2674,N_2563,N_2587);
nand U2675 (N_2675,N_2552,N_2504);
or U2676 (N_2676,N_2569,N_2544);
or U2677 (N_2677,N_2500,N_2503);
nor U2678 (N_2678,N_2502,N_2573);
nand U2679 (N_2679,N_2548,N_2587);
nor U2680 (N_2680,N_2588,N_2553);
nand U2681 (N_2681,N_2503,N_2590);
nand U2682 (N_2682,N_2502,N_2503);
xor U2683 (N_2683,N_2582,N_2563);
nand U2684 (N_2684,N_2556,N_2593);
nand U2685 (N_2685,N_2590,N_2523);
and U2686 (N_2686,N_2541,N_2560);
xnor U2687 (N_2687,N_2523,N_2579);
nor U2688 (N_2688,N_2537,N_2527);
and U2689 (N_2689,N_2537,N_2576);
xor U2690 (N_2690,N_2516,N_2505);
or U2691 (N_2691,N_2526,N_2550);
xnor U2692 (N_2692,N_2576,N_2550);
or U2693 (N_2693,N_2578,N_2531);
nand U2694 (N_2694,N_2549,N_2510);
nor U2695 (N_2695,N_2575,N_2582);
xor U2696 (N_2696,N_2587,N_2542);
xnor U2697 (N_2697,N_2530,N_2540);
and U2698 (N_2698,N_2530,N_2525);
and U2699 (N_2699,N_2529,N_2539);
and U2700 (N_2700,N_2636,N_2655);
xnor U2701 (N_2701,N_2649,N_2615);
xnor U2702 (N_2702,N_2686,N_2628);
and U2703 (N_2703,N_2602,N_2644);
or U2704 (N_2704,N_2684,N_2633);
nand U2705 (N_2705,N_2677,N_2604);
or U2706 (N_2706,N_2605,N_2648);
nand U2707 (N_2707,N_2687,N_2632);
and U2708 (N_2708,N_2606,N_2607);
and U2709 (N_2709,N_2613,N_2690);
xnor U2710 (N_2710,N_2631,N_2647);
or U2711 (N_2711,N_2614,N_2622);
or U2712 (N_2712,N_2641,N_2671);
xor U2713 (N_2713,N_2663,N_2689);
and U2714 (N_2714,N_2661,N_2662);
nand U2715 (N_2715,N_2629,N_2674);
xor U2716 (N_2716,N_2653,N_2603);
nor U2717 (N_2717,N_2695,N_2640);
nor U2718 (N_2718,N_2650,N_2639);
nor U2719 (N_2719,N_2652,N_2688);
nor U2720 (N_2720,N_2645,N_2668);
or U2721 (N_2721,N_2691,N_2685);
and U2722 (N_2722,N_2610,N_2620);
nand U2723 (N_2723,N_2680,N_2609);
nand U2724 (N_2724,N_2676,N_2697);
xnor U2725 (N_2725,N_2630,N_2600);
or U2726 (N_2726,N_2651,N_2623);
or U2727 (N_2727,N_2658,N_2643);
and U2728 (N_2728,N_2694,N_2679);
nor U2729 (N_2729,N_2678,N_2621);
xnor U2730 (N_2730,N_2637,N_2635);
and U2731 (N_2731,N_2692,N_2681);
and U2732 (N_2732,N_2612,N_2611);
nor U2733 (N_2733,N_2667,N_2617);
and U2734 (N_2734,N_2619,N_2642);
nand U2735 (N_2735,N_2601,N_2665);
nand U2736 (N_2736,N_2682,N_2616);
xnor U2737 (N_2737,N_2654,N_2627);
and U2738 (N_2738,N_2660,N_2624);
nand U2739 (N_2739,N_2673,N_2659);
and U2740 (N_2740,N_2657,N_2656);
nor U2741 (N_2741,N_2634,N_2693);
or U2742 (N_2742,N_2683,N_2698);
or U2743 (N_2743,N_2608,N_2646);
or U2744 (N_2744,N_2626,N_2625);
or U2745 (N_2745,N_2638,N_2670);
and U2746 (N_2746,N_2666,N_2699);
and U2747 (N_2747,N_2696,N_2675);
or U2748 (N_2748,N_2669,N_2664);
and U2749 (N_2749,N_2672,N_2618);
nor U2750 (N_2750,N_2681,N_2633);
nor U2751 (N_2751,N_2609,N_2611);
nor U2752 (N_2752,N_2640,N_2603);
nand U2753 (N_2753,N_2640,N_2683);
and U2754 (N_2754,N_2698,N_2699);
or U2755 (N_2755,N_2681,N_2631);
xnor U2756 (N_2756,N_2661,N_2627);
and U2757 (N_2757,N_2606,N_2641);
xnor U2758 (N_2758,N_2680,N_2699);
nand U2759 (N_2759,N_2649,N_2679);
nor U2760 (N_2760,N_2639,N_2609);
and U2761 (N_2761,N_2604,N_2647);
nor U2762 (N_2762,N_2648,N_2679);
and U2763 (N_2763,N_2697,N_2633);
and U2764 (N_2764,N_2689,N_2618);
and U2765 (N_2765,N_2628,N_2682);
or U2766 (N_2766,N_2648,N_2634);
xnor U2767 (N_2767,N_2631,N_2621);
or U2768 (N_2768,N_2621,N_2604);
and U2769 (N_2769,N_2699,N_2656);
xor U2770 (N_2770,N_2603,N_2632);
nand U2771 (N_2771,N_2695,N_2676);
xnor U2772 (N_2772,N_2644,N_2666);
xnor U2773 (N_2773,N_2684,N_2646);
xnor U2774 (N_2774,N_2688,N_2651);
nor U2775 (N_2775,N_2681,N_2605);
xnor U2776 (N_2776,N_2671,N_2644);
or U2777 (N_2777,N_2615,N_2628);
nand U2778 (N_2778,N_2603,N_2671);
xor U2779 (N_2779,N_2676,N_2659);
xnor U2780 (N_2780,N_2647,N_2624);
nand U2781 (N_2781,N_2670,N_2697);
and U2782 (N_2782,N_2621,N_2608);
and U2783 (N_2783,N_2607,N_2679);
nand U2784 (N_2784,N_2640,N_2631);
nor U2785 (N_2785,N_2648,N_2660);
or U2786 (N_2786,N_2663,N_2693);
nand U2787 (N_2787,N_2688,N_2612);
or U2788 (N_2788,N_2644,N_2616);
nand U2789 (N_2789,N_2655,N_2653);
nand U2790 (N_2790,N_2665,N_2676);
nand U2791 (N_2791,N_2643,N_2676);
and U2792 (N_2792,N_2696,N_2657);
nand U2793 (N_2793,N_2611,N_2667);
and U2794 (N_2794,N_2638,N_2667);
xnor U2795 (N_2795,N_2659,N_2657);
and U2796 (N_2796,N_2630,N_2666);
and U2797 (N_2797,N_2657,N_2649);
and U2798 (N_2798,N_2651,N_2660);
nor U2799 (N_2799,N_2645,N_2604);
xor U2800 (N_2800,N_2796,N_2791);
nand U2801 (N_2801,N_2751,N_2734);
nand U2802 (N_2802,N_2773,N_2739);
and U2803 (N_2803,N_2785,N_2788);
or U2804 (N_2804,N_2787,N_2766);
xnor U2805 (N_2805,N_2742,N_2752);
xor U2806 (N_2806,N_2714,N_2760);
and U2807 (N_2807,N_2781,N_2706);
nand U2808 (N_2808,N_2786,N_2733);
xor U2809 (N_2809,N_2792,N_2703);
nand U2810 (N_2810,N_2719,N_2789);
xor U2811 (N_2811,N_2731,N_2748);
and U2812 (N_2812,N_2780,N_2782);
or U2813 (N_2813,N_2778,N_2741);
and U2814 (N_2814,N_2736,N_2710);
xnor U2815 (N_2815,N_2737,N_2756);
and U2816 (N_2816,N_2723,N_2716);
and U2817 (N_2817,N_2728,N_2761);
or U2818 (N_2818,N_2771,N_2758);
xor U2819 (N_2819,N_2777,N_2718);
xor U2820 (N_2820,N_2774,N_2764);
nor U2821 (N_2821,N_2783,N_2762);
xnor U2822 (N_2822,N_2717,N_2772);
or U2823 (N_2823,N_2702,N_2747);
nand U2824 (N_2824,N_2738,N_2799);
and U2825 (N_2825,N_2744,N_2779);
nand U2826 (N_2826,N_2767,N_2784);
nor U2827 (N_2827,N_2732,N_2735);
nor U2828 (N_2828,N_2770,N_2749);
nand U2829 (N_2829,N_2720,N_2726);
nand U2830 (N_2830,N_2750,N_2798);
and U2831 (N_2831,N_2740,N_2765);
nor U2832 (N_2832,N_2709,N_2707);
and U2833 (N_2833,N_2793,N_2775);
nand U2834 (N_2834,N_2753,N_2759);
or U2835 (N_2835,N_2729,N_2743);
nand U2836 (N_2836,N_2755,N_2790);
and U2837 (N_2837,N_2711,N_2730);
and U2838 (N_2838,N_2700,N_2722);
nor U2839 (N_2839,N_2705,N_2754);
xor U2840 (N_2840,N_2708,N_2701);
xnor U2841 (N_2841,N_2724,N_2794);
or U2842 (N_2842,N_2712,N_2797);
nand U2843 (N_2843,N_2769,N_2757);
xor U2844 (N_2844,N_2725,N_2795);
nand U2845 (N_2845,N_2776,N_2745);
nor U2846 (N_2846,N_2721,N_2713);
nor U2847 (N_2847,N_2727,N_2704);
or U2848 (N_2848,N_2746,N_2763);
nand U2849 (N_2849,N_2768,N_2715);
xnor U2850 (N_2850,N_2750,N_2723);
xnor U2851 (N_2851,N_2741,N_2703);
or U2852 (N_2852,N_2701,N_2736);
nand U2853 (N_2853,N_2718,N_2757);
xnor U2854 (N_2854,N_2722,N_2712);
xor U2855 (N_2855,N_2714,N_2708);
nor U2856 (N_2856,N_2761,N_2772);
nor U2857 (N_2857,N_2744,N_2723);
nor U2858 (N_2858,N_2743,N_2756);
and U2859 (N_2859,N_2763,N_2743);
or U2860 (N_2860,N_2788,N_2744);
xor U2861 (N_2861,N_2773,N_2796);
and U2862 (N_2862,N_2740,N_2786);
xor U2863 (N_2863,N_2718,N_2753);
and U2864 (N_2864,N_2748,N_2705);
nand U2865 (N_2865,N_2768,N_2778);
nor U2866 (N_2866,N_2770,N_2738);
and U2867 (N_2867,N_2749,N_2715);
and U2868 (N_2868,N_2700,N_2772);
nor U2869 (N_2869,N_2716,N_2707);
or U2870 (N_2870,N_2751,N_2705);
nor U2871 (N_2871,N_2745,N_2732);
xnor U2872 (N_2872,N_2757,N_2715);
xor U2873 (N_2873,N_2756,N_2774);
or U2874 (N_2874,N_2736,N_2787);
and U2875 (N_2875,N_2708,N_2775);
xor U2876 (N_2876,N_2728,N_2731);
and U2877 (N_2877,N_2759,N_2710);
xor U2878 (N_2878,N_2753,N_2762);
xnor U2879 (N_2879,N_2792,N_2709);
xor U2880 (N_2880,N_2798,N_2738);
nand U2881 (N_2881,N_2754,N_2701);
nor U2882 (N_2882,N_2748,N_2728);
nand U2883 (N_2883,N_2710,N_2772);
and U2884 (N_2884,N_2738,N_2720);
xnor U2885 (N_2885,N_2759,N_2737);
xnor U2886 (N_2886,N_2721,N_2761);
xnor U2887 (N_2887,N_2723,N_2793);
and U2888 (N_2888,N_2782,N_2774);
and U2889 (N_2889,N_2709,N_2701);
and U2890 (N_2890,N_2792,N_2742);
nor U2891 (N_2891,N_2732,N_2777);
and U2892 (N_2892,N_2758,N_2798);
xnor U2893 (N_2893,N_2743,N_2726);
or U2894 (N_2894,N_2777,N_2719);
or U2895 (N_2895,N_2713,N_2754);
nor U2896 (N_2896,N_2760,N_2742);
or U2897 (N_2897,N_2768,N_2746);
nor U2898 (N_2898,N_2702,N_2721);
xnor U2899 (N_2899,N_2724,N_2763);
xnor U2900 (N_2900,N_2850,N_2818);
nand U2901 (N_2901,N_2896,N_2880);
xnor U2902 (N_2902,N_2851,N_2886);
and U2903 (N_2903,N_2856,N_2877);
nor U2904 (N_2904,N_2853,N_2835);
xnor U2905 (N_2905,N_2876,N_2800);
nor U2906 (N_2906,N_2803,N_2892);
or U2907 (N_2907,N_2887,N_2844);
and U2908 (N_2908,N_2820,N_2861);
nand U2909 (N_2909,N_2825,N_2866);
nor U2910 (N_2910,N_2859,N_2841);
nor U2911 (N_2911,N_2895,N_2806);
xor U2912 (N_2912,N_2874,N_2897);
or U2913 (N_2913,N_2873,N_2813);
or U2914 (N_2914,N_2831,N_2816);
nand U2915 (N_2915,N_2833,N_2815);
xnor U2916 (N_2916,N_2805,N_2890);
or U2917 (N_2917,N_2821,N_2827);
or U2918 (N_2918,N_2888,N_2898);
xor U2919 (N_2919,N_2801,N_2867);
and U2920 (N_2920,N_2839,N_2875);
nor U2921 (N_2921,N_2817,N_2894);
or U2922 (N_2922,N_2863,N_2872);
or U2923 (N_2923,N_2864,N_2845);
nor U2924 (N_2924,N_2865,N_2854);
or U2925 (N_2925,N_2878,N_2807);
xnor U2926 (N_2926,N_2836,N_2871);
xor U2927 (N_2927,N_2829,N_2840);
and U2928 (N_2928,N_2834,N_2869);
nand U2929 (N_2929,N_2852,N_2843);
nor U2930 (N_2930,N_2870,N_2838);
xor U2931 (N_2931,N_2828,N_2885);
nand U2932 (N_2932,N_2819,N_2824);
and U2933 (N_2933,N_2889,N_2893);
xnor U2934 (N_2934,N_2868,N_2809);
nand U2935 (N_2935,N_2830,N_2881);
or U2936 (N_2936,N_2826,N_2855);
nand U2937 (N_2937,N_2860,N_2883);
xor U2938 (N_2938,N_2822,N_2812);
xor U2939 (N_2939,N_2810,N_2823);
or U2940 (N_2940,N_2802,N_2884);
nand U2941 (N_2941,N_2832,N_2814);
and U2942 (N_2942,N_2879,N_2846);
nand U2943 (N_2943,N_2882,N_2858);
nand U2944 (N_2944,N_2847,N_2849);
xnor U2945 (N_2945,N_2862,N_2842);
or U2946 (N_2946,N_2804,N_2811);
or U2947 (N_2947,N_2891,N_2808);
and U2948 (N_2948,N_2899,N_2848);
and U2949 (N_2949,N_2837,N_2857);
and U2950 (N_2950,N_2809,N_2824);
xor U2951 (N_2951,N_2898,N_2806);
nor U2952 (N_2952,N_2866,N_2875);
nand U2953 (N_2953,N_2857,N_2886);
and U2954 (N_2954,N_2858,N_2878);
and U2955 (N_2955,N_2835,N_2839);
nor U2956 (N_2956,N_2839,N_2815);
nor U2957 (N_2957,N_2857,N_2826);
or U2958 (N_2958,N_2878,N_2822);
nor U2959 (N_2959,N_2854,N_2805);
xor U2960 (N_2960,N_2809,N_2892);
xnor U2961 (N_2961,N_2825,N_2823);
nor U2962 (N_2962,N_2876,N_2898);
xnor U2963 (N_2963,N_2855,N_2857);
or U2964 (N_2964,N_2807,N_2877);
nand U2965 (N_2965,N_2822,N_2815);
and U2966 (N_2966,N_2885,N_2853);
or U2967 (N_2967,N_2856,N_2805);
nor U2968 (N_2968,N_2821,N_2856);
and U2969 (N_2969,N_2878,N_2803);
nand U2970 (N_2970,N_2869,N_2810);
or U2971 (N_2971,N_2885,N_2854);
xor U2972 (N_2972,N_2854,N_2800);
nand U2973 (N_2973,N_2850,N_2803);
and U2974 (N_2974,N_2859,N_2846);
xnor U2975 (N_2975,N_2862,N_2894);
nand U2976 (N_2976,N_2862,N_2872);
and U2977 (N_2977,N_2875,N_2846);
nor U2978 (N_2978,N_2895,N_2884);
xnor U2979 (N_2979,N_2847,N_2810);
xor U2980 (N_2980,N_2864,N_2813);
nor U2981 (N_2981,N_2820,N_2805);
nor U2982 (N_2982,N_2817,N_2846);
nand U2983 (N_2983,N_2825,N_2815);
and U2984 (N_2984,N_2816,N_2806);
nor U2985 (N_2985,N_2805,N_2858);
xor U2986 (N_2986,N_2884,N_2853);
nand U2987 (N_2987,N_2810,N_2854);
xnor U2988 (N_2988,N_2888,N_2878);
or U2989 (N_2989,N_2832,N_2853);
and U2990 (N_2990,N_2819,N_2809);
and U2991 (N_2991,N_2817,N_2821);
nand U2992 (N_2992,N_2873,N_2899);
nand U2993 (N_2993,N_2876,N_2860);
or U2994 (N_2994,N_2826,N_2880);
or U2995 (N_2995,N_2840,N_2896);
nor U2996 (N_2996,N_2867,N_2890);
or U2997 (N_2997,N_2866,N_2889);
nor U2998 (N_2998,N_2864,N_2804);
or U2999 (N_2999,N_2886,N_2840);
xnor UO_0 (O_0,N_2992,N_2959);
nand UO_1 (O_1,N_2975,N_2955);
nand UO_2 (O_2,N_2964,N_2919);
or UO_3 (O_3,N_2935,N_2914);
nor UO_4 (O_4,N_2981,N_2968);
and UO_5 (O_5,N_2904,N_2913);
or UO_6 (O_6,N_2976,N_2940);
nand UO_7 (O_7,N_2910,N_2949);
and UO_8 (O_8,N_2998,N_2988);
nand UO_9 (O_9,N_2980,N_2957);
and UO_10 (O_10,N_2983,N_2995);
xor UO_11 (O_11,N_2990,N_2954);
nor UO_12 (O_12,N_2979,N_2965);
nor UO_13 (O_13,N_2911,N_2908);
nand UO_14 (O_14,N_2978,N_2984);
nor UO_15 (O_15,N_2929,N_2912);
nand UO_16 (O_16,N_2991,N_2977);
and UO_17 (O_17,N_2921,N_2952);
nand UO_18 (O_18,N_2969,N_2924);
xnor UO_19 (O_19,N_2994,N_2934);
nand UO_20 (O_20,N_2997,N_2945);
nand UO_21 (O_21,N_2928,N_2989);
xor UO_22 (O_22,N_2966,N_2986);
xnor UO_23 (O_23,N_2956,N_2901);
nor UO_24 (O_24,N_2905,N_2999);
and UO_25 (O_25,N_2951,N_2923);
and UO_26 (O_26,N_2932,N_2939);
xor UO_27 (O_27,N_2922,N_2920);
nor UO_28 (O_28,N_2925,N_2953);
nand UO_29 (O_29,N_2907,N_2915);
nor UO_30 (O_30,N_2947,N_2900);
and UO_31 (O_31,N_2960,N_2931);
and UO_32 (O_32,N_2906,N_2973);
and UO_33 (O_33,N_2970,N_2902);
nor UO_34 (O_34,N_2936,N_2903);
nor UO_35 (O_35,N_2962,N_2950);
nor UO_36 (O_36,N_2933,N_2944);
or UO_37 (O_37,N_2930,N_2948);
or UO_38 (O_38,N_2958,N_2961);
and UO_39 (O_39,N_2937,N_2926);
nor UO_40 (O_40,N_2943,N_2917);
or UO_41 (O_41,N_2918,N_2963);
nor UO_42 (O_42,N_2927,N_2916);
xor UO_43 (O_43,N_2941,N_2909);
or UO_44 (O_44,N_2942,N_2946);
or UO_45 (O_45,N_2971,N_2974);
nor UO_46 (O_46,N_2985,N_2996);
and UO_47 (O_47,N_2938,N_2987);
nor UO_48 (O_48,N_2993,N_2982);
nor UO_49 (O_49,N_2972,N_2967);
xor UO_50 (O_50,N_2922,N_2956);
xnor UO_51 (O_51,N_2922,N_2946);
nand UO_52 (O_52,N_2976,N_2980);
or UO_53 (O_53,N_2959,N_2972);
and UO_54 (O_54,N_2935,N_2915);
nor UO_55 (O_55,N_2900,N_2958);
or UO_56 (O_56,N_2996,N_2905);
and UO_57 (O_57,N_2937,N_2999);
or UO_58 (O_58,N_2951,N_2928);
xor UO_59 (O_59,N_2968,N_2921);
or UO_60 (O_60,N_2961,N_2923);
xor UO_61 (O_61,N_2963,N_2956);
nor UO_62 (O_62,N_2957,N_2947);
or UO_63 (O_63,N_2957,N_2963);
xor UO_64 (O_64,N_2948,N_2987);
or UO_65 (O_65,N_2913,N_2995);
and UO_66 (O_66,N_2914,N_2906);
xnor UO_67 (O_67,N_2959,N_2908);
nor UO_68 (O_68,N_2956,N_2975);
and UO_69 (O_69,N_2933,N_2977);
or UO_70 (O_70,N_2978,N_2946);
or UO_71 (O_71,N_2924,N_2994);
xor UO_72 (O_72,N_2905,N_2990);
and UO_73 (O_73,N_2982,N_2937);
or UO_74 (O_74,N_2949,N_2990);
nor UO_75 (O_75,N_2970,N_2951);
nor UO_76 (O_76,N_2952,N_2931);
nor UO_77 (O_77,N_2921,N_2944);
nor UO_78 (O_78,N_2921,N_2940);
nor UO_79 (O_79,N_2943,N_2951);
nor UO_80 (O_80,N_2979,N_2911);
and UO_81 (O_81,N_2919,N_2963);
nor UO_82 (O_82,N_2965,N_2966);
or UO_83 (O_83,N_2935,N_2902);
and UO_84 (O_84,N_2989,N_2945);
xnor UO_85 (O_85,N_2912,N_2923);
or UO_86 (O_86,N_2986,N_2923);
nand UO_87 (O_87,N_2941,N_2980);
nand UO_88 (O_88,N_2929,N_2943);
nand UO_89 (O_89,N_2974,N_2994);
and UO_90 (O_90,N_2923,N_2972);
nor UO_91 (O_91,N_2996,N_2909);
or UO_92 (O_92,N_2959,N_2935);
xor UO_93 (O_93,N_2960,N_2946);
and UO_94 (O_94,N_2906,N_2988);
and UO_95 (O_95,N_2968,N_2944);
xnor UO_96 (O_96,N_2924,N_2983);
nand UO_97 (O_97,N_2996,N_2932);
xor UO_98 (O_98,N_2927,N_2991);
and UO_99 (O_99,N_2976,N_2986);
nand UO_100 (O_100,N_2912,N_2917);
xor UO_101 (O_101,N_2955,N_2911);
and UO_102 (O_102,N_2995,N_2985);
nand UO_103 (O_103,N_2996,N_2902);
or UO_104 (O_104,N_2938,N_2994);
xor UO_105 (O_105,N_2985,N_2960);
and UO_106 (O_106,N_2989,N_2988);
nor UO_107 (O_107,N_2950,N_2926);
nand UO_108 (O_108,N_2911,N_2994);
xor UO_109 (O_109,N_2920,N_2983);
xor UO_110 (O_110,N_2969,N_2967);
or UO_111 (O_111,N_2971,N_2993);
xor UO_112 (O_112,N_2949,N_2978);
nor UO_113 (O_113,N_2920,N_2901);
or UO_114 (O_114,N_2991,N_2974);
nor UO_115 (O_115,N_2954,N_2918);
xnor UO_116 (O_116,N_2922,N_2910);
and UO_117 (O_117,N_2957,N_2976);
and UO_118 (O_118,N_2907,N_2938);
nor UO_119 (O_119,N_2909,N_2994);
or UO_120 (O_120,N_2970,N_2969);
nand UO_121 (O_121,N_2970,N_2931);
nand UO_122 (O_122,N_2992,N_2901);
or UO_123 (O_123,N_2965,N_2941);
nand UO_124 (O_124,N_2922,N_2915);
xor UO_125 (O_125,N_2995,N_2924);
and UO_126 (O_126,N_2918,N_2926);
and UO_127 (O_127,N_2966,N_2967);
xor UO_128 (O_128,N_2907,N_2936);
nor UO_129 (O_129,N_2997,N_2927);
or UO_130 (O_130,N_2941,N_2986);
nor UO_131 (O_131,N_2934,N_2933);
nor UO_132 (O_132,N_2943,N_2990);
or UO_133 (O_133,N_2990,N_2911);
or UO_134 (O_134,N_2944,N_2966);
nand UO_135 (O_135,N_2931,N_2916);
and UO_136 (O_136,N_2967,N_2991);
and UO_137 (O_137,N_2967,N_2962);
nor UO_138 (O_138,N_2906,N_2972);
nand UO_139 (O_139,N_2949,N_2938);
nand UO_140 (O_140,N_2958,N_2915);
nor UO_141 (O_141,N_2997,N_2998);
nand UO_142 (O_142,N_2916,N_2992);
xor UO_143 (O_143,N_2919,N_2947);
and UO_144 (O_144,N_2994,N_2987);
or UO_145 (O_145,N_2980,N_2989);
and UO_146 (O_146,N_2906,N_2951);
xor UO_147 (O_147,N_2991,N_2965);
nand UO_148 (O_148,N_2948,N_2906);
and UO_149 (O_149,N_2911,N_2924);
nand UO_150 (O_150,N_2978,N_2957);
nor UO_151 (O_151,N_2935,N_2934);
or UO_152 (O_152,N_2992,N_2943);
and UO_153 (O_153,N_2911,N_2961);
or UO_154 (O_154,N_2944,N_2995);
xnor UO_155 (O_155,N_2921,N_2926);
nor UO_156 (O_156,N_2917,N_2976);
nor UO_157 (O_157,N_2983,N_2992);
nor UO_158 (O_158,N_2923,N_2905);
nand UO_159 (O_159,N_2924,N_2964);
nor UO_160 (O_160,N_2944,N_2973);
nor UO_161 (O_161,N_2970,N_2948);
and UO_162 (O_162,N_2950,N_2957);
or UO_163 (O_163,N_2957,N_2953);
nor UO_164 (O_164,N_2962,N_2986);
xor UO_165 (O_165,N_2940,N_2914);
xor UO_166 (O_166,N_2948,N_2911);
nand UO_167 (O_167,N_2988,N_2929);
nor UO_168 (O_168,N_2964,N_2963);
nand UO_169 (O_169,N_2953,N_2907);
nor UO_170 (O_170,N_2915,N_2992);
nand UO_171 (O_171,N_2913,N_2991);
nor UO_172 (O_172,N_2954,N_2991);
and UO_173 (O_173,N_2904,N_2971);
nand UO_174 (O_174,N_2945,N_2948);
nand UO_175 (O_175,N_2994,N_2981);
xor UO_176 (O_176,N_2981,N_2911);
or UO_177 (O_177,N_2921,N_2993);
nor UO_178 (O_178,N_2931,N_2927);
nor UO_179 (O_179,N_2909,N_2999);
nand UO_180 (O_180,N_2909,N_2961);
or UO_181 (O_181,N_2934,N_2982);
and UO_182 (O_182,N_2907,N_2980);
or UO_183 (O_183,N_2961,N_2993);
xor UO_184 (O_184,N_2959,N_2948);
nand UO_185 (O_185,N_2958,N_2963);
and UO_186 (O_186,N_2975,N_2977);
xnor UO_187 (O_187,N_2901,N_2981);
or UO_188 (O_188,N_2931,N_2995);
and UO_189 (O_189,N_2992,N_2977);
nor UO_190 (O_190,N_2938,N_2930);
or UO_191 (O_191,N_2936,N_2923);
xnor UO_192 (O_192,N_2903,N_2923);
or UO_193 (O_193,N_2917,N_2989);
xnor UO_194 (O_194,N_2973,N_2908);
nand UO_195 (O_195,N_2998,N_2948);
xnor UO_196 (O_196,N_2960,N_2936);
or UO_197 (O_197,N_2982,N_2954);
nor UO_198 (O_198,N_2925,N_2907);
xor UO_199 (O_199,N_2943,N_2994);
nand UO_200 (O_200,N_2941,N_2935);
nor UO_201 (O_201,N_2922,N_2900);
nor UO_202 (O_202,N_2922,N_2919);
or UO_203 (O_203,N_2952,N_2959);
nor UO_204 (O_204,N_2990,N_2931);
nand UO_205 (O_205,N_2995,N_2908);
nor UO_206 (O_206,N_2963,N_2916);
nor UO_207 (O_207,N_2953,N_2954);
and UO_208 (O_208,N_2961,N_2926);
and UO_209 (O_209,N_2914,N_2953);
nand UO_210 (O_210,N_2903,N_2940);
nor UO_211 (O_211,N_2956,N_2989);
or UO_212 (O_212,N_2902,N_2985);
xnor UO_213 (O_213,N_2988,N_2951);
nor UO_214 (O_214,N_2937,N_2940);
xnor UO_215 (O_215,N_2977,N_2990);
nand UO_216 (O_216,N_2946,N_2902);
nor UO_217 (O_217,N_2950,N_2984);
nor UO_218 (O_218,N_2976,N_2973);
nand UO_219 (O_219,N_2984,N_2917);
nand UO_220 (O_220,N_2996,N_2961);
nand UO_221 (O_221,N_2976,N_2990);
xor UO_222 (O_222,N_2942,N_2972);
or UO_223 (O_223,N_2934,N_2917);
and UO_224 (O_224,N_2957,N_2964);
nand UO_225 (O_225,N_2976,N_2933);
or UO_226 (O_226,N_2910,N_2920);
nand UO_227 (O_227,N_2909,N_2911);
nor UO_228 (O_228,N_2925,N_2979);
and UO_229 (O_229,N_2934,N_2993);
xnor UO_230 (O_230,N_2980,N_2925);
nand UO_231 (O_231,N_2933,N_2930);
or UO_232 (O_232,N_2908,N_2954);
xor UO_233 (O_233,N_2918,N_2919);
and UO_234 (O_234,N_2916,N_2988);
or UO_235 (O_235,N_2964,N_2978);
nand UO_236 (O_236,N_2930,N_2980);
xnor UO_237 (O_237,N_2953,N_2923);
xnor UO_238 (O_238,N_2979,N_2912);
nor UO_239 (O_239,N_2994,N_2955);
xnor UO_240 (O_240,N_2957,N_2930);
nor UO_241 (O_241,N_2927,N_2960);
nor UO_242 (O_242,N_2984,N_2945);
nor UO_243 (O_243,N_2949,N_2904);
and UO_244 (O_244,N_2940,N_2944);
xor UO_245 (O_245,N_2980,N_2948);
xnor UO_246 (O_246,N_2945,N_2912);
or UO_247 (O_247,N_2955,N_2922);
xor UO_248 (O_248,N_2968,N_2967);
and UO_249 (O_249,N_2982,N_2968);
xnor UO_250 (O_250,N_2943,N_2987);
or UO_251 (O_251,N_2940,N_2934);
nand UO_252 (O_252,N_2980,N_2995);
nor UO_253 (O_253,N_2902,N_2977);
and UO_254 (O_254,N_2963,N_2945);
nor UO_255 (O_255,N_2948,N_2946);
and UO_256 (O_256,N_2960,N_2967);
or UO_257 (O_257,N_2964,N_2988);
and UO_258 (O_258,N_2945,N_2904);
and UO_259 (O_259,N_2984,N_2957);
and UO_260 (O_260,N_2995,N_2916);
nand UO_261 (O_261,N_2956,N_2983);
or UO_262 (O_262,N_2954,N_2970);
nor UO_263 (O_263,N_2906,N_2954);
nor UO_264 (O_264,N_2949,N_2927);
or UO_265 (O_265,N_2933,N_2915);
and UO_266 (O_266,N_2963,N_2903);
xor UO_267 (O_267,N_2966,N_2984);
or UO_268 (O_268,N_2948,N_2922);
and UO_269 (O_269,N_2922,N_2913);
or UO_270 (O_270,N_2955,N_2917);
nor UO_271 (O_271,N_2989,N_2923);
and UO_272 (O_272,N_2965,N_2918);
or UO_273 (O_273,N_2906,N_2999);
nand UO_274 (O_274,N_2972,N_2978);
nor UO_275 (O_275,N_2914,N_2909);
nand UO_276 (O_276,N_2932,N_2938);
nor UO_277 (O_277,N_2994,N_2946);
nand UO_278 (O_278,N_2930,N_2958);
or UO_279 (O_279,N_2956,N_2940);
or UO_280 (O_280,N_2946,N_2914);
nand UO_281 (O_281,N_2968,N_2960);
nand UO_282 (O_282,N_2951,N_2932);
xnor UO_283 (O_283,N_2985,N_2998);
and UO_284 (O_284,N_2959,N_2961);
nand UO_285 (O_285,N_2936,N_2943);
and UO_286 (O_286,N_2989,N_2931);
xor UO_287 (O_287,N_2993,N_2989);
and UO_288 (O_288,N_2947,N_2980);
nor UO_289 (O_289,N_2910,N_2986);
and UO_290 (O_290,N_2966,N_2924);
or UO_291 (O_291,N_2947,N_2970);
nand UO_292 (O_292,N_2994,N_2932);
nand UO_293 (O_293,N_2918,N_2941);
or UO_294 (O_294,N_2977,N_2956);
nor UO_295 (O_295,N_2932,N_2902);
nor UO_296 (O_296,N_2991,N_2988);
nor UO_297 (O_297,N_2921,N_2917);
and UO_298 (O_298,N_2989,N_2908);
or UO_299 (O_299,N_2921,N_2958);
or UO_300 (O_300,N_2936,N_2955);
or UO_301 (O_301,N_2982,N_2996);
or UO_302 (O_302,N_2958,N_2919);
nand UO_303 (O_303,N_2977,N_2921);
xnor UO_304 (O_304,N_2971,N_2944);
or UO_305 (O_305,N_2925,N_2995);
and UO_306 (O_306,N_2905,N_2973);
xnor UO_307 (O_307,N_2956,N_2919);
xor UO_308 (O_308,N_2976,N_2979);
or UO_309 (O_309,N_2928,N_2923);
nand UO_310 (O_310,N_2956,N_2942);
xor UO_311 (O_311,N_2901,N_2998);
and UO_312 (O_312,N_2910,N_2916);
nor UO_313 (O_313,N_2983,N_2964);
nand UO_314 (O_314,N_2924,N_2998);
and UO_315 (O_315,N_2972,N_2937);
nand UO_316 (O_316,N_2986,N_2913);
nor UO_317 (O_317,N_2906,N_2961);
xor UO_318 (O_318,N_2915,N_2986);
and UO_319 (O_319,N_2911,N_2951);
xor UO_320 (O_320,N_2917,N_2968);
nand UO_321 (O_321,N_2949,N_2964);
nand UO_322 (O_322,N_2926,N_2923);
and UO_323 (O_323,N_2977,N_2903);
nor UO_324 (O_324,N_2999,N_2930);
xor UO_325 (O_325,N_2932,N_2948);
xor UO_326 (O_326,N_2992,N_2919);
and UO_327 (O_327,N_2977,N_2945);
or UO_328 (O_328,N_2962,N_2947);
nand UO_329 (O_329,N_2942,N_2959);
xor UO_330 (O_330,N_2913,N_2925);
nor UO_331 (O_331,N_2958,N_2927);
nand UO_332 (O_332,N_2955,N_2933);
xnor UO_333 (O_333,N_2991,N_2958);
xor UO_334 (O_334,N_2971,N_2990);
or UO_335 (O_335,N_2981,N_2967);
or UO_336 (O_336,N_2964,N_2922);
and UO_337 (O_337,N_2998,N_2923);
xor UO_338 (O_338,N_2914,N_2911);
xor UO_339 (O_339,N_2976,N_2901);
or UO_340 (O_340,N_2994,N_2957);
xnor UO_341 (O_341,N_2971,N_2948);
nand UO_342 (O_342,N_2902,N_2939);
nor UO_343 (O_343,N_2967,N_2925);
and UO_344 (O_344,N_2981,N_2943);
nor UO_345 (O_345,N_2976,N_2932);
nor UO_346 (O_346,N_2907,N_2993);
and UO_347 (O_347,N_2910,N_2903);
or UO_348 (O_348,N_2926,N_2993);
xor UO_349 (O_349,N_2994,N_2914);
xor UO_350 (O_350,N_2990,N_2956);
nand UO_351 (O_351,N_2982,N_2930);
and UO_352 (O_352,N_2935,N_2909);
and UO_353 (O_353,N_2964,N_2936);
and UO_354 (O_354,N_2912,N_2913);
nor UO_355 (O_355,N_2952,N_2998);
or UO_356 (O_356,N_2949,N_2958);
and UO_357 (O_357,N_2932,N_2992);
or UO_358 (O_358,N_2942,N_2951);
or UO_359 (O_359,N_2961,N_2991);
nor UO_360 (O_360,N_2994,N_2915);
nand UO_361 (O_361,N_2934,N_2931);
xor UO_362 (O_362,N_2940,N_2906);
nor UO_363 (O_363,N_2967,N_2988);
or UO_364 (O_364,N_2930,N_2909);
or UO_365 (O_365,N_2958,N_2998);
nor UO_366 (O_366,N_2971,N_2969);
xnor UO_367 (O_367,N_2912,N_2973);
or UO_368 (O_368,N_2961,N_2914);
xnor UO_369 (O_369,N_2917,N_2964);
nor UO_370 (O_370,N_2916,N_2959);
and UO_371 (O_371,N_2929,N_2999);
or UO_372 (O_372,N_2947,N_2933);
nor UO_373 (O_373,N_2976,N_2960);
xnor UO_374 (O_374,N_2907,N_2987);
and UO_375 (O_375,N_2978,N_2968);
nor UO_376 (O_376,N_2919,N_2959);
and UO_377 (O_377,N_2983,N_2985);
and UO_378 (O_378,N_2947,N_2987);
or UO_379 (O_379,N_2915,N_2947);
nand UO_380 (O_380,N_2922,N_2995);
and UO_381 (O_381,N_2987,N_2964);
and UO_382 (O_382,N_2925,N_2963);
or UO_383 (O_383,N_2928,N_2996);
or UO_384 (O_384,N_2963,N_2927);
or UO_385 (O_385,N_2973,N_2982);
nand UO_386 (O_386,N_2921,N_2980);
and UO_387 (O_387,N_2976,N_2963);
nor UO_388 (O_388,N_2917,N_2949);
nor UO_389 (O_389,N_2920,N_2985);
and UO_390 (O_390,N_2973,N_2986);
nor UO_391 (O_391,N_2994,N_2908);
xor UO_392 (O_392,N_2984,N_2942);
or UO_393 (O_393,N_2979,N_2927);
nand UO_394 (O_394,N_2967,N_2978);
or UO_395 (O_395,N_2912,N_2978);
and UO_396 (O_396,N_2927,N_2983);
nand UO_397 (O_397,N_2960,N_2996);
and UO_398 (O_398,N_2994,N_2939);
or UO_399 (O_399,N_2913,N_2900);
or UO_400 (O_400,N_2925,N_2986);
or UO_401 (O_401,N_2938,N_2952);
xnor UO_402 (O_402,N_2985,N_2999);
nor UO_403 (O_403,N_2929,N_2939);
nor UO_404 (O_404,N_2959,N_2907);
nor UO_405 (O_405,N_2947,N_2983);
and UO_406 (O_406,N_2995,N_2982);
xnor UO_407 (O_407,N_2906,N_2958);
and UO_408 (O_408,N_2999,N_2919);
and UO_409 (O_409,N_2969,N_2947);
xnor UO_410 (O_410,N_2962,N_2980);
xnor UO_411 (O_411,N_2985,N_2931);
nand UO_412 (O_412,N_2905,N_2935);
nand UO_413 (O_413,N_2991,N_2959);
xnor UO_414 (O_414,N_2948,N_2964);
xor UO_415 (O_415,N_2941,N_2930);
and UO_416 (O_416,N_2962,N_2917);
xor UO_417 (O_417,N_2969,N_2932);
nand UO_418 (O_418,N_2941,N_2922);
nor UO_419 (O_419,N_2924,N_2937);
xor UO_420 (O_420,N_2947,N_2916);
nor UO_421 (O_421,N_2908,N_2992);
nand UO_422 (O_422,N_2916,N_2914);
and UO_423 (O_423,N_2909,N_2937);
or UO_424 (O_424,N_2950,N_2940);
nand UO_425 (O_425,N_2959,N_2999);
xor UO_426 (O_426,N_2937,N_2976);
nand UO_427 (O_427,N_2909,N_2926);
xnor UO_428 (O_428,N_2999,N_2920);
nor UO_429 (O_429,N_2992,N_2946);
or UO_430 (O_430,N_2942,N_2965);
xor UO_431 (O_431,N_2950,N_2959);
nor UO_432 (O_432,N_2949,N_2940);
or UO_433 (O_433,N_2928,N_2957);
and UO_434 (O_434,N_2903,N_2951);
xnor UO_435 (O_435,N_2947,N_2951);
or UO_436 (O_436,N_2901,N_2928);
xor UO_437 (O_437,N_2920,N_2956);
and UO_438 (O_438,N_2986,N_2965);
and UO_439 (O_439,N_2945,N_2972);
nand UO_440 (O_440,N_2972,N_2948);
nand UO_441 (O_441,N_2934,N_2948);
or UO_442 (O_442,N_2967,N_2953);
nor UO_443 (O_443,N_2986,N_2994);
xnor UO_444 (O_444,N_2983,N_2904);
or UO_445 (O_445,N_2953,N_2939);
nor UO_446 (O_446,N_2902,N_2922);
or UO_447 (O_447,N_2903,N_2965);
nor UO_448 (O_448,N_2949,N_2970);
xor UO_449 (O_449,N_2954,N_2902);
or UO_450 (O_450,N_2999,N_2949);
nor UO_451 (O_451,N_2938,N_2970);
nand UO_452 (O_452,N_2943,N_2942);
xnor UO_453 (O_453,N_2928,N_2929);
nor UO_454 (O_454,N_2967,N_2915);
xnor UO_455 (O_455,N_2979,N_2961);
and UO_456 (O_456,N_2908,N_2943);
nand UO_457 (O_457,N_2968,N_2908);
and UO_458 (O_458,N_2943,N_2980);
nor UO_459 (O_459,N_2949,N_2922);
and UO_460 (O_460,N_2978,N_2954);
nand UO_461 (O_461,N_2994,N_2982);
nor UO_462 (O_462,N_2921,N_2932);
or UO_463 (O_463,N_2915,N_2944);
xor UO_464 (O_464,N_2920,N_2931);
xnor UO_465 (O_465,N_2941,N_2981);
xor UO_466 (O_466,N_2918,N_2958);
and UO_467 (O_467,N_2960,N_2993);
xnor UO_468 (O_468,N_2946,N_2917);
nand UO_469 (O_469,N_2928,N_2970);
nand UO_470 (O_470,N_2955,N_2960);
nor UO_471 (O_471,N_2994,N_2963);
xnor UO_472 (O_472,N_2966,N_2973);
and UO_473 (O_473,N_2986,N_2920);
xor UO_474 (O_474,N_2933,N_2935);
or UO_475 (O_475,N_2916,N_2969);
nor UO_476 (O_476,N_2974,N_2917);
and UO_477 (O_477,N_2942,N_2988);
xnor UO_478 (O_478,N_2965,N_2972);
and UO_479 (O_479,N_2928,N_2959);
and UO_480 (O_480,N_2999,N_2902);
nor UO_481 (O_481,N_2977,N_2993);
nor UO_482 (O_482,N_2908,N_2913);
xor UO_483 (O_483,N_2940,N_2912);
nor UO_484 (O_484,N_2953,N_2904);
nand UO_485 (O_485,N_2957,N_2917);
and UO_486 (O_486,N_2915,N_2969);
xor UO_487 (O_487,N_2936,N_2929);
xnor UO_488 (O_488,N_2992,N_2993);
xnor UO_489 (O_489,N_2994,N_2942);
nor UO_490 (O_490,N_2931,N_2986);
xor UO_491 (O_491,N_2936,N_2918);
or UO_492 (O_492,N_2937,N_2970);
and UO_493 (O_493,N_2929,N_2987);
or UO_494 (O_494,N_2941,N_2931);
and UO_495 (O_495,N_2939,N_2937);
nor UO_496 (O_496,N_2910,N_2963);
nand UO_497 (O_497,N_2913,N_2967);
and UO_498 (O_498,N_2992,N_2928);
nand UO_499 (O_499,N_2965,N_2951);
endmodule